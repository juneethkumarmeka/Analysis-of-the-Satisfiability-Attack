module basic_1500_15000_2000_5_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
xnor U0 (N_0,In_409,In_1365);
nor U1 (N_1,In_251,In_576);
nand U2 (N_2,In_694,In_296);
xnor U3 (N_3,In_242,In_1180);
or U4 (N_4,In_984,In_515);
nor U5 (N_5,In_56,In_1078);
nand U6 (N_6,In_110,In_1252);
and U7 (N_7,In_434,In_592);
nand U8 (N_8,In_224,In_819);
nor U9 (N_9,In_315,In_64);
nor U10 (N_10,In_747,In_989);
nor U11 (N_11,In_259,In_1087);
nor U12 (N_12,In_1002,In_857);
xor U13 (N_13,In_377,In_640);
nor U14 (N_14,In_1219,In_117);
nand U15 (N_15,In_1428,In_379);
nand U16 (N_16,In_286,In_436);
nor U17 (N_17,In_650,In_712);
or U18 (N_18,In_1028,In_1303);
nand U19 (N_19,In_1275,In_417);
or U20 (N_20,In_871,In_624);
nand U21 (N_21,In_44,In_481);
nor U22 (N_22,In_388,In_1030);
nand U23 (N_23,In_865,In_328);
nor U24 (N_24,In_872,In_1478);
nand U25 (N_25,In_189,In_429);
nor U26 (N_26,In_266,In_510);
nand U27 (N_27,In_825,In_460);
nor U28 (N_28,In_1240,In_1264);
nand U29 (N_29,In_1396,In_759);
nor U30 (N_30,In_758,In_1339);
and U31 (N_31,In_1268,In_913);
xor U32 (N_32,In_413,In_1415);
xor U33 (N_33,In_98,In_212);
or U34 (N_34,In_4,In_1439);
nor U35 (N_35,In_1257,In_391);
and U36 (N_36,In_835,In_967);
xnor U37 (N_37,In_34,In_214);
and U38 (N_38,In_1077,In_578);
nor U39 (N_39,In_794,In_172);
nor U40 (N_40,In_288,In_868);
nor U41 (N_41,In_438,In_154);
nand U42 (N_42,In_79,In_962);
and U43 (N_43,In_180,In_127);
nand U44 (N_44,In_580,In_244);
and U45 (N_45,In_749,In_211);
and U46 (N_46,In_325,In_561);
and U47 (N_47,In_1473,In_1476);
nor U48 (N_48,In_1097,In_699);
nor U49 (N_49,In_1061,In_729);
or U50 (N_50,In_1270,In_599);
xnor U51 (N_51,In_126,In_866);
or U52 (N_52,In_1470,In_1004);
nor U53 (N_53,In_430,In_904);
xor U54 (N_54,In_1132,In_139);
nor U55 (N_55,In_1261,In_1050);
nor U56 (N_56,In_682,In_703);
and U57 (N_57,In_1133,In_1360);
or U58 (N_58,In_1461,In_734);
nor U59 (N_59,In_457,In_621);
or U60 (N_60,In_1272,In_517);
nor U61 (N_61,In_1242,In_641);
nand U62 (N_62,In_1115,In_671);
nand U63 (N_63,In_1361,In_870);
nand U64 (N_64,In_635,In_18);
xor U65 (N_65,In_804,In_1335);
and U66 (N_66,In_46,In_1094);
or U67 (N_67,In_750,In_90);
or U68 (N_68,In_771,In_947);
nor U69 (N_69,In_797,In_411);
or U70 (N_70,In_550,In_1312);
nor U71 (N_71,In_387,In_1244);
nand U72 (N_72,In_191,In_1232);
nor U73 (N_73,In_1391,In_277);
or U74 (N_74,In_1246,In_676);
and U75 (N_75,In_28,In_1041);
and U76 (N_76,In_831,In_558);
and U77 (N_77,In_176,In_385);
or U78 (N_78,In_1285,In_1025);
and U79 (N_79,In_92,In_594);
and U80 (N_80,In_744,In_1202);
nor U81 (N_81,In_1214,In_1157);
nor U82 (N_82,In_13,In_291);
or U83 (N_83,In_169,In_338);
nand U84 (N_84,In_602,In_99);
and U85 (N_85,In_1072,In_1297);
nor U86 (N_86,In_596,In_336);
nand U87 (N_87,In_678,In_41);
nor U88 (N_88,In_944,In_1300);
or U89 (N_89,In_193,In_1422);
nor U90 (N_90,In_454,In_1369);
or U91 (N_91,In_71,In_809);
nor U92 (N_92,In_1457,In_1340);
and U93 (N_93,In_1353,In_252);
xor U94 (N_94,In_497,In_76);
nor U95 (N_95,In_1225,In_516);
nor U96 (N_96,In_914,In_321);
nand U97 (N_97,In_665,In_1372);
and U98 (N_98,In_318,In_1319);
nand U99 (N_99,In_226,In_828);
xor U100 (N_100,In_1450,In_726);
nand U101 (N_101,In_492,In_1059);
and U102 (N_102,In_538,In_358);
nor U103 (N_103,In_269,In_1175);
or U104 (N_104,In_610,In_1455);
nor U105 (N_105,In_299,In_293);
and U106 (N_106,In_312,In_1018);
nand U107 (N_107,In_930,In_1222);
nor U108 (N_108,In_1306,In_1003);
nand U109 (N_109,In_415,In_767);
nor U110 (N_110,In_1276,In_82);
and U111 (N_111,In_752,In_1484);
or U112 (N_112,In_68,In_1235);
nor U113 (N_113,In_1141,In_929);
nand U114 (N_114,In_1314,In_1490);
or U115 (N_115,In_710,In_822);
and U116 (N_116,In_850,In_183);
nand U117 (N_117,In_170,In_143);
or U118 (N_118,In_1152,In_1421);
or U119 (N_119,In_1084,In_875);
nor U120 (N_120,In_485,In_570);
or U121 (N_121,In_642,In_271);
or U122 (N_122,In_604,In_416);
xor U123 (N_123,In_258,In_581);
and U124 (N_124,In_966,In_1237);
xnor U125 (N_125,In_833,In_1071);
nor U126 (N_126,In_628,In_1343);
nor U127 (N_127,In_996,In_689);
nand U128 (N_128,In_499,In_958);
and U129 (N_129,In_792,In_419);
nand U130 (N_130,In_826,In_348);
nand U131 (N_131,In_491,In_856);
nor U132 (N_132,In_213,In_209);
or U133 (N_133,In_884,In_339);
xor U134 (N_134,In_302,In_294);
nand U135 (N_135,In_1298,In_637);
nor U136 (N_136,In_1221,In_607);
nor U137 (N_137,In_74,In_1048);
xor U138 (N_138,In_1196,In_48);
and U139 (N_139,In_651,In_1350);
xnor U140 (N_140,In_1345,In_761);
or U141 (N_141,In_1435,In_129);
or U142 (N_142,In_1393,In_52);
or U143 (N_143,In_1169,In_199);
xor U144 (N_144,In_796,In_840);
or U145 (N_145,In_498,In_472);
nor U146 (N_146,In_1096,In_204);
and U147 (N_147,In_1438,In_124);
and U148 (N_148,In_1430,In_1248);
xor U149 (N_149,In_688,In_1354);
or U150 (N_150,In_784,In_210);
nor U151 (N_151,In_1099,In_330);
nor U152 (N_152,In_1493,In_471);
nor U153 (N_153,In_32,In_575);
nand U154 (N_154,In_440,In_462);
nand U155 (N_155,In_1182,In_839);
nor U156 (N_156,In_687,In_990);
nor U157 (N_157,In_1333,In_1104);
or U158 (N_158,In_335,In_344);
nor U159 (N_159,In_185,In_902);
or U160 (N_160,In_731,In_69);
or U161 (N_161,In_85,In_1281);
or U162 (N_162,In_933,In_45);
nand U163 (N_163,In_182,In_1427);
and U164 (N_164,In_1256,In_1015);
nand U165 (N_165,In_428,In_443);
xnor U166 (N_166,In_322,In_686);
nor U167 (N_167,In_995,In_1321);
nor U168 (N_168,In_733,In_577);
xor U169 (N_169,In_369,In_541);
nor U170 (N_170,In_220,In_1486);
nand U171 (N_171,In_77,In_632);
nand U172 (N_172,In_1447,In_205);
nor U173 (N_173,In_166,In_368);
nor U174 (N_174,In_431,In_201);
xor U175 (N_175,In_149,In_389);
nor U176 (N_176,In_347,In_463);
and U177 (N_177,In_292,In_873);
and U178 (N_178,In_614,In_847);
or U179 (N_179,In_1446,In_1459);
or U180 (N_180,In_384,In_700);
and U181 (N_181,In_598,In_151);
xnor U182 (N_182,In_623,In_134);
nor U183 (N_183,In_1352,In_745);
and U184 (N_184,In_1024,In_101);
and U185 (N_185,In_874,In_1198);
and U186 (N_186,In_692,In_1379);
nand U187 (N_187,In_1146,In_309);
or U188 (N_188,In_760,In_1082);
and U189 (N_189,In_1075,In_1398);
xor U190 (N_190,In_821,In_346);
xnor U191 (N_191,In_367,In_1187);
and U192 (N_192,In_298,In_636);
nor U193 (N_193,In_529,In_1035);
nor U194 (N_194,In_290,In_1249);
nand U195 (N_195,In_1234,In_107);
nand U196 (N_196,In_780,In_1452);
nand U197 (N_197,In_403,In_737);
xnor U198 (N_198,In_1496,In_1332);
nand U199 (N_199,In_748,In_43);
nor U200 (N_200,In_1009,In_969);
or U201 (N_201,In_1480,In_1184);
nor U202 (N_202,In_114,In_1109);
or U203 (N_203,In_219,In_53);
nand U204 (N_204,In_333,In_222);
nor U205 (N_205,In_1358,In_102);
and U206 (N_206,In_1411,In_863);
nand U207 (N_207,In_1116,In_352);
nor U208 (N_208,In_588,In_736);
nand U209 (N_209,In_265,In_707);
xor U210 (N_210,In_412,In_135);
nand U211 (N_211,In_1117,In_803);
nor U212 (N_212,In_960,In_532);
nand U213 (N_213,In_1051,In_1029);
and U214 (N_214,In_1086,In_1218);
or U215 (N_215,In_63,In_546);
nor U216 (N_216,In_727,In_281);
nand U217 (N_217,In_397,In_530);
or U218 (N_218,In_1395,In_1014);
or U219 (N_219,In_609,In_569);
nor U220 (N_220,In_1211,In_533);
nor U221 (N_221,In_1049,In_10);
nand U222 (N_222,In_1194,In_1057);
nand U223 (N_223,In_983,In_1027);
and U224 (N_224,In_42,In_1047);
nand U225 (N_225,In_168,In_1236);
and U226 (N_226,In_317,In_525);
or U227 (N_227,In_879,In_1073);
or U228 (N_228,In_1482,In_1227);
and U229 (N_229,In_477,In_61);
and U230 (N_230,In_545,In_590);
nand U231 (N_231,In_240,In_218);
and U232 (N_232,In_813,In_920);
nand U233 (N_233,In_754,In_223);
or U234 (N_234,In_993,In_1195);
nand U235 (N_235,In_938,In_1188);
and U236 (N_236,In_320,In_1463);
or U237 (N_237,In_319,In_1323);
nor U238 (N_238,In_661,In_843);
nand U239 (N_239,In_978,In_480);
and U240 (N_240,In_741,In_583);
and U241 (N_241,In_1036,In_1420);
nor U242 (N_242,In_111,In_1220);
nor U243 (N_243,In_130,In_732);
or U244 (N_244,In_1216,In_1380);
nand U245 (N_245,In_1193,In_364);
or U246 (N_246,In_939,In_356);
and U247 (N_247,In_494,In_946);
or U248 (N_248,In_29,In_653);
or U249 (N_249,In_1417,In_763);
nand U250 (N_250,In_233,In_1449);
xnor U251 (N_251,In_442,In_394);
nor U252 (N_252,In_297,In_772);
xor U253 (N_253,In_793,In_612);
nor U254 (N_254,In_1044,In_420);
and U255 (N_255,In_560,In_746);
xor U256 (N_256,In_730,In_489);
or U257 (N_257,In_125,In_836);
nand U258 (N_258,In_961,In_1147);
xnor U259 (N_259,In_70,In_57);
nand U260 (N_260,In_502,In_1255);
nand U261 (N_261,In_1007,In_192);
nor U262 (N_262,In_1171,In_559);
or U263 (N_263,In_1055,In_805);
and U264 (N_264,In_812,In_261);
and U265 (N_265,In_1183,In_698);
nand U266 (N_266,In_706,In_359);
nor U267 (N_267,In_1226,In_1357);
or U268 (N_268,In_1081,In_1381);
nor U269 (N_269,In_743,In_777);
xnor U270 (N_270,In_683,In_1181);
or U271 (N_271,In_1224,In_1178);
nor U272 (N_272,In_907,In_310);
nor U273 (N_273,In_0,In_1042);
and U274 (N_274,In_1349,In_662);
nor U275 (N_275,In_885,In_400);
and U276 (N_276,In_165,In_217);
xnor U277 (N_277,In_1093,In_848);
nand U278 (N_278,In_1383,In_1129);
and U279 (N_279,In_1467,In_402);
nand U280 (N_280,In_1108,In_1172);
or U281 (N_281,In_1331,In_1245);
nor U282 (N_282,In_235,In_1229);
or U283 (N_283,In_991,In_116);
nor U284 (N_284,In_672,In_1305);
and U285 (N_285,In_324,In_898);
or U286 (N_286,In_307,In_791);
or U287 (N_287,In_1017,In_1160);
nand U288 (N_288,In_751,In_345);
xor U289 (N_289,In_514,In_1023);
or U290 (N_290,In_618,In_1233);
or U291 (N_291,In_361,In_790);
or U292 (N_292,In_87,In_631);
nor U293 (N_293,In_877,In_216);
or U294 (N_294,In_264,In_1138);
xnor U295 (N_295,In_501,In_660);
nor U296 (N_296,In_509,In_1091);
xnor U297 (N_297,In_256,In_519);
nor U298 (N_298,In_1090,In_584);
and U299 (N_299,In_283,In_1013);
and U300 (N_300,In_1403,In_25);
or U301 (N_301,In_329,In_1282);
or U302 (N_302,In_1389,In_1151);
xor U303 (N_303,In_1342,In_1161);
or U304 (N_304,In_770,In_1274);
nand U305 (N_305,In_490,In_171);
and U306 (N_306,In_1377,In_928);
nand U307 (N_307,In_753,In_518);
and U308 (N_308,In_287,In_764);
and U309 (N_309,In_1006,In_1148);
or U310 (N_310,In_1310,In_1067);
nand U311 (N_311,In_625,In_1280);
or U312 (N_312,In_1070,In_466);
xor U313 (N_313,In_72,In_888);
and U314 (N_314,In_1021,In_274);
or U315 (N_315,In_781,In_215);
nor U316 (N_316,In_253,In_629);
nor U317 (N_317,In_1477,In_1469);
or U318 (N_318,In_1414,In_128);
xnor U319 (N_319,In_940,In_1454);
xor U320 (N_320,In_1238,In_1304);
and U321 (N_321,In_375,In_556);
nor U322 (N_322,In_1192,In_1176);
nor U323 (N_323,In_1165,In_854);
nand U324 (N_324,In_395,In_202);
nand U325 (N_325,In_782,In_1499);
nand U326 (N_326,In_279,In_1155);
nor U327 (N_327,In_691,In_951);
and U328 (N_328,In_713,In_236);
and U329 (N_329,In_316,In_198);
or U330 (N_330,In_1026,In_399);
nor U331 (N_331,In_657,In_1136);
and U332 (N_332,In_355,In_2);
nand U333 (N_333,In_950,In_1355);
nor U334 (N_334,In_351,In_1037);
nor U335 (N_335,In_1170,In_896);
nor U336 (N_336,In_1487,In_314);
or U337 (N_337,In_374,In_73);
nor U338 (N_338,In_721,In_622);
nand U339 (N_339,In_1154,In_798);
nor U340 (N_340,In_40,In_19);
xnor U341 (N_341,In_1267,In_893);
nand U342 (N_342,In_230,In_103);
or U343 (N_343,In_304,In_513);
nor U344 (N_344,In_511,In_1142);
or U345 (N_345,In_1005,In_799);
nor U346 (N_346,In_147,In_540);
and U347 (N_347,In_1110,In_62);
or U348 (N_348,In_88,In_450);
and U349 (N_349,In_257,In_1283);
nand U350 (N_350,In_181,In_1120);
nand U351 (N_351,In_987,In_1311);
or U352 (N_352,In_231,In_1173);
and U353 (N_353,In_861,In_909);
or U354 (N_354,In_362,In_1258);
nor U355 (N_355,In_949,In_638);
nor U356 (N_356,In_468,In_300);
and U357 (N_357,In_832,In_65);
nand U358 (N_358,In_901,In_1458);
and U359 (N_359,In_675,In_1105);
or U360 (N_360,In_1284,In_1066);
and U361 (N_361,In_980,In_486);
nor U362 (N_362,In_479,In_1210);
and U363 (N_363,In_1000,In_1400);
nor U364 (N_364,In_406,In_534);
or U365 (N_365,In_976,In_229);
or U366 (N_366,In_1118,In_284);
and U367 (N_367,In_112,In_897);
and U368 (N_368,In_643,In_1293);
nor U369 (N_369,In_1223,In_627);
and U370 (N_370,In_838,In_1189);
xnor U371 (N_371,In_1168,In_1359);
nor U372 (N_372,In_900,In_401);
and U373 (N_373,In_435,In_120);
and U374 (N_374,In_91,In_33);
and U375 (N_375,In_977,In_1318);
nor U376 (N_376,In_864,In_1494);
xnor U377 (N_377,In_701,In_927);
nor U378 (N_378,In_273,In_719);
and U379 (N_379,In_932,In_912);
and U380 (N_380,In_152,In_998);
nor U381 (N_381,In_882,In_1112);
or U382 (N_382,In_679,In_109);
nor U383 (N_383,In_572,In_820);
and U384 (N_384,In_1069,In_1368);
nor U385 (N_385,In_1315,In_704);
nor U386 (N_386,In_725,In_167);
and U387 (N_387,In_118,In_27);
nand U388 (N_388,In_766,In_783);
nor U389 (N_389,In_988,In_1301);
and U390 (N_390,In_841,In_327);
or U391 (N_391,In_1063,In_1289);
and U392 (N_392,In_808,In_1166);
or U393 (N_393,In_1128,In_227);
and U394 (N_394,In_407,In_1032);
xnor U395 (N_395,In_816,In_883);
nor U396 (N_396,In_488,In_1408);
and U397 (N_397,In_1443,In_921);
or U398 (N_398,In_475,In_282);
and U399 (N_399,In_423,In_272);
nand U400 (N_400,In_270,In_1008);
nor U401 (N_401,In_999,In_289);
nor U402 (N_402,In_1062,In_1076);
or U403 (N_403,In_1040,In_232);
or U404 (N_404,In_959,In_1456);
nand U405 (N_405,In_157,In_1204);
or U406 (N_406,In_881,In_1327);
nand U407 (N_407,In_1140,In_895);
nor U408 (N_408,In_383,In_78);
nor U409 (N_409,In_887,In_241);
and U410 (N_410,In_630,In_1174);
and U411 (N_411,In_179,In_1418);
nand U412 (N_412,In_587,In_451);
nand U413 (N_413,In_1046,In_408);
nand U414 (N_414,In_1472,In_544);
or U415 (N_415,In_554,In_943);
nor U416 (N_416,In_444,In_1206);
nand U417 (N_417,In_196,In_802);
nor U418 (N_418,In_404,In_1497);
nor U419 (N_419,In_842,In_267);
nand U420 (N_420,In_446,In_178);
and U421 (N_421,In_906,In_133);
or U422 (N_422,In_859,In_762);
and U423 (N_423,In_773,In_552);
or U424 (N_424,In_817,In_852);
nor U425 (N_425,In_1378,In_371);
and U426 (N_426,In_551,In_155);
nor U427 (N_427,In_337,In_908);
nand U428 (N_428,In_1344,In_862);
and U429 (N_429,In_935,In_1095);
and U430 (N_430,In_1001,In_1336);
xor U431 (N_431,In_1167,In_207);
or U432 (N_432,In_1462,In_1405);
nor U433 (N_433,In_953,In_439);
nor U434 (N_434,In_160,In_557);
nand U435 (N_435,In_565,In_810);
xnor U436 (N_436,In_620,In_1371);
and U437 (N_437,In_1409,In_23);
nand U438 (N_438,In_1130,In_424);
nand U439 (N_439,In_156,In_1150);
xnor U440 (N_440,In_67,In_1277);
and U441 (N_441,In_696,In_350);
nand U442 (N_442,In_360,In_1424);
or U443 (N_443,In_97,In_526);
and U444 (N_444,In_1366,In_1286);
nand U445 (N_445,In_164,In_326);
and U446 (N_446,In_593,In_894);
nand U447 (N_447,In_849,In_1481);
or U448 (N_448,In_184,In_823);
or U449 (N_449,In_373,In_1269);
nand U450 (N_450,In_603,In_11);
nand U451 (N_451,In_717,In_634);
or U452 (N_452,In_889,In_141);
nor U453 (N_453,In_925,In_646);
nand U454 (N_454,In_145,In_705);
nand U455 (N_455,In_1127,In_432);
xnor U456 (N_456,In_1060,In_964);
xor U457 (N_457,In_425,In_30);
nand U458 (N_458,In_945,In_8);
and U459 (N_459,In_1228,In_942);
nor U460 (N_460,In_956,In_426);
and U461 (N_461,In_452,In_1330);
and U462 (N_462,In_973,In_437);
nand U463 (N_463,In_123,In_24);
and U464 (N_464,In_1253,In_668);
nor U465 (N_465,In_1351,In_779);
or U466 (N_466,In_1364,In_601);
nor U467 (N_467,In_1068,In_1208);
and U468 (N_468,In_1460,In_1019);
xor U469 (N_469,In_1292,In_1058);
nand U470 (N_470,In_343,In_1341);
nand U471 (N_471,In_786,In_1362);
nor U472 (N_472,In_396,In_1213);
or U473 (N_473,In_714,In_1334);
and U474 (N_474,In_937,In_1394);
nor U475 (N_475,In_382,In_611);
nand U476 (N_476,In_331,In_136);
or U477 (N_477,In_1011,In_1052);
xor U478 (N_478,In_1387,In_684);
or U479 (N_479,In_1149,In_354);
nor U480 (N_480,In_441,In_1346);
or U481 (N_481,In_765,In_177);
or U482 (N_482,In_564,In_1278);
or U483 (N_483,In_1471,In_681);
or U484 (N_484,In_482,In_1367);
and U485 (N_485,In_194,In_1489);
nor U486 (N_486,In_1074,In_262);
nand U487 (N_487,In_1416,In_1134);
nand U488 (N_488,In_778,In_918);
and U489 (N_489,In_1488,In_459);
xor U490 (N_490,In_476,In_974);
nor U491 (N_491,In_617,In_1207);
or U492 (N_492,In_455,In_1266);
nor U493 (N_493,In_96,In_237);
and U494 (N_494,In_880,In_693);
nor U495 (N_495,In_495,In_3);
and U496 (N_496,In_206,In_1325);
or U497 (N_497,In_456,In_1106);
and U498 (N_498,In_886,In_1122);
nor U499 (N_499,In_1190,In_1392);
or U500 (N_500,In_571,In_1143);
nor U501 (N_501,In_89,In_249);
and U502 (N_502,In_1433,In_504);
or U503 (N_503,In_146,In_647);
or U504 (N_504,In_851,In_245);
nor U505 (N_505,In_1031,In_1);
and U506 (N_506,In_1111,In_740);
xor U507 (N_507,In_1374,In_7);
nor U508 (N_508,In_876,In_890);
xnor U509 (N_509,In_1429,In_716);
and U510 (N_510,In_106,In_1444);
and U511 (N_511,In_1033,In_228);
or U512 (N_512,In_648,In_1363);
and U513 (N_513,In_86,In_591);
nand U514 (N_514,In_386,In_1137);
or U515 (N_515,In_246,In_12);
nor U516 (N_516,In_639,In_1162);
nor U517 (N_517,In_1022,In_574);
or U518 (N_518,In_911,In_680);
or U519 (N_519,In_595,In_474);
and U520 (N_520,In_174,In_563);
nor U521 (N_521,In_507,In_555);
xnor U522 (N_522,In_243,In_162);
or U523 (N_523,In_1251,In_524);
and U524 (N_524,In_1491,In_1139);
or U525 (N_525,In_979,In_238);
nand U526 (N_526,In_709,In_119);
nor U527 (N_527,In_138,In_398);
or U528 (N_528,In_239,In_891);
nand U529 (N_529,In_878,In_248);
nor U530 (N_530,In_1328,In_834);
nor U531 (N_531,In_586,In_225);
xor U532 (N_532,In_1230,In_1442);
xnor U533 (N_533,In_132,In_21);
or U534 (N_534,In_769,In_1434);
or U535 (N_535,In_536,In_806);
and U536 (N_536,In_418,In_774);
nor U537 (N_537,In_1465,In_113);
and U538 (N_538,In_142,In_553);
or U539 (N_539,In_1243,In_789);
xnor U540 (N_540,In_1468,In_702);
nand U541 (N_541,In_1100,In_311);
nand U542 (N_542,In_531,In_685);
nor U543 (N_543,In_1356,In_1492);
and U544 (N_544,In_673,In_49);
and U545 (N_545,In_860,In_380);
or U546 (N_546,In_458,In_405);
xor U547 (N_547,In_853,In_1474);
nand U548 (N_548,In_1156,In_1291);
and U549 (N_549,In_100,In_1479);
or U550 (N_550,In_1186,In_659);
and U551 (N_551,In_390,In_449);
nand U552 (N_552,In_1413,In_1250);
or U553 (N_553,In_1397,In_500);
nand U554 (N_554,In_1475,In_1101);
nor U555 (N_555,In_144,In_305);
nor U556 (N_556,In_1114,In_1159);
and U557 (N_557,In_278,In_992);
or U558 (N_558,In_697,In_208);
nor U559 (N_559,In_795,In_785);
nor U560 (N_560,In_1338,In_616);
nor U561 (N_561,In_715,In_955);
and U562 (N_562,In_801,In_787);
and U563 (N_563,In_58,In_473);
nand U564 (N_564,In_1495,In_105);
nand U565 (N_565,In_669,In_1288);
and U566 (N_566,In_31,In_645);
xor U567 (N_567,In_1205,In_903);
nand U568 (N_568,In_1419,In_512);
and U569 (N_569,In_971,In_140);
nand U570 (N_570,In_667,In_975);
nand U571 (N_571,In_800,In_357);
or U572 (N_572,In_899,In_414);
nor U573 (N_573,In_487,In_1177);
nor U574 (N_574,In_15,In_742);
or U575 (N_575,In_1329,In_1012);
nor U576 (N_576,In_453,In_1313);
or U577 (N_577,In_1010,In_372);
nand U578 (N_578,In_1337,In_363);
xnor U579 (N_579,In_1126,In_250);
nor U580 (N_580,In_1440,In_963);
nand U581 (N_581,In_566,In_582);
or U582 (N_582,In_1247,In_59);
or U583 (N_583,In_1273,In_1039);
and U584 (N_584,In_1259,In_922);
and U585 (N_585,In_1302,In_957);
nor U586 (N_586,In_1212,In_845);
nand U587 (N_587,In_814,In_916);
and U588 (N_588,In_1426,In_585);
or U589 (N_589,In_470,In_664);
nor U590 (N_590,In_365,In_1386);
nand U591 (N_591,In_150,In_1308);
nand U592 (N_592,In_66,In_1287);
nor U593 (N_593,In_910,In_970);
xnor U594 (N_594,In_478,In_1085);
and U595 (N_595,In_75,In_81);
nand U596 (N_596,In_1448,In_656);
nand U597 (N_597,In_654,In_427);
or U598 (N_598,In_523,In_724);
nor U599 (N_599,In_674,In_954);
and U600 (N_600,In_1092,In_234);
nand U601 (N_601,In_1483,In_711);
nand U602 (N_602,In_1348,In_378);
and U603 (N_603,In_1445,In_757);
and U604 (N_604,In_738,In_549);
or U605 (N_605,In_341,In_188);
nand U606 (N_606,In_60,In_187);
nand U607 (N_607,In_934,In_370);
nand U608 (N_608,In_548,In_505);
or U609 (N_609,In_670,In_1083);
nor U610 (N_610,In_433,In_756);
nor U611 (N_611,In_926,In_115);
xor U612 (N_612,In_1053,In_422);
nand U613 (N_613,In_858,In_108);
and U614 (N_614,In_1382,In_924);
and U615 (N_615,In_1054,In_994);
nand U616 (N_616,In_755,In_38);
nor U617 (N_617,In_55,In_1431);
and U618 (N_618,In_1199,In_1179);
nor U619 (N_619,In_1385,In_1399);
xor U620 (N_620,In_254,In_1125);
nor U621 (N_621,In_708,In_652);
and U622 (N_622,In_658,In_619);
or U623 (N_623,In_35,In_1326);
nand U624 (N_624,In_815,In_268);
or U625 (N_625,In_376,In_1423);
or U626 (N_626,In_1020,In_952);
or U627 (N_627,In_94,In_735);
or U628 (N_628,In_1347,In_1317);
nor U629 (N_629,In_158,In_195);
nand U630 (N_630,In_606,In_1135);
or U631 (N_631,In_1376,In_986);
nand U632 (N_632,In_827,In_1451);
and U633 (N_633,In_159,In_39);
or U634 (N_634,In_600,In_506);
or U635 (N_635,In_824,In_818);
and U636 (N_636,In_1185,In_1260);
or U637 (N_637,In_1038,In_1375);
nor U638 (N_638,In_104,In_535);
and U639 (N_639,In_1254,In_1464);
nor U640 (N_640,In_26,In_666);
or U641 (N_641,In_788,In_867);
nor U642 (N_642,In_50,In_80);
or U643 (N_643,In_1045,In_190);
or U644 (N_644,In_175,In_844);
xor U645 (N_645,In_301,In_1144);
and U646 (N_646,In_1263,In_260);
nor U647 (N_647,In_1485,In_1241);
nor U648 (N_648,In_22,In_122);
nand U649 (N_649,In_1239,In_527);
and U650 (N_650,In_567,In_931);
or U651 (N_651,In_5,In_467);
nor U652 (N_652,In_1197,In_1164);
and U653 (N_653,In_776,In_522);
nor U654 (N_654,In_308,In_1324);
and U655 (N_655,In_461,In_1373);
nand U656 (N_656,In_247,In_276);
nand U657 (N_657,In_1370,In_1034);
xor U658 (N_658,In_508,In_1158);
and U659 (N_659,In_1209,In_342);
and U660 (N_660,In_936,In_1407);
and U661 (N_661,In_1453,In_410);
nand U662 (N_662,In_917,In_340);
and U663 (N_663,In_982,In_1123);
xnor U664 (N_664,In_1119,In_1262);
nor U665 (N_665,In_421,In_720);
and U666 (N_666,In_1065,In_985);
nor U667 (N_667,In_203,In_280);
xor U668 (N_668,In_285,In_972);
and U669 (N_669,In_811,In_137);
xnor U670 (N_670,In_221,In_306);
or U671 (N_671,In_539,In_1309);
nor U672 (N_672,In_93,In_1390);
nand U673 (N_673,In_1271,In_153);
xnor U674 (N_674,In_1437,In_47);
xnor U675 (N_675,In_464,In_353);
and U676 (N_676,In_718,In_6);
xnor U677 (N_677,In_1215,In_1432);
and U678 (N_678,In_197,In_445);
and U679 (N_679,In_846,In_644);
or U680 (N_680,In_9,In_83);
and U681 (N_681,In_366,In_1098);
nand U682 (N_682,In_14,In_349);
nand U683 (N_683,In_1404,In_633);
nor U684 (N_684,In_323,In_573);
nor U685 (N_685,In_51,In_1089);
xor U686 (N_686,In_1294,In_520);
and U687 (N_687,In_829,In_1322);
nor U688 (N_688,In_981,In_54);
or U689 (N_689,In_20,In_528);
or U690 (N_690,In_1412,In_830);
nor U691 (N_691,In_695,In_1121);
and U692 (N_692,In_579,In_1124);
and U693 (N_693,In_677,In_521);
and U694 (N_694,In_690,In_1388);
or U695 (N_695,In_1200,In_1425);
and U696 (N_696,In_1316,In_1203);
nand U697 (N_697,In_393,In_613);
or U698 (N_698,In_722,In_1103);
nand U699 (N_699,In_1088,In_892);
nor U700 (N_700,In_1113,In_615);
or U701 (N_701,In_186,In_173);
nor U702 (N_702,In_392,In_1016);
nand U703 (N_703,In_313,In_1296);
nor U704 (N_704,In_1279,In_837);
nand U705 (N_705,In_295,In_484);
or U706 (N_706,In_303,In_381);
nor U707 (N_707,In_941,In_1056);
nor U708 (N_708,In_923,In_965);
and U709 (N_709,In_1290,In_775);
nor U710 (N_710,In_1043,In_768);
and U711 (N_711,In_869,In_1498);
or U712 (N_712,In_1080,In_728);
and U713 (N_713,In_626,In_95);
or U714 (N_714,In_1217,In_1064);
and U715 (N_715,In_537,In_1131);
xnor U716 (N_716,In_131,In_1145);
or U717 (N_717,In_1406,In_855);
nor U718 (N_718,In_503,In_1402);
nor U719 (N_719,In_448,In_568);
or U720 (N_720,In_723,In_543);
or U721 (N_721,In_1265,In_332);
or U722 (N_722,In_547,In_608);
nor U723 (N_723,In_1466,In_493);
xor U724 (N_724,In_597,In_275);
or U725 (N_725,In_465,In_1107);
or U726 (N_726,In_200,In_562);
nor U727 (N_727,In_663,In_148);
and U728 (N_728,In_1163,In_1231);
and U729 (N_729,In_605,In_1299);
nor U730 (N_730,In_915,In_948);
xor U731 (N_731,In_589,In_1441);
nor U732 (N_732,In_334,In_1153);
nand U733 (N_733,In_1201,In_649);
nand U734 (N_734,In_1079,In_1401);
and U735 (N_735,In_17,In_469);
and U736 (N_736,In_968,In_1295);
or U737 (N_737,In_1384,In_447);
and U738 (N_738,In_483,In_161);
nor U739 (N_739,In_37,In_542);
nand U740 (N_740,In_919,In_84);
or U741 (N_741,In_739,In_1410);
or U742 (N_742,In_1307,In_121);
nand U743 (N_743,In_496,In_1191);
or U744 (N_744,In_807,In_36);
and U745 (N_745,In_1102,In_263);
nand U746 (N_746,In_16,In_905);
nor U747 (N_747,In_997,In_255);
and U748 (N_748,In_1320,In_655);
or U749 (N_749,In_163,In_1436);
nand U750 (N_750,In_323,In_910);
nor U751 (N_751,In_1479,In_1398);
nor U752 (N_752,In_1082,In_130);
nor U753 (N_753,In_1325,In_534);
nand U754 (N_754,In_1032,In_1060);
and U755 (N_755,In_546,In_87);
xor U756 (N_756,In_221,In_1220);
nor U757 (N_757,In_479,In_893);
nor U758 (N_758,In_392,In_901);
nand U759 (N_759,In_25,In_168);
nor U760 (N_760,In_109,In_451);
nor U761 (N_761,In_1324,In_613);
and U762 (N_762,In_459,In_375);
and U763 (N_763,In_947,In_1086);
or U764 (N_764,In_64,In_594);
nand U765 (N_765,In_1170,In_584);
nand U766 (N_766,In_577,In_199);
or U767 (N_767,In_674,In_733);
or U768 (N_768,In_7,In_1033);
nor U769 (N_769,In_938,In_1360);
nor U770 (N_770,In_524,In_42);
nor U771 (N_771,In_644,In_60);
nand U772 (N_772,In_1128,In_1127);
or U773 (N_773,In_1398,In_1446);
xnor U774 (N_774,In_1311,In_1178);
and U775 (N_775,In_1278,In_508);
nand U776 (N_776,In_1264,In_950);
or U777 (N_777,In_325,In_1487);
and U778 (N_778,In_1473,In_504);
nor U779 (N_779,In_860,In_1151);
nand U780 (N_780,In_1055,In_955);
nand U781 (N_781,In_1460,In_1268);
xnor U782 (N_782,In_897,In_1486);
and U783 (N_783,In_598,In_404);
nand U784 (N_784,In_18,In_1446);
or U785 (N_785,In_1133,In_1113);
xnor U786 (N_786,In_712,In_1434);
xor U787 (N_787,In_800,In_144);
and U788 (N_788,In_937,In_737);
nand U789 (N_789,In_1190,In_690);
and U790 (N_790,In_426,In_668);
and U791 (N_791,In_175,In_853);
nand U792 (N_792,In_1371,In_454);
and U793 (N_793,In_778,In_1288);
nor U794 (N_794,In_494,In_783);
or U795 (N_795,In_1297,In_529);
or U796 (N_796,In_531,In_523);
nor U797 (N_797,In_138,In_579);
nand U798 (N_798,In_1233,In_765);
nor U799 (N_799,In_465,In_656);
xnor U800 (N_800,In_1066,In_131);
nor U801 (N_801,In_496,In_443);
xor U802 (N_802,In_606,In_667);
or U803 (N_803,In_546,In_1289);
and U804 (N_804,In_1447,In_405);
nor U805 (N_805,In_6,In_185);
and U806 (N_806,In_1300,In_1221);
nor U807 (N_807,In_1281,In_72);
or U808 (N_808,In_1296,In_83);
or U809 (N_809,In_1033,In_190);
xnor U810 (N_810,In_1086,In_1311);
nand U811 (N_811,In_414,In_572);
or U812 (N_812,In_595,In_1192);
or U813 (N_813,In_246,In_1214);
nor U814 (N_814,In_127,In_1212);
nand U815 (N_815,In_337,In_1305);
nand U816 (N_816,In_96,In_1343);
and U817 (N_817,In_239,In_547);
nor U818 (N_818,In_1030,In_1276);
or U819 (N_819,In_1102,In_428);
nor U820 (N_820,In_1112,In_105);
or U821 (N_821,In_82,In_915);
or U822 (N_822,In_890,In_710);
and U823 (N_823,In_1407,In_979);
nor U824 (N_824,In_42,In_440);
and U825 (N_825,In_229,In_222);
or U826 (N_826,In_199,In_350);
nand U827 (N_827,In_618,In_1436);
nor U828 (N_828,In_33,In_1284);
or U829 (N_829,In_1137,In_1422);
or U830 (N_830,In_964,In_1163);
and U831 (N_831,In_847,In_622);
or U832 (N_832,In_847,In_1377);
xnor U833 (N_833,In_1242,In_12);
nor U834 (N_834,In_671,In_445);
nor U835 (N_835,In_551,In_1312);
nand U836 (N_836,In_972,In_413);
or U837 (N_837,In_910,In_1285);
and U838 (N_838,In_748,In_337);
and U839 (N_839,In_307,In_899);
xnor U840 (N_840,In_132,In_194);
and U841 (N_841,In_665,In_586);
nor U842 (N_842,In_810,In_1010);
and U843 (N_843,In_369,In_725);
nand U844 (N_844,In_714,In_1482);
nand U845 (N_845,In_325,In_504);
nor U846 (N_846,In_905,In_715);
or U847 (N_847,In_721,In_823);
or U848 (N_848,In_769,In_808);
xnor U849 (N_849,In_689,In_546);
or U850 (N_850,In_417,In_907);
and U851 (N_851,In_10,In_411);
nor U852 (N_852,In_1176,In_869);
xnor U853 (N_853,In_900,In_233);
or U854 (N_854,In_152,In_797);
and U855 (N_855,In_1120,In_1113);
and U856 (N_856,In_1322,In_1040);
nand U857 (N_857,In_1467,In_1270);
nand U858 (N_858,In_599,In_1049);
nand U859 (N_859,In_1184,In_1317);
nand U860 (N_860,In_290,In_767);
nor U861 (N_861,In_38,In_1189);
or U862 (N_862,In_1152,In_1368);
nand U863 (N_863,In_327,In_201);
xnor U864 (N_864,In_1120,In_530);
nor U865 (N_865,In_291,In_765);
or U866 (N_866,In_1307,In_1112);
and U867 (N_867,In_742,In_959);
nor U868 (N_868,In_1294,In_797);
and U869 (N_869,In_654,In_38);
or U870 (N_870,In_900,In_957);
nand U871 (N_871,In_1251,In_1323);
nor U872 (N_872,In_459,In_774);
and U873 (N_873,In_146,In_831);
and U874 (N_874,In_917,In_250);
or U875 (N_875,In_163,In_674);
and U876 (N_876,In_563,In_1008);
nor U877 (N_877,In_541,In_430);
and U878 (N_878,In_1074,In_610);
nand U879 (N_879,In_620,In_684);
or U880 (N_880,In_1288,In_1223);
nand U881 (N_881,In_225,In_1306);
or U882 (N_882,In_678,In_1317);
and U883 (N_883,In_1191,In_960);
xor U884 (N_884,In_1486,In_1187);
or U885 (N_885,In_1007,In_555);
or U886 (N_886,In_1156,In_1393);
or U887 (N_887,In_11,In_989);
or U888 (N_888,In_219,In_1431);
or U889 (N_889,In_217,In_1071);
and U890 (N_890,In_1324,In_305);
nor U891 (N_891,In_530,In_1168);
nor U892 (N_892,In_822,In_1366);
and U893 (N_893,In_823,In_1143);
nand U894 (N_894,In_914,In_385);
nand U895 (N_895,In_680,In_1453);
nand U896 (N_896,In_1330,In_512);
nand U897 (N_897,In_30,In_1429);
nor U898 (N_898,In_1424,In_1353);
xnor U899 (N_899,In_553,In_293);
or U900 (N_900,In_582,In_35);
nand U901 (N_901,In_625,In_811);
xnor U902 (N_902,In_895,In_821);
nor U903 (N_903,In_1482,In_1171);
nor U904 (N_904,In_662,In_932);
or U905 (N_905,In_355,In_1136);
or U906 (N_906,In_1361,In_78);
or U907 (N_907,In_55,In_1491);
xor U908 (N_908,In_1256,In_255);
nand U909 (N_909,In_656,In_11);
xor U910 (N_910,In_282,In_955);
or U911 (N_911,In_796,In_561);
nand U912 (N_912,In_6,In_812);
and U913 (N_913,In_556,In_1015);
nor U914 (N_914,In_589,In_371);
xnor U915 (N_915,In_1085,In_709);
or U916 (N_916,In_61,In_485);
or U917 (N_917,In_1389,In_350);
nand U918 (N_918,In_1142,In_28);
nand U919 (N_919,In_164,In_690);
and U920 (N_920,In_1026,In_288);
nor U921 (N_921,In_293,In_727);
and U922 (N_922,In_1239,In_553);
xnor U923 (N_923,In_594,In_1348);
nand U924 (N_924,In_1494,In_1099);
nor U925 (N_925,In_1096,In_1057);
and U926 (N_926,In_1379,In_433);
xnor U927 (N_927,In_167,In_808);
or U928 (N_928,In_161,In_887);
nand U929 (N_929,In_1395,In_532);
xor U930 (N_930,In_1104,In_819);
nand U931 (N_931,In_191,In_1073);
and U932 (N_932,In_627,In_836);
nand U933 (N_933,In_781,In_65);
nand U934 (N_934,In_1002,In_884);
and U935 (N_935,In_1429,In_1272);
nor U936 (N_936,In_541,In_1351);
nor U937 (N_937,In_586,In_605);
nor U938 (N_938,In_271,In_1113);
xor U939 (N_939,In_1289,In_646);
and U940 (N_940,In_335,In_94);
and U941 (N_941,In_288,In_1105);
nor U942 (N_942,In_122,In_1309);
and U943 (N_943,In_1109,In_331);
or U944 (N_944,In_914,In_171);
xnor U945 (N_945,In_230,In_860);
nor U946 (N_946,In_568,In_1107);
nor U947 (N_947,In_136,In_383);
nor U948 (N_948,In_497,In_999);
or U949 (N_949,In_617,In_780);
xnor U950 (N_950,In_682,In_185);
or U951 (N_951,In_1241,In_13);
nand U952 (N_952,In_388,In_1162);
or U953 (N_953,In_173,In_623);
or U954 (N_954,In_1045,In_785);
nor U955 (N_955,In_974,In_415);
nand U956 (N_956,In_767,In_137);
nor U957 (N_957,In_1259,In_823);
nor U958 (N_958,In_894,In_750);
or U959 (N_959,In_1218,In_1030);
and U960 (N_960,In_589,In_1217);
and U961 (N_961,In_881,In_309);
nand U962 (N_962,In_42,In_1013);
nor U963 (N_963,In_217,In_224);
or U964 (N_964,In_204,In_426);
or U965 (N_965,In_1062,In_1200);
nand U966 (N_966,In_1180,In_1182);
and U967 (N_967,In_1444,In_202);
nor U968 (N_968,In_1116,In_505);
nor U969 (N_969,In_1430,In_1244);
nand U970 (N_970,In_1482,In_785);
or U971 (N_971,In_113,In_81);
or U972 (N_972,In_1147,In_1476);
nand U973 (N_973,In_615,In_542);
or U974 (N_974,In_356,In_1205);
nor U975 (N_975,In_8,In_730);
nand U976 (N_976,In_504,In_905);
nor U977 (N_977,In_1478,In_183);
or U978 (N_978,In_460,In_806);
nor U979 (N_979,In_933,In_1373);
and U980 (N_980,In_337,In_438);
xnor U981 (N_981,In_1060,In_571);
and U982 (N_982,In_347,In_841);
and U983 (N_983,In_670,In_1049);
xor U984 (N_984,In_97,In_914);
and U985 (N_985,In_50,In_9);
nand U986 (N_986,In_10,In_841);
and U987 (N_987,In_1493,In_1106);
xor U988 (N_988,In_1090,In_930);
and U989 (N_989,In_910,In_1333);
or U990 (N_990,In_1336,In_597);
xor U991 (N_991,In_703,In_1278);
nand U992 (N_992,In_1358,In_442);
or U993 (N_993,In_285,In_1098);
and U994 (N_994,In_326,In_443);
nand U995 (N_995,In_1356,In_150);
nor U996 (N_996,In_1270,In_284);
nand U997 (N_997,In_1050,In_1497);
or U998 (N_998,In_594,In_1205);
nand U999 (N_999,In_1277,In_1132);
and U1000 (N_1000,In_1018,In_1347);
or U1001 (N_1001,In_899,In_600);
or U1002 (N_1002,In_841,In_689);
or U1003 (N_1003,In_510,In_652);
nand U1004 (N_1004,In_388,In_1224);
nand U1005 (N_1005,In_838,In_1042);
and U1006 (N_1006,In_303,In_1161);
nor U1007 (N_1007,In_115,In_1204);
or U1008 (N_1008,In_754,In_1285);
and U1009 (N_1009,In_523,In_546);
nor U1010 (N_1010,In_389,In_1212);
and U1011 (N_1011,In_590,In_382);
or U1012 (N_1012,In_798,In_1414);
nand U1013 (N_1013,In_1334,In_1176);
or U1014 (N_1014,In_989,In_329);
nand U1015 (N_1015,In_525,In_572);
or U1016 (N_1016,In_679,In_1017);
nor U1017 (N_1017,In_1114,In_1112);
nor U1018 (N_1018,In_1401,In_548);
xor U1019 (N_1019,In_508,In_1015);
xnor U1020 (N_1020,In_1149,In_1078);
and U1021 (N_1021,In_663,In_420);
xor U1022 (N_1022,In_565,In_395);
and U1023 (N_1023,In_471,In_785);
or U1024 (N_1024,In_253,In_1094);
and U1025 (N_1025,In_655,In_1422);
or U1026 (N_1026,In_483,In_366);
or U1027 (N_1027,In_267,In_1179);
nor U1028 (N_1028,In_477,In_517);
and U1029 (N_1029,In_744,In_831);
and U1030 (N_1030,In_740,In_1122);
and U1031 (N_1031,In_1066,In_804);
or U1032 (N_1032,In_904,In_580);
or U1033 (N_1033,In_868,In_1172);
or U1034 (N_1034,In_62,In_1132);
nand U1035 (N_1035,In_561,In_1327);
nand U1036 (N_1036,In_1066,In_471);
nand U1037 (N_1037,In_101,In_565);
and U1038 (N_1038,In_883,In_749);
nand U1039 (N_1039,In_32,In_264);
or U1040 (N_1040,In_784,In_890);
or U1041 (N_1041,In_117,In_214);
nor U1042 (N_1042,In_374,In_1023);
and U1043 (N_1043,In_195,In_773);
nor U1044 (N_1044,In_200,In_207);
or U1045 (N_1045,In_859,In_617);
nand U1046 (N_1046,In_1399,In_1332);
nor U1047 (N_1047,In_982,In_828);
nand U1048 (N_1048,In_681,In_836);
or U1049 (N_1049,In_1288,In_287);
and U1050 (N_1050,In_741,In_902);
and U1051 (N_1051,In_543,In_1011);
or U1052 (N_1052,In_633,In_938);
nand U1053 (N_1053,In_1121,In_263);
and U1054 (N_1054,In_1217,In_78);
or U1055 (N_1055,In_933,In_158);
or U1056 (N_1056,In_1494,In_970);
or U1057 (N_1057,In_1099,In_90);
and U1058 (N_1058,In_312,In_684);
nand U1059 (N_1059,In_130,In_1462);
and U1060 (N_1060,In_652,In_338);
and U1061 (N_1061,In_624,In_198);
or U1062 (N_1062,In_716,In_742);
nor U1063 (N_1063,In_942,In_896);
nor U1064 (N_1064,In_903,In_1019);
or U1065 (N_1065,In_1032,In_7);
or U1066 (N_1066,In_666,In_561);
xor U1067 (N_1067,In_180,In_165);
or U1068 (N_1068,In_440,In_684);
or U1069 (N_1069,In_954,In_567);
xnor U1070 (N_1070,In_1296,In_418);
nand U1071 (N_1071,In_373,In_284);
and U1072 (N_1072,In_333,In_637);
nand U1073 (N_1073,In_685,In_1484);
nor U1074 (N_1074,In_1463,In_677);
and U1075 (N_1075,In_825,In_1389);
nand U1076 (N_1076,In_1087,In_433);
and U1077 (N_1077,In_339,In_1249);
xor U1078 (N_1078,In_256,In_1332);
nand U1079 (N_1079,In_1113,In_1157);
nor U1080 (N_1080,In_1357,In_1328);
nand U1081 (N_1081,In_71,In_1366);
xnor U1082 (N_1082,In_397,In_1035);
nor U1083 (N_1083,In_578,In_1208);
or U1084 (N_1084,In_81,In_288);
and U1085 (N_1085,In_215,In_1423);
or U1086 (N_1086,In_18,In_1326);
and U1087 (N_1087,In_494,In_806);
and U1088 (N_1088,In_1034,In_775);
nand U1089 (N_1089,In_434,In_1368);
and U1090 (N_1090,In_447,In_90);
and U1091 (N_1091,In_648,In_550);
nor U1092 (N_1092,In_648,In_1072);
nand U1093 (N_1093,In_764,In_1403);
and U1094 (N_1094,In_1459,In_691);
or U1095 (N_1095,In_1127,In_697);
or U1096 (N_1096,In_1179,In_152);
xor U1097 (N_1097,In_703,In_814);
or U1098 (N_1098,In_904,In_1185);
and U1099 (N_1099,In_490,In_1044);
nor U1100 (N_1100,In_855,In_1126);
nand U1101 (N_1101,In_1127,In_116);
nor U1102 (N_1102,In_927,In_666);
nand U1103 (N_1103,In_992,In_231);
or U1104 (N_1104,In_574,In_133);
nor U1105 (N_1105,In_1378,In_118);
or U1106 (N_1106,In_1083,In_1348);
nor U1107 (N_1107,In_827,In_1128);
and U1108 (N_1108,In_1334,In_621);
xnor U1109 (N_1109,In_651,In_943);
nor U1110 (N_1110,In_163,In_488);
or U1111 (N_1111,In_377,In_523);
nand U1112 (N_1112,In_434,In_1194);
and U1113 (N_1113,In_1244,In_959);
nand U1114 (N_1114,In_634,In_122);
nor U1115 (N_1115,In_1184,In_68);
or U1116 (N_1116,In_636,In_635);
xor U1117 (N_1117,In_82,In_1474);
nand U1118 (N_1118,In_55,In_603);
nand U1119 (N_1119,In_97,In_617);
nand U1120 (N_1120,In_590,In_607);
nand U1121 (N_1121,In_1074,In_219);
xor U1122 (N_1122,In_105,In_1417);
nor U1123 (N_1123,In_923,In_901);
and U1124 (N_1124,In_44,In_189);
and U1125 (N_1125,In_917,In_988);
nand U1126 (N_1126,In_718,In_141);
nor U1127 (N_1127,In_552,In_1345);
nor U1128 (N_1128,In_589,In_1494);
xnor U1129 (N_1129,In_627,In_736);
and U1130 (N_1130,In_1232,In_1429);
nor U1131 (N_1131,In_231,In_165);
or U1132 (N_1132,In_1056,In_737);
or U1133 (N_1133,In_24,In_892);
and U1134 (N_1134,In_844,In_1222);
xnor U1135 (N_1135,In_823,In_218);
or U1136 (N_1136,In_1081,In_1355);
xnor U1137 (N_1137,In_830,In_1452);
nor U1138 (N_1138,In_804,In_592);
nor U1139 (N_1139,In_617,In_1055);
nor U1140 (N_1140,In_504,In_326);
or U1141 (N_1141,In_1401,In_1000);
or U1142 (N_1142,In_1466,In_1011);
and U1143 (N_1143,In_1383,In_681);
nor U1144 (N_1144,In_146,In_1159);
or U1145 (N_1145,In_1188,In_247);
nand U1146 (N_1146,In_706,In_509);
or U1147 (N_1147,In_222,In_669);
or U1148 (N_1148,In_568,In_1031);
or U1149 (N_1149,In_183,In_1113);
or U1150 (N_1150,In_19,In_256);
xor U1151 (N_1151,In_130,In_607);
or U1152 (N_1152,In_162,In_751);
nand U1153 (N_1153,In_686,In_1175);
nand U1154 (N_1154,In_369,In_195);
nor U1155 (N_1155,In_1058,In_382);
or U1156 (N_1156,In_515,In_1429);
and U1157 (N_1157,In_120,In_878);
nand U1158 (N_1158,In_589,In_1134);
and U1159 (N_1159,In_1361,In_491);
nor U1160 (N_1160,In_1396,In_623);
nor U1161 (N_1161,In_34,In_496);
xnor U1162 (N_1162,In_569,In_375);
and U1163 (N_1163,In_1229,In_404);
and U1164 (N_1164,In_164,In_643);
or U1165 (N_1165,In_931,In_789);
and U1166 (N_1166,In_1135,In_113);
and U1167 (N_1167,In_616,In_1099);
and U1168 (N_1168,In_935,In_117);
nand U1169 (N_1169,In_1105,In_227);
nand U1170 (N_1170,In_1104,In_291);
nor U1171 (N_1171,In_1493,In_860);
or U1172 (N_1172,In_383,In_53);
xnor U1173 (N_1173,In_821,In_673);
nor U1174 (N_1174,In_48,In_538);
and U1175 (N_1175,In_127,In_1169);
xnor U1176 (N_1176,In_1313,In_119);
and U1177 (N_1177,In_174,In_812);
nand U1178 (N_1178,In_448,In_530);
nand U1179 (N_1179,In_812,In_71);
or U1180 (N_1180,In_188,In_1249);
nor U1181 (N_1181,In_356,In_384);
and U1182 (N_1182,In_869,In_644);
or U1183 (N_1183,In_496,In_468);
and U1184 (N_1184,In_1493,In_1225);
and U1185 (N_1185,In_397,In_1420);
and U1186 (N_1186,In_913,In_48);
and U1187 (N_1187,In_1287,In_307);
nand U1188 (N_1188,In_1228,In_872);
or U1189 (N_1189,In_1472,In_740);
nand U1190 (N_1190,In_84,In_1348);
and U1191 (N_1191,In_73,In_1463);
nand U1192 (N_1192,In_251,In_973);
and U1193 (N_1193,In_37,In_105);
and U1194 (N_1194,In_563,In_55);
and U1195 (N_1195,In_1132,In_243);
and U1196 (N_1196,In_95,In_1152);
xnor U1197 (N_1197,In_561,In_275);
and U1198 (N_1198,In_1372,In_742);
nor U1199 (N_1199,In_1329,In_1220);
and U1200 (N_1200,In_1132,In_596);
nand U1201 (N_1201,In_1471,In_1054);
nand U1202 (N_1202,In_1311,In_278);
xnor U1203 (N_1203,In_341,In_818);
or U1204 (N_1204,In_807,In_727);
nor U1205 (N_1205,In_247,In_198);
nand U1206 (N_1206,In_81,In_443);
nand U1207 (N_1207,In_1245,In_1052);
nor U1208 (N_1208,In_27,In_347);
or U1209 (N_1209,In_1397,In_36);
or U1210 (N_1210,In_558,In_477);
nor U1211 (N_1211,In_1124,In_383);
xnor U1212 (N_1212,In_1296,In_427);
nand U1213 (N_1213,In_115,In_895);
or U1214 (N_1214,In_1152,In_454);
xor U1215 (N_1215,In_345,In_1413);
or U1216 (N_1216,In_1403,In_684);
nor U1217 (N_1217,In_1064,In_711);
or U1218 (N_1218,In_562,In_1467);
and U1219 (N_1219,In_488,In_1297);
nor U1220 (N_1220,In_295,In_251);
and U1221 (N_1221,In_1450,In_1146);
and U1222 (N_1222,In_209,In_269);
and U1223 (N_1223,In_863,In_2);
nand U1224 (N_1224,In_154,In_1048);
nor U1225 (N_1225,In_233,In_1035);
nand U1226 (N_1226,In_941,In_765);
nor U1227 (N_1227,In_1290,In_277);
xor U1228 (N_1228,In_1097,In_1265);
nor U1229 (N_1229,In_232,In_1127);
or U1230 (N_1230,In_622,In_682);
or U1231 (N_1231,In_1200,In_566);
or U1232 (N_1232,In_46,In_422);
xor U1233 (N_1233,In_586,In_1060);
or U1234 (N_1234,In_940,In_797);
or U1235 (N_1235,In_536,In_1258);
nor U1236 (N_1236,In_553,In_412);
nand U1237 (N_1237,In_300,In_603);
and U1238 (N_1238,In_45,In_47);
or U1239 (N_1239,In_892,In_796);
nor U1240 (N_1240,In_29,In_675);
and U1241 (N_1241,In_1235,In_365);
xnor U1242 (N_1242,In_979,In_960);
or U1243 (N_1243,In_1208,In_195);
and U1244 (N_1244,In_1059,In_116);
or U1245 (N_1245,In_1010,In_162);
nand U1246 (N_1246,In_1051,In_955);
nand U1247 (N_1247,In_206,In_1391);
and U1248 (N_1248,In_1029,In_845);
and U1249 (N_1249,In_1229,In_1275);
xnor U1250 (N_1250,In_607,In_1249);
nand U1251 (N_1251,In_281,In_261);
or U1252 (N_1252,In_1302,In_938);
nor U1253 (N_1253,In_1054,In_1236);
and U1254 (N_1254,In_333,In_601);
nor U1255 (N_1255,In_709,In_1079);
nor U1256 (N_1256,In_1495,In_1336);
nand U1257 (N_1257,In_451,In_162);
or U1258 (N_1258,In_525,In_1412);
and U1259 (N_1259,In_871,In_337);
or U1260 (N_1260,In_1279,In_1355);
and U1261 (N_1261,In_1021,In_465);
nor U1262 (N_1262,In_1448,In_1390);
or U1263 (N_1263,In_163,In_874);
nand U1264 (N_1264,In_1449,In_1138);
or U1265 (N_1265,In_317,In_225);
nor U1266 (N_1266,In_771,In_975);
or U1267 (N_1267,In_1263,In_1416);
and U1268 (N_1268,In_433,In_497);
and U1269 (N_1269,In_604,In_742);
or U1270 (N_1270,In_1396,In_903);
and U1271 (N_1271,In_1478,In_368);
nor U1272 (N_1272,In_259,In_1447);
xnor U1273 (N_1273,In_1472,In_1380);
xor U1274 (N_1274,In_1335,In_313);
or U1275 (N_1275,In_1460,In_340);
and U1276 (N_1276,In_791,In_1408);
nor U1277 (N_1277,In_1360,In_1229);
and U1278 (N_1278,In_1353,In_247);
or U1279 (N_1279,In_1205,In_196);
nor U1280 (N_1280,In_1473,In_193);
or U1281 (N_1281,In_161,In_584);
nor U1282 (N_1282,In_365,In_718);
nand U1283 (N_1283,In_482,In_445);
xnor U1284 (N_1284,In_144,In_1188);
or U1285 (N_1285,In_966,In_1002);
xnor U1286 (N_1286,In_233,In_200);
xnor U1287 (N_1287,In_139,In_565);
nor U1288 (N_1288,In_1371,In_215);
nand U1289 (N_1289,In_1204,In_137);
nor U1290 (N_1290,In_939,In_144);
and U1291 (N_1291,In_1425,In_458);
and U1292 (N_1292,In_625,In_643);
nor U1293 (N_1293,In_1494,In_823);
and U1294 (N_1294,In_685,In_639);
nand U1295 (N_1295,In_308,In_428);
nand U1296 (N_1296,In_388,In_1453);
or U1297 (N_1297,In_671,In_1460);
nand U1298 (N_1298,In_785,In_1329);
or U1299 (N_1299,In_248,In_10);
nor U1300 (N_1300,In_196,In_696);
and U1301 (N_1301,In_565,In_711);
or U1302 (N_1302,In_141,In_602);
and U1303 (N_1303,In_283,In_412);
nand U1304 (N_1304,In_536,In_308);
or U1305 (N_1305,In_634,In_281);
nor U1306 (N_1306,In_1356,In_508);
and U1307 (N_1307,In_810,In_175);
nand U1308 (N_1308,In_662,In_1172);
nand U1309 (N_1309,In_499,In_1291);
and U1310 (N_1310,In_660,In_1171);
and U1311 (N_1311,In_1335,In_430);
nor U1312 (N_1312,In_490,In_1346);
nand U1313 (N_1313,In_379,In_518);
nand U1314 (N_1314,In_501,In_562);
and U1315 (N_1315,In_66,In_754);
or U1316 (N_1316,In_1430,In_1362);
nor U1317 (N_1317,In_1027,In_134);
nand U1318 (N_1318,In_1355,In_852);
and U1319 (N_1319,In_1310,In_344);
nand U1320 (N_1320,In_1183,In_1333);
nand U1321 (N_1321,In_681,In_655);
nand U1322 (N_1322,In_862,In_474);
nor U1323 (N_1323,In_796,In_160);
or U1324 (N_1324,In_430,In_823);
nand U1325 (N_1325,In_882,In_1074);
nand U1326 (N_1326,In_1329,In_1112);
and U1327 (N_1327,In_1197,In_1380);
nand U1328 (N_1328,In_1279,In_149);
or U1329 (N_1329,In_60,In_652);
xnor U1330 (N_1330,In_268,In_872);
and U1331 (N_1331,In_605,In_20);
or U1332 (N_1332,In_1458,In_120);
or U1333 (N_1333,In_1319,In_33);
nand U1334 (N_1334,In_121,In_431);
nand U1335 (N_1335,In_671,In_1194);
and U1336 (N_1336,In_873,In_397);
xnor U1337 (N_1337,In_376,In_576);
nand U1338 (N_1338,In_41,In_963);
xor U1339 (N_1339,In_460,In_174);
nand U1340 (N_1340,In_616,In_731);
or U1341 (N_1341,In_906,In_1419);
or U1342 (N_1342,In_1318,In_699);
and U1343 (N_1343,In_1088,In_350);
nand U1344 (N_1344,In_483,In_1194);
nand U1345 (N_1345,In_1016,In_1163);
nor U1346 (N_1346,In_21,In_547);
and U1347 (N_1347,In_939,In_1443);
or U1348 (N_1348,In_1232,In_634);
or U1349 (N_1349,In_160,In_69);
or U1350 (N_1350,In_165,In_335);
and U1351 (N_1351,In_1403,In_1079);
or U1352 (N_1352,In_518,In_198);
and U1353 (N_1353,In_825,In_532);
and U1354 (N_1354,In_1284,In_1292);
nor U1355 (N_1355,In_862,In_851);
nand U1356 (N_1356,In_736,In_484);
nand U1357 (N_1357,In_786,In_524);
xor U1358 (N_1358,In_364,In_81);
nor U1359 (N_1359,In_1228,In_1338);
nor U1360 (N_1360,In_1046,In_1017);
nand U1361 (N_1361,In_38,In_371);
or U1362 (N_1362,In_926,In_48);
nor U1363 (N_1363,In_1481,In_767);
and U1364 (N_1364,In_744,In_1325);
xnor U1365 (N_1365,In_187,In_876);
and U1366 (N_1366,In_509,In_401);
nand U1367 (N_1367,In_560,In_1107);
nand U1368 (N_1368,In_1311,In_783);
and U1369 (N_1369,In_814,In_1089);
and U1370 (N_1370,In_916,In_817);
xor U1371 (N_1371,In_1323,In_1176);
or U1372 (N_1372,In_1026,In_9);
nand U1373 (N_1373,In_521,In_997);
nand U1374 (N_1374,In_766,In_1332);
nor U1375 (N_1375,In_97,In_501);
nand U1376 (N_1376,In_772,In_356);
nand U1377 (N_1377,In_240,In_895);
nor U1378 (N_1378,In_120,In_1153);
and U1379 (N_1379,In_545,In_913);
or U1380 (N_1380,In_1383,In_1421);
or U1381 (N_1381,In_832,In_705);
or U1382 (N_1382,In_424,In_972);
nor U1383 (N_1383,In_408,In_1416);
nand U1384 (N_1384,In_722,In_502);
nand U1385 (N_1385,In_619,In_827);
nor U1386 (N_1386,In_376,In_226);
xor U1387 (N_1387,In_1282,In_1292);
or U1388 (N_1388,In_681,In_61);
nand U1389 (N_1389,In_288,In_365);
and U1390 (N_1390,In_821,In_1279);
or U1391 (N_1391,In_931,In_1020);
and U1392 (N_1392,In_223,In_194);
and U1393 (N_1393,In_1480,In_513);
xnor U1394 (N_1394,In_237,In_153);
nand U1395 (N_1395,In_366,In_577);
nand U1396 (N_1396,In_808,In_1234);
or U1397 (N_1397,In_737,In_931);
or U1398 (N_1398,In_938,In_705);
nor U1399 (N_1399,In_82,In_1478);
or U1400 (N_1400,In_810,In_958);
or U1401 (N_1401,In_574,In_1068);
nor U1402 (N_1402,In_764,In_766);
or U1403 (N_1403,In_777,In_1028);
or U1404 (N_1404,In_284,In_1169);
and U1405 (N_1405,In_181,In_927);
nor U1406 (N_1406,In_380,In_557);
or U1407 (N_1407,In_1076,In_190);
nor U1408 (N_1408,In_1248,In_625);
or U1409 (N_1409,In_538,In_1130);
nor U1410 (N_1410,In_964,In_588);
and U1411 (N_1411,In_330,In_654);
nand U1412 (N_1412,In_229,In_392);
nor U1413 (N_1413,In_646,In_338);
nor U1414 (N_1414,In_432,In_1187);
and U1415 (N_1415,In_536,In_987);
nand U1416 (N_1416,In_221,In_917);
nor U1417 (N_1417,In_941,In_502);
nor U1418 (N_1418,In_1110,In_224);
nand U1419 (N_1419,In_1173,In_1165);
and U1420 (N_1420,In_1254,In_74);
nor U1421 (N_1421,In_1297,In_687);
nand U1422 (N_1422,In_412,In_423);
and U1423 (N_1423,In_465,In_89);
and U1424 (N_1424,In_886,In_1155);
nand U1425 (N_1425,In_547,In_395);
and U1426 (N_1426,In_632,In_645);
and U1427 (N_1427,In_1425,In_1102);
nor U1428 (N_1428,In_698,In_94);
nand U1429 (N_1429,In_407,In_1431);
or U1430 (N_1430,In_196,In_337);
nor U1431 (N_1431,In_107,In_769);
and U1432 (N_1432,In_337,In_313);
and U1433 (N_1433,In_466,In_360);
xnor U1434 (N_1434,In_609,In_438);
or U1435 (N_1435,In_515,In_315);
nor U1436 (N_1436,In_667,In_40);
and U1437 (N_1437,In_991,In_48);
or U1438 (N_1438,In_592,In_80);
nor U1439 (N_1439,In_1472,In_719);
or U1440 (N_1440,In_1432,In_368);
xor U1441 (N_1441,In_1192,In_1499);
and U1442 (N_1442,In_921,In_530);
or U1443 (N_1443,In_671,In_237);
nor U1444 (N_1444,In_218,In_1253);
and U1445 (N_1445,In_1270,In_805);
or U1446 (N_1446,In_1305,In_422);
nor U1447 (N_1447,In_1079,In_1262);
nor U1448 (N_1448,In_1085,In_296);
nor U1449 (N_1449,In_473,In_1385);
xor U1450 (N_1450,In_345,In_926);
nand U1451 (N_1451,In_385,In_442);
or U1452 (N_1452,In_1018,In_1231);
xnor U1453 (N_1453,In_1330,In_617);
or U1454 (N_1454,In_846,In_1053);
and U1455 (N_1455,In_266,In_1031);
nor U1456 (N_1456,In_11,In_1394);
and U1457 (N_1457,In_666,In_749);
or U1458 (N_1458,In_26,In_1449);
nand U1459 (N_1459,In_876,In_111);
nor U1460 (N_1460,In_998,In_192);
nor U1461 (N_1461,In_1296,In_116);
or U1462 (N_1462,In_596,In_141);
nand U1463 (N_1463,In_563,In_217);
nand U1464 (N_1464,In_650,In_1217);
nor U1465 (N_1465,In_951,In_1030);
nor U1466 (N_1466,In_1303,In_809);
or U1467 (N_1467,In_371,In_211);
and U1468 (N_1468,In_1004,In_834);
nand U1469 (N_1469,In_1337,In_883);
and U1470 (N_1470,In_1114,In_1350);
or U1471 (N_1471,In_327,In_862);
nand U1472 (N_1472,In_44,In_194);
or U1473 (N_1473,In_836,In_740);
or U1474 (N_1474,In_147,In_952);
nand U1475 (N_1475,In_998,In_598);
nand U1476 (N_1476,In_1040,In_1044);
or U1477 (N_1477,In_523,In_83);
and U1478 (N_1478,In_108,In_1243);
nand U1479 (N_1479,In_1215,In_445);
xnor U1480 (N_1480,In_573,In_565);
nor U1481 (N_1481,In_627,In_1220);
or U1482 (N_1482,In_396,In_221);
xnor U1483 (N_1483,In_433,In_1444);
nand U1484 (N_1484,In_1186,In_944);
nand U1485 (N_1485,In_1467,In_1389);
and U1486 (N_1486,In_1387,In_1148);
nor U1487 (N_1487,In_162,In_354);
and U1488 (N_1488,In_1016,In_1242);
and U1489 (N_1489,In_63,In_1443);
nor U1490 (N_1490,In_615,In_901);
nor U1491 (N_1491,In_798,In_487);
and U1492 (N_1492,In_776,In_663);
or U1493 (N_1493,In_587,In_340);
or U1494 (N_1494,In_588,In_1397);
or U1495 (N_1495,In_654,In_1227);
xor U1496 (N_1496,In_260,In_327);
or U1497 (N_1497,In_1247,In_534);
and U1498 (N_1498,In_887,In_1097);
nor U1499 (N_1499,In_1120,In_599);
or U1500 (N_1500,In_1348,In_125);
nand U1501 (N_1501,In_705,In_53);
or U1502 (N_1502,In_494,In_673);
and U1503 (N_1503,In_995,In_1219);
nand U1504 (N_1504,In_147,In_843);
and U1505 (N_1505,In_189,In_1175);
and U1506 (N_1506,In_654,In_1398);
xor U1507 (N_1507,In_1195,In_869);
and U1508 (N_1508,In_791,In_306);
nand U1509 (N_1509,In_771,In_1387);
nor U1510 (N_1510,In_742,In_469);
and U1511 (N_1511,In_858,In_1044);
or U1512 (N_1512,In_1038,In_1000);
nand U1513 (N_1513,In_1252,In_96);
xnor U1514 (N_1514,In_1464,In_1396);
or U1515 (N_1515,In_168,In_424);
nand U1516 (N_1516,In_1051,In_519);
or U1517 (N_1517,In_981,In_188);
nand U1518 (N_1518,In_948,In_283);
and U1519 (N_1519,In_535,In_265);
xor U1520 (N_1520,In_127,In_930);
nand U1521 (N_1521,In_383,In_70);
and U1522 (N_1522,In_1485,In_673);
and U1523 (N_1523,In_63,In_1499);
xnor U1524 (N_1524,In_704,In_1397);
xor U1525 (N_1525,In_271,In_130);
nor U1526 (N_1526,In_312,In_275);
and U1527 (N_1527,In_223,In_444);
and U1528 (N_1528,In_66,In_854);
nand U1529 (N_1529,In_1170,In_954);
or U1530 (N_1530,In_1149,In_805);
or U1531 (N_1531,In_1415,In_642);
nand U1532 (N_1532,In_284,In_879);
or U1533 (N_1533,In_1050,In_643);
nand U1534 (N_1534,In_524,In_897);
or U1535 (N_1535,In_408,In_1465);
nand U1536 (N_1536,In_1223,In_739);
nand U1537 (N_1537,In_476,In_1452);
nor U1538 (N_1538,In_864,In_259);
or U1539 (N_1539,In_457,In_237);
nor U1540 (N_1540,In_496,In_314);
xor U1541 (N_1541,In_1143,In_414);
or U1542 (N_1542,In_837,In_280);
nor U1543 (N_1543,In_992,In_347);
and U1544 (N_1544,In_900,In_899);
nand U1545 (N_1545,In_15,In_1417);
and U1546 (N_1546,In_1454,In_1292);
and U1547 (N_1547,In_1263,In_993);
xor U1548 (N_1548,In_1305,In_770);
xor U1549 (N_1549,In_1426,In_1086);
xnor U1550 (N_1550,In_190,In_17);
nor U1551 (N_1551,In_882,In_1157);
or U1552 (N_1552,In_653,In_107);
and U1553 (N_1553,In_128,In_55);
nand U1554 (N_1554,In_1376,In_607);
nand U1555 (N_1555,In_409,In_744);
nor U1556 (N_1556,In_143,In_1203);
nand U1557 (N_1557,In_355,In_487);
nor U1558 (N_1558,In_428,In_229);
or U1559 (N_1559,In_762,In_1411);
nor U1560 (N_1560,In_1016,In_1138);
or U1561 (N_1561,In_1331,In_991);
nand U1562 (N_1562,In_721,In_1029);
nand U1563 (N_1563,In_1277,In_277);
xor U1564 (N_1564,In_23,In_1235);
nand U1565 (N_1565,In_1107,In_385);
nor U1566 (N_1566,In_293,In_65);
nor U1567 (N_1567,In_1382,In_660);
and U1568 (N_1568,In_746,In_163);
nand U1569 (N_1569,In_839,In_842);
nand U1570 (N_1570,In_1248,In_77);
and U1571 (N_1571,In_688,In_1400);
nor U1572 (N_1572,In_1170,In_205);
nor U1573 (N_1573,In_386,In_1465);
and U1574 (N_1574,In_1385,In_110);
nor U1575 (N_1575,In_1445,In_604);
xor U1576 (N_1576,In_294,In_1026);
nand U1577 (N_1577,In_800,In_1481);
or U1578 (N_1578,In_616,In_1157);
nor U1579 (N_1579,In_33,In_1123);
or U1580 (N_1580,In_1387,In_122);
and U1581 (N_1581,In_254,In_580);
nor U1582 (N_1582,In_1001,In_1452);
nor U1583 (N_1583,In_1474,In_1310);
and U1584 (N_1584,In_537,In_216);
xor U1585 (N_1585,In_201,In_898);
nor U1586 (N_1586,In_1170,In_556);
xor U1587 (N_1587,In_1028,In_789);
nand U1588 (N_1588,In_764,In_39);
xor U1589 (N_1589,In_508,In_1471);
nor U1590 (N_1590,In_1286,In_1272);
or U1591 (N_1591,In_1028,In_440);
or U1592 (N_1592,In_111,In_669);
nor U1593 (N_1593,In_850,In_311);
xor U1594 (N_1594,In_1410,In_818);
or U1595 (N_1595,In_1330,In_865);
nor U1596 (N_1596,In_266,In_971);
nor U1597 (N_1597,In_709,In_531);
nand U1598 (N_1598,In_497,In_1059);
nand U1599 (N_1599,In_1253,In_659);
nand U1600 (N_1600,In_706,In_689);
nand U1601 (N_1601,In_1395,In_416);
and U1602 (N_1602,In_879,In_363);
or U1603 (N_1603,In_1077,In_506);
xor U1604 (N_1604,In_763,In_727);
xnor U1605 (N_1605,In_1269,In_1425);
xnor U1606 (N_1606,In_1182,In_825);
nor U1607 (N_1607,In_146,In_1416);
and U1608 (N_1608,In_668,In_481);
and U1609 (N_1609,In_511,In_291);
nor U1610 (N_1610,In_551,In_1133);
nand U1611 (N_1611,In_1038,In_1489);
or U1612 (N_1612,In_237,In_914);
or U1613 (N_1613,In_449,In_970);
nand U1614 (N_1614,In_267,In_526);
nor U1615 (N_1615,In_897,In_478);
and U1616 (N_1616,In_1474,In_226);
nand U1617 (N_1617,In_283,In_297);
and U1618 (N_1618,In_1263,In_549);
and U1619 (N_1619,In_506,In_1245);
nand U1620 (N_1620,In_107,In_809);
nor U1621 (N_1621,In_234,In_857);
nand U1622 (N_1622,In_1046,In_199);
xnor U1623 (N_1623,In_1305,In_1224);
xor U1624 (N_1624,In_725,In_514);
or U1625 (N_1625,In_1024,In_1191);
nand U1626 (N_1626,In_894,In_1243);
nor U1627 (N_1627,In_739,In_730);
xnor U1628 (N_1628,In_633,In_704);
nor U1629 (N_1629,In_378,In_949);
and U1630 (N_1630,In_355,In_1465);
xnor U1631 (N_1631,In_1259,In_749);
nor U1632 (N_1632,In_1282,In_219);
and U1633 (N_1633,In_131,In_389);
nor U1634 (N_1634,In_628,In_443);
or U1635 (N_1635,In_296,In_1428);
xnor U1636 (N_1636,In_1456,In_541);
nand U1637 (N_1637,In_409,In_1490);
nand U1638 (N_1638,In_1229,In_323);
xnor U1639 (N_1639,In_129,In_1069);
or U1640 (N_1640,In_1230,In_475);
and U1641 (N_1641,In_1088,In_554);
and U1642 (N_1642,In_415,In_873);
or U1643 (N_1643,In_600,In_584);
or U1644 (N_1644,In_1389,In_44);
and U1645 (N_1645,In_1228,In_1452);
or U1646 (N_1646,In_649,In_578);
xor U1647 (N_1647,In_490,In_1236);
nand U1648 (N_1648,In_449,In_578);
nor U1649 (N_1649,In_137,In_985);
and U1650 (N_1650,In_1304,In_1458);
nor U1651 (N_1651,In_1149,In_1498);
nor U1652 (N_1652,In_161,In_720);
or U1653 (N_1653,In_630,In_1371);
or U1654 (N_1654,In_419,In_347);
or U1655 (N_1655,In_1118,In_6);
nand U1656 (N_1656,In_1069,In_952);
xnor U1657 (N_1657,In_1098,In_109);
or U1658 (N_1658,In_859,In_1479);
or U1659 (N_1659,In_1139,In_524);
and U1660 (N_1660,In_50,In_943);
nand U1661 (N_1661,In_1132,In_1352);
nand U1662 (N_1662,In_1481,In_415);
and U1663 (N_1663,In_236,In_1109);
nor U1664 (N_1664,In_774,In_255);
nor U1665 (N_1665,In_1011,In_776);
and U1666 (N_1666,In_1350,In_575);
or U1667 (N_1667,In_909,In_176);
nand U1668 (N_1668,In_712,In_453);
nor U1669 (N_1669,In_1381,In_1324);
and U1670 (N_1670,In_821,In_1135);
nor U1671 (N_1671,In_815,In_454);
nor U1672 (N_1672,In_117,In_981);
nand U1673 (N_1673,In_899,In_671);
and U1674 (N_1674,In_1140,In_1391);
nand U1675 (N_1675,In_196,In_1123);
or U1676 (N_1676,In_821,In_859);
nand U1677 (N_1677,In_1301,In_1045);
and U1678 (N_1678,In_194,In_849);
and U1679 (N_1679,In_526,In_1146);
xor U1680 (N_1680,In_47,In_288);
nor U1681 (N_1681,In_598,In_737);
and U1682 (N_1682,In_1195,In_1155);
or U1683 (N_1683,In_859,In_674);
nand U1684 (N_1684,In_1485,In_1035);
nand U1685 (N_1685,In_814,In_16);
and U1686 (N_1686,In_227,In_282);
nand U1687 (N_1687,In_21,In_639);
or U1688 (N_1688,In_988,In_713);
nand U1689 (N_1689,In_519,In_791);
nor U1690 (N_1690,In_1259,In_836);
xor U1691 (N_1691,In_235,In_1179);
or U1692 (N_1692,In_1211,In_1334);
and U1693 (N_1693,In_1009,In_952);
and U1694 (N_1694,In_280,In_1203);
nor U1695 (N_1695,In_858,In_1397);
and U1696 (N_1696,In_544,In_1419);
or U1697 (N_1697,In_745,In_1144);
or U1698 (N_1698,In_637,In_910);
or U1699 (N_1699,In_454,In_788);
xnor U1700 (N_1700,In_156,In_299);
nor U1701 (N_1701,In_261,In_1002);
nor U1702 (N_1702,In_303,In_391);
or U1703 (N_1703,In_955,In_921);
xor U1704 (N_1704,In_495,In_982);
nand U1705 (N_1705,In_1353,In_753);
xor U1706 (N_1706,In_515,In_1025);
or U1707 (N_1707,In_578,In_182);
or U1708 (N_1708,In_1416,In_582);
nor U1709 (N_1709,In_544,In_433);
xor U1710 (N_1710,In_525,In_956);
nand U1711 (N_1711,In_665,In_93);
nor U1712 (N_1712,In_1370,In_496);
nand U1713 (N_1713,In_640,In_652);
or U1714 (N_1714,In_1026,In_583);
nand U1715 (N_1715,In_624,In_889);
nor U1716 (N_1716,In_812,In_448);
xor U1717 (N_1717,In_991,In_999);
nand U1718 (N_1718,In_1165,In_1187);
or U1719 (N_1719,In_287,In_296);
nor U1720 (N_1720,In_745,In_1401);
nand U1721 (N_1721,In_1446,In_775);
xor U1722 (N_1722,In_849,In_1467);
or U1723 (N_1723,In_743,In_1062);
or U1724 (N_1724,In_250,In_519);
nor U1725 (N_1725,In_929,In_1035);
nor U1726 (N_1726,In_729,In_510);
nand U1727 (N_1727,In_1399,In_1398);
and U1728 (N_1728,In_1250,In_576);
or U1729 (N_1729,In_253,In_1266);
or U1730 (N_1730,In_1145,In_1120);
nand U1731 (N_1731,In_93,In_25);
nor U1732 (N_1732,In_143,In_300);
or U1733 (N_1733,In_857,In_1479);
xnor U1734 (N_1734,In_418,In_72);
nor U1735 (N_1735,In_1214,In_1072);
nor U1736 (N_1736,In_547,In_1020);
and U1737 (N_1737,In_1347,In_626);
nand U1738 (N_1738,In_1481,In_73);
or U1739 (N_1739,In_513,In_850);
and U1740 (N_1740,In_940,In_1382);
nand U1741 (N_1741,In_838,In_1322);
nand U1742 (N_1742,In_19,In_127);
xnor U1743 (N_1743,In_143,In_841);
and U1744 (N_1744,In_560,In_506);
or U1745 (N_1745,In_177,In_451);
nor U1746 (N_1746,In_1417,In_1090);
and U1747 (N_1747,In_162,In_310);
or U1748 (N_1748,In_1059,In_910);
nand U1749 (N_1749,In_24,In_506);
or U1750 (N_1750,In_1423,In_0);
nand U1751 (N_1751,In_957,In_527);
nor U1752 (N_1752,In_908,In_121);
and U1753 (N_1753,In_566,In_1039);
nand U1754 (N_1754,In_311,In_465);
nor U1755 (N_1755,In_1291,In_1126);
and U1756 (N_1756,In_801,In_565);
or U1757 (N_1757,In_941,In_936);
nand U1758 (N_1758,In_1313,In_858);
or U1759 (N_1759,In_307,In_61);
xor U1760 (N_1760,In_1155,In_1033);
or U1761 (N_1761,In_444,In_329);
or U1762 (N_1762,In_179,In_174);
or U1763 (N_1763,In_1040,In_585);
nand U1764 (N_1764,In_285,In_1395);
nor U1765 (N_1765,In_1494,In_201);
xnor U1766 (N_1766,In_414,In_312);
or U1767 (N_1767,In_613,In_435);
or U1768 (N_1768,In_845,In_1097);
nand U1769 (N_1769,In_983,In_667);
or U1770 (N_1770,In_283,In_849);
xnor U1771 (N_1771,In_404,In_543);
and U1772 (N_1772,In_724,In_1355);
nor U1773 (N_1773,In_237,In_298);
and U1774 (N_1774,In_751,In_322);
xnor U1775 (N_1775,In_862,In_1346);
xor U1776 (N_1776,In_637,In_576);
or U1777 (N_1777,In_1025,In_276);
nor U1778 (N_1778,In_1181,In_1005);
nor U1779 (N_1779,In_708,In_467);
nand U1780 (N_1780,In_1024,In_1084);
xor U1781 (N_1781,In_564,In_998);
nand U1782 (N_1782,In_691,In_737);
nand U1783 (N_1783,In_1214,In_954);
nor U1784 (N_1784,In_39,In_266);
or U1785 (N_1785,In_344,In_511);
and U1786 (N_1786,In_71,In_1475);
or U1787 (N_1787,In_1113,In_181);
or U1788 (N_1788,In_613,In_547);
xnor U1789 (N_1789,In_969,In_1167);
nand U1790 (N_1790,In_1460,In_1328);
nand U1791 (N_1791,In_213,In_916);
and U1792 (N_1792,In_682,In_708);
nor U1793 (N_1793,In_895,In_478);
xor U1794 (N_1794,In_193,In_577);
and U1795 (N_1795,In_769,In_41);
nor U1796 (N_1796,In_499,In_978);
nand U1797 (N_1797,In_1331,In_1147);
or U1798 (N_1798,In_131,In_1037);
or U1799 (N_1799,In_882,In_181);
xnor U1800 (N_1800,In_44,In_471);
xor U1801 (N_1801,In_142,In_431);
and U1802 (N_1802,In_160,In_98);
nor U1803 (N_1803,In_1256,In_1376);
nand U1804 (N_1804,In_1195,In_395);
or U1805 (N_1805,In_365,In_190);
or U1806 (N_1806,In_646,In_1436);
nand U1807 (N_1807,In_827,In_867);
and U1808 (N_1808,In_863,In_1123);
nand U1809 (N_1809,In_1438,In_1209);
nor U1810 (N_1810,In_1495,In_293);
or U1811 (N_1811,In_545,In_758);
or U1812 (N_1812,In_1497,In_1416);
or U1813 (N_1813,In_1053,In_1366);
and U1814 (N_1814,In_811,In_859);
or U1815 (N_1815,In_1490,In_798);
nor U1816 (N_1816,In_919,In_1084);
or U1817 (N_1817,In_1062,In_921);
nand U1818 (N_1818,In_519,In_1369);
nor U1819 (N_1819,In_1144,In_391);
nor U1820 (N_1820,In_1227,In_285);
xor U1821 (N_1821,In_1091,In_758);
xor U1822 (N_1822,In_926,In_1161);
and U1823 (N_1823,In_955,In_894);
and U1824 (N_1824,In_199,In_468);
nand U1825 (N_1825,In_1219,In_492);
nor U1826 (N_1826,In_731,In_235);
or U1827 (N_1827,In_1285,In_186);
or U1828 (N_1828,In_925,In_63);
xor U1829 (N_1829,In_1156,In_581);
or U1830 (N_1830,In_483,In_1335);
nand U1831 (N_1831,In_222,In_1384);
xor U1832 (N_1832,In_928,In_290);
nand U1833 (N_1833,In_1087,In_1261);
nor U1834 (N_1834,In_611,In_487);
nand U1835 (N_1835,In_704,In_1257);
xor U1836 (N_1836,In_233,In_906);
and U1837 (N_1837,In_1324,In_1406);
nand U1838 (N_1838,In_78,In_626);
and U1839 (N_1839,In_888,In_238);
or U1840 (N_1840,In_579,In_1177);
and U1841 (N_1841,In_1042,In_1303);
nor U1842 (N_1842,In_542,In_782);
or U1843 (N_1843,In_1073,In_819);
nand U1844 (N_1844,In_880,In_764);
nor U1845 (N_1845,In_1234,In_1492);
and U1846 (N_1846,In_1480,In_1316);
xnor U1847 (N_1847,In_44,In_353);
or U1848 (N_1848,In_796,In_669);
or U1849 (N_1849,In_1477,In_1415);
and U1850 (N_1850,In_1399,In_1045);
xnor U1851 (N_1851,In_1472,In_917);
or U1852 (N_1852,In_448,In_824);
nor U1853 (N_1853,In_495,In_265);
nor U1854 (N_1854,In_1119,In_335);
nand U1855 (N_1855,In_740,In_281);
nand U1856 (N_1856,In_1141,In_912);
or U1857 (N_1857,In_212,In_1028);
nand U1858 (N_1858,In_1098,In_383);
and U1859 (N_1859,In_573,In_1332);
or U1860 (N_1860,In_1096,In_1125);
and U1861 (N_1861,In_478,In_1115);
and U1862 (N_1862,In_1495,In_269);
nand U1863 (N_1863,In_120,In_884);
and U1864 (N_1864,In_1256,In_895);
or U1865 (N_1865,In_205,In_977);
nand U1866 (N_1866,In_45,In_21);
nor U1867 (N_1867,In_431,In_125);
or U1868 (N_1868,In_1083,In_1335);
or U1869 (N_1869,In_64,In_192);
nand U1870 (N_1870,In_1158,In_671);
nand U1871 (N_1871,In_487,In_643);
and U1872 (N_1872,In_248,In_1338);
nand U1873 (N_1873,In_687,In_67);
xnor U1874 (N_1874,In_92,In_366);
or U1875 (N_1875,In_1446,In_483);
nor U1876 (N_1876,In_1413,In_190);
or U1877 (N_1877,In_183,In_385);
nand U1878 (N_1878,In_87,In_1012);
and U1879 (N_1879,In_1295,In_798);
nand U1880 (N_1880,In_635,In_1224);
nor U1881 (N_1881,In_1075,In_625);
nand U1882 (N_1882,In_6,In_1290);
nand U1883 (N_1883,In_699,In_1446);
nor U1884 (N_1884,In_103,In_1472);
xor U1885 (N_1885,In_817,In_33);
nor U1886 (N_1886,In_648,In_858);
nor U1887 (N_1887,In_1240,In_163);
or U1888 (N_1888,In_651,In_422);
xnor U1889 (N_1889,In_1341,In_941);
or U1890 (N_1890,In_445,In_514);
or U1891 (N_1891,In_995,In_379);
xor U1892 (N_1892,In_1296,In_364);
or U1893 (N_1893,In_1483,In_1290);
nor U1894 (N_1894,In_79,In_1486);
nand U1895 (N_1895,In_300,In_591);
xnor U1896 (N_1896,In_255,In_1036);
and U1897 (N_1897,In_1270,In_1109);
or U1898 (N_1898,In_575,In_648);
xor U1899 (N_1899,In_1119,In_482);
nor U1900 (N_1900,In_1364,In_737);
and U1901 (N_1901,In_444,In_818);
nand U1902 (N_1902,In_957,In_772);
xnor U1903 (N_1903,In_343,In_723);
and U1904 (N_1904,In_35,In_318);
nand U1905 (N_1905,In_1053,In_54);
or U1906 (N_1906,In_393,In_1181);
nand U1907 (N_1907,In_112,In_1322);
and U1908 (N_1908,In_728,In_286);
xor U1909 (N_1909,In_745,In_548);
nor U1910 (N_1910,In_632,In_680);
nor U1911 (N_1911,In_105,In_455);
and U1912 (N_1912,In_901,In_1268);
xnor U1913 (N_1913,In_1278,In_1309);
or U1914 (N_1914,In_152,In_422);
or U1915 (N_1915,In_564,In_262);
nand U1916 (N_1916,In_1107,In_98);
and U1917 (N_1917,In_817,In_1310);
nand U1918 (N_1918,In_515,In_1414);
and U1919 (N_1919,In_749,In_861);
or U1920 (N_1920,In_541,In_213);
nor U1921 (N_1921,In_864,In_214);
nor U1922 (N_1922,In_1087,In_507);
and U1923 (N_1923,In_1018,In_895);
nor U1924 (N_1924,In_748,In_269);
nand U1925 (N_1925,In_1468,In_1115);
nand U1926 (N_1926,In_175,In_1335);
or U1927 (N_1927,In_278,In_1436);
nor U1928 (N_1928,In_1288,In_903);
nor U1929 (N_1929,In_1371,In_727);
and U1930 (N_1930,In_680,In_574);
nand U1931 (N_1931,In_754,In_1480);
nand U1932 (N_1932,In_1084,In_1206);
nor U1933 (N_1933,In_124,In_1385);
nand U1934 (N_1934,In_1411,In_643);
nor U1935 (N_1935,In_268,In_577);
and U1936 (N_1936,In_904,In_645);
nand U1937 (N_1937,In_179,In_15);
nand U1938 (N_1938,In_254,In_1000);
nor U1939 (N_1939,In_466,In_723);
nor U1940 (N_1940,In_1433,In_1290);
nor U1941 (N_1941,In_442,In_975);
nor U1942 (N_1942,In_771,In_1101);
nand U1943 (N_1943,In_396,In_503);
nand U1944 (N_1944,In_688,In_536);
and U1945 (N_1945,In_3,In_260);
nor U1946 (N_1946,In_138,In_334);
nand U1947 (N_1947,In_1332,In_157);
nand U1948 (N_1948,In_1317,In_804);
nor U1949 (N_1949,In_865,In_1322);
nor U1950 (N_1950,In_1028,In_1322);
and U1951 (N_1951,In_473,In_968);
nand U1952 (N_1952,In_1170,In_293);
nor U1953 (N_1953,In_515,In_493);
nand U1954 (N_1954,In_665,In_1404);
nor U1955 (N_1955,In_172,In_272);
xor U1956 (N_1956,In_810,In_52);
and U1957 (N_1957,In_1385,In_1383);
xor U1958 (N_1958,In_1130,In_805);
or U1959 (N_1959,In_1404,In_1328);
and U1960 (N_1960,In_1375,In_1016);
or U1961 (N_1961,In_350,In_991);
and U1962 (N_1962,In_202,In_654);
or U1963 (N_1963,In_517,In_1136);
and U1964 (N_1964,In_139,In_541);
or U1965 (N_1965,In_1120,In_1368);
and U1966 (N_1966,In_291,In_1202);
xor U1967 (N_1967,In_575,In_482);
and U1968 (N_1968,In_785,In_398);
or U1969 (N_1969,In_1352,In_1166);
nand U1970 (N_1970,In_53,In_831);
or U1971 (N_1971,In_1489,In_642);
or U1972 (N_1972,In_1278,In_310);
nand U1973 (N_1973,In_143,In_158);
nor U1974 (N_1974,In_1101,In_703);
nor U1975 (N_1975,In_1360,In_264);
nor U1976 (N_1976,In_852,In_774);
nor U1977 (N_1977,In_1249,In_1232);
nand U1978 (N_1978,In_1301,In_1373);
nor U1979 (N_1979,In_1145,In_567);
and U1980 (N_1980,In_1213,In_1013);
and U1981 (N_1981,In_214,In_1365);
and U1982 (N_1982,In_1324,In_184);
or U1983 (N_1983,In_571,In_547);
nand U1984 (N_1984,In_298,In_1466);
nor U1985 (N_1985,In_1143,In_336);
or U1986 (N_1986,In_738,In_242);
nand U1987 (N_1987,In_440,In_997);
nand U1988 (N_1988,In_377,In_1350);
nor U1989 (N_1989,In_184,In_309);
nor U1990 (N_1990,In_1253,In_1125);
or U1991 (N_1991,In_178,In_1394);
and U1992 (N_1992,In_1006,In_795);
nand U1993 (N_1993,In_988,In_1403);
or U1994 (N_1994,In_437,In_829);
xnor U1995 (N_1995,In_230,In_1413);
nor U1996 (N_1996,In_390,In_964);
nor U1997 (N_1997,In_175,In_874);
or U1998 (N_1998,In_889,In_1139);
nor U1999 (N_1999,In_341,In_416);
and U2000 (N_2000,In_564,In_123);
or U2001 (N_2001,In_421,In_1093);
and U2002 (N_2002,In_647,In_470);
and U2003 (N_2003,In_832,In_1333);
nor U2004 (N_2004,In_47,In_320);
and U2005 (N_2005,In_1190,In_447);
and U2006 (N_2006,In_802,In_941);
xnor U2007 (N_2007,In_0,In_1289);
nand U2008 (N_2008,In_1235,In_1181);
and U2009 (N_2009,In_54,In_217);
xor U2010 (N_2010,In_174,In_1089);
or U2011 (N_2011,In_1457,In_51);
nor U2012 (N_2012,In_1168,In_1278);
nand U2013 (N_2013,In_816,In_1270);
or U2014 (N_2014,In_1288,In_706);
nand U2015 (N_2015,In_912,In_212);
and U2016 (N_2016,In_112,In_170);
or U2017 (N_2017,In_411,In_71);
and U2018 (N_2018,In_310,In_610);
xnor U2019 (N_2019,In_581,In_106);
nor U2020 (N_2020,In_228,In_1315);
and U2021 (N_2021,In_594,In_162);
nand U2022 (N_2022,In_750,In_1052);
or U2023 (N_2023,In_1290,In_281);
nor U2024 (N_2024,In_1189,In_1201);
nand U2025 (N_2025,In_778,In_372);
or U2026 (N_2026,In_1140,In_978);
or U2027 (N_2027,In_1321,In_882);
xnor U2028 (N_2028,In_738,In_188);
or U2029 (N_2029,In_168,In_1387);
and U2030 (N_2030,In_1319,In_273);
or U2031 (N_2031,In_917,In_1209);
xnor U2032 (N_2032,In_1040,In_1449);
xor U2033 (N_2033,In_1141,In_63);
and U2034 (N_2034,In_1253,In_652);
nor U2035 (N_2035,In_378,In_470);
nor U2036 (N_2036,In_1290,In_579);
nand U2037 (N_2037,In_844,In_613);
nor U2038 (N_2038,In_545,In_708);
nand U2039 (N_2039,In_515,In_477);
nand U2040 (N_2040,In_1449,In_1114);
xor U2041 (N_2041,In_1171,In_1375);
nor U2042 (N_2042,In_112,In_436);
and U2043 (N_2043,In_96,In_879);
and U2044 (N_2044,In_71,In_566);
and U2045 (N_2045,In_405,In_822);
nor U2046 (N_2046,In_1101,In_1363);
and U2047 (N_2047,In_354,In_349);
nor U2048 (N_2048,In_1486,In_1276);
nand U2049 (N_2049,In_9,In_1178);
nor U2050 (N_2050,In_1404,In_587);
nor U2051 (N_2051,In_318,In_911);
nor U2052 (N_2052,In_436,In_789);
nor U2053 (N_2053,In_805,In_1186);
nand U2054 (N_2054,In_1068,In_1403);
and U2055 (N_2055,In_551,In_1253);
nor U2056 (N_2056,In_925,In_721);
nor U2057 (N_2057,In_828,In_480);
nand U2058 (N_2058,In_409,In_498);
or U2059 (N_2059,In_910,In_1138);
and U2060 (N_2060,In_1282,In_452);
xnor U2061 (N_2061,In_1468,In_1016);
nand U2062 (N_2062,In_227,In_751);
and U2063 (N_2063,In_252,In_1229);
and U2064 (N_2064,In_586,In_640);
nor U2065 (N_2065,In_1020,In_1126);
or U2066 (N_2066,In_1303,In_959);
and U2067 (N_2067,In_808,In_24);
nor U2068 (N_2068,In_836,In_508);
and U2069 (N_2069,In_898,In_1338);
and U2070 (N_2070,In_1181,In_937);
and U2071 (N_2071,In_434,In_1326);
nor U2072 (N_2072,In_1384,In_1177);
and U2073 (N_2073,In_1138,In_215);
or U2074 (N_2074,In_967,In_395);
nand U2075 (N_2075,In_685,In_670);
nand U2076 (N_2076,In_901,In_902);
nand U2077 (N_2077,In_50,In_868);
nand U2078 (N_2078,In_1398,In_43);
nor U2079 (N_2079,In_901,In_278);
or U2080 (N_2080,In_291,In_1025);
and U2081 (N_2081,In_65,In_312);
nand U2082 (N_2082,In_237,In_1119);
nor U2083 (N_2083,In_713,In_690);
xor U2084 (N_2084,In_664,In_463);
nor U2085 (N_2085,In_771,In_496);
and U2086 (N_2086,In_1254,In_742);
nand U2087 (N_2087,In_851,In_885);
and U2088 (N_2088,In_1152,In_906);
nand U2089 (N_2089,In_174,In_1499);
nand U2090 (N_2090,In_79,In_327);
or U2091 (N_2091,In_772,In_173);
nor U2092 (N_2092,In_1072,In_1195);
or U2093 (N_2093,In_893,In_89);
nand U2094 (N_2094,In_386,In_990);
nor U2095 (N_2095,In_526,In_885);
and U2096 (N_2096,In_1093,In_709);
xnor U2097 (N_2097,In_61,In_1017);
nand U2098 (N_2098,In_1206,In_1168);
nor U2099 (N_2099,In_135,In_662);
or U2100 (N_2100,In_609,In_1483);
and U2101 (N_2101,In_751,In_1300);
and U2102 (N_2102,In_1356,In_1212);
nand U2103 (N_2103,In_1087,In_1177);
or U2104 (N_2104,In_626,In_386);
nand U2105 (N_2105,In_510,In_439);
nor U2106 (N_2106,In_49,In_1126);
nor U2107 (N_2107,In_1090,In_257);
and U2108 (N_2108,In_498,In_82);
nand U2109 (N_2109,In_116,In_1241);
nor U2110 (N_2110,In_1354,In_1010);
nor U2111 (N_2111,In_848,In_381);
and U2112 (N_2112,In_689,In_638);
and U2113 (N_2113,In_1331,In_1129);
nand U2114 (N_2114,In_649,In_81);
or U2115 (N_2115,In_1176,In_614);
nand U2116 (N_2116,In_30,In_1412);
nand U2117 (N_2117,In_872,In_939);
xnor U2118 (N_2118,In_1003,In_90);
and U2119 (N_2119,In_761,In_1296);
nor U2120 (N_2120,In_955,In_502);
nor U2121 (N_2121,In_1258,In_1488);
nor U2122 (N_2122,In_1418,In_761);
nor U2123 (N_2123,In_312,In_1316);
nand U2124 (N_2124,In_1270,In_181);
nand U2125 (N_2125,In_1177,In_796);
nor U2126 (N_2126,In_852,In_551);
nand U2127 (N_2127,In_1074,In_13);
or U2128 (N_2128,In_1402,In_1480);
and U2129 (N_2129,In_1007,In_1069);
or U2130 (N_2130,In_885,In_1008);
nand U2131 (N_2131,In_808,In_67);
and U2132 (N_2132,In_523,In_682);
and U2133 (N_2133,In_869,In_916);
and U2134 (N_2134,In_1005,In_1400);
nor U2135 (N_2135,In_475,In_1038);
nor U2136 (N_2136,In_327,In_333);
and U2137 (N_2137,In_210,In_731);
and U2138 (N_2138,In_45,In_727);
nand U2139 (N_2139,In_622,In_1472);
nor U2140 (N_2140,In_828,In_939);
nand U2141 (N_2141,In_253,In_620);
nand U2142 (N_2142,In_935,In_992);
xor U2143 (N_2143,In_1437,In_1251);
nand U2144 (N_2144,In_1037,In_1192);
nand U2145 (N_2145,In_128,In_694);
or U2146 (N_2146,In_592,In_1444);
nand U2147 (N_2147,In_1391,In_413);
nor U2148 (N_2148,In_1443,In_769);
nor U2149 (N_2149,In_917,In_573);
nand U2150 (N_2150,In_546,In_1118);
or U2151 (N_2151,In_774,In_613);
nor U2152 (N_2152,In_426,In_387);
and U2153 (N_2153,In_954,In_274);
and U2154 (N_2154,In_515,In_137);
and U2155 (N_2155,In_979,In_980);
or U2156 (N_2156,In_1384,In_88);
nand U2157 (N_2157,In_986,In_664);
or U2158 (N_2158,In_601,In_754);
or U2159 (N_2159,In_898,In_48);
xor U2160 (N_2160,In_1032,In_113);
and U2161 (N_2161,In_823,In_445);
nand U2162 (N_2162,In_83,In_503);
nor U2163 (N_2163,In_505,In_428);
xor U2164 (N_2164,In_1024,In_341);
nand U2165 (N_2165,In_1024,In_1437);
nand U2166 (N_2166,In_1209,In_1284);
or U2167 (N_2167,In_603,In_268);
or U2168 (N_2168,In_1204,In_165);
nand U2169 (N_2169,In_302,In_452);
xnor U2170 (N_2170,In_240,In_4);
xor U2171 (N_2171,In_782,In_816);
xnor U2172 (N_2172,In_1103,In_1010);
and U2173 (N_2173,In_1134,In_892);
xor U2174 (N_2174,In_1430,In_30);
xnor U2175 (N_2175,In_263,In_1437);
nor U2176 (N_2176,In_848,In_605);
or U2177 (N_2177,In_1369,In_444);
nand U2178 (N_2178,In_1313,In_738);
and U2179 (N_2179,In_1161,In_1458);
and U2180 (N_2180,In_603,In_1398);
nor U2181 (N_2181,In_515,In_1118);
and U2182 (N_2182,In_308,In_852);
nor U2183 (N_2183,In_217,In_594);
nor U2184 (N_2184,In_805,In_488);
or U2185 (N_2185,In_1299,In_1389);
nand U2186 (N_2186,In_798,In_239);
nand U2187 (N_2187,In_700,In_559);
nand U2188 (N_2188,In_669,In_23);
nand U2189 (N_2189,In_1083,In_214);
xor U2190 (N_2190,In_822,In_1420);
nand U2191 (N_2191,In_1411,In_494);
nor U2192 (N_2192,In_287,In_1400);
nand U2193 (N_2193,In_246,In_70);
nor U2194 (N_2194,In_1108,In_1170);
and U2195 (N_2195,In_1335,In_956);
xnor U2196 (N_2196,In_448,In_279);
nand U2197 (N_2197,In_74,In_457);
or U2198 (N_2198,In_1155,In_908);
nor U2199 (N_2199,In_551,In_310);
nand U2200 (N_2200,In_1175,In_29);
nand U2201 (N_2201,In_1210,In_263);
nand U2202 (N_2202,In_664,In_1381);
and U2203 (N_2203,In_1030,In_720);
and U2204 (N_2204,In_117,In_182);
or U2205 (N_2205,In_356,In_1124);
nor U2206 (N_2206,In_548,In_677);
and U2207 (N_2207,In_830,In_11);
nand U2208 (N_2208,In_401,In_130);
xor U2209 (N_2209,In_111,In_1481);
or U2210 (N_2210,In_505,In_1402);
or U2211 (N_2211,In_757,In_457);
or U2212 (N_2212,In_1007,In_849);
nand U2213 (N_2213,In_939,In_561);
nor U2214 (N_2214,In_853,In_85);
xnor U2215 (N_2215,In_153,In_77);
or U2216 (N_2216,In_886,In_494);
and U2217 (N_2217,In_1015,In_936);
nor U2218 (N_2218,In_469,In_1369);
and U2219 (N_2219,In_31,In_1103);
nand U2220 (N_2220,In_138,In_1493);
and U2221 (N_2221,In_290,In_731);
nor U2222 (N_2222,In_50,In_670);
nor U2223 (N_2223,In_1312,In_599);
nand U2224 (N_2224,In_902,In_437);
and U2225 (N_2225,In_257,In_1490);
and U2226 (N_2226,In_1070,In_701);
or U2227 (N_2227,In_742,In_543);
and U2228 (N_2228,In_532,In_141);
or U2229 (N_2229,In_515,In_1395);
or U2230 (N_2230,In_309,In_714);
nand U2231 (N_2231,In_173,In_327);
nor U2232 (N_2232,In_379,In_1465);
nand U2233 (N_2233,In_1057,In_1107);
nand U2234 (N_2234,In_460,In_508);
nor U2235 (N_2235,In_286,In_419);
nand U2236 (N_2236,In_875,In_1223);
nand U2237 (N_2237,In_872,In_1467);
and U2238 (N_2238,In_1128,In_69);
nand U2239 (N_2239,In_381,In_71);
nand U2240 (N_2240,In_158,In_589);
nand U2241 (N_2241,In_1187,In_53);
nor U2242 (N_2242,In_192,In_1015);
and U2243 (N_2243,In_726,In_1488);
or U2244 (N_2244,In_742,In_739);
nor U2245 (N_2245,In_510,In_396);
nor U2246 (N_2246,In_1235,In_692);
nor U2247 (N_2247,In_1485,In_896);
nor U2248 (N_2248,In_724,In_925);
xnor U2249 (N_2249,In_980,In_427);
nor U2250 (N_2250,In_674,In_603);
or U2251 (N_2251,In_1014,In_553);
nor U2252 (N_2252,In_516,In_154);
or U2253 (N_2253,In_1059,In_532);
nand U2254 (N_2254,In_816,In_33);
nand U2255 (N_2255,In_964,In_883);
and U2256 (N_2256,In_958,In_981);
nand U2257 (N_2257,In_1087,In_1026);
or U2258 (N_2258,In_851,In_1401);
xor U2259 (N_2259,In_1216,In_1158);
or U2260 (N_2260,In_945,In_1289);
nor U2261 (N_2261,In_902,In_365);
and U2262 (N_2262,In_1351,In_1399);
xnor U2263 (N_2263,In_214,In_56);
nand U2264 (N_2264,In_611,In_1420);
nand U2265 (N_2265,In_451,In_636);
or U2266 (N_2266,In_1478,In_166);
nand U2267 (N_2267,In_1188,In_95);
nand U2268 (N_2268,In_1057,In_1022);
nor U2269 (N_2269,In_1241,In_977);
and U2270 (N_2270,In_1298,In_132);
xor U2271 (N_2271,In_1426,In_6);
nand U2272 (N_2272,In_1343,In_467);
or U2273 (N_2273,In_179,In_135);
or U2274 (N_2274,In_727,In_1393);
nand U2275 (N_2275,In_254,In_1431);
and U2276 (N_2276,In_494,In_420);
and U2277 (N_2277,In_350,In_923);
nand U2278 (N_2278,In_1208,In_1472);
nand U2279 (N_2279,In_49,In_349);
nor U2280 (N_2280,In_136,In_1252);
nor U2281 (N_2281,In_629,In_1269);
nor U2282 (N_2282,In_1218,In_1213);
and U2283 (N_2283,In_699,In_1152);
or U2284 (N_2284,In_1155,In_1200);
or U2285 (N_2285,In_1487,In_500);
nand U2286 (N_2286,In_656,In_619);
nand U2287 (N_2287,In_279,In_593);
and U2288 (N_2288,In_290,In_1058);
or U2289 (N_2289,In_71,In_377);
nand U2290 (N_2290,In_1062,In_1077);
and U2291 (N_2291,In_323,In_518);
nor U2292 (N_2292,In_255,In_1154);
nand U2293 (N_2293,In_1092,In_1021);
nor U2294 (N_2294,In_1178,In_241);
or U2295 (N_2295,In_287,In_220);
and U2296 (N_2296,In_469,In_950);
xnor U2297 (N_2297,In_522,In_241);
nand U2298 (N_2298,In_519,In_1055);
nand U2299 (N_2299,In_1484,In_267);
xor U2300 (N_2300,In_196,In_517);
and U2301 (N_2301,In_983,In_513);
xnor U2302 (N_2302,In_823,In_607);
nand U2303 (N_2303,In_465,In_803);
nor U2304 (N_2304,In_1497,In_1143);
nand U2305 (N_2305,In_1430,In_760);
or U2306 (N_2306,In_185,In_210);
and U2307 (N_2307,In_531,In_648);
xor U2308 (N_2308,In_776,In_851);
and U2309 (N_2309,In_584,In_705);
nor U2310 (N_2310,In_193,In_1261);
xor U2311 (N_2311,In_93,In_498);
nor U2312 (N_2312,In_29,In_418);
nor U2313 (N_2313,In_591,In_78);
or U2314 (N_2314,In_1416,In_1271);
nand U2315 (N_2315,In_27,In_881);
xnor U2316 (N_2316,In_1086,In_1435);
nor U2317 (N_2317,In_487,In_1341);
and U2318 (N_2318,In_840,In_718);
nor U2319 (N_2319,In_702,In_325);
nor U2320 (N_2320,In_78,In_351);
xnor U2321 (N_2321,In_443,In_286);
xnor U2322 (N_2322,In_743,In_1071);
nand U2323 (N_2323,In_742,In_228);
and U2324 (N_2324,In_668,In_1498);
and U2325 (N_2325,In_148,In_1249);
and U2326 (N_2326,In_1254,In_33);
nand U2327 (N_2327,In_209,In_1146);
or U2328 (N_2328,In_706,In_801);
nand U2329 (N_2329,In_401,In_379);
or U2330 (N_2330,In_1198,In_725);
or U2331 (N_2331,In_1076,In_45);
and U2332 (N_2332,In_1344,In_593);
or U2333 (N_2333,In_1016,In_308);
nor U2334 (N_2334,In_226,In_370);
nand U2335 (N_2335,In_757,In_805);
nand U2336 (N_2336,In_190,In_866);
and U2337 (N_2337,In_873,In_426);
nand U2338 (N_2338,In_703,In_783);
and U2339 (N_2339,In_796,In_1309);
or U2340 (N_2340,In_881,In_777);
or U2341 (N_2341,In_918,In_1299);
nand U2342 (N_2342,In_622,In_665);
xnor U2343 (N_2343,In_24,In_200);
or U2344 (N_2344,In_623,In_395);
nor U2345 (N_2345,In_1318,In_1203);
xor U2346 (N_2346,In_1135,In_1126);
nor U2347 (N_2347,In_1247,In_1256);
nand U2348 (N_2348,In_1472,In_43);
or U2349 (N_2349,In_344,In_395);
or U2350 (N_2350,In_774,In_487);
or U2351 (N_2351,In_134,In_1270);
or U2352 (N_2352,In_601,In_850);
and U2353 (N_2353,In_1196,In_1077);
or U2354 (N_2354,In_154,In_631);
nor U2355 (N_2355,In_1309,In_567);
and U2356 (N_2356,In_506,In_174);
nor U2357 (N_2357,In_858,In_1069);
or U2358 (N_2358,In_1008,In_1253);
nor U2359 (N_2359,In_654,In_701);
and U2360 (N_2360,In_229,In_1044);
xor U2361 (N_2361,In_32,In_774);
nor U2362 (N_2362,In_121,In_1225);
nand U2363 (N_2363,In_945,In_1128);
and U2364 (N_2364,In_100,In_535);
and U2365 (N_2365,In_1363,In_192);
nor U2366 (N_2366,In_932,In_1188);
xnor U2367 (N_2367,In_433,In_596);
nand U2368 (N_2368,In_827,In_1444);
nor U2369 (N_2369,In_1068,In_577);
or U2370 (N_2370,In_615,In_692);
and U2371 (N_2371,In_430,In_279);
and U2372 (N_2372,In_382,In_253);
nand U2373 (N_2373,In_541,In_1112);
and U2374 (N_2374,In_1176,In_335);
nand U2375 (N_2375,In_1025,In_423);
or U2376 (N_2376,In_43,In_933);
nand U2377 (N_2377,In_573,In_207);
or U2378 (N_2378,In_861,In_1046);
nor U2379 (N_2379,In_1026,In_1333);
or U2380 (N_2380,In_1050,In_920);
and U2381 (N_2381,In_232,In_482);
and U2382 (N_2382,In_952,In_1383);
or U2383 (N_2383,In_33,In_1460);
nor U2384 (N_2384,In_267,In_568);
and U2385 (N_2385,In_979,In_379);
or U2386 (N_2386,In_1042,In_1366);
nand U2387 (N_2387,In_1289,In_1310);
xnor U2388 (N_2388,In_85,In_1368);
nand U2389 (N_2389,In_6,In_595);
and U2390 (N_2390,In_155,In_1258);
xnor U2391 (N_2391,In_308,In_273);
or U2392 (N_2392,In_179,In_238);
nand U2393 (N_2393,In_461,In_404);
xnor U2394 (N_2394,In_39,In_131);
or U2395 (N_2395,In_784,In_903);
nor U2396 (N_2396,In_476,In_702);
and U2397 (N_2397,In_300,In_86);
nor U2398 (N_2398,In_483,In_231);
nand U2399 (N_2399,In_1439,In_678);
nor U2400 (N_2400,In_1147,In_82);
and U2401 (N_2401,In_593,In_1321);
nand U2402 (N_2402,In_198,In_1214);
nand U2403 (N_2403,In_641,In_827);
and U2404 (N_2404,In_1189,In_181);
and U2405 (N_2405,In_702,In_481);
nand U2406 (N_2406,In_540,In_880);
or U2407 (N_2407,In_36,In_666);
nor U2408 (N_2408,In_876,In_739);
or U2409 (N_2409,In_4,In_377);
and U2410 (N_2410,In_543,In_754);
or U2411 (N_2411,In_811,In_1345);
and U2412 (N_2412,In_421,In_1494);
nor U2413 (N_2413,In_829,In_927);
and U2414 (N_2414,In_350,In_1482);
and U2415 (N_2415,In_312,In_671);
nand U2416 (N_2416,In_1443,In_470);
and U2417 (N_2417,In_1153,In_980);
and U2418 (N_2418,In_356,In_1242);
nand U2419 (N_2419,In_1254,In_189);
and U2420 (N_2420,In_1318,In_938);
nor U2421 (N_2421,In_313,In_270);
or U2422 (N_2422,In_163,In_1040);
nor U2423 (N_2423,In_426,In_631);
nor U2424 (N_2424,In_769,In_432);
nand U2425 (N_2425,In_405,In_806);
or U2426 (N_2426,In_168,In_908);
xnor U2427 (N_2427,In_362,In_545);
and U2428 (N_2428,In_283,In_1287);
nand U2429 (N_2429,In_626,In_505);
or U2430 (N_2430,In_358,In_611);
or U2431 (N_2431,In_994,In_855);
or U2432 (N_2432,In_431,In_483);
and U2433 (N_2433,In_762,In_500);
and U2434 (N_2434,In_267,In_737);
nor U2435 (N_2435,In_959,In_603);
and U2436 (N_2436,In_218,In_1275);
xnor U2437 (N_2437,In_654,In_880);
or U2438 (N_2438,In_616,In_993);
and U2439 (N_2439,In_636,In_325);
or U2440 (N_2440,In_280,In_528);
and U2441 (N_2441,In_1396,In_814);
nor U2442 (N_2442,In_936,In_669);
and U2443 (N_2443,In_67,In_1468);
and U2444 (N_2444,In_1447,In_997);
nand U2445 (N_2445,In_494,In_136);
nor U2446 (N_2446,In_1307,In_1276);
nor U2447 (N_2447,In_338,In_798);
and U2448 (N_2448,In_991,In_224);
nand U2449 (N_2449,In_574,In_73);
nand U2450 (N_2450,In_860,In_582);
or U2451 (N_2451,In_1180,In_1155);
nor U2452 (N_2452,In_827,In_900);
and U2453 (N_2453,In_1493,In_191);
nor U2454 (N_2454,In_1356,In_1407);
or U2455 (N_2455,In_463,In_307);
or U2456 (N_2456,In_1199,In_1423);
nand U2457 (N_2457,In_248,In_254);
nand U2458 (N_2458,In_1103,In_762);
xor U2459 (N_2459,In_442,In_1282);
and U2460 (N_2460,In_904,In_1454);
xor U2461 (N_2461,In_482,In_1252);
nand U2462 (N_2462,In_1133,In_1388);
nand U2463 (N_2463,In_574,In_348);
xor U2464 (N_2464,In_1465,In_1466);
nor U2465 (N_2465,In_399,In_4);
xor U2466 (N_2466,In_269,In_821);
or U2467 (N_2467,In_358,In_1262);
xnor U2468 (N_2468,In_1178,In_709);
or U2469 (N_2469,In_644,In_423);
and U2470 (N_2470,In_1402,In_519);
or U2471 (N_2471,In_1102,In_133);
or U2472 (N_2472,In_143,In_1482);
nor U2473 (N_2473,In_1259,In_1215);
xor U2474 (N_2474,In_945,In_729);
or U2475 (N_2475,In_796,In_651);
or U2476 (N_2476,In_292,In_1302);
nor U2477 (N_2477,In_515,In_1403);
nand U2478 (N_2478,In_572,In_1257);
xnor U2479 (N_2479,In_1189,In_1343);
nor U2480 (N_2480,In_74,In_43);
and U2481 (N_2481,In_1286,In_846);
and U2482 (N_2482,In_498,In_816);
and U2483 (N_2483,In_686,In_249);
xnor U2484 (N_2484,In_1403,In_1459);
or U2485 (N_2485,In_1234,In_386);
and U2486 (N_2486,In_392,In_1175);
or U2487 (N_2487,In_560,In_228);
nand U2488 (N_2488,In_545,In_1479);
nor U2489 (N_2489,In_978,In_367);
nor U2490 (N_2490,In_1109,In_225);
or U2491 (N_2491,In_818,In_684);
and U2492 (N_2492,In_60,In_1187);
or U2493 (N_2493,In_503,In_1371);
nor U2494 (N_2494,In_1433,In_1387);
or U2495 (N_2495,In_1365,In_1108);
nand U2496 (N_2496,In_1347,In_119);
nor U2497 (N_2497,In_696,In_1369);
xor U2498 (N_2498,In_140,In_532);
or U2499 (N_2499,In_1442,In_147);
nand U2500 (N_2500,In_1294,In_728);
nor U2501 (N_2501,In_760,In_992);
and U2502 (N_2502,In_1484,In_1148);
or U2503 (N_2503,In_407,In_1291);
or U2504 (N_2504,In_1410,In_1123);
nor U2505 (N_2505,In_351,In_988);
or U2506 (N_2506,In_1342,In_316);
nand U2507 (N_2507,In_1059,In_1019);
nor U2508 (N_2508,In_315,In_10);
nand U2509 (N_2509,In_741,In_717);
and U2510 (N_2510,In_319,In_722);
and U2511 (N_2511,In_826,In_485);
nor U2512 (N_2512,In_786,In_1330);
or U2513 (N_2513,In_39,In_1437);
or U2514 (N_2514,In_502,In_1024);
and U2515 (N_2515,In_1265,In_687);
or U2516 (N_2516,In_485,In_1203);
and U2517 (N_2517,In_154,In_916);
or U2518 (N_2518,In_646,In_597);
or U2519 (N_2519,In_838,In_1372);
nand U2520 (N_2520,In_877,In_115);
or U2521 (N_2521,In_304,In_485);
nand U2522 (N_2522,In_274,In_1173);
or U2523 (N_2523,In_66,In_336);
or U2524 (N_2524,In_437,In_1248);
nand U2525 (N_2525,In_1310,In_1312);
xnor U2526 (N_2526,In_1442,In_1203);
nand U2527 (N_2527,In_1231,In_1381);
or U2528 (N_2528,In_581,In_365);
xor U2529 (N_2529,In_337,In_1462);
or U2530 (N_2530,In_120,In_160);
nand U2531 (N_2531,In_107,In_267);
and U2532 (N_2532,In_1486,In_199);
or U2533 (N_2533,In_683,In_277);
nor U2534 (N_2534,In_26,In_1348);
or U2535 (N_2535,In_398,In_731);
nor U2536 (N_2536,In_364,In_559);
and U2537 (N_2537,In_1456,In_939);
xor U2538 (N_2538,In_565,In_980);
xor U2539 (N_2539,In_634,In_1496);
nor U2540 (N_2540,In_1342,In_1049);
or U2541 (N_2541,In_344,In_819);
and U2542 (N_2542,In_1082,In_544);
nor U2543 (N_2543,In_891,In_983);
nor U2544 (N_2544,In_33,In_407);
or U2545 (N_2545,In_7,In_828);
and U2546 (N_2546,In_491,In_970);
or U2547 (N_2547,In_37,In_532);
nand U2548 (N_2548,In_99,In_660);
nand U2549 (N_2549,In_574,In_1133);
nor U2550 (N_2550,In_1137,In_1208);
and U2551 (N_2551,In_1146,In_356);
nand U2552 (N_2552,In_1486,In_1443);
or U2553 (N_2553,In_1270,In_668);
nor U2554 (N_2554,In_160,In_550);
nor U2555 (N_2555,In_386,In_700);
and U2556 (N_2556,In_36,In_1274);
nor U2557 (N_2557,In_526,In_1478);
nand U2558 (N_2558,In_693,In_239);
and U2559 (N_2559,In_677,In_1149);
or U2560 (N_2560,In_165,In_1307);
or U2561 (N_2561,In_511,In_236);
nor U2562 (N_2562,In_630,In_728);
or U2563 (N_2563,In_954,In_923);
or U2564 (N_2564,In_837,In_1112);
or U2565 (N_2565,In_813,In_1437);
and U2566 (N_2566,In_618,In_407);
xnor U2567 (N_2567,In_1250,In_781);
nor U2568 (N_2568,In_137,In_1073);
or U2569 (N_2569,In_553,In_182);
nor U2570 (N_2570,In_1266,In_1317);
nand U2571 (N_2571,In_336,In_1081);
and U2572 (N_2572,In_505,In_44);
and U2573 (N_2573,In_1138,In_842);
nand U2574 (N_2574,In_52,In_1088);
nand U2575 (N_2575,In_1194,In_1219);
nand U2576 (N_2576,In_679,In_705);
nand U2577 (N_2577,In_33,In_995);
nor U2578 (N_2578,In_365,In_526);
nor U2579 (N_2579,In_738,In_1442);
and U2580 (N_2580,In_658,In_1253);
nor U2581 (N_2581,In_103,In_1146);
or U2582 (N_2582,In_598,In_127);
and U2583 (N_2583,In_1105,In_785);
or U2584 (N_2584,In_86,In_1222);
or U2585 (N_2585,In_571,In_1470);
and U2586 (N_2586,In_263,In_108);
and U2587 (N_2587,In_555,In_1203);
xnor U2588 (N_2588,In_1168,In_224);
or U2589 (N_2589,In_839,In_1250);
and U2590 (N_2590,In_532,In_659);
or U2591 (N_2591,In_51,In_859);
xnor U2592 (N_2592,In_977,In_502);
and U2593 (N_2593,In_321,In_1288);
nand U2594 (N_2594,In_575,In_1203);
nand U2595 (N_2595,In_93,In_904);
nand U2596 (N_2596,In_1207,In_1297);
and U2597 (N_2597,In_1099,In_712);
or U2598 (N_2598,In_516,In_1152);
and U2599 (N_2599,In_305,In_539);
or U2600 (N_2600,In_215,In_814);
and U2601 (N_2601,In_747,In_991);
and U2602 (N_2602,In_274,In_1403);
nor U2603 (N_2603,In_630,In_1401);
and U2604 (N_2604,In_1421,In_896);
nor U2605 (N_2605,In_1031,In_1170);
nor U2606 (N_2606,In_1129,In_922);
nand U2607 (N_2607,In_1289,In_579);
or U2608 (N_2608,In_273,In_327);
and U2609 (N_2609,In_257,In_923);
nor U2610 (N_2610,In_1375,In_1308);
nand U2611 (N_2611,In_816,In_724);
nand U2612 (N_2612,In_341,In_1373);
nor U2613 (N_2613,In_220,In_943);
nor U2614 (N_2614,In_944,In_300);
nand U2615 (N_2615,In_639,In_230);
xor U2616 (N_2616,In_1080,In_63);
and U2617 (N_2617,In_679,In_1325);
nand U2618 (N_2618,In_724,In_224);
nand U2619 (N_2619,In_346,In_1039);
or U2620 (N_2620,In_333,In_362);
nand U2621 (N_2621,In_1382,In_829);
xnor U2622 (N_2622,In_973,In_1145);
and U2623 (N_2623,In_403,In_546);
nand U2624 (N_2624,In_19,In_1075);
and U2625 (N_2625,In_640,In_154);
nor U2626 (N_2626,In_957,In_267);
nor U2627 (N_2627,In_661,In_803);
or U2628 (N_2628,In_1193,In_1189);
or U2629 (N_2629,In_1182,In_266);
nor U2630 (N_2630,In_142,In_1050);
xnor U2631 (N_2631,In_570,In_264);
nor U2632 (N_2632,In_35,In_255);
or U2633 (N_2633,In_689,In_121);
or U2634 (N_2634,In_1153,In_794);
nor U2635 (N_2635,In_38,In_607);
or U2636 (N_2636,In_633,In_728);
nand U2637 (N_2637,In_807,In_642);
nor U2638 (N_2638,In_526,In_1269);
or U2639 (N_2639,In_807,In_271);
and U2640 (N_2640,In_1334,In_1006);
nor U2641 (N_2641,In_1324,In_897);
nand U2642 (N_2642,In_661,In_92);
nor U2643 (N_2643,In_14,In_590);
nor U2644 (N_2644,In_511,In_1441);
and U2645 (N_2645,In_706,In_1461);
and U2646 (N_2646,In_1039,In_931);
and U2647 (N_2647,In_1313,In_1175);
and U2648 (N_2648,In_155,In_71);
xor U2649 (N_2649,In_351,In_69);
or U2650 (N_2650,In_990,In_1484);
nand U2651 (N_2651,In_78,In_1325);
nor U2652 (N_2652,In_1129,In_1146);
or U2653 (N_2653,In_1213,In_878);
nor U2654 (N_2654,In_408,In_352);
nand U2655 (N_2655,In_49,In_139);
and U2656 (N_2656,In_423,In_1028);
or U2657 (N_2657,In_267,In_320);
or U2658 (N_2658,In_1422,In_1239);
and U2659 (N_2659,In_86,In_43);
nor U2660 (N_2660,In_279,In_892);
and U2661 (N_2661,In_470,In_491);
nand U2662 (N_2662,In_1326,In_1098);
and U2663 (N_2663,In_666,In_941);
or U2664 (N_2664,In_526,In_1224);
nand U2665 (N_2665,In_97,In_38);
xnor U2666 (N_2666,In_291,In_685);
xor U2667 (N_2667,In_1466,In_485);
nand U2668 (N_2668,In_920,In_807);
or U2669 (N_2669,In_75,In_1066);
nand U2670 (N_2670,In_663,In_352);
nand U2671 (N_2671,In_637,In_585);
nor U2672 (N_2672,In_928,In_1277);
or U2673 (N_2673,In_327,In_65);
nor U2674 (N_2674,In_729,In_1172);
xor U2675 (N_2675,In_1069,In_1485);
xor U2676 (N_2676,In_761,In_793);
or U2677 (N_2677,In_177,In_8);
or U2678 (N_2678,In_566,In_570);
and U2679 (N_2679,In_504,In_1205);
nor U2680 (N_2680,In_522,In_966);
nand U2681 (N_2681,In_639,In_665);
and U2682 (N_2682,In_1028,In_672);
nor U2683 (N_2683,In_560,In_1097);
and U2684 (N_2684,In_530,In_655);
and U2685 (N_2685,In_1294,In_1196);
nand U2686 (N_2686,In_647,In_755);
or U2687 (N_2687,In_1344,In_937);
or U2688 (N_2688,In_30,In_563);
nand U2689 (N_2689,In_799,In_88);
or U2690 (N_2690,In_299,In_516);
nor U2691 (N_2691,In_1114,In_847);
nor U2692 (N_2692,In_254,In_56);
nand U2693 (N_2693,In_810,In_291);
nor U2694 (N_2694,In_745,In_951);
nand U2695 (N_2695,In_1014,In_405);
nor U2696 (N_2696,In_1117,In_380);
or U2697 (N_2697,In_949,In_459);
nor U2698 (N_2698,In_227,In_857);
nor U2699 (N_2699,In_357,In_1282);
and U2700 (N_2700,In_420,In_510);
or U2701 (N_2701,In_757,In_130);
and U2702 (N_2702,In_24,In_814);
and U2703 (N_2703,In_784,In_1112);
and U2704 (N_2704,In_199,In_1423);
and U2705 (N_2705,In_282,In_23);
nand U2706 (N_2706,In_1388,In_373);
nand U2707 (N_2707,In_1361,In_1359);
or U2708 (N_2708,In_975,In_767);
nand U2709 (N_2709,In_436,In_1205);
and U2710 (N_2710,In_944,In_1324);
or U2711 (N_2711,In_591,In_1078);
and U2712 (N_2712,In_365,In_141);
nor U2713 (N_2713,In_1018,In_1462);
nor U2714 (N_2714,In_1283,In_543);
xnor U2715 (N_2715,In_770,In_349);
nor U2716 (N_2716,In_68,In_1145);
and U2717 (N_2717,In_128,In_669);
or U2718 (N_2718,In_390,In_447);
nand U2719 (N_2719,In_258,In_559);
nand U2720 (N_2720,In_1259,In_776);
nand U2721 (N_2721,In_1263,In_516);
nand U2722 (N_2722,In_1154,In_245);
nand U2723 (N_2723,In_912,In_1047);
and U2724 (N_2724,In_591,In_1253);
and U2725 (N_2725,In_917,In_367);
or U2726 (N_2726,In_695,In_10);
xnor U2727 (N_2727,In_986,In_1496);
nand U2728 (N_2728,In_1192,In_1010);
or U2729 (N_2729,In_1112,In_467);
xnor U2730 (N_2730,In_1382,In_1207);
and U2731 (N_2731,In_955,In_1347);
xor U2732 (N_2732,In_780,In_137);
and U2733 (N_2733,In_1228,In_1493);
and U2734 (N_2734,In_441,In_777);
nand U2735 (N_2735,In_1108,In_309);
or U2736 (N_2736,In_1146,In_1274);
nand U2737 (N_2737,In_1022,In_1085);
and U2738 (N_2738,In_1457,In_200);
nor U2739 (N_2739,In_627,In_176);
and U2740 (N_2740,In_1297,In_157);
or U2741 (N_2741,In_791,In_200);
or U2742 (N_2742,In_1481,In_374);
xnor U2743 (N_2743,In_1165,In_15);
nor U2744 (N_2744,In_449,In_1269);
xor U2745 (N_2745,In_157,In_1047);
nor U2746 (N_2746,In_916,In_1241);
or U2747 (N_2747,In_247,In_705);
nor U2748 (N_2748,In_558,In_1193);
nor U2749 (N_2749,In_173,In_530);
nand U2750 (N_2750,In_1367,In_419);
and U2751 (N_2751,In_1101,In_643);
nand U2752 (N_2752,In_368,In_442);
or U2753 (N_2753,In_1497,In_85);
and U2754 (N_2754,In_86,In_627);
and U2755 (N_2755,In_411,In_825);
and U2756 (N_2756,In_555,In_978);
or U2757 (N_2757,In_925,In_603);
or U2758 (N_2758,In_618,In_327);
or U2759 (N_2759,In_2,In_1186);
or U2760 (N_2760,In_626,In_649);
and U2761 (N_2761,In_393,In_1266);
nor U2762 (N_2762,In_878,In_1192);
and U2763 (N_2763,In_1319,In_652);
xnor U2764 (N_2764,In_949,In_657);
or U2765 (N_2765,In_97,In_1250);
and U2766 (N_2766,In_1035,In_900);
nor U2767 (N_2767,In_1472,In_771);
or U2768 (N_2768,In_1245,In_68);
nand U2769 (N_2769,In_563,In_157);
and U2770 (N_2770,In_1265,In_17);
or U2771 (N_2771,In_182,In_153);
nand U2772 (N_2772,In_161,In_1132);
nor U2773 (N_2773,In_333,In_818);
nand U2774 (N_2774,In_226,In_915);
nor U2775 (N_2775,In_81,In_612);
and U2776 (N_2776,In_424,In_1109);
nand U2777 (N_2777,In_1215,In_1160);
nand U2778 (N_2778,In_25,In_480);
or U2779 (N_2779,In_1083,In_588);
and U2780 (N_2780,In_437,In_240);
and U2781 (N_2781,In_532,In_641);
nor U2782 (N_2782,In_759,In_1260);
nand U2783 (N_2783,In_1265,In_799);
nand U2784 (N_2784,In_1217,In_153);
or U2785 (N_2785,In_1137,In_312);
xor U2786 (N_2786,In_703,In_1366);
nor U2787 (N_2787,In_1347,In_673);
or U2788 (N_2788,In_1340,In_24);
and U2789 (N_2789,In_1323,In_298);
xnor U2790 (N_2790,In_1038,In_789);
nor U2791 (N_2791,In_915,In_352);
and U2792 (N_2792,In_483,In_1498);
nor U2793 (N_2793,In_351,In_902);
or U2794 (N_2794,In_1278,In_275);
nand U2795 (N_2795,In_1152,In_701);
nor U2796 (N_2796,In_307,In_1172);
nand U2797 (N_2797,In_355,In_1070);
or U2798 (N_2798,In_1436,In_938);
nand U2799 (N_2799,In_157,In_794);
and U2800 (N_2800,In_384,In_835);
or U2801 (N_2801,In_403,In_577);
and U2802 (N_2802,In_1385,In_1055);
nand U2803 (N_2803,In_382,In_1138);
or U2804 (N_2804,In_1328,In_1246);
and U2805 (N_2805,In_1490,In_515);
and U2806 (N_2806,In_1369,In_1068);
xor U2807 (N_2807,In_1165,In_407);
xor U2808 (N_2808,In_226,In_1455);
and U2809 (N_2809,In_1257,In_1028);
nor U2810 (N_2810,In_654,In_1036);
nor U2811 (N_2811,In_711,In_1079);
xnor U2812 (N_2812,In_964,In_169);
nand U2813 (N_2813,In_1069,In_1231);
or U2814 (N_2814,In_1459,In_88);
and U2815 (N_2815,In_1327,In_166);
and U2816 (N_2816,In_757,In_584);
nor U2817 (N_2817,In_1461,In_1134);
or U2818 (N_2818,In_277,In_1321);
xnor U2819 (N_2819,In_171,In_1432);
nor U2820 (N_2820,In_969,In_186);
nand U2821 (N_2821,In_767,In_159);
nor U2822 (N_2822,In_1388,In_648);
nand U2823 (N_2823,In_322,In_1414);
and U2824 (N_2824,In_435,In_1135);
nand U2825 (N_2825,In_180,In_1299);
nor U2826 (N_2826,In_852,In_450);
or U2827 (N_2827,In_752,In_269);
and U2828 (N_2828,In_480,In_142);
nand U2829 (N_2829,In_807,In_1109);
nand U2830 (N_2830,In_170,In_1308);
nor U2831 (N_2831,In_1441,In_745);
and U2832 (N_2832,In_276,In_732);
xnor U2833 (N_2833,In_518,In_1220);
xor U2834 (N_2834,In_767,In_754);
nand U2835 (N_2835,In_1353,In_5);
or U2836 (N_2836,In_271,In_799);
and U2837 (N_2837,In_1052,In_65);
nand U2838 (N_2838,In_965,In_609);
nand U2839 (N_2839,In_1026,In_533);
xor U2840 (N_2840,In_873,In_942);
nand U2841 (N_2841,In_842,In_767);
or U2842 (N_2842,In_872,In_885);
xnor U2843 (N_2843,In_1454,In_447);
and U2844 (N_2844,In_686,In_343);
nor U2845 (N_2845,In_61,In_914);
and U2846 (N_2846,In_394,In_93);
and U2847 (N_2847,In_1138,In_265);
or U2848 (N_2848,In_548,In_638);
and U2849 (N_2849,In_520,In_174);
nand U2850 (N_2850,In_286,In_633);
or U2851 (N_2851,In_830,In_119);
or U2852 (N_2852,In_146,In_996);
nor U2853 (N_2853,In_1028,In_1180);
nand U2854 (N_2854,In_1074,In_466);
and U2855 (N_2855,In_267,In_428);
xnor U2856 (N_2856,In_9,In_1401);
or U2857 (N_2857,In_440,In_755);
xnor U2858 (N_2858,In_207,In_1144);
or U2859 (N_2859,In_258,In_450);
and U2860 (N_2860,In_1336,In_842);
nand U2861 (N_2861,In_17,In_57);
and U2862 (N_2862,In_1371,In_227);
nor U2863 (N_2863,In_332,In_867);
or U2864 (N_2864,In_297,In_865);
nand U2865 (N_2865,In_687,In_493);
or U2866 (N_2866,In_833,In_54);
nor U2867 (N_2867,In_128,In_471);
nor U2868 (N_2868,In_288,In_426);
xor U2869 (N_2869,In_1481,In_353);
nand U2870 (N_2870,In_210,In_60);
nand U2871 (N_2871,In_1015,In_123);
nor U2872 (N_2872,In_346,In_1348);
nand U2873 (N_2873,In_491,In_1234);
nand U2874 (N_2874,In_812,In_499);
or U2875 (N_2875,In_535,In_1382);
nand U2876 (N_2876,In_25,In_1177);
or U2877 (N_2877,In_661,In_616);
or U2878 (N_2878,In_649,In_929);
or U2879 (N_2879,In_321,In_505);
nor U2880 (N_2880,In_1155,In_498);
or U2881 (N_2881,In_374,In_1349);
and U2882 (N_2882,In_547,In_1142);
nand U2883 (N_2883,In_764,In_147);
nor U2884 (N_2884,In_648,In_751);
and U2885 (N_2885,In_959,In_1084);
or U2886 (N_2886,In_587,In_336);
and U2887 (N_2887,In_614,In_42);
nand U2888 (N_2888,In_1019,In_210);
or U2889 (N_2889,In_490,In_475);
nand U2890 (N_2890,In_738,In_125);
nor U2891 (N_2891,In_1410,In_1327);
xnor U2892 (N_2892,In_1256,In_1431);
and U2893 (N_2893,In_468,In_561);
or U2894 (N_2894,In_433,In_484);
and U2895 (N_2895,In_1,In_133);
and U2896 (N_2896,In_882,In_380);
and U2897 (N_2897,In_1149,In_23);
xnor U2898 (N_2898,In_470,In_1227);
or U2899 (N_2899,In_302,In_905);
xor U2900 (N_2900,In_444,In_406);
or U2901 (N_2901,In_347,In_1296);
xnor U2902 (N_2902,In_1127,In_1336);
and U2903 (N_2903,In_1163,In_1183);
and U2904 (N_2904,In_415,In_677);
and U2905 (N_2905,In_84,In_93);
nand U2906 (N_2906,In_1113,In_435);
nor U2907 (N_2907,In_1182,In_1128);
nand U2908 (N_2908,In_609,In_71);
and U2909 (N_2909,In_1085,In_1071);
nor U2910 (N_2910,In_715,In_192);
xnor U2911 (N_2911,In_703,In_686);
or U2912 (N_2912,In_699,In_199);
xor U2913 (N_2913,In_1417,In_634);
xnor U2914 (N_2914,In_771,In_199);
nand U2915 (N_2915,In_1247,In_551);
and U2916 (N_2916,In_1263,In_159);
and U2917 (N_2917,In_264,In_848);
nand U2918 (N_2918,In_783,In_451);
nand U2919 (N_2919,In_164,In_406);
nor U2920 (N_2920,In_1048,In_1223);
or U2921 (N_2921,In_1294,In_494);
or U2922 (N_2922,In_355,In_816);
or U2923 (N_2923,In_1463,In_380);
and U2924 (N_2924,In_835,In_1438);
or U2925 (N_2925,In_635,In_990);
and U2926 (N_2926,In_1464,In_1327);
nor U2927 (N_2927,In_168,In_1159);
nand U2928 (N_2928,In_1491,In_242);
or U2929 (N_2929,In_1047,In_960);
nand U2930 (N_2930,In_381,In_705);
nor U2931 (N_2931,In_502,In_1392);
and U2932 (N_2932,In_902,In_758);
or U2933 (N_2933,In_1062,In_78);
nand U2934 (N_2934,In_483,In_1172);
nand U2935 (N_2935,In_608,In_636);
nand U2936 (N_2936,In_903,In_340);
and U2937 (N_2937,In_1330,In_942);
nor U2938 (N_2938,In_417,In_1163);
and U2939 (N_2939,In_1350,In_987);
nor U2940 (N_2940,In_1417,In_1459);
nand U2941 (N_2941,In_1449,In_351);
and U2942 (N_2942,In_464,In_661);
and U2943 (N_2943,In_77,In_215);
xnor U2944 (N_2944,In_1138,In_167);
nand U2945 (N_2945,In_1265,In_76);
and U2946 (N_2946,In_154,In_227);
nor U2947 (N_2947,In_1139,In_1112);
or U2948 (N_2948,In_880,In_802);
nor U2949 (N_2949,In_760,In_204);
or U2950 (N_2950,In_1360,In_484);
nand U2951 (N_2951,In_272,In_113);
nand U2952 (N_2952,In_246,In_830);
xnor U2953 (N_2953,In_639,In_1491);
and U2954 (N_2954,In_1279,In_423);
nor U2955 (N_2955,In_205,In_453);
nor U2956 (N_2956,In_1008,In_652);
and U2957 (N_2957,In_389,In_331);
nand U2958 (N_2958,In_104,In_1066);
or U2959 (N_2959,In_126,In_962);
nand U2960 (N_2960,In_1387,In_107);
nor U2961 (N_2961,In_395,In_615);
xnor U2962 (N_2962,In_281,In_857);
nor U2963 (N_2963,In_50,In_97);
and U2964 (N_2964,In_640,In_10);
nor U2965 (N_2965,In_1110,In_497);
nand U2966 (N_2966,In_1105,In_395);
nand U2967 (N_2967,In_594,In_962);
nand U2968 (N_2968,In_857,In_570);
xor U2969 (N_2969,In_979,In_800);
nor U2970 (N_2970,In_626,In_1220);
nand U2971 (N_2971,In_663,In_1000);
nand U2972 (N_2972,In_1402,In_1353);
or U2973 (N_2973,In_1281,In_549);
nor U2974 (N_2974,In_1206,In_988);
or U2975 (N_2975,In_574,In_712);
nor U2976 (N_2976,In_1050,In_209);
or U2977 (N_2977,In_992,In_897);
and U2978 (N_2978,In_639,In_977);
and U2979 (N_2979,In_647,In_339);
nor U2980 (N_2980,In_705,In_942);
nand U2981 (N_2981,In_466,In_282);
or U2982 (N_2982,In_681,In_490);
or U2983 (N_2983,In_800,In_161);
nand U2984 (N_2984,In_1047,In_96);
nor U2985 (N_2985,In_1125,In_1299);
and U2986 (N_2986,In_1281,In_1101);
or U2987 (N_2987,In_1425,In_254);
nor U2988 (N_2988,In_764,In_190);
nand U2989 (N_2989,In_335,In_1152);
nor U2990 (N_2990,In_238,In_1404);
nor U2991 (N_2991,In_434,In_1210);
nor U2992 (N_2992,In_916,In_908);
or U2993 (N_2993,In_41,In_1162);
or U2994 (N_2994,In_334,In_617);
or U2995 (N_2995,In_173,In_1115);
nor U2996 (N_2996,In_165,In_903);
and U2997 (N_2997,In_905,In_1371);
nand U2998 (N_2998,In_79,In_1037);
nor U2999 (N_2999,In_731,In_43);
and U3000 (N_3000,N_1744,N_969);
nand U3001 (N_3001,N_2741,N_1531);
xor U3002 (N_3002,N_2020,N_1316);
nand U3003 (N_3003,N_812,N_2866);
xnor U3004 (N_3004,N_913,N_1692);
nor U3005 (N_3005,N_1721,N_1218);
and U3006 (N_3006,N_307,N_1805);
nand U3007 (N_3007,N_617,N_2422);
or U3008 (N_3008,N_1048,N_1802);
or U3009 (N_3009,N_1090,N_1831);
or U3010 (N_3010,N_1340,N_2049);
nand U3011 (N_3011,N_710,N_1987);
nand U3012 (N_3012,N_1346,N_511);
and U3013 (N_3013,N_1251,N_1247);
and U3014 (N_3014,N_1973,N_1573);
nor U3015 (N_3015,N_286,N_323);
and U3016 (N_3016,N_2805,N_292);
nand U3017 (N_3017,N_94,N_1659);
nor U3018 (N_3018,N_2554,N_165);
and U3019 (N_3019,N_52,N_2197);
or U3020 (N_3020,N_2025,N_862);
and U3021 (N_3021,N_2100,N_1915);
nor U3022 (N_3022,N_99,N_2346);
or U3023 (N_3023,N_927,N_688);
or U3024 (N_3024,N_2870,N_2395);
or U3025 (N_3025,N_2759,N_2340);
nand U3026 (N_3026,N_379,N_1804);
and U3027 (N_3027,N_2970,N_818);
nor U3028 (N_3028,N_938,N_48);
xnor U3029 (N_3029,N_437,N_2338);
and U3030 (N_3030,N_470,N_2596);
nor U3031 (N_3031,N_126,N_1164);
or U3032 (N_3032,N_169,N_2743);
and U3033 (N_3033,N_2221,N_2914);
nand U3034 (N_3034,N_0,N_1555);
and U3035 (N_3035,N_721,N_1442);
and U3036 (N_3036,N_2522,N_289);
or U3037 (N_3037,N_1897,N_2061);
nor U3038 (N_3038,N_2872,N_860);
or U3039 (N_3039,N_2074,N_541);
nor U3040 (N_3040,N_1956,N_1623);
nand U3041 (N_3041,N_1731,N_751);
or U3042 (N_3042,N_76,N_1726);
and U3043 (N_3043,N_1628,N_1222);
nor U3044 (N_3044,N_162,N_895);
nand U3045 (N_3045,N_2463,N_919);
nor U3046 (N_3046,N_2862,N_1453);
nand U3047 (N_3047,N_728,N_1200);
or U3048 (N_3048,N_213,N_987);
nand U3049 (N_3049,N_1195,N_2719);
nand U3050 (N_3050,N_1756,N_2246);
nand U3051 (N_3051,N_2734,N_472);
nand U3052 (N_3052,N_2644,N_431);
nor U3053 (N_3053,N_610,N_448);
or U3054 (N_3054,N_2259,N_1906);
nor U3055 (N_3055,N_2194,N_426);
nand U3056 (N_3056,N_1097,N_168);
and U3057 (N_3057,N_2302,N_1064);
nor U3058 (N_3058,N_2566,N_2236);
nand U3059 (N_3059,N_1369,N_2528);
and U3060 (N_3060,N_2934,N_2956);
and U3061 (N_3061,N_2264,N_1053);
or U3062 (N_3062,N_1440,N_2949);
nor U3063 (N_3063,N_2313,N_1554);
nor U3064 (N_3064,N_1753,N_800);
nand U3065 (N_3065,N_1852,N_257);
and U3066 (N_3066,N_641,N_2411);
nor U3067 (N_3067,N_2048,N_1790);
nand U3068 (N_3068,N_2986,N_1381);
nor U3069 (N_3069,N_1888,N_2925);
and U3070 (N_3070,N_1201,N_424);
and U3071 (N_3071,N_604,N_329);
nand U3072 (N_3072,N_2916,N_1544);
and U3073 (N_3073,N_67,N_2114);
xnor U3074 (N_3074,N_759,N_1770);
nor U3075 (N_3075,N_2928,N_1035);
and U3076 (N_3076,N_2184,N_857);
and U3077 (N_3077,N_79,N_1158);
or U3078 (N_3078,N_1582,N_2900);
nor U3079 (N_3079,N_1191,N_2877);
nor U3080 (N_3080,N_2372,N_1058);
and U3081 (N_3081,N_1073,N_2014);
xor U3082 (N_3082,N_348,N_1905);
nor U3083 (N_3083,N_504,N_1745);
and U3084 (N_3084,N_907,N_106);
nand U3085 (N_3085,N_2398,N_1287);
xor U3086 (N_3086,N_1822,N_135);
and U3087 (N_3087,N_1597,N_219);
nor U3088 (N_3088,N_497,N_2849);
nand U3089 (N_3089,N_1736,N_1685);
nand U3090 (N_3090,N_1416,N_1793);
xor U3091 (N_3091,N_941,N_2193);
xor U3092 (N_3092,N_455,N_1909);
nand U3093 (N_3093,N_2196,N_225);
or U3094 (N_3094,N_130,N_2035);
nor U3095 (N_3095,N_2881,N_2141);
xnor U3096 (N_3096,N_4,N_1787);
and U3097 (N_3097,N_844,N_193);
and U3098 (N_3098,N_397,N_2843);
nand U3099 (N_3099,N_360,N_1147);
or U3100 (N_3100,N_1611,N_2195);
and U3101 (N_3101,N_2278,N_2590);
xor U3102 (N_3102,N_833,N_77);
and U3103 (N_3103,N_897,N_625);
nand U3104 (N_3104,N_2433,N_2892);
nand U3105 (N_3105,N_1275,N_2825);
nand U3106 (N_3106,N_117,N_2845);
xor U3107 (N_3107,N_2107,N_2532);
and U3108 (N_3108,N_354,N_2387);
nand U3109 (N_3109,N_2146,N_2622);
and U3110 (N_3110,N_1705,N_295);
nor U3111 (N_3111,N_2527,N_1403);
nand U3112 (N_3112,N_1496,N_1697);
and U3113 (N_3113,N_2455,N_847);
or U3114 (N_3114,N_1036,N_140);
and U3115 (N_3115,N_2242,N_246);
nand U3116 (N_3116,N_1478,N_2327);
and U3117 (N_3117,N_2469,N_1245);
or U3118 (N_3118,N_105,N_2669);
nand U3119 (N_3119,N_316,N_2772);
and U3120 (N_3120,N_1872,N_2628);
nor U3121 (N_3121,N_2329,N_2738);
nand U3122 (N_3122,N_935,N_2751);
nor U3123 (N_3123,N_1886,N_731);
or U3124 (N_3124,N_1690,N_807);
and U3125 (N_3125,N_946,N_2075);
or U3126 (N_3126,N_1710,N_43);
and U3127 (N_3127,N_1171,N_1389);
nor U3128 (N_3128,N_1278,N_1627);
nand U3129 (N_3129,N_414,N_1684);
and U3130 (N_3130,N_1625,N_1314);
or U3131 (N_3131,N_1299,N_1165);
or U3132 (N_3132,N_2247,N_221);
or U3133 (N_3133,N_757,N_1142);
nor U3134 (N_3134,N_2295,N_1920);
and U3135 (N_3135,N_1312,N_2981);
xnor U3136 (N_3136,N_2686,N_1012);
or U3137 (N_3137,N_2478,N_1994);
nand U3138 (N_3138,N_944,N_365);
nand U3139 (N_3139,N_532,N_2535);
nand U3140 (N_3140,N_2477,N_1493);
or U3141 (N_3141,N_1373,N_2919);
xor U3142 (N_3142,N_1564,N_1594);
nor U3143 (N_3143,N_963,N_1491);
nand U3144 (N_3144,N_803,N_1683);
xor U3145 (N_3145,N_409,N_1460);
or U3146 (N_3146,N_2178,N_2303);
or U3147 (N_3147,N_1211,N_1999);
or U3148 (N_3148,N_551,N_2063);
nor U3149 (N_3149,N_1452,N_264);
nor U3150 (N_3150,N_765,N_420);
nor U3151 (N_3151,N_2572,N_2248);
xnor U3152 (N_3152,N_110,N_2471);
or U3153 (N_3153,N_1724,N_367);
or U3154 (N_3154,N_2503,N_1118);
and U3155 (N_3155,N_2638,N_708);
and U3156 (N_3156,N_2036,N_1370);
and U3157 (N_3157,N_603,N_2655);
nor U3158 (N_3158,N_1830,N_1434);
and U3159 (N_3159,N_1159,N_1656);
and U3160 (N_3160,N_1993,N_1444);
and U3161 (N_3161,N_1576,N_934);
or U3162 (N_3162,N_239,N_700);
and U3163 (N_3163,N_2988,N_100);
nand U3164 (N_3164,N_1034,N_1655);
or U3165 (N_3165,N_911,N_2022);
and U3166 (N_3166,N_328,N_1031);
or U3167 (N_3167,N_1672,N_2488);
nor U3168 (N_3168,N_1483,N_482);
and U3169 (N_3169,N_2267,N_1382);
nor U3170 (N_3170,N_1912,N_549);
xor U3171 (N_3171,N_748,N_306);
and U3172 (N_3172,N_872,N_1621);
xnor U3173 (N_3173,N_98,N_386);
nor U3174 (N_3174,N_271,N_2320);
or U3175 (N_3175,N_33,N_2089);
or U3176 (N_3176,N_716,N_2162);
and U3177 (N_3177,N_754,N_2927);
nor U3178 (N_3178,N_1936,N_121);
nand U3179 (N_3179,N_1873,N_2721);
nand U3180 (N_3180,N_1928,N_1739);
nor U3181 (N_3181,N_794,N_650);
nor U3182 (N_3182,N_2679,N_498);
or U3183 (N_3183,N_815,N_2834);
or U3184 (N_3184,N_1867,N_2860);
and U3185 (N_3185,N_703,N_1182);
or U3186 (N_3186,N_1521,N_285);
or U3187 (N_3187,N_1931,N_997);
and U3188 (N_3188,N_2332,N_2869);
nand U3189 (N_3189,N_1348,N_2873);
xor U3190 (N_3190,N_2182,N_1466);
and U3191 (N_3191,N_1155,N_875);
and U3192 (N_3192,N_1860,N_396);
and U3193 (N_3193,N_2219,N_1894);
nor U3194 (N_3194,N_172,N_1789);
and U3195 (N_3195,N_2637,N_2487);
nand U3196 (N_3196,N_45,N_1168);
nand U3197 (N_3197,N_2363,N_1589);
and U3198 (N_3198,N_839,N_1797);
and U3199 (N_3199,N_1061,N_2428);
and U3200 (N_3200,N_2567,N_2533);
or U3201 (N_3201,N_419,N_693);
or U3202 (N_3202,N_977,N_324);
or U3203 (N_3203,N_107,N_2967);
nand U3204 (N_3204,N_2462,N_1242);
and U3205 (N_3205,N_988,N_1652);
nor U3206 (N_3206,N_1341,N_2524);
or U3207 (N_3207,N_1429,N_910);
and U3208 (N_3208,N_1832,N_903);
nor U3209 (N_3209,N_1911,N_2360);
and U3210 (N_3210,N_2798,N_799);
and U3211 (N_3211,N_2672,N_1244);
or U3212 (N_3212,N_1393,N_2552);
nand U3213 (N_3213,N_341,N_1096);
nand U3214 (N_3214,N_590,N_901);
nor U3215 (N_3215,N_2895,N_2274);
and U3216 (N_3216,N_1292,N_620);
or U3217 (N_3217,N_567,N_2476);
or U3218 (N_3218,N_1448,N_1954);
nand U3219 (N_3219,N_114,N_1908);
nor U3220 (N_3220,N_745,N_1820);
nand U3221 (N_3221,N_444,N_2085);
nor U3222 (N_3222,N_667,N_1698);
and U3223 (N_3223,N_854,N_1892);
and U3224 (N_3224,N_273,N_1577);
or U3225 (N_3225,N_411,N_2775);
nand U3226 (N_3226,N_1835,N_572);
nor U3227 (N_3227,N_1866,N_2982);
nand U3228 (N_3228,N_2727,N_960);
or U3229 (N_3229,N_186,N_123);
or U3230 (N_3230,N_203,N_2262);
xnor U3231 (N_3231,N_493,N_142);
nand U3232 (N_3232,N_364,N_2296);
nand U3233 (N_3233,N_563,N_1113);
or U3234 (N_3234,N_2570,N_1713);
xor U3235 (N_3235,N_160,N_2565);
xor U3236 (N_3236,N_2850,N_326);
or U3237 (N_3237,N_90,N_1547);
nand U3238 (N_3238,N_291,N_2814);
or U3239 (N_3239,N_1047,N_993);
or U3240 (N_3240,N_654,N_2073);
nor U3241 (N_3241,N_2199,N_2763);
nor U3242 (N_3242,N_2865,N_91);
or U3243 (N_3243,N_653,N_2890);
nand U3244 (N_3244,N_525,N_1210);
nor U3245 (N_3245,N_2731,N_1005);
xor U3246 (N_3246,N_2645,N_446);
and U3247 (N_3247,N_2786,N_163);
nand U3248 (N_3248,N_133,N_2514);
nand U3249 (N_3249,N_599,N_2012);
xnor U3250 (N_3250,N_1425,N_1354);
xnor U3251 (N_3251,N_317,N_2801);
nand U3252 (N_3252,N_579,N_2762);
or U3253 (N_3253,N_920,N_2641);
nand U3254 (N_3254,N_2209,N_2044);
or U3255 (N_3255,N_1502,N_128);
xnor U3256 (N_3256,N_1996,N_2712);
or U3257 (N_3257,N_2132,N_1534);
nor U3258 (N_3258,N_2795,N_2019);
xor U3259 (N_3259,N_1421,N_2407);
or U3260 (N_3260,N_2081,N_1718);
nand U3261 (N_3261,N_1653,N_1116);
xnor U3262 (N_3262,N_1068,N_609);
and U3263 (N_3263,N_1431,N_1043);
or U3264 (N_3264,N_2308,N_931);
or U3265 (N_3265,N_2946,N_1426);
and U3266 (N_3266,N_1223,N_1809);
nor U3267 (N_3267,N_113,N_2349);
or U3268 (N_3268,N_202,N_527);
nor U3269 (N_3269,N_1612,N_2716);
or U3270 (N_3270,N_1654,N_1600);
or U3271 (N_3271,N_2750,N_2173);
nor U3272 (N_3272,N_2660,N_2060);
and U3273 (N_3273,N_209,N_1461);
nor U3274 (N_3274,N_1719,N_1458);
and U3275 (N_3275,N_2177,N_971);
xnor U3276 (N_3276,N_1439,N_119);
nor U3277 (N_3277,N_1940,N_1548);
nand U3278 (N_3278,N_1380,N_1896);
and U3279 (N_3279,N_2458,N_722);
nand U3280 (N_3280,N_2116,N_631);
or U3281 (N_3281,N_959,N_1467);
or U3282 (N_3282,N_711,N_1330);
and U3283 (N_3283,N_2347,N_1203);
or U3284 (N_3284,N_2508,N_509);
nor U3285 (N_3285,N_580,N_1870);
nand U3286 (N_3286,N_2656,N_1163);
nand U3287 (N_3287,N_683,N_2984);
and U3288 (N_3288,N_1841,N_2290);
xor U3289 (N_3289,N_2909,N_640);
nand U3290 (N_3290,N_164,N_2737);
and U3291 (N_3291,N_215,N_245);
or U3292 (N_3292,N_2551,N_1941);
nor U3293 (N_3293,N_47,N_2234);
nor U3294 (N_3294,N_1219,N_2930);
nand U3295 (N_3295,N_1405,N_55);
or U3296 (N_3296,N_909,N_1070);
nor U3297 (N_3297,N_1863,N_1591);
nor U3298 (N_3298,N_2440,N_2723);
or U3299 (N_3299,N_1844,N_2067);
or U3300 (N_3300,N_2220,N_924);
xor U3301 (N_3301,N_2942,N_974);
and U3302 (N_3302,N_1497,N_395);
or U3303 (N_3303,N_2192,N_972);
xnor U3304 (N_3304,N_1707,N_1855);
nor U3305 (N_3305,N_1711,N_2664);
or U3306 (N_3306,N_2013,N_2539);
nor U3307 (N_3307,N_1392,N_1332);
or U3308 (N_3308,N_1420,N_2657);
xor U3309 (N_3309,N_495,N_1456);
nand U3310 (N_3310,N_336,N_1136);
nand U3311 (N_3311,N_2200,N_1366);
xor U3312 (N_3312,N_2091,N_361);
or U3313 (N_3313,N_561,N_2926);
nor U3314 (N_3314,N_2228,N_1361);
and U3315 (N_3315,N_1230,N_1102);
nand U3316 (N_3316,N_2159,N_2382);
nor U3317 (N_3317,N_20,N_357);
and U3318 (N_3318,N_170,N_894);
nor U3319 (N_3319,N_2310,N_878);
and U3320 (N_3320,N_736,N_1984);
xnor U3321 (N_3321,N_2764,N_1174);
xnor U3322 (N_3322,N_1723,N_1372);
and U3323 (N_3323,N_837,N_2855);
nor U3324 (N_3324,N_531,N_2500);
xnor U3325 (N_3325,N_828,N_2465);
and U3326 (N_3326,N_2708,N_238);
and U3327 (N_3327,N_2709,N_2652);
nand U3328 (N_3328,N_1138,N_1678);
xor U3329 (N_3329,N_887,N_914);
nand U3330 (N_3330,N_2125,N_565);
nor U3331 (N_3331,N_1365,N_1030);
nor U3332 (N_3332,N_1350,N_1180);
or U3333 (N_3333,N_2612,N_1281);
or U3334 (N_3334,N_1500,N_2042);
or U3335 (N_3335,N_758,N_2187);
and U3336 (N_3336,N_252,N_756);
or U3337 (N_3337,N_1249,N_368);
nand U3338 (N_3338,N_192,N_2907);
and U3339 (N_3339,N_1666,N_2520);
xnor U3340 (N_3340,N_265,N_363);
and U3341 (N_3341,N_922,N_908);
nand U3342 (N_3342,N_59,N_115);
and U3343 (N_3343,N_450,N_2490);
nor U3344 (N_3344,N_1193,N_1749);
nand U3345 (N_3345,N_1122,N_1760);
nand U3346 (N_3346,N_1668,N_1995);
or U3347 (N_3347,N_2482,N_1585);
and U3348 (N_3348,N_1482,N_1949);
xor U3349 (N_3349,N_2856,N_1764);
nor U3350 (N_3350,N_2156,N_853);
nor U3351 (N_3351,N_380,N_1932);
nor U3352 (N_3352,N_524,N_1402);
nor U3353 (N_3353,N_836,N_2874);
xnor U3354 (N_3354,N_2375,N_1981);
or U3355 (N_3355,N_1781,N_744);
nand U3356 (N_3356,N_2714,N_372);
or U3357 (N_3357,N_218,N_2541);
nand U3358 (N_3358,N_967,N_902);
or U3359 (N_3359,N_1052,N_1812);
nor U3360 (N_3360,N_21,N_2083);
nor U3361 (N_3361,N_2413,N_1488);
nand U3362 (N_3362,N_224,N_1851);
or U3363 (N_3363,N_886,N_2837);
and U3364 (N_3364,N_2434,N_1085);
xor U3365 (N_3365,N_548,N_1103);
nor U3366 (N_3366,N_2037,N_2380);
nand U3367 (N_3367,N_2625,N_536);
nand U3368 (N_3368,N_2386,N_1955);
nor U3369 (N_3369,N_464,N_884);
and U3370 (N_3370,N_984,N_1066);
and U3371 (N_3371,N_280,N_429);
or U3372 (N_3372,N_1878,N_2113);
and U3373 (N_3373,N_267,N_2088);
nor U3374 (N_3374,N_999,N_1094);
and U3375 (N_3375,N_1379,N_1919);
nand U3376 (N_3376,N_1447,N_1100);
and U3377 (N_3377,N_2618,N_2505);
nand U3378 (N_3378,N_2486,N_662);
nor U3379 (N_3379,N_928,N_1811);
nor U3380 (N_3380,N_244,N_652);
nor U3381 (N_3381,N_787,N_2148);
nor U3382 (N_3382,N_241,N_322);
or U3383 (N_3383,N_262,N_190);
or U3384 (N_3384,N_1759,N_1111);
xor U3385 (N_3385,N_2766,N_2384);
nand U3386 (N_3386,N_1015,N_578);
nor U3387 (N_3387,N_2754,N_1227);
or U3388 (N_3388,N_2268,N_254);
nand U3389 (N_3389,N_449,N_1092);
nor U3390 (N_3390,N_510,N_2077);
nor U3391 (N_3391,N_356,N_427);
xor U3392 (N_3392,N_2852,N_1798);
nor U3393 (N_3393,N_2253,N_2365);
or U3394 (N_3394,N_212,N_2255);
or U3395 (N_3395,N_2168,N_739);
nand U3396 (N_3396,N_2442,N_1602);
or U3397 (N_3397,N_2050,N_1974);
nor U3398 (N_3398,N_1826,N_2968);
or U3399 (N_3399,N_2201,N_2677);
or U3400 (N_3400,N_1579,N_2039);
and U3401 (N_3401,N_2328,N_2740);
and U3402 (N_3402,N_2710,N_1128);
xnor U3403 (N_3403,N_992,N_1261);
nand U3404 (N_3404,N_2480,N_668);
nor U3405 (N_3405,N_1243,N_1950);
nor U3406 (N_3406,N_1963,N_1767);
nor U3407 (N_3407,N_1260,N_575);
nor U3408 (N_3408,N_523,N_1335);
and U3409 (N_3409,N_1948,N_643);
and U3410 (N_3410,N_933,N_2871);
nand U3411 (N_3411,N_584,N_1333);
nor U3412 (N_3412,N_1924,N_1410);
nand U3413 (N_3413,N_29,N_2103);
nand U3414 (N_3414,N_2630,N_622);
or U3415 (N_3415,N_964,N_2448);
or U3416 (N_3416,N_1008,N_125);
and U3417 (N_3417,N_1686,N_2207);
and U3418 (N_3418,N_1454,N_2693);
or U3419 (N_3419,N_2831,N_649);
xor U3420 (N_3420,N_321,N_2745);
nor U3421 (N_3421,N_775,N_473);
xor U3422 (N_3422,N_1490,N_2828);
nor U3423 (N_3423,N_1563,N_1838);
nor U3424 (N_3424,N_806,N_2931);
nor U3425 (N_3425,N_242,N_2359);
xnor U3426 (N_3426,N_1834,N_2033);
or U3427 (N_3427,N_2560,N_1971);
nor U3428 (N_3428,N_413,N_1042);
and U3429 (N_3429,N_2883,N_2393);
nand U3430 (N_3430,N_277,N_1451);
xor U3431 (N_3431,N_1303,N_2429);
nor U3432 (N_3432,N_597,N_1353);
nand U3433 (N_3433,N_2602,N_1875);
and U3434 (N_3434,N_1796,N_2249);
and U3435 (N_3435,N_2378,N_1825);
or U3436 (N_3436,N_642,N_841);
nor U3437 (N_3437,N_589,N_1693);
nor U3438 (N_3438,N_1004,N_1549);
or U3439 (N_3439,N_2474,N_829);
nor U3440 (N_3440,N_741,N_634);
and U3441 (N_3441,N_1120,N_223);
nand U3442 (N_3442,N_1587,N_1326);
and U3443 (N_3443,N_2229,N_2771);
xor U3444 (N_3444,N_2553,N_2886);
and U3445 (N_3445,N_1337,N_2582);
nor U3446 (N_3446,N_961,N_1022);
and U3447 (N_3447,N_2188,N_1485);
nand U3448 (N_3448,N_50,N_255);
and U3449 (N_3449,N_2120,N_1807);
and U3450 (N_3450,N_491,N_2127);
nor U3451 (N_3451,N_2893,N_1687);
nor U3452 (N_3452,N_2402,N_556);
or U3453 (N_3453,N_2975,N_1619);
nand U3454 (N_3454,N_461,N_1307);
nor U3455 (N_3455,N_2348,N_1728);
or U3456 (N_3456,N_2121,N_2726);
xor U3457 (N_3457,N_266,N_2951);
or U3458 (N_3458,N_1091,N_2041);
nor U3459 (N_3459,N_412,N_1757);
or U3460 (N_3460,N_69,N_766);
nor U3461 (N_3461,N_2932,N_12);
or U3462 (N_3462,N_2293,N_611);
xor U3463 (N_3463,N_606,N_2356);
nor U3464 (N_3464,N_989,N_702);
nand U3465 (N_3465,N_2810,N_2105);
and U3466 (N_3466,N_1637,N_453);
and U3467 (N_3467,N_1708,N_159);
xnor U3468 (N_3468,N_2822,N_2214);
and U3469 (N_3469,N_1327,N_674);
or U3470 (N_3470,N_715,N_1412);
or U3471 (N_3471,N_1509,N_1649);
xnor U3472 (N_3472,N_2286,N_767);
nor U3473 (N_3473,N_1647,N_1185);
and U3474 (N_3474,N_1065,N_2062);
nand U3475 (N_3475,N_2696,N_2435);
and U3476 (N_3476,N_467,N_229);
nor U3477 (N_3477,N_1153,N_1151);
or U3478 (N_3478,N_2096,N_982);
or U3479 (N_3479,N_342,N_2588);
or U3480 (N_3480,N_2773,N_1268);
and U3481 (N_3481,N_1527,N_2711);
or U3482 (N_3482,N_1651,N_1422);
xor U3483 (N_3483,N_2369,N_1917);
and U3484 (N_3484,N_216,N_2181);
nor U3485 (N_3485,N_1988,N_1902);
or U3486 (N_3486,N_2648,N_65);
nand U3487 (N_3487,N_687,N_2158);
nand U3488 (N_3488,N_2543,N_1028);
or U3489 (N_3489,N_2426,N_278);
nor U3490 (N_3490,N_2003,N_438);
or U3491 (N_3491,N_661,N_750);
or U3492 (N_3492,N_1057,N_535);
nor U3493 (N_3493,N_2854,N_2667);
or U3494 (N_3494,N_2017,N_1038);
nor U3495 (N_3495,N_808,N_1252);
nand U3496 (N_3496,N_2732,N_2307);
or U3497 (N_3497,N_970,N_2430);
nor U3498 (N_3498,N_2270,N_1140);
xor U3499 (N_3499,N_330,N_842);
nor U3500 (N_3500,N_331,N_1177);
or U3501 (N_3501,N_1978,N_1695);
nor U3502 (N_3502,N_2451,N_2343);
and U3503 (N_3503,N_2111,N_2492);
and U3504 (N_3504,N_1480,N_1965);
nand U3505 (N_3505,N_2544,N_2281);
nand U3506 (N_3506,N_651,N_2510);
and U3507 (N_3507,N_1847,N_1846);
and U3508 (N_3508,N_339,N_23);
and U3509 (N_3509,N_2636,N_184);
or U3510 (N_3510,N_663,N_2705);
nand U3511 (N_3511,N_75,N_2587);
or U3512 (N_3512,N_696,N_1593);
nand U3513 (N_3513,N_1550,N_279);
and U3514 (N_3514,N_299,N_1438);
and U3515 (N_3515,N_2634,N_15);
or U3516 (N_3516,N_868,N_2941);
and U3517 (N_3517,N_1259,N_2817);
or U3518 (N_3518,N_519,N_1682);
or U3519 (N_3519,N_2546,N_287);
or U3520 (N_3520,N_1428,N_2969);
and U3521 (N_3521,N_150,N_1119);
or U3522 (N_3522,N_1408,N_2604);
nand U3523 (N_3523,N_393,N_1725);
and U3524 (N_3524,N_51,N_2787);
nand U3525 (N_3525,N_263,N_2227);
xnor U3526 (N_3526,N_1712,N_2110);
nor U3527 (N_3527,N_188,N_1615);
or U3528 (N_3528,N_2506,N_780);
and U3529 (N_3529,N_2597,N_856);
or U3530 (N_3530,N_2231,N_645);
nand U3531 (N_3531,N_1143,N_2922);
nor U3532 (N_3532,N_2479,N_1856);
nand U3533 (N_3533,N_189,N_1418);
and U3534 (N_3534,N_425,N_2812);
nand U3535 (N_3535,N_2821,N_2432);
nand U3536 (N_3536,N_1212,N_1743);
nor U3537 (N_3537,N_161,N_529);
and U3538 (N_3538,N_846,N_1702);
nand U3539 (N_3539,N_647,N_293);
nor U3540 (N_3540,N_1514,N_2598);
and U3541 (N_3541,N_2397,N_309);
and U3542 (N_3542,N_1339,N_740);
nor U3543 (N_3543,N_592,N_2957);
and U3544 (N_3544,N_585,N_1877);
nand U3545 (N_3545,N_1300,N_1315);
or U3546 (N_3546,N_1964,N_2321);
and U3547 (N_3547,N_2939,N_1417);
nand U3548 (N_3548,N_1343,N_2918);
or U3549 (N_3549,N_870,N_1598);
nand U3550 (N_3550,N_619,N_699);
or U3551 (N_3551,N_891,N_103);
or U3552 (N_3552,N_2592,N_1127);
and U3553 (N_3553,N_1196,N_2903);
nor U3554 (N_3554,N_1779,N_2568);
or U3555 (N_3555,N_1238,N_1648);
nand U3556 (N_3556,N_1289,N_180);
nor U3557 (N_3557,N_2436,N_1293);
xor U3558 (N_3558,N_1101,N_174);
nand U3559 (N_3559,N_771,N_194);
and U3560 (N_3560,N_350,N_564);
and U3561 (N_3561,N_801,N_2747);
nand U3562 (N_3562,N_232,N_2216);
nor U3563 (N_3563,N_2999,N_1562);
nor U3564 (N_3564,N_937,N_2620);
or U3565 (N_3565,N_435,N_2779);
nor U3566 (N_3566,N_2796,N_433);
nand U3567 (N_3567,N_2300,N_777);
or U3568 (N_3568,N_352,N_2124);
xor U3569 (N_3569,N_1050,N_546);
nand U3570 (N_3570,N_14,N_1129);
and U3571 (N_3571,N_1443,N_2578);
nor U3572 (N_3572,N_1310,N_1938);
or U3573 (N_3573,N_714,N_2867);
or U3574 (N_3574,N_1487,N_2040);
and U3575 (N_3575,N_863,N_1041);
nand U3576 (N_3576,N_2818,N_1977);
nand U3577 (N_3577,N_2868,N_261);
or U3578 (N_3578,N_1586,N_2368);
nand U3579 (N_3579,N_1395,N_1572);
nor U3580 (N_3580,N_2322,N_1414);
or U3581 (N_3581,N_2211,N_2640);
xor U3582 (N_3582,N_792,N_2137);
or U3583 (N_3583,N_2288,N_2454);
and U3584 (N_3584,N_486,N_2392);
xor U3585 (N_3585,N_2767,N_659);
nand U3586 (N_3586,N_87,N_57);
nor U3587 (N_3587,N_2609,N_867);
and U3588 (N_3588,N_2752,N_2550);
or U3589 (N_3589,N_2678,N_2298);
or U3590 (N_3590,N_1617,N_1040);
nand U3591 (N_3591,N_2412,N_1663);
nand U3592 (N_3592,N_1895,N_2509);
or U3593 (N_3593,N_858,N_518);
or U3594 (N_3594,N_1730,N_677);
or U3595 (N_3595,N_2717,N_222);
or U3596 (N_3596,N_1763,N_1755);
nor U3597 (N_3597,N_544,N_921);
xnor U3598 (N_3598,N_543,N_1062);
nor U3599 (N_3599,N_1391,N_1255);
nand U3600 (N_3600,N_802,N_1161);
nor U3601 (N_3601,N_1900,N_1098);
or U3602 (N_3602,N_2904,N_571);
and U3603 (N_3603,N_92,N_1657);
nor U3604 (N_3604,N_2953,N_1975);
and U3605 (N_3605,N_1720,N_1236);
and U3606 (N_3606,N_1489,N_2791);
or U3607 (N_3607,N_1601,N_1513);
and U3608 (N_3608,N_2065,N_1729);
nand U3609 (N_3609,N_2542,N_2449);
nand U3610 (N_3610,N_282,N_2275);
nand U3611 (N_3611,N_197,N_2055);
nand U3612 (N_3612,N_1882,N_2571);
nor U3613 (N_3613,N_2806,N_1803);
or U3614 (N_3614,N_1112,N_1699);
and U3615 (N_3615,N_1939,N_2210);
or U3616 (N_3616,N_1459,N_2962);
nand U3617 (N_3617,N_1689,N_2792);
and U3618 (N_3618,N_581,N_2150);
xor U3619 (N_3619,N_1819,N_375);
nor U3620 (N_3620,N_253,N_976);
or U3621 (N_3621,N_2026,N_781);
nand U3622 (N_3622,N_2153,N_2163);
and U3623 (N_3623,N_2742,N_349);
and U3624 (N_3624,N_227,N_669);
or U3625 (N_3625,N_1121,N_2241);
nor U3626 (N_3626,N_2353,N_1229);
and U3627 (N_3627,N_2203,N_2965);
and U3628 (N_3628,N_864,N_2933);
and U3629 (N_3629,N_146,N_2815);
nand U3630 (N_3630,N_2936,N_2235);
and U3631 (N_3631,N_996,N_134);
nand U3632 (N_3632,N_2038,N_1788);
nand U3633 (N_3633,N_1157,N_1921);
or U3634 (N_3634,N_2339,N_2170);
nand U3635 (N_3635,N_547,N_1643);
or U3636 (N_3636,N_2902,N_1842);
xor U3637 (N_3637,N_268,N_2651);
xnor U3638 (N_3638,N_2314,N_2312);
nand U3639 (N_3639,N_2057,N_1786);
or U3640 (N_3640,N_2547,N_2912);
xnor U3641 (N_3641,N_346,N_72);
and U3642 (N_3642,N_2250,N_2489);
nand U3643 (N_3643,N_1477,N_506);
or U3644 (N_3644,N_727,N_2059);
or U3645 (N_3645,N_2483,N_2827);
nand U3646 (N_3646,N_400,N_2682);
or U3647 (N_3647,N_2108,N_769);
xor U3648 (N_3648,N_2087,N_1178);
or U3649 (N_3649,N_2718,N_2586);
or U3650 (N_3650,N_1701,N_768);
nor U3651 (N_3651,N_882,N_1800);
and U3652 (N_3652,N_1291,N_1578);
nand U3653 (N_3653,N_2481,N_1202);
and U3654 (N_3654,N_1575,N_602);
nor U3655 (N_3655,N_1324,N_1172);
or U3656 (N_3656,N_2915,N_74);
and U3657 (N_3657,N_2016,N_1910);
nor U3658 (N_3658,N_742,N_657);
and U3659 (N_3659,N_2118,N_1317);
nor U3660 (N_3660,N_1703,N_1321);
or U3661 (N_3661,N_904,N_1017);
and U3662 (N_3662,N_1507,N_2668);
xor U3663 (N_3663,N_2878,N_2109);
or U3664 (N_3664,N_1435,N_1990);
and U3665 (N_3665,N_1616,N_2989);
nor U3666 (N_3666,N_1003,N_939);
nor U3667 (N_3667,N_2145,N_62);
xnor U3668 (N_3668,N_626,N_614);
and U3669 (N_3669,N_1484,N_1640);
xor U3670 (N_3670,N_481,N_2576);
and U3671 (N_3671,N_834,N_2002);
xnor U3672 (N_3672,N_1854,N_717);
or U3673 (N_3673,N_1262,N_35);
nor U3674 (N_3674,N_1109,N_644);
and U3675 (N_3675,N_145,N_1495);
or U3676 (N_3676,N_298,N_1751);
nand U3677 (N_3677,N_2943,N_1634);
and U3678 (N_3678,N_1397,N_1588);
and U3679 (N_3679,N_2245,N_480);
or U3680 (N_3680,N_2364,N_817);
or U3681 (N_3681,N_2995,N_204);
or U3682 (N_3682,N_8,N_2830);
nand U3683 (N_3683,N_2987,N_1469);
or U3684 (N_3684,N_2749,N_1857);
and U3685 (N_3685,N_2217,N_2736);
nor U3686 (N_3686,N_1865,N_1893);
xnor U3687 (N_3687,N_1325,N_1499);
and U3688 (N_3688,N_2846,N_2098);
and U3689 (N_3689,N_1874,N_459);
nor U3690 (N_3690,N_40,N_1541);
and U3691 (N_3691,N_2920,N_441);
nor U3692 (N_3692,N_208,N_2615);
xnor U3693 (N_3693,N_2832,N_2218);
nor U3694 (N_3694,N_2318,N_1007);
nand U3695 (N_3695,N_2001,N_725);
and U3696 (N_3696,N_1777,N_2777);
nor U3697 (N_3697,N_1836,N_2152);
nand U3698 (N_3698,N_313,N_1970);
or U3699 (N_3699,N_1605,N_1075);
xor U3700 (N_3700,N_851,N_1953);
or U3701 (N_3701,N_2015,N_1144);
and U3702 (N_3702,N_2265,N_1824);
and U3703 (N_3703,N_2494,N_1378);
and U3704 (N_3704,N_1115,N_945);
or U3705 (N_3705,N_2324,N_2706);
nor U3706 (N_3706,N_866,N_10);
nand U3707 (N_3707,N_1795,N_2921);
nand U3708 (N_3708,N_1868,N_2557);
nor U3709 (N_3709,N_2937,N_1419);
nand U3710 (N_3710,N_2289,N_1709);
or U3711 (N_3711,N_2082,N_1638);
xor U3712 (N_3712,N_1,N_1887);
xor U3713 (N_3713,N_410,N_861);
and U3714 (N_3714,N_1622,N_1504);
nand U3715 (N_3715,N_2102,N_2238);
or U3716 (N_3716,N_1437,N_958);
nor U3717 (N_3717,N_681,N_2129);
or U3718 (N_3718,N_1944,N_770);
nand U3719 (N_3719,N_97,N_948);
or U3720 (N_3720,N_2826,N_1265);
nand U3721 (N_3721,N_1818,N_608);
or U3722 (N_3722,N_445,N_2690);
nor U3723 (N_3723,N_2122,N_421);
or U3724 (N_3724,N_484,N_1093);
and U3725 (N_3725,N_2007,N_1228);
xor U3726 (N_3726,N_804,N_1134);
nor U3727 (N_3727,N_1046,N_2534);
or U3728 (N_3728,N_2820,N_2186);
and U3729 (N_3729,N_1558,N_952);
nand U3730 (N_3730,N_1849,N_2164);
nor U3731 (N_3731,N_1957,N_1780);
nand U3732 (N_3732,N_26,N_850);
and U3733 (N_3733,N_1603,N_1626);
xnor U3734 (N_3734,N_2823,N_598);
nand U3735 (N_3735,N_1859,N_111);
nand U3736 (N_3736,N_1752,N_1256);
nor U3737 (N_3737,N_1188,N_1274);
or U3738 (N_3738,N_900,N_1850);
and U3739 (N_3739,N_2273,N_2415);
and U3740 (N_3740,N_1301,N_1441);
and U3741 (N_3741,N_515,N_1498);
or U3742 (N_3742,N_1220,N_166);
xnor U3743 (N_3743,N_2819,N_1375);
or U3744 (N_3744,N_1475,N_2467);
nor U3745 (N_3745,N_311,N_1890);
nor U3746 (N_3746,N_552,N_2758);
and U3747 (N_3747,N_1067,N_838);
and U3748 (N_3748,N_2366,N_2099);
and U3749 (N_3749,N_1002,N_1349);
and U3750 (N_3750,N_2607,N_1536);
nor U3751 (N_3751,N_1510,N_1532);
nor U3752 (N_3752,N_2172,N_2069);
and U3753 (N_3753,N_628,N_2009);
and U3754 (N_3754,N_507,N_2973);
or U3755 (N_3755,N_880,N_2344);
nand U3756 (N_3756,N_2115,N_2964);
nand U3757 (N_3757,N_147,N_1671);
and U3758 (N_3758,N_2680,N_1283);
nand U3759 (N_3759,N_2996,N_1642);
nand U3760 (N_3760,N_2496,N_2990);
and U3761 (N_3761,N_2610,N_1636);
or U3762 (N_3762,N_975,N_1765);
nor U3763 (N_3763,N_2799,N_2809);
nand U3764 (N_3764,N_2780,N_1608);
nand U3765 (N_3765,N_1880,N_1918);
and U3766 (N_3766,N_2460,N_1571);
nand U3767 (N_3767,N_1204,N_2092);
and U3768 (N_3768,N_732,N_690);
xor U3769 (N_3769,N_1545,N_917);
nor U3770 (N_3770,N_1552,N_810);
or U3771 (N_3771,N_2459,N_1945);
nor U3772 (N_3772,N_1016,N_207);
nand U3773 (N_3773,N_762,N_335);
or U3774 (N_3774,N_1923,N_2418);
and U3775 (N_3775,N_1750,N_2094);
or U3776 (N_3776,N_2470,N_2600);
xor U3777 (N_3777,N_816,N_2885);
nor U3778 (N_3778,N_1862,N_483);
nor U3779 (N_3779,N_1404,N_475);
or U3780 (N_3780,N_233,N_16);
and U3781 (N_3781,N_2954,N_1427);
or U3782 (N_3782,N_434,N_1610);
nand U3783 (N_3783,N_1481,N_2704);
or U3784 (N_3784,N_2663,N_1679);
xnor U3785 (N_3785,N_385,N_2213);
and U3786 (N_3786,N_327,N_1105);
nor U3787 (N_3787,N_2284,N_1492);
nor U3788 (N_3788,N_962,N_2021);
nand U3789 (N_3789,N_2755,N_1433);
or U3790 (N_3790,N_2537,N_2744);
nor U3791 (N_3791,N_2357,N_1806);
nor U3792 (N_3792,N_452,N_417);
or U3793 (N_3793,N_240,N_2438);
and U3794 (N_3794,N_1192,N_2446);
and U3795 (N_3795,N_2848,N_2515);
nand U3796 (N_3796,N_1082,N_2569);
and U3797 (N_3797,N_191,N_990);
and U3798 (N_3798,N_1179,N_1304);
or U3799 (N_3799,N_574,N_275);
and U3800 (N_3800,N_370,N_85);
nor U3801 (N_3801,N_1662,N_2450);
or U3802 (N_3802,N_2493,N_1899);
nor U3803 (N_3803,N_726,N_790);
nand U3804 (N_3804,N_2844,N_621);
or U3805 (N_3805,N_1099,N_2361);
nor U3806 (N_3806,N_1828,N_735);
nor U3807 (N_3807,N_1523,N_2097);
nand U3808 (N_3808,N_2390,N_881);
xor U3809 (N_3809,N_627,N_522);
nor U3810 (N_3810,N_2106,N_2257);
and U3811 (N_3811,N_2581,N_1253);
or U3812 (N_3812,N_1074,N_2410);
or U3813 (N_3813,N_2325,N_2306);
or U3814 (N_3814,N_1476,N_2748);
nor U3815 (N_3815,N_1286,N_276);
nand U3816 (N_3816,N_1186,N_25);
or U3817 (N_3817,N_141,N_709);
and U3818 (N_3818,N_3,N_1776);
and U3819 (N_3819,N_2670,N_494);
and U3820 (N_3820,N_88,N_474);
or U3821 (N_3821,N_428,N_2613);
and U3822 (N_3822,N_811,N_2627);
nand U3823 (N_3823,N_2377,N_1078);
nand U3824 (N_3824,N_2076,N_734);
xnor U3825 (N_3825,N_2400,N_1409);
and U3826 (N_3826,N_1423,N_2080);
xnor U3827 (N_3827,N_86,N_553);
and U3828 (N_3828,N_2047,N_2689);
or U3829 (N_3829,N_2394,N_2305);
and U3830 (N_3830,N_670,N_2739);
nor U3831 (N_3831,N_1072,N_2064);
nand U3832 (N_3832,N_2561,N_1907);
xnor U3833 (N_3833,N_1817,N_2028);
nor U3834 (N_3834,N_675,N_2142);
nand U3835 (N_3835,N_2126,N_315);
nor U3836 (N_3836,N_2342,N_1515);
or U3837 (N_3837,N_2445,N_2804);
nor U3838 (N_3838,N_513,N_296);
nand U3839 (N_3839,N_1966,N_1746);
or U3840 (N_3840,N_865,N_1010);
xor U3841 (N_3841,N_1876,N_995);
or U3842 (N_3842,N_1991,N_260);
nand U3843 (N_3843,N_1525,N_2468);
nand U3844 (N_3844,N_1371,N_2945);
and U3845 (N_3845,N_1359,N_2691);
nor U3846 (N_3846,N_986,N_956);
nand U3847 (N_3847,N_1486,N_1691);
and U3848 (N_3848,N_1386,N_2564);
and U3849 (N_3849,N_684,N_2206);
nor U3850 (N_3850,N_569,N_1059);
nand U3851 (N_3851,N_1149,N_2884);
xnor U3852 (N_3852,N_211,N_11);
and U3853 (N_3853,N_925,N_664);
nand U3854 (N_3854,N_243,N_2594);
nor U3855 (N_3855,N_502,N_2725);
or U3856 (N_3856,N_805,N_2616);
or U3857 (N_3857,N_2841,N_2518);
nand U3858 (N_3858,N_60,N_228);
nor U3859 (N_3859,N_2224,N_2271);
and U3860 (N_3860,N_723,N_1084);
and U3861 (N_3861,N_408,N_831);
nand U3862 (N_3862,N_686,N_220);
or U3863 (N_3863,N_1269,N_2138);
nor U3864 (N_3864,N_1290,N_568);
or U3865 (N_3865,N_389,N_2154);
nand U3866 (N_3866,N_138,N_1967);
and U3867 (N_3867,N_1951,N_2233);
nor U3868 (N_3868,N_2917,N_719);
nand U3869 (N_3869,N_2464,N_1479);
or U3870 (N_3870,N_718,N_1468);
nor U3871 (N_3871,N_1583,N_22);
nor U3872 (N_3872,N_679,N_1131);
nand U3873 (N_3873,N_1733,N_418);
or U3874 (N_3874,N_64,N_200);
nor U3875 (N_3875,N_2139,N_1011);
or U3876 (N_3876,N_129,N_528);
and U3877 (N_3877,N_1704,N_1706);
and U3878 (N_3878,N_122,N_2501);
nand U3879 (N_3879,N_730,N_81);
or U3880 (N_3880,N_305,N_1823);
or U3881 (N_3881,N_1960,N_1595);
nand U3882 (N_3882,N_673,N_2788);
nand U3883 (N_3883,N_929,N_594);
or U3884 (N_3884,N_1538,N_2183);
xor U3885 (N_3885,N_954,N_1104);
nor U3886 (N_3886,N_451,N_639);
and U3887 (N_3887,N_1569,N_2354);
and U3888 (N_3888,N_300,N_1727);
and U3889 (N_3889,N_2416,N_1288);
nor U3890 (N_3890,N_1152,N_1450);
nor U3891 (N_3891,N_566,N_2525);
and U3892 (N_3892,N_966,N_1998);
nor U3893 (N_3893,N_236,N_1197);
or U3894 (N_3894,N_1606,N_1049);
or U3895 (N_3895,N_2051,N_559);
or U3896 (N_3896,N_2431,N_2447);
nand U3897 (N_3897,N_2639,N_923);
nand U3898 (N_3898,N_1284,N_2237);
nand U3899 (N_3899,N_2665,N_871);
nand U3900 (N_3900,N_2133,N_2757);
or U3901 (N_3901,N_635,N_1107);
nand U3902 (N_3902,N_199,N_1023);
and U3903 (N_3903,N_1904,N_2263);
or U3904 (N_3904,N_104,N_554);
and U3905 (N_3905,N_855,N_1374);
nor U3906 (N_3906,N_1044,N_2940);
nand U3907 (N_3907,N_73,N_1156);
xnor U3908 (N_3908,N_672,N_248);
nor U3909 (N_3909,N_2778,N_2653);
xnor U3910 (N_3910,N_701,N_1947);
nor U3911 (N_3911,N_830,N_694);
and U3912 (N_3912,N_888,N_1135);
or U3913 (N_3913,N_2891,N_526);
or U3914 (N_3914,N_1318,N_733);
or U3915 (N_3915,N_2839,N_2713);
or U3916 (N_3916,N_2155,N_2702);
and U3917 (N_3917,N_2389,N_859);
nand U3918 (N_3918,N_2068,N_2283);
xor U3919 (N_3919,N_1522,N_1154);
xor U3920 (N_3920,N_1060,N_371);
nor U3921 (N_3921,N_753,N_2783);
nand U3922 (N_3922,N_570,N_2101);
nor U3923 (N_3923,N_1840,N_692);
nand U3924 (N_3924,N_406,N_1553);
xor U3925 (N_3925,N_1766,N_1929);
and U3926 (N_3926,N_2005,N_334);
and U3927 (N_3927,N_1114,N_196);
or U3928 (N_3928,N_1801,N_1614);
and U3929 (N_3929,N_1254,N_1221);
or U3930 (N_3930,N_2526,N_2519);
or U3931 (N_3931,N_2053,N_151);
nor U3932 (N_3932,N_1885,N_2908);
nand U3933 (N_3933,N_1982,N_1632);
and U3934 (N_3934,N_1266,N_2030);
nand U3935 (N_3935,N_2223,N_183);
or U3936 (N_3936,N_198,N_2504);
nor U3937 (N_3937,N_1302,N_2379);
nand U3938 (N_3938,N_632,N_2134);
nor U3939 (N_3939,N_2385,N_1792);
and U3940 (N_3940,N_258,N_2529);
xor U3941 (N_3941,N_555,N_1869);
nor U3942 (N_3942,N_382,N_179);
nor U3943 (N_3943,N_521,N_2697);
nor U3944 (N_3944,N_1088,N_1530);
xnor U3945 (N_3945,N_1629,N_1362);
nand U3946 (N_3946,N_2169,N_2495);
nor U3947 (N_3947,N_1927,N_2345);
nand U3948 (N_3948,N_776,N_577);
nand U3949 (N_3949,N_2675,N_2419);
nor U3950 (N_3950,N_1406,N_355);
nand U3951 (N_3951,N_832,N_666);
or U3952 (N_3952,N_2976,N_2171);
or U3953 (N_3953,N_2929,N_353);
xor U3954 (N_3954,N_1889,N_2559);
or U3955 (N_3955,N_1056,N_2160);
nand U3956 (N_3956,N_1871,N_2790);
or U3957 (N_3957,N_2955,N_182);
or U3958 (N_3958,N_1282,N_214);
xnor U3959 (N_3959,N_2456,N_1342);
nand U3960 (N_3960,N_1400,N_873);
and U3961 (N_3961,N_1297,N_2161);
nor U3962 (N_3962,N_601,N_1183);
nor U3963 (N_3963,N_2078,N_1635);
nand U3964 (N_3964,N_1773,N_1347);
or U3965 (N_3965,N_468,N_68);
or U3966 (N_3966,N_2383,N_676);
xnor U3967 (N_3967,N_1922,N_423);
or U3968 (N_3968,N_2299,N_2498);
or U3969 (N_3969,N_1473,N_1309);
xnor U3970 (N_3970,N_1137,N_2948);
nand U3971 (N_3971,N_1471,N_2621);
or U3972 (N_3972,N_2517,N_378);
or U3973 (N_3973,N_2294,N_540);
nor U3974 (N_3974,N_1716,N_562);
nor U3975 (N_3975,N_1722,N_950);
nor U3976 (N_3976,N_1209,N_1401);
nor U3977 (N_3977,N_2593,N_724);
or U3978 (N_3978,N_695,N_1080);
xor U3979 (N_3979,N_2683,N_1529);
or U3980 (N_3980,N_1740,N_2315);
or U3981 (N_3981,N_2864,N_707);
nand U3982 (N_3982,N_177,N_2086);
nor U3983 (N_3983,N_185,N_1173);
nand U3984 (N_3984,N_320,N_1574);
nand U3985 (N_3985,N_1879,N_1968);
or U3986 (N_3986,N_102,N_2688);
nand U3987 (N_3987,N_2417,N_2735);
and U3988 (N_3988,N_2147,N_1735);
xor U3989 (N_3989,N_1364,N_978);
and U3990 (N_3990,N_2232,N_2010);
nor U3991 (N_3991,N_1542,N_1319);
nand U3992 (N_3992,N_80,N_596);
nor U3993 (N_3993,N_2880,N_2441);
or U3994 (N_3994,N_304,N_665);
or U3995 (N_3995,N_2575,N_1858);
or U3996 (N_3996,N_915,N_2654);
and U3997 (N_3997,N_456,N_70);
and U3998 (N_3998,N_2491,N_2733);
nor U3999 (N_3999,N_2277,N_2351);
or U4000 (N_4000,N_2240,N_1224);
or U4001 (N_4001,N_1688,N_351);
nand U4002 (N_4002,N_1032,N_824);
nand U4003 (N_4003,N_345,N_1233);
nand U4004 (N_4004,N_2374,N_2254);
nand U4005 (N_4005,N_2266,N_201);
nand U4006 (N_4006,N_1079,N_1566);
nor U4007 (N_4007,N_1396,N_1388);
or U4008 (N_4008,N_1272,N_1581);
nor U4009 (N_4009,N_774,N_2599);
nand U4010 (N_4010,N_1742,N_985);
or U4011 (N_4011,N_1216,N_2782);
or U4012 (N_4012,N_500,N_2681);
xor U4013 (N_4013,N_2341,N_2960);
nand U4014 (N_4014,N_994,N_1959);
and U4015 (N_4015,N_144,N_1399);
or U4016 (N_4016,N_2730,N_1992);
or U4017 (N_4017,N_1024,N_2176);
and U4018 (N_4018,N_2899,N_247);
or U4019 (N_4019,N_1306,N_991);
or U4020 (N_4020,N_2326,N_1081);
nand U4021 (N_4021,N_1754,N_1714);
or U4022 (N_4022,N_2808,N_2004);
xor U4023 (N_4023,N_2584,N_843);
nand U4024 (N_4024,N_689,N_1462);
nor U4025 (N_4025,N_1972,N_2466);
nor U4026 (N_4026,N_1296,N_1778);
nor U4027 (N_4027,N_9,N_2056);
xor U4028 (N_4028,N_1665,N_2023);
nand U4029 (N_4029,N_388,N_1631);
or U4030 (N_4030,N_1661,N_2853);
nor U4031 (N_4031,N_303,N_2980);
or U4032 (N_4032,N_2728,N_2549);
and U4033 (N_4033,N_2516,N_1351);
nand U4034 (N_4034,N_432,N_2276);
and U4035 (N_4035,N_633,N_1644);
nand U4036 (N_4036,N_981,N_1323);
nand U4037 (N_4037,N_998,N_2851);
or U4038 (N_4038,N_1676,N_2906);
and U4039 (N_4039,N_127,N_1398);
or U4040 (N_4040,N_415,N_605);
or U4041 (N_4041,N_1472,N_796);
nor U4042 (N_4042,N_1025,N_1071);
nand U4043 (N_4043,N_1607,N_108);
nand U4044 (N_4044,N_1519,N_465);
and U4045 (N_4045,N_120,N_764);
nor U4046 (N_4046,N_2166,N_499);
or U4047 (N_4047,N_2095,N_2);
nand U4048 (N_4048,N_637,N_1524);
nor U4049 (N_4049,N_638,N_874);
nor U4050 (N_4050,N_2331,N_112);
or U4051 (N_4051,N_376,N_1557);
or U4052 (N_4052,N_2776,N_1848);
or U4053 (N_4053,N_560,N_1700);
nor U4054 (N_4054,N_19,N_2323);
nor U4055 (N_4055,N_471,N_1263);
nand U4056 (N_4056,N_1772,N_783);
nor U4057 (N_4057,N_46,N_1368);
and U4058 (N_4058,N_1356,N_1799);
and U4059 (N_4059,N_1748,N_1355);
nor U4060 (N_4060,N_2974,N_2189);
and U4061 (N_4061,N_195,N_2309);
nor U4062 (N_4062,N_2334,N_2029);
and U4063 (N_4063,N_1599,N_89);
or U4064 (N_4064,N_1501,N_391);
nor U4065 (N_4065,N_84,N_1051);
xor U4066 (N_4066,N_1540,N_778);
and U4067 (N_4067,N_2208,N_1205);
or U4068 (N_4068,N_398,N_1639);
nand U4069 (N_4069,N_890,N_251);
nor U4070 (N_4070,N_283,N_1320);
nor U4071 (N_4071,N_2256,N_139);
and U4072 (N_4072,N_1430,N_1285);
and U4073 (N_4073,N_2802,N_2966);
nand U4074 (N_4074,N_2425,N_2404);
xnor U4075 (N_4075,N_1148,N_1677);
nor U4076 (N_4076,N_234,N_440);
or U4077 (N_4077,N_109,N_49);
nand U4078 (N_4078,N_1774,N_2157);
and U4079 (N_4079,N_2457,N_612);
nand U4080 (N_4080,N_318,N_501);
nor U4081 (N_4081,N_42,N_1641);
nor U4082 (N_4082,N_2720,N_2633);
and U4083 (N_4083,N_176,N_1208);
and U4084 (N_4084,N_2258,N_2058);
and U4085 (N_4085,N_2753,N_957);
nor U4086 (N_4086,N_2054,N_2198);
and U4087 (N_4087,N_301,N_1658);
or U4088 (N_4088,N_809,N_2924);
or U4089 (N_4089,N_132,N_1305);
or U4090 (N_4090,N_2991,N_2993);
and U4091 (N_4091,N_1785,N_713);
and U4092 (N_4092,N_898,N_1808);
nor U4093 (N_4093,N_1747,N_1226);
or U4094 (N_4094,N_430,N_520);
and U4095 (N_4095,N_2694,N_344);
nor U4096 (N_4096,N_789,N_582);
nand U4097 (N_4097,N_2531,N_624);
or U4098 (N_4098,N_2136,N_747);
nor U4099 (N_4099,N_447,N_2512);
xor U4100 (N_4100,N_1901,N_2128);
or U4101 (N_4101,N_359,N_206);
nor U4102 (N_4102,N_416,N_2913);
nand U4103 (N_4103,N_512,N_704);
nand U4104 (N_4104,N_1199,N_2676);
and U4105 (N_4105,N_2079,N_2350);
xnor U4106 (N_4106,N_821,N_2626);
or U4107 (N_4107,N_314,N_1667);
nand U4108 (N_4108,N_2140,N_2540);
or U4109 (N_4109,N_2863,N_616);
and U4110 (N_4110,N_1344,N_1132);
and U4111 (N_4111,N_2746,N_2355);
and U4112 (N_4112,N_439,N_2882);
and U4113 (N_4113,N_1546,N_1916);
or U4114 (N_4114,N_503,N_340);
or U4115 (N_4115,N_951,N_743);
and U4116 (N_4116,N_648,N_586);
xor U4117 (N_4117,N_1027,N_786);
nor U4118 (N_4118,N_61,N_2887);
nand U4119 (N_4119,N_2439,N_2376);
or U4120 (N_4120,N_2985,N_5);
nand U4121 (N_4121,N_2977,N_1827);
or U4122 (N_4122,N_1584,N_2765);
or U4123 (N_4123,N_595,N_1814);
nor U4124 (N_4124,N_2838,N_791);
nor U4125 (N_4125,N_2280,N_2507);
and U4126 (N_4126,N_1039,N_1298);
and U4127 (N_4127,N_2180,N_2530);
nand U4128 (N_4128,N_2032,N_2144);
or U4129 (N_4129,N_2997,N_2292);
xor U4130 (N_4130,N_1231,N_965);
xnor U4131 (N_4131,N_231,N_1783);
nand U4132 (N_4132,N_2807,N_155);
nand U4133 (N_4133,N_1526,N_826);
xor U4134 (N_4134,N_940,N_178);
or U4135 (N_4135,N_2769,N_2824);
and U4136 (N_4136,N_2403,N_1313);
nand U4137 (N_4137,N_1518,N_755);
xor U4138 (N_4138,N_1925,N_1055);
and U4139 (N_4139,N_1190,N_436);
nand U4140 (N_4140,N_2243,N_557);
nand U4141 (N_4141,N_2858,N_156);
or U4142 (N_4142,N_1962,N_2971);
nor U4143 (N_4143,N_1881,N_593);
or U4144 (N_4144,N_256,N_1837);
nor U4145 (N_4145,N_1660,N_2251);
nor U4146 (N_4146,N_2052,N_2760);
nor U4147 (N_4147,N_784,N_399);
or U4148 (N_4148,N_2729,N_1568);
nand U4149 (N_4149,N_2408,N_2629);
or U4150 (N_4150,N_1997,N_845);
or U4151 (N_4151,N_1076,N_1741);
xnor U4152 (N_4152,N_1187,N_54);
nor U4153 (N_4153,N_2901,N_1198);
or U4154 (N_4154,N_1311,N_623);
xnor U4155 (N_4155,N_2135,N_2179);
and U4156 (N_4156,N_333,N_205);
or U4157 (N_4157,N_1207,N_1839);
nor U4158 (N_4158,N_1533,N_2684);
nand U4159 (N_4159,N_926,N_2185);
nand U4160 (N_4160,N_1567,N_697);
nand U4161 (N_4161,N_2905,N_1273);
nand U4162 (N_4162,N_30,N_2658);
nor U4163 (N_4163,N_154,N_1845);
and U4164 (N_4164,N_2963,N_1794);
and U4165 (N_4165,N_2230,N_1217);
or U4166 (N_4166,N_980,N_738);
or U4167 (N_4167,N_2632,N_1650);
and U4168 (N_4168,N_840,N_1258);
nand U4169 (N_4169,N_797,N_137);
nand U4170 (N_4170,N_1160,N_545);
nand U4171 (N_4171,N_2123,N_1077);
nor U4172 (N_4172,N_319,N_1415);
nand U4173 (N_4173,N_53,N_71);
nand U4174 (N_4174,N_2538,N_403);
nor U4175 (N_4175,N_1411,N_1539);
or U4176 (N_4176,N_2829,N_1511);
xnor U4177 (N_4177,N_83,N_1241);
nor U4178 (N_4178,N_1775,N_2046);
or U4179 (N_4179,N_712,N_2006);
and U4180 (N_4180,N_2424,N_1358);
nor U4181 (N_4181,N_32,N_2646);
nand U4182 (N_4182,N_534,N_2992);
nor U4183 (N_4183,N_2797,N_2473);
and U4184 (N_4184,N_2649,N_2297);
nor U4185 (N_4185,N_2335,N_2842);
or U4186 (N_4186,N_2577,N_533);
nand U4187 (N_4187,N_1019,N_1013);
or U4188 (N_4188,N_1590,N_294);
nand U4189 (N_4189,N_2287,N_2774);
nor U4190 (N_4190,N_2475,N_2619);
nor U4191 (N_4191,N_36,N_1095);
and U4192 (N_4192,N_2715,N_2427);
nand U4193 (N_4193,N_1934,N_387);
nor U4194 (N_4194,N_377,N_1239);
nor U4195 (N_4195,N_152,N_7);
nand U4196 (N_4196,N_2695,N_1506);
nand U4197 (N_4197,N_1063,N_479);
nand U4198 (N_4198,N_1271,N_2611);
or U4199 (N_4199,N_746,N_2024);
or U4200 (N_4200,N_2143,N_1913);
nor U4201 (N_4201,N_1213,N_2204);
nand U4202 (N_4202,N_2585,N_2562);
or U4203 (N_4203,N_31,N_660);
nand U4204 (N_4204,N_1861,N_2724);
or U4205 (N_4205,N_63,N_849);
nor U4206 (N_4206,N_422,N_2011);
nand U4207 (N_4207,N_1432,N_290);
or U4208 (N_4208,N_508,N_2800);
nand U4209 (N_4209,N_1280,N_883);
and U4210 (N_4210,N_1436,N_274);
and U4211 (N_4211,N_2225,N_1089);
or U4212 (N_4212,N_2317,N_629);
or U4213 (N_4213,N_2045,N_487);
and U4214 (N_4214,N_17,N_2034);
nand U4215 (N_4215,N_1006,N_885);
and U4216 (N_4216,N_1181,N_1108);
nor U4217 (N_4217,N_955,N_2285);
and U4218 (N_4218,N_685,N_1761);
and U4219 (N_4219,N_2282,N_2311);
or U4220 (N_4220,N_2215,N_259);
or U4221 (N_4221,N_729,N_1014);
nand U4222 (N_4222,N_2650,N_782);
or U4223 (N_4223,N_82,N_2452);
and U4224 (N_4224,N_1821,N_1470);
nand U4225 (N_4225,N_2617,N_1246);
nor U4226 (N_4226,N_1646,N_210);
nor U4227 (N_4227,N_1125,N_788);
nor U4228 (N_4228,N_2624,N_772);
and U4229 (N_4229,N_1813,N_760);
and U4230 (N_4230,N_1214,N_390);
or U4231 (N_4231,N_1465,N_171);
nor U4232 (N_4232,N_1976,N_124);
or U4233 (N_4233,N_1175,N_1279);
or U4234 (N_4234,N_1738,N_893);
nor U4235 (N_4235,N_462,N_1235);
nor U4236 (N_4236,N_143,N_1782);
and U4237 (N_4237,N_2722,N_2222);
xor U4238 (N_4238,N_2043,N_1935);
nand U4239 (N_4239,N_2789,N_1952);
nor U4240 (N_4240,N_877,N_2833);
nand U4241 (N_4241,N_1715,N_41);
nand U4242 (N_4242,N_6,N_2423);
nand U4243 (N_4243,N_1816,N_1494);
or U4244 (N_4244,N_288,N_820);
or U4245 (N_4245,N_550,N_1117);
nor U4246 (N_4246,N_2659,N_2938);
nor U4247 (N_4247,N_405,N_1596);
nand U4248 (N_4248,N_78,N_793);
xor U4249 (N_4249,N_607,N_250);
or U4250 (N_4250,N_272,N_1696);
nand U4251 (N_4251,N_2606,N_1455);
and U4252 (N_4252,N_338,N_1124);
and U4253 (N_4253,N_1946,N_656);
and U4254 (N_4254,N_1001,N_1083);
or U4255 (N_4255,N_968,N_38);
and U4256 (N_4256,N_2370,N_1609);
xnor U4257 (N_4257,N_869,N_2443);
or U4258 (N_4258,N_325,N_1139);
and U4259 (N_4259,N_1257,N_1508);
nand U4260 (N_4260,N_889,N_2879);
nor U4261 (N_4261,N_2396,N_2405);
nand U4262 (N_4262,N_1000,N_761);
or U4263 (N_4263,N_892,N_1732);
nand U4264 (N_4264,N_157,N_947);
nor U4265 (N_4265,N_44,N_2816);
xor U4266 (N_4266,N_2811,N_116);
and U4267 (N_4267,N_2511,N_2401);
or U4268 (N_4268,N_1505,N_2558);
nand U4269 (N_4269,N_1517,N_2269);
or U4270 (N_4270,N_1385,N_2894);
and U4271 (N_4271,N_1264,N_1989);
or U4272 (N_4272,N_1167,N_1215);
nand U4273 (N_4273,N_655,N_1930);
or U4274 (N_4274,N_1194,N_18);
or U4275 (N_4275,N_2279,N_478);
nor U4276 (N_4276,N_953,N_1270);
and U4277 (N_4277,N_269,N_217);
or U4278 (N_4278,N_153,N_2781);
nor U4279 (N_4279,N_24,N_2556);
and U4280 (N_4280,N_1674,N_2202);
and U4281 (N_4281,N_558,N_514);
nor U4282 (N_4282,N_2605,N_1267);
or U4283 (N_4283,N_469,N_1758);
xnor U4284 (N_4284,N_2388,N_691);
nand U4285 (N_4285,N_1503,N_1768);
nand U4286 (N_4286,N_463,N_2104);
and U4287 (N_4287,N_2835,N_1734);
nand U4288 (N_4288,N_1240,N_916);
and U4289 (N_4289,N_1943,N_2072);
and U4290 (N_4290,N_347,N_187);
nand U4291 (N_4291,N_1891,N_1033);
nand U4292 (N_4292,N_1054,N_2367);
nand U4293 (N_4293,N_1914,N_773);
and U4294 (N_4294,N_779,N_2671);
or U4295 (N_4295,N_1681,N_1294);
nor U4296 (N_4296,N_2614,N_28);
nor U4297 (N_4297,N_496,N_2420);
and U4298 (N_4298,N_1762,N_1980);
nand U4299 (N_4299,N_1363,N_2008);
and U4300 (N_4300,N_1328,N_705);
or U4301 (N_4301,N_281,N_2661);
nor U4302 (N_4302,N_1377,N_1884);
nand U4303 (N_4303,N_983,N_343);
or U4304 (N_4304,N_1367,N_1009);
nor U4305 (N_4305,N_576,N_1018);
and U4306 (N_4306,N_2190,N_2484);
or U4307 (N_4307,N_905,N_2896);
nand U4308 (N_4308,N_181,N_2947);
nand U4309 (N_4309,N_2642,N_630);
nor U4310 (N_4310,N_505,N_1087);
nand U4311 (N_4311,N_930,N_1670);
and U4312 (N_4312,N_477,N_1474);
nand U4313 (N_4313,N_1141,N_1086);
or U4314 (N_4314,N_2910,N_404);
or U4315 (N_4315,N_2698,N_2261);
or U4316 (N_4316,N_2444,N_763);
or U4317 (N_4317,N_2499,N_34);
nor U4318 (N_4318,N_798,N_1979);
nor U4319 (N_4319,N_1942,N_2911);
nand U4320 (N_4320,N_2381,N_2692);
or U4321 (N_4321,N_2861,N_2635);
nand U4322 (N_4322,N_2961,N_2437);
nand U4323 (N_4323,N_2485,N_1334);
or U4324 (N_4324,N_95,N_822);
and U4325 (N_4325,N_530,N_2813);
and U4326 (N_4326,N_56,N_2330);
nand U4327 (N_4327,N_457,N_2784);
nor U4328 (N_4328,N_2272,N_2859);
xor U4329 (N_4329,N_2521,N_1833);
xor U4330 (N_4330,N_2244,N_2591);
or U4331 (N_4331,N_1110,N_1516);
or U4332 (N_4332,N_2972,N_785);
and U4333 (N_4333,N_671,N_848);
nand U4334 (N_4334,N_2112,N_2131);
nor U4335 (N_4335,N_175,N_358);
xor U4336 (N_4336,N_2226,N_383);
xor U4337 (N_4337,N_542,N_2935);
nand U4338 (N_4338,N_2391,N_460);
nor U4339 (N_4339,N_2291,N_615);
and U4340 (N_4340,N_2998,N_2239);
or U4341 (N_4341,N_1184,N_2319);
nand U4342 (N_4342,N_454,N_827);
and U4343 (N_4343,N_1986,N_96);
and U4344 (N_4344,N_1926,N_749);
nand U4345 (N_4345,N_825,N_1383);
or U4346 (N_4346,N_2687,N_1150);
xor U4347 (N_4347,N_1645,N_2603);
nand U4348 (N_4348,N_1556,N_2950);
or U4349 (N_4349,N_2130,N_1633);
or U4350 (N_4350,N_1413,N_1958);
xnor U4351 (N_4351,N_332,N_600);
or U4352 (N_4352,N_1618,N_2703);
or U4353 (N_4353,N_1248,N_1225);
nor U4354 (N_4354,N_2959,N_148);
nand U4355 (N_4355,N_226,N_297);
or U4356 (N_4356,N_1026,N_2794);
or U4357 (N_4357,N_2583,N_2674);
nand U4358 (N_4358,N_1130,N_2358);
nand U4359 (N_4359,N_1933,N_2700);
or U4360 (N_4360,N_973,N_835);
nand U4361 (N_4361,N_814,N_362);
nor U4362 (N_4362,N_2352,N_2371);
nor U4363 (N_4363,N_402,N_2768);
and U4364 (N_4364,N_1937,N_490);
xor U4365 (N_4365,N_646,N_1407);
nand U4366 (N_4366,N_230,N_2093);
or U4367 (N_4367,N_1580,N_2066);
and U4368 (N_4368,N_2958,N_2573);
xor U4369 (N_4369,N_2952,N_2888);
nand U4370 (N_4370,N_2084,N_1560);
or U4371 (N_4371,N_1559,N_2631);
or U4372 (N_4372,N_2151,N_2175);
or U4373 (N_4373,N_2336,N_698);
xor U4374 (N_4374,N_1883,N_879);
or U4375 (N_4375,N_118,N_1384);
and U4376 (N_4376,N_488,N_13);
or U4377 (N_4377,N_284,N_1189);
and U4378 (N_4378,N_1445,N_1570);
nor U4379 (N_4379,N_1387,N_2167);
nor U4380 (N_4380,N_591,N_1162);
or U4381 (N_4381,N_2574,N_2027);
and U4382 (N_4382,N_2174,N_2090);
or U4383 (N_4383,N_752,N_2875);
and U4384 (N_4384,N_538,N_823);
or U4385 (N_4385,N_2362,N_1810);
xnor U4386 (N_4386,N_1126,N_813);
nand U4387 (N_4387,N_1829,N_2536);
nand U4388 (N_4388,N_795,N_1604);
or U4389 (N_4389,N_682,N_720);
xor U4390 (N_4390,N_2983,N_2117);
nor U4391 (N_4391,N_2497,N_2502);
nor U4392 (N_4392,N_270,N_1983);
nor U4393 (N_4393,N_2563,N_2205);
and U4394 (N_4394,N_476,N_588);
and U4395 (N_4395,N_1969,N_1769);
or U4396 (N_4396,N_2601,N_942);
and U4397 (N_4397,N_2761,N_2979);
nor U4398 (N_4398,N_2793,N_1322);
xnor U4399 (N_4399,N_1146,N_2666);
nand U4400 (N_4400,N_173,N_337);
nand U4401 (N_4401,N_1551,N_1843);
and U4402 (N_4402,N_2414,N_539);
nand U4403 (N_4403,N_1357,N_1680);
and U4404 (N_4404,N_1376,N_537);
or U4405 (N_4405,N_1771,N_39);
nor U4406 (N_4406,N_1624,N_1424);
nand U4407 (N_4407,N_2898,N_1232);
nand U4408 (N_4408,N_392,N_1390);
and U4409 (N_4409,N_2453,N_1276);
and U4410 (N_4410,N_2836,N_2857);
and U4411 (N_4411,N_706,N_1360);
nand U4412 (N_4412,N_401,N_1853);
or U4413 (N_4413,N_2260,N_1020);
nor U4414 (N_4414,N_489,N_1565);
and U4415 (N_4415,N_1237,N_2409);
and U4416 (N_4416,N_587,N_167);
nand U4417 (N_4417,N_1345,N_2373);
nand U4418 (N_4418,N_2840,N_249);
and U4419 (N_4419,N_2018,N_2555);
nor U4420 (N_4420,N_2421,N_1133);
nand U4421 (N_4421,N_443,N_1561);
or U4422 (N_4422,N_374,N_407);
nand U4423 (N_4423,N_2472,N_1394);
nor U4424 (N_4424,N_2944,N_1669);
and U4425 (N_4425,N_896,N_2756);
nor U4426 (N_4426,N_1277,N_2406);
nor U4427 (N_4427,N_852,N_485);
nand U4428 (N_4428,N_1166,N_932);
nand U4429 (N_4429,N_1961,N_737);
and U4430 (N_4430,N_2647,N_1331);
and U4431 (N_4431,N_2337,N_2165);
or U4432 (N_4432,N_1449,N_658);
or U4433 (N_4433,N_899,N_2316);
or U4434 (N_4434,N_1815,N_517);
nor U4435 (N_4435,N_1308,N_2191);
and U4436 (N_4436,N_2589,N_2847);
or U4437 (N_4437,N_1620,N_2770);
and U4438 (N_4438,N_1630,N_1528);
and U4439 (N_4439,N_1250,N_2662);
and U4440 (N_4440,N_1717,N_373);
or U4441 (N_4441,N_2070,N_2333);
nand U4442 (N_4442,N_1069,N_1206);
or U4443 (N_4443,N_1864,N_1903);
nand U4444 (N_4444,N_1898,N_1675);
nor U4445 (N_4445,N_2548,N_1537);
and U4446 (N_4446,N_1234,N_583);
xnor U4447 (N_4447,N_2545,N_384);
xnor U4448 (N_4448,N_2000,N_1464);
nor U4449 (N_4449,N_906,N_1021);
or U4450 (N_4450,N_2643,N_1045);
nand U4451 (N_4451,N_2978,N_1463);
or U4452 (N_4452,N_2513,N_1145);
nand U4453 (N_4453,N_394,N_2031);
xnor U4454 (N_4454,N_101,N_66);
and U4455 (N_4455,N_58,N_2685);
or U4456 (N_4456,N_1123,N_2699);
and U4457 (N_4457,N_1664,N_1352);
nand U4458 (N_4458,N_2889,N_312);
or U4459 (N_4459,N_1169,N_458);
or U4460 (N_4460,N_1029,N_912);
nand U4461 (N_4461,N_876,N_1037);
or U4462 (N_4462,N_136,N_366);
xnor U4463 (N_4463,N_943,N_2304);
nor U4464 (N_4464,N_381,N_131);
nand U4465 (N_4465,N_1520,N_2461);
nand U4466 (N_4466,N_918,N_618);
nand U4467 (N_4467,N_1512,N_936);
and U4468 (N_4468,N_1613,N_613);
nor U4469 (N_4469,N_2579,N_2623);
xor U4470 (N_4470,N_308,N_2707);
nor U4471 (N_4471,N_2876,N_1694);
xor U4472 (N_4472,N_2897,N_1457);
nor U4473 (N_4473,N_1295,N_2785);
xor U4474 (N_4474,N_2212,N_1176);
and U4475 (N_4475,N_1543,N_516);
nor U4476 (N_4476,N_636,N_949);
and U4477 (N_4477,N_1338,N_2673);
and U4478 (N_4478,N_302,N_1336);
nor U4479 (N_4479,N_1535,N_1592);
nand U4480 (N_4480,N_2301,N_1985);
xnor U4481 (N_4481,N_1106,N_678);
or U4482 (N_4482,N_1784,N_2119);
nand U4483 (N_4483,N_680,N_2252);
nand U4484 (N_4484,N_442,N_2071);
nor U4485 (N_4485,N_158,N_310);
and U4486 (N_4486,N_819,N_2399);
or U4487 (N_4487,N_235,N_466);
nand U4488 (N_4488,N_2701,N_1329);
nor U4489 (N_4489,N_1170,N_2608);
or U4490 (N_4490,N_492,N_1673);
or U4491 (N_4491,N_2994,N_573);
and U4492 (N_4492,N_369,N_1737);
xnor U4493 (N_4493,N_2595,N_1791);
nor U4494 (N_4494,N_2923,N_237);
nand U4495 (N_4495,N_979,N_2523);
and U4496 (N_4496,N_93,N_27);
nor U4497 (N_4497,N_2149,N_2803);
nand U4498 (N_4498,N_149,N_2580);
and U4499 (N_4499,N_37,N_1446);
xor U4500 (N_4500,N_2732,N_1841);
and U4501 (N_4501,N_210,N_293);
nand U4502 (N_4502,N_1766,N_1136);
or U4503 (N_4503,N_2393,N_1637);
xnor U4504 (N_4504,N_287,N_957);
and U4505 (N_4505,N_1287,N_2520);
or U4506 (N_4506,N_1975,N_1541);
or U4507 (N_4507,N_38,N_771);
or U4508 (N_4508,N_1863,N_2355);
nor U4509 (N_4509,N_1,N_625);
or U4510 (N_4510,N_612,N_2171);
nor U4511 (N_4511,N_343,N_1512);
nor U4512 (N_4512,N_1907,N_247);
nor U4513 (N_4513,N_2105,N_2104);
nand U4514 (N_4514,N_1681,N_916);
nor U4515 (N_4515,N_79,N_1329);
xor U4516 (N_4516,N_1475,N_1068);
and U4517 (N_4517,N_2235,N_1480);
nand U4518 (N_4518,N_2249,N_1875);
nor U4519 (N_4519,N_1004,N_1575);
or U4520 (N_4520,N_2174,N_1498);
nand U4521 (N_4521,N_1432,N_1079);
or U4522 (N_4522,N_750,N_1508);
nand U4523 (N_4523,N_2835,N_621);
or U4524 (N_4524,N_2451,N_622);
nor U4525 (N_4525,N_2888,N_2388);
nand U4526 (N_4526,N_673,N_2085);
and U4527 (N_4527,N_1671,N_2502);
and U4528 (N_4528,N_2438,N_2891);
xnor U4529 (N_4529,N_2771,N_1676);
xor U4530 (N_4530,N_2921,N_2419);
and U4531 (N_4531,N_1377,N_83);
and U4532 (N_4532,N_994,N_1515);
and U4533 (N_4533,N_604,N_2041);
xor U4534 (N_4534,N_2372,N_2044);
xor U4535 (N_4535,N_1538,N_1880);
xor U4536 (N_4536,N_718,N_2034);
or U4537 (N_4537,N_553,N_335);
nor U4538 (N_4538,N_1359,N_2637);
nor U4539 (N_4539,N_1075,N_2383);
or U4540 (N_4540,N_124,N_161);
nor U4541 (N_4541,N_565,N_125);
nor U4542 (N_4542,N_1794,N_60);
and U4543 (N_4543,N_1196,N_1503);
xnor U4544 (N_4544,N_1186,N_2719);
and U4545 (N_4545,N_1144,N_2895);
xor U4546 (N_4546,N_2125,N_1638);
nand U4547 (N_4547,N_2353,N_239);
nand U4548 (N_4548,N_2076,N_1309);
or U4549 (N_4549,N_1278,N_1950);
nand U4550 (N_4550,N_1397,N_377);
or U4551 (N_4551,N_756,N_2527);
nor U4552 (N_4552,N_2903,N_1581);
xor U4553 (N_4553,N_2712,N_2897);
nand U4554 (N_4554,N_295,N_32);
nor U4555 (N_4555,N_1626,N_439);
nor U4556 (N_4556,N_2436,N_564);
or U4557 (N_4557,N_2969,N_2826);
or U4558 (N_4558,N_1920,N_2970);
nand U4559 (N_4559,N_680,N_1595);
nand U4560 (N_4560,N_53,N_909);
nand U4561 (N_4561,N_2163,N_899);
and U4562 (N_4562,N_2677,N_2351);
or U4563 (N_4563,N_2801,N_717);
or U4564 (N_4564,N_2348,N_1825);
nor U4565 (N_4565,N_225,N_1218);
nor U4566 (N_4566,N_2901,N_2956);
or U4567 (N_4567,N_2098,N_2528);
nand U4568 (N_4568,N_2295,N_2009);
xnor U4569 (N_4569,N_2585,N_799);
and U4570 (N_4570,N_613,N_173);
nand U4571 (N_4571,N_2402,N_1206);
or U4572 (N_4572,N_1600,N_2328);
nor U4573 (N_4573,N_1742,N_1099);
and U4574 (N_4574,N_1778,N_2007);
and U4575 (N_4575,N_983,N_404);
or U4576 (N_4576,N_255,N_2222);
and U4577 (N_4577,N_948,N_686);
and U4578 (N_4578,N_1340,N_2008);
xnor U4579 (N_4579,N_859,N_2824);
nand U4580 (N_4580,N_1110,N_2649);
nand U4581 (N_4581,N_1312,N_2797);
and U4582 (N_4582,N_1664,N_15);
and U4583 (N_4583,N_2867,N_2000);
nand U4584 (N_4584,N_244,N_1341);
nand U4585 (N_4585,N_162,N_2555);
or U4586 (N_4586,N_2386,N_1189);
xor U4587 (N_4587,N_429,N_2425);
xor U4588 (N_4588,N_2112,N_1119);
or U4589 (N_4589,N_1768,N_434);
or U4590 (N_4590,N_812,N_1812);
nor U4591 (N_4591,N_1072,N_2985);
or U4592 (N_4592,N_139,N_1055);
nand U4593 (N_4593,N_2971,N_2940);
nor U4594 (N_4594,N_614,N_2753);
and U4595 (N_4595,N_1842,N_252);
or U4596 (N_4596,N_981,N_1796);
and U4597 (N_4597,N_526,N_1674);
xnor U4598 (N_4598,N_739,N_59);
nor U4599 (N_4599,N_1710,N_1913);
or U4600 (N_4600,N_1457,N_2499);
and U4601 (N_4601,N_1028,N_2609);
and U4602 (N_4602,N_1975,N_2718);
or U4603 (N_4603,N_105,N_2645);
and U4604 (N_4604,N_1775,N_454);
or U4605 (N_4605,N_126,N_179);
xor U4606 (N_4606,N_268,N_430);
or U4607 (N_4607,N_1402,N_1369);
xnor U4608 (N_4608,N_70,N_416);
nor U4609 (N_4609,N_45,N_1266);
or U4610 (N_4610,N_1056,N_2865);
xnor U4611 (N_4611,N_1243,N_299);
nor U4612 (N_4612,N_2512,N_2585);
nor U4613 (N_4613,N_2826,N_1075);
and U4614 (N_4614,N_1163,N_2097);
nor U4615 (N_4615,N_14,N_2155);
and U4616 (N_4616,N_2404,N_287);
nor U4617 (N_4617,N_243,N_2837);
xor U4618 (N_4618,N_1599,N_1886);
nand U4619 (N_4619,N_541,N_2718);
nand U4620 (N_4620,N_2443,N_2776);
nand U4621 (N_4621,N_1679,N_1553);
and U4622 (N_4622,N_2365,N_2271);
or U4623 (N_4623,N_937,N_517);
nor U4624 (N_4624,N_2101,N_1285);
nor U4625 (N_4625,N_1245,N_1677);
or U4626 (N_4626,N_2696,N_1232);
nor U4627 (N_4627,N_2576,N_131);
nand U4628 (N_4628,N_2536,N_1624);
or U4629 (N_4629,N_2698,N_2350);
or U4630 (N_4630,N_883,N_2717);
xor U4631 (N_4631,N_2698,N_2288);
or U4632 (N_4632,N_1496,N_2813);
nor U4633 (N_4633,N_740,N_399);
or U4634 (N_4634,N_1504,N_2706);
nand U4635 (N_4635,N_2441,N_1569);
nand U4636 (N_4636,N_2989,N_1096);
nor U4637 (N_4637,N_2251,N_1151);
xnor U4638 (N_4638,N_911,N_1221);
nand U4639 (N_4639,N_135,N_2781);
nand U4640 (N_4640,N_1262,N_2925);
nand U4641 (N_4641,N_1044,N_1854);
and U4642 (N_4642,N_1344,N_1654);
or U4643 (N_4643,N_498,N_27);
and U4644 (N_4644,N_571,N_1539);
and U4645 (N_4645,N_591,N_2561);
or U4646 (N_4646,N_1081,N_1390);
and U4647 (N_4647,N_2871,N_1205);
nor U4648 (N_4648,N_2618,N_1974);
and U4649 (N_4649,N_2913,N_2526);
xnor U4650 (N_4650,N_897,N_414);
or U4651 (N_4651,N_1353,N_1484);
and U4652 (N_4652,N_2858,N_1717);
xor U4653 (N_4653,N_1698,N_276);
nand U4654 (N_4654,N_116,N_491);
xnor U4655 (N_4655,N_379,N_49);
nor U4656 (N_4656,N_494,N_1615);
or U4657 (N_4657,N_795,N_2193);
and U4658 (N_4658,N_1900,N_157);
or U4659 (N_4659,N_1899,N_2569);
or U4660 (N_4660,N_1328,N_2096);
and U4661 (N_4661,N_1057,N_1602);
nor U4662 (N_4662,N_384,N_2684);
nor U4663 (N_4663,N_2888,N_2517);
or U4664 (N_4664,N_2658,N_1323);
and U4665 (N_4665,N_2657,N_413);
and U4666 (N_4666,N_152,N_2557);
or U4667 (N_4667,N_1257,N_1977);
and U4668 (N_4668,N_669,N_2069);
nand U4669 (N_4669,N_678,N_1671);
and U4670 (N_4670,N_2349,N_1387);
nor U4671 (N_4671,N_424,N_779);
or U4672 (N_4672,N_431,N_2131);
or U4673 (N_4673,N_369,N_287);
nor U4674 (N_4674,N_1398,N_2183);
nor U4675 (N_4675,N_1644,N_1836);
nand U4676 (N_4676,N_1552,N_1833);
nor U4677 (N_4677,N_1790,N_998);
and U4678 (N_4678,N_1663,N_2321);
nor U4679 (N_4679,N_2886,N_2791);
and U4680 (N_4680,N_323,N_1652);
nor U4681 (N_4681,N_2091,N_2770);
nand U4682 (N_4682,N_191,N_584);
nand U4683 (N_4683,N_652,N_2055);
and U4684 (N_4684,N_1658,N_2961);
nand U4685 (N_4685,N_2129,N_2871);
or U4686 (N_4686,N_878,N_1998);
nor U4687 (N_4687,N_797,N_1851);
nand U4688 (N_4688,N_2148,N_2489);
xor U4689 (N_4689,N_762,N_966);
nand U4690 (N_4690,N_973,N_2446);
and U4691 (N_4691,N_2459,N_506);
nor U4692 (N_4692,N_1644,N_501);
or U4693 (N_4693,N_737,N_349);
and U4694 (N_4694,N_338,N_792);
nand U4695 (N_4695,N_2325,N_819);
or U4696 (N_4696,N_2476,N_762);
nand U4697 (N_4697,N_1546,N_1788);
nand U4698 (N_4698,N_1068,N_2889);
and U4699 (N_4699,N_2753,N_339);
and U4700 (N_4700,N_472,N_474);
and U4701 (N_4701,N_938,N_666);
and U4702 (N_4702,N_2197,N_27);
nor U4703 (N_4703,N_1360,N_1498);
xor U4704 (N_4704,N_55,N_1241);
and U4705 (N_4705,N_1320,N_1714);
and U4706 (N_4706,N_35,N_977);
nand U4707 (N_4707,N_2048,N_2340);
nand U4708 (N_4708,N_1196,N_2179);
or U4709 (N_4709,N_1960,N_251);
nor U4710 (N_4710,N_2819,N_1092);
and U4711 (N_4711,N_1590,N_1201);
and U4712 (N_4712,N_769,N_649);
and U4713 (N_4713,N_2614,N_1199);
or U4714 (N_4714,N_1525,N_2672);
nand U4715 (N_4715,N_1064,N_1563);
and U4716 (N_4716,N_2494,N_1812);
nor U4717 (N_4717,N_2275,N_840);
and U4718 (N_4718,N_1390,N_38);
and U4719 (N_4719,N_56,N_1985);
nand U4720 (N_4720,N_2368,N_1527);
or U4721 (N_4721,N_2959,N_416);
nand U4722 (N_4722,N_323,N_2362);
or U4723 (N_4723,N_2182,N_1923);
xor U4724 (N_4724,N_2318,N_2016);
nor U4725 (N_4725,N_2266,N_991);
or U4726 (N_4726,N_2120,N_1120);
nor U4727 (N_4727,N_2747,N_279);
or U4728 (N_4728,N_2162,N_94);
xnor U4729 (N_4729,N_1019,N_325);
or U4730 (N_4730,N_2522,N_1512);
nand U4731 (N_4731,N_656,N_329);
nand U4732 (N_4732,N_316,N_979);
nor U4733 (N_4733,N_839,N_332);
nor U4734 (N_4734,N_1801,N_300);
nor U4735 (N_4735,N_758,N_2603);
and U4736 (N_4736,N_370,N_53);
or U4737 (N_4737,N_2370,N_2259);
nand U4738 (N_4738,N_1815,N_768);
nand U4739 (N_4739,N_1004,N_976);
nand U4740 (N_4740,N_2668,N_2407);
and U4741 (N_4741,N_1035,N_560);
nand U4742 (N_4742,N_2348,N_156);
nor U4743 (N_4743,N_2074,N_472);
nor U4744 (N_4744,N_2720,N_2050);
and U4745 (N_4745,N_190,N_788);
and U4746 (N_4746,N_2475,N_70);
and U4747 (N_4747,N_1074,N_1842);
and U4748 (N_4748,N_1176,N_2373);
nand U4749 (N_4749,N_1035,N_1618);
nor U4750 (N_4750,N_1253,N_234);
or U4751 (N_4751,N_1281,N_1707);
or U4752 (N_4752,N_1814,N_2869);
or U4753 (N_4753,N_2314,N_1693);
nand U4754 (N_4754,N_832,N_302);
nand U4755 (N_4755,N_2548,N_1983);
nand U4756 (N_4756,N_1673,N_1382);
nor U4757 (N_4757,N_1887,N_1472);
or U4758 (N_4758,N_2735,N_2824);
and U4759 (N_4759,N_733,N_2358);
or U4760 (N_4760,N_2740,N_568);
and U4761 (N_4761,N_2006,N_2737);
or U4762 (N_4762,N_822,N_2358);
nand U4763 (N_4763,N_1958,N_2911);
and U4764 (N_4764,N_1573,N_2910);
or U4765 (N_4765,N_2207,N_1099);
or U4766 (N_4766,N_484,N_2240);
nor U4767 (N_4767,N_1371,N_1477);
nor U4768 (N_4768,N_1342,N_286);
or U4769 (N_4769,N_703,N_58);
nand U4770 (N_4770,N_1749,N_219);
nand U4771 (N_4771,N_2472,N_253);
or U4772 (N_4772,N_812,N_1737);
nand U4773 (N_4773,N_237,N_2700);
or U4774 (N_4774,N_2052,N_806);
nor U4775 (N_4775,N_1966,N_308);
nand U4776 (N_4776,N_541,N_1093);
or U4777 (N_4777,N_2253,N_2922);
and U4778 (N_4778,N_252,N_1800);
xor U4779 (N_4779,N_463,N_2095);
and U4780 (N_4780,N_1566,N_2656);
xnor U4781 (N_4781,N_2009,N_867);
or U4782 (N_4782,N_1085,N_2885);
nor U4783 (N_4783,N_1385,N_134);
nor U4784 (N_4784,N_2813,N_1756);
or U4785 (N_4785,N_2918,N_1324);
or U4786 (N_4786,N_2261,N_528);
or U4787 (N_4787,N_1363,N_2669);
and U4788 (N_4788,N_2887,N_2586);
nor U4789 (N_4789,N_1961,N_1394);
nand U4790 (N_4790,N_2043,N_499);
nor U4791 (N_4791,N_439,N_1665);
and U4792 (N_4792,N_2486,N_199);
nor U4793 (N_4793,N_905,N_2932);
or U4794 (N_4794,N_171,N_1711);
xor U4795 (N_4795,N_2217,N_1535);
and U4796 (N_4796,N_591,N_1174);
nor U4797 (N_4797,N_902,N_366);
nor U4798 (N_4798,N_1590,N_2492);
and U4799 (N_4799,N_1208,N_2517);
nor U4800 (N_4800,N_555,N_1327);
and U4801 (N_4801,N_2926,N_1244);
and U4802 (N_4802,N_2158,N_2868);
nor U4803 (N_4803,N_941,N_933);
or U4804 (N_4804,N_802,N_2109);
and U4805 (N_4805,N_1013,N_2633);
and U4806 (N_4806,N_2147,N_890);
nor U4807 (N_4807,N_177,N_1984);
and U4808 (N_4808,N_992,N_176);
or U4809 (N_4809,N_902,N_29);
or U4810 (N_4810,N_189,N_401);
and U4811 (N_4811,N_233,N_1335);
and U4812 (N_4812,N_427,N_577);
nor U4813 (N_4813,N_1579,N_866);
or U4814 (N_4814,N_1094,N_2073);
and U4815 (N_4815,N_1896,N_1781);
xor U4816 (N_4816,N_2653,N_979);
nand U4817 (N_4817,N_857,N_2425);
and U4818 (N_4818,N_2272,N_934);
xor U4819 (N_4819,N_661,N_1579);
or U4820 (N_4820,N_2061,N_1908);
or U4821 (N_4821,N_527,N_2616);
and U4822 (N_4822,N_1350,N_586);
nor U4823 (N_4823,N_2497,N_870);
nor U4824 (N_4824,N_1159,N_221);
xor U4825 (N_4825,N_2855,N_392);
xnor U4826 (N_4826,N_362,N_2374);
or U4827 (N_4827,N_1439,N_2818);
or U4828 (N_4828,N_2789,N_1791);
or U4829 (N_4829,N_27,N_765);
nand U4830 (N_4830,N_2480,N_2514);
or U4831 (N_4831,N_1277,N_452);
or U4832 (N_4832,N_2349,N_2516);
or U4833 (N_4833,N_1866,N_779);
nand U4834 (N_4834,N_655,N_2707);
xnor U4835 (N_4835,N_1447,N_707);
and U4836 (N_4836,N_2343,N_2004);
or U4837 (N_4837,N_2925,N_1823);
xnor U4838 (N_4838,N_2017,N_523);
or U4839 (N_4839,N_576,N_567);
and U4840 (N_4840,N_2498,N_2468);
nand U4841 (N_4841,N_623,N_2829);
or U4842 (N_4842,N_2951,N_542);
or U4843 (N_4843,N_19,N_148);
nand U4844 (N_4844,N_1214,N_202);
nor U4845 (N_4845,N_1867,N_2067);
or U4846 (N_4846,N_720,N_2801);
and U4847 (N_4847,N_1145,N_1603);
nand U4848 (N_4848,N_2699,N_976);
nand U4849 (N_4849,N_715,N_2796);
nand U4850 (N_4850,N_1267,N_1653);
and U4851 (N_4851,N_1690,N_2073);
or U4852 (N_4852,N_2961,N_334);
or U4853 (N_4853,N_657,N_773);
nand U4854 (N_4854,N_2901,N_786);
nor U4855 (N_4855,N_801,N_2033);
nand U4856 (N_4856,N_2082,N_2489);
nand U4857 (N_4857,N_36,N_1471);
nor U4858 (N_4858,N_1170,N_2521);
nor U4859 (N_4859,N_1243,N_2572);
or U4860 (N_4860,N_830,N_802);
and U4861 (N_4861,N_1684,N_2771);
nor U4862 (N_4862,N_2389,N_73);
nand U4863 (N_4863,N_509,N_2043);
and U4864 (N_4864,N_2905,N_200);
xor U4865 (N_4865,N_2919,N_1627);
and U4866 (N_4866,N_1363,N_327);
and U4867 (N_4867,N_981,N_2775);
nor U4868 (N_4868,N_304,N_2802);
xor U4869 (N_4869,N_1754,N_2344);
nand U4870 (N_4870,N_420,N_1099);
or U4871 (N_4871,N_1869,N_3);
nor U4872 (N_4872,N_1883,N_1506);
nand U4873 (N_4873,N_2809,N_1608);
nand U4874 (N_4874,N_2595,N_2022);
xnor U4875 (N_4875,N_446,N_358);
nor U4876 (N_4876,N_1513,N_2104);
and U4877 (N_4877,N_2559,N_535);
nor U4878 (N_4878,N_2924,N_1158);
or U4879 (N_4879,N_771,N_2131);
or U4880 (N_4880,N_800,N_2350);
nor U4881 (N_4881,N_524,N_2969);
and U4882 (N_4882,N_2183,N_1065);
nor U4883 (N_4883,N_2594,N_2092);
or U4884 (N_4884,N_2045,N_1222);
nand U4885 (N_4885,N_1593,N_1355);
nand U4886 (N_4886,N_1587,N_2608);
xnor U4887 (N_4887,N_2134,N_2322);
nand U4888 (N_4888,N_420,N_639);
nor U4889 (N_4889,N_1801,N_1487);
and U4890 (N_4890,N_289,N_1371);
or U4891 (N_4891,N_1089,N_2571);
nor U4892 (N_4892,N_80,N_1625);
xor U4893 (N_4893,N_2708,N_2370);
nand U4894 (N_4894,N_2727,N_1398);
or U4895 (N_4895,N_274,N_2842);
or U4896 (N_4896,N_1357,N_2129);
and U4897 (N_4897,N_713,N_2470);
nor U4898 (N_4898,N_918,N_132);
or U4899 (N_4899,N_1344,N_1220);
or U4900 (N_4900,N_599,N_842);
nor U4901 (N_4901,N_810,N_1173);
xor U4902 (N_4902,N_2260,N_2797);
or U4903 (N_4903,N_435,N_22);
or U4904 (N_4904,N_1979,N_724);
or U4905 (N_4905,N_603,N_316);
nand U4906 (N_4906,N_1598,N_219);
nor U4907 (N_4907,N_1606,N_1696);
nor U4908 (N_4908,N_2868,N_1263);
nor U4909 (N_4909,N_753,N_289);
nor U4910 (N_4910,N_1662,N_1026);
nor U4911 (N_4911,N_2899,N_1324);
nor U4912 (N_4912,N_262,N_2623);
nand U4913 (N_4913,N_296,N_729);
nand U4914 (N_4914,N_2755,N_590);
nor U4915 (N_4915,N_936,N_1563);
or U4916 (N_4916,N_326,N_2543);
or U4917 (N_4917,N_2568,N_939);
nand U4918 (N_4918,N_712,N_2298);
nor U4919 (N_4919,N_2271,N_718);
nor U4920 (N_4920,N_2976,N_2285);
nand U4921 (N_4921,N_2341,N_2538);
nor U4922 (N_4922,N_1748,N_2080);
and U4923 (N_4923,N_733,N_1242);
or U4924 (N_4924,N_2981,N_2048);
or U4925 (N_4925,N_2809,N_776);
and U4926 (N_4926,N_2303,N_1885);
nand U4927 (N_4927,N_2656,N_1180);
nor U4928 (N_4928,N_873,N_748);
nand U4929 (N_4929,N_622,N_1736);
nor U4930 (N_4930,N_2700,N_428);
xnor U4931 (N_4931,N_1647,N_2188);
or U4932 (N_4932,N_211,N_1565);
xnor U4933 (N_4933,N_431,N_907);
and U4934 (N_4934,N_1008,N_1838);
or U4935 (N_4935,N_1202,N_1089);
nand U4936 (N_4936,N_29,N_117);
nor U4937 (N_4937,N_2975,N_202);
or U4938 (N_4938,N_2025,N_1117);
and U4939 (N_4939,N_2631,N_2952);
nand U4940 (N_4940,N_2476,N_2960);
nand U4941 (N_4941,N_1710,N_2848);
or U4942 (N_4942,N_780,N_1966);
nand U4943 (N_4943,N_1690,N_1162);
or U4944 (N_4944,N_1983,N_2617);
or U4945 (N_4945,N_736,N_1518);
nand U4946 (N_4946,N_1390,N_1026);
nand U4947 (N_4947,N_28,N_1841);
nor U4948 (N_4948,N_1276,N_449);
and U4949 (N_4949,N_491,N_2562);
or U4950 (N_4950,N_753,N_1351);
nor U4951 (N_4951,N_2582,N_2868);
nor U4952 (N_4952,N_983,N_2341);
nor U4953 (N_4953,N_498,N_2003);
nor U4954 (N_4954,N_191,N_1442);
nor U4955 (N_4955,N_2065,N_2016);
or U4956 (N_4956,N_1508,N_2339);
or U4957 (N_4957,N_1213,N_1153);
or U4958 (N_4958,N_2377,N_2757);
and U4959 (N_4959,N_2228,N_2028);
nand U4960 (N_4960,N_2895,N_2410);
nor U4961 (N_4961,N_1325,N_948);
and U4962 (N_4962,N_37,N_322);
nand U4963 (N_4963,N_298,N_774);
nor U4964 (N_4964,N_927,N_72);
or U4965 (N_4965,N_1119,N_734);
nor U4966 (N_4966,N_2686,N_578);
and U4967 (N_4967,N_2698,N_399);
or U4968 (N_4968,N_1537,N_252);
and U4969 (N_4969,N_1541,N_2345);
or U4970 (N_4970,N_2626,N_2304);
nor U4971 (N_4971,N_2610,N_1215);
or U4972 (N_4972,N_396,N_2148);
nor U4973 (N_4973,N_98,N_836);
nand U4974 (N_4974,N_2999,N_455);
and U4975 (N_4975,N_742,N_2134);
or U4976 (N_4976,N_1666,N_1968);
or U4977 (N_4977,N_1155,N_179);
or U4978 (N_4978,N_741,N_1289);
nand U4979 (N_4979,N_758,N_402);
nand U4980 (N_4980,N_807,N_492);
nand U4981 (N_4981,N_679,N_1919);
nand U4982 (N_4982,N_391,N_1011);
nor U4983 (N_4983,N_769,N_2471);
and U4984 (N_4984,N_2484,N_193);
xnor U4985 (N_4985,N_367,N_1401);
nor U4986 (N_4986,N_1779,N_2580);
or U4987 (N_4987,N_1306,N_18);
nor U4988 (N_4988,N_1231,N_2343);
or U4989 (N_4989,N_934,N_1651);
or U4990 (N_4990,N_899,N_2990);
nor U4991 (N_4991,N_1615,N_2303);
nand U4992 (N_4992,N_260,N_1820);
xnor U4993 (N_4993,N_1220,N_2271);
nand U4994 (N_4994,N_2461,N_675);
and U4995 (N_4995,N_824,N_985);
xor U4996 (N_4996,N_2644,N_214);
or U4997 (N_4997,N_2553,N_982);
or U4998 (N_4998,N_1339,N_2361);
and U4999 (N_4999,N_1982,N_1071);
or U5000 (N_5000,N_1572,N_1267);
nor U5001 (N_5001,N_2634,N_1218);
nand U5002 (N_5002,N_353,N_973);
and U5003 (N_5003,N_1128,N_797);
nand U5004 (N_5004,N_2407,N_2286);
nand U5005 (N_5005,N_2597,N_1064);
and U5006 (N_5006,N_335,N_2376);
xor U5007 (N_5007,N_728,N_2687);
nor U5008 (N_5008,N_2149,N_2628);
and U5009 (N_5009,N_2096,N_1463);
nand U5010 (N_5010,N_1150,N_2182);
and U5011 (N_5011,N_622,N_879);
or U5012 (N_5012,N_2454,N_1833);
and U5013 (N_5013,N_1382,N_1868);
nor U5014 (N_5014,N_2325,N_2645);
or U5015 (N_5015,N_677,N_231);
nand U5016 (N_5016,N_1682,N_2941);
nor U5017 (N_5017,N_2694,N_2230);
xnor U5018 (N_5018,N_2925,N_266);
and U5019 (N_5019,N_2652,N_1492);
nand U5020 (N_5020,N_1375,N_2650);
nand U5021 (N_5021,N_2883,N_833);
and U5022 (N_5022,N_218,N_814);
nand U5023 (N_5023,N_2188,N_581);
xor U5024 (N_5024,N_2959,N_2059);
and U5025 (N_5025,N_1406,N_1925);
or U5026 (N_5026,N_2948,N_465);
or U5027 (N_5027,N_2028,N_1842);
and U5028 (N_5028,N_952,N_739);
xor U5029 (N_5029,N_1156,N_644);
or U5030 (N_5030,N_1075,N_2816);
nor U5031 (N_5031,N_141,N_1752);
nand U5032 (N_5032,N_587,N_775);
and U5033 (N_5033,N_1027,N_1012);
nand U5034 (N_5034,N_717,N_2371);
nand U5035 (N_5035,N_1144,N_683);
nor U5036 (N_5036,N_2760,N_2172);
nand U5037 (N_5037,N_1610,N_2918);
or U5038 (N_5038,N_172,N_1712);
and U5039 (N_5039,N_1079,N_2463);
or U5040 (N_5040,N_1160,N_1082);
xor U5041 (N_5041,N_1257,N_1762);
or U5042 (N_5042,N_160,N_2219);
or U5043 (N_5043,N_2126,N_369);
nand U5044 (N_5044,N_2378,N_1971);
nand U5045 (N_5045,N_355,N_2693);
nor U5046 (N_5046,N_2286,N_2624);
nor U5047 (N_5047,N_291,N_2928);
or U5048 (N_5048,N_641,N_1563);
or U5049 (N_5049,N_1794,N_1480);
nand U5050 (N_5050,N_2963,N_1872);
xor U5051 (N_5051,N_206,N_1325);
and U5052 (N_5052,N_1345,N_439);
or U5053 (N_5053,N_2802,N_958);
and U5054 (N_5054,N_1284,N_1590);
and U5055 (N_5055,N_586,N_1325);
and U5056 (N_5056,N_2073,N_634);
nor U5057 (N_5057,N_2961,N_2719);
nand U5058 (N_5058,N_1080,N_2862);
xor U5059 (N_5059,N_2863,N_2075);
xor U5060 (N_5060,N_116,N_963);
nor U5061 (N_5061,N_2205,N_174);
nor U5062 (N_5062,N_46,N_1939);
nor U5063 (N_5063,N_1611,N_2976);
and U5064 (N_5064,N_1377,N_1670);
and U5065 (N_5065,N_2449,N_1980);
or U5066 (N_5066,N_1394,N_1517);
nor U5067 (N_5067,N_2906,N_1697);
nand U5068 (N_5068,N_1005,N_1324);
nand U5069 (N_5069,N_1699,N_969);
nor U5070 (N_5070,N_1394,N_777);
and U5071 (N_5071,N_808,N_734);
nand U5072 (N_5072,N_1620,N_301);
nand U5073 (N_5073,N_1515,N_2124);
and U5074 (N_5074,N_1285,N_1422);
and U5075 (N_5075,N_1995,N_2830);
nor U5076 (N_5076,N_1654,N_2492);
or U5077 (N_5077,N_739,N_2541);
and U5078 (N_5078,N_2984,N_2192);
xnor U5079 (N_5079,N_2173,N_2820);
nor U5080 (N_5080,N_70,N_1834);
nand U5081 (N_5081,N_1923,N_2452);
nand U5082 (N_5082,N_494,N_1415);
or U5083 (N_5083,N_1567,N_694);
nand U5084 (N_5084,N_48,N_549);
or U5085 (N_5085,N_1063,N_1629);
nor U5086 (N_5086,N_1393,N_1953);
or U5087 (N_5087,N_384,N_544);
nor U5088 (N_5088,N_1032,N_2431);
xor U5089 (N_5089,N_2086,N_1451);
nand U5090 (N_5090,N_397,N_2000);
nand U5091 (N_5091,N_42,N_2508);
or U5092 (N_5092,N_833,N_1928);
or U5093 (N_5093,N_1147,N_2424);
nand U5094 (N_5094,N_1504,N_2084);
or U5095 (N_5095,N_790,N_2327);
or U5096 (N_5096,N_2657,N_1782);
or U5097 (N_5097,N_2372,N_2201);
xor U5098 (N_5098,N_2118,N_2975);
nor U5099 (N_5099,N_1817,N_952);
nand U5100 (N_5100,N_330,N_2037);
nor U5101 (N_5101,N_738,N_671);
and U5102 (N_5102,N_2650,N_2733);
nand U5103 (N_5103,N_204,N_1537);
and U5104 (N_5104,N_573,N_2793);
or U5105 (N_5105,N_1299,N_564);
and U5106 (N_5106,N_82,N_1495);
nand U5107 (N_5107,N_776,N_1945);
and U5108 (N_5108,N_2366,N_41);
xnor U5109 (N_5109,N_605,N_2987);
and U5110 (N_5110,N_832,N_2868);
nor U5111 (N_5111,N_1030,N_107);
and U5112 (N_5112,N_987,N_541);
nor U5113 (N_5113,N_1547,N_1302);
nor U5114 (N_5114,N_1665,N_1143);
or U5115 (N_5115,N_2039,N_2151);
or U5116 (N_5116,N_2721,N_2820);
nor U5117 (N_5117,N_361,N_146);
nor U5118 (N_5118,N_257,N_446);
nand U5119 (N_5119,N_2276,N_1657);
nand U5120 (N_5120,N_924,N_2578);
nand U5121 (N_5121,N_1658,N_2834);
nor U5122 (N_5122,N_2153,N_2339);
nand U5123 (N_5123,N_2538,N_1266);
or U5124 (N_5124,N_508,N_1060);
or U5125 (N_5125,N_665,N_2227);
nand U5126 (N_5126,N_879,N_2039);
or U5127 (N_5127,N_1158,N_2443);
or U5128 (N_5128,N_2359,N_62);
nor U5129 (N_5129,N_1260,N_1290);
nand U5130 (N_5130,N_786,N_2741);
or U5131 (N_5131,N_1349,N_2562);
nor U5132 (N_5132,N_2366,N_828);
and U5133 (N_5133,N_2757,N_1127);
xnor U5134 (N_5134,N_794,N_1870);
xor U5135 (N_5135,N_1336,N_1603);
and U5136 (N_5136,N_1722,N_212);
or U5137 (N_5137,N_1436,N_283);
and U5138 (N_5138,N_2907,N_655);
nand U5139 (N_5139,N_1641,N_825);
nor U5140 (N_5140,N_2079,N_1363);
and U5141 (N_5141,N_1608,N_1471);
and U5142 (N_5142,N_2566,N_1777);
and U5143 (N_5143,N_292,N_1988);
nor U5144 (N_5144,N_2682,N_773);
or U5145 (N_5145,N_701,N_2658);
or U5146 (N_5146,N_884,N_772);
and U5147 (N_5147,N_2501,N_2006);
and U5148 (N_5148,N_1457,N_2617);
or U5149 (N_5149,N_821,N_2550);
xor U5150 (N_5150,N_2971,N_2430);
or U5151 (N_5151,N_2860,N_2065);
and U5152 (N_5152,N_2874,N_1518);
or U5153 (N_5153,N_375,N_30);
or U5154 (N_5154,N_1477,N_2185);
and U5155 (N_5155,N_608,N_1649);
nand U5156 (N_5156,N_608,N_588);
nor U5157 (N_5157,N_83,N_97);
and U5158 (N_5158,N_1637,N_1277);
xnor U5159 (N_5159,N_814,N_2143);
nor U5160 (N_5160,N_182,N_27);
and U5161 (N_5161,N_2003,N_552);
or U5162 (N_5162,N_1833,N_1416);
or U5163 (N_5163,N_131,N_2271);
nor U5164 (N_5164,N_171,N_2179);
or U5165 (N_5165,N_305,N_1301);
nor U5166 (N_5166,N_2309,N_2643);
and U5167 (N_5167,N_1148,N_2424);
nor U5168 (N_5168,N_1340,N_1816);
or U5169 (N_5169,N_1957,N_467);
and U5170 (N_5170,N_478,N_1545);
and U5171 (N_5171,N_2635,N_1295);
xnor U5172 (N_5172,N_183,N_2656);
nand U5173 (N_5173,N_1615,N_1359);
nand U5174 (N_5174,N_2451,N_1320);
or U5175 (N_5175,N_1098,N_2576);
xor U5176 (N_5176,N_1748,N_2882);
xor U5177 (N_5177,N_987,N_2061);
nor U5178 (N_5178,N_1367,N_1958);
xor U5179 (N_5179,N_724,N_2040);
or U5180 (N_5180,N_1389,N_2478);
or U5181 (N_5181,N_2623,N_1368);
or U5182 (N_5182,N_1673,N_445);
nor U5183 (N_5183,N_1039,N_197);
nor U5184 (N_5184,N_2398,N_872);
xnor U5185 (N_5185,N_1140,N_1321);
or U5186 (N_5186,N_786,N_1164);
or U5187 (N_5187,N_1322,N_2177);
nand U5188 (N_5188,N_595,N_2485);
or U5189 (N_5189,N_597,N_2697);
and U5190 (N_5190,N_911,N_1234);
nor U5191 (N_5191,N_1371,N_56);
and U5192 (N_5192,N_2812,N_2230);
nand U5193 (N_5193,N_2261,N_1482);
nor U5194 (N_5194,N_2105,N_1028);
nand U5195 (N_5195,N_181,N_1159);
nor U5196 (N_5196,N_2598,N_2582);
xor U5197 (N_5197,N_1014,N_1383);
nand U5198 (N_5198,N_392,N_2255);
and U5199 (N_5199,N_158,N_399);
and U5200 (N_5200,N_2568,N_2722);
and U5201 (N_5201,N_1061,N_1702);
xor U5202 (N_5202,N_1175,N_1806);
nand U5203 (N_5203,N_1135,N_1281);
and U5204 (N_5204,N_110,N_741);
and U5205 (N_5205,N_2319,N_2442);
and U5206 (N_5206,N_1679,N_1285);
or U5207 (N_5207,N_759,N_1854);
and U5208 (N_5208,N_624,N_1188);
nor U5209 (N_5209,N_776,N_1254);
and U5210 (N_5210,N_1494,N_2526);
nand U5211 (N_5211,N_2493,N_709);
nor U5212 (N_5212,N_2000,N_76);
or U5213 (N_5213,N_718,N_1371);
or U5214 (N_5214,N_2282,N_1315);
or U5215 (N_5215,N_2429,N_897);
and U5216 (N_5216,N_1207,N_224);
or U5217 (N_5217,N_1227,N_1327);
nand U5218 (N_5218,N_974,N_1844);
nor U5219 (N_5219,N_911,N_1544);
or U5220 (N_5220,N_2934,N_1205);
and U5221 (N_5221,N_1049,N_752);
or U5222 (N_5222,N_2406,N_2526);
xor U5223 (N_5223,N_1348,N_172);
nand U5224 (N_5224,N_2183,N_2955);
nand U5225 (N_5225,N_502,N_802);
nand U5226 (N_5226,N_498,N_814);
xor U5227 (N_5227,N_148,N_1029);
nand U5228 (N_5228,N_581,N_1777);
and U5229 (N_5229,N_2838,N_1211);
or U5230 (N_5230,N_1740,N_496);
and U5231 (N_5231,N_2355,N_1856);
nor U5232 (N_5232,N_1326,N_2182);
and U5233 (N_5233,N_1269,N_2603);
xor U5234 (N_5234,N_689,N_2184);
and U5235 (N_5235,N_1237,N_882);
nand U5236 (N_5236,N_345,N_121);
nand U5237 (N_5237,N_2985,N_2802);
nand U5238 (N_5238,N_452,N_280);
nand U5239 (N_5239,N_493,N_2599);
nor U5240 (N_5240,N_522,N_1745);
or U5241 (N_5241,N_2118,N_765);
and U5242 (N_5242,N_2703,N_580);
or U5243 (N_5243,N_2257,N_1649);
and U5244 (N_5244,N_2069,N_2162);
and U5245 (N_5245,N_2910,N_2955);
and U5246 (N_5246,N_1325,N_916);
nand U5247 (N_5247,N_1030,N_806);
nand U5248 (N_5248,N_1585,N_835);
xnor U5249 (N_5249,N_2315,N_1321);
nor U5250 (N_5250,N_724,N_2614);
nand U5251 (N_5251,N_485,N_301);
xor U5252 (N_5252,N_1939,N_1968);
nor U5253 (N_5253,N_2135,N_2671);
nor U5254 (N_5254,N_285,N_923);
or U5255 (N_5255,N_1203,N_1931);
nand U5256 (N_5256,N_2058,N_2338);
or U5257 (N_5257,N_2627,N_301);
or U5258 (N_5258,N_2028,N_1407);
and U5259 (N_5259,N_2058,N_53);
nor U5260 (N_5260,N_2723,N_152);
nor U5261 (N_5261,N_2609,N_1542);
or U5262 (N_5262,N_249,N_661);
nor U5263 (N_5263,N_2584,N_2671);
xnor U5264 (N_5264,N_785,N_51);
nand U5265 (N_5265,N_293,N_192);
or U5266 (N_5266,N_484,N_2810);
or U5267 (N_5267,N_2294,N_1524);
nor U5268 (N_5268,N_1451,N_214);
nand U5269 (N_5269,N_1781,N_706);
nor U5270 (N_5270,N_1164,N_1862);
and U5271 (N_5271,N_721,N_2015);
and U5272 (N_5272,N_1909,N_252);
and U5273 (N_5273,N_1284,N_557);
nand U5274 (N_5274,N_2858,N_1387);
nor U5275 (N_5275,N_1382,N_2242);
or U5276 (N_5276,N_2235,N_2110);
nand U5277 (N_5277,N_501,N_1268);
or U5278 (N_5278,N_1882,N_60);
nand U5279 (N_5279,N_336,N_1463);
nor U5280 (N_5280,N_16,N_673);
nand U5281 (N_5281,N_2140,N_308);
nand U5282 (N_5282,N_184,N_2624);
nor U5283 (N_5283,N_2021,N_393);
or U5284 (N_5284,N_2985,N_597);
or U5285 (N_5285,N_2121,N_1934);
xor U5286 (N_5286,N_1535,N_726);
nor U5287 (N_5287,N_671,N_1437);
or U5288 (N_5288,N_973,N_2075);
or U5289 (N_5289,N_655,N_2621);
nand U5290 (N_5290,N_1296,N_2031);
and U5291 (N_5291,N_1542,N_52);
nand U5292 (N_5292,N_2328,N_412);
nor U5293 (N_5293,N_1707,N_2699);
nor U5294 (N_5294,N_1316,N_1679);
xor U5295 (N_5295,N_1083,N_491);
xor U5296 (N_5296,N_73,N_971);
nand U5297 (N_5297,N_2947,N_2516);
nor U5298 (N_5298,N_27,N_1726);
or U5299 (N_5299,N_2144,N_1427);
nor U5300 (N_5300,N_1885,N_2643);
and U5301 (N_5301,N_1896,N_2364);
nand U5302 (N_5302,N_1181,N_466);
or U5303 (N_5303,N_716,N_598);
and U5304 (N_5304,N_285,N_313);
nor U5305 (N_5305,N_1027,N_75);
nor U5306 (N_5306,N_158,N_594);
and U5307 (N_5307,N_1504,N_319);
xor U5308 (N_5308,N_2394,N_1544);
xnor U5309 (N_5309,N_787,N_1407);
xnor U5310 (N_5310,N_2740,N_2231);
and U5311 (N_5311,N_1498,N_1605);
or U5312 (N_5312,N_420,N_2149);
or U5313 (N_5313,N_501,N_2327);
or U5314 (N_5314,N_856,N_696);
or U5315 (N_5315,N_503,N_1758);
or U5316 (N_5316,N_1082,N_1570);
nand U5317 (N_5317,N_541,N_1005);
xor U5318 (N_5318,N_1019,N_457);
nor U5319 (N_5319,N_1830,N_1293);
nor U5320 (N_5320,N_555,N_2108);
or U5321 (N_5321,N_1204,N_1067);
nor U5322 (N_5322,N_564,N_544);
nor U5323 (N_5323,N_2553,N_1925);
xor U5324 (N_5324,N_1014,N_2123);
nor U5325 (N_5325,N_231,N_1007);
and U5326 (N_5326,N_863,N_522);
nor U5327 (N_5327,N_1413,N_428);
nor U5328 (N_5328,N_1019,N_1409);
or U5329 (N_5329,N_401,N_2755);
or U5330 (N_5330,N_627,N_383);
nand U5331 (N_5331,N_572,N_1243);
and U5332 (N_5332,N_955,N_573);
xor U5333 (N_5333,N_600,N_2332);
and U5334 (N_5334,N_2199,N_466);
and U5335 (N_5335,N_656,N_2718);
nand U5336 (N_5336,N_1202,N_256);
nor U5337 (N_5337,N_2457,N_1037);
or U5338 (N_5338,N_2936,N_2923);
xnor U5339 (N_5339,N_953,N_1970);
or U5340 (N_5340,N_2429,N_2567);
or U5341 (N_5341,N_2763,N_2589);
or U5342 (N_5342,N_2660,N_2926);
nor U5343 (N_5343,N_634,N_742);
nand U5344 (N_5344,N_1475,N_1032);
and U5345 (N_5345,N_2474,N_362);
or U5346 (N_5346,N_1328,N_376);
and U5347 (N_5347,N_1957,N_2938);
and U5348 (N_5348,N_712,N_1436);
nor U5349 (N_5349,N_216,N_326);
and U5350 (N_5350,N_1822,N_2285);
nor U5351 (N_5351,N_314,N_207);
nor U5352 (N_5352,N_2424,N_1174);
or U5353 (N_5353,N_278,N_2519);
nor U5354 (N_5354,N_2597,N_174);
nand U5355 (N_5355,N_2645,N_832);
nor U5356 (N_5356,N_1754,N_2421);
nor U5357 (N_5357,N_84,N_2870);
nand U5358 (N_5358,N_1530,N_2326);
or U5359 (N_5359,N_1413,N_479);
nor U5360 (N_5360,N_366,N_2531);
nor U5361 (N_5361,N_2364,N_1263);
or U5362 (N_5362,N_2660,N_1727);
nor U5363 (N_5363,N_1719,N_1657);
nand U5364 (N_5364,N_2148,N_1629);
and U5365 (N_5365,N_1210,N_2256);
xnor U5366 (N_5366,N_1936,N_1551);
xnor U5367 (N_5367,N_2628,N_176);
nand U5368 (N_5368,N_1927,N_1200);
nand U5369 (N_5369,N_2922,N_2898);
nand U5370 (N_5370,N_2914,N_773);
xor U5371 (N_5371,N_2622,N_522);
nor U5372 (N_5372,N_1816,N_1333);
and U5373 (N_5373,N_773,N_2167);
nor U5374 (N_5374,N_1680,N_2935);
and U5375 (N_5375,N_56,N_2981);
nand U5376 (N_5376,N_330,N_1210);
and U5377 (N_5377,N_791,N_1859);
and U5378 (N_5378,N_2357,N_377);
and U5379 (N_5379,N_956,N_1792);
nand U5380 (N_5380,N_1651,N_472);
or U5381 (N_5381,N_2755,N_832);
nand U5382 (N_5382,N_998,N_1238);
and U5383 (N_5383,N_373,N_2617);
or U5384 (N_5384,N_225,N_1640);
xnor U5385 (N_5385,N_845,N_1615);
nor U5386 (N_5386,N_1130,N_2308);
nor U5387 (N_5387,N_1285,N_2930);
and U5388 (N_5388,N_2392,N_778);
nor U5389 (N_5389,N_1693,N_2746);
nand U5390 (N_5390,N_2028,N_33);
or U5391 (N_5391,N_927,N_1923);
and U5392 (N_5392,N_2264,N_1618);
and U5393 (N_5393,N_2257,N_1899);
nand U5394 (N_5394,N_467,N_1572);
nand U5395 (N_5395,N_474,N_1272);
nand U5396 (N_5396,N_2462,N_2324);
nand U5397 (N_5397,N_1857,N_2115);
or U5398 (N_5398,N_812,N_2724);
nor U5399 (N_5399,N_454,N_2871);
and U5400 (N_5400,N_2663,N_1784);
or U5401 (N_5401,N_2055,N_1410);
nor U5402 (N_5402,N_1256,N_1849);
nor U5403 (N_5403,N_2191,N_193);
nand U5404 (N_5404,N_729,N_2396);
nor U5405 (N_5405,N_1906,N_2691);
xor U5406 (N_5406,N_701,N_2752);
or U5407 (N_5407,N_2133,N_2300);
and U5408 (N_5408,N_2216,N_2647);
and U5409 (N_5409,N_1233,N_1190);
or U5410 (N_5410,N_299,N_549);
and U5411 (N_5411,N_2069,N_1568);
nor U5412 (N_5412,N_2022,N_2814);
nand U5413 (N_5413,N_1999,N_1945);
nand U5414 (N_5414,N_2545,N_1477);
nor U5415 (N_5415,N_734,N_804);
xnor U5416 (N_5416,N_839,N_981);
nand U5417 (N_5417,N_930,N_1188);
nor U5418 (N_5418,N_1588,N_1052);
or U5419 (N_5419,N_818,N_2552);
and U5420 (N_5420,N_847,N_1568);
and U5421 (N_5421,N_2102,N_2917);
nand U5422 (N_5422,N_1738,N_2367);
nand U5423 (N_5423,N_2408,N_2561);
nand U5424 (N_5424,N_135,N_2146);
nor U5425 (N_5425,N_887,N_2449);
nand U5426 (N_5426,N_1062,N_1450);
and U5427 (N_5427,N_2628,N_48);
or U5428 (N_5428,N_1704,N_1935);
nor U5429 (N_5429,N_874,N_2902);
or U5430 (N_5430,N_497,N_1673);
or U5431 (N_5431,N_1287,N_2797);
xor U5432 (N_5432,N_2964,N_807);
or U5433 (N_5433,N_1661,N_2127);
and U5434 (N_5434,N_1837,N_2868);
nor U5435 (N_5435,N_2958,N_857);
xor U5436 (N_5436,N_964,N_916);
nand U5437 (N_5437,N_573,N_338);
or U5438 (N_5438,N_376,N_1769);
xor U5439 (N_5439,N_2960,N_1496);
nor U5440 (N_5440,N_2954,N_2802);
or U5441 (N_5441,N_1101,N_2144);
nand U5442 (N_5442,N_1081,N_2687);
nor U5443 (N_5443,N_1107,N_2170);
nor U5444 (N_5444,N_1436,N_2125);
or U5445 (N_5445,N_1367,N_2629);
nand U5446 (N_5446,N_2076,N_1851);
xnor U5447 (N_5447,N_726,N_1762);
nand U5448 (N_5448,N_1055,N_41);
or U5449 (N_5449,N_2025,N_2804);
nor U5450 (N_5450,N_2691,N_1720);
nand U5451 (N_5451,N_1868,N_2727);
and U5452 (N_5452,N_342,N_2549);
nor U5453 (N_5453,N_2884,N_992);
nand U5454 (N_5454,N_2817,N_208);
or U5455 (N_5455,N_987,N_2880);
and U5456 (N_5456,N_833,N_1542);
or U5457 (N_5457,N_2731,N_1422);
nand U5458 (N_5458,N_2026,N_2894);
nand U5459 (N_5459,N_791,N_1343);
or U5460 (N_5460,N_83,N_2675);
and U5461 (N_5461,N_241,N_2974);
or U5462 (N_5462,N_2035,N_2679);
nand U5463 (N_5463,N_1665,N_1328);
and U5464 (N_5464,N_1970,N_1814);
nand U5465 (N_5465,N_1901,N_584);
nor U5466 (N_5466,N_1073,N_2201);
and U5467 (N_5467,N_2586,N_2073);
nand U5468 (N_5468,N_775,N_2968);
or U5469 (N_5469,N_1587,N_145);
and U5470 (N_5470,N_457,N_1716);
nor U5471 (N_5471,N_414,N_1856);
nor U5472 (N_5472,N_1856,N_2580);
or U5473 (N_5473,N_1396,N_977);
nor U5474 (N_5474,N_1480,N_226);
nand U5475 (N_5475,N_2401,N_106);
xor U5476 (N_5476,N_334,N_602);
nor U5477 (N_5477,N_2359,N_292);
nand U5478 (N_5478,N_789,N_974);
nor U5479 (N_5479,N_183,N_221);
or U5480 (N_5480,N_778,N_1050);
nor U5481 (N_5481,N_290,N_1032);
and U5482 (N_5482,N_889,N_2660);
and U5483 (N_5483,N_726,N_2529);
nand U5484 (N_5484,N_51,N_272);
or U5485 (N_5485,N_920,N_214);
or U5486 (N_5486,N_2368,N_2135);
or U5487 (N_5487,N_1881,N_941);
xor U5488 (N_5488,N_363,N_304);
nor U5489 (N_5489,N_524,N_1659);
nor U5490 (N_5490,N_2700,N_2221);
nand U5491 (N_5491,N_1983,N_349);
nand U5492 (N_5492,N_2476,N_2457);
and U5493 (N_5493,N_609,N_260);
nand U5494 (N_5494,N_80,N_64);
xnor U5495 (N_5495,N_1411,N_2637);
and U5496 (N_5496,N_613,N_103);
and U5497 (N_5497,N_2106,N_959);
nor U5498 (N_5498,N_303,N_1963);
nor U5499 (N_5499,N_1392,N_2593);
or U5500 (N_5500,N_1601,N_2728);
nor U5501 (N_5501,N_2511,N_2701);
nor U5502 (N_5502,N_456,N_1493);
nor U5503 (N_5503,N_383,N_2374);
xnor U5504 (N_5504,N_1287,N_1746);
nor U5505 (N_5505,N_1864,N_1766);
and U5506 (N_5506,N_504,N_1882);
or U5507 (N_5507,N_620,N_2221);
and U5508 (N_5508,N_1018,N_1084);
nand U5509 (N_5509,N_1950,N_405);
nand U5510 (N_5510,N_2502,N_703);
nand U5511 (N_5511,N_2262,N_2495);
and U5512 (N_5512,N_1407,N_1230);
xor U5513 (N_5513,N_163,N_348);
and U5514 (N_5514,N_2566,N_601);
nand U5515 (N_5515,N_2815,N_1331);
xnor U5516 (N_5516,N_2150,N_946);
nand U5517 (N_5517,N_2872,N_8);
nor U5518 (N_5518,N_1874,N_1956);
nor U5519 (N_5519,N_2379,N_441);
or U5520 (N_5520,N_1734,N_2586);
nand U5521 (N_5521,N_2290,N_364);
nor U5522 (N_5522,N_2307,N_31);
or U5523 (N_5523,N_1429,N_1395);
nor U5524 (N_5524,N_944,N_816);
and U5525 (N_5525,N_1015,N_63);
nand U5526 (N_5526,N_1302,N_263);
nand U5527 (N_5527,N_2846,N_2539);
nand U5528 (N_5528,N_1178,N_1829);
nand U5529 (N_5529,N_195,N_1560);
or U5530 (N_5530,N_1633,N_2187);
xnor U5531 (N_5531,N_1266,N_1276);
nor U5532 (N_5532,N_199,N_1422);
and U5533 (N_5533,N_2288,N_2057);
or U5534 (N_5534,N_434,N_1450);
nand U5535 (N_5535,N_2836,N_2536);
nand U5536 (N_5536,N_22,N_2223);
xnor U5537 (N_5537,N_673,N_521);
or U5538 (N_5538,N_2103,N_247);
or U5539 (N_5539,N_996,N_742);
nand U5540 (N_5540,N_453,N_1007);
nor U5541 (N_5541,N_1578,N_146);
nor U5542 (N_5542,N_1498,N_2028);
nand U5543 (N_5543,N_2031,N_1198);
or U5544 (N_5544,N_2982,N_2820);
and U5545 (N_5545,N_6,N_17);
or U5546 (N_5546,N_2442,N_1287);
nor U5547 (N_5547,N_1510,N_1059);
or U5548 (N_5548,N_56,N_1952);
nand U5549 (N_5549,N_1027,N_2665);
and U5550 (N_5550,N_155,N_1026);
nor U5551 (N_5551,N_2287,N_1780);
xnor U5552 (N_5552,N_2007,N_1826);
nand U5553 (N_5553,N_1587,N_2530);
nand U5554 (N_5554,N_2426,N_807);
xnor U5555 (N_5555,N_621,N_1302);
and U5556 (N_5556,N_1553,N_1294);
nor U5557 (N_5557,N_1152,N_1299);
nor U5558 (N_5558,N_1188,N_1640);
nor U5559 (N_5559,N_1105,N_2280);
or U5560 (N_5560,N_2276,N_2132);
nand U5561 (N_5561,N_793,N_1438);
nor U5562 (N_5562,N_798,N_1450);
or U5563 (N_5563,N_1676,N_650);
or U5564 (N_5564,N_2753,N_887);
and U5565 (N_5565,N_1492,N_2261);
nor U5566 (N_5566,N_2139,N_430);
and U5567 (N_5567,N_1952,N_2594);
xnor U5568 (N_5568,N_1087,N_2364);
or U5569 (N_5569,N_2120,N_2266);
and U5570 (N_5570,N_583,N_2825);
nor U5571 (N_5571,N_1174,N_2980);
nor U5572 (N_5572,N_984,N_2370);
and U5573 (N_5573,N_724,N_271);
nand U5574 (N_5574,N_851,N_1327);
nor U5575 (N_5575,N_2471,N_1);
nand U5576 (N_5576,N_23,N_724);
and U5577 (N_5577,N_2281,N_647);
nor U5578 (N_5578,N_1465,N_1775);
and U5579 (N_5579,N_935,N_2019);
nand U5580 (N_5580,N_2346,N_1601);
xnor U5581 (N_5581,N_1661,N_2929);
and U5582 (N_5582,N_2190,N_2798);
or U5583 (N_5583,N_129,N_2683);
nand U5584 (N_5584,N_254,N_1022);
and U5585 (N_5585,N_770,N_729);
and U5586 (N_5586,N_1701,N_126);
xor U5587 (N_5587,N_766,N_414);
or U5588 (N_5588,N_1273,N_60);
nand U5589 (N_5589,N_47,N_225);
and U5590 (N_5590,N_2798,N_278);
nor U5591 (N_5591,N_2162,N_2348);
xor U5592 (N_5592,N_1285,N_548);
nor U5593 (N_5593,N_2874,N_2312);
or U5594 (N_5594,N_2922,N_2067);
nor U5595 (N_5595,N_2569,N_2168);
and U5596 (N_5596,N_2950,N_2117);
xnor U5597 (N_5597,N_2572,N_2457);
and U5598 (N_5598,N_1086,N_2270);
or U5599 (N_5599,N_42,N_1085);
and U5600 (N_5600,N_1495,N_1165);
and U5601 (N_5601,N_133,N_2453);
and U5602 (N_5602,N_2183,N_1141);
or U5603 (N_5603,N_2439,N_1399);
or U5604 (N_5604,N_2967,N_486);
nor U5605 (N_5605,N_678,N_2547);
nor U5606 (N_5606,N_22,N_2736);
or U5607 (N_5607,N_502,N_1117);
nor U5608 (N_5608,N_1869,N_617);
nand U5609 (N_5609,N_590,N_2825);
nand U5610 (N_5610,N_1333,N_1659);
and U5611 (N_5611,N_1339,N_2614);
nor U5612 (N_5612,N_2544,N_1163);
nor U5613 (N_5613,N_42,N_412);
nand U5614 (N_5614,N_380,N_1519);
nor U5615 (N_5615,N_1241,N_783);
or U5616 (N_5616,N_1458,N_1815);
nor U5617 (N_5617,N_2274,N_472);
xnor U5618 (N_5618,N_1552,N_1404);
nor U5619 (N_5619,N_1240,N_8);
nand U5620 (N_5620,N_631,N_82);
and U5621 (N_5621,N_1032,N_2886);
nor U5622 (N_5622,N_1497,N_2890);
and U5623 (N_5623,N_767,N_1084);
and U5624 (N_5624,N_532,N_393);
xnor U5625 (N_5625,N_420,N_2607);
nand U5626 (N_5626,N_1255,N_614);
and U5627 (N_5627,N_2087,N_882);
nand U5628 (N_5628,N_1463,N_1477);
and U5629 (N_5629,N_518,N_2289);
nand U5630 (N_5630,N_53,N_1269);
and U5631 (N_5631,N_1047,N_1654);
nand U5632 (N_5632,N_2781,N_1419);
nor U5633 (N_5633,N_2143,N_2519);
nand U5634 (N_5634,N_2473,N_1260);
nand U5635 (N_5635,N_1867,N_2688);
nand U5636 (N_5636,N_203,N_1315);
nor U5637 (N_5637,N_1269,N_1908);
nand U5638 (N_5638,N_1424,N_731);
and U5639 (N_5639,N_2613,N_880);
and U5640 (N_5640,N_742,N_2817);
xor U5641 (N_5641,N_2734,N_1894);
and U5642 (N_5642,N_429,N_377);
and U5643 (N_5643,N_1574,N_219);
nand U5644 (N_5644,N_4,N_191);
and U5645 (N_5645,N_1454,N_9);
and U5646 (N_5646,N_2466,N_2225);
nor U5647 (N_5647,N_2458,N_2451);
xnor U5648 (N_5648,N_747,N_2497);
and U5649 (N_5649,N_1314,N_1196);
xor U5650 (N_5650,N_1814,N_1336);
or U5651 (N_5651,N_1154,N_628);
nor U5652 (N_5652,N_1589,N_2665);
nand U5653 (N_5653,N_1843,N_1397);
nand U5654 (N_5654,N_2156,N_1103);
and U5655 (N_5655,N_2552,N_1319);
xor U5656 (N_5656,N_1984,N_543);
or U5657 (N_5657,N_526,N_1172);
xor U5658 (N_5658,N_522,N_1168);
nor U5659 (N_5659,N_442,N_2558);
nor U5660 (N_5660,N_34,N_1064);
and U5661 (N_5661,N_731,N_1982);
nor U5662 (N_5662,N_553,N_120);
xor U5663 (N_5663,N_2863,N_2039);
and U5664 (N_5664,N_804,N_1263);
or U5665 (N_5665,N_1380,N_2755);
xor U5666 (N_5666,N_1369,N_2188);
or U5667 (N_5667,N_2627,N_2053);
nor U5668 (N_5668,N_1087,N_43);
and U5669 (N_5669,N_1967,N_394);
nand U5670 (N_5670,N_2527,N_455);
or U5671 (N_5671,N_2747,N_1182);
xor U5672 (N_5672,N_2371,N_2238);
nand U5673 (N_5673,N_1554,N_1019);
nand U5674 (N_5674,N_2895,N_1088);
or U5675 (N_5675,N_1402,N_611);
nor U5676 (N_5676,N_1048,N_1508);
and U5677 (N_5677,N_1308,N_2386);
and U5678 (N_5678,N_654,N_2847);
and U5679 (N_5679,N_1261,N_2895);
or U5680 (N_5680,N_2955,N_2391);
and U5681 (N_5681,N_2815,N_412);
nand U5682 (N_5682,N_2912,N_746);
nor U5683 (N_5683,N_2252,N_1763);
xor U5684 (N_5684,N_2751,N_2372);
and U5685 (N_5685,N_366,N_259);
nor U5686 (N_5686,N_2249,N_2713);
or U5687 (N_5687,N_193,N_1999);
nand U5688 (N_5688,N_2050,N_2727);
and U5689 (N_5689,N_1387,N_2458);
nor U5690 (N_5690,N_364,N_2590);
or U5691 (N_5691,N_2329,N_784);
nor U5692 (N_5692,N_560,N_186);
or U5693 (N_5693,N_2925,N_160);
nor U5694 (N_5694,N_2688,N_2598);
or U5695 (N_5695,N_904,N_12);
and U5696 (N_5696,N_2227,N_686);
xnor U5697 (N_5697,N_1294,N_950);
nand U5698 (N_5698,N_1357,N_1940);
nor U5699 (N_5699,N_1802,N_2655);
nand U5700 (N_5700,N_236,N_2862);
nand U5701 (N_5701,N_2524,N_2808);
or U5702 (N_5702,N_936,N_1405);
nor U5703 (N_5703,N_502,N_868);
xnor U5704 (N_5704,N_652,N_94);
nor U5705 (N_5705,N_2473,N_1014);
or U5706 (N_5706,N_2228,N_1508);
nor U5707 (N_5707,N_2182,N_1308);
nor U5708 (N_5708,N_1237,N_200);
xor U5709 (N_5709,N_397,N_2031);
nand U5710 (N_5710,N_2815,N_793);
xnor U5711 (N_5711,N_2446,N_880);
nor U5712 (N_5712,N_431,N_1291);
nor U5713 (N_5713,N_156,N_2955);
nand U5714 (N_5714,N_2520,N_1221);
or U5715 (N_5715,N_2957,N_2680);
nor U5716 (N_5716,N_1583,N_48);
or U5717 (N_5717,N_806,N_478);
or U5718 (N_5718,N_187,N_443);
xnor U5719 (N_5719,N_755,N_158);
or U5720 (N_5720,N_1295,N_2990);
or U5721 (N_5721,N_1173,N_2875);
xnor U5722 (N_5722,N_110,N_1541);
or U5723 (N_5723,N_2200,N_2196);
nor U5724 (N_5724,N_970,N_155);
nor U5725 (N_5725,N_2889,N_1350);
nor U5726 (N_5726,N_1106,N_471);
xor U5727 (N_5727,N_420,N_1585);
and U5728 (N_5728,N_778,N_317);
nand U5729 (N_5729,N_429,N_821);
nand U5730 (N_5730,N_2401,N_338);
nor U5731 (N_5731,N_2236,N_508);
nand U5732 (N_5732,N_2797,N_919);
nor U5733 (N_5733,N_2541,N_1127);
and U5734 (N_5734,N_2753,N_2848);
nand U5735 (N_5735,N_978,N_2641);
or U5736 (N_5736,N_2419,N_1966);
nor U5737 (N_5737,N_392,N_2276);
nand U5738 (N_5738,N_2314,N_1002);
nand U5739 (N_5739,N_1733,N_439);
and U5740 (N_5740,N_444,N_182);
and U5741 (N_5741,N_1102,N_2592);
nor U5742 (N_5742,N_2307,N_659);
and U5743 (N_5743,N_2668,N_600);
nor U5744 (N_5744,N_2485,N_902);
nand U5745 (N_5745,N_1790,N_2218);
or U5746 (N_5746,N_2029,N_197);
and U5747 (N_5747,N_1046,N_688);
xnor U5748 (N_5748,N_1343,N_2030);
or U5749 (N_5749,N_948,N_2634);
nand U5750 (N_5750,N_2236,N_1348);
or U5751 (N_5751,N_2211,N_953);
nor U5752 (N_5752,N_674,N_1084);
or U5753 (N_5753,N_986,N_2057);
and U5754 (N_5754,N_414,N_2750);
or U5755 (N_5755,N_897,N_2935);
xnor U5756 (N_5756,N_135,N_1402);
nand U5757 (N_5757,N_1057,N_2742);
and U5758 (N_5758,N_2846,N_2288);
and U5759 (N_5759,N_1492,N_974);
and U5760 (N_5760,N_78,N_1652);
nor U5761 (N_5761,N_1337,N_2707);
nor U5762 (N_5762,N_2696,N_81);
nor U5763 (N_5763,N_1158,N_681);
or U5764 (N_5764,N_1440,N_232);
or U5765 (N_5765,N_214,N_1227);
and U5766 (N_5766,N_229,N_1067);
and U5767 (N_5767,N_1639,N_2182);
and U5768 (N_5768,N_2022,N_2041);
nor U5769 (N_5769,N_2876,N_1379);
nor U5770 (N_5770,N_1419,N_653);
xor U5771 (N_5771,N_719,N_223);
or U5772 (N_5772,N_2566,N_2060);
xor U5773 (N_5773,N_1426,N_2143);
nand U5774 (N_5774,N_1277,N_1407);
nand U5775 (N_5775,N_1686,N_2449);
or U5776 (N_5776,N_1844,N_1048);
nand U5777 (N_5777,N_1061,N_649);
nand U5778 (N_5778,N_2430,N_1382);
and U5779 (N_5779,N_1603,N_1445);
nor U5780 (N_5780,N_2908,N_1165);
or U5781 (N_5781,N_237,N_286);
or U5782 (N_5782,N_2642,N_1185);
xnor U5783 (N_5783,N_2948,N_1643);
or U5784 (N_5784,N_2037,N_68);
nor U5785 (N_5785,N_172,N_1770);
xor U5786 (N_5786,N_2545,N_1695);
nand U5787 (N_5787,N_1300,N_1566);
and U5788 (N_5788,N_2841,N_2945);
xor U5789 (N_5789,N_809,N_1886);
and U5790 (N_5790,N_739,N_673);
or U5791 (N_5791,N_1603,N_2544);
nor U5792 (N_5792,N_1542,N_1062);
nand U5793 (N_5793,N_536,N_1126);
nor U5794 (N_5794,N_1190,N_1467);
and U5795 (N_5795,N_729,N_1277);
or U5796 (N_5796,N_145,N_1701);
or U5797 (N_5797,N_562,N_582);
nor U5798 (N_5798,N_1256,N_1833);
nor U5799 (N_5799,N_2533,N_175);
xnor U5800 (N_5800,N_2013,N_2513);
nor U5801 (N_5801,N_1510,N_2120);
nor U5802 (N_5802,N_373,N_37);
nand U5803 (N_5803,N_1279,N_2451);
or U5804 (N_5804,N_327,N_963);
or U5805 (N_5805,N_383,N_1172);
or U5806 (N_5806,N_2343,N_1562);
or U5807 (N_5807,N_351,N_2061);
nand U5808 (N_5808,N_71,N_2576);
xnor U5809 (N_5809,N_278,N_210);
nor U5810 (N_5810,N_1849,N_2557);
nor U5811 (N_5811,N_1606,N_404);
or U5812 (N_5812,N_1839,N_878);
and U5813 (N_5813,N_2505,N_194);
nand U5814 (N_5814,N_1658,N_1309);
and U5815 (N_5815,N_1155,N_2838);
xor U5816 (N_5816,N_1138,N_2648);
or U5817 (N_5817,N_3,N_1598);
nor U5818 (N_5818,N_664,N_2177);
and U5819 (N_5819,N_2900,N_1271);
and U5820 (N_5820,N_1485,N_54);
xnor U5821 (N_5821,N_989,N_2688);
nor U5822 (N_5822,N_1923,N_2416);
nand U5823 (N_5823,N_307,N_2438);
or U5824 (N_5824,N_530,N_1052);
xnor U5825 (N_5825,N_858,N_125);
nor U5826 (N_5826,N_5,N_1277);
xnor U5827 (N_5827,N_980,N_2746);
and U5828 (N_5828,N_2575,N_2887);
nor U5829 (N_5829,N_1649,N_277);
nand U5830 (N_5830,N_1361,N_278);
or U5831 (N_5831,N_1795,N_784);
xnor U5832 (N_5832,N_444,N_2824);
nor U5833 (N_5833,N_848,N_1317);
nor U5834 (N_5834,N_1339,N_2572);
nand U5835 (N_5835,N_1063,N_2030);
nor U5836 (N_5836,N_554,N_1369);
nor U5837 (N_5837,N_534,N_1054);
nand U5838 (N_5838,N_1736,N_2907);
or U5839 (N_5839,N_79,N_310);
or U5840 (N_5840,N_1440,N_265);
nor U5841 (N_5841,N_1921,N_95);
or U5842 (N_5842,N_1186,N_2393);
or U5843 (N_5843,N_2146,N_114);
nor U5844 (N_5844,N_2437,N_935);
nand U5845 (N_5845,N_2974,N_1980);
and U5846 (N_5846,N_715,N_869);
and U5847 (N_5847,N_916,N_1493);
nand U5848 (N_5848,N_64,N_686);
and U5849 (N_5849,N_1257,N_1874);
and U5850 (N_5850,N_553,N_1788);
nand U5851 (N_5851,N_110,N_1021);
and U5852 (N_5852,N_2490,N_2234);
or U5853 (N_5853,N_1413,N_836);
and U5854 (N_5854,N_270,N_512);
xnor U5855 (N_5855,N_8,N_235);
nor U5856 (N_5856,N_596,N_749);
nand U5857 (N_5857,N_640,N_2368);
nor U5858 (N_5858,N_751,N_781);
xnor U5859 (N_5859,N_2230,N_807);
and U5860 (N_5860,N_1833,N_84);
nand U5861 (N_5861,N_75,N_1069);
nor U5862 (N_5862,N_2617,N_2202);
nand U5863 (N_5863,N_2415,N_694);
nand U5864 (N_5864,N_575,N_2902);
nand U5865 (N_5865,N_326,N_1211);
or U5866 (N_5866,N_191,N_1942);
nor U5867 (N_5867,N_2590,N_2458);
nor U5868 (N_5868,N_621,N_910);
nor U5869 (N_5869,N_1687,N_584);
nand U5870 (N_5870,N_1134,N_1432);
nand U5871 (N_5871,N_626,N_1190);
or U5872 (N_5872,N_1608,N_1083);
or U5873 (N_5873,N_2543,N_250);
nand U5874 (N_5874,N_893,N_57);
and U5875 (N_5875,N_1477,N_1748);
xnor U5876 (N_5876,N_40,N_2639);
nor U5877 (N_5877,N_1923,N_2263);
nor U5878 (N_5878,N_42,N_323);
or U5879 (N_5879,N_2641,N_2482);
xnor U5880 (N_5880,N_2356,N_872);
or U5881 (N_5881,N_844,N_1252);
xnor U5882 (N_5882,N_376,N_1897);
and U5883 (N_5883,N_1748,N_2677);
or U5884 (N_5884,N_1771,N_2870);
nand U5885 (N_5885,N_763,N_2400);
and U5886 (N_5886,N_1158,N_1066);
nand U5887 (N_5887,N_1240,N_2448);
nand U5888 (N_5888,N_572,N_2786);
nor U5889 (N_5889,N_2233,N_101);
xor U5890 (N_5890,N_640,N_1710);
and U5891 (N_5891,N_2669,N_627);
or U5892 (N_5892,N_447,N_2106);
and U5893 (N_5893,N_1508,N_1318);
nand U5894 (N_5894,N_1080,N_1274);
nand U5895 (N_5895,N_1500,N_1927);
or U5896 (N_5896,N_1959,N_394);
and U5897 (N_5897,N_2477,N_832);
and U5898 (N_5898,N_1596,N_1440);
nor U5899 (N_5899,N_859,N_1301);
nand U5900 (N_5900,N_307,N_578);
nand U5901 (N_5901,N_2373,N_2251);
or U5902 (N_5902,N_496,N_1349);
xnor U5903 (N_5903,N_2896,N_2763);
nand U5904 (N_5904,N_1104,N_1523);
or U5905 (N_5905,N_914,N_1071);
and U5906 (N_5906,N_1982,N_853);
nor U5907 (N_5907,N_341,N_2648);
or U5908 (N_5908,N_2789,N_1861);
nor U5909 (N_5909,N_1175,N_2547);
and U5910 (N_5910,N_1810,N_2711);
or U5911 (N_5911,N_1916,N_2643);
or U5912 (N_5912,N_2827,N_785);
nor U5913 (N_5913,N_1886,N_33);
nand U5914 (N_5914,N_918,N_869);
and U5915 (N_5915,N_2148,N_1881);
or U5916 (N_5916,N_1963,N_917);
nand U5917 (N_5917,N_425,N_1657);
nand U5918 (N_5918,N_1885,N_1418);
and U5919 (N_5919,N_1050,N_1694);
and U5920 (N_5920,N_1286,N_943);
xnor U5921 (N_5921,N_2697,N_1963);
and U5922 (N_5922,N_1391,N_961);
or U5923 (N_5923,N_2906,N_363);
nand U5924 (N_5924,N_626,N_2772);
nor U5925 (N_5925,N_461,N_2949);
xor U5926 (N_5926,N_1969,N_1368);
xor U5927 (N_5927,N_912,N_1119);
nand U5928 (N_5928,N_1046,N_1497);
nand U5929 (N_5929,N_1668,N_2851);
nand U5930 (N_5930,N_793,N_1137);
nand U5931 (N_5931,N_1270,N_1538);
or U5932 (N_5932,N_2659,N_2090);
or U5933 (N_5933,N_157,N_2084);
nor U5934 (N_5934,N_2146,N_2651);
nor U5935 (N_5935,N_2357,N_2006);
or U5936 (N_5936,N_796,N_1737);
or U5937 (N_5937,N_2912,N_2721);
nand U5938 (N_5938,N_775,N_650);
nand U5939 (N_5939,N_942,N_128);
nor U5940 (N_5940,N_6,N_2030);
and U5941 (N_5941,N_1861,N_1551);
nor U5942 (N_5942,N_1141,N_632);
nor U5943 (N_5943,N_20,N_1725);
nand U5944 (N_5944,N_2262,N_118);
nand U5945 (N_5945,N_2984,N_1251);
nand U5946 (N_5946,N_716,N_563);
nor U5947 (N_5947,N_2544,N_1175);
or U5948 (N_5948,N_1520,N_1128);
nor U5949 (N_5949,N_2291,N_2583);
or U5950 (N_5950,N_2608,N_2760);
nor U5951 (N_5951,N_2772,N_1310);
nand U5952 (N_5952,N_1278,N_2185);
and U5953 (N_5953,N_1878,N_1984);
nor U5954 (N_5954,N_1614,N_985);
or U5955 (N_5955,N_1304,N_701);
xnor U5956 (N_5956,N_346,N_363);
nor U5957 (N_5957,N_2416,N_2041);
nor U5958 (N_5958,N_1927,N_997);
or U5959 (N_5959,N_1286,N_661);
nor U5960 (N_5960,N_2726,N_2972);
or U5961 (N_5961,N_1835,N_2910);
xnor U5962 (N_5962,N_593,N_1806);
nor U5963 (N_5963,N_1360,N_2891);
xor U5964 (N_5964,N_1688,N_55);
and U5965 (N_5965,N_2388,N_80);
nand U5966 (N_5966,N_1948,N_598);
xnor U5967 (N_5967,N_530,N_549);
and U5968 (N_5968,N_2415,N_455);
or U5969 (N_5969,N_2390,N_2540);
and U5970 (N_5970,N_2610,N_2931);
nand U5971 (N_5971,N_1487,N_1259);
and U5972 (N_5972,N_1074,N_2766);
and U5973 (N_5973,N_349,N_1780);
or U5974 (N_5974,N_1401,N_2650);
nand U5975 (N_5975,N_2475,N_1196);
xor U5976 (N_5976,N_1571,N_2436);
nand U5977 (N_5977,N_2738,N_2517);
nor U5978 (N_5978,N_219,N_1991);
nand U5979 (N_5979,N_2228,N_551);
nor U5980 (N_5980,N_301,N_1743);
nand U5981 (N_5981,N_1386,N_2741);
nand U5982 (N_5982,N_2994,N_2421);
and U5983 (N_5983,N_1553,N_791);
nand U5984 (N_5984,N_1135,N_2806);
and U5985 (N_5985,N_1573,N_2542);
nor U5986 (N_5986,N_636,N_444);
or U5987 (N_5987,N_32,N_2536);
and U5988 (N_5988,N_1176,N_1194);
nand U5989 (N_5989,N_2259,N_957);
nand U5990 (N_5990,N_2830,N_1196);
or U5991 (N_5991,N_1682,N_891);
and U5992 (N_5992,N_2968,N_1934);
or U5993 (N_5993,N_1064,N_2094);
xor U5994 (N_5994,N_2578,N_863);
nor U5995 (N_5995,N_2049,N_799);
nor U5996 (N_5996,N_1101,N_2807);
and U5997 (N_5997,N_1078,N_2914);
nand U5998 (N_5998,N_2797,N_2548);
and U5999 (N_5999,N_621,N_1932);
and U6000 (N_6000,N_4308,N_4149);
nand U6001 (N_6001,N_4634,N_3194);
and U6002 (N_6002,N_3728,N_5992);
and U6003 (N_6003,N_4258,N_3958);
nor U6004 (N_6004,N_3892,N_5615);
or U6005 (N_6005,N_4107,N_5398);
or U6006 (N_6006,N_3817,N_5850);
or U6007 (N_6007,N_4850,N_5065);
and U6008 (N_6008,N_4586,N_5784);
nor U6009 (N_6009,N_4075,N_3718);
nor U6010 (N_6010,N_5549,N_5369);
nor U6011 (N_6011,N_3212,N_5002);
nand U6012 (N_6012,N_5883,N_3582);
xnor U6013 (N_6013,N_3167,N_5930);
nand U6014 (N_6014,N_5163,N_3477);
nor U6015 (N_6015,N_5162,N_3013);
nand U6016 (N_6016,N_4895,N_5942);
and U6017 (N_6017,N_5351,N_4282);
and U6018 (N_6018,N_5121,N_4576);
or U6019 (N_6019,N_3573,N_4709);
or U6020 (N_6020,N_3229,N_3150);
and U6021 (N_6021,N_4114,N_5757);
nor U6022 (N_6022,N_4867,N_4876);
xnor U6023 (N_6023,N_4838,N_4321);
nor U6024 (N_6024,N_5200,N_5935);
and U6025 (N_6025,N_4715,N_3609);
xor U6026 (N_6026,N_3327,N_5439);
xnor U6027 (N_6027,N_4824,N_4920);
nor U6028 (N_6028,N_5299,N_4507);
xor U6029 (N_6029,N_4285,N_5462);
nand U6030 (N_6030,N_5035,N_3767);
nand U6031 (N_6031,N_3702,N_5740);
nand U6032 (N_6032,N_5262,N_3562);
nor U6033 (N_6033,N_4869,N_3207);
and U6034 (N_6034,N_4662,N_5073);
and U6035 (N_6035,N_5739,N_5920);
or U6036 (N_6036,N_3084,N_3317);
nand U6037 (N_6037,N_5683,N_4029);
nor U6038 (N_6038,N_4394,N_5341);
or U6039 (N_6039,N_5018,N_3657);
and U6040 (N_6040,N_4427,N_3650);
nor U6041 (N_6041,N_4874,N_4121);
and U6042 (N_6042,N_4601,N_5653);
nand U6043 (N_6043,N_4994,N_3070);
and U6044 (N_6044,N_4015,N_4133);
and U6045 (N_6045,N_4281,N_4698);
and U6046 (N_6046,N_4857,N_5787);
and U6047 (N_6047,N_3022,N_3060);
xnor U6048 (N_6048,N_3242,N_4080);
nand U6049 (N_6049,N_4441,N_4305);
or U6050 (N_6050,N_3587,N_5958);
and U6051 (N_6051,N_4273,N_4078);
nor U6052 (N_6052,N_5088,N_5005);
and U6053 (N_6053,N_3062,N_5959);
nor U6054 (N_6054,N_4521,N_3899);
nor U6055 (N_6055,N_3680,N_3162);
and U6056 (N_6056,N_3402,N_4546);
nand U6057 (N_6057,N_5913,N_5168);
and U6058 (N_6058,N_3119,N_3190);
nand U6059 (N_6059,N_4971,N_3875);
nand U6060 (N_6060,N_3638,N_4620);
or U6061 (N_6061,N_3542,N_5633);
nor U6062 (N_6062,N_5180,N_3646);
nor U6063 (N_6063,N_3482,N_5228);
and U6064 (N_6064,N_4729,N_4203);
nand U6065 (N_6065,N_4645,N_3129);
xnor U6066 (N_6066,N_4218,N_3637);
nor U6067 (N_6067,N_4678,N_4239);
and U6068 (N_6068,N_3065,N_4062);
or U6069 (N_6069,N_5489,N_4621);
nand U6070 (N_6070,N_3803,N_4598);
and U6071 (N_6071,N_4828,N_5310);
and U6072 (N_6072,N_3806,N_4243);
nand U6073 (N_6073,N_4437,N_5177);
nor U6074 (N_6074,N_4201,N_3641);
nor U6075 (N_6075,N_5790,N_3854);
and U6076 (N_6076,N_5379,N_5526);
and U6077 (N_6077,N_3350,N_4632);
nand U6078 (N_6078,N_4884,N_4152);
nand U6079 (N_6079,N_3225,N_3669);
nor U6080 (N_6080,N_3213,N_5902);
nor U6081 (N_6081,N_5539,N_5225);
or U6082 (N_6082,N_5700,N_5105);
nand U6083 (N_6083,N_3157,N_3300);
xnor U6084 (N_6084,N_5270,N_3965);
or U6085 (N_6085,N_3451,N_5258);
and U6086 (N_6086,N_4405,N_5721);
nand U6087 (N_6087,N_5362,N_5662);
nor U6088 (N_6088,N_3596,N_5911);
nand U6089 (N_6089,N_5976,N_3253);
nor U6090 (N_6090,N_4271,N_4186);
and U6091 (N_6091,N_4949,N_4241);
nand U6092 (N_6092,N_5785,N_4446);
or U6093 (N_6093,N_5630,N_3987);
and U6094 (N_6094,N_3309,N_4060);
or U6095 (N_6095,N_5160,N_5907);
nand U6096 (N_6096,N_4820,N_3860);
or U6097 (N_6097,N_3107,N_5422);
nand U6098 (N_6098,N_4347,N_3967);
and U6099 (N_6099,N_5954,N_3124);
nand U6100 (N_6100,N_3238,N_4624);
nor U6101 (N_6101,N_3090,N_5860);
and U6102 (N_6102,N_5857,N_5754);
xor U6103 (N_6103,N_5839,N_3307);
and U6104 (N_6104,N_5364,N_5540);
or U6105 (N_6105,N_5557,N_5908);
or U6106 (N_6106,N_4848,N_3594);
nand U6107 (N_6107,N_5309,N_4320);
xnor U6108 (N_6108,N_5034,N_4140);
xnor U6109 (N_6109,N_4897,N_4061);
and U6110 (N_6110,N_5553,N_3962);
and U6111 (N_6111,N_4980,N_4726);
nand U6112 (N_6112,N_5933,N_3068);
nand U6113 (N_6113,N_4623,N_3362);
nand U6114 (N_6114,N_3017,N_3618);
nand U6115 (N_6115,N_4786,N_5014);
nor U6116 (N_6116,N_4115,N_3106);
nand U6117 (N_6117,N_3290,N_4333);
nor U6118 (N_6118,N_5409,N_5676);
nor U6119 (N_6119,N_3230,N_4537);
or U6120 (N_6120,N_4759,N_3308);
nand U6121 (N_6121,N_3600,N_3415);
nand U6122 (N_6122,N_5811,N_5519);
xor U6123 (N_6123,N_4111,N_4083);
or U6124 (N_6124,N_3649,N_3580);
and U6125 (N_6125,N_3864,N_4192);
and U6126 (N_6126,N_5000,N_3531);
xor U6127 (N_6127,N_5010,N_5273);
and U6128 (N_6128,N_5244,N_5541);
nor U6129 (N_6129,N_4360,N_3581);
or U6130 (N_6130,N_4068,N_3012);
nor U6131 (N_6131,N_5871,N_4932);
nor U6132 (N_6132,N_3489,N_5891);
nor U6133 (N_6133,N_3696,N_5607);
or U6134 (N_6134,N_4292,N_4578);
nor U6135 (N_6135,N_4334,N_5516);
nor U6136 (N_6136,N_3087,N_3622);
nand U6137 (N_6137,N_5138,N_5900);
nor U6138 (N_6138,N_4113,N_4081);
nor U6139 (N_6139,N_3935,N_5190);
xnor U6140 (N_6140,N_3683,N_3430);
xor U6141 (N_6141,N_5484,N_3786);
and U6142 (N_6142,N_3567,N_4556);
or U6143 (N_6143,N_5815,N_5695);
nor U6144 (N_6144,N_4501,N_3282);
xnor U6145 (N_6145,N_5142,N_4633);
nor U6146 (N_6146,N_4010,N_3839);
nor U6147 (N_6147,N_4480,N_3697);
nor U6148 (N_6148,N_3805,N_5550);
or U6149 (N_6149,N_3976,N_5892);
and U6150 (N_6150,N_3333,N_5674);
and U6151 (N_6151,N_3994,N_4675);
nor U6152 (N_6152,N_5361,N_3170);
and U6153 (N_6153,N_4278,N_4942);
nor U6154 (N_6154,N_4963,N_3037);
nand U6155 (N_6155,N_4640,N_3069);
nand U6156 (N_6156,N_5703,N_3930);
or U6157 (N_6157,N_4102,N_5631);
nand U6158 (N_6158,N_5457,N_4560);
or U6159 (N_6159,N_5473,N_4513);
nor U6160 (N_6160,N_4154,N_5347);
nand U6161 (N_6161,N_4159,N_4772);
and U6162 (N_6162,N_3050,N_5094);
xnor U6163 (N_6163,N_3841,N_5611);
nor U6164 (N_6164,N_4065,N_4390);
or U6165 (N_6165,N_4656,N_5461);
nand U6166 (N_6166,N_3948,N_3874);
and U6167 (N_6167,N_4177,N_5146);
xnor U6168 (N_6168,N_3432,N_4082);
and U6169 (N_6169,N_4473,N_5029);
nor U6170 (N_6170,N_5050,N_5229);
xor U6171 (N_6171,N_5127,N_4315);
and U6172 (N_6172,N_4089,N_3706);
and U6173 (N_6173,N_3957,N_3407);
and U6174 (N_6174,N_5720,N_5944);
nor U6175 (N_6175,N_5020,N_4479);
and U6176 (N_6176,N_3329,N_3387);
nor U6177 (N_6177,N_5603,N_5292);
or U6178 (N_6178,N_5670,N_4855);
xor U6179 (N_6179,N_5922,N_5556);
nor U6180 (N_6180,N_5036,N_5904);
and U6181 (N_6181,N_4485,N_5325);
xnor U6182 (N_6182,N_5885,N_3919);
nand U6183 (N_6183,N_5288,N_4749);
nand U6184 (N_6184,N_5305,N_5404);
nand U6185 (N_6185,N_5338,N_3501);
or U6186 (N_6186,N_3078,N_5345);
or U6187 (N_6187,N_4276,N_5008);
nand U6188 (N_6188,N_5421,N_4669);
nand U6189 (N_6189,N_4727,N_3742);
and U6190 (N_6190,N_4930,N_5108);
nor U6191 (N_6191,N_4907,N_5781);
xor U6192 (N_6192,N_3131,N_3274);
and U6193 (N_6193,N_5972,N_4033);
nor U6194 (N_6194,N_4288,N_3708);
or U6195 (N_6195,N_3798,N_4826);
nand U6196 (N_6196,N_3373,N_4407);
or U6197 (N_6197,N_3104,N_5934);
nor U6198 (N_6198,N_3904,N_3031);
nand U6199 (N_6199,N_4805,N_5834);
and U6200 (N_6200,N_5508,N_5803);
nor U6201 (N_6201,N_5284,N_4468);
and U6202 (N_6202,N_5434,N_5620);
xnor U6203 (N_6203,N_3406,N_5775);
nor U6204 (N_6204,N_4522,N_5873);
nand U6205 (N_6205,N_4377,N_4067);
nand U6206 (N_6206,N_4782,N_5593);
or U6207 (N_6207,N_5650,N_4684);
and U6208 (N_6208,N_3054,N_3789);
nand U6209 (N_6209,N_5322,N_4500);
or U6210 (N_6210,N_3115,N_5753);
or U6211 (N_6211,N_4663,N_3419);
xor U6212 (N_6212,N_3156,N_4565);
xor U6213 (N_6213,N_3003,N_5329);
or U6214 (N_6214,N_3142,N_5802);
or U6215 (N_6215,N_5081,N_4999);
nor U6216 (N_6216,N_5965,N_3945);
nand U6217 (N_6217,N_5664,N_4156);
nor U6218 (N_6218,N_3660,N_5818);
or U6219 (N_6219,N_3818,N_5690);
xor U6220 (N_6220,N_3335,N_3429);
nor U6221 (N_6221,N_3653,N_4451);
nand U6222 (N_6222,N_5101,N_4572);
or U6223 (N_6223,N_3296,N_5048);
or U6224 (N_6224,N_3952,N_3859);
nor U6225 (N_6225,N_3739,N_5246);
nor U6226 (N_6226,N_4969,N_5814);
or U6227 (N_6227,N_3145,N_5438);
or U6228 (N_6228,N_4412,N_5278);
or U6229 (N_6229,N_3399,N_5788);
nand U6230 (N_6230,N_4584,N_4738);
nand U6231 (N_6231,N_4606,N_4246);
or U6232 (N_6232,N_3937,N_4331);
and U6233 (N_6233,N_5232,N_4872);
or U6234 (N_6234,N_3357,N_5012);
and U6235 (N_6235,N_5715,N_4823);
or U6236 (N_6236,N_5576,N_3487);
nor U6237 (N_6237,N_5429,N_3584);
nand U6238 (N_6238,N_4048,N_5119);
nand U6239 (N_6239,N_5668,N_5241);
or U6240 (N_6240,N_3227,N_5209);
nor U6241 (N_6241,N_4696,N_5170);
nor U6242 (N_6242,N_5497,N_4854);
xnor U6243 (N_6243,N_5819,N_3990);
and U6244 (N_6244,N_4842,N_5365);
nor U6245 (N_6245,N_5263,N_5730);
nor U6246 (N_6246,N_5779,N_5875);
nor U6247 (N_6247,N_3291,N_4797);
or U6248 (N_6248,N_3187,N_3098);
nand U6249 (N_6249,N_3725,N_4732);
nor U6250 (N_6250,N_3809,N_5331);
nor U6251 (N_6251,N_5407,N_4743);
xor U6252 (N_6252,N_5382,N_4450);
nand U6253 (N_6253,N_4227,N_5182);
xor U6254 (N_6254,N_4520,N_5712);
nor U6255 (N_6255,N_3030,N_3143);
nor U6256 (N_6256,N_3160,N_4349);
nand U6257 (N_6257,N_5054,N_4958);
nor U6258 (N_6258,N_5713,N_5978);
or U6259 (N_6259,N_5886,N_4922);
nor U6260 (N_6260,N_4224,N_3738);
and U6261 (N_6261,N_4351,N_5584);
and U6262 (N_6262,N_5371,N_3393);
nand U6263 (N_6263,N_3521,N_5183);
and U6264 (N_6264,N_4272,N_5966);
xor U6265 (N_6265,N_4938,N_3993);
xor U6266 (N_6266,N_3231,N_4919);
or U6267 (N_6267,N_3627,N_5080);
or U6268 (N_6268,N_4814,N_3804);
or U6269 (N_6269,N_3729,N_5264);
and U6270 (N_6270,N_5372,N_3223);
nand U6271 (N_6271,N_5558,N_4723);
nand U6272 (N_6272,N_4187,N_4466);
nand U6273 (N_6273,N_5657,N_3502);
and U6274 (N_6274,N_4505,N_4460);
nand U6275 (N_6275,N_3028,N_4040);
and U6276 (N_6276,N_3204,N_4753);
and U6277 (N_6277,N_5570,N_4983);
and U6278 (N_6278,N_4801,N_3960);
and U6279 (N_6279,N_4209,N_4178);
nor U6280 (N_6280,N_5103,N_3845);
and U6281 (N_6281,N_4045,N_5145);
or U6282 (N_6282,N_4184,N_5019);
nor U6283 (N_6283,N_5301,N_3447);
or U6284 (N_6284,N_5252,N_5004);
xnor U6285 (N_6285,N_4954,N_5852);
or U6286 (N_6286,N_4052,N_4936);
nor U6287 (N_6287,N_5076,N_5465);
or U6288 (N_6288,N_5193,N_3799);
nand U6289 (N_6289,N_3422,N_4204);
and U6290 (N_6290,N_4998,N_5843);
and U6291 (N_6291,N_4385,N_4366);
nor U6292 (N_6292,N_5166,N_4103);
and U6293 (N_6293,N_3464,N_4885);
and U6294 (N_6294,N_3936,N_3511);
nor U6295 (N_6295,N_3108,N_4170);
or U6296 (N_6296,N_5504,N_5043);
and U6297 (N_6297,N_3975,N_5426);
nand U6298 (N_6298,N_3360,N_5537);
nand U6299 (N_6299,N_5996,N_3826);
or U6300 (N_6300,N_4087,N_5280);
nand U6301 (N_6301,N_4094,N_4299);
or U6302 (N_6302,N_3908,N_4235);
or U6303 (N_6303,N_3568,N_4055);
nor U6304 (N_6304,N_3716,N_4134);
and U6305 (N_6305,N_4760,N_3301);
or U6306 (N_6306,N_5923,N_3754);
nor U6307 (N_6307,N_3916,N_5235);
nor U6308 (N_6308,N_5172,N_3825);
nor U6309 (N_6309,N_4582,N_5468);
and U6310 (N_6310,N_3304,N_5092);
or U6311 (N_6311,N_5981,N_4311);
nor U6312 (N_6312,N_5420,N_3286);
or U6313 (N_6313,N_3784,N_3883);
or U6314 (N_6314,N_3232,N_4242);
and U6315 (N_6315,N_5027,N_4099);
and U6316 (N_6316,N_5799,N_3785);
and U6317 (N_6317,N_4918,N_3113);
nand U6318 (N_6318,N_5955,N_4791);
and U6319 (N_6319,N_5298,N_4630);
nor U6320 (N_6320,N_5805,N_3214);
nor U6321 (N_6321,N_4843,N_3514);
nand U6322 (N_6322,N_4910,N_3695);
nor U6323 (N_6323,N_3436,N_4042);
nand U6324 (N_6324,N_4637,N_3281);
and U6325 (N_6325,N_3849,N_3614);
or U6326 (N_6326,N_3759,N_3893);
or U6327 (N_6327,N_5718,N_3135);
or U6328 (N_6328,N_3118,N_5711);
nand U6329 (N_6329,N_3338,N_5868);
or U6330 (N_6330,N_3655,N_4792);
xnor U6331 (N_6331,N_3966,N_5095);
or U6332 (N_6332,N_4638,N_4141);
or U6333 (N_6333,N_3540,N_4497);
and U6334 (N_6334,N_5865,N_5964);
or U6335 (N_6335,N_3733,N_5949);
nand U6336 (N_6336,N_4966,N_5068);
xnor U6337 (N_6337,N_5245,N_4325);
nor U6338 (N_6338,N_5030,N_3983);
or U6339 (N_6339,N_4336,N_3457);
xor U6340 (N_6340,N_3671,N_4771);
xor U6341 (N_6341,N_4145,N_5460);
nand U6342 (N_6342,N_3132,N_4266);
nand U6343 (N_6343,N_3101,N_4551);
or U6344 (N_6344,N_4472,N_3710);
nand U6345 (N_6345,N_3195,N_3424);
nor U6346 (N_6346,N_3389,N_5303);
nand U6347 (N_6347,N_4986,N_3298);
nor U6348 (N_6348,N_5872,N_3698);
nand U6349 (N_6349,N_5137,N_4197);
xnor U6350 (N_6350,N_4532,N_4138);
and U6351 (N_6351,N_5474,N_4515);
nor U6352 (N_6352,N_3868,N_4713);
nor U6353 (N_6353,N_3985,N_4364);
xor U6354 (N_6354,N_4737,N_5893);
nand U6355 (N_6355,N_5842,N_3134);
or U6356 (N_6356,N_5941,N_3867);
xnor U6357 (N_6357,N_4461,N_4914);
nand U6358 (N_6358,N_3814,N_3063);
nor U6359 (N_6359,N_5637,N_3963);
and U6360 (N_6360,N_4379,N_5367);
or U6361 (N_6361,N_3557,N_3171);
or U6362 (N_6362,N_3446,N_3210);
and U6363 (N_6363,N_3968,N_4761);
or U6364 (N_6364,N_3626,N_3316);
xor U6365 (N_6365,N_5441,N_3388);
nand U6366 (N_6366,N_3326,N_5988);
and U6367 (N_6367,N_3492,N_5275);
nor U6368 (N_6368,N_4395,N_3876);
xor U6369 (N_6369,N_5250,N_4649);
xnor U6370 (N_6370,N_3576,N_5311);
and U6371 (N_6371,N_3163,N_3510);
xnor U6372 (N_6372,N_3005,N_5074);
and U6373 (N_6373,N_3828,N_3894);
nor U6374 (N_6374,N_4552,N_3746);
and U6375 (N_6375,N_4193,N_5414);
nand U6376 (N_6376,N_3041,N_3349);
nor U6377 (N_6377,N_3453,N_3973);
or U6378 (N_6378,N_4039,N_5026);
nor U6379 (N_6379,N_3148,N_4631);
and U6380 (N_6380,N_5247,N_4350);
or U6381 (N_6381,N_3233,N_3589);
xnor U6382 (N_6382,N_4063,N_4000);
or U6383 (N_6383,N_4416,N_5614);
nand U6384 (N_6384,N_5751,N_4007);
nor U6385 (N_6385,N_4886,N_4686);
or U6386 (N_6386,N_4770,N_4345);
xnor U6387 (N_6387,N_3268,N_3885);
nand U6388 (N_6388,N_3097,N_4400);
nand U6389 (N_6389,N_4973,N_3775);
and U6390 (N_6390,N_4355,N_5684);
or U6391 (N_6391,N_5406,N_3761);
nor U6392 (N_6392,N_5878,N_5906);
xor U6393 (N_6393,N_4027,N_3052);
xnor U6394 (N_6394,N_3992,N_4112);
or U6395 (N_6395,N_4362,N_5268);
and U6396 (N_6396,N_3656,N_5510);
or U6397 (N_6397,N_3982,N_5658);
and U6398 (N_6398,N_5534,N_4084);
nand U6399 (N_6399,N_5667,N_4579);
nor U6400 (N_6400,N_3321,N_4525);
or U6401 (N_6401,N_3459,N_5741);
nor U6402 (N_6402,N_3259,N_3408);
nor U6403 (N_6403,N_4744,N_4066);
or U6404 (N_6404,N_5506,N_3347);
nand U6405 (N_6405,N_3640,N_5673);
nor U6406 (N_6406,N_4859,N_3048);
or U6407 (N_6407,N_3400,N_5618);
or U6408 (N_6408,N_5496,N_5525);
xnor U6409 (N_6409,N_4787,N_5300);
nor U6410 (N_6410,N_3159,N_3203);
nand U6411 (N_6411,N_5638,N_5986);
nor U6412 (N_6412,N_5249,N_4896);
nor U6413 (N_6413,N_3155,N_3959);
or U6414 (N_6414,N_4798,N_5478);
nand U6415 (N_6415,N_3625,N_5471);
and U6416 (N_6416,N_3865,N_5479);
or U6417 (N_6417,N_3125,N_5122);
and U6418 (N_6418,N_5223,N_5380);
nor U6419 (N_6419,N_4636,N_5354);
nand U6420 (N_6420,N_3763,N_4599);
and U6421 (N_6421,N_4322,N_4674);
or U6422 (N_6422,N_4987,N_3032);
or U6423 (N_6423,N_3917,N_4875);
and U6424 (N_6424,N_3319,N_3271);
or U6425 (N_6425,N_4455,N_5493);
nor U6426 (N_6426,N_4766,N_5449);
and U6427 (N_6427,N_5856,N_3096);
and U6428 (N_6428,N_5387,N_3503);
nand U6429 (N_6429,N_3218,N_3964);
nor U6430 (N_6430,N_3216,N_3456);
nor U6431 (N_6431,N_3416,N_3010);
nor U6432 (N_6432,N_5574,N_4701);
nor U6433 (N_6433,N_5109,N_5957);
nor U6434 (N_6434,N_3234,N_5780);
and U6435 (N_6435,N_4244,N_3621);
nand U6436 (N_6436,N_3256,N_5987);
nor U6437 (N_6437,N_3025,N_5656);
nor U6438 (N_6438,N_3693,N_3377);
nand U6439 (N_6439,N_3020,N_5825);
nand U6440 (N_6440,N_3991,N_4700);
or U6441 (N_6441,N_4297,N_3297);
and U6442 (N_6442,N_5271,N_3493);
and U6443 (N_6443,N_4712,N_4799);
or U6444 (N_6444,N_3922,N_3394);
and U6445 (N_6445,N_4423,N_5107);
nand U6446 (N_6446,N_4035,N_3033);
nor U6447 (N_6447,N_5764,N_3659);
or U6448 (N_6448,N_4452,N_4720);
nor U6449 (N_6449,N_3665,N_3942);
nor U6450 (N_6450,N_5343,N_4736);
nand U6451 (N_6451,N_4238,N_3611);
and U6452 (N_6452,N_5204,N_3343);
or U6453 (N_6453,N_4871,N_5702);
and U6454 (N_6454,N_3490,N_5359);
and U6455 (N_6455,N_5123,N_5100);
and U6456 (N_6456,N_5577,N_5686);
nor U6457 (N_6457,N_5826,N_5905);
nor U6458 (N_6458,N_4458,N_3586);
nand U6459 (N_6459,N_3925,N_4495);
or U6460 (N_6460,N_4742,N_4264);
nor U6461 (N_6461,N_4383,N_3369);
and U6462 (N_6462,N_3314,N_4563);
nand U6463 (N_6463,N_4758,N_4221);
or U6464 (N_6464,N_3497,N_3367);
nor U6465 (N_6465,N_4142,N_5151);
and U6466 (N_6466,N_5175,N_3224);
nor U6467 (N_6467,N_4573,N_3591);
or U6468 (N_6468,N_4290,N_4677);
xnor U6469 (N_6469,N_5219,N_5486);
and U6470 (N_6470,N_3525,N_5091);
and U6471 (N_6471,N_3024,N_4536);
and U6472 (N_6472,N_3601,N_3872);
nand U6473 (N_6473,N_5357,N_4526);
nor U6474 (N_6474,N_5112,N_5897);
nor U6475 (N_6475,N_4506,N_5234);
nand U6476 (N_6476,N_3452,N_3133);
or U6477 (N_6477,N_3272,N_3687);
or U6478 (N_6478,N_4157,N_4931);
nand U6479 (N_6479,N_3743,N_3642);
nand U6480 (N_6480,N_4127,N_4550);
or U6481 (N_6481,N_4471,N_3014);
or U6482 (N_6482,N_4916,N_4459);
nor U6483 (N_6483,N_3535,N_3479);
nand U6484 (N_6484,N_3427,N_4207);
and U6485 (N_6485,N_5423,N_5220);
or U6486 (N_6486,N_5257,N_4194);
nor U6487 (N_6487,N_5385,N_3509);
and U6488 (N_6488,N_5613,N_3411);
nor U6489 (N_6489,N_5833,N_4449);
nand U6490 (N_6490,N_4891,N_3774);
and U6491 (N_6491,N_3284,N_3295);
nor U6492 (N_6492,N_4893,N_5882);
and U6493 (N_6493,N_3154,N_5279);
and U6494 (N_6494,N_3252,N_4417);
and U6495 (N_6495,N_5679,N_4047);
nor U6496 (N_6496,N_3907,N_3927);
xor U6497 (N_6497,N_3658,N_3720);
or U6498 (N_6498,N_5417,N_5015);
or U6499 (N_6499,N_4981,N_5645);
and U6500 (N_6500,N_5946,N_3328);
and U6501 (N_6501,N_5236,N_5055);
or U6502 (N_6502,N_4924,N_4293);
or U6503 (N_6503,N_3353,N_4212);
and U6504 (N_6504,N_4167,N_3635);
nand U6505 (N_6505,N_4804,N_3201);
nand U6506 (N_6506,N_4935,N_5596);
or U6507 (N_6507,N_5761,N_3794);
nand U6508 (N_6508,N_5635,N_4927);
xor U6509 (N_6509,N_4323,N_5436);
and U6510 (N_6510,N_5836,N_4289);
or U6511 (N_6511,N_4251,N_4868);
and U6512 (N_6512,N_4908,N_3534);
and U6513 (N_6513,N_3895,N_5625);
nor U6514 (N_6514,N_5410,N_5016);
nor U6515 (N_6515,N_5998,N_3473);
nand U6516 (N_6516,N_3643,N_4332);
nand U6517 (N_6517,N_4830,N_5876);
nor U6518 (N_6518,N_4368,N_4044);
xor U6519 (N_6519,N_5349,N_3138);
and U6520 (N_6520,N_5492,N_3546);
nor U6521 (N_6521,N_5624,N_4540);
or U6522 (N_6522,N_5156,N_3007);
nor U6523 (N_6523,N_5710,N_3206);
nand U6524 (N_6524,N_5879,N_3910);
nor U6525 (N_6525,N_5824,N_5744);
nor U6526 (N_6526,N_5148,N_3448);
nand U6527 (N_6527,N_3293,N_5810);
nand U6528 (N_6528,N_4101,N_4327);
nand U6529 (N_6529,N_4268,N_4024);
nand U6530 (N_6530,N_5291,N_5502);
and U6531 (N_6531,N_5444,N_3325);
nand U6532 (N_6532,N_3782,N_5125);
nand U6533 (N_6533,N_5859,N_5213);
and U6534 (N_6534,N_3320,N_3029);
or U6535 (N_6535,N_4605,N_3015);
and U6536 (N_6536,N_4642,N_4151);
and U6537 (N_6537,N_5045,N_5256);
and U6538 (N_6538,N_3661,N_3873);
and U6539 (N_6539,N_4953,N_4757);
and U6540 (N_6540,N_3740,N_3246);
nand U6541 (N_6541,N_3258,N_3812);
nor U6542 (N_6542,N_4511,N_5945);
xnor U6543 (N_6543,N_3644,N_4093);
nor U6544 (N_6544,N_5595,N_4488);
and U6545 (N_6545,N_5165,N_3276);
nor U6546 (N_6546,N_3009,N_3467);
nand U6547 (N_6547,N_5565,N_3183);
nor U6548 (N_6548,N_4120,N_3613);
nor U6549 (N_6549,N_4202,N_5960);
or U6550 (N_6550,N_5538,N_4341);
xor U6551 (N_6551,N_5494,N_5217);
or U6552 (N_6552,N_4625,N_5575);
xnor U6553 (N_6553,N_5621,N_5281);
and U6554 (N_6554,N_5578,N_4106);
nor U6555 (N_6555,N_3100,N_5060);
xor U6556 (N_6556,N_4808,N_3372);
xor U6557 (N_6557,N_4879,N_5968);
nand U6558 (N_6558,N_5829,N_3188);
or U6559 (N_6559,N_5445,N_3186);
xor U6560 (N_6560,N_4493,N_3879);
xor U6561 (N_6561,N_5150,N_3802);
or U6562 (N_6562,N_3288,N_4597);
or U6563 (N_6563,N_5543,N_4104);
nand U6564 (N_6564,N_4382,N_5333);
and U6565 (N_6565,N_4781,N_5195);
or U6566 (N_6566,N_4964,N_5210);
and U6567 (N_6567,N_5919,N_4160);
and U6568 (N_6568,N_4627,N_3726);
nand U6569 (N_6569,N_4812,N_5806);
or U6570 (N_6570,N_3882,N_4494);
nor U6571 (N_6571,N_5381,N_3519);
nand U6572 (N_6572,N_4492,N_4976);
and U6573 (N_6573,N_5734,N_4960);
nand U6574 (N_6574,N_4648,N_5466);
and U6575 (N_6575,N_4123,N_3924);
nand U6576 (N_6576,N_4248,N_5062);
and U6577 (N_6577,N_5755,N_3332);
and U6578 (N_6578,N_5157,N_4974);
nand U6579 (N_6579,N_5675,N_4585);
xor U6580 (N_6580,N_5090,N_5191);
and U6581 (N_6581,N_3470,N_3198);
and U6582 (N_6582,N_4502,N_5552);
nand U6583 (N_6583,N_4231,N_3663);
or U6584 (N_6584,N_4852,N_4925);
nand U6585 (N_6585,N_5336,N_4600);
nand U6586 (N_6586,N_5529,N_3506);
nand U6587 (N_6587,N_5726,N_3578);
xor U6588 (N_6588,N_3496,N_3381);
nor U6589 (N_6589,N_4509,N_3773);
or U6590 (N_6590,N_5373,N_4304);
nor U6591 (N_6591,N_4533,N_5979);
nand U6592 (N_6592,N_3694,N_4912);
nor U6593 (N_6593,N_4769,N_3000);
nor U6594 (N_6594,N_3179,N_5370);
and U6595 (N_6595,N_4426,N_4414);
or U6596 (N_6596,N_4851,N_5267);
xor U6597 (N_6597,N_3103,N_5463);
nor U6598 (N_6598,N_5588,N_5971);
or U6599 (N_6599,N_3652,N_4014);
and U6600 (N_6600,N_3354,N_5344);
and U6601 (N_6601,N_4219,N_5598);
nand U6602 (N_6602,N_4448,N_4049);
or U6603 (N_6603,N_4432,N_5007);
and U6604 (N_6604,N_3278,N_3593);
and U6605 (N_6605,N_4535,N_5601);
nor U6606 (N_6606,N_3262,N_4541);
and U6607 (N_6607,N_4714,N_5446);
or U6608 (N_6608,N_5517,N_4837);
nand U6609 (N_6609,N_4373,N_3890);
nand U6610 (N_6610,N_5984,N_4359);
or U6611 (N_6611,N_3523,N_4764);
or U6612 (N_6612,N_4343,N_5783);
and U6613 (N_6613,N_5390,N_3832);
nor U6614 (N_6614,N_5069,N_5568);
or U6615 (N_6615,N_4070,N_5242);
nand U6616 (N_6616,N_5139,N_3998);
nor U6617 (N_6617,N_3499,N_4022);
nand U6618 (N_6618,N_3631,N_5314);
or U6619 (N_6619,N_3912,N_5704);
nor U6620 (N_6620,N_3639,N_5769);
and U6621 (N_6621,N_5355,N_4137);
nand U6622 (N_6622,N_4880,N_3026);
nand U6623 (N_6623,N_3645,N_3330);
nand U6624 (N_6624,N_5427,N_3468);
xnor U6625 (N_6625,N_3494,N_4086);
and U6626 (N_6626,N_4402,N_3152);
and U6627 (N_6627,N_4660,N_3302);
nor U6628 (N_6628,N_4929,N_4318);
or U6629 (N_6629,N_4574,N_5910);
and U6630 (N_6630,N_3310,N_3215);
nand U6631 (N_6631,N_3707,N_5049);
nand U6632 (N_6632,N_3943,N_3228);
nor U6633 (N_6633,N_4124,N_4381);
and U6634 (N_6634,N_4263,N_5207);
and U6635 (N_6635,N_3455,N_4337);
or U6636 (N_6636,N_4756,N_5845);
nor U6637 (N_6637,N_4046,N_4169);
nand U6638 (N_6638,N_5693,N_3889);
xnor U6639 (N_6639,N_5187,N_4478);
nor U6640 (N_6640,N_4583,N_5149);
xnor U6641 (N_6641,N_5837,N_4261);
nand U6642 (N_6642,N_4477,N_5424);
nor U6643 (N_6643,N_4317,N_3292);
and U6644 (N_6644,N_5059,N_5286);
nand U6645 (N_6645,N_3781,N_4945);
or U6646 (N_6646,N_5792,N_4233);
nand U6647 (N_6647,N_3954,N_5722);
xnor U6648 (N_6648,N_3376,N_5993);
or U6649 (N_6649,N_4490,N_3219);
xnor U6650 (N_6650,N_3361,N_3602);
nor U6651 (N_6651,N_3672,N_5915);
nor U6652 (N_6652,N_4646,N_3127);
nand U6653 (N_6653,N_3984,N_3001);
xnor U6654 (N_6654,N_4071,N_5374);
nand U6655 (N_6655,N_5530,N_3551);
or U6656 (N_6656,N_5639,N_3891);
nand U6657 (N_6657,N_5569,N_3654);
nand U6658 (N_6658,N_5605,N_4528);
nor U6659 (N_6659,N_3458,N_5176);
or U6660 (N_6660,N_3527,N_4012);
and U6661 (N_6661,N_5745,N_5535);
nand U6662 (N_6662,N_4984,N_4371);
or U6663 (N_6663,N_4796,N_5481);
and U6664 (N_6664,N_4129,N_4687);
or U6665 (N_6665,N_4229,N_5039);
nor U6666 (N_6666,N_3768,N_3112);
nand U6667 (N_6667,N_3862,N_3870);
or U6668 (N_6668,N_4780,N_3553);
nor U6669 (N_6669,N_5991,N_4594);
or U6670 (N_6670,N_3371,N_5353);
nand U6671 (N_6671,N_3444,N_3002);
or U6672 (N_6672,N_3732,N_5640);
or U6673 (N_6673,N_5707,N_4353);
nand U6674 (N_6674,N_3059,N_3239);
xor U6675 (N_6675,N_4326,N_4447);
and U6676 (N_6676,N_3844,N_5393);
or U6677 (N_6677,N_4467,N_5732);
or U6678 (N_6678,N_4328,N_3633);
nor U6679 (N_6679,N_4610,N_4109);
nor U6680 (N_6680,N_3064,N_5999);
or U6681 (N_6681,N_4148,N_4267);
and U6682 (N_6682,N_5527,N_5452);
nor U6683 (N_6683,N_5778,N_4122);
nand U6684 (N_6684,N_3712,N_4982);
nand U6685 (N_6685,N_3264,N_5580);
nand U6686 (N_6686,N_4190,N_3331);
and U6687 (N_6687,N_4979,N_3704);
nand U6688 (N_6688,N_4554,N_4750);
xnor U6689 (N_6689,N_5626,N_4581);
or U6690 (N_6690,N_4608,N_3403);
nand U6691 (N_6691,N_4673,N_3486);
nor U6692 (N_6692,N_3928,N_4064);
nor U6693 (N_6693,N_4735,N_5866);
nand U6694 (N_6694,N_5947,N_4456);
nand U6695 (N_6695,N_4659,N_5951);
and U6696 (N_6696,N_4972,N_4286);
nand U6697 (N_6697,N_3840,N_5064);
nor U6698 (N_6698,N_4864,N_5586);
or U6699 (N_6699,N_5495,N_5936);
or U6700 (N_6700,N_3684,N_4489);
nor U6701 (N_6701,N_4776,N_5518);
xnor U6702 (N_6702,N_4728,N_4312);
nor U6703 (N_6703,N_3934,N_3083);
xnor U6704 (N_6704,N_3260,N_4523);
or U6705 (N_6705,N_4813,N_3846);
nand U6706 (N_6706,N_3173,N_5867);
nand U6707 (N_6707,N_4882,N_3255);
nand U6708 (N_6708,N_5587,N_5937);
or U6709 (N_6709,N_5820,N_4378);
nand U6710 (N_6710,N_3197,N_5666);
and U6711 (N_6711,N_4730,N_3056);
or U6712 (N_6712,N_3556,N_4421);
or U6713 (N_6713,N_5623,N_4411);
nor U6714 (N_6714,N_5290,N_4915);
or U6715 (N_6715,N_5317,N_5399);
and U6716 (N_6716,N_5482,N_5340);
and U6717 (N_6717,N_3549,N_3714);
nor U6718 (N_6718,N_4774,N_4475);
or U6719 (N_6719,N_3480,N_5366);
nand U6720 (N_6720,N_3939,N_4165);
or U6721 (N_6721,N_4719,N_5144);
nor U6722 (N_6722,N_4356,N_4978);
or U6723 (N_6723,N_5685,N_4845);
nand U6724 (N_6724,N_3737,N_5854);
nor U6725 (N_6725,N_3088,N_4985);
nor U6726 (N_6726,N_5881,N_3095);
xnor U6727 (N_6727,N_5980,N_4144);
nor U6728 (N_6728,N_4794,N_3835);
xor U6729 (N_6729,N_3550,N_4762);
and U6730 (N_6730,N_4635,N_5660);
nor U6731 (N_6731,N_4018,N_3505);
and U6732 (N_6732,N_4126,N_3604);
nand U6733 (N_6733,N_4434,N_4291);
nor U6734 (N_6734,N_5283,N_3058);
and U6735 (N_6735,N_5077,N_4208);
nand U6736 (N_6736,N_3797,N_3688);
or U6737 (N_6737,N_5738,N_5437);
and U6738 (N_6738,N_3988,N_5476);
nor U6739 (N_6739,N_4346,N_5567);
nor U6740 (N_6740,N_3404,N_3947);
and U6741 (N_6741,N_4135,N_5022);
or U6742 (N_6742,N_5078,N_4653);
nand U6743 (N_6743,N_5500,N_4622);
and U6744 (N_6744,N_5430,N_5224);
nand U6745 (N_6745,N_5714,N_5431);
nor U6746 (N_6746,N_5521,N_4444);
or U6747 (N_6747,N_4652,N_4543);
xor U6748 (N_6748,N_4185,N_5940);
and U6749 (N_6749,N_5472,N_4549);
or U6750 (N_6750,N_5402,N_3753);
or U6751 (N_6751,N_5723,N_5167);
nand U6752 (N_6752,N_3630,N_3944);
xnor U6753 (N_6753,N_4741,N_5388);
nand U6754 (N_6754,N_4257,N_4639);
and U6755 (N_6755,N_3670,N_4833);
or U6756 (N_6756,N_4006,N_3322);
or U6757 (N_6757,N_5042,N_3166);
nand U6758 (N_6758,N_3192,N_3508);
xor U6759 (N_6759,N_3450,N_3995);
or U6760 (N_6760,N_3554,N_5644);
or U6761 (N_6761,N_4245,N_5698);
nand U6762 (N_6762,N_3780,N_3472);
nor U6763 (N_6763,N_5330,N_5831);
nor U6764 (N_6764,N_3495,N_4300);
or U6765 (N_6765,N_4789,N_4161);
nand U6766 (N_6766,N_3760,N_5276);
and U6767 (N_6767,N_3109,N_4038);
or U6768 (N_6768,N_3417,N_3175);
xor U6769 (N_6769,N_4146,N_4846);
xnor U6770 (N_6770,N_5360,N_3086);
nor U6771 (N_6771,N_3583,N_3039);
and U6772 (N_6772,N_4173,N_4195);
nand U6773 (N_6773,N_5888,N_4335);
or U6774 (N_6774,N_3816,N_5841);
and U6775 (N_6775,N_4399,N_3136);
xnor U6776 (N_6776,N_4739,N_3747);
and U6777 (N_6777,N_4074,N_4894);
and U6778 (N_6778,N_3045,N_4150);
or U6779 (N_6779,N_5287,N_3678);
xor U6780 (N_6780,N_4329,N_4172);
nor U6781 (N_6781,N_5599,N_4072);
xnor U6782 (N_6782,N_4365,N_4542);
and U6783 (N_6783,N_5428,N_5997);
or U6784 (N_6784,N_4821,N_5890);
nand U6785 (N_6785,N_3923,N_4508);
nor U6786 (N_6786,N_4968,N_5308);
nand U6787 (N_6787,N_5513,N_5318);
nor U6788 (N_6788,N_4363,N_3800);
and U6789 (N_6789,N_3364,N_3275);
nor U6790 (N_6790,N_3561,N_5773);
or U6791 (N_6791,N_4962,N_5498);
and U6792 (N_6792,N_5216,N_4724);
and U6793 (N_6793,N_4457,N_4557);
or U6794 (N_6794,N_5272,N_3397);
or U6795 (N_6795,N_5801,N_5724);
or U6796 (N_6796,N_4547,N_4283);
nor U6797 (N_6797,N_4431,N_5124);
xnor U6798 (N_6798,N_4408,N_5197);
and U6799 (N_6799,N_3902,N_5763);
and U6800 (N_6800,N_5211,N_4763);
and U6801 (N_6801,N_3067,N_3597);
or U6802 (N_6802,N_5032,N_4118);
and U6803 (N_6803,N_3560,N_3414);
xor U6804 (N_6804,N_5041,N_3465);
nand U6805 (N_6805,N_4051,N_3076);
nand U6806 (N_6806,N_5572,N_4117);
or U6807 (N_6807,N_3823,N_3863);
xnor U6808 (N_6808,N_4892,N_3023);
nor U6809 (N_6809,N_3191,N_5798);
xor U6810 (N_6810,N_3843,N_5134);
xor U6811 (N_6811,N_4386,N_5038);
and U6812 (N_6812,N_4778,N_3820);
and U6813 (N_6813,N_5408,N_3185);
and U6814 (N_6814,N_3705,N_4695);
and U6815 (N_6815,N_4904,N_4319);
nand U6816 (N_6816,N_3530,N_4143);
and U6817 (N_6817,N_5990,N_5259);
and U6818 (N_6818,N_3196,N_5037);
nand U6819 (N_6819,N_4013,N_4189);
nand U6820 (N_6820,N_4819,N_3261);
nand U6821 (N_6821,N_5969,N_4096);
nand U6822 (N_6822,N_3340,N_5786);
xnor U6823 (N_6823,N_3040,N_4618);
nand U6824 (N_6824,N_4254,N_5307);
or U6825 (N_6825,N_3701,N_4693);
and U6826 (N_6826,N_3463,N_3881);
nor U6827 (N_6827,N_5312,N_3897);
and U6828 (N_6828,N_3792,N_3117);
and U6829 (N_6829,N_4722,N_3813);
nor U6830 (N_6830,N_4439,N_5293);
and U6831 (N_6831,N_3409,N_5503);
and U6832 (N_6832,N_4518,N_5411);
or U6833 (N_6833,N_5324,N_3769);
nand U6834 (N_6834,N_3336,N_4788);
or U6835 (N_6835,N_3829,N_5164);
and U6836 (N_6836,N_4664,N_3731);
or U6837 (N_6837,N_4878,N_4504);
nor U6838 (N_6838,N_5956,N_5320);
nand U6839 (N_6839,N_3199,N_5277);
nand U6840 (N_6840,N_3711,N_4793);
nor U6841 (N_6841,N_4499,N_4992);
and U6842 (N_6842,N_4951,N_4795);
nor U6843 (N_6843,N_5804,N_5855);
and U6844 (N_6844,N_4975,N_4628);
nor U6845 (N_6845,N_3566,N_3481);
or U6846 (N_6846,N_5470,N_5089);
or U6847 (N_6847,N_4593,N_5289);
xnor U6848 (N_6848,N_3819,N_5058);
or U6849 (N_6849,N_5161,N_5571);
and U6850 (N_6850,N_3857,N_4571);
and U6851 (N_6851,N_4374,N_4617);
or U6852 (N_6852,N_5709,N_3791);
nor U6853 (N_6853,N_5202,N_4703);
nand U6854 (N_6854,N_5083,N_5475);
nor U6855 (N_6855,N_5454,N_4903);
nor U6856 (N_6856,N_5442,N_4196);
nor U6857 (N_6857,N_5334,N_3245);
and U6858 (N_6858,N_3955,N_3847);
nand U6859 (N_6859,N_3949,N_5681);
nand U6860 (N_6860,N_4110,N_3808);
xnor U6861 (N_6861,N_5448,N_5196);
nor U6862 (N_6862,N_4171,N_5024);
nand U6863 (N_6863,N_3116,N_3736);
nand U6864 (N_6864,N_3552,N_5874);
xor U6865 (N_6865,N_5418,N_3518);
or U6866 (N_6866,N_4262,N_5895);
or U6867 (N_6867,N_4181,N_5609);
nand U6868 (N_6868,N_4484,N_3842);
and U6869 (N_6869,N_4767,N_3529);
xor U6870 (N_6870,N_5795,N_3043);
and U6871 (N_6871,N_4232,N_5924);
or U6872 (N_6872,N_4021,N_3378);
nor U6873 (N_6873,N_5199,N_5115);
xnor U6874 (N_6874,N_3344,N_5178);
nand U6875 (N_6875,N_5395,N_4561);
xnor U6876 (N_6876,N_4939,N_3541);
or U6877 (N_6877,N_4883,N_4153);
nor U6878 (N_6878,N_3572,N_5208);
nor U6879 (N_6879,N_3770,N_4105);
nand U6880 (N_6880,N_3211,N_3801);
xnor U6881 (N_6881,N_4961,N_4166);
xnor U6882 (N_6882,N_5689,N_3778);
or U6883 (N_6883,N_5063,N_5304);
nand U6884 (N_6884,N_5828,N_3144);
or U6885 (N_6885,N_4338,N_4538);
nor U6886 (N_6886,N_3950,N_3522);
xor U6887 (N_6887,N_4957,N_5383);
xor U6888 (N_6888,N_5085,N_4077);
or U6889 (N_6889,N_5622,N_4706);
or U6890 (N_6890,N_4681,N_5742);
or U6891 (N_6891,N_3042,N_4944);
or U6892 (N_6892,N_5152,N_4970);
nor U6893 (N_6893,N_4934,N_4956);
and U6894 (N_6894,N_3834,N_3285);
and U6895 (N_6895,N_4188,N_3283);
or U6896 (N_6896,N_5735,N_3439);
nor U6897 (N_6897,N_3676,N_4921);
xnor U6898 (N_6898,N_3011,N_3592);
and U6899 (N_6899,N_4844,N_5894);
and U6900 (N_6900,N_3339,N_5499);
nand U6901 (N_6901,N_4853,N_3046);
and U6902 (N_6902,N_4534,N_5731);
nor U6903 (N_6903,N_4754,N_3544);
nor U6904 (N_6904,N_3648,N_4658);
nand U6905 (N_6905,N_4265,N_5564);
or U6906 (N_6906,N_3263,N_3545);
nor U6907 (N_6907,N_3395,N_3926);
nor U6908 (N_6908,N_4887,N_5053);
or U6909 (N_6909,N_5677,N_3664);
nand U6910 (N_6910,N_5589,N_3850);
nand U6911 (N_6911,N_4454,N_4784);
or U6912 (N_6912,N_5759,N_3741);
nand U6913 (N_6913,N_4026,N_5903);
xor U6914 (N_6914,N_5983,N_4252);
nand U6915 (N_6915,N_3174,N_3355);
nand U6916 (N_6916,N_4531,N_4375);
or U6917 (N_6917,N_5655,N_3681);
or U6918 (N_6918,N_5953,N_3236);
or U6919 (N_6919,N_3777,N_3500);
and U6920 (N_6920,N_3730,N_4147);
and U6921 (N_6921,N_5717,N_4442);
nand U6922 (N_6922,N_5485,N_3240);
nor U6923 (N_6923,N_4626,N_4725);
xnor U6924 (N_6924,N_4155,N_5729);
and U6925 (N_6925,N_3717,N_5522);
or U6926 (N_6926,N_5155,N_5129);
nor U6927 (N_6927,N_4591,N_5342);
nand U6928 (N_6928,N_5253,N_3289);
xnor U6929 (N_6929,N_3177,N_5602);
xor U6930 (N_6930,N_5948,N_3051);
nor U6931 (N_6931,N_5017,N_4707);
and U6932 (N_6932,N_3140,N_4530);
and U6933 (N_6933,N_4430,N_5222);
and U6934 (N_6934,N_3675,N_4902);
or U6935 (N_6935,N_5830,N_5056);
and U6936 (N_6936,N_3169,N_5363);
nor U6937 (N_6937,N_3123,N_4002);
nor U6938 (N_6938,N_5415,N_3351);
nor U6939 (N_6939,N_4294,N_3267);
nor U6940 (N_6940,N_4544,N_4917);
xor U6941 (N_6941,N_3722,N_3158);
and U6942 (N_6942,N_4384,N_4691);
xnor U6943 (N_6943,N_3636,N_3368);
nor U6944 (N_6944,N_4367,N_5179);
and U6945 (N_6945,N_5040,N_3685);
nor U6946 (N_6946,N_4008,N_4694);
xor U6947 (N_6947,N_4198,N_5082);
and U6948 (N_6948,N_3608,N_5840);
or U6949 (N_6949,N_3205,N_3172);
and U6950 (N_6950,N_4711,N_4555);
or U6951 (N_6951,N_4139,N_4498);
or U6952 (N_6952,N_4775,N_3526);
and U6953 (N_6953,N_4933,N_3724);
nor U6954 (N_6954,N_4005,N_5524);
and U6955 (N_6955,N_3412,N_5928);
nand U6956 (N_6956,N_5265,N_5455);
xnor U6957 (N_6957,N_3858,N_4710);
and U6958 (N_6958,N_3667,N_3565);
nor U6959 (N_6959,N_5583,N_3691);
nor U6960 (N_6960,N_5128,N_5116);
and U6961 (N_6961,N_3877,N_3006);
nand U6962 (N_6962,N_5817,N_3209);
nor U6963 (N_6963,N_3249,N_5532);
nor U6964 (N_6964,N_5985,N_5313);
nand U6965 (N_6965,N_3077,N_5464);
nor U6966 (N_6966,N_4339,N_5912);
and U6967 (N_6967,N_3703,N_4348);
or U6968 (N_6968,N_3932,N_4418);
or U6969 (N_6969,N_3543,N_5412);
nor U6970 (N_6970,N_3385,N_5651);
or U6971 (N_6971,N_3248,N_4401);
and U6972 (N_6972,N_3946,N_3365);
or U6973 (N_6973,N_3838,N_5376);
nor U6974 (N_6974,N_5215,N_4287);
nor U6975 (N_6975,N_5970,N_4747);
nor U6976 (N_6976,N_3940,N_5938);
nor U6977 (N_6977,N_5047,N_4685);
nand U6978 (N_6978,N_5590,N_3294);
or U6979 (N_6979,N_4548,N_3788);
and U6980 (N_6980,N_3824,N_5629);
nor U6981 (N_6981,N_3689,N_5563);
nand U6982 (N_6982,N_4031,N_5627);
xor U6983 (N_6983,N_5901,N_5597);
or U6984 (N_6984,N_3413,N_3018);
and U6985 (N_6985,N_5652,N_3222);
or U6986 (N_6986,N_4108,N_3517);
nand U6987 (N_6987,N_3269,N_3682);
or U6988 (N_6988,N_3606,N_3647);
and U6989 (N_6989,N_3513,N_4119);
or U6990 (N_6990,N_4419,N_4249);
or U6991 (N_6991,N_3315,N_3807);
and U6992 (N_6992,N_3570,N_4174);
nor U6993 (N_6993,N_3765,N_3034);
nor U6994 (N_6994,N_5963,N_5158);
or U6995 (N_6995,N_4073,N_5326);
or U6996 (N_6996,N_3235,N_5274);
or U6997 (N_6997,N_3564,N_3723);
xor U6998 (N_6998,N_5212,N_3483);
nand U6999 (N_6999,N_3851,N_4667);
nand U7000 (N_7000,N_4704,N_4440);
or U7001 (N_7001,N_5719,N_5663);
or U7002 (N_7002,N_4517,N_5746);
and U7003 (N_7003,N_3122,N_3418);
nand U7004 (N_7004,N_3536,N_4420);
xnor U7005 (N_7005,N_5086,N_4463);
or U7006 (N_7006,N_4054,N_5346);
or U7007 (N_7007,N_5239,N_3305);
nand U7008 (N_7008,N_5181,N_3398);
or U7009 (N_7009,N_4748,N_5750);
or U7010 (N_7010,N_3607,N_5862);
nand U7011 (N_7011,N_4568,N_3380);
nand U7012 (N_7012,N_4810,N_5743);
or U7013 (N_7013,N_4361,N_5932);
nand U7014 (N_7014,N_4053,N_4011);
xnor U7015 (N_7015,N_5433,N_4512);
nor U7016 (N_7016,N_3342,N_3528);
and U7017 (N_7017,N_5691,N_4870);
xnor U7018 (N_7018,N_3053,N_4866);
nor U7019 (N_7019,N_3120,N_3004);
nor U7020 (N_7020,N_5628,N_5591);
and U7021 (N_7021,N_3914,N_5542);
and U7022 (N_7022,N_3366,N_5682);
and U7023 (N_7023,N_5405,N_3715);
and U7024 (N_7024,N_5760,N_4807);
and U7025 (N_7025,N_3280,N_4873);
and U7026 (N_7026,N_5899,N_3745);
nand U7027 (N_7027,N_5416,N_3830);
nor U7028 (N_7028,N_4993,N_5070);
nor U7029 (N_7029,N_5716,N_3462);
nand U7030 (N_7030,N_5084,N_5827);
nand U7031 (N_7031,N_5392,N_5643);
and U7032 (N_7032,N_5218,N_3038);
or U7033 (N_7033,N_5701,N_3318);
nor U7034 (N_7034,N_4425,N_4900);
and U7035 (N_7035,N_4303,N_5447);
or U7036 (N_7036,N_5809,N_4657);
nor U7037 (N_7037,N_5075,N_5251);
and U7038 (N_7038,N_4860,N_5776);
and U7039 (N_7039,N_3762,N_4650);
xnor U7040 (N_7040,N_5813,N_4746);
nand U7041 (N_7041,N_5770,N_4716);
or U7042 (N_7042,N_5725,N_4755);
nand U7043 (N_7043,N_5511,N_5821);
nand U7044 (N_7044,N_4595,N_5184);
or U7045 (N_7045,N_5848,N_4206);
nor U7046 (N_7046,N_3265,N_3035);
nand U7047 (N_7047,N_3016,N_4946);
nor U7048 (N_7048,N_4487,N_4397);
nand U7049 (N_7049,N_5548,N_3221);
nand U7050 (N_7050,N_5391,N_3146);
and U7051 (N_7051,N_5295,N_5389);
nand U7052 (N_7052,N_3512,N_5962);
nor U7053 (N_7053,N_4130,N_3454);
and U7054 (N_7054,N_4269,N_5612);
nor U7055 (N_7055,N_4613,N_5642);
or U7056 (N_7056,N_4841,N_5678);
nor U7057 (N_7057,N_4596,N_4809);
or U7058 (N_7058,N_5610,N_4768);
nor U7059 (N_7059,N_5523,N_3833);
nand U7060 (N_7060,N_4314,N_3110);
nand U7061 (N_7061,N_4510,N_5477);
nand U7062 (N_7062,N_3250,N_5604);
and U7063 (N_7063,N_3352,N_3577);
or U7064 (N_7064,N_4023,N_4214);
nand U7065 (N_7065,N_3431,N_3886);
and U7066 (N_7066,N_3257,N_4940);
or U7067 (N_7067,N_5488,N_3903);
nand U7068 (N_7068,N_4176,N_5687);
nor U7069 (N_7069,N_3312,N_4016);
and U7070 (N_7070,N_3072,N_4091);
nor U7071 (N_7071,N_4403,N_4858);
nor U7072 (N_7072,N_5021,N_4566);
and U7073 (N_7073,N_5419,N_3111);
or U7074 (N_7074,N_3200,N_4616);
xor U7075 (N_7075,N_5205,N_4811);
nor U7076 (N_7076,N_4465,N_3287);
nor U7077 (N_7077,N_5294,N_5147);
nor U7078 (N_7078,N_3303,N_3913);
nor U7079 (N_7079,N_3396,N_5617);
nor U7080 (N_7080,N_5943,N_4132);
and U7081 (N_7081,N_3237,N_3382);
xnor U7082 (N_7082,N_3102,N_5114);
nor U7083 (N_7083,N_5952,N_4164);
and U7084 (N_7084,N_3027,N_5555);
nor U7085 (N_7085,N_5118,N_4923);
nor U7086 (N_7086,N_3375,N_3978);
nand U7087 (N_7087,N_5566,N_3036);
nand U7088 (N_7088,N_4228,N_4832);
nor U7089 (N_7089,N_4615,N_5727);
or U7090 (N_7090,N_4529,N_4705);
nand U7091 (N_7091,N_5051,N_4223);
or U7092 (N_7092,N_4898,N_4553);
nor U7093 (N_7093,N_4226,N_4025);
nor U7094 (N_7094,N_4671,N_3999);
nor U7095 (N_7095,N_5796,N_4802);
or U7096 (N_7096,N_5140,N_5733);
or U7097 (N_7097,N_5141,N_5672);
nand U7098 (N_7098,N_5554,N_4009);
and U7099 (N_7099,N_4803,N_3692);
nand U7100 (N_7100,N_4100,N_5079);
and U7101 (N_7101,N_5844,N_5400);
nor U7102 (N_7102,N_5671,N_3476);
or U7103 (N_7103,N_5028,N_4205);
nor U7104 (N_7104,N_3220,N_4877);
or U7105 (N_7105,N_4302,N_4928);
and U7106 (N_7106,N_3900,N_4057);
and U7107 (N_7107,N_5975,N_5560);
nand U7108 (N_7108,N_4570,N_3771);
nand U7109 (N_7109,N_5130,N_5237);
nand U7110 (N_7110,N_3979,N_3673);
or U7111 (N_7111,N_3363,N_5403);
nand U7112 (N_7112,N_5120,N_5846);
and U7113 (N_7113,N_3989,N_4240);
and U7114 (N_7114,N_4436,N_4020);
nand U7115 (N_7115,N_4745,N_3776);
nand U7116 (N_7116,N_3790,N_4831);
nand U7117 (N_7117,N_3972,N_4230);
xnor U7118 (N_7118,N_5483,N_4296);
and U7119 (N_7119,N_5561,N_4881);
or U7120 (N_7120,N_4815,N_5545);
nand U7121 (N_7121,N_5531,N_5132);
nand U7122 (N_7122,N_3426,N_4310);
nand U7123 (N_7123,N_5104,N_4655);
nor U7124 (N_7124,N_4217,N_5533);
or U7125 (N_7125,N_4692,N_5044);
nand U7126 (N_7126,N_3126,N_5243);
nand U7127 (N_7127,N_5378,N_3337);
and U7128 (N_7128,N_4688,N_4255);
or U7129 (N_7129,N_3764,N_5774);
nor U7130 (N_7130,N_5851,N_3498);
nor U7131 (N_7131,N_4977,N_4592);
nand U7132 (N_7132,N_4085,N_5939);
and U7133 (N_7133,N_3475,N_5973);
or U7134 (N_7134,N_3254,N_3810);
nand U7135 (N_7135,N_3153,N_4679);
or U7136 (N_7136,N_3066,N_4965);
nor U7137 (N_7137,N_4603,N_5669);
and U7138 (N_7138,N_4279,N_3861);
or U7139 (N_7139,N_3938,N_3165);
xnor U7140 (N_7140,N_4672,N_4580);
or U7141 (N_7141,N_3440,N_3909);
nor U7142 (N_7142,N_5728,N_3178);
nor U7143 (N_7143,N_3713,N_3815);
and U7144 (N_7144,N_4050,N_3251);
nor U7145 (N_7145,N_5413,N_3080);
and U7146 (N_7146,N_3266,N_3524);
or U7147 (N_7147,N_3208,N_5490);
xnor U7148 (N_7148,N_4340,N_5093);
and U7149 (N_7149,N_3306,N_4215);
nor U7150 (N_7150,N_4587,N_5352);
and U7151 (N_7151,N_4481,N_4865);
nand U7152 (N_7152,N_3837,N_3139);
xor U7153 (N_7153,N_3980,N_5507);
or U7154 (N_7154,N_5171,N_4247);
nand U7155 (N_7155,N_4028,N_5961);
and U7156 (N_7156,N_5918,N_3202);
and U7157 (N_7157,N_4996,N_5240);
and U7158 (N_7158,N_4702,N_5337);
nor U7159 (N_7159,N_5377,N_3074);
nand U7160 (N_7160,N_4733,N_5768);
nand U7161 (N_7161,N_4611,N_4443);
and U7162 (N_7162,N_3410,N_4313);
xnor U7163 (N_7163,N_5159,N_5238);
or U7164 (N_7164,N_4225,N_4643);
nand U7165 (N_7165,N_4825,N_5269);
or U7166 (N_7166,N_4519,N_4476);
and U7167 (N_7167,N_3057,N_5562);
or U7168 (N_7168,N_4380,N_5254);
nor U7169 (N_7169,N_5046,N_3021);
nand U7170 (N_7170,N_5057,N_5432);
and U7171 (N_7171,N_4785,N_4751);
or U7172 (N_7172,N_5665,N_5749);
and U7173 (N_7173,N_4740,N_4950);
or U7174 (N_7174,N_3299,N_5106);
and U7175 (N_7175,N_5440,N_3906);
nor U7176 (N_7176,N_5375,N_3184);
nand U7177 (N_7177,N_4564,N_3313);
nand U7178 (N_7178,N_5214,N_4577);
or U7179 (N_7179,N_3585,N_3401);
nor U7180 (N_7180,N_4856,N_4911);
nand U7181 (N_7181,N_5869,N_3073);
nand U7182 (N_7182,N_3474,N_5072);
nor U7183 (N_7183,N_4913,N_5994);
nand U7184 (N_7184,N_4469,N_3766);
xnor U7185 (N_7185,N_5995,N_5737);
and U7186 (N_7186,N_3956,N_5762);
and U7187 (N_7187,N_5169,N_5061);
nor U7188 (N_7188,N_5315,N_4717);
xnor U7189 (N_7189,N_3374,N_3478);
xnor U7190 (N_7190,N_5608,N_4990);
xnor U7191 (N_7191,N_4388,N_4721);
nor U7192 (N_7192,N_4158,N_4839);
or U7193 (N_7193,N_4773,N_4734);
and U7194 (N_7194,N_5925,N_4588);
nor U7195 (N_7195,N_4424,N_3887);
and U7196 (N_7196,N_4295,N_4524);
xor U7197 (N_7197,N_4835,N_5989);
and U7198 (N_7198,N_4614,N_5356);
or U7199 (N_7199,N_5368,N_5648);
or U7200 (N_7200,N_3055,N_5927);
nor U7201 (N_7201,N_5011,N_4004);
or U7202 (N_7202,N_5194,N_3044);
nand U7203 (N_7203,N_3384,N_5067);
xor U7204 (N_7204,N_3595,N_3905);
xnor U7205 (N_7205,N_5579,N_4849);
and U7206 (N_7206,N_3756,N_3421);
nor U7207 (N_7207,N_5982,N_5800);
and U7208 (N_7208,N_5230,N_4357);
nor U7209 (N_7209,N_5302,N_3933);
nor U7210 (N_7210,N_4682,N_3445);
or U7211 (N_7211,N_3491,N_4765);
and U7212 (N_7212,N_5480,N_3442);
xor U7213 (N_7213,N_3666,N_3193);
and U7214 (N_7214,N_3969,N_5772);
nand U7215 (N_7215,N_3180,N_3181);
and U7216 (N_7216,N_5838,N_4539);
nand U7217 (N_7217,N_5110,N_5174);
nand U7218 (N_7218,N_5096,N_4358);
or U7219 (N_7219,N_5227,N_4342);
and U7220 (N_7220,N_3758,N_3147);
nor U7221 (N_7221,N_5397,N_5425);
nor U7222 (N_7222,N_5131,N_3515);
or U7223 (N_7223,N_5606,N_4676);
or U7224 (N_7224,N_3931,N_3383);
xnor U7225 (N_7225,N_5758,N_5198);
and U7226 (N_7226,N_3270,N_5133);
nor U7227 (N_7227,N_5006,N_4058);
nand U7228 (N_7228,N_3575,N_3182);
and U7229 (N_7229,N_5696,N_4413);
and U7230 (N_7230,N_3548,N_5616);
nor U7231 (N_7231,N_3538,N_5505);
and U7232 (N_7232,N_3677,N_3751);
nand U7233 (N_7233,N_3547,N_3822);
nand U7234 (N_7234,N_3793,N_5636);
or U7235 (N_7235,N_3099,N_3460);
nand U7236 (N_7236,N_4816,N_4183);
nor U7237 (N_7237,N_3634,N_4090);
and U7238 (N_7238,N_5926,N_3920);
or U7239 (N_7239,N_5255,N_4116);
nor U7240 (N_7240,N_5515,N_4211);
nand U7241 (N_7241,N_5394,N_3516);
or U7242 (N_7242,N_5547,N_4392);
nor U7243 (N_7243,N_5861,N_4665);
nand U7244 (N_7244,N_3599,N_5111);
and U7245 (N_7245,N_4428,N_3856);
nand U7246 (N_7246,N_5559,N_5812);
nor U7247 (N_7247,N_3092,N_5832);
xor U7248 (N_7248,N_5880,N_4861);
and U7249 (N_7249,N_3241,N_4863);
nor U7250 (N_7250,N_5931,N_3821);
nand U7251 (N_7251,N_3273,N_3466);
xnor U7252 (N_7252,N_4840,N_4162);
or U7253 (N_7253,N_3189,N_5282);
or U7254 (N_7254,N_4527,N_4906);
nand U7255 (N_7255,N_3390,N_3977);
nand U7256 (N_7256,N_3612,N_4690);
or U7257 (N_7257,N_4668,N_4567);
or U7258 (N_7258,N_5009,N_5600);
nor U7259 (N_7259,N_4516,N_3348);
nand U7260 (N_7260,N_5887,N_4995);
and U7261 (N_7261,N_4641,N_4496);
and U7262 (N_7262,N_4947,N_4034);
and U7263 (N_7263,N_3757,N_5646);
and U7264 (N_7264,N_3748,N_4683);
nand U7265 (N_7265,N_3915,N_4503);
xnor U7266 (N_7266,N_5929,N_5864);
nand U7267 (N_7267,N_3598,N_4079);
nor U7268 (N_7268,N_3085,N_3615);
or U7269 (N_7269,N_5748,N_5808);
and U7270 (N_7270,N_3744,N_5585);
and U7271 (N_7271,N_3082,N_4306);
nand U7272 (N_7272,N_5573,N_4098);
nor U7273 (N_7273,N_4818,N_5789);
nand U7274 (N_7274,N_4128,N_4708);
xor U7275 (N_7275,N_5544,N_3151);
nand U7276 (N_7276,N_5173,N_4569);
and U7277 (N_7277,N_5708,N_4391);
nor U7278 (N_7278,N_5332,N_5536);
and U7279 (N_7279,N_4817,N_3831);
or U7280 (N_7280,N_5261,N_3779);
nand U7281 (N_7281,N_3105,N_4404);
nor U7282 (N_7282,N_3488,N_3795);
nand U7283 (N_7283,N_4210,N_4575);
and U7284 (N_7284,N_4352,N_3662);
and U7285 (N_7285,N_5456,N_4429);
nor U7286 (N_7286,N_4125,N_5546);
and U7287 (N_7287,N_5491,N_4589);
nand U7288 (N_7288,N_3668,N_4234);
or U7289 (N_7289,N_4369,N_4474);
and U7290 (N_7290,N_5297,N_5025);
nor U7291 (N_7291,N_4396,N_3379);
nor U7292 (N_7292,N_5189,N_5870);
nand U7293 (N_7293,N_5023,N_3884);
nand U7294 (N_7294,N_4030,N_3953);
or U7295 (N_7295,N_5203,N_3168);
nor U7296 (N_7296,N_5136,N_4822);
nor U7297 (N_7297,N_3359,N_5692);
nand U7298 (N_7298,N_4559,N_5767);
and U7299 (N_7299,N_5135,N_5396);
or U7300 (N_7300,N_3571,N_4056);
and U7301 (N_7301,N_4354,N_4370);
and U7302 (N_7302,N_5823,N_4644);
or U7303 (N_7303,N_3537,N_4834);
nand U7304 (N_7304,N_5097,N_5884);
nand U7305 (N_7305,N_5248,N_4237);
nor U7306 (N_7306,N_3709,N_3345);
nor U7307 (N_7307,N_5659,N_5514);
nor U7308 (N_7308,N_3358,N_3019);
or U7309 (N_7309,N_4389,N_3437);
or U7310 (N_7310,N_3901,N_3918);
nand U7311 (N_7311,N_4800,N_3008);
and U7312 (N_7312,N_3507,N_4001);
and U7313 (N_7313,N_3279,N_3075);
and U7314 (N_7314,N_5647,N_4619);
nor U7315 (N_7315,N_5641,N_4076);
or U7316 (N_7316,N_4393,N_3217);
nor U7317 (N_7317,N_4376,N_3853);
or U7318 (N_7318,N_3755,N_5098);
nor U7319 (N_7319,N_5797,N_3616);
or U7320 (N_7320,N_3700,N_3787);
nor U7321 (N_7321,N_4590,N_4909);
or U7322 (N_7322,N_4309,N_5528);
and U7323 (N_7323,N_3699,N_3094);
and U7324 (N_7324,N_4612,N_3433);
and U7325 (N_7325,N_4988,N_5699);
nor U7326 (N_7326,N_3749,N_5226);
nor U7327 (N_7327,N_3356,N_4260);
nor U7328 (N_7328,N_4175,N_5328);
nand U7329 (N_7329,N_5896,N_4445);
or U7330 (N_7330,N_4200,N_5450);
or U7331 (N_7331,N_4901,N_4280);
nand U7332 (N_7332,N_5154,N_3651);
nand U7333 (N_7333,N_5113,N_4036);
nor U7334 (N_7334,N_5512,N_4836);
and U7335 (N_7335,N_3852,N_4888);
nand U7336 (N_7336,N_3244,N_3855);
nor U7337 (N_7337,N_3391,N_4097);
nor U7338 (N_7338,N_3324,N_5285);
or U7339 (N_7339,N_5835,N_3721);
or U7340 (N_7340,N_3370,N_5697);
or U7341 (N_7341,N_4967,N_5384);
and U7342 (N_7342,N_4275,N_4387);
and U7343 (N_7343,N_3690,N_4482);
or U7344 (N_7344,N_3888,N_4491);
nand U7345 (N_7345,N_3997,N_3827);
or U7346 (N_7346,N_3971,N_4435);
nor U7347 (N_7347,N_5453,N_5306);
nor U7348 (N_7348,N_3624,N_5153);
or U7349 (N_7349,N_4422,N_4298);
and U7350 (N_7350,N_4486,N_5551);
or U7351 (N_7351,N_3164,N_5977);
nand U7352 (N_7352,N_5706,N_5756);
nand U7353 (N_7353,N_5632,N_4220);
or U7354 (N_7354,N_5335,N_5459);
and U7355 (N_7355,N_4718,N_5126);
nor U7356 (N_7356,N_3504,N_4827);
nor U7357 (N_7357,N_3161,N_5296);
and U7358 (N_7358,N_3866,N_5771);
and U7359 (N_7359,N_3911,N_4697);
and U7360 (N_7360,N_3226,N_4179);
or U7361 (N_7361,N_4959,N_5323);
or U7362 (N_7362,N_3986,N_4136);
or U7363 (N_7363,N_3869,N_4059);
and U7364 (N_7364,N_3605,N_4330);
nand U7365 (N_7365,N_4862,N_4182);
nor U7366 (N_7366,N_4250,N_3674);
or U7367 (N_7367,N_3137,N_3563);
nand U7368 (N_7368,N_4003,N_3428);
xnor U7369 (N_7369,N_5143,N_5321);
xor U7370 (N_7370,N_3796,N_4256);
nand U7371 (N_7371,N_5467,N_5582);
nor U7372 (N_7372,N_5680,N_5186);
nor U7373 (N_7373,N_4829,N_5863);
nor U7374 (N_7374,N_4406,N_3247);
nand U7375 (N_7375,N_4191,N_5752);
and U7376 (N_7376,N_4905,N_5013);
nand U7377 (N_7377,N_5458,N_3141);
nor U7378 (N_7378,N_3346,N_3996);
nand U7379 (N_7379,N_3772,N_5231);
xor U7380 (N_7380,N_3735,N_5661);
nand U7381 (N_7381,N_3558,N_3727);
xnor U7382 (N_7382,N_5443,N_5316);
nand U7383 (N_7383,N_5435,N_3485);
nor U7384 (N_7384,N_4433,N_4790);
xor U7385 (N_7385,N_3617,N_4661);
and U7386 (N_7386,N_4017,N_5451);
and U7387 (N_7387,N_3574,N_5766);
nand U7388 (N_7388,N_4783,N_4464);
or U7389 (N_7389,N_4019,N_5877);
nor U7390 (N_7390,N_4470,N_4943);
xnor U7391 (N_7391,N_4415,N_5849);
or U7392 (N_7392,N_4647,N_4955);
or U7393 (N_7393,N_4037,N_3783);
or U7394 (N_7394,N_4410,N_5898);
and U7395 (N_7395,N_3049,N_3061);
nor U7396 (N_7396,N_3629,N_3951);
nor U7397 (N_7397,N_3089,N_3539);
xor U7398 (N_7398,N_5807,N_3520);
and U7399 (N_7399,N_4462,N_4699);
nand U7400 (N_7400,N_3438,N_5765);
nor U7401 (N_7401,N_3620,N_4041);
or U7402 (N_7402,N_3484,N_3811);
or U7403 (N_7403,N_3149,N_3623);
and U7404 (N_7404,N_4274,N_4438);
and U7405 (N_7405,N_3392,N_4629);
nand U7406 (N_7406,N_4236,N_3974);
nor U7407 (N_7407,N_4372,N_3836);
and U7408 (N_7408,N_5917,N_5386);
or U7409 (N_7409,N_4180,N_5858);
or U7410 (N_7410,N_5594,N_5592);
nand U7411 (N_7411,N_3921,N_4301);
nor U7412 (N_7412,N_4307,N_4259);
and U7413 (N_7413,N_3632,N_3311);
nor U7414 (N_7414,N_3590,N_3420);
and U7415 (N_7415,N_5188,N_5487);
nor U7416 (N_7416,N_5052,N_4088);
xor U7417 (N_7417,N_4607,N_3970);
or U7418 (N_7418,N_3628,N_5266);
or U7419 (N_7419,N_5358,N_4752);
and U7420 (N_7420,N_3471,N_5581);
or U7421 (N_7421,N_4670,N_3961);
nand U7422 (N_7422,N_3750,N_5348);
or U7423 (N_7423,N_4890,N_3425);
nand U7424 (N_7424,N_4095,N_4806);
and U7425 (N_7425,N_3734,N_3871);
and U7426 (N_7426,N_4937,N_5974);
nand U7427 (N_7427,N_4253,N_4777);
and U7428 (N_7428,N_4316,N_3533);
and U7429 (N_7429,N_4199,N_4277);
xnor U7430 (N_7430,N_4092,N_3423);
nor U7431 (N_7431,N_3878,N_3610);
and U7432 (N_7432,N_5649,N_4731);
and U7433 (N_7433,N_3176,N_3081);
nand U7434 (N_7434,N_4216,N_3896);
xnor U7435 (N_7435,N_3848,N_3435);
and U7436 (N_7436,N_4453,N_3569);
nand U7437 (N_7437,N_5401,N_5520);
nand U7438 (N_7438,N_3386,N_3334);
nor U7439 (N_7439,N_5102,N_4989);
or U7440 (N_7440,N_4941,N_3941);
or U7441 (N_7441,N_4680,N_4689);
nand U7442 (N_7442,N_4602,N_5099);
nor U7443 (N_7443,N_3121,N_5736);
nand U7444 (N_7444,N_4398,N_3880);
or U7445 (N_7445,N_5889,N_5688);
nor U7446 (N_7446,N_3341,N_5705);
and U7447 (N_7447,N_5816,N_5782);
and U7448 (N_7448,N_3752,N_3434);
nor U7449 (N_7449,N_4779,N_3929);
or U7450 (N_7450,N_5914,N_5793);
and U7451 (N_7451,N_4558,N_5087);
xnor U7452 (N_7452,N_4899,N_4032);
nor U7453 (N_7453,N_3079,N_3405);
nor U7454 (N_7454,N_4270,N_5192);
nand U7455 (N_7455,N_3277,N_3469);
and U7456 (N_7456,N_4514,N_4069);
and U7457 (N_7457,N_5501,N_3461);
nand U7458 (N_7458,N_5003,N_4284);
nand U7459 (N_7459,N_4666,N_3532);
nand U7460 (N_7460,N_3603,N_3619);
nor U7461 (N_7461,N_5791,N_5319);
and U7462 (N_7462,N_5634,N_4213);
nor U7463 (N_7463,N_4889,N_3588);
and U7464 (N_7464,N_5509,N_4654);
nor U7465 (N_7465,N_4222,N_4163);
nor U7466 (N_7466,N_3686,N_4651);
nor U7467 (N_7467,N_3114,N_5794);
nand U7468 (N_7468,N_5921,N_5350);
xnor U7469 (N_7469,N_5747,N_3898);
nor U7470 (N_7470,N_4483,N_5071);
or U7471 (N_7471,N_3441,N_4952);
nor U7472 (N_7472,N_5909,N_5619);
nor U7473 (N_7473,N_5916,N_3128);
and U7474 (N_7474,N_5221,N_5001);
or U7475 (N_7475,N_4131,N_5066);
or U7476 (N_7476,N_3093,N_4997);
xnor U7477 (N_7477,N_3449,N_5853);
nand U7478 (N_7478,N_3323,N_4324);
and U7479 (N_7479,N_4847,N_4604);
and U7480 (N_7480,N_5339,N_3555);
nor U7481 (N_7481,N_5654,N_4948);
nor U7482 (N_7482,N_5117,N_3047);
and U7483 (N_7483,N_5201,N_5033);
xnor U7484 (N_7484,N_4043,N_5822);
nor U7485 (N_7485,N_5777,N_3443);
nor U7486 (N_7486,N_4562,N_5031);
nor U7487 (N_7487,N_4409,N_3559);
and U7488 (N_7488,N_3579,N_3091);
nor U7489 (N_7489,N_5847,N_3130);
nand U7490 (N_7490,N_3071,N_5694);
nor U7491 (N_7491,N_3679,N_5185);
nor U7492 (N_7492,N_4609,N_3719);
or U7493 (N_7493,N_5950,N_4545);
nor U7494 (N_7494,N_5327,N_4344);
nor U7495 (N_7495,N_4991,N_5233);
nand U7496 (N_7496,N_5469,N_3981);
nand U7497 (N_7497,N_3243,N_5260);
nor U7498 (N_7498,N_4168,N_5206);
xnor U7499 (N_7499,N_5967,N_4926);
or U7500 (N_7500,N_4234,N_3021);
nand U7501 (N_7501,N_3984,N_3561);
or U7502 (N_7502,N_4586,N_4780);
or U7503 (N_7503,N_4284,N_3584);
or U7504 (N_7504,N_5909,N_5997);
nand U7505 (N_7505,N_3167,N_3058);
or U7506 (N_7506,N_5825,N_3307);
nor U7507 (N_7507,N_5603,N_3173);
or U7508 (N_7508,N_5936,N_5419);
nor U7509 (N_7509,N_4912,N_5008);
nand U7510 (N_7510,N_5482,N_3592);
and U7511 (N_7511,N_4353,N_3583);
and U7512 (N_7512,N_4232,N_4427);
or U7513 (N_7513,N_5295,N_4199);
xnor U7514 (N_7514,N_4081,N_5459);
or U7515 (N_7515,N_3839,N_5158);
xnor U7516 (N_7516,N_4365,N_3545);
or U7517 (N_7517,N_5985,N_3721);
nor U7518 (N_7518,N_3732,N_5981);
and U7519 (N_7519,N_4076,N_5252);
or U7520 (N_7520,N_3249,N_4610);
nand U7521 (N_7521,N_5363,N_5662);
nand U7522 (N_7522,N_3944,N_5271);
nor U7523 (N_7523,N_3183,N_4353);
nand U7524 (N_7524,N_4320,N_4094);
nor U7525 (N_7525,N_3656,N_5268);
or U7526 (N_7526,N_5045,N_3476);
and U7527 (N_7527,N_4212,N_5451);
or U7528 (N_7528,N_5388,N_3827);
and U7529 (N_7529,N_3695,N_5747);
nand U7530 (N_7530,N_5170,N_5835);
nand U7531 (N_7531,N_4539,N_4095);
nor U7532 (N_7532,N_5031,N_4619);
xnor U7533 (N_7533,N_3492,N_3621);
or U7534 (N_7534,N_4310,N_3827);
xor U7535 (N_7535,N_4203,N_4896);
nor U7536 (N_7536,N_5487,N_3162);
nor U7537 (N_7537,N_5460,N_5958);
or U7538 (N_7538,N_4828,N_4513);
or U7539 (N_7539,N_5142,N_4779);
and U7540 (N_7540,N_3385,N_3746);
and U7541 (N_7541,N_4188,N_5447);
and U7542 (N_7542,N_4846,N_3159);
and U7543 (N_7543,N_5342,N_5686);
or U7544 (N_7544,N_5662,N_3316);
xnor U7545 (N_7545,N_5819,N_4341);
nor U7546 (N_7546,N_4851,N_5473);
and U7547 (N_7547,N_5052,N_4602);
nor U7548 (N_7548,N_3641,N_5108);
or U7549 (N_7549,N_5485,N_4516);
nand U7550 (N_7550,N_3499,N_4805);
or U7551 (N_7551,N_4733,N_5554);
xnor U7552 (N_7552,N_4014,N_5401);
or U7553 (N_7553,N_5436,N_4408);
nor U7554 (N_7554,N_4010,N_3916);
nand U7555 (N_7555,N_3066,N_3236);
xor U7556 (N_7556,N_3282,N_3883);
or U7557 (N_7557,N_3524,N_5313);
nor U7558 (N_7558,N_3967,N_5685);
nor U7559 (N_7559,N_4630,N_3386);
nor U7560 (N_7560,N_5688,N_4752);
nor U7561 (N_7561,N_3421,N_4170);
and U7562 (N_7562,N_5177,N_3480);
nor U7563 (N_7563,N_3307,N_4596);
xnor U7564 (N_7564,N_5763,N_5192);
or U7565 (N_7565,N_3992,N_5829);
or U7566 (N_7566,N_4567,N_4632);
nor U7567 (N_7567,N_4109,N_5064);
or U7568 (N_7568,N_4144,N_3216);
and U7569 (N_7569,N_4942,N_4505);
xor U7570 (N_7570,N_3862,N_4738);
nor U7571 (N_7571,N_5599,N_4785);
and U7572 (N_7572,N_3556,N_4143);
xor U7573 (N_7573,N_3117,N_4672);
or U7574 (N_7574,N_3011,N_4022);
and U7575 (N_7575,N_4012,N_5640);
or U7576 (N_7576,N_3824,N_3589);
or U7577 (N_7577,N_4627,N_4676);
and U7578 (N_7578,N_4572,N_5373);
nor U7579 (N_7579,N_5372,N_5439);
and U7580 (N_7580,N_4439,N_3613);
nor U7581 (N_7581,N_5783,N_4270);
nand U7582 (N_7582,N_3291,N_3073);
nor U7583 (N_7583,N_4223,N_3977);
nor U7584 (N_7584,N_4515,N_3283);
nor U7585 (N_7585,N_4770,N_4378);
nand U7586 (N_7586,N_5420,N_3887);
nand U7587 (N_7587,N_5190,N_5091);
nand U7588 (N_7588,N_3402,N_3609);
nand U7589 (N_7589,N_4479,N_5897);
and U7590 (N_7590,N_4618,N_5392);
and U7591 (N_7591,N_5877,N_5828);
xnor U7592 (N_7592,N_4362,N_3932);
nand U7593 (N_7593,N_4930,N_4709);
and U7594 (N_7594,N_3806,N_4597);
or U7595 (N_7595,N_4639,N_4829);
nand U7596 (N_7596,N_3267,N_5362);
or U7597 (N_7597,N_5614,N_4598);
nand U7598 (N_7598,N_4501,N_4515);
nor U7599 (N_7599,N_5738,N_4270);
nand U7600 (N_7600,N_5993,N_5207);
or U7601 (N_7601,N_5066,N_3372);
and U7602 (N_7602,N_5433,N_3536);
nor U7603 (N_7603,N_3853,N_5322);
or U7604 (N_7604,N_5920,N_4801);
nand U7605 (N_7605,N_4485,N_3046);
nand U7606 (N_7606,N_3008,N_3048);
and U7607 (N_7607,N_4631,N_3741);
and U7608 (N_7608,N_3745,N_5564);
nand U7609 (N_7609,N_4518,N_4269);
or U7610 (N_7610,N_3014,N_3605);
or U7611 (N_7611,N_4138,N_4176);
nand U7612 (N_7612,N_3407,N_4173);
nor U7613 (N_7613,N_5333,N_4275);
and U7614 (N_7614,N_5054,N_4421);
nor U7615 (N_7615,N_5960,N_3719);
or U7616 (N_7616,N_3814,N_4204);
or U7617 (N_7617,N_3340,N_3142);
and U7618 (N_7618,N_5021,N_5201);
xor U7619 (N_7619,N_3500,N_5011);
nor U7620 (N_7620,N_3167,N_4609);
or U7621 (N_7621,N_4771,N_4652);
or U7622 (N_7622,N_3314,N_5777);
or U7623 (N_7623,N_5522,N_4369);
nor U7624 (N_7624,N_5088,N_5939);
nor U7625 (N_7625,N_5607,N_4991);
and U7626 (N_7626,N_4970,N_4406);
nor U7627 (N_7627,N_5456,N_3480);
or U7628 (N_7628,N_4166,N_4263);
nor U7629 (N_7629,N_3069,N_3950);
and U7630 (N_7630,N_5795,N_3750);
or U7631 (N_7631,N_3552,N_5222);
nor U7632 (N_7632,N_3172,N_4839);
nand U7633 (N_7633,N_5350,N_3806);
nand U7634 (N_7634,N_4648,N_3100);
or U7635 (N_7635,N_4327,N_5693);
or U7636 (N_7636,N_4561,N_3127);
nand U7637 (N_7637,N_4592,N_5374);
nand U7638 (N_7638,N_5792,N_3001);
and U7639 (N_7639,N_3508,N_4657);
xnor U7640 (N_7640,N_5599,N_3658);
nand U7641 (N_7641,N_3587,N_5288);
or U7642 (N_7642,N_4201,N_3652);
nor U7643 (N_7643,N_3781,N_4617);
nor U7644 (N_7644,N_4813,N_3313);
or U7645 (N_7645,N_5752,N_4838);
and U7646 (N_7646,N_3942,N_4779);
or U7647 (N_7647,N_5117,N_4737);
nand U7648 (N_7648,N_5164,N_3505);
nor U7649 (N_7649,N_5059,N_4367);
nor U7650 (N_7650,N_5544,N_5489);
or U7651 (N_7651,N_3012,N_4677);
nand U7652 (N_7652,N_4460,N_5456);
and U7653 (N_7653,N_4405,N_3595);
nor U7654 (N_7654,N_3748,N_4061);
nand U7655 (N_7655,N_5170,N_5961);
nand U7656 (N_7656,N_4472,N_5305);
nor U7657 (N_7657,N_3544,N_3411);
or U7658 (N_7658,N_3732,N_5801);
or U7659 (N_7659,N_3640,N_3986);
xnor U7660 (N_7660,N_3369,N_5664);
xor U7661 (N_7661,N_3999,N_5081);
nor U7662 (N_7662,N_5439,N_4776);
and U7663 (N_7663,N_4105,N_4302);
or U7664 (N_7664,N_3844,N_4048);
nand U7665 (N_7665,N_3530,N_3013);
or U7666 (N_7666,N_4259,N_4506);
nand U7667 (N_7667,N_4904,N_5619);
nor U7668 (N_7668,N_4275,N_4510);
and U7669 (N_7669,N_4606,N_5773);
xnor U7670 (N_7670,N_4403,N_4899);
or U7671 (N_7671,N_3162,N_3692);
and U7672 (N_7672,N_3314,N_4993);
nor U7673 (N_7673,N_4949,N_5323);
nor U7674 (N_7674,N_3726,N_5748);
nor U7675 (N_7675,N_4553,N_5243);
nand U7676 (N_7676,N_3119,N_3543);
nor U7677 (N_7677,N_3619,N_5085);
xor U7678 (N_7678,N_3366,N_4363);
or U7679 (N_7679,N_5162,N_5032);
nor U7680 (N_7680,N_4701,N_5667);
xnor U7681 (N_7681,N_5753,N_4813);
nand U7682 (N_7682,N_4180,N_3356);
and U7683 (N_7683,N_4736,N_4689);
nand U7684 (N_7684,N_3305,N_4941);
nor U7685 (N_7685,N_4244,N_5535);
nand U7686 (N_7686,N_4589,N_3136);
or U7687 (N_7687,N_5001,N_5642);
nand U7688 (N_7688,N_4342,N_3243);
nand U7689 (N_7689,N_3918,N_3442);
and U7690 (N_7690,N_4874,N_4184);
nand U7691 (N_7691,N_3919,N_4957);
nor U7692 (N_7692,N_3004,N_4291);
and U7693 (N_7693,N_4452,N_3025);
nor U7694 (N_7694,N_4890,N_3243);
nor U7695 (N_7695,N_4669,N_5660);
and U7696 (N_7696,N_3938,N_4953);
xor U7697 (N_7697,N_3747,N_3673);
and U7698 (N_7698,N_4735,N_4255);
or U7699 (N_7699,N_5198,N_5848);
and U7700 (N_7700,N_5539,N_4423);
nand U7701 (N_7701,N_5222,N_3111);
nor U7702 (N_7702,N_3902,N_4269);
nand U7703 (N_7703,N_3402,N_5116);
or U7704 (N_7704,N_5834,N_5906);
nor U7705 (N_7705,N_4040,N_3035);
nor U7706 (N_7706,N_5058,N_4256);
xnor U7707 (N_7707,N_3219,N_4934);
or U7708 (N_7708,N_3918,N_4207);
xor U7709 (N_7709,N_5324,N_3029);
nor U7710 (N_7710,N_4683,N_5154);
nand U7711 (N_7711,N_4186,N_4615);
and U7712 (N_7712,N_5985,N_3523);
xor U7713 (N_7713,N_4997,N_3682);
or U7714 (N_7714,N_3140,N_4319);
and U7715 (N_7715,N_5304,N_3580);
xor U7716 (N_7716,N_5464,N_5091);
and U7717 (N_7717,N_5157,N_4364);
and U7718 (N_7718,N_3522,N_4623);
or U7719 (N_7719,N_5207,N_4150);
nand U7720 (N_7720,N_5367,N_4518);
nor U7721 (N_7721,N_4215,N_3927);
nor U7722 (N_7722,N_4010,N_4773);
xnor U7723 (N_7723,N_4054,N_4669);
nor U7724 (N_7724,N_3675,N_5833);
nand U7725 (N_7725,N_3584,N_5989);
or U7726 (N_7726,N_4991,N_5573);
or U7727 (N_7727,N_4887,N_3156);
nand U7728 (N_7728,N_3470,N_4462);
xnor U7729 (N_7729,N_3251,N_5487);
xor U7730 (N_7730,N_3123,N_5864);
and U7731 (N_7731,N_3096,N_3975);
xor U7732 (N_7732,N_3877,N_3225);
and U7733 (N_7733,N_3330,N_5610);
nand U7734 (N_7734,N_4040,N_3546);
or U7735 (N_7735,N_3559,N_4838);
or U7736 (N_7736,N_3687,N_5493);
nand U7737 (N_7737,N_4626,N_4882);
nand U7738 (N_7738,N_4403,N_3500);
nand U7739 (N_7739,N_3374,N_5777);
or U7740 (N_7740,N_4833,N_3849);
nand U7741 (N_7741,N_4727,N_4945);
nor U7742 (N_7742,N_4794,N_4376);
nor U7743 (N_7743,N_5216,N_5652);
and U7744 (N_7744,N_3919,N_3800);
or U7745 (N_7745,N_3777,N_5672);
or U7746 (N_7746,N_4038,N_3522);
and U7747 (N_7747,N_5874,N_3819);
nor U7748 (N_7748,N_5530,N_3525);
nor U7749 (N_7749,N_4660,N_5931);
nand U7750 (N_7750,N_3440,N_4747);
xor U7751 (N_7751,N_4967,N_5275);
nand U7752 (N_7752,N_5614,N_5162);
or U7753 (N_7753,N_4343,N_4764);
nand U7754 (N_7754,N_3602,N_4589);
nor U7755 (N_7755,N_3375,N_4492);
nand U7756 (N_7756,N_5533,N_4876);
and U7757 (N_7757,N_3501,N_3342);
nor U7758 (N_7758,N_3870,N_4883);
nand U7759 (N_7759,N_3266,N_5284);
nor U7760 (N_7760,N_3807,N_3738);
nand U7761 (N_7761,N_5060,N_5937);
and U7762 (N_7762,N_4538,N_3774);
nand U7763 (N_7763,N_3158,N_3236);
nor U7764 (N_7764,N_4055,N_4162);
or U7765 (N_7765,N_4775,N_5573);
nor U7766 (N_7766,N_3581,N_3278);
nand U7767 (N_7767,N_3808,N_5709);
nor U7768 (N_7768,N_4346,N_5312);
xor U7769 (N_7769,N_5169,N_4758);
or U7770 (N_7770,N_3761,N_3133);
or U7771 (N_7771,N_4392,N_4696);
nor U7772 (N_7772,N_3959,N_4211);
nor U7773 (N_7773,N_5461,N_4281);
and U7774 (N_7774,N_3339,N_3047);
xnor U7775 (N_7775,N_4838,N_3599);
or U7776 (N_7776,N_5948,N_3031);
and U7777 (N_7777,N_5938,N_4380);
and U7778 (N_7778,N_4555,N_4227);
and U7779 (N_7779,N_4789,N_4681);
or U7780 (N_7780,N_4043,N_5759);
nand U7781 (N_7781,N_3156,N_5915);
and U7782 (N_7782,N_4078,N_5454);
xor U7783 (N_7783,N_5122,N_4793);
and U7784 (N_7784,N_4194,N_5990);
or U7785 (N_7785,N_5782,N_5369);
or U7786 (N_7786,N_3482,N_5925);
nor U7787 (N_7787,N_5737,N_5409);
nand U7788 (N_7788,N_3308,N_5211);
and U7789 (N_7789,N_5802,N_4566);
nand U7790 (N_7790,N_3677,N_5858);
or U7791 (N_7791,N_4163,N_4891);
nor U7792 (N_7792,N_5251,N_5376);
nand U7793 (N_7793,N_4411,N_5939);
or U7794 (N_7794,N_5246,N_4499);
nand U7795 (N_7795,N_3334,N_5740);
and U7796 (N_7796,N_3490,N_4839);
or U7797 (N_7797,N_5781,N_4291);
or U7798 (N_7798,N_3990,N_3777);
or U7799 (N_7799,N_3977,N_3712);
nand U7800 (N_7800,N_5381,N_4585);
nor U7801 (N_7801,N_4062,N_3120);
xor U7802 (N_7802,N_3828,N_3006);
or U7803 (N_7803,N_4301,N_3691);
nand U7804 (N_7804,N_3198,N_4692);
and U7805 (N_7805,N_4690,N_3008);
xnor U7806 (N_7806,N_3443,N_4418);
nand U7807 (N_7807,N_3327,N_4195);
nor U7808 (N_7808,N_3963,N_3578);
nor U7809 (N_7809,N_5064,N_5274);
and U7810 (N_7810,N_3448,N_5610);
nor U7811 (N_7811,N_5973,N_4216);
xnor U7812 (N_7812,N_3615,N_3556);
nand U7813 (N_7813,N_4788,N_3055);
nor U7814 (N_7814,N_4835,N_5234);
nor U7815 (N_7815,N_5551,N_5998);
nand U7816 (N_7816,N_3525,N_3728);
and U7817 (N_7817,N_3796,N_3961);
nand U7818 (N_7818,N_5493,N_5548);
nor U7819 (N_7819,N_3073,N_3662);
or U7820 (N_7820,N_4460,N_5764);
nor U7821 (N_7821,N_4592,N_3037);
nand U7822 (N_7822,N_3118,N_5644);
nor U7823 (N_7823,N_3538,N_4976);
nand U7824 (N_7824,N_4855,N_4560);
nor U7825 (N_7825,N_4022,N_4244);
or U7826 (N_7826,N_4091,N_5881);
nand U7827 (N_7827,N_3584,N_5485);
or U7828 (N_7828,N_5214,N_3573);
and U7829 (N_7829,N_5999,N_3162);
nand U7830 (N_7830,N_3698,N_4746);
or U7831 (N_7831,N_4325,N_5498);
nand U7832 (N_7832,N_4989,N_4129);
and U7833 (N_7833,N_3981,N_4470);
or U7834 (N_7834,N_5546,N_3258);
nor U7835 (N_7835,N_5609,N_5875);
and U7836 (N_7836,N_3688,N_5062);
and U7837 (N_7837,N_3958,N_4257);
nand U7838 (N_7838,N_5901,N_3302);
or U7839 (N_7839,N_4038,N_3449);
and U7840 (N_7840,N_5412,N_4079);
nand U7841 (N_7841,N_3360,N_5091);
or U7842 (N_7842,N_4786,N_4325);
or U7843 (N_7843,N_5308,N_4130);
nor U7844 (N_7844,N_5520,N_4918);
and U7845 (N_7845,N_4952,N_3637);
or U7846 (N_7846,N_4867,N_4500);
nor U7847 (N_7847,N_3813,N_3391);
nor U7848 (N_7848,N_4551,N_4286);
nand U7849 (N_7849,N_5217,N_5510);
and U7850 (N_7850,N_4077,N_3917);
nand U7851 (N_7851,N_4196,N_5228);
or U7852 (N_7852,N_5179,N_4011);
nor U7853 (N_7853,N_3696,N_3709);
and U7854 (N_7854,N_5164,N_4424);
or U7855 (N_7855,N_4287,N_3695);
nand U7856 (N_7856,N_5999,N_3741);
nor U7857 (N_7857,N_3857,N_4442);
and U7858 (N_7858,N_3453,N_4635);
nand U7859 (N_7859,N_3842,N_3265);
xor U7860 (N_7860,N_4094,N_3886);
xnor U7861 (N_7861,N_5637,N_5003);
or U7862 (N_7862,N_5345,N_3318);
nor U7863 (N_7863,N_5164,N_3542);
nor U7864 (N_7864,N_3398,N_3208);
nor U7865 (N_7865,N_4899,N_5738);
and U7866 (N_7866,N_5360,N_4689);
or U7867 (N_7867,N_4053,N_3697);
and U7868 (N_7868,N_3658,N_3215);
and U7869 (N_7869,N_5578,N_5920);
or U7870 (N_7870,N_3540,N_3725);
or U7871 (N_7871,N_3998,N_5332);
nand U7872 (N_7872,N_5371,N_3814);
and U7873 (N_7873,N_3740,N_4410);
nand U7874 (N_7874,N_3920,N_3758);
or U7875 (N_7875,N_4637,N_3801);
nor U7876 (N_7876,N_3095,N_3842);
nor U7877 (N_7877,N_5391,N_5350);
nor U7878 (N_7878,N_4876,N_5575);
nor U7879 (N_7879,N_3904,N_4671);
nor U7880 (N_7880,N_4475,N_3642);
or U7881 (N_7881,N_4159,N_5515);
or U7882 (N_7882,N_5289,N_4658);
and U7883 (N_7883,N_5437,N_3239);
or U7884 (N_7884,N_4898,N_5892);
nor U7885 (N_7885,N_3541,N_4001);
nor U7886 (N_7886,N_5742,N_5834);
nand U7887 (N_7887,N_5009,N_3411);
and U7888 (N_7888,N_3942,N_4791);
or U7889 (N_7889,N_4429,N_4265);
nand U7890 (N_7890,N_3345,N_4730);
nand U7891 (N_7891,N_4732,N_3273);
or U7892 (N_7892,N_5035,N_4798);
nor U7893 (N_7893,N_4203,N_5115);
or U7894 (N_7894,N_5509,N_4125);
nand U7895 (N_7895,N_3119,N_3624);
and U7896 (N_7896,N_3273,N_3599);
nor U7897 (N_7897,N_4319,N_5119);
nand U7898 (N_7898,N_4451,N_3408);
nand U7899 (N_7899,N_4621,N_4095);
nor U7900 (N_7900,N_3995,N_5833);
and U7901 (N_7901,N_4783,N_4542);
or U7902 (N_7902,N_4586,N_4743);
nor U7903 (N_7903,N_4283,N_4498);
or U7904 (N_7904,N_3232,N_3158);
or U7905 (N_7905,N_3820,N_4545);
and U7906 (N_7906,N_4831,N_4076);
and U7907 (N_7907,N_4832,N_5230);
nand U7908 (N_7908,N_5364,N_5793);
and U7909 (N_7909,N_3662,N_3191);
nand U7910 (N_7910,N_5887,N_5215);
or U7911 (N_7911,N_3299,N_5242);
and U7912 (N_7912,N_5896,N_5340);
nand U7913 (N_7913,N_5179,N_4680);
or U7914 (N_7914,N_5745,N_3670);
and U7915 (N_7915,N_4793,N_4980);
or U7916 (N_7916,N_5826,N_5232);
and U7917 (N_7917,N_5029,N_5910);
nand U7918 (N_7918,N_3771,N_4242);
or U7919 (N_7919,N_5077,N_4939);
or U7920 (N_7920,N_5638,N_3519);
nor U7921 (N_7921,N_4035,N_5942);
and U7922 (N_7922,N_4078,N_5424);
and U7923 (N_7923,N_3503,N_4596);
nand U7924 (N_7924,N_5465,N_5707);
and U7925 (N_7925,N_3458,N_4531);
and U7926 (N_7926,N_4295,N_3559);
nor U7927 (N_7927,N_4466,N_3282);
nor U7928 (N_7928,N_4885,N_4894);
nor U7929 (N_7929,N_3177,N_3742);
nor U7930 (N_7930,N_4778,N_3539);
or U7931 (N_7931,N_5314,N_4157);
or U7932 (N_7932,N_3964,N_4608);
nand U7933 (N_7933,N_3419,N_5461);
nand U7934 (N_7934,N_3744,N_3521);
xor U7935 (N_7935,N_5923,N_4378);
nor U7936 (N_7936,N_3064,N_4652);
nor U7937 (N_7937,N_3354,N_3431);
and U7938 (N_7938,N_3073,N_3370);
nor U7939 (N_7939,N_3498,N_4065);
nor U7940 (N_7940,N_4696,N_4038);
and U7941 (N_7941,N_3657,N_4194);
nand U7942 (N_7942,N_3956,N_3076);
nand U7943 (N_7943,N_5136,N_3492);
xnor U7944 (N_7944,N_3972,N_4468);
or U7945 (N_7945,N_4889,N_3972);
nor U7946 (N_7946,N_5976,N_4674);
nor U7947 (N_7947,N_4833,N_5182);
nand U7948 (N_7948,N_3422,N_5154);
nand U7949 (N_7949,N_3940,N_4595);
and U7950 (N_7950,N_5552,N_4999);
and U7951 (N_7951,N_5376,N_4844);
xor U7952 (N_7952,N_3779,N_4871);
and U7953 (N_7953,N_5663,N_5241);
xnor U7954 (N_7954,N_4665,N_4130);
nor U7955 (N_7955,N_4899,N_3928);
and U7956 (N_7956,N_5343,N_3164);
and U7957 (N_7957,N_4094,N_4934);
xnor U7958 (N_7958,N_5330,N_5609);
nand U7959 (N_7959,N_4409,N_4544);
nor U7960 (N_7960,N_3353,N_4489);
or U7961 (N_7961,N_5149,N_4067);
or U7962 (N_7962,N_3300,N_4071);
xor U7963 (N_7963,N_4673,N_4841);
nand U7964 (N_7964,N_5140,N_3789);
nor U7965 (N_7965,N_3672,N_4392);
and U7966 (N_7966,N_4761,N_3897);
nor U7967 (N_7967,N_5253,N_3046);
or U7968 (N_7968,N_4065,N_3767);
and U7969 (N_7969,N_4380,N_4878);
nand U7970 (N_7970,N_5587,N_4992);
nand U7971 (N_7971,N_3200,N_4765);
or U7972 (N_7972,N_4606,N_5040);
nand U7973 (N_7973,N_5142,N_5778);
nor U7974 (N_7974,N_5923,N_4029);
nand U7975 (N_7975,N_5951,N_4871);
or U7976 (N_7976,N_3000,N_3621);
nand U7977 (N_7977,N_4976,N_4067);
or U7978 (N_7978,N_3798,N_3555);
nand U7979 (N_7979,N_5289,N_3056);
nand U7980 (N_7980,N_3014,N_5223);
or U7981 (N_7981,N_5700,N_3698);
and U7982 (N_7982,N_5757,N_4419);
or U7983 (N_7983,N_4627,N_4532);
xnor U7984 (N_7984,N_5311,N_4555);
or U7985 (N_7985,N_5165,N_4848);
and U7986 (N_7986,N_3107,N_3192);
xnor U7987 (N_7987,N_3065,N_5343);
or U7988 (N_7988,N_5946,N_4432);
or U7989 (N_7989,N_3728,N_4604);
nor U7990 (N_7990,N_5265,N_4784);
nor U7991 (N_7991,N_3192,N_5950);
nand U7992 (N_7992,N_5767,N_3707);
xor U7993 (N_7993,N_3244,N_4927);
nor U7994 (N_7994,N_4760,N_5163);
nor U7995 (N_7995,N_4218,N_5370);
or U7996 (N_7996,N_4187,N_3324);
or U7997 (N_7997,N_5773,N_5604);
nand U7998 (N_7998,N_5668,N_5349);
nor U7999 (N_7999,N_5959,N_3566);
nand U8000 (N_8000,N_5045,N_4508);
nor U8001 (N_8001,N_5410,N_5836);
nor U8002 (N_8002,N_5486,N_5382);
and U8003 (N_8003,N_4288,N_4976);
or U8004 (N_8004,N_4832,N_5353);
or U8005 (N_8005,N_3285,N_5352);
nor U8006 (N_8006,N_3460,N_4708);
and U8007 (N_8007,N_3889,N_4100);
or U8008 (N_8008,N_4641,N_5274);
or U8009 (N_8009,N_5866,N_3535);
and U8010 (N_8010,N_3703,N_5345);
or U8011 (N_8011,N_4403,N_4822);
nand U8012 (N_8012,N_4857,N_3753);
nand U8013 (N_8013,N_3786,N_4477);
or U8014 (N_8014,N_4914,N_3793);
and U8015 (N_8015,N_4039,N_5762);
nand U8016 (N_8016,N_4979,N_5825);
or U8017 (N_8017,N_4805,N_3625);
nand U8018 (N_8018,N_4466,N_5250);
nor U8019 (N_8019,N_3283,N_3659);
and U8020 (N_8020,N_3770,N_3422);
nand U8021 (N_8021,N_4938,N_4275);
nand U8022 (N_8022,N_4431,N_4600);
nand U8023 (N_8023,N_3721,N_4469);
xor U8024 (N_8024,N_4228,N_5325);
or U8025 (N_8025,N_5866,N_5174);
nor U8026 (N_8026,N_3023,N_4409);
nand U8027 (N_8027,N_4812,N_5695);
nand U8028 (N_8028,N_3287,N_5602);
or U8029 (N_8029,N_5239,N_4975);
and U8030 (N_8030,N_4842,N_3550);
nor U8031 (N_8031,N_3662,N_3558);
nand U8032 (N_8032,N_4531,N_4409);
nand U8033 (N_8033,N_4590,N_5132);
nand U8034 (N_8034,N_4803,N_4164);
or U8035 (N_8035,N_5872,N_4664);
nor U8036 (N_8036,N_3657,N_3712);
nand U8037 (N_8037,N_3584,N_4939);
nand U8038 (N_8038,N_4129,N_4816);
nor U8039 (N_8039,N_4483,N_4118);
or U8040 (N_8040,N_4153,N_3537);
or U8041 (N_8041,N_3347,N_5237);
nor U8042 (N_8042,N_3163,N_3758);
or U8043 (N_8043,N_5276,N_3758);
and U8044 (N_8044,N_4884,N_5679);
nor U8045 (N_8045,N_3580,N_3606);
nand U8046 (N_8046,N_4569,N_3424);
nand U8047 (N_8047,N_4058,N_4663);
and U8048 (N_8048,N_5530,N_3846);
or U8049 (N_8049,N_4335,N_3699);
nor U8050 (N_8050,N_4011,N_3150);
nor U8051 (N_8051,N_3027,N_5915);
and U8052 (N_8052,N_5036,N_3110);
and U8053 (N_8053,N_5490,N_4633);
and U8054 (N_8054,N_3637,N_3199);
and U8055 (N_8055,N_3511,N_4924);
nor U8056 (N_8056,N_3636,N_5586);
nand U8057 (N_8057,N_4826,N_5449);
nand U8058 (N_8058,N_4884,N_3446);
or U8059 (N_8059,N_4638,N_4582);
nand U8060 (N_8060,N_5734,N_4602);
nor U8061 (N_8061,N_4998,N_4322);
nand U8062 (N_8062,N_5752,N_4904);
nor U8063 (N_8063,N_3326,N_5018);
nor U8064 (N_8064,N_4822,N_3501);
or U8065 (N_8065,N_3032,N_4144);
and U8066 (N_8066,N_4112,N_4831);
xor U8067 (N_8067,N_4222,N_3161);
nor U8068 (N_8068,N_3261,N_5140);
nor U8069 (N_8069,N_4698,N_5739);
and U8070 (N_8070,N_5996,N_4535);
and U8071 (N_8071,N_3270,N_3211);
and U8072 (N_8072,N_3850,N_3521);
and U8073 (N_8073,N_4402,N_3405);
and U8074 (N_8074,N_4381,N_3778);
and U8075 (N_8075,N_5162,N_4523);
nand U8076 (N_8076,N_4247,N_3392);
and U8077 (N_8077,N_5340,N_4795);
nor U8078 (N_8078,N_5168,N_4892);
nor U8079 (N_8079,N_4216,N_3729);
or U8080 (N_8080,N_4596,N_5773);
or U8081 (N_8081,N_3178,N_4228);
and U8082 (N_8082,N_4967,N_4715);
xor U8083 (N_8083,N_5885,N_4270);
nand U8084 (N_8084,N_4157,N_3337);
nand U8085 (N_8085,N_5582,N_4266);
nor U8086 (N_8086,N_5919,N_4695);
and U8087 (N_8087,N_5571,N_4009);
or U8088 (N_8088,N_3904,N_4444);
and U8089 (N_8089,N_4255,N_3704);
nor U8090 (N_8090,N_5804,N_5430);
nor U8091 (N_8091,N_4716,N_5121);
nor U8092 (N_8092,N_3866,N_4476);
and U8093 (N_8093,N_4727,N_4795);
or U8094 (N_8094,N_3654,N_4596);
nand U8095 (N_8095,N_5288,N_5203);
or U8096 (N_8096,N_4601,N_5952);
xor U8097 (N_8097,N_3103,N_4786);
xnor U8098 (N_8098,N_5636,N_4908);
and U8099 (N_8099,N_4544,N_4956);
xnor U8100 (N_8100,N_4996,N_3493);
xnor U8101 (N_8101,N_3053,N_5315);
and U8102 (N_8102,N_4311,N_4301);
nand U8103 (N_8103,N_5635,N_4040);
and U8104 (N_8104,N_5566,N_4615);
nand U8105 (N_8105,N_5994,N_3665);
nor U8106 (N_8106,N_5051,N_5370);
nand U8107 (N_8107,N_4698,N_3568);
nor U8108 (N_8108,N_3324,N_4142);
nand U8109 (N_8109,N_5937,N_5223);
nand U8110 (N_8110,N_4945,N_3847);
nor U8111 (N_8111,N_3902,N_3569);
nand U8112 (N_8112,N_3103,N_4595);
nand U8113 (N_8113,N_3789,N_5265);
nor U8114 (N_8114,N_5678,N_3856);
and U8115 (N_8115,N_5270,N_5981);
and U8116 (N_8116,N_3362,N_5022);
nor U8117 (N_8117,N_5900,N_5892);
nand U8118 (N_8118,N_3029,N_4234);
nand U8119 (N_8119,N_4567,N_3227);
nor U8120 (N_8120,N_3359,N_3531);
nor U8121 (N_8121,N_3885,N_5040);
and U8122 (N_8122,N_5042,N_5231);
or U8123 (N_8123,N_5456,N_3630);
nand U8124 (N_8124,N_4975,N_4545);
and U8125 (N_8125,N_5928,N_5702);
nand U8126 (N_8126,N_3608,N_5802);
and U8127 (N_8127,N_3834,N_3959);
nor U8128 (N_8128,N_5483,N_5875);
or U8129 (N_8129,N_5484,N_5344);
nand U8130 (N_8130,N_4520,N_4020);
nand U8131 (N_8131,N_4384,N_5539);
or U8132 (N_8132,N_4521,N_3082);
xnor U8133 (N_8133,N_5120,N_4617);
xor U8134 (N_8134,N_4560,N_3509);
xor U8135 (N_8135,N_3771,N_3210);
and U8136 (N_8136,N_3940,N_4900);
nand U8137 (N_8137,N_5846,N_3677);
and U8138 (N_8138,N_3769,N_3238);
xor U8139 (N_8139,N_3156,N_4423);
or U8140 (N_8140,N_3739,N_3849);
and U8141 (N_8141,N_5339,N_3939);
or U8142 (N_8142,N_5608,N_5209);
nor U8143 (N_8143,N_3167,N_3873);
or U8144 (N_8144,N_3445,N_4862);
and U8145 (N_8145,N_3253,N_5770);
nor U8146 (N_8146,N_3021,N_3459);
nor U8147 (N_8147,N_3890,N_5412);
or U8148 (N_8148,N_5690,N_4585);
or U8149 (N_8149,N_4373,N_4603);
or U8150 (N_8150,N_4773,N_5301);
and U8151 (N_8151,N_3110,N_3502);
nand U8152 (N_8152,N_3554,N_4488);
nand U8153 (N_8153,N_5644,N_4524);
and U8154 (N_8154,N_5769,N_5563);
nor U8155 (N_8155,N_4616,N_3207);
xor U8156 (N_8156,N_5539,N_5927);
and U8157 (N_8157,N_3839,N_5393);
nand U8158 (N_8158,N_3777,N_3310);
or U8159 (N_8159,N_4671,N_4646);
and U8160 (N_8160,N_4922,N_3067);
nand U8161 (N_8161,N_4950,N_4460);
or U8162 (N_8162,N_4915,N_4920);
and U8163 (N_8163,N_4671,N_3023);
nor U8164 (N_8164,N_3170,N_3223);
or U8165 (N_8165,N_5750,N_3562);
xnor U8166 (N_8166,N_3038,N_3092);
nand U8167 (N_8167,N_5732,N_4860);
or U8168 (N_8168,N_4820,N_4308);
or U8169 (N_8169,N_5087,N_3113);
nor U8170 (N_8170,N_3822,N_4712);
or U8171 (N_8171,N_3609,N_3798);
nand U8172 (N_8172,N_4450,N_5424);
nor U8173 (N_8173,N_3836,N_5542);
nand U8174 (N_8174,N_5975,N_4115);
or U8175 (N_8175,N_5765,N_5268);
or U8176 (N_8176,N_4795,N_4523);
nor U8177 (N_8177,N_3668,N_4623);
nor U8178 (N_8178,N_4973,N_3741);
nor U8179 (N_8179,N_3980,N_3452);
and U8180 (N_8180,N_5290,N_5243);
nor U8181 (N_8181,N_4184,N_4394);
xnor U8182 (N_8182,N_5095,N_4112);
and U8183 (N_8183,N_5918,N_4950);
or U8184 (N_8184,N_3121,N_3559);
or U8185 (N_8185,N_3638,N_5609);
or U8186 (N_8186,N_5761,N_3401);
and U8187 (N_8187,N_5711,N_3144);
nand U8188 (N_8188,N_3067,N_5195);
and U8189 (N_8189,N_4257,N_3661);
and U8190 (N_8190,N_5156,N_5940);
or U8191 (N_8191,N_3635,N_4376);
nor U8192 (N_8192,N_5429,N_3056);
or U8193 (N_8193,N_3155,N_3137);
or U8194 (N_8194,N_4523,N_5112);
and U8195 (N_8195,N_3267,N_3000);
nor U8196 (N_8196,N_4921,N_3475);
nor U8197 (N_8197,N_3170,N_5701);
nor U8198 (N_8198,N_4868,N_5392);
xor U8199 (N_8199,N_4302,N_5562);
and U8200 (N_8200,N_5914,N_5452);
nand U8201 (N_8201,N_3646,N_5435);
nor U8202 (N_8202,N_5484,N_3960);
nand U8203 (N_8203,N_3403,N_5295);
and U8204 (N_8204,N_5471,N_5150);
or U8205 (N_8205,N_3261,N_4112);
or U8206 (N_8206,N_3181,N_5833);
nor U8207 (N_8207,N_5917,N_4613);
or U8208 (N_8208,N_4193,N_5819);
nor U8209 (N_8209,N_4642,N_5399);
and U8210 (N_8210,N_4588,N_4039);
or U8211 (N_8211,N_3727,N_3746);
and U8212 (N_8212,N_5213,N_4468);
and U8213 (N_8213,N_5271,N_3568);
and U8214 (N_8214,N_5235,N_3055);
xnor U8215 (N_8215,N_4667,N_5540);
and U8216 (N_8216,N_5264,N_3019);
nand U8217 (N_8217,N_4224,N_5017);
or U8218 (N_8218,N_5496,N_5400);
and U8219 (N_8219,N_5163,N_4599);
or U8220 (N_8220,N_3793,N_5858);
nor U8221 (N_8221,N_5067,N_4439);
and U8222 (N_8222,N_5293,N_3289);
or U8223 (N_8223,N_3540,N_4055);
or U8224 (N_8224,N_5541,N_5249);
or U8225 (N_8225,N_4747,N_5657);
nand U8226 (N_8226,N_4713,N_5634);
or U8227 (N_8227,N_5264,N_4638);
nor U8228 (N_8228,N_5528,N_3531);
and U8229 (N_8229,N_4373,N_5046);
or U8230 (N_8230,N_5735,N_5292);
or U8231 (N_8231,N_3407,N_3109);
xnor U8232 (N_8232,N_3389,N_5707);
nand U8233 (N_8233,N_5301,N_4223);
nor U8234 (N_8234,N_4636,N_3070);
nor U8235 (N_8235,N_4346,N_3063);
and U8236 (N_8236,N_3964,N_3446);
nor U8237 (N_8237,N_4752,N_4696);
and U8238 (N_8238,N_3851,N_3962);
nor U8239 (N_8239,N_3630,N_3128);
or U8240 (N_8240,N_4232,N_4004);
and U8241 (N_8241,N_4969,N_5887);
nand U8242 (N_8242,N_4780,N_3301);
or U8243 (N_8243,N_3829,N_5380);
nor U8244 (N_8244,N_3098,N_4484);
xnor U8245 (N_8245,N_5583,N_5647);
nand U8246 (N_8246,N_3115,N_5734);
and U8247 (N_8247,N_3014,N_3011);
and U8248 (N_8248,N_5903,N_3811);
nand U8249 (N_8249,N_4744,N_3847);
and U8250 (N_8250,N_5984,N_4873);
and U8251 (N_8251,N_5769,N_3652);
nor U8252 (N_8252,N_4453,N_3456);
nor U8253 (N_8253,N_3846,N_3906);
and U8254 (N_8254,N_3733,N_5979);
and U8255 (N_8255,N_3028,N_4903);
nor U8256 (N_8256,N_5456,N_4856);
and U8257 (N_8257,N_4854,N_3116);
or U8258 (N_8258,N_4491,N_3478);
nor U8259 (N_8259,N_5358,N_5351);
nor U8260 (N_8260,N_5335,N_4453);
nand U8261 (N_8261,N_3959,N_4277);
nor U8262 (N_8262,N_4319,N_5225);
nand U8263 (N_8263,N_4715,N_3186);
and U8264 (N_8264,N_4690,N_3555);
and U8265 (N_8265,N_4428,N_4607);
and U8266 (N_8266,N_4208,N_3197);
and U8267 (N_8267,N_3896,N_4124);
or U8268 (N_8268,N_4104,N_4286);
nand U8269 (N_8269,N_5771,N_3736);
nor U8270 (N_8270,N_5499,N_3095);
nor U8271 (N_8271,N_5225,N_3918);
xnor U8272 (N_8272,N_4661,N_4211);
or U8273 (N_8273,N_5262,N_4545);
nand U8274 (N_8274,N_3605,N_3688);
or U8275 (N_8275,N_5157,N_4233);
or U8276 (N_8276,N_3993,N_3678);
nand U8277 (N_8277,N_4240,N_3701);
and U8278 (N_8278,N_3997,N_4430);
or U8279 (N_8279,N_5496,N_5797);
nand U8280 (N_8280,N_4510,N_5548);
nand U8281 (N_8281,N_4177,N_4528);
nor U8282 (N_8282,N_3136,N_5629);
and U8283 (N_8283,N_4806,N_5691);
or U8284 (N_8284,N_3741,N_5205);
and U8285 (N_8285,N_5619,N_5220);
or U8286 (N_8286,N_5353,N_3846);
nor U8287 (N_8287,N_3230,N_4845);
and U8288 (N_8288,N_3967,N_5898);
nor U8289 (N_8289,N_4953,N_4975);
and U8290 (N_8290,N_5826,N_5224);
or U8291 (N_8291,N_5123,N_5252);
xor U8292 (N_8292,N_5783,N_5009);
nor U8293 (N_8293,N_5669,N_3977);
or U8294 (N_8294,N_4262,N_4677);
nand U8295 (N_8295,N_4901,N_4200);
or U8296 (N_8296,N_3310,N_5102);
nor U8297 (N_8297,N_5452,N_5984);
nand U8298 (N_8298,N_5310,N_3540);
or U8299 (N_8299,N_3018,N_4786);
nand U8300 (N_8300,N_5219,N_3163);
nand U8301 (N_8301,N_4471,N_5044);
nand U8302 (N_8302,N_4079,N_3666);
xnor U8303 (N_8303,N_4817,N_3754);
nor U8304 (N_8304,N_5706,N_5354);
and U8305 (N_8305,N_5102,N_3099);
nand U8306 (N_8306,N_4466,N_3757);
nand U8307 (N_8307,N_4347,N_5572);
nor U8308 (N_8308,N_3105,N_3420);
or U8309 (N_8309,N_3769,N_3997);
nor U8310 (N_8310,N_4198,N_5091);
nor U8311 (N_8311,N_5281,N_4054);
and U8312 (N_8312,N_4821,N_4697);
nor U8313 (N_8313,N_4322,N_4427);
nand U8314 (N_8314,N_5697,N_4491);
and U8315 (N_8315,N_4326,N_3233);
xor U8316 (N_8316,N_4309,N_4286);
and U8317 (N_8317,N_5875,N_5964);
nor U8318 (N_8318,N_3854,N_5610);
nand U8319 (N_8319,N_3742,N_4360);
or U8320 (N_8320,N_5285,N_4447);
and U8321 (N_8321,N_5851,N_5115);
and U8322 (N_8322,N_4301,N_4629);
nor U8323 (N_8323,N_5323,N_4668);
nor U8324 (N_8324,N_5925,N_3202);
or U8325 (N_8325,N_5056,N_3900);
or U8326 (N_8326,N_3271,N_3662);
or U8327 (N_8327,N_5106,N_5789);
nand U8328 (N_8328,N_3091,N_4368);
and U8329 (N_8329,N_5073,N_3899);
nor U8330 (N_8330,N_5377,N_3264);
or U8331 (N_8331,N_4745,N_3313);
or U8332 (N_8332,N_5736,N_4874);
or U8333 (N_8333,N_5056,N_4568);
nor U8334 (N_8334,N_3985,N_4091);
or U8335 (N_8335,N_5326,N_3428);
nor U8336 (N_8336,N_3009,N_3221);
nor U8337 (N_8337,N_4213,N_4677);
and U8338 (N_8338,N_3585,N_4630);
nand U8339 (N_8339,N_3519,N_5844);
nand U8340 (N_8340,N_5613,N_3356);
nor U8341 (N_8341,N_5478,N_5002);
xnor U8342 (N_8342,N_5871,N_4080);
nor U8343 (N_8343,N_5379,N_4482);
xor U8344 (N_8344,N_4119,N_5544);
xor U8345 (N_8345,N_3080,N_3743);
and U8346 (N_8346,N_5310,N_4325);
and U8347 (N_8347,N_5870,N_4689);
nor U8348 (N_8348,N_4161,N_4987);
nand U8349 (N_8349,N_4048,N_3743);
or U8350 (N_8350,N_5784,N_3207);
and U8351 (N_8351,N_5279,N_4570);
nor U8352 (N_8352,N_5328,N_4621);
nor U8353 (N_8353,N_4645,N_4592);
and U8354 (N_8354,N_5407,N_3951);
nand U8355 (N_8355,N_5186,N_5749);
and U8356 (N_8356,N_3067,N_3913);
or U8357 (N_8357,N_3653,N_5116);
or U8358 (N_8358,N_5102,N_4294);
xnor U8359 (N_8359,N_4516,N_4427);
and U8360 (N_8360,N_5836,N_3989);
or U8361 (N_8361,N_5730,N_5443);
or U8362 (N_8362,N_4411,N_4014);
or U8363 (N_8363,N_3015,N_5631);
and U8364 (N_8364,N_3389,N_4329);
or U8365 (N_8365,N_4048,N_4368);
nor U8366 (N_8366,N_5507,N_5992);
or U8367 (N_8367,N_4810,N_4350);
nor U8368 (N_8368,N_4986,N_4546);
nor U8369 (N_8369,N_5465,N_3181);
or U8370 (N_8370,N_4125,N_3296);
or U8371 (N_8371,N_3257,N_5812);
xor U8372 (N_8372,N_4769,N_3578);
nor U8373 (N_8373,N_3235,N_4547);
or U8374 (N_8374,N_4378,N_4005);
xor U8375 (N_8375,N_3470,N_5707);
or U8376 (N_8376,N_3683,N_4675);
or U8377 (N_8377,N_3277,N_3333);
nand U8378 (N_8378,N_3229,N_4140);
nand U8379 (N_8379,N_3119,N_5821);
and U8380 (N_8380,N_4542,N_5885);
and U8381 (N_8381,N_3031,N_4567);
or U8382 (N_8382,N_4195,N_5529);
nor U8383 (N_8383,N_4465,N_3547);
nand U8384 (N_8384,N_5587,N_3976);
nor U8385 (N_8385,N_3887,N_4243);
nand U8386 (N_8386,N_3906,N_5872);
or U8387 (N_8387,N_5896,N_3503);
and U8388 (N_8388,N_3850,N_5474);
nor U8389 (N_8389,N_5462,N_5796);
nand U8390 (N_8390,N_3250,N_3555);
or U8391 (N_8391,N_4423,N_4085);
and U8392 (N_8392,N_5168,N_4210);
nand U8393 (N_8393,N_3052,N_4443);
xnor U8394 (N_8394,N_4588,N_4001);
nor U8395 (N_8395,N_4288,N_3753);
nor U8396 (N_8396,N_3795,N_4591);
and U8397 (N_8397,N_4534,N_3152);
nor U8398 (N_8398,N_3587,N_3654);
nand U8399 (N_8399,N_4076,N_5285);
nand U8400 (N_8400,N_5826,N_3759);
or U8401 (N_8401,N_5792,N_5640);
nor U8402 (N_8402,N_4905,N_4034);
xnor U8403 (N_8403,N_3096,N_4189);
nand U8404 (N_8404,N_5642,N_5716);
and U8405 (N_8405,N_4648,N_3616);
or U8406 (N_8406,N_5776,N_5092);
nand U8407 (N_8407,N_4799,N_3357);
and U8408 (N_8408,N_3751,N_5833);
nor U8409 (N_8409,N_4599,N_3925);
nor U8410 (N_8410,N_3886,N_5491);
nor U8411 (N_8411,N_3705,N_4391);
nand U8412 (N_8412,N_5685,N_4477);
nor U8413 (N_8413,N_5836,N_4858);
nor U8414 (N_8414,N_5898,N_5066);
and U8415 (N_8415,N_3147,N_4786);
xnor U8416 (N_8416,N_3998,N_4498);
and U8417 (N_8417,N_4235,N_4829);
nand U8418 (N_8418,N_5776,N_4054);
nand U8419 (N_8419,N_3630,N_5349);
or U8420 (N_8420,N_5422,N_3633);
or U8421 (N_8421,N_3744,N_5426);
or U8422 (N_8422,N_4707,N_5095);
or U8423 (N_8423,N_4992,N_4337);
xnor U8424 (N_8424,N_3936,N_3695);
or U8425 (N_8425,N_5982,N_5001);
nand U8426 (N_8426,N_5354,N_5785);
or U8427 (N_8427,N_3786,N_3553);
and U8428 (N_8428,N_3870,N_3480);
nor U8429 (N_8429,N_4807,N_4416);
xor U8430 (N_8430,N_5785,N_3842);
nor U8431 (N_8431,N_5404,N_3454);
and U8432 (N_8432,N_3743,N_4751);
nor U8433 (N_8433,N_4508,N_5367);
nand U8434 (N_8434,N_5452,N_5251);
and U8435 (N_8435,N_3238,N_4765);
or U8436 (N_8436,N_4253,N_3257);
nor U8437 (N_8437,N_3716,N_5669);
xor U8438 (N_8438,N_5565,N_4965);
xnor U8439 (N_8439,N_5225,N_3686);
or U8440 (N_8440,N_3925,N_4957);
nand U8441 (N_8441,N_4071,N_5609);
or U8442 (N_8442,N_4225,N_3636);
nor U8443 (N_8443,N_3973,N_5106);
nor U8444 (N_8444,N_5767,N_3326);
and U8445 (N_8445,N_5688,N_4944);
nand U8446 (N_8446,N_5038,N_5194);
nand U8447 (N_8447,N_5854,N_5922);
and U8448 (N_8448,N_3046,N_5087);
nor U8449 (N_8449,N_5959,N_5419);
nand U8450 (N_8450,N_4171,N_3868);
nor U8451 (N_8451,N_4452,N_5446);
or U8452 (N_8452,N_5990,N_5941);
or U8453 (N_8453,N_3509,N_5485);
and U8454 (N_8454,N_4503,N_3659);
and U8455 (N_8455,N_4275,N_3911);
nor U8456 (N_8456,N_4543,N_5423);
nand U8457 (N_8457,N_5034,N_3120);
nor U8458 (N_8458,N_5605,N_4069);
and U8459 (N_8459,N_5548,N_3579);
or U8460 (N_8460,N_4880,N_5542);
nor U8461 (N_8461,N_5690,N_3235);
and U8462 (N_8462,N_4037,N_3786);
and U8463 (N_8463,N_3152,N_3353);
nor U8464 (N_8464,N_4725,N_4278);
nor U8465 (N_8465,N_4868,N_5170);
or U8466 (N_8466,N_3408,N_3973);
nand U8467 (N_8467,N_5944,N_5188);
nor U8468 (N_8468,N_3054,N_5974);
nand U8469 (N_8469,N_5302,N_4494);
nor U8470 (N_8470,N_4536,N_3718);
and U8471 (N_8471,N_5785,N_4739);
or U8472 (N_8472,N_4417,N_4858);
nor U8473 (N_8473,N_4090,N_5613);
nand U8474 (N_8474,N_5715,N_4847);
nor U8475 (N_8475,N_4139,N_3236);
and U8476 (N_8476,N_3814,N_3894);
and U8477 (N_8477,N_3637,N_3386);
and U8478 (N_8478,N_3822,N_4975);
and U8479 (N_8479,N_5599,N_5495);
nand U8480 (N_8480,N_4156,N_3199);
and U8481 (N_8481,N_4299,N_5821);
and U8482 (N_8482,N_5246,N_3759);
or U8483 (N_8483,N_3325,N_4091);
nor U8484 (N_8484,N_3289,N_4083);
nor U8485 (N_8485,N_4055,N_4985);
nor U8486 (N_8486,N_4568,N_5400);
or U8487 (N_8487,N_4033,N_3915);
nand U8488 (N_8488,N_4585,N_5273);
and U8489 (N_8489,N_4281,N_4302);
nor U8490 (N_8490,N_4159,N_4331);
nand U8491 (N_8491,N_4514,N_3770);
nand U8492 (N_8492,N_5552,N_3424);
and U8493 (N_8493,N_3143,N_3396);
xor U8494 (N_8494,N_3813,N_3897);
or U8495 (N_8495,N_5075,N_3179);
or U8496 (N_8496,N_3958,N_5683);
nor U8497 (N_8497,N_3041,N_5712);
and U8498 (N_8498,N_4535,N_3656);
or U8499 (N_8499,N_4653,N_3710);
xnor U8500 (N_8500,N_4636,N_3566);
nand U8501 (N_8501,N_4401,N_5438);
nor U8502 (N_8502,N_5121,N_4368);
and U8503 (N_8503,N_5614,N_4590);
nor U8504 (N_8504,N_5569,N_4264);
nor U8505 (N_8505,N_5518,N_4503);
or U8506 (N_8506,N_3353,N_5934);
and U8507 (N_8507,N_4113,N_4926);
xor U8508 (N_8508,N_3887,N_4390);
nand U8509 (N_8509,N_3529,N_4156);
xor U8510 (N_8510,N_3398,N_5646);
nand U8511 (N_8511,N_3705,N_4166);
and U8512 (N_8512,N_4755,N_4118);
or U8513 (N_8513,N_4137,N_4689);
nor U8514 (N_8514,N_5332,N_3269);
nand U8515 (N_8515,N_4891,N_4611);
nor U8516 (N_8516,N_4721,N_5535);
or U8517 (N_8517,N_4831,N_3636);
nor U8518 (N_8518,N_3986,N_3072);
nand U8519 (N_8519,N_3278,N_5189);
or U8520 (N_8520,N_3845,N_5913);
nor U8521 (N_8521,N_4255,N_5936);
nand U8522 (N_8522,N_4442,N_4002);
and U8523 (N_8523,N_5114,N_4024);
or U8524 (N_8524,N_5082,N_4984);
and U8525 (N_8525,N_3452,N_3639);
nor U8526 (N_8526,N_3583,N_3963);
nand U8527 (N_8527,N_4168,N_4026);
and U8528 (N_8528,N_3715,N_3086);
xnor U8529 (N_8529,N_3227,N_3681);
and U8530 (N_8530,N_4874,N_3020);
or U8531 (N_8531,N_4296,N_5830);
nand U8532 (N_8532,N_3157,N_5791);
and U8533 (N_8533,N_3468,N_3907);
and U8534 (N_8534,N_4420,N_4703);
or U8535 (N_8535,N_5380,N_5209);
and U8536 (N_8536,N_4484,N_3299);
nand U8537 (N_8537,N_5593,N_3169);
xnor U8538 (N_8538,N_5143,N_5254);
or U8539 (N_8539,N_5513,N_3815);
and U8540 (N_8540,N_3320,N_4529);
or U8541 (N_8541,N_3781,N_4081);
and U8542 (N_8542,N_5470,N_4337);
nor U8543 (N_8543,N_3072,N_4661);
nor U8544 (N_8544,N_4537,N_5257);
and U8545 (N_8545,N_4694,N_5301);
or U8546 (N_8546,N_4400,N_3967);
nand U8547 (N_8547,N_3071,N_3832);
and U8548 (N_8548,N_3516,N_5575);
nor U8549 (N_8549,N_4660,N_5891);
nor U8550 (N_8550,N_3222,N_3152);
or U8551 (N_8551,N_4055,N_4811);
and U8552 (N_8552,N_5030,N_3264);
nand U8553 (N_8553,N_5188,N_5170);
nand U8554 (N_8554,N_4138,N_4697);
or U8555 (N_8555,N_5964,N_3183);
nand U8556 (N_8556,N_5621,N_5625);
nand U8557 (N_8557,N_5584,N_5039);
or U8558 (N_8558,N_4911,N_5407);
nand U8559 (N_8559,N_5331,N_5068);
and U8560 (N_8560,N_4520,N_3453);
or U8561 (N_8561,N_5268,N_5904);
nand U8562 (N_8562,N_5208,N_5401);
and U8563 (N_8563,N_3844,N_3337);
or U8564 (N_8564,N_4667,N_4062);
nor U8565 (N_8565,N_4160,N_5435);
nor U8566 (N_8566,N_4843,N_3319);
nand U8567 (N_8567,N_5474,N_3502);
and U8568 (N_8568,N_3989,N_4331);
nor U8569 (N_8569,N_5738,N_3636);
nand U8570 (N_8570,N_4450,N_5800);
or U8571 (N_8571,N_3901,N_3006);
or U8572 (N_8572,N_5635,N_4695);
nor U8573 (N_8573,N_5453,N_3526);
and U8574 (N_8574,N_4976,N_4190);
nand U8575 (N_8575,N_4719,N_5868);
xnor U8576 (N_8576,N_4569,N_4657);
and U8577 (N_8577,N_5097,N_5051);
or U8578 (N_8578,N_3064,N_3578);
xor U8579 (N_8579,N_4840,N_3861);
and U8580 (N_8580,N_4724,N_5658);
and U8581 (N_8581,N_3866,N_4247);
nor U8582 (N_8582,N_4191,N_5386);
nand U8583 (N_8583,N_4794,N_3450);
xnor U8584 (N_8584,N_4988,N_4077);
or U8585 (N_8585,N_3570,N_5999);
xnor U8586 (N_8586,N_5891,N_4296);
nor U8587 (N_8587,N_3862,N_4748);
or U8588 (N_8588,N_5682,N_3817);
xnor U8589 (N_8589,N_3219,N_3613);
or U8590 (N_8590,N_5132,N_3489);
xor U8591 (N_8591,N_4073,N_3664);
or U8592 (N_8592,N_3414,N_4187);
or U8593 (N_8593,N_3870,N_5588);
nand U8594 (N_8594,N_4642,N_3908);
and U8595 (N_8595,N_3556,N_4128);
and U8596 (N_8596,N_5769,N_4521);
and U8597 (N_8597,N_5874,N_3155);
or U8598 (N_8598,N_4704,N_4140);
nand U8599 (N_8599,N_5858,N_3241);
nand U8600 (N_8600,N_3139,N_4672);
nand U8601 (N_8601,N_4145,N_5926);
and U8602 (N_8602,N_4372,N_4193);
or U8603 (N_8603,N_5222,N_4288);
and U8604 (N_8604,N_5693,N_3020);
and U8605 (N_8605,N_3422,N_3156);
nand U8606 (N_8606,N_4006,N_4668);
nor U8607 (N_8607,N_3748,N_3871);
or U8608 (N_8608,N_4704,N_5844);
and U8609 (N_8609,N_4964,N_5640);
and U8610 (N_8610,N_3810,N_4960);
and U8611 (N_8611,N_5599,N_3381);
or U8612 (N_8612,N_3232,N_4581);
nor U8613 (N_8613,N_4197,N_5466);
xnor U8614 (N_8614,N_3907,N_3699);
or U8615 (N_8615,N_5121,N_3565);
nand U8616 (N_8616,N_5427,N_4441);
and U8617 (N_8617,N_3372,N_4723);
nand U8618 (N_8618,N_5287,N_3426);
nand U8619 (N_8619,N_5258,N_3957);
and U8620 (N_8620,N_5165,N_3964);
xnor U8621 (N_8621,N_3179,N_5797);
and U8622 (N_8622,N_4635,N_5996);
nor U8623 (N_8623,N_5981,N_3135);
or U8624 (N_8624,N_3021,N_3887);
or U8625 (N_8625,N_3528,N_5993);
nand U8626 (N_8626,N_5926,N_5446);
nand U8627 (N_8627,N_3323,N_5186);
nor U8628 (N_8628,N_3683,N_4328);
xor U8629 (N_8629,N_4321,N_3300);
nand U8630 (N_8630,N_3001,N_5496);
and U8631 (N_8631,N_5019,N_5083);
xor U8632 (N_8632,N_5584,N_5435);
nand U8633 (N_8633,N_4145,N_5681);
xnor U8634 (N_8634,N_5465,N_5326);
nor U8635 (N_8635,N_5866,N_5743);
or U8636 (N_8636,N_5989,N_5430);
nor U8637 (N_8637,N_3425,N_5764);
or U8638 (N_8638,N_4394,N_5732);
or U8639 (N_8639,N_3318,N_4152);
and U8640 (N_8640,N_4299,N_5694);
and U8641 (N_8641,N_4425,N_4962);
nand U8642 (N_8642,N_3511,N_5594);
nor U8643 (N_8643,N_5399,N_5567);
xnor U8644 (N_8644,N_5468,N_5341);
or U8645 (N_8645,N_5174,N_3714);
nand U8646 (N_8646,N_5876,N_5864);
or U8647 (N_8647,N_5491,N_5560);
xnor U8648 (N_8648,N_3132,N_4400);
nand U8649 (N_8649,N_3104,N_5125);
or U8650 (N_8650,N_5847,N_3721);
nand U8651 (N_8651,N_5082,N_4619);
and U8652 (N_8652,N_5011,N_3696);
and U8653 (N_8653,N_5129,N_4806);
nand U8654 (N_8654,N_4429,N_5281);
or U8655 (N_8655,N_4612,N_4428);
nand U8656 (N_8656,N_4589,N_3089);
and U8657 (N_8657,N_4184,N_5831);
nand U8658 (N_8658,N_3879,N_5301);
nor U8659 (N_8659,N_4185,N_5372);
nand U8660 (N_8660,N_5152,N_5888);
nor U8661 (N_8661,N_3253,N_5094);
xnor U8662 (N_8662,N_3149,N_5595);
nand U8663 (N_8663,N_4045,N_3617);
and U8664 (N_8664,N_5992,N_3634);
or U8665 (N_8665,N_5641,N_3867);
nand U8666 (N_8666,N_3133,N_3609);
or U8667 (N_8667,N_4674,N_4402);
and U8668 (N_8668,N_3686,N_3606);
nand U8669 (N_8669,N_3482,N_4592);
nor U8670 (N_8670,N_3976,N_3010);
nor U8671 (N_8671,N_3736,N_3179);
and U8672 (N_8672,N_3513,N_5679);
xnor U8673 (N_8673,N_3436,N_5005);
nand U8674 (N_8674,N_5879,N_5071);
and U8675 (N_8675,N_5634,N_3802);
nand U8676 (N_8676,N_4657,N_4232);
nand U8677 (N_8677,N_5046,N_5976);
or U8678 (N_8678,N_5252,N_5983);
nand U8679 (N_8679,N_4970,N_3958);
nand U8680 (N_8680,N_3339,N_4378);
or U8681 (N_8681,N_3375,N_4255);
xor U8682 (N_8682,N_3081,N_4365);
nand U8683 (N_8683,N_5134,N_4903);
nand U8684 (N_8684,N_4827,N_5770);
nor U8685 (N_8685,N_4350,N_5086);
and U8686 (N_8686,N_4935,N_4348);
nand U8687 (N_8687,N_5523,N_3663);
and U8688 (N_8688,N_4259,N_5293);
or U8689 (N_8689,N_5644,N_3567);
nor U8690 (N_8690,N_5876,N_5966);
or U8691 (N_8691,N_3544,N_4312);
or U8692 (N_8692,N_3734,N_4160);
nand U8693 (N_8693,N_4969,N_5212);
nor U8694 (N_8694,N_5650,N_4454);
nand U8695 (N_8695,N_3421,N_5740);
or U8696 (N_8696,N_3389,N_5844);
and U8697 (N_8697,N_3689,N_3846);
or U8698 (N_8698,N_3864,N_3693);
nand U8699 (N_8699,N_4649,N_3974);
xnor U8700 (N_8700,N_3860,N_5422);
nand U8701 (N_8701,N_3329,N_3566);
and U8702 (N_8702,N_5038,N_4460);
and U8703 (N_8703,N_3055,N_5753);
nor U8704 (N_8704,N_5030,N_5595);
nor U8705 (N_8705,N_4234,N_3469);
or U8706 (N_8706,N_5539,N_4634);
or U8707 (N_8707,N_4239,N_4422);
or U8708 (N_8708,N_3244,N_3548);
or U8709 (N_8709,N_4454,N_4267);
or U8710 (N_8710,N_5791,N_3328);
nand U8711 (N_8711,N_5978,N_3098);
nand U8712 (N_8712,N_5714,N_4310);
and U8713 (N_8713,N_3540,N_3374);
and U8714 (N_8714,N_3701,N_5079);
nand U8715 (N_8715,N_5701,N_4282);
or U8716 (N_8716,N_3786,N_5358);
and U8717 (N_8717,N_3932,N_4479);
and U8718 (N_8718,N_4737,N_5654);
nor U8719 (N_8719,N_3423,N_5146);
nand U8720 (N_8720,N_5200,N_5160);
xor U8721 (N_8721,N_5778,N_5174);
nand U8722 (N_8722,N_5079,N_5100);
nand U8723 (N_8723,N_4423,N_5775);
or U8724 (N_8724,N_4533,N_4298);
and U8725 (N_8725,N_4911,N_4807);
and U8726 (N_8726,N_3425,N_3293);
and U8727 (N_8727,N_4514,N_4438);
nand U8728 (N_8728,N_4684,N_4705);
or U8729 (N_8729,N_4755,N_5947);
xor U8730 (N_8730,N_3813,N_3500);
or U8731 (N_8731,N_3133,N_3443);
and U8732 (N_8732,N_5030,N_3910);
or U8733 (N_8733,N_4037,N_3471);
and U8734 (N_8734,N_5910,N_5521);
nor U8735 (N_8735,N_5270,N_3969);
and U8736 (N_8736,N_5058,N_5872);
nand U8737 (N_8737,N_3403,N_5107);
and U8738 (N_8738,N_5651,N_4017);
or U8739 (N_8739,N_4483,N_5281);
nor U8740 (N_8740,N_4143,N_4978);
nor U8741 (N_8741,N_4514,N_5497);
nand U8742 (N_8742,N_3806,N_4786);
and U8743 (N_8743,N_3007,N_4306);
nor U8744 (N_8744,N_5402,N_4670);
nor U8745 (N_8745,N_5377,N_4546);
xnor U8746 (N_8746,N_5445,N_3535);
nor U8747 (N_8747,N_4842,N_4963);
or U8748 (N_8748,N_4106,N_4205);
and U8749 (N_8749,N_4651,N_3163);
and U8750 (N_8750,N_4508,N_4141);
nor U8751 (N_8751,N_4749,N_5455);
xnor U8752 (N_8752,N_5895,N_5568);
nor U8753 (N_8753,N_3797,N_4582);
or U8754 (N_8754,N_5409,N_3270);
or U8755 (N_8755,N_3877,N_3686);
nor U8756 (N_8756,N_4989,N_5050);
and U8757 (N_8757,N_5965,N_4565);
and U8758 (N_8758,N_4055,N_3053);
and U8759 (N_8759,N_4049,N_3001);
and U8760 (N_8760,N_3312,N_4979);
nor U8761 (N_8761,N_4127,N_3205);
and U8762 (N_8762,N_4077,N_5281);
or U8763 (N_8763,N_3556,N_4611);
nor U8764 (N_8764,N_4020,N_3529);
nand U8765 (N_8765,N_4236,N_4876);
or U8766 (N_8766,N_3029,N_3555);
and U8767 (N_8767,N_5545,N_3189);
nand U8768 (N_8768,N_3678,N_4176);
and U8769 (N_8769,N_4274,N_5944);
nor U8770 (N_8770,N_4085,N_5106);
or U8771 (N_8771,N_4649,N_3817);
or U8772 (N_8772,N_4722,N_5048);
xnor U8773 (N_8773,N_3022,N_5430);
or U8774 (N_8774,N_5806,N_3985);
nor U8775 (N_8775,N_3670,N_5010);
nor U8776 (N_8776,N_3043,N_5897);
xor U8777 (N_8777,N_3785,N_4339);
or U8778 (N_8778,N_3527,N_3142);
nand U8779 (N_8779,N_4708,N_4268);
nand U8780 (N_8780,N_5383,N_5730);
nor U8781 (N_8781,N_3871,N_5694);
nand U8782 (N_8782,N_4969,N_3349);
nor U8783 (N_8783,N_3439,N_4514);
or U8784 (N_8784,N_5241,N_3378);
nand U8785 (N_8785,N_4292,N_3923);
xor U8786 (N_8786,N_4779,N_3104);
or U8787 (N_8787,N_4602,N_4462);
or U8788 (N_8788,N_4223,N_3360);
and U8789 (N_8789,N_4189,N_4906);
and U8790 (N_8790,N_5416,N_5963);
or U8791 (N_8791,N_5359,N_4367);
or U8792 (N_8792,N_3538,N_5371);
nor U8793 (N_8793,N_5139,N_5266);
xor U8794 (N_8794,N_4075,N_3922);
and U8795 (N_8795,N_5414,N_4762);
and U8796 (N_8796,N_5450,N_3784);
nand U8797 (N_8797,N_4083,N_4852);
nand U8798 (N_8798,N_3088,N_3024);
nor U8799 (N_8799,N_4748,N_3314);
nor U8800 (N_8800,N_4805,N_3654);
xnor U8801 (N_8801,N_5408,N_5681);
or U8802 (N_8802,N_3371,N_4335);
nor U8803 (N_8803,N_4342,N_5688);
nor U8804 (N_8804,N_4619,N_3821);
nand U8805 (N_8805,N_4375,N_5710);
or U8806 (N_8806,N_5027,N_5164);
nand U8807 (N_8807,N_3581,N_4236);
nand U8808 (N_8808,N_5353,N_4654);
nand U8809 (N_8809,N_5449,N_4371);
nand U8810 (N_8810,N_5462,N_4665);
and U8811 (N_8811,N_4942,N_4042);
nand U8812 (N_8812,N_4127,N_3666);
nor U8813 (N_8813,N_4201,N_3808);
or U8814 (N_8814,N_4242,N_5470);
and U8815 (N_8815,N_3030,N_3653);
xor U8816 (N_8816,N_4940,N_3269);
xor U8817 (N_8817,N_4869,N_5107);
or U8818 (N_8818,N_4115,N_5947);
or U8819 (N_8819,N_3316,N_3852);
nor U8820 (N_8820,N_5548,N_3344);
nand U8821 (N_8821,N_4132,N_3572);
nand U8822 (N_8822,N_3498,N_4394);
nor U8823 (N_8823,N_4875,N_3730);
xnor U8824 (N_8824,N_3695,N_5822);
or U8825 (N_8825,N_3357,N_4500);
and U8826 (N_8826,N_4164,N_4170);
xnor U8827 (N_8827,N_3211,N_4538);
and U8828 (N_8828,N_5411,N_5685);
nor U8829 (N_8829,N_5700,N_4701);
nor U8830 (N_8830,N_5020,N_4917);
nor U8831 (N_8831,N_5729,N_5088);
and U8832 (N_8832,N_3663,N_3425);
or U8833 (N_8833,N_3815,N_3279);
nor U8834 (N_8834,N_3672,N_5445);
or U8835 (N_8835,N_3003,N_3166);
nor U8836 (N_8836,N_4051,N_5845);
nand U8837 (N_8837,N_4519,N_5934);
nand U8838 (N_8838,N_5126,N_3564);
nor U8839 (N_8839,N_4067,N_5503);
nor U8840 (N_8840,N_5274,N_3690);
and U8841 (N_8841,N_4118,N_3552);
or U8842 (N_8842,N_4997,N_3350);
nand U8843 (N_8843,N_3658,N_4869);
xnor U8844 (N_8844,N_5720,N_3715);
nand U8845 (N_8845,N_3528,N_3624);
and U8846 (N_8846,N_3776,N_3478);
or U8847 (N_8847,N_5777,N_4052);
nand U8848 (N_8848,N_5914,N_4675);
nor U8849 (N_8849,N_3656,N_4750);
nand U8850 (N_8850,N_3930,N_5357);
and U8851 (N_8851,N_3573,N_5199);
or U8852 (N_8852,N_3239,N_3125);
nor U8853 (N_8853,N_3293,N_3985);
nand U8854 (N_8854,N_3013,N_3446);
and U8855 (N_8855,N_4962,N_3653);
nand U8856 (N_8856,N_4097,N_3027);
nand U8857 (N_8857,N_5121,N_3193);
or U8858 (N_8858,N_5360,N_5626);
nor U8859 (N_8859,N_4120,N_5149);
nand U8860 (N_8860,N_3936,N_5973);
nand U8861 (N_8861,N_3291,N_5841);
nor U8862 (N_8862,N_4313,N_5348);
nor U8863 (N_8863,N_4269,N_4936);
and U8864 (N_8864,N_3728,N_4405);
nand U8865 (N_8865,N_4606,N_3825);
nor U8866 (N_8866,N_3110,N_3535);
nand U8867 (N_8867,N_4080,N_5724);
nand U8868 (N_8868,N_4552,N_4534);
nor U8869 (N_8869,N_5637,N_3959);
nand U8870 (N_8870,N_5787,N_4426);
nand U8871 (N_8871,N_3223,N_5866);
and U8872 (N_8872,N_4708,N_5456);
or U8873 (N_8873,N_5776,N_3204);
or U8874 (N_8874,N_5999,N_3186);
nand U8875 (N_8875,N_4284,N_4843);
nand U8876 (N_8876,N_3984,N_5494);
or U8877 (N_8877,N_3963,N_4843);
xnor U8878 (N_8878,N_5250,N_3944);
or U8879 (N_8879,N_5202,N_3185);
nor U8880 (N_8880,N_3746,N_4940);
and U8881 (N_8881,N_5281,N_3309);
or U8882 (N_8882,N_4105,N_5527);
nand U8883 (N_8883,N_5082,N_4100);
nor U8884 (N_8884,N_4951,N_5047);
and U8885 (N_8885,N_3577,N_4854);
nand U8886 (N_8886,N_4702,N_3659);
nand U8887 (N_8887,N_4372,N_4313);
xnor U8888 (N_8888,N_5518,N_3378);
nand U8889 (N_8889,N_5574,N_5226);
xor U8890 (N_8890,N_4072,N_3436);
xor U8891 (N_8891,N_5349,N_3599);
or U8892 (N_8892,N_4600,N_5551);
or U8893 (N_8893,N_5694,N_3457);
nor U8894 (N_8894,N_4448,N_4469);
xor U8895 (N_8895,N_3315,N_3482);
nand U8896 (N_8896,N_3039,N_4150);
nand U8897 (N_8897,N_4343,N_5253);
or U8898 (N_8898,N_3393,N_5702);
or U8899 (N_8899,N_5180,N_4485);
and U8900 (N_8900,N_3773,N_5447);
and U8901 (N_8901,N_4720,N_5179);
nand U8902 (N_8902,N_4927,N_4731);
xnor U8903 (N_8903,N_3047,N_3687);
or U8904 (N_8904,N_4336,N_4930);
and U8905 (N_8905,N_5933,N_3168);
nand U8906 (N_8906,N_4211,N_5962);
nand U8907 (N_8907,N_4776,N_4286);
nor U8908 (N_8908,N_3033,N_5378);
or U8909 (N_8909,N_3763,N_3981);
or U8910 (N_8910,N_3384,N_4785);
and U8911 (N_8911,N_5328,N_4253);
or U8912 (N_8912,N_3656,N_3766);
and U8913 (N_8913,N_3232,N_5408);
and U8914 (N_8914,N_5210,N_3424);
or U8915 (N_8915,N_5783,N_3161);
or U8916 (N_8916,N_5741,N_3725);
nor U8917 (N_8917,N_4276,N_3377);
and U8918 (N_8918,N_5685,N_5690);
nor U8919 (N_8919,N_3360,N_4732);
and U8920 (N_8920,N_4588,N_5154);
or U8921 (N_8921,N_5966,N_5964);
or U8922 (N_8922,N_4355,N_3960);
or U8923 (N_8923,N_4018,N_3008);
nor U8924 (N_8924,N_5817,N_4345);
xor U8925 (N_8925,N_5255,N_5391);
nor U8926 (N_8926,N_3497,N_5553);
and U8927 (N_8927,N_3330,N_4155);
or U8928 (N_8928,N_4927,N_4799);
xnor U8929 (N_8929,N_4356,N_3262);
and U8930 (N_8930,N_5171,N_4528);
nand U8931 (N_8931,N_4246,N_4435);
nand U8932 (N_8932,N_5030,N_5570);
nor U8933 (N_8933,N_4402,N_3903);
nand U8934 (N_8934,N_3311,N_5427);
nand U8935 (N_8935,N_5257,N_5070);
nor U8936 (N_8936,N_5766,N_5410);
nand U8937 (N_8937,N_3625,N_5241);
and U8938 (N_8938,N_3028,N_3584);
and U8939 (N_8939,N_5399,N_3542);
and U8940 (N_8940,N_4678,N_5444);
nor U8941 (N_8941,N_3220,N_3824);
and U8942 (N_8942,N_3704,N_4964);
nor U8943 (N_8943,N_4197,N_4741);
xor U8944 (N_8944,N_5664,N_5579);
and U8945 (N_8945,N_4349,N_3984);
and U8946 (N_8946,N_5679,N_5145);
xnor U8947 (N_8947,N_5127,N_5945);
xor U8948 (N_8948,N_5654,N_5818);
nor U8949 (N_8949,N_5560,N_5372);
nor U8950 (N_8950,N_5329,N_3917);
nand U8951 (N_8951,N_5759,N_4470);
or U8952 (N_8952,N_5328,N_4271);
xor U8953 (N_8953,N_3797,N_5721);
nor U8954 (N_8954,N_3080,N_3459);
and U8955 (N_8955,N_4029,N_5437);
nand U8956 (N_8956,N_4568,N_5508);
nand U8957 (N_8957,N_5792,N_4089);
nand U8958 (N_8958,N_3230,N_5982);
or U8959 (N_8959,N_3550,N_3407);
and U8960 (N_8960,N_5749,N_4598);
nand U8961 (N_8961,N_4066,N_3057);
nand U8962 (N_8962,N_3005,N_3922);
nor U8963 (N_8963,N_3122,N_4184);
or U8964 (N_8964,N_3716,N_4899);
xor U8965 (N_8965,N_5521,N_4102);
nand U8966 (N_8966,N_4226,N_5127);
xnor U8967 (N_8967,N_4492,N_5881);
and U8968 (N_8968,N_3130,N_5556);
nor U8969 (N_8969,N_4755,N_3692);
nand U8970 (N_8970,N_4515,N_4333);
and U8971 (N_8971,N_5832,N_4350);
nand U8972 (N_8972,N_5159,N_4217);
nor U8973 (N_8973,N_3834,N_5956);
or U8974 (N_8974,N_4578,N_5627);
nor U8975 (N_8975,N_4528,N_4016);
or U8976 (N_8976,N_4068,N_5321);
nor U8977 (N_8977,N_4669,N_4081);
or U8978 (N_8978,N_5519,N_3371);
and U8979 (N_8979,N_4778,N_5013);
and U8980 (N_8980,N_4162,N_3432);
or U8981 (N_8981,N_5899,N_4402);
and U8982 (N_8982,N_5172,N_3103);
xnor U8983 (N_8983,N_4959,N_5501);
nand U8984 (N_8984,N_3510,N_3964);
and U8985 (N_8985,N_3793,N_4875);
xnor U8986 (N_8986,N_5974,N_5914);
or U8987 (N_8987,N_4435,N_5878);
nand U8988 (N_8988,N_5535,N_5331);
nand U8989 (N_8989,N_4890,N_3739);
nand U8990 (N_8990,N_3613,N_5265);
or U8991 (N_8991,N_4369,N_3259);
nand U8992 (N_8992,N_5742,N_5938);
nor U8993 (N_8993,N_3180,N_4454);
xor U8994 (N_8994,N_4639,N_3106);
nand U8995 (N_8995,N_5376,N_5970);
nand U8996 (N_8996,N_4867,N_3213);
and U8997 (N_8997,N_3734,N_5211);
nand U8998 (N_8998,N_5327,N_3619);
nor U8999 (N_8999,N_4366,N_3598);
nand U9000 (N_9000,N_8240,N_8502);
nand U9001 (N_9001,N_7018,N_8136);
or U9002 (N_9002,N_7891,N_8423);
or U9003 (N_9003,N_8115,N_7400);
and U9004 (N_9004,N_6080,N_7740);
xor U9005 (N_9005,N_8865,N_8858);
nand U9006 (N_9006,N_7720,N_6721);
or U9007 (N_9007,N_7823,N_7119);
nand U9008 (N_9008,N_7775,N_8400);
nand U9009 (N_9009,N_6201,N_6778);
nor U9010 (N_9010,N_8007,N_7777);
nand U9011 (N_9011,N_6441,N_6338);
nand U9012 (N_9012,N_8834,N_6865);
nor U9013 (N_9013,N_6930,N_7630);
or U9014 (N_9014,N_7910,N_6713);
and U9015 (N_9015,N_6158,N_6000);
nand U9016 (N_9016,N_7181,N_7693);
nand U9017 (N_9017,N_8170,N_8134);
or U9018 (N_9018,N_8767,N_6983);
or U9019 (N_9019,N_8307,N_7407);
nand U9020 (N_9020,N_6092,N_7277);
or U9021 (N_9021,N_7444,N_7873);
nand U9022 (N_9022,N_8605,N_8758);
nand U9023 (N_9023,N_6958,N_8390);
nor U9024 (N_9024,N_7782,N_6732);
nor U9025 (N_9025,N_7022,N_8312);
or U9026 (N_9026,N_7074,N_7129);
or U9027 (N_9027,N_7058,N_8025);
nor U9028 (N_9028,N_8002,N_6844);
nand U9029 (N_9029,N_7763,N_7009);
nor U9030 (N_9030,N_6668,N_8492);
or U9031 (N_9031,N_6645,N_7028);
xor U9032 (N_9032,N_7158,N_8925);
or U9033 (N_9033,N_7362,N_7170);
or U9034 (N_9034,N_8268,N_7858);
and U9035 (N_9035,N_7324,N_6527);
and U9036 (N_9036,N_6119,N_8163);
or U9037 (N_9037,N_6822,N_7943);
xnor U9038 (N_9038,N_7088,N_6138);
and U9039 (N_9039,N_6323,N_6973);
xnor U9040 (N_9040,N_7530,N_8071);
xnor U9041 (N_9041,N_6387,N_6694);
or U9042 (N_9042,N_6188,N_7801);
nor U9043 (N_9043,N_8033,N_6041);
nor U9044 (N_9044,N_7653,N_8179);
nand U9045 (N_9045,N_8284,N_8777);
xnor U9046 (N_9046,N_7734,N_8577);
xor U9047 (N_9047,N_6141,N_6061);
nand U9048 (N_9048,N_6505,N_8408);
or U9049 (N_9049,N_7112,N_6510);
nor U9050 (N_9050,N_6334,N_8957);
nand U9051 (N_9051,N_6813,N_7625);
and U9052 (N_9052,N_7041,N_7645);
and U9053 (N_9053,N_6969,N_7947);
or U9054 (N_9054,N_6491,N_8806);
nor U9055 (N_9055,N_7526,N_8624);
nand U9056 (N_9056,N_7266,N_8601);
or U9057 (N_9057,N_6295,N_8412);
and U9058 (N_9058,N_8874,N_6727);
nor U9059 (N_9059,N_6555,N_7717);
or U9060 (N_9060,N_7748,N_6465);
or U9061 (N_9061,N_7854,N_6917);
xnor U9062 (N_9062,N_6619,N_7497);
and U9063 (N_9063,N_6600,N_7410);
and U9064 (N_9064,N_7118,N_8885);
nor U9065 (N_9065,N_7884,N_8964);
and U9066 (N_9066,N_6927,N_7273);
xor U9067 (N_9067,N_6557,N_7002);
nand U9068 (N_9068,N_6671,N_6972);
or U9069 (N_9069,N_6664,N_7728);
or U9070 (N_9070,N_6082,N_7632);
or U9071 (N_9071,N_6234,N_7951);
nand U9072 (N_9072,N_8581,N_7219);
and U9073 (N_9073,N_6956,N_7014);
and U9074 (N_9074,N_8591,N_7877);
and U9075 (N_9075,N_7974,N_7121);
or U9076 (N_9076,N_8528,N_8039);
nor U9077 (N_9077,N_6352,N_8602);
or U9078 (N_9078,N_7606,N_7244);
and U9079 (N_9079,N_6626,N_6752);
and U9080 (N_9080,N_6538,N_8667);
nor U9081 (N_9081,N_7930,N_7867);
and U9082 (N_9082,N_6533,N_8373);
nor U9083 (N_9083,N_7200,N_8419);
and U9084 (N_9084,N_7965,N_6477);
and U9085 (N_9085,N_8882,N_6076);
nand U9086 (N_9086,N_8856,N_6634);
nor U9087 (N_9087,N_6405,N_6891);
or U9088 (N_9088,N_6427,N_7189);
nor U9089 (N_9089,N_6191,N_7684);
or U9090 (N_9090,N_8529,N_6679);
nor U9091 (N_9091,N_8967,N_7475);
nand U9092 (N_9092,N_6209,N_8036);
and U9093 (N_9093,N_6877,N_6878);
nor U9094 (N_9094,N_8918,N_7073);
nor U9095 (N_9095,N_6616,N_7150);
or U9096 (N_9096,N_6094,N_6860);
nand U9097 (N_9097,N_7706,N_7817);
or U9098 (N_9098,N_8143,N_8366);
and U9099 (N_9099,N_6636,N_7286);
and U9100 (N_9100,N_7998,N_6202);
xnor U9101 (N_9101,N_7205,N_8573);
and U9102 (N_9102,N_8593,N_7992);
nand U9103 (N_9103,N_7233,N_8812);
nor U9104 (N_9104,N_7185,N_8067);
or U9105 (N_9105,N_8424,N_7633);
and U9106 (N_9106,N_6319,N_7667);
or U9107 (N_9107,N_6605,N_6269);
or U9108 (N_9108,N_7264,N_7476);
and U9109 (N_9109,N_8384,N_7703);
nor U9110 (N_9110,N_8642,N_8098);
nand U9111 (N_9111,N_7599,N_8206);
nor U9112 (N_9112,N_6929,N_7924);
or U9113 (N_9113,N_6750,N_7870);
or U9114 (N_9114,N_8316,N_6419);
or U9115 (N_9115,N_7689,N_8130);
and U9116 (N_9116,N_7203,N_8364);
or U9117 (N_9117,N_8140,N_8022);
or U9118 (N_9118,N_8448,N_8970);
or U9119 (N_9119,N_7934,N_7345);
and U9120 (N_9120,N_6838,N_8301);
and U9121 (N_9121,N_8550,N_6475);
nor U9122 (N_9122,N_6134,N_7287);
nand U9123 (N_9123,N_7169,N_8173);
xnor U9124 (N_9124,N_7876,N_6374);
nor U9125 (N_9125,N_7591,N_8907);
or U9126 (N_9126,N_6585,N_8501);
nor U9127 (N_9127,N_6013,N_8505);
and U9128 (N_9128,N_7566,N_7695);
nand U9129 (N_9129,N_6697,N_8676);
and U9130 (N_9130,N_8458,N_8406);
nand U9131 (N_9131,N_6857,N_7552);
nand U9132 (N_9132,N_8138,N_6971);
nand U9133 (N_9133,N_6086,N_6122);
xor U9134 (N_9134,N_6035,N_7839);
nor U9135 (N_9135,N_8447,N_8056);
and U9136 (N_9136,N_6689,N_8841);
and U9137 (N_9137,N_7956,N_8347);
nand U9138 (N_9138,N_6712,N_8641);
and U9139 (N_9139,N_7191,N_7524);
nand U9140 (N_9140,N_7096,N_6568);
or U9141 (N_9141,N_7253,N_7042);
nand U9142 (N_9142,N_6455,N_6582);
and U9143 (N_9143,N_6839,N_7749);
and U9144 (N_9144,N_6536,N_8122);
nor U9145 (N_9145,N_7292,N_7802);
or U9146 (N_9146,N_6793,N_8818);
nor U9147 (N_9147,N_7837,N_8768);
and U9148 (N_9148,N_8234,N_7791);
nor U9149 (N_9149,N_6925,N_8220);
and U9150 (N_9150,N_6445,N_6125);
or U9151 (N_9151,N_7577,N_6272);
xnor U9152 (N_9152,N_8755,N_7060);
nand U9153 (N_9153,N_6322,N_8973);
and U9154 (N_9154,N_7289,N_7384);
or U9155 (N_9155,N_8819,N_7386);
nand U9156 (N_9156,N_7739,N_7729);
nor U9157 (N_9157,N_7565,N_6836);
or U9158 (N_9158,N_6054,N_6719);
nand U9159 (N_9159,N_6497,N_8315);
and U9160 (N_9160,N_6494,N_7994);
nand U9161 (N_9161,N_8992,N_7932);
nor U9162 (N_9162,N_8042,N_6699);
nand U9163 (N_9163,N_6753,N_8625);
and U9164 (N_9164,N_7710,N_6489);
xnor U9165 (N_9165,N_8280,N_6566);
nor U9166 (N_9166,N_7660,N_6556);
nand U9167 (N_9167,N_6299,N_7117);
and U9168 (N_9168,N_8653,N_7855);
nand U9169 (N_9169,N_6402,N_7807);
nand U9170 (N_9170,N_6896,N_8461);
and U9171 (N_9171,N_8432,N_8146);
nor U9172 (N_9172,N_6591,N_6456);
or U9173 (N_9173,N_8935,N_6296);
nor U9174 (N_9174,N_7333,N_8254);
nor U9175 (N_9175,N_6792,N_7545);
xnor U9176 (N_9176,N_7414,N_8333);
or U9177 (N_9177,N_8431,N_7025);
xor U9178 (N_9178,N_6314,N_8728);
or U9179 (N_9179,N_7366,N_7767);
and U9180 (N_9180,N_8621,N_7351);
nor U9181 (N_9181,N_8020,N_8380);
xor U9182 (N_9182,N_8521,N_7307);
and U9183 (N_9183,N_7019,N_8200);
and U9184 (N_9184,N_6245,N_6084);
or U9185 (N_9185,N_6207,N_8389);
or U9186 (N_9186,N_7367,N_7923);
nand U9187 (N_9187,N_8449,N_8889);
and U9188 (N_9188,N_7111,N_7109);
nor U9189 (N_9189,N_6143,N_7243);
xnor U9190 (N_9190,N_7600,N_8799);
and U9191 (N_9191,N_6598,N_8162);
xor U9192 (N_9192,N_6607,N_8207);
and U9193 (N_9193,N_6415,N_7935);
and U9194 (N_9194,N_6170,N_6867);
nor U9195 (N_9195,N_8804,N_8994);
nand U9196 (N_9196,N_8786,N_7655);
xnor U9197 (N_9197,N_7370,N_6227);
and U9198 (N_9198,N_7852,N_6952);
nand U9199 (N_9199,N_6248,N_8244);
or U9200 (N_9200,N_8990,N_7179);
and U9201 (N_9201,N_7776,N_8356);
nor U9202 (N_9202,N_8944,N_6832);
or U9203 (N_9203,N_8672,N_6757);
or U9204 (N_9204,N_6666,N_7670);
or U9205 (N_9205,N_8187,N_6931);
nor U9206 (N_9206,N_7869,N_6263);
or U9207 (N_9207,N_6611,N_8250);
and U9208 (N_9208,N_6660,N_6683);
nand U9209 (N_9209,N_8982,N_8780);
and U9210 (N_9210,N_8375,N_8582);
nand U9211 (N_9211,N_8091,N_8879);
nand U9212 (N_9212,N_7824,N_8464);
nor U9213 (N_9213,N_8494,N_6926);
nand U9214 (N_9214,N_7328,N_7644);
or U9215 (N_9215,N_6604,N_8741);
and U9216 (N_9216,N_8063,N_7330);
nand U9217 (N_9217,N_8231,N_6412);
and U9218 (N_9218,N_6534,N_8747);
nand U9219 (N_9219,N_6071,N_6022);
nand U9220 (N_9220,N_7172,N_6121);
nor U9221 (N_9221,N_6291,N_7385);
nand U9222 (N_9222,N_8855,N_7601);
nand U9223 (N_9223,N_6550,N_8185);
nor U9224 (N_9224,N_6286,N_6883);
nand U9225 (N_9225,N_6389,N_8626);
nand U9226 (N_9226,N_6223,N_8714);
and U9227 (N_9227,N_6488,N_7135);
nand U9228 (N_9228,N_8236,N_8241);
nor U9229 (N_9229,N_6253,N_7394);
and U9230 (N_9230,N_6769,N_8842);
or U9231 (N_9231,N_6663,N_6336);
or U9232 (N_9232,N_7482,N_6975);
nor U9233 (N_9233,N_7318,N_8409);
nand U9234 (N_9234,N_8168,N_7144);
or U9235 (N_9235,N_8319,N_6725);
or U9236 (N_9236,N_7418,N_6482);
nor U9237 (N_9237,N_7469,N_6995);
or U9238 (N_9238,N_7602,N_6171);
or U9239 (N_9239,N_8608,N_8652);
or U9240 (N_9240,N_6365,N_7449);
nor U9241 (N_9241,N_8727,N_8807);
nand U9242 (N_9242,N_8435,N_8734);
nand U9243 (N_9243,N_8705,N_6770);
nor U9244 (N_9244,N_6357,N_7723);
and U9245 (N_9245,N_7509,N_8515);
and U9246 (N_9246,N_7881,N_8800);
or U9247 (N_9247,N_7340,N_6820);
nor U9248 (N_9248,N_8868,N_7716);
nand U9249 (N_9249,N_8015,N_8480);
nand U9250 (N_9250,N_6474,N_6045);
and U9251 (N_9251,N_7933,N_6326);
or U9252 (N_9252,N_8945,N_8579);
nand U9253 (N_9253,N_8508,N_8607);
nand U9254 (N_9254,N_8884,N_8118);
nand U9255 (N_9255,N_7850,N_6216);
nor U9256 (N_9256,N_6083,N_6088);
or U9257 (N_9257,N_7473,N_6690);
and U9258 (N_9258,N_8346,N_7461);
or U9259 (N_9259,N_8846,N_6457);
nand U9260 (N_9260,N_8451,N_8597);
or U9261 (N_9261,N_8142,N_6351);
and U9262 (N_9262,N_7308,N_7747);
or U9263 (N_9263,N_6051,N_7033);
and U9264 (N_9264,N_6936,N_7215);
nor U9265 (N_9265,N_6833,N_6243);
nand U9266 (N_9266,N_7982,N_6341);
nand U9267 (N_9267,N_7561,N_7329);
or U9268 (N_9268,N_8829,N_8989);
or U9269 (N_9269,N_6362,N_7211);
and U9270 (N_9270,N_6939,N_7420);
xnor U9271 (N_9271,N_7495,N_7288);
nand U9272 (N_9272,N_7553,N_7709);
nand U9273 (N_9273,N_7458,N_6458);
and U9274 (N_9274,N_7113,N_8956);
nor U9275 (N_9275,N_8857,N_8701);
or U9276 (N_9276,N_7132,N_6775);
and U9277 (N_9277,N_6224,N_7976);
and U9278 (N_9278,N_8271,N_8993);
and U9279 (N_9279,N_8564,N_6882);
nor U9280 (N_9280,N_7166,N_7589);
nand U9281 (N_9281,N_8255,N_7068);
nand U9282 (N_9282,N_8554,N_7023);
nor U9283 (N_9283,N_6642,N_8756);
and U9284 (N_9284,N_7276,N_7434);
xor U9285 (N_9285,N_6578,N_7293);
or U9286 (N_9286,N_6379,N_6019);
xor U9287 (N_9287,N_8282,N_6916);
and U9288 (N_9288,N_8239,N_8736);
or U9289 (N_9289,N_8825,N_7492);
or U9290 (N_9290,N_8078,N_6359);
nor U9291 (N_9291,N_8403,N_7522);
or U9292 (N_9292,N_7339,N_7477);
and U9293 (N_9293,N_7234,N_6961);
and U9294 (N_9294,N_7503,N_6677);
and U9295 (N_9295,N_6440,N_8444);
nand U9296 (N_9296,N_7206,N_6064);
nand U9297 (N_9297,N_8568,N_8272);
and U9298 (N_9298,N_7527,N_8222);
nor U9299 (N_9299,N_6115,N_7236);
or U9300 (N_9300,N_6347,N_7409);
nand U9301 (N_9301,N_6811,N_6547);
nand U9302 (N_9302,N_7387,N_7905);
xnor U9303 (N_9303,N_8835,N_8471);
nor U9304 (N_9304,N_8126,N_6992);
nor U9305 (N_9305,N_8183,N_6580);
or U9306 (N_9306,N_8097,N_8520);
xnor U9307 (N_9307,N_7498,N_7610);
xor U9308 (N_9308,N_8668,N_7618);
or U9309 (N_9309,N_8177,N_7505);
and U9310 (N_9310,N_7569,N_8981);
or U9311 (N_9311,N_7779,N_8571);
nand U9312 (N_9312,N_7608,N_7224);
or U9313 (N_9313,N_7911,N_6260);
or U9314 (N_9314,N_8311,N_6986);
nand U9315 (N_9315,N_7262,N_8455);
or U9316 (N_9316,N_6530,N_8805);
or U9317 (N_9317,N_8659,N_8960);
xor U9318 (N_9318,N_6782,N_8947);
nand U9319 (N_9319,N_6633,N_8425);
nand U9320 (N_9320,N_7299,N_7195);
and U9321 (N_9321,N_7928,N_6430);
and U9322 (N_9322,N_7658,N_8649);
and U9323 (N_9323,N_7356,N_7275);
xor U9324 (N_9324,N_6553,N_6169);
nand U9325 (N_9325,N_6442,N_6340);
nor U9326 (N_9326,N_6845,N_6764);
nand U9327 (N_9327,N_7742,N_7134);
nor U9328 (N_9328,N_7280,N_6384);
and U9329 (N_9329,N_7668,N_7327);
and U9330 (N_9330,N_6066,N_6552);
and U9331 (N_9331,N_7471,N_6197);
or U9332 (N_9332,N_7395,N_8106);
nor U9333 (N_9333,N_7937,N_7652);
or U9334 (N_9334,N_8418,N_8644);
nand U9335 (N_9335,N_6342,N_6572);
nand U9336 (N_9336,N_8260,N_7666);
nor U9337 (N_9337,N_6966,N_7103);
nand U9338 (N_9338,N_7972,N_6237);
nor U9339 (N_9339,N_7188,N_8584);
nand U9340 (N_9340,N_6797,N_8703);
or U9341 (N_9341,N_7325,N_6674);
and U9342 (N_9342,N_8490,N_7548);
and U9343 (N_9343,N_7744,N_7916);
nand U9344 (N_9344,N_6065,N_8779);
and U9345 (N_9345,N_8149,N_8660);
or U9346 (N_9346,N_7550,N_6062);
and U9347 (N_9347,N_8420,N_8764);
or U9348 (N_9348,N_8083,N_7764);
xnor U9349 (N_9349,N_8578,N_6696);
nor U9350 (N_9350,N_8365,N_6250);
or U9351 (N_9351,N_8229,N_7541);
nand U9352 (N_9352,N_6354,N_6543);
nand U9353 (N_9353,N_6606,N_8295);
nor U9354 (N_9354,N_6609,N_8395);
or U9355 (N_9355,N_7013,N_7544);
nand U9356 (N_9356,N_6398,N_6371);
or U9357 (N_9357,N_6308,N_8481);
nor U9358 (N_9358,N_8986,N_7460);
nor U9359 (N_9359,N_7603,N_6004);
nor U9360 (N_9360,N_6337,N_6754);
or U9361 (N_9361,N_7525,N_8332);
or U9362 (N_9362,N_7004,N_6853);
xnor U9363 (N_9363,N_6964,N_6922);
nor U9364 (N_9364,N_6462,N_8038);
nand U9365 (N_9365,N_8911,N_7297);
and U9366 (N_9366,N_8084,N_8963);
and U9367 (N_9367,N_6344,N_6498);
xor U9368 (N_9368,N_8833,N_7153);
nor U9369 (N_9369,N_7057,N_7353);
xor U9370 (N_9370,N_6998,N_6020);
xor U9371 (N_9371,N_8585,N_6638);
or U9372 (N_9372,N_8853,N_7398);
or U9373 (N_9373,N_6404,N_7361);
and U9374 (N_9374,N_7183,N_6739);
nor U9375 (N_9375,N_8849,N_6861);
and U9376 (N_9376,N_7892,N_8987);
or U9377 (N_9377,N_8158,N_6343);
or U9378 (N_9378,N_6040,N_8771);
and U9379 (N_9379,N_7897,N_6241);
or U9380 (N_9380,N_7197,N_6603);
and U9381 (N_9381,N_6548,N_6394);
nand U9382 (N_9382,N_7040,N_8298);
nand U9383 (N_9383,N_7510,N_7048);
or U9384 (N_9384,N_8186,N_6864);
nand U9385 (N_9385,N_7246,N_8631);
nand U9386 (N_9386,N_8344,N_6274);
or U9387 (N_9387,N_8309,N_6070);
and U9388 (N_9388,N_7194,N_8479);
nand U9389 (N_9389,N_6508,N_8544);
or U9390 (N_9390,N_8367,N_8402);
nor U9391 (N_9391,N_7470,N_7904);
nand U9392 (N_9392,N_6742,N_8802);
or U9393 (N_9393,N_6843,N_6225);
or U9394 (N_9394,N_7065,N_7719);
and U9395 (N_9395,N_6196,N_6933);
nor U9396 (N_9396,N_7316,N_6819);
nor U9397 (N_9397,N_8830,N_8252);
or U9398 (N_9398,N_8297,N_6108);
nand U9399 (N_9399,N_8937,N_7388);
and U9400 (N_9400,N_8718,N_6109);
and U9401 (N_9401,N_8700,N_8283);
nor U9402 (N_9402,N_7549,N_8167);
nor U9403 (N_9403,N_8066,N_8870);
nand U9404 (N_9404,N_6174,N_6252);
nor U9405 (N_9405,N_6963,N_8751);
nand U9406 (N_9406,N_6211,N_6277);
or U9407 (N_9407,N_8349,N_7752);
and U9408 (N_9408,N_7543,N_8748);
or U9409 (N_9409,N_7402,N_6385);
and U9410 (N_9410,N_8513,N_7399);
nor U9411 (N_9411,N_8662,N_7771);
nand U9412 (N_9412,N_7826,N_7788);
nor U9413 (N_9413,N_6399,N_7936);
or U9414 (N_9414,N_8536,N_7439);
or U9415 (N_9415,N_7741,N_7502);
or U9416 (N_9416,N_8509,N_8157);
nand U9417 (N_9417,N_7862,N_6266);
nand U9418 (N_9418,N_6943,N_8417);
xor U9419 (N_9419,N_8489,N_8345);
nor U9420 (N_9420,N_7560,N_8029);
nand U9421 (N_9421,N_7092,N_8090);
xnor U9422 (N_9422,N_8230,N_8046);
xnor U9423 (N_9423,N_8915,N_7404);
nand U9424 (N_9424,N_7975,N_7347);
and U9425 (N_9425,N_6281,N_7240);
and U9426 (N_9426,N_6029,N_8011);
and U9427 (N_9427,N_7152,N_8991);
and U9428 (N_9428,N_6574,N_8620);
and U9429 (N_9429,N_8511,N_6329);
nand U9430 (N_9430,N_6400,N_8691);
nand U9431 (N_9431,N_7466,N_6653);
or U9432 (N_9432,N_7301,N_8196);
nand U9433 (N_9433,N_7769,N_6849);
xor U9434 (N_9434,N_8306,N_8933);
or U9435 (N_9435,N_6651,N_6976);
or U9436 (N_9436,N_7130,N_8160);
nor U9437 (N_9437,N_8000,N_7563);
nor U9438 (N_9438,N_7713,N_7416);
nand U9439 (N_9439,N_7320,N_7690);
nor U9440 (N_9440,N_8276,N_6060);
or U9441 (N_9441,N_7459,N_7762);
xor U9442 (N_9442,N_8460,N_7629);
and U9443 (N_9443,N_8010,N_7371);
or U9444 (N_9444,N_7627,N_8437);
or U9445 (N_9445,N_8617,N_7467);
or U9446 (N_9446,N_7151,N_6788);
xor U9447 (N_9447,N_6009,N_7016);
nor U9448 (N_9448,N_7506,N_7496);
or U9449 (N_9449,N_8761,N_8338);
and U9450 (N_9450,N_6688,N_8517);
nor U9451 (N_9451,N_8934,N_6847);
and U9452 (N_9452,N_6230,N_8685);
and U9453 (N_9453,N_8815,N_8181);
and U9454 (N_9454,N_7047,N_6144);
and U9455 (N_9455,N_8145,N_6625);
nor U9456 (N_9456,N_8687,N_7437);
or U9457 (N_9457,N_6814,N_7746);
or U9458 (N_9458,N_7091,N_7305);
and U9459 (N_9459,N_6424,N_8916);
nor U9460 (N_9460,N_6672,N_6306);
nand U9461 (N_9461,N_8760,N_6622);
nand U9462 (N_9462,N_8796,N_8221);
nand U9463 (N_9463,N_8996,N_7484);
xnor U9464 (N_9464,N_7222,N_8101);
nor U9465 (N_9465,N_8671,N_8401);
nor U9466 (N_9466,N_7614,N_8488);
nand U9467 (N_9467,N_6073,N_6686);
and U9468 (N_9468,N_6661,N_6873);
nor U9469 (N_9469,N_6081,N_7705);
nand U9470 (N_9470,N_8131,N_6863);
nand U9471 (N_9471,N_7082,N_8811);
and U9472 (N_9472,N_7411,N_8600);
nor U9473 (N_9473,N_7210,N_7774);
and U9474 (N_9474,N_8358,N_6214);
and U9475 (N_9475,N_7355,N_7207);
and U9476 (N_9476,N_8599,N_7647);
nand U9477 (N_9477,N_7232,N_6231);
nor U9478 (N_9478,N_6087,N_7008);
or U9479 (N_9479,N_8637,N_7489);
or U9480 (N_9480,N_8698,N_8051);
or U9481 (N_9481,N_7587,N_6413);
or U9482 (N_9482,N_8785,N_6588);
and U9483 (N_9483,N_7906,N_7472);
and U9484 (N_9484,N_7265,N_7260);
nand U9485 (N_9485,N_7036,N_7405);
xnor U9486 (N_9486,N_7512,N_6648);
nor U9487 (N_9487,N_6584,N_7798);
or U9488 (N_9488,N_7805,N_6561);
or U9489 (N_9489,N_8968,N_8580);
and U9490 (N_9490,N_7570,N_7303);
nor U9491 (N_9491,N_7793,N_7350);
or U9492 (N_9492,N_8452,N_7612);
nand U9493 (N_9493,N_6485,N_7268);
nor U9494 (N_9494,N_6748,N_7607);
nand U9495 (N_9495,N_7256,N_7745);
and U9496 (N_9496,N_8863,N_7687);
and U9497 (N_9497,N_7247,N_7958);
and U9498 (N_9498,N_6236,N_6478);
and U9499 (N_9499,N_7201,N_7754);
nor U9500 (N_9500,N_6830,N_8095);
or U9501 (N_9501,N_7733,N_7397);
nand U9502 (N_9502,N_6514,N_8150);
nand U9503 (N_9503,N_8891,N_7086);
nand U9504 (N_9504,N_7491,N_6831);
or U9505 (N_9505,N_7819,N_6545);
nand U9506 (N_9506,N_6738,N_8318);
or U9507 (N_9507,N_8661,N_6273);
xnor U9508 (N_9508,N_7619,N_7160);
and U9509 (N_9509,N_8049,N_6678);
xor U9510 (N_9510,N_6573,N_8474);
and U9511 (N_9511,N_7961,N_7980);
and U9512 (N_9512,N_8790,N_8931);
nand U9513 (N_9513,N_7372,N_7863);
or U9514 (N_9514,N_7248,N_8226);
or U9515 (N_9515,N_7927,N_6152);
nor U9516 (N_9516,N_7343,N_7828);
or U9517 (N_9517,N_6554,N_6518);
or U9518 (N_9518,N_6637,N_8330);
or U9519 (N_9519,N_7392,N_7504);
or U9520 (N_9520,N_8946,N_6390);
or U9521 (N_9521,N_7750,N_8610);
or U9522 (N_9522,N_7564,N_8077);
and U9523 (N_9523,N_7954,N_8279);
nand U9524 (N_9524,N_7620,N_6294);
and U9525 (N_9525,N_7722,N_7225);
nor U9526 (N_9526,N_7836,N_6452);
and U9527 (N_9527,N_6284,N_7657);
or U9528 (N_9528,N_8040,N_8657);
nor U9529 (N_9529,N_7783,N_8438);
nor U9530 (N_9530,N_8299,N_6249);
nor U9531 (N_9531,N_8331,N_8125);
or U9532 (N_9532,N_6136,N_7124);
nor U9533 (N_9533,N_6991,N_6150);
xor U9534 (N_9534,N_6640,N_7230);
and U9535 (N_9535,N_7966,N_6382);
nor U9536 (N_9536,N_8430,N_8909);
and U9537 (N_9537,N_7611,N_8053);
nor U9538 (N_9538,N_8476,N_8538);
nor U9539 (N_9539,N_7737,N_6195);
and U9540 (N_9540,N_6002,N_8245);
nand U9541 (N_9541,N_7841,N_7173);
and U9542 (N_9542,N_8753,N_6068);
nor U9543 (N_9543,N_7669,N_7202);
nor U9544 (N_9544,N_6407,N_7698);
or U9545 (N_9545,N_7708,N_6037);
nand U9546 (N_9546,N_7914,N_8439);
nand U9547 (N_9547,N_8072,N_6282);
nor U9548 (N_9548,N_8171,N_6047);
nand U9549 (N_9549,N_6923,N_7613);
nand U9550 (N_9550,N_6824,N_6967);
nor U9551 (N_9551,N_6057,N_8523);
or U9552 (N_9552,N_6470,N_7797);
nand U9553 (N_9553,N_7665,N_7164);
nand U9554 (N_9554,N_7080,N_8243);
nand U9555 (N_9555,N_8035,N_6148);
and U9556 (N_9556,N_8343,N_8281);
and U9557 (N_9557,N_6624,N_7597);
nor U9558 (N_9558,N_7396,N_7533);
nor U9559 (N_9559,N_6984,N_6851);
nand U9560 (N_9560,N_7269,N_6300);
nand U9561 (N_9561,N_8251,N_7237);
nor U9562 (N_9562,N_7486,N_7678);
nand U9563 (N_9563,N_8518,N_6397);
or U9564 (N_9564,N_8547,N_6189);
and U9565 (N_9565,N_6386,N_6669);
nor U9566 (N_9566,N_6466,N_8305);
nand U9567 (N_9567,N_7365,N_6244);
or U9568 (N_9568,N_8754,N_6215);
and U9569 (N_9569,N_6043,N_8706);
and U9570 (N_9570,N_8636,N_6024);
nor U9571 (N_9571,N_8496,N_8218);
or U9572 (N_9572,N_7738,N_8522);
nor U9573 (N_9573,N_8396,N_7856);
nand U9574 (N_9574,N_8503,N_8724);
or U9575 (N_9575,N_7809,N_6515);
xor U9576 (N_9576,N_7860,N_8596);
and U9577 (N_9577,N_6521,N_8546);
and U9578 (N_9578,N_8456,N_6618);
xor U9579 (N_9579,N_6126,N_6546);
xnor U9580 (N_9580,N_7309,N_7794);
or U9581 (N_9581,N_7813,N_6565);
and U9582 (N_9582,N_7377,N_6178);
xor U9583 (N_9583,N_8675,N_8765);
xnor U9584 (N_9584,N_6483,N_6114);
or U9585 (N_9585,N_6210,N_8827);
xor U9586 (N_9586,N_6502,N_8740);
or U9587 (N_9587,N_7701,N_6693);
xor U9588 (N_9588,N_7845,N_7926);
and U9589 (N_9589,N_7635,N_8495);
nor U9590 (N_9590,N_8939,N_8725);
nor U9591 (N_9591,N_6181,N_6781);
nor U9592 (N_9592,N_7226,N_6828);
nor U9593 (N_9593,N_7726,N_7948);
nor U9594 (N_9594,N_7582,N_6799);
nand U9595 (N_9595,N_6011,N_8211);
and U9596 (N_9596,N_8936,N_8735);
nor U9597 (N_9597,N_7284,N_7790);
nand U9598 (N_9598,N_7326,N_6460);
nor U9599 (N_9599,N_8559,N_6228);
nand U9600 (N_9600,N_8152,N_6434);
or U9601 (N_9601,N_8587,N_7623);
nor U9602 (N_9602,N_7663,N_8290);
or U9603 (N_9603,N_6639,N_8789);
nor U9604 (N_9604,N_6380,N_6194);
nand U9605 (N_9605,N_8616,N_7430);
or U9606 (N_9606,N_7148,N_6190);
or U9607 (N_9607,N_6912,N_6476);
nor U9608 (N_9608,N_7214,N_7515);
nand U9609 (N_9609,N_8658,N_7429);
nand U9610 (N_9610,N_6246,N_6461);
and U9611 (N_9611,N_8782,N_8368);
nand U9612 (N_9612,N_7945,N_7922);
and U9613 (N_9613,N_6238,N_6451);
nor U9614 (N_9614,N_8781,N_7304);
or U9615 (N_9615,N_8440,N_8656);
or U9616 (N_9616,N_8962,N_8826);
and U9617 (N_9617,N_8711,N_7700);
and U9618 (N_9618,N_7006,N_8708);
and U9619 (N_9619,N_8560,N_8638);
xor U9620 (N_9620,N_8362,N_8822);
and U9621 (N_9621,N_6056,N_7517);
nor U9622 (N_9622,N_6911,N_8681);
nor U9623 (N_9623,N_8598,N_7571);
nor U9624 (N_9624,N_7531,N_7358);
and U9625 (N_9625,N_8924,N_8021);
or U9626 (N_9626,N_6420,N_7990);
or U9627 (N_9627,N_6999,N_6028);
xor U9628 (N_9628,N_6501,N_7108);
nand U9629 (N_9629,N_6620,N_7886);
nor U9630 (N_9630,N_6172,N_8139);
or U9631 (N_9631,N_7131,N_7382);
and U9632 (N_9632,N_7037,N_8633);
nor U9633 (N_9633,N_7714,N_7743);
and U9634 (N_9634,N_6876,N_6468);
and U9635 (N_9635,N_6472,N_8861);
nand U9636 (N_9636,N_6920,N_7331);
xor U9637 (N_9637,N_8096,N_8843);
or U9638 (N_9638,N_8467,N_6111);
and U9639 (N_9639,N_8859,N_7490);
xnor U9640 (N_9640,N_7692,N_8974);
nand U9641 (N_9641,N_8064,N_8809);
or U9642 (N_9642,N_6898,N_7894);
or U9643 (N_9643,N_7513,N_6575);
and U9644 (N_9644,N_7997,N_7063);
xnor U9645 (N_9645,N_8902,N_7454);
or U9646 (N_9646,N_8942,N_6220);
nand U9647 (N_9647,N_8429,N_8845);
nand U9648 (N_9648,N_7448,N_7196);
nor U9649 (N_9649,N_6356,N_6840);
xnor U9650 (N_9650,N_7271,N_6425);
nand U9651 (N_9651,N_8575,N_6889);
xnor U9652 (N_9652,N_7431,N_7554);
nor U9653 (N_9653,N_6628,N_6417);
nor U9654 (N_9654,N_6325,N_6776);
or U9655 (N_9655,N_7731,N_8640);
and U9656 (N_9656,N_8959,N_6212);
or U9657 (N_9657,N_6315,N_6367);
and U9658 (N_9658,N_6980,N_8537);
and U9659 (N_9659,N_8385,N_7508);
or U9660 (N_9660,N_6747,N_6265);
or U9661 (N_9661,N_8159,N_7908);
nand U9662 (N_9662,N_8762,N_6509);
or U9663 (N_9663,N_7622,N_8562);
or U9664 (N_9664,N_8533,N_6676);
nor U9665 (N_9665,N_6506,N_7536);
or U9666 (N_9666,N_7302,N_6304);
nor U9667 (N_9667,N_8112,N_8697);
or U9668 (N_9668,N_8732,N_8632);
or U9669 (N_9669,N_8277,N_7501);
and U9670 (N_9670,N_8905,N_7507);
and U9671 (N_9671,N_8377,N_7178);
and U9672 (N_9672,N_6469,N_7278);
nor U9673 (N_9673,N_8073,N_8985);
nand U9674 (N_9674,N_8198,N_7168);
nor U9675 (N_9675,N_7919,N_6285);
and U9676 (N_9676,N_6801,N_8952);
and U9677 (N_9677,N_6499,N_6151);
and U9678 (N_9678,N_7311,N_6007);
or U9679 (N_9679,N_6859,N_6751);
nor U9680 (N_9680,N_6540,N_8374);
nor U9681 (N_9681,N_6446,N_6708);
nor U9682 (N_9682,N_6368,N_7156);
and U9683 (N_9683,N_8086,N_6256);
and U9684 (N_9684,N_6948,N_8137);
and U9685 (N_9685,N_8264,N_7557);
and U9686 (N_9686,N_7115,N_6522);
nor U9687 (N_9687,N_8583,N_7039);
nand U9688 (N_9688,N_8721,N_7986);
nand U9689 (N_9689,N_6892,N_6532);
or U9690 (N_9690,N_7772,N_8940);
xor U9691 (N_9691,N_6480,N_8752);
and U9692 (N_9692,N_8526,N_6159);
and U9693 (N_9693,N_8746,N_6773);
nor U9694 (N_9694,N_7252,N_7962);
or U9695 (N_9695,N_6067,N_6104);
xnor U9696 (N_9696,N_8124,N_6724);
and U9697 (N_9697,N_7518,N_8174);
nor U9698 (N_9698,N_7251,N_8715);
nor U9699 (N_9699,N_8387,N_6481);
nor U9700 (N_9700,N_8770,N_8908);
or U9701 (N_9701,N_8238,N_8766);
nand U9702 (N_9702,N_7055,N_6353);
or U9703 (N_9703,N_6915,N_8216);
nor U9704 (N_9704,N_8965,N_7753);
nor U9705 (N_9705,N_6383,N_6077);
nand U9706 (N_9706,N_6133,N_6960);
nand U9707 (N_9707,N_7021,N_6528);
and U9708 (N_9708,N_6180,N_8976);
or U9709 (N_9709,N_8850,N_8913);
and U9710 (N_9710,N_8074,N_6232);
xor U9711 (N_9711,N_6728,N_7087);
nand U9712 (N_9712,N_6680,N_7139);
nor U9713 (N_9713,N_7673,N_8603);
or U9714 (N_9714,N_6730,N_7281);
or U9715 (N_9715,N_7766,N_7447);
or U9716 (N_9716,N_6705,N_7639);
nor U9717 (N_9717,N_6492,N_8713);
or U9718 (N_9718,N_6968,N_6156);
or U9719 (N_9719,N_6226,N_7071);
and U9720 (N_9720,N_6052,N_8670);
nor U9721 (N_9721,N_6103,N_6842);
nand U9722 (N_9722,N_8784,N_7376);
or U9723 (N_9723,N_7175,N_7417);
nor U9724 (N_9724,N_8213,N_8619);
nand U9725 (N_9725,N_7540,N_7451);
nor U9726 (N_9726,N_7159,N_7641);
nor U9727 (N_9727,N_7617,N_7500);
xor U9728 (N_9728,N_7101,N_6903);
xnor U9729 (N_9729,N_6695,N_6795);
and U9730 (N_9730,N_7751,N_6500);
nand U9731 (N_9731,N_6722,N_7848);
nand U9732 (N_9732,N_7049,N_8034);
and U9733 (N_9733,N_6261,N_6785);
xor U9734 (N_9734,N_8553,N_7245);
xor U9735 (N_9735,N_7294,N_6803);
and U9736 (N_9736,N_8249,N_8563);
and U9737 (N_9737,N_8912,N_7964);
and U9738 (N_9738,N_8540,N_8872);
and U9739 (N_9739,N_8949,N_6551);
xor U9740 (N_9740,N_7100,N_6887);
or U9741 (N_9741,N_7707,N_7996);
and U9742 (N_9742,N_7176,N_6146);
nor U9743 (N_9743,N_6437,N_7084);
nor U9744 (N_9744,N_6075,N_8310);
and U9745 (N_9745,N_7291,N_8288);
nand U9746 (N_9746,N_6529,N_7859);
nor U9747 (N_9747,N_8082,N_6085);
or U9748 (N_9748,N_8258,N_8048);
nand U9749 (N_9749,N_6837,N_7315);
or U9750 (N_9750,N_6979,N_6177);
nand U9751 (N_9751,N_6139,N_7574);
and U9752 (N_9752,N_7487,N_6978);
nor U9753 (N_9753,N_8823,N_7463);
nand U9754 (N_9754,N_8890,N_8837);
and U9755 (N_9755,N_8274,N_8214);
or U9756 (N_9756,N_7624,N_6802);
or U9757 (N_9757,N_6710,N_7321);
or U9758 (N_9758,N_7373,N_6423);
or U9759 (N_9759,N_6381,N_7069);
nand U9760 (N_9760,N_7427,N_8041);
nor U9761 (N_9761,N_6403,N_8742);
or U9762 (N_9762,N_6953,N_7921);
nor U9763 (N_9763,N_8498,N_6848);
or U9764 (N_9764,N_8704,N_8273);
or U9765 (N_9765,N_8686,N_7978);
nand U9766 (N_9766,N_7450,N_7369);
nand U9767 (N_9767,N_6032,N_7184);
and U9768 (N_9768,N_6443,N_8682);
nand U9769 (N_9769,N_6247,N_6259);
or U9770 (N_9770,N_7795,N_6667);
nand U9771 (N_9771,N_8465,N_7648);
and U9772 (N_9772,N_8209,N_7971);
or U9773 (N_9773,N_6590,N_6063);
and U9774 (N_9774,N_7968,N_7865);
nand U9775 (N_9775,N_8966,N_7842);
nand U9776 (N_9776,N_7846,N_7136);
xnor U9777 (N_9777,N_7337,N_7572);
nand U9778 (N_9778,N_7290,N_7963);
or U9779 (N_9779,N_6715,N_7806);
nand U9780 (N_9780,N_7511,N_6033);
nor U9781 (N_9781,N_8132,N_7883);
or U9782 (N_9782,N_8267,N_8763);
nor U9783 (N_9783,N_7154,N_8749);
and U9784 (N_9784,N_7909,N_7568);
nand U9785 (N_9785,N_8103,N_6426);
nor U9786 (N_9786,N_7831,N_8178);
or U9787 (N_9787,N_8031,N_6128);
nand U9788 (N_9788,N_8712,N_6760);
nor U9789 (N_9789,N_7270,N_6989);
or U9790 (N_9790,N_8917,N_7401);
and U9791 (N_9791,N_6621,N_7480);
or U9792 (N_9792,N_6222,N_8953);
and U9793 (N_9793,N_7940,N_7981);
nor U9794 (N_9794,N_7844,N_8275);
nand U9795 (N_9795,N_6806,N_7238);
nand U9796 (N_9796,N_8180,N_8541);
or U9797 (N_9797,N_7977,N_6762);
nor U9798 (N_9798,N_7900,N_7821);
nand U9799 (N_9799,N_8262,N_6855);
and U9800 (N_9800,N_6657,N_8392);
xor U9801 (N_9801,N_8397,N_6255);
or U9802 (N_9802,N_8027,N_7580);
nand U9803 (N_9803,N_7987,N_7903);
nor U9804 (N_9804,N_7592,N_7585);
or U9805 (N_9805,N_7171,N_7590);
nor U9806 (N_9806,N_8047,N_6894);
or U9807 (N_9807,N_8111,N_8510);
nor U9808 (N_9808,N_6535,N_7534);
nor U9809 (N_9809,N_8897,N_6331);
or U9810 (N_9810,N_7985,N_6447);
or U9811 (N_9811,N_6023,N_6106);
and U9812 (N_9812,N_8454,N_6825);
nor U9813 (N_9813,N_6800,N_7097);
xnor U9814 (N_9814,N_6895,N_8433);
or U9815 (N_9815,N_7499,N_6320);
and U9816 (N_9816,N_6558,N_6631);
nor U9817 (N_9817,N_7258,N_7456);
nor U9818 (N_9818,N_6432,N_6870);
nor U9819 (N_9819,N_8416,N_7093);
nand U9820 (N_9820,N_7162,N_7379);
xor U9821 (N_9821,N_8951,N_7581);
and U9822 (N_9822,N_8707,N_6145);
xor U9823 (N_9823,N_8778,N_7650);
and U9824 (N_9824,N_6749,N_6030);
nand U9825 (N_9825,N_8499,N_6623);
xor U9826 (N_9826,N_6317,N_6823);
xnor U9827 (N_9827,N_6059,N_8651);
and U9828 (N_9828,N_8665,N_7685);
or U9829 (N_9829,N_7944,N_8147);
nand U9830 (N_9830,N_6595,N_6997);
or U9831 (N_9831,N_7786,N_8422);
or U9832 (N_9832,N_6025,N_8069);
nor U9833 (N_9833,N_8883,N_6852);
nor U9834 (N_9834,N_6003,N_8405);
and U9835 (N_9835,N_6723,N_8363);
and U9836 (N_9836,N_7691,N_8117);
or U9837 (N_9837,N_6436,N_8353);
nand U9838 (N_9838,N_7757,N_6994);
nor U9839 (N_9839,N_8151,N_7866);
and U9840 (N_9840,N_8927,N_8199);
and U9841 (N_9841,N_8516,N_6946);
or U9842 (N_9842,N_7279,N_7180);
nor U9843 (N_9843,N_6761,N_6736);
or U9844 (N_9844,N_6132,N_6416);
or U9845 (N_9845,N_7000,N_7221);
nand U9846 (N_9846,N_7474,N_8326);
and U9847 (N_9847,N_6001,N_8611);
nand U9848 (N_9848,N_8204,N_6901);
and U9849 (N_9849,N_6366,N_6691);
nand U9850 (N_9850,N_7075,N_7917);
and U9851 (N_9851,N_6871,N_6289);
and U9852 (N_9852,N_7342,N_6630);
nand U9853 (N_9853,N_6560,N_7651);
nor U9854 (N_9854,N_8296,N_8709);
or U9855 (N_9855,N_7682,N_6129);
nand U9856 (N_9856,N_6318,N_8009);
or U9857 (N_9857,N_8376,N_8839);
or U9858 (N_9858,N_7521,N_7198);
nor U9859 (N_9859,N_7081,N_6433);
nor U9860 (N_9860,N_6487,N_6632);
nand U9861 (N_9861,N_8165,N_8524);
nand U9862 (N_9862,N_7584,N_8108);
or U9863 (N_9863,N_6112,N_8854);
and U9864 (N_9864,N_8016,N_6906);
nor U9865 (N_9865,N_8983,N_8979);
nor U9866 (N_9866,N_6021,N_7811);
nor U9867 (N_9867,N_7547,N_6601);
and U9868 (N_9868,N_8128,N_8032);
or U9869 (N_9869,N_6904,N_8977);
and U9870 (N_9870,N_8190,N_7773);
nor U9871 (N_9871,N_7419,N_7020);
nor U9872 (N_9872,N_7830,N_7679);
and U9873 (N_9873,N_8370,N_7149);
xor U9874 (N_9874,N_7878,N_7812);
nor U9875 (N_9875,N_8606,N_7902);
or U9876 (N_9876,N_8189,N_8327);
and U9877 (N_9877,N_7755,N_8613);
nand U9878 (N_9878,N_7983,N_7626);
or U9879 (N_9879,N_8388,N_8246);
nand U9880 (N_9880,N_8975,N_8469);
or U9881 (N_9881,N_8472,N_7893);
nor U9882 (N_9882,N_6049,N_6467);
and U9883 (N_9883,N_8294,N_6886);
nand U9884 (N_9884,N_7078,N_8722);
or U9885 (N_9885,N_8669,N_7478);
or U9886 (N_9886,N_7970,N_6635);
or U9887 (N_9887,N_6155,N_6777);
and U9888 (N_9888,N_7537,N_6267);
nor U9889 (N_9889,N_7885,N_6784);
nand U9890 (N_9890,N_6942,N_8237);
nor U9891 (N_9891,N_7493,N_6829);
and U9892 (N_9892,N_7636,N_8415);
nand U9893 (N_9893,N_6921,N_8500);
and U9894 (N_9894,N_6408,N_7575);
or U9895 (N_9895,N_8769,N_6615);
or U9896 (N_9896,N_8680,N_6647);
nand U9897 (N_9897,N_8325,N_6213);
nor U9898 (N_9898,N_6641,N_6698);
and U9899 (N_9899,N_7960,N_8080);
and U9900 (N_9900,N_6941,N_8300);
and U9901 (N_9901,N_7889,N_7003);
and U9902 (N_9902,N_6817,N_7556);
xnor U9903 (N_9903,N_7274,N_6100);
or U9904 (N_9904,N_8381,N_8351);
nor U9905 (N_9905,N_8576,N_8192);
nor U9906 (N_9906,N_8569,N_7029);
nor U9907 (N_9907,N_7438,N_8923);
nor U9908 (N_9908,N_6496,N_7412);
and U9909 (N_9909,N_6909,N_6962);
and U9910 (N_9910,N_7578,N_8175);
nor U9911 (N_9911,N_7145,N_8594);
nand U9912 (N_9912,N_8359,N_8876);
or U9913 (N_9913,N_7389,N_8323);
or U9914 (N_9914,N_8135,N_8689);
nor U9915 (N_9915,N_7586,N_6206);
or U9916 (N_9916,N_7688,N_7725);
nor U9917 (N_9917,N_6646,N_7847);
nand U9918 (N_9918,N_7616,N_7140);
xor U9919 (N_9919,N_6610,N_6453);
nand U9920 (N_9920,N_7896,N_8813);
or U9921 (N_9921,N_6311,N_6703);
nand U9922 (N_9922,N_6303,N_8759);
nand U9923 (N_9923,N_7229,N_7468);
nor U9924 (N_9924,N_8930,N_7770);
or U9925 (N_9925,N_6928,N_6718);
or U9926 (N_9926,N_6484,N_6741);
or U9927 (N_9927,N_8816,N_8666);
nand U9928 (N_9928,N_8572,N_6885);
nor U9929 (N_9929,N_8427,N_7780);
nand U9930 (N_9930,N_8075,N_8184);
or U9931 (N_9931,N_6704,N_6709);
xor U9932 (N_9932,N_6018,N_8028);
or U9933 (N_9933,N_8589,N_7838);
or U9934 (N_9934,N_7792,N_7851);
or U9935 (N_9935,N_7223,N_8107);
or U9936 (N_9936,N_8329,N_6774);
xor U9937 (N_9937,N_8840,N_8932);
xor U9938 (N_9938,N_8466,N_7479);
xnor U9939 (N_9939,N_8903,N_6239);
and U9940 (N_9940,N_7596,N_7217);
and U9941 (N_9941,N_6401,N_7621);
nand U9942 (N_9942,N_6332,N_6316);
nand U9943 (N_9943,N_6924,N_6970);
nor U9944 (N_9944,N_7843,N_6217);
or U9945 (N_9945,N_8129,N_8341);
or U9946 (N_9946,N_8468,N_8085);
nor U9947 (N_9947,N_8485,N_6808);
nor U9948 (N_9948,N_8548,N_8774);
and U9949 (N_9949,N_7697,N_7070);
or U9950 (N_9950,N_8791,N_6422);
nand U9951 (N_9951,N_8477,N_6576);
and U9952 (N_9952,N_6388,N_7094);
and U9953 (N_9953,N_7259,N_7999);
nand U9954 (N_9954,N_8969,N_8287);
and U9955 (N_9955,N_7804,N_7123);
and U9956 (N_9956,N_8997,N_6746);
or U9957 (N_9957,N_6350,N_8869);
nor U9958 (N_9958,N_6503,N_6349);
or U9959 (N_9959,N_8848,N_8894);
and U9960 (N_9960,N_8293,N_6884);
and U9961 (N_9961,N_7263,N_6026);
or U9962 (N_9962,N_8906,N_6053);
or U9963 (N_9963,N_8878,N_8941);
nor U9964 (N_9964,N_8674,N_8814);
nand U9965 (N_9965,N_7849,N_8948);
nor U9966 (N_9966,N_7423,N_6675);
nor U9967 (N_9967,N_6659,N_8643);
xor U9968 (N_9968,N_6581,N_7929);
or U9969 (N_9969,N_8215,N_8493);
nand U9970 (N_9970,N_8411,N_8525);
nor U9971 (N_9971,N_7857,N_6735);
and U9972 (N_9972,N_7542,N_6039);
nor U9973 (N_9973,N_7696,N_6687);
nand U9974 (N_9974,N_7989,N_8399);
xor U9975 (N_9975,N_6596,N_6662);
and U9976 (N_9976,N_8161,N_7861);
or U9977 (N_9977,N_6012,N_6879);
or U9978 (N_9978,N_6944,N_6321);
or U9979 (N_9979,N_8308,N_6810);
nor U9980 (N_9980,N_8217,N_8068);
or U9981 (N_9981,N_8156,N_6981);
nand U9982 (N_9982,N_8684,N_8817);
nor U9983 (N_9983,N_8414,N_8862);
and U9984 (N_9984,N_7672,N_6221);
nand U9985 (N_9985,N_8773,N_7015);
nor U9986 (N_9986,N_7167,N_8693);
nand U9987 (N_9987,N_6954,N_8487);
nand U9988 (N_9988,N_7680,N_7283);
or U9989 (N_9989,N_8026,N_7443);
xor U9990 (N_9990,N_7334,N_8831);
xor U9991 (N_9991,N_7095,N_8954);
and U9992 (N_9992,N_7993,N_8486);
or U9993 (N_9993,N_6805,N_6804);
and U9994 (N_9994,N_7677,N_8797);
nand U9995 (N_9995,N_7519,N_6335);
nand U9996 (N_9996,N_8497,N_8731);
nor U9997 (N_9997,N_7335,N_6411);
or U9998 (N_9998,N_7915,N_7546);
xor U9999 (N_9999,N_6116,N_8210);
and U10000 (N_10000,N_6330,N_6559);
nor U10001 (N_10001,N_6617,N_7044);
nand U10002 (N_10002,N_8892,N_8470);
nand U10003 (N_10003,N_7317,N_7721);
or U10004 (N_10004,N_8629,N_6791);
nand U10005 (N_10005,N_6048,N_6010);
nand U10006 (N_10006,N_8808,N_7694);
and U10007 (N_10007,N_7913,N_7895);
nand U10008 (N_10008,N_8482,N_8650);
and U10009 (N_10009,N_7314,N_6395);
xnor U10010 (N_10010,N_8720,N_6815);
or U10011 (N_10011,N_7864,N_6377);
nand U10012 (N_10012,N_8081,N_7105);
or U10013 (N_10013,N_6301,N_8391);
nor U10014 (N_10014,N_8928,N_7141);
and U10015 (N_10015,N_7785,N_7637);
or U10016 (N_10016,N_7920,N_6613);
and U10017 (N_10017,N_7686,N_6888);
or U10018 (N_10018,N_7674,N_6932);
nand U10019 (N_10019,N_6937,N_7142);
nor U10020 (N_10020,N_8588,N_6198);
nor U10021 (N_10021,N_6182,N_7662);
nand U10022 (N_10022,N_8793,N_6772);
nand U10023 (N_10023,N_6219,N_8507);
or U10024 (N_10024,N_6091,N_6866);
or U10025 (N_10025,N_7352,N_7031);
nand U10026 (N_10026,N_7453,N_8899);
nand U10027 (N_10027,N_6734,N_8017);
nor U10028 (N_10028,N_8193,N_8094);
and U10029 (N_10029,N_8114,N_7348);
nor U10030 (N_10030,N_6187,N_6717);
nor U10031 (N_10031,N_6834,N_6093);
nand U10032 (N_10032,N_8212,N_8776);
nor U10033 (N_10033,N_7089,N_6726);
and U10034 (N_10034,N_7374,N_6107);
and U10035 (N_10035,N_8743,N_6302);
and U10036 (N_10036,N_7735,N_6165);
nor U10037 (N_10037,N_7991,N_7539);
and U10038 (N_10038,N_8875,N_8772);
nor U10039 (N_10039,N_7413,N_6450);
xor U10040 (N_10040,N_6755,N_7249);
xor U10041 (N_10041,N_7638,N_7912);
nand U10042 (N_10042,N_6856,N_6593);
nor U10043 (N_10043,N_7104,N_8795);
or U10044 (N_10044,N_8888,N_8860);
and U10045 (N_10045,N_7106,N_8590);
or U10046 (N_10046,N_7661,N_7216);
or U10047 (N_10047,N_8694,N_7250);
or U10048 (N_10048,N_8723,N_8302);
nor U10049 (N_10049,N_7001,N_7760);
nand U10050 (N_10050,N_7789,N_7664);
and U10051 (N_10051,N_6307,N_7988);
nand U10052 (N_10052,N_8360,N_8618);
nand U10053 (N_10053,N_8169,N_6745);
nand U10054 (N_10054,N_6826,N_6428);
nand U10055 (N_10055,N_7890,N_8076);
nor U10056 (N_10056,N_7818,N_6541);
nand U10057 (N_10057,N_6905,N_7349);
or U10058 (N_10058,N_6862,N_7967);
and U10059 (N_10059,N_8257,N_7059);
or U10060 (N_10060,N_7035,N_7126);
and U10061 (N_10061,N_7209,N_8110);
nand U10062 (N_10062,N_6579,N_8176);
or U10063 (N_10063,N_6105,N_6328);
nor U10064 (N_10064,N_8164,N_6731);
nand U10065 (N_10065,N_8062,N_7024);
nor U10066 (N_10066,N_6652,N_6421);
or U10067 (N_10067,N_6597,N_8059);
nand U10068 (N_10068,N_6714,N_6444);
or U10069 (N_10069,N_7888,N_6110);
nor U10070 (N_10070,N_7360,N_6131);
and U10071 (N_10071,N_6949,N_7272);
nand U10072 (N_10072,N_8233,N_8702);
nor U10073 (N_10073,N_7803,N_6288);
or U10074 (N_10074,N_7640,N_6046);
xor U10075 (N_10075,N_6279,N_6410);
nand U10076 (N_10076,N_7535,N_8014);
nand U10077 (N_10077,N_6205,N_6897);
or U10078 (N_10078,N_8043,N_6786);
xor U10079 (N_10079,N_7114,N_8442);
xnor U10080 (N_10080,N_8219,N_8867);
nand U10081 (N_10081,N_7296,N_6184);
or U10082 (N_10082,N_7177,N_7704);
and U10083 (N_10083,N_6486,N_7671);
nor U10084 (N_10084,N_8832,N_7192);
and U10085 (N_10085,N_7941,N_6361);
and U10086 (N_10086,N_6160,N_7026);
and U10087 (N_10087,N_8896,N_8628);
nor U10088 (N_10088,N_6183,N_7257);
or U10089 (N_10089,N_6124,N_6313);
and U10090 (N_10090,N_8463,N_6278);
or U10091 (N_10091,N_8289,N_8037);
nand U10092 (N_10092,N_7241,N_8386);
nand U10093 (N_10093,N_8013,N_6996);
and U10094 (N_10094,N_6310,N_8824);
nor U10095 (N_10095,N_6096,N_7573);
and U10096 (N_10096,N_7649,N_6756);
nand U10097 (N_10097,N_7143,N_6473);
or U10098 (N_10098,N_6355,N_7344);
nand U10099 (N_10099,N_6759,N_6324);
or U10100 (N_10100,N_6692,N_8342);
and U10101 (N_10101,N_8393,N_8092);
or U10102 (N_10102,N_8088,N_8030);
or U10103 (N_10103,N_7699,N_8079);
or U10104 (N_10104,N_6016,N_6955);
or U10105 (N_10105,N_7732,N_8278);
and U10106 (N_10106,N_8922,N_7426);
or U10107 (N_10107,N_8292,N_7875);
and U10108 (N_10108,N_6038,N_7727);
nor U10109 (N_10109,N_8887,N_7403);
and U10110 (N_10110,N_8205,N_7516);
and U10111 (N_10111,N_6542,N_6463);
nor U10112 (N_10112,N_8929,N_7157);
and U10113 (N_10113,N_6577,N_8336);
and U10114 (N_10114,N_7133,N_7408);
xor U10115 (N_10115,N_7711,N_6102);
nand U10116 (N_10116,N_8148,N_6644);
and U10117 (N_10117,N_8291,N_8004);
nand U10118 (N_10118,N_8303,N_8847);
nor U10119 (N_10119,N_8044,N_6913);
nand U10120 (N_10120,N_6015,N_6950);
or U10121 (N_10121,N_8355,N_7050);
nand U10122 (N_10122,N_7393,N_6185);
nand U10123 (N_10123,N_7186,N_8441);
xor U10124 (N_10124,N_7642,N_8227);
nor U10125 (N_10125,N_7759,N_7076);
or U10126 (N_10126,N_8886,N_6173);
or U10127 (N_10127,N_8133,N_8100);
nor U10128 (N_10128,N_7643,N_7583);
nor U10129 (N_10129,N_6531,N_6841);
nor U10130 (N_10130,N_6846,N_6120);
nand U10131 (N_10131,N_6459,N_7381);
and U10132 (N_10132,N_6396,N_6985);
nor U10133 (N_10133,N_7341,N_7323);
nand U10134 (N_10134,N_7218,N_6290);
or U10135 (N_10135,N_6526,N_6200);
and U10136 (N_10136,N_8445,N_8567);
xnor U10137 (N_10137,N_7446,N_8655);
or U10138 (N_10138,N_7079,N_6235);
nor U10139 (N_10139,N_7567,N_6987);
nand U10140 (N_10140,N_6090,N_7765);
or U10141 (N_10141,N_8750,N_7127);
or U10142 (N_10142,N_7887,N_8337);
or U10143 (N_10143,N_7261,N_7067);
nor U10144 (N_10144,N_6251,N_7212);
or U10145 (N_10145,N_7285,N_6907);
nand U10146 (N_10146,N_8127,N_7520);
nor U10147 (N_10147,N_8726,N_8794);
and U10148 (N_10148,N_7718,N_8371);
nand U10149 (N_10149,N_6298,N_7122);
nand U10150 (N_10150,N_8436,N_8314);
and U10151 (N_10151,N_7457,N_8943);
xnor U10152 (N_10152,N_6370,N_8253);
and U10153 (N_10153,N_6977,N_7955);
and U10154 (N_10154,N_6835,N_8426);
nand U10155 (N_10155,N_7465,N_8121);
nor U10156 (N_10156,N_8191,N_8881);
and U10157 (N_10157,N_7098,N_6562);
and U10158 (N_10158,N_8089,N_8304);
nor U10159 (N_10159,N_6512,N_8995);
nand U10160 (N_10160,N_8484,N_7822);
xnor U10161 (N_10161,N_8248,N_8654);
nand U10162 (N_10162,N_7681,N_6771);
nand U10163 (N_10163,N_6364,N_7593);
nand U10164 (N_10164,N_8919,N_7609);
or U10165 (N_10165,N_8141,N_8900);
nor U10166 (N_10166,N_7882,N_7820);
xor U10167 (N_10167,N_7138,N_8877);
xnor U10168 (N_10168,N_6275,N_6287);
and U10169 (N_10169,N_8673,N_7931);
or U10170 (N_10170,N_7483,N_8561);
nand U10171 (N_10171,N_8005,N_6438);
or U10172 (N_10172,N_8322,N_6268);
and U10173 (N_10173,N_8352,N_8348);
and U10174 (N_10174,N_8201,N_7187);
and U10175 (N_10175,N_6567,N_7125);
and U10176 (N_10176,N_7428,N_6262);
and U10177 (N_10177,N_6821,N_6767);
nor U10178 (N_10178,N_6599,N_7595);
or U10179 (N_10179,N_8688,N_8195);
nand U10180 (N_10180,N_8265,N_6740);
nand U10181 (N_10181,N_7984,N_6448);
nor U10182 (N_10182,N_7784,N_8203);
nand U10183 (N_10183,N_8895,N_6504);
and U10184 (N_10184,N_8999,N_8473);
and U10185 (N_10185,N_7808,N_8153);
nor U10186 (N_10186,N_6965,N_8443);
and U10187 (N_10187,N_7282,N_7062);
and U10188 (N_10188,N_8938,N_8519);
and U10189 (N_10189,N_7406,N_6794);
nand U10190 (N_10190,N_8978,N_8627);
or U10191 (N_10191,N_6700,N_7712);
or U10192 (N_10192,N_6592,N_8551);
and U10193 (N_10193,N_8357,N_7052);
and U10194 (N_10194,N_6874,N_8866);
and U10195 (N_10195,N_8194,N_7364);
xor U10196 (N_10196,N_8172,N_7594);
or U10197 (N_10197,N_6242,N_6945);
nor U10198 (N_10198,N_6406,N_8093);
or U10199 (N_10199,N_8552,N_8534);
nand U10200 (N_10200,N_7072,N_6140);
nor U10201 (N_10201,N_6516,N_7946);
nand U10202 (N_10202,N_6643,N_6375);
nand U10203 (N_10203,N_8428,N_7853);
nand U10204 (N_10204,N_8060,N_7357);
or U10205 (N_10205,N_8462,N_7827);
and U10206 (N_10206,N_7562,N_8450);
nand U10207 (N_10207,N_6614,N_8269);
and U10208 (N_10208,N_7034,N_7435);
xnor U10209 (N_10209,N_8648,N_6658);
nor U10210 (N_10210,N_7017,N_6240);
nor U10211 (N_10211,N_7045,N_6058);
nor U10212 (N_10212,N_6339,N_6520);
nand U10213 (N_10213,N_7874,N_6034);
nor U10214 (N_10214,N_6017,N_6449);
xor U10215 (N_10215,N_8738,N_8050);
or U10216 (N_10216,N_8893,N_7514);
nand U10217 (N_10217,N_8259,N_8340);
nand U10218 (N_10218,N_6101,N_8612);
nor U10219 (N_10219,N_7829,N_6780);
nor U10220 (N_10220,N_8873,N_6346);
or U10221 (N_10221,N_8057,N_6935);
and U10222 (N_10222,N_8223,N_7959);
nor U10223 (N_10223,N_7085,N_7781);
or U10224 (N_10224,N_8690,N_8266);
and U10225 (N_10225,N_6327,N_6893);
nor U10226 (N_10226,N_6031,N_7953);
nor U10227 (N_10227,N_7066,N_7675);
nor U10228 (N_10228,N_7715,N_7155);
nand U10229 (N_10229,N_8144,N_6157);
nand U10230 (N_10230,N_6392,N_6650);
nand U10231 (N_10231,N_6684,N_6258);
or U10232 (N_10232,N_7038,N_7825);
nor U10233 (N_10233,N_6539,N_6982);
nand U10234 (N_10234,N_6345,N_8102);
xnor U10235 (N_10235,N_8733,N_6796);
or U10236 (N_10236,N_8378,N_6154);
or U10237 (N_10237,N_7814,N_8744);
or U10238 (N_10238,N_7267,N_6271);
nor U10239 (N_10239,N_8926,N_8166);
nor U10240 (N_10240,N_6570,N_7656);
nor U10241 (N_10241,N_7871,N_8155);
xor U10242 (N_10242,N_6149,N_7056);
nand U10243 (N_10243,N_7116,N_6363);
and U10244 (N_10244,N_7907,N_8099);
nor U10245 (N_10245,N_7835,N_6789);
or U10246 (N_10246,N_7077,N_8595);
nand U10247 (N_10247,N_6947,N_8379);
or U10248 (N_10248,N_6940,N_8334);
and U10249 (N_10249,N_7208,N_8609);
nand U10250 (N_10250,N_6670,N_7102);
nor U10251 (N_10251,N_6229,N_6276);
nor U10252 (N_10252,N_6283,N_8116);
or U10253 (N_10253,N_6312,N_7204);
and U10254 (N_10254,N_6716,N_8070);
xor U10255 (N_10255,N_6779,N_8054);
nand U10256 (N_10256,N_6168,N_6280);
and U10257 (N_10257,N_7872,N_6292);
nor U10258 (N_10258,N_8798,N_8052);
xor U10259 (N_10259,N_8113,N_6649);
and U10260 (N_10260,N_7702,N_7332);
xor U10261 (N_10261,N_6113,N_6701);
and U10262 (N_10262,N_6868,N_8801);
nor U10263 (N_10263,N_7758,N_7440);
nand U10264 (N_10264,N_6089,N_8635);
and U10265 (N_10265,N_6414,N_6507);
nor U10266 (N_10266,N_7054,N_7558);
nor U10267 (N_10267,N_8512,N_6418);
and U10268 (N_10268,N_7012,N_6858);
xnor U10269 (N_10269,N_7391,N_8188);
nand U10270 (N_10270,N_7973,N_6147);
nand U10271 (N_10271,N_6524,N_7899);
nand U10272 (N_10272,N_6373,N_7736);
nand U10273 (N_10273,N_7005,N_6908);
nand U10274 (N_10274,N_6493,N_7676);
or U10275 (N_10275,N_6130,N_7346);
nor U10276 (N_10276,N_8630,N_7756);
nor U10277 (N_10277,N_7051,N_6464);
xnor U10278 (N_10278,N_6563,N_8810);
or U10279 (N_10279,N_8530,N_6006);
or U10280 (N_10280,N_8555,N_8592);
and U10281 (N_10281,N_6270,N_8852);
nor U10282 (N_10282,N_7634,N_8984);
nand U10283 (N_10283,N_6074,N_6050);
nor U10284 (N_10284,N_8545,N_6587);
nor U10285 (N_10285,N_8504,N_6720);
nand U10286 (N_10286,N_7833,N_8350);
xor U10287 (N_10287,N_6525,N_6665);
nand U10288 (N_10288,N_7654,N_8775);
nor U10289 (N_10289,N_7312,N_7494);
and U10290 (N_10290,N_7182,N_7555);
or U10291 (N_10291,N_8998,N_7380);
nand U10292 (N_10292,N_6685,N_6988);
nand U10293 (N_10293,N_8622,N_6490);
and U10294 (N_10294,N_7445,N_8407);
nor U10295 (N_10295,N_7128,N_6164);
or U10296 (N_10296,N_8001,N_7918);
and U10297 (N_10297,N_7061,N_8235);
or U10298 (N_10298,N_6055,N_8413);
nor U10299 (N_10299,N_7538,N_6257);
xnor U10300 (N_10300,N_8535,N_7422);
nand U10301 (N_10301,N_7235,N_6208);
nand U10302 (N_10302,N_7242,N_6594);
or U10303 (N_10303,N_6629,N_8514);
nor U10304 (N_10304,N_6589,N_8645);
nand U10305 (N_10305,N_8019,N_8792);
and U10306 (N_10306,N_8394,N_6818);
nor U10307 (N_10307,N_7027,N_7432);
nor U10308 (N_10308,N_6519,N_7815);
nand U10309 (N_10309,N_8361,N_8012);
or U10310 (N_10310,N_6743,N_7952);
nor U10311 (N_10311,N_8566,N_8398);
and U10312 (N_10312,N_7107,N_8531);
and U10313 (N_10313,N_6809,N_7659);
nand U10314 (N_10314,N_6027,N_7796);
nor U10315 (N_10315,N_8614,N_8539);
or U10316 (N_10316,N_7099,N_8737);
nor U10317 (N_10317,N_6435,N_7174);
and U10318 (N_10318,N_8717,N_8446);
and U10319 (N_10319,N_8224,N_6881);
nor U10320 (N_10320,N_6517,N_8898);
and U10321 (N_10321,N_6179,N_7046);
nand U10322 (N_10322,N_7979,N_8972);
nor U10323 (N_10323,N_6899,N_7481);
nand U10324 (N_10324,N_8023,N_7436);
nand U10325 (N_10325,N_6787,N_8586);
or U10326 (N_10326,N_7043,N_8285);
nor U10327 (N_10327,N_6993,N_6854);
and U10328 (N_10328,N_8901,N_6117);
and U10329 (N_10329,N_7147,N_8120);
nand U10330 (N_10330,N_8634,N_6627);
or U10331 (N_10331,N_6766,N_8202);
and U10332 (N_10332,N_8061,N_8335);
nand U10333 (N_10333,N_7761,N_8557);
nand U10334 (N_10334,N_8527,N_6305);
nor U10335 (N_10335,N_6358,N_7007);
nand U10336 (N_10336,N_7239,N_6309);
or U10337 (N_10337,N_8757,N_6044);
or U10338 (N_10338,N_6166,N_8208);
and U10339 (N_10339,N_6333,N_8745);
and U10340 (N_10340,N_8604,N_8828);
nor U10341 (N_10341,N_8421,N_8263);
nor U10342 (N_10342,N_6042,N_6914);
xnor U10343 (N_10343,N_7110,N_6372);
nor U10344 (N_10344,N_6163,N_6439);
or U10345 (N_10345,N_6707,N_6711);
or U10346 (N_10346,N_8549,N_8491);
nor U10347 (N_10347,N_7724,N_8008);
xnor U10348 (N_10348,N_7298,N_6850);
nand U10349 (N_10349,N_6974,N_8679);
or U10350 (N_10350,N_7425,N_6254);
and U10351 (N_10351,N_8739,N_8006);
or U10352 (N_10352,N_7295,N_8321);
and U10353 (N_10353,N_7228,N_8055);
or U10354 (N_10354,N_7452,N_8317);
nor U10355 (N_10355,N_6990,N_6153);
nand U10356 (N_10356,N_7010,N_8197);
nand U10357 (N_10357,N_8328,N_6768);
nand U10358 (N_10358,N_6654,N_6097);
nand U10359 (N_10359,N_6471,N_7064);
nand U10360 (N_10360,N_6608,N_7137);
nand U10361 (N_10361,N_6069,N_7254);
nand U10362 (N_10362,N_6571,N_7995);
or U10363 (N_10363,N_7810,N_6079);
nor U10364 (N_10364,N_6827,N_6175);
nand U10365 (N_10365,N_6495,N_8696);
and U10366 (N_10366,N_7816,N_6391);
nand U10367 (N_10367,N_7939,N_6872);
nor U10368 (N_10368,N_7030,N_6036);
or U10369 (N_10369,N_7799,N_6602);
and U10370 (N_10370,N_6919,N_6656);
nand U10371 (N_10371,N_7319,N_7421);
nor U10372 (N_10372,N_8871,N_6682);
or U10373 (N_10373,N_7949,N_7957);
and U10374 (N_10374,N_8677,N_7532);
nand U10375 (N_10375,N_8639,N_8453);
nand U10376 (N_10376,N_8483,N_8506);
nand U10377 (N_10377,N_8955,N_8664);
and U10378 (N_10378,N_8615,N_6199);
or U10379 (N_10379,N_7190,N_6431);
and U10380 (N_10380,N_6393,N_8372);
or U10381 (N_10381,N_6014,N_7090);
nand U10382 (N_10382,N_7354,N_6902);
and U10383 (N_10383,N_8232,N_6123);
nor U10384 (N_10384,N_6204,N_8730);
or U10385 (N_10385,N_6008,N_8270);
nand U10386 (N_10386,N_8065,N_8024);
or U10387 (N_10387,N_8109,N_7424);
nand U10388 (N_10388,N_7950,N_8565);
xnor U10389 (N_10389,N_7879,N_6959);
and U10390 (N_10390,N_6118,N_7880);
nand U10391 (N_10391,N_8844,N_8286);
nand U10392 (N_10392,N_8558,N_8457);
nor U10393 (N_10393,N_8683,N_6005);
or U10394 (N_10394,N_6537,N_6733);
and U10395 (N_10395,N_7778,N_7213);
or U10396 (N_10396,N_8719,N_7083);
nand U10397 (N_10397,N_7834,N_8313);
and U10398 (N_10398,N_6511,N_6376);
or U10399 (N_10399,N_8382,N_6513);
or U10400 (N_10400,N_6569,N_6297);
nand U10401 (N_10401,N_6348,N_6890);
or U10402 (N_10402,N_8678,N_7441);
or U10403 (N_10403,N_7336,N_7255);
nor U10404 (N_10404,N_6706,N_8369);
nor U10405 (N_10405,N_7313,N_8783);
nand U10406 (N_10406,N_6203,N_8647);
nor U10407 (N_10407,N_8695,N_6744);
nor U10408 (N_10408,N_6783,N_7868);
xor U10409 (N_10409,N_8904,N_7300);
and U10410 (N_10410,N_7969,N_8574);
nor U10411 (N_10411,N_7464,N_8803);
nor U10412 (N_10412,N_7368,N_7898);
nand U10413 (N_10413,N_6218,N_8710);
and U10414 (N_10414,N_7485,N_6729);
and U10415 (N_10415,N_7800,N_8729);
and U10416 (N_10416,N_6378,N_7615);
or U10417 (N_10417,N_7375,N_7199);
nand U10418 (N_10418,N_8958,N_8154);
nand U10419 (N_10419,N_6454,N_7455);
or U10420 (N_10420,N_6758,N_8354);
nand U10421 (N_10421,N_8880,N_7942);
or U10422 (N_10422,N_6737,N_8123);
or U10423 (N_10423,N_7646,N_7383);
nor U10424 (N_10424,N_8980,N_7631);
xor U10425 (N_10425,N_6142,N_7488);
or U10426 (N_10426,N_8910,N_8971);
xor U10427 (N_10427,N_7559,N_7787);
nor U10428 (N_10428,N_6702,N_7415);
and U10429 (N_10429,N_6957,N_8105);
and U10430 (N_10430,N_8261,N_6193);
and U10431 (N_10431,N_6951,N_7442);
nor U10432 (N_10432,N_8225,N_6807);
and U10433 (N_10433,N_6544,N_8119);
nor U10434 (N_10434,N_8459,N_7604);
and U10435 (N_10435,N_8532,N_8950);
and U10436 (N_10436,N_6798,N_7840);
and U10437 (N_10437,N_6078,N_8623);
nor U10438 (N_10438,N_6869,N_6765);
or U10439 (N_10439,N_6293,N_8556);
nor U10440 (N_10440,N_6900,N_8788);
xnor U10441 (N_10441,N_6586,N_6812);
and U10442 (N_10442,N_6681,N_8104);
and U10443 (N_10443,N_8543,N_8663);
nor U10444 (N_10444,N_7161,N_6099);
xor U10445 (N_10445,N_6192,N_6790);
nand U10446 (N_10446,N_7529,N_6369);
nand U10447 (N_10447,N_6934,N_6918);
nor U10448 (N_10448,N_8434,N_6167);
xor U10449 (N_10449,N_7925,N_6880);
nand U10450 (N_10450,N_7220,N_7227);
nand U10451 (N_10451,N_7683,N_8383);
nand U10452 (N_10452,N_6098,N_7901);
and U10453 (N_10453,N_7011,N_8256);
xor U10454 (N_10454,N_8542,N_8247);
or U10455 (N_10455,N_7359,N_8692);
or U10456 (N_10456,N_7576,N_8058);
nand U10457 (N_10457,N_6429,N_7231);
or U10458 (N_10458,N_8851,N_6763);
and U10459 (N_10459,N_7551,N_8228);
and U10460 (N_10460,N_8821,N_8003);
and U10461 (N_10461,N_6549,N_6161);
nand U10462 (N_10462,N_7338,N_7523);
or U10463 (N_10463,N_7193,N_7605);
and U10464 (N_10464,N_7628,N_8716);
nand U10465 (N_10465,N_8914,N_6162);
or U10466 (N_10466,N_8699,N_6523);
or U10467 (N_10467,N_8820,N_8045);
nor U10468 (N_10468,N_7032,N_6137);
xnor U10469 (N_10469,N_7390,N_8787);
or U10470 (N_10470,N_6095,N_6655);
nand U10471 (N_10471,N_6135,N_6360);
and U10472 (N_10472,N_8838,N_8478);
and U10473 (N_10473,N_6938,N_8404);
nor U10474 (N_10474,N_7938,N_8864);
or U10475 (N_10475,N_8570,N_6127);
or U10476 (N_10476,N_7053,N_8320);
xor U10477 (N_10477,N_6564,N_6816);
xnor U10478 (N_10478,N_6264,N_7462);
or U10479 (N_10479,N_6910,N_6186);
or U10480 (N_10480,N_7579,N_7768);
nand U10481 (N_10481,N_7310,N_7588);
and U10482 (N_10482,N_6233,N_7146);
or U10483 (N_10483,N_8087,N_7598);
nor U10484 (N_10484,N_6072,N_8921);
nand U10485 (N_10485,N_7163,N_6176);
nor U10486 (N_10486,N_6875,N_8324);
nand U10487 (N_10487,N_7322,N_8410);
nor U10488 (N_10488,N_8646,N_7165);
or U10489 (N_10489,N_7120,N_6673);
and U10490 (N_10490,N_7378,N_6612);
and U10491 (N_10491,N_6583,N_7306);
and U10492 (N_10492,N_8182,N_7832);
nand U10493 (N_10493,N_7363,N_6479);
nand U10494 (N_10494,N_6409,N_8339);
nor U10495 (N_10495,N_8242,N_8836);
nand U10496 (N_10496,N_7730,N_7433);
nand U10497 (N_10497,N_8475,N_7528);
or U10498 (N_10498,N_8018,N_8920);
and U10499 (N_10499,N_8961,N_8988);
and U10500 (N_10500,N_8968,N_7536);
nand U10501 (N_10501,N_8423,N_6661);
xnor U10502 (N_10502,N_7808,N_8331);
or U10503 (N_10503,N_8127,N_8912);
or U10504 (N_10504,N_8902,N_7962);
nor U10505 (N_10505,N_6343,N_6850);
nor U10506 (N_10506,N_7343,N_6145);
nand U10507 (N_10507,N_8867,N_8247);
xnor U10508 (N_10508,N_8630,N_7879);
nor U10509 (N_10509,N_6318,N_8690);
or U10510 (N_10510,N_8058,N_6179);
nor U10511 (N_10511,N_6429,N_8357);
nor U10512 (N_10512,N_6590,N_7924);
nand U10513 (N_10513,N_8823,N_7333);
or U10514 (N_10514,N_7997,N_7313);
nor U10515 (N_10515,N_8401,N_6548);
nor U10516 (N_10516,N_7682,N_8050);
nand U10517 (N_10517,N_6502,N_7234);
and U10518 (N_10518,N_7073,N_8296);
nand U10519 (N_10519,N_7205,N_8015);
and U10520 (N_10520,N_8877,N_6100);
nand U10521 (N_10521,N_6829,N_7388);
nor U10522 (N_10522,N_8530,N_8546);
xor U10523 (N_10523,N_6214,N_6913);
nor U10524 (N_10524,N_8532,N_8723);
or U10525 (N_10525,N_8029,N_7146);
nor U10526 (N_10526,N_7445,N_8247);
nor U10527 (N_10527,N_8128,N_7563);
nor U10528 (N_10528,N_8213,N_7927);
and U10529 (N_10529,N_6071,N_7790);
nor U10530 (N_10530,N_8375,N_6493);
xnor U10531 (N_10531,N_7311,N_6736);
nor U10532 (N_10532,N_7096,N_6110);
or U10533 (N_10533,N_6700,N_8376);
xnor U10534 (N_10534,N_8043,N_7390);
nand U10535 (N_10535,N_7221,N_6491);
nand U10536 (N_10536,N_8477,N_7326);
nand U10537 (N_10537,N_6716,N_7886);
and U10538 (N_10538,N_7807,N_7689);
nor U10539 (N_10539,N_6111,N_7005);
and U10540 (N_10540,N_8606,N_7813);
or U10541 (N_10541,N_8741,N_7040);
xor U10542 (N_10542,N_7600,N_7106);
nor U10543 (N_10543,N_8455,N_8377);
and U10544 (N_10544,N_6190,N_8652);
nand U10545 (N_10545,N_6668,N_8702);
and U10546 (N_10546,N_6745,N_8450);
nand U10547 (N_10547,N_8870,N_7904);
nor U10548 (N_10548,N_6496,N_7255);
nand U10549 (N_10549,N_7571,N_7757);
and U10550 (N_10550,N_8977,N_7134);
nor U10551 (N_10551,N_6081,N_6393);
and U10552 (N_10552,N_7377,N_6974);
or U10553 (N_10553,N_7024,N_6855);
and U10554 (N_10554,N_6988,N_7184);
xnor U10555 (N_10555,N_8579,N_7492);
nor U10556 (N_10556,N_6859,N_6116);
or U10557 (N_10557,N_8546,N_6864);
or U10558 (N_10558,N_8068,N_6280);
or U10559 (N_10559,N_7629,N_6450);
or U10560 (N_10560,N_6262,N_7204);
nand U10561 (N_10561,N_6523,N_6877);
xnor U10562 (N_10562,N_6759,N_7231);
nand U10563 (N_10563,N_8734,N_7526);
and U10564 (N_10564,N_8435,N_7769);
nor U10565 (N_10565,N_7214,N_7679);
nor U10566 (N_10566,N_8706,N_6244);
nor U10567 (N_10567,N_7659,N_8102);
or U10568 (N_10568,N_7164,N_6666);
nor U10569 (N_10569,N_8820,N_8654);
nand U10570 (N_10570,N_8653,N_8020);
nand U10571 (N_10571,N_7225,N_6376);
and U10572 (N_10572,N_7356,N_8229);
nand U10573 (N_10573,N_6299,N_7732);
nand U10574 (N_10574,N_8095,N_6158);
nor U10575 (N_10575,N_6496,N_7129);
and U10576 (N_10576,N_6420,N_7218);
nor U10577 (N_10577,N_6615,N_7758);
xnor U10578 (N_10578,N_8365,N_7230);
nor U10579 (N_10579,N_6567,N_6577);
xnor U10580 (N_10580,N_6980,N_8001);
nand U10581 (N_10581,N_8072,N_8299);
xor U10582 (N_10582,N_7637,N_8995);
and U10583 (N_10583,N_8744,N_6941);
xor U10584 (N_10584,N_6702,N_8627);
nor U10585 (N_10585,N_6913,N_7739);
and U10586 (N_10586,N_6505,N_7783);
and U10587 (N_10587,N_8494,N_7649);
nand U10588 (N_10588,N_6125,N_8991);
nand U10589 (N_10589,N_8701,N_7208);
nor U10590 (N_10590,N_8096,N_8507);
xor U10591 (N_10591,N_7146,N_6675);
nor U10592 (N_10592,N_6723,N_6391);
nor U10593 (N_10593,N_6109,N_8265);
nand U10594 (N_10594,N_6457,N_6430);
or U10595 (N_10595,N_7559,N_8607);
nand U10596 (N_10596,N_6655,N_7393);
and U10597 (N_10597,N_7783,N_6023);
nor U10598 (N_10598,N_6516,N_6040);
and U10599 (N_10599,N_6820,N_8426);
or U10600 (N_10600,N_6436,N_8873);
nor U10601 (N_10601,N_6320,N_7890);
nand U10602 (N_10602,N_8731,N_8172);
nand U10603 (N_10603,N_8346,N_7548);
and U10604 (N_10604,N_8857,N_8591);
and U10605 (N_10605,N_6256,N_7928);
nor U10606 (N_10606,N_8427,N_8359);
or U10607 (N_10607,N_6745,N_7266);
or U10608 (N_10608,N_7474,N_6586);
and U10609 (N_10609,N_8983,N_6881);
nor U10610 (N_10610,N_7970,N_8180);
nor U10611 (N_10611,N_8407,N_8504);
nor U10612 (N_10612,N_7594,N_6914);
or U10613 (N_10613,N_8938,N_7024);
or U10614 (N_10614,N_6709,N_7895);
and U10615 (N_10615,N_8096,N_8803);
nor U10616 (N_10616,N_7579,N_7480);
nor U10617 (N_10617,N_8804,N_8888);
nor U10618 (N_10618,N_7554,N_7850);
nor U10619 (N_10619,N_7377,N_8459);
and U10620 (N_10620,N_8261,N_6303);
nand U10621 (N_10621,N_6988,N_6827);
or U10622 (N_10622,N_6873,N_7201);
nor U10623 (N_10623,N_8015,N_7731);
nor U10624 (N_10624,N_7897,N_7327);
nand U10625 (N_10625,N_6062,N_7956);
or U10626 (N_10626,N_7531,N_7657);
nor U10627 (N_10627,N_6282,N_7137);
and U10628 (N_10628,N_8340,N_8369);
nand U10629 (N_10629,N_6292,N_7006);
nand U10630 (N_10630,N_7577,N_7155);
and U10631 (N_10631,N_7156,N_7796);
nand U10632 (N_10632,N_7379,N_6367);
nand U10633 (N_10633,N_6336,N_8534);
and U10634 (N_10634,N_6893,N_7388);
nor U10635 (N_10635,N_7510,N_6389);
or U10636 (N_10636,N_8419,N_7652);
nor U10637 (N_10637,N_6729,N_6469);
or U10638 (N_10638,N_8333,N_8769);
nand U10639 (N_10639,N_6757,N_6498);
and U10640 (N_10640,N_8117,N_7216);
nor U10641 (N_10641,N_6895,N_6653);
and U10642 (N_10642,N_7116,N_7885);
nor U10643 (N_10643,N_7905,N_6293);
nor U10644 (N_10644,N_7666,N_8702);
or U10645 (N_10645,N_7912,N_7172);
nor U10646 (N_10646,N_6250,N_8334);
nor U10647 (N_10647,N_8674,N_8442);
nor U10648 (N_10648,N_7218,N_6559);
or U10649 (N_10649,N_8117,N_6169);
or U10650 (N_10650,N_8006,N_7354);
nor U10651 (N_10651,N_7960,N_8001);
or U10652 (N_10652,N_8968,N_6638);
nor U10653 (N_10653,N_8182,N_6492);
nor U10654 (N_10654,N_6412,N_8253);
nand U10655 (N_10655,N_8057,N_7455);
and U10656 (N_10656,N_6045,N_6319);
xnor U10657 (N_10657,N_6572,N_8873);
nand U10658 (N_10658,N_8380,N_7189);
or U10659 (N_10659,N_8438,N_6901);
and U10660 (N_10660,N_8975,N_6691);
and U10661 (N_10661,N_6621,N_7439);
and U10662 (N_10662,N_6471,N_8217);
xor U10663 (N_10663,N_6445,N_7896);
or U10664 (N_10664,N_8205,N_6977);
nor U10665 (N_10665,N_8165,N_8160);
nor U10666 (N_10666,N_7529,N_6981);
nand U10667 (N_10667,N_6903,N_6231);
nor U10668 (N_10668,N_6511,N_7907);
nor U10669 (N_10669,N_6076,N_8459);
nor U10670 (N_10670,N_8722,N_8955);
nand U10671 (N_10671,N_6170,N_7674);
nor U10672 (N_10672,N_7757,N_8097);
xor U10673 (N_10673,N_8615,N_7933);
and U10674 (N_10674,N_7269,N_6842);
xnor U10675 (N_10675,N_7780,N_7836);
xor U10676 (N_10676,N_7253,N_7878);
and U10677 (N_10677,N_6402,N_7336);
nor U10678 (N_10678,N_7581,N_7289);
and U10679 (N_10679,N_8446,N_6393);
xnor U10680 (N_10680,N_7978,N_6605);
and U10681 (N_10681,N_8129,N_8343);
nand U10682 (N_10682,N_6946,N_7505);
xnor U10683 (N_10683,N_6242,N_7494);
nor U10684 (N_10684,N_6119,N_8208);
and U10685 (N_10685,N_8481,N_7611);
xor U10686 (N_10686,N_6208,N_7334);
nand U10687 (N_10687,N_6303,N_6580);
and U10688 (N_10688,N_6512,N_8689);
or U10689 (N_10689,N_8254,N_7993);
and U10690 (N_10690,N_6749,N_8820);
xnor U10691 (N_10691,N_6933,N_6117);
nor U10692 (N_10692,N_6030,N_8375);
or U10693 (N_10693,N_7307,N_7873);
or U10694 (N_10694,N_6712,N_8807);
or U10695 (N_10695,N_7812,N_6437);
and U10696 (N_10696,N_6706,N_6681);
and U10697 (N_10697,N_7018,N_8958);
and U10698 (N_10698,N_6275,N_7253);
nand U10699 (N_10699,N_7133,N_8486);
and U10700 (N_10700,N_6566,N_7321);
or U10701 (N_10701,N_6136,N_7364);
nand U10702 (N_10702,N_7204,N_8291);
nor U10703 (N_10703,N_7709,N_8248);
nand U10704 (N_10704,N_8854,N_7372);
nor U10705 (N_10705,N_6748,N_6148);
xnor U10706 (N_10706,N_6839,N_6930);
nor U10707 (N_10707,N_8432,N_8439);
and U10708 (N_10708,N_6689,N_7621);
and U10709 (N_10709,N_8233,N_7268);
xor U10710 (N_10710,N_7500,N_7007);
nor U10711 (N_10711,N_6917,N_8529);
nor U10712 (N_10712,N_6213,N_7356);
and U10713 (N_10713,N_7030,N_6882);
or U10714 (N_10714,N_8337,N_6119);
nand U10715 (N_10715,N_6219,N_6794);
nand U10716 (N_10716,N_6959,N_6597);
and U10717 (N_10717,N_6353,N_8377);
nand U10718 (N_10718,N_6193,N_7653);
and U10719 (N_10719,N_8968,N_6356);
or U10720 (N_10720,N_6929,N_6782);
and U10721 (N_10721,N_6260,N_6334);
nand U10722 (N_10722,N_8355,N_8624);
or U10723 (N_10723,N_7110,N_7617);
nor U10724 (N_10724,N_6804,N_8764);
nor U10725 (N_10725,N_8658,N_6589);
and U10726 (N_10726,N_7635,N_7251);
nor U10727 (N_10727,N_8660,N_7774);
xnor U10728 (N_10728,N_6161,N_8198);
xor U10729 (N_10729,N_6863,N_6886);
or U10730 (N_10730,N_7629,N_8808);
xor U10731 (N_10731,N_7104,N_8293);
nand U10732 (N_10732,N_8774,N_6049);
nor U10733 (N_10733,N_8622,N_7924);
nand U10734 (N_10734,N_7231,N_7648);
and U10735 (N_10735,N_8643,N_6350);
nand U10736 (N_10736,N_7628,N_8612);
or U10737 (N_10737,N_6601,N_6808);
or U10738 (N_10738,N_8057,N_7833);
nor U10739 (N_10739,N_7903,N_8532);
nand U10740 (N_10740,N_7327,N_8814);
and U10741 (N_10741,N_8535,N_6172);
nor U10742 (N_10742,N_7243,N_7491);
or U10743 (N_10743,N_7695,N_7747);
nor U10744 (N_10744,N_8929,N_6980);
nor U10745 (N_10745,N_7694,N_7440);
or U10746 (N_10746,N_8412,N_7658);
nand U10747 (N_10747,N_7390,N_8516);
or U10748 (N_10748,N_8222,N_7890);
or U10749 (N_10749,N_8766,N_8638);
or U10750 (N_10750,N_8107,N_6750);
and U10751 (N_10751,N_7866,N_6125);
nor U10752 (N_10752,N_8283,N_8864);
or U10753 (N_10753,N_7146,N_7308);
xor U10754 (N_10754,N_7743,N_8384);
nor U10755 (N_10755,N_8707,N_6680);
xor U10756 (N_10756,N_7052,N_8696);
nor U10757 (N_10757,N_8071,N_8280);
nor U10758 (N_10758,N_7583,N_7622);
or U10759 (N_10759,N_7480,N_6667);
xor U10760 (N_10760,N_8862,N_7015);
and U10761 (N_10761,N_8384,N_6986);
and U10762 (N_10762,N_6672,N_6284);
or U10763 (N_10763,N_6852,N_7531);
and U10764 (N_10764,N_8265,N_6497);
or U10765 (N_10765,N_7441,N_7580);
and U10766 (N_10766,N_8885,N_7050);
nand U10767 (N_10767,N_8822,N_6772);
nand U10768 (N_10768,N_7976,N_7822);
nor U10769 (N_10769,N_8747,N_8516);
and U10770 (N_10770,N_6011,N_8338);
and U10771 (N_10771,N_8985,N_8155);
nor U10772 (N_10772,N_8470,N_6073);
nor U10773 (N_10773,N_7761,N_7964);
nor U10774 (N_10774,N_8154,N_8459);
nor U10775 (N_10775,N_7340,N_6536);
nand U10776 (N_10776,N_7531,N_7752);
or U10777 (N_10777,N_7876,N_6729);
nor U10778 (N_10778,N_6009,N_7538);
and U10779 (N_10779,N_7167,N_7223);
or U10780 (N_10780,N_8354,N_6463);
or U10781 (N_10781,N_7501,N_6139);
nor U10782 (N_10782,N_8783,N_7055);
nand U10783 (N_10783,N_6715,N_7888);
xor U10784 (N_10784,N_6225,N_6175);
and U10785 (N_10785,N_8833,N_8037);
xnor U10786 (N_10786,N_7243,N_7594);
or U10787 (N_10787,N_6042,N_8138);
or U10788 (N_10788,N_6238,N_7410);
xnor U10789 (N_10789,N_8285,N_7330);
nand U10790 (N_10790,N_7203,N_6212);
nand U10791 (N_10791,N_7286,N_7131);
nor U10792 (N_10792,N_7356,N_8660);
nand U10793 (N_10793,N_7421,N_8247);
nand U10794 (N_10794,N_6143,N_6322);
nor U10795 (N_10795,N_6076,N_7495);
nor U10796 (N_10796,N_8439,N_8342);
nand U10797 (N_10797,N_6038,N_8018);
and U10798 (N_10798,N_6223,N_8553);
xnor U10799 (N_10799,N_8369,N_6300);
nand U10800 (N_10800,N_6582,N_7821);
and U10801 (N_10801,N_7577,N_8561);
and U10802 (N_10802,N_7600,N_7078);
or U10803 (N_10803,N_6251,N_7389);
or U10804 (N_10804,N_7951,N_7039);
and U10805 (N_10805,N_7188,N_6505);
and U10806 (N_10806,N_6420,N_8497);
nor U10807 (N_10807,N_8912,N_8451);
nor U10808 (N_10808,N_8654,N_7704);
or U10809 (N_10809,N_6974,N_8462);
or U10810 (N_10810,N_8924,N_6360);
nor U10811 (N_10811,N_6790,N_8782);
nor U10812 (N_10812,N_7746,N_8161);
or U10813 (N_10813,N_6384,N_7903);
or U10814 (N_10814,N_7249,N_6240);
nor U10815 (N_10815,N_7937,N_6500);
xnor U10816 (N_10816,N_6932,N_7049);
xor U10817 (N_10817,N_6679,N_8167);
and U10818 (N_10818,N_8019,N_6792);
and U10819 (N_10819,N_7250,N_8056);
or U10820 (N_10820,N_6868,N_8380);
or U10821 (N_10821,N_7478,N_6757);
nor U10822 (N_10822,N_6114,N_7606);
nand U10823 (N_10823,N_8842,N_8596);
nor U10824 (N_10824,N_6662,N_7682);
nand U10825 (N_10825,N_7809,N_6068);
nand U10826 (N_10826,N_7914,N_6159);
nor U10827 (N_10827,N_7407,N_6471);
nor U10828 (N_10828,N_7956,N_6576);
nand U10829 (N_10829,N_6091,N_7206);
or U10830 (N_10830,N_8082,N_6144);
xor U10831 (N_10831,N_6409,N_8435);
or U10832 (N_10832,N_6420,N_6625);
nor U10833 (N_10833,N_6798,N_8793);
xor U10834 (N_10834,N_8350,N_8417);
nor U10835 (N_10835,N_6339,N_8615);
nand U10836 (N_10836,N_7713,N_6057);
or U10837 (N_10837,N_8669,N_6814);
nand U10838 (N_10838,N_8685,N_8453);
nand U10839 (N_10839,N_6765,N_8455);
xnor U10840 (N_10840,N_6987,N_6674);
nor U10841 (N_10841,N_8542,N_8283);
nor U10842 (N_10842,N_7194,N_7826);
and U10843 (N_10843,N_8659,N_6128);
xor U10844 (N_10844,N_6581,N_6387);
nand U10845 (N_10845,N_7099,N_7278);
nand U10846 (N_10846,N_6258,N_8659);
xor U10847 (N_10847,N_8641,N_8384);
or U10848 (N_10848,N_7042,N_6320);
nor U10849 (N_10849,N_8301,N_7336);
nor U10850 (N_10850,N_8122,N_8789);
or U10851 (N_10851,N_7523,N_8420);
nand U10852 (N_10852,N_8667,N_6400);
nor U10853 (N_10853,N_6494,N_6671);
xor U10854 (N_10854,N_7792,N_6936);
and U10855 (N_10855,N_6254,N_6214);
nand U10856 (N_10856,N_8662,N_8463);
or U10857 (N_10857,N_6739,N_7027);
or U10858 (N_10858,N_7530,N_6787);
and U10859 (N_10859,N_7152,N_7525);
and U10860 (N_10860,N_7276,N_7052);
and U10861 (N_10861,N_7115,N_6007);
nor U10862 (N_10862,N_8383,N_7623);
nand U10863 (N_10863,N_6481,N_8462);
or U10864 (N_10864,N_8644,N_8319);
nand U10865 (N_10865,N_6251,N_8624);
nand U10866 (N_10866,N_8424,N_7424);
or U10867 (N_10867,N_7261,N_6900);
and U10868 (N_10868,N_6972,N_7387);
and U10869 (N_10869,N_6646,N_8149);
and U10870 (N_10870,N_6071,N_8382);
nor U10871 (N_10871,N_6994,N_8811);
xor U10872 (N_10872,N_7289,N_8624);
nor U10873 (N_10873,N_6350,N_8438);
nand U10874 (N_10874,N_8052,N_6742);
nor U10875 (N_10875,N_6745,N_7273);
xnor U10876 (N_10876,N_8347,N_7601);
or U10877 (N_10877,N_6471,N_8391);
and U10878 (N_10878,N_8984,N_7423);
nor U10879 (N_10879,N_8663,N_8628);
nor U10880 (N_10880,N_6028,N_8480);
nor U10881 (N_10881,N_7012,N_6880);
nor U10882 (N_10882,N_6462,N_8354);
nand U10883 (N_10883,N_6490,N_6746);
or U10884 (N_10884,N_6259,N_8089);
nor U10885 (N_10885,N_6110,N_6906);
and U10886 (N_10886,N_6571,N_7880);
nor U10887 (N_10887,N_7863,N_6345);
or U10888 (N_10888,N_8285,N_8016);
nand U10889 (N_10889,N_6357,N_6726);
nor U10890 (N_10890,N_8746,N_6180);
or U10891 (N_10891,N_7964,N_8085);
and U10892 (N_10892,N_7409,N_6948);
nand U10893 (N_10893,N_7911,N_7872);
nor U10894 (N_10894,N_7738,N_8551);
nor U10895 (N_10895,N_7790,N_8152);
nand U10896 (N_10896,N_7414,N_6152);
and U10897 (N_10897,N_6549,N_7307);
nor U10898 (N_10898,N_7832,N_7231);
nand U10899 (N_10899,N_6994,N_7789);
and U10900 (N_10900,N_6266,N_6609);
or U10901 (N_10901,N_8135,N_8581);
nor U10902 (N_10902,N_8416,N_7817);
nor U10903 (N_10903,N_8596,N_8641);
and U10904 (N_10904,N_8197,N_6409);
nor U10905 (N_10905,N_7383,N_6010);
nand U10906 (N_10906,N_7121,N_8456);
or U10907 (N_10907,N_8066,N_7120);
and U10908 (N_10908,N_8481,N_8359);
or U10909 (N_10909,N_8001,N_7198);
and U10910 (N_10910,N_8980,N_8654);
and U10911 (N_10911,N_8451,N_7353);
nand U10912 (N_10912,N_7458,N_8925);
nand U10913 (N_10913,N_7537,N_6008);
nand U10914 (N_10914,N_6911,N_7483);
nor U10915 (N_10915,N_8593,N_6043);
or U10916 (N_10916,N_8280,N_8338);
nand U10917 (N_10917,N_7904,N_8413);
or U10918 (N_10918,N_6566,N_6474);
and U10919 (N_10919,N_8176,N_6554);
nor U10920 (N_10920,N_8520,N_6492);
and U10921 (N_10921,N_6613,N_8957);
nand U10922 (N_10922,N_7631,N_7487);
nand U10923 (N_10923,N_6124,N_6321);
and U10924 (N_10924,N_8281,N_6481);
nor U10925 (N_10925,N_8033,N_7746);
or U10926 (N_10926,N_8279,N_6088);
and U10927 (N_10927,N_6869,N_8534);
or U10928 (N_10928,N_8274,N_8325);
and U10929 (N_10929,N_7366,N_8110);
and U10930 (N_10930,N_7516,N_7824);
and U10931 (N_10931,N_7420,N_6578);
and U10932 (N_10932,N_7434,N_6588);
nor U10933 (N_10933,N_7851,N_8273);
nor U10934 (N_10934,N_8974,N_8286);
or U10935 (N_10935,N_6352,N_8179);
nand U10936 (N_10936,N_8869,N_8670);
and U10937 (N_10937,N_7625,N_8078);
nor U10938 (N_10938,N_7185,N_8561);
or U10939 (N_10939,N_7852,N_7516);
nand U10940 (N_10940,N_6564,N_8137);
or U10941 (N_10941,N_8182,N_8359);
nor U10942 (N_10942,N_7003,N_6388);
or U10943 (N_10943,N_6958,N_7657);
xor U10944 (N_10944,N_7464,N_6921);
and U10945 (N_10945,N_6831,N_7689);
nor U10946 (N_10946,N_7725,N_7994);
and U10947 (N_10947,N_7839,N_7854);
and U10948 (N_10948,N_6759,N_7797);
or U10949 (N_10949,N_6589,N_7053);
xnor U10950 (N_10950,N_8420,N_7588);
and U10951 (N_10951,N_7433,N_8410);
or U10952 (N_10952,N_8472,N_8932);
nor U10953 (N_10953,N_8409,N_6057);
nand U10954 (N_10954,N_8141,N_8185);
nand U10955 (N_10955,N_7462,N_7693);
nor U10956 (N_10956,N_8718,N_8921);
nor U10957 (N_10957,N_8712,N_6055);
nor U10958 (N_10958,N_6346,N_7144);
nor U10959 (N_10959,N_8613,N_7763);
nand U10960 (N_10960,N_6473,N_6834);
nand U10961 (N_10961,N_7263,N_8011);
and U10962 (N_10962,N_7334,N_8632);
xor U10963 (N_10963,N_7503,N_7441);
or U10964 (N_10964,N_6975,N_7859);
and U10965 (N_10965,N_7975,N_6568);
and U10966 (N_10966,N_6415,N_7162);
or U10967 (N_10967,N_7658,N_7897);
nor U10968 (N_10968,N_6156,N_6505);
nand U10969 (N_10969,N_8618,N_7197);
nand U10970 (N_10970,N_8846,N_7803);
and U10971 (N_10971,N_7310,N_8383);
or U10972 (N_10972,N_7638,N_8142);
or U10973 (N_10973,N_6861,N_7859);
nand U10974 (N_10974,N_7997,N_6404);
nand U10975 (N_10975,N_6812,N_7098);
nand U10976 (N_10976,N_6018,N_7599);
nand U10977 (N_10977,N_6061,N_6419);
nand U10978 (N_10978,N_6249,N_6330);
and U10979 (N_10979,N_6496,N_7190);
nand U10980 (N_10980,N_7954,N_8913);
nand U10981 (N_10981,N_8340,N_7343);
and U10982 (N_10982,N_6799,N_8493);
and U10983 (N_10983,N_8771,N_7287);
xnor U10984 (N_10984,N_7755,N_6664);
nand U10985 (N_10985,N_8892,N_8176);
xnor U10986 (N_10986,N_7065,N_7744);
nor U10987 (N_10987,N_8377,N_7407);
or U10988 (N_10988,N_8483,N_8794);
nand U10989 (N_10989,N_7283,N_6128);
or U10990 (N_10990,N_7484,N_6214);
nor U10991 (N_10991,N_6633,N_8363);
xnor U10992 (N_10992,N_7201,N_8869);
nand U10993 (N_10993,N_7375,N_8827);
and U10994 (N_10994,N_8730,N_6003);
nor U10995 (N_10995,N_8313,N_8111);
nand U10996 (N_10996,N_7210,N_6785);
nand U10997 (N_10997,N_8146,N_6248);
or U10998 (N_10998,N_6139,N_6873);
nor U10999 (N_10999,N_8093,N_7007);
nor U11000 (N_11000,N_7704,N_7846);
nor U11001 (N_11001,N_6346,N_8171);
or U11002 (N_11002,N_8069,N_7688);
and U11003 (N_11003,N_8140,N_6721);
nor U11004 (N_11004,N_8862,N_8874);
or U11005 (N_11005,N_8409,N_7167);
or U11006 (N_11006,N_6630,N_6045);
and U11007 (N_11007,N_8632,N_6002);
xor U11008 (N_11008,N_6458,N_6042);
and U11009 (N_11009,N_8003,N_7181);
nand U11010 (N_11010,N_8943,N_6924);
xnor U11011 (N_11011,N_7115,N_8172);
nand U11012 (N_11012,N_7933,N_6287);
nand U11013 (N_11013,N_6651,N_7284);
nand U11014 (N_11014,N_7988,N_6213);
or U11015 (N_11015,N_7207,N_6733);
and U11016 (N_11016,N_6944,N_6533);
or U11017 (N_11017,N_6506,N_6279);
nand U11018 (N_11018,N_7404,N_8407);
or U11019 (N_11019,N_8446,N_8303);
nand U11020 (N_11020,N_7686,N_6365);
nand U11021 (N_11021,N_6578,N_7970);
xnor U11022 (N_11022,N_8620,N_8213);
or U11023 (N_11023,N_8573,N_7526);
nor U11024 (N_11024,N_7013,N_7031);
and U11025 (N_11025,N_8708,N_6211);
or U11026 (N_11026,N_6122,N_8740);
nor U11027 (N_11027,N_8932,N_8585);
nor U11028 (N_11028,N_6569,N_8761);
xnor U11029 (N_11029,N_6936,N_8248);
nor U11030 (N_11030,N_6266,N_6877);
and U11031 (N_11031,N_8173,N_7011);
nand U11032 (N_11032,N_8728,N_7889);
nor U11033 (N_11033,N_8568,N_8825);
or U11034 (N_11034,N_7137,N_7971);
and U11035 (N_11035,N_6401,N_6217);
nor U11036 (N_11036,N_8187,N_8136);
xor U11037 (N_11037,N_7604,N_8854);
and U11038 (N_11038,N_8237,N_6410);
nand U11039 (N_11039,N_8429,N_6285);
nand U11040 (N_11040,N_6075,N_7881);
xor U11041 (N_11041,N_7466,N_7609);
xor U11042 (N_11042,N_6703,N_7273);
nand U11043 (N_11043,N_6093,N_6394);
or U11044 (N_11044,N_8847,N_6976);
or U11045 (N_11045,N_6753,N_6632);
and U11046 (N_11046,N_8986,N_8071);
or U11047 (N_11047,N_8868,N_8687);
and U11048 (N_11048,N_6965,N_8924);
nand U11049 (N_11049,N_7083,N_6471);
and U11050 (N_11050,N_6060,N_6801);
nor U11051 (N_11051,N_7978,N_6334);
nand U11052 (N_11052,N_7365,N_8203);
and U11053 (N_11053,N_6457,N_7384);
nor U11054 (N_11054,N_8178,N_8104);
xor U11055 (N_11055,N_6283,N_8354);
or U11056 (N_11056,N_8838,N_7317);
xnor U11057 (N_11057,N_6106,N_8885);
and U11058 (N_11058,N_7595,N_6813);
or U11059 (N_11059,N_8238,N_6959);
nor U11060 (N_11060,N_7476,N_6427);
nor U11061 (N_11061,N_7579,N_6728);
or U11062 (N_11062,N_6167,N_8989);
or U11063 (N_11063,N_8386,N_7259);
or U11064 (N_11064,N_7519,N_7441);
nor U11065 (N_11065,N_7208,N_6291);
xnor U11066 (N_11066,N_6453,N_8613);
or U11067 (N_11067,N_6805,N_6761);
nand U11068 (N_11068,N_6641,N_7376);
and U11069 (N_11069,N_8964,N_6967);
and U11070 (N_11070,N_7003,N_8087);
or U11071 (N_11071,N_7229,N_6462);
nor U11072 (N_11072,N_6411,N_8588);
nand U11073 (N_11073,N_8829,N_8149);
and U11074 (N_11074,N_8496,N_7570);
xor U11075 (N_11075,N_8785,N_6179);
or U11076 (N_11076,N_7176,N_6010);
and U11077 (N_11077,N_8228,N_7335);
and U11078 (N_11078,N_8068,N_7015);
or U11079 (N_11079,N_6204,N_6481);
nor U11080 (N_11080,N_8756,N_8197);
and U11081 (N_11081,N_6244,N_6603);
nand U11082 (N_11082,N_7187,N_7341);
nor U11083 (N_11083,N_7835,N_6261);
xor U11084 (N_11084,N_8993,N_6392);
xor U11085 (N_11085,N_6374,N_8594);
and U11086 (N_11086,N_8816,N_6081);
or U11087 (N_11087,N_6275,N_7298);
nand U11088 (N_11088,N_7137,N_7147);
or U11089 (N_11089,N_7875,N_8165);
or U11090 (N_11090,N_8770,N_7402);
and U11091 (N_11091,N_8510,N_8515);
or U11092 (N_11092,N_6284,N_7047);
nor U11093 (N_11093,N_6619,N_8449);
xnor U11094 (N_11094,N_8988,N_8815);
nor U11095 (N_11095,N_8695,N_8476);
xnor U11096 (N_11096,N_6769,N_6967);
nand U11097 (N_11097,N_8267,N_7005);
nor U11098 (N_11098,N_6721,N_7184);
nand U11099 (N_11099,N_6839,N_8486);
and U11100 (N_11100,N_6712,N_6427);
and U11101 (N_11101,N_6574,N_7113);
nor U11102 (N_11102,N_6879,N_8848);
nor U11103 (N_11103,N_8969,N_8557);
nand U11104 (N_11104,N_7814,N_7223);
nand U11105 (N_11105,N_7658,N_6670);
nor U11106 (N_11106,N_8864,N_8920);
nand U11107 (N_11107,N_8359,N_7206);
nand U11108 (N_11108,N_7382,N_8206);
nand U11109 (N_11109,N_7400,N_6397);
or U11110 (N_11110,N_7888,N_7095);
and U11111 (N_11111,N_6530,N_8149);
xnor U11112 (N_11112,N_8203,N_6513);
and U11113 (N_11113,N_7309,N_7286);
or U11114 (N_11114,N_7166,N_8324);
nor U11115 (N_11115,N_6452,N_7789);
nand U11116 (N_11116,N_7733,N_8773);
xor U11117 (N_11117,N_7506,N_8690);
or U11118 (N_11118,N_7977,N_8882);
and U11119 (N_11119,N_6431,N_8653);
and U11120 (N_11120,N_7507,N_6081);
nand U11121 (N_11121,N_7504,N_8455);
nand U11122 (N_11122,N_6058,N_8103);
or U11123 (N_11123,N_7627,N_7439);
nand U11124 (N_11124,N_8908,N_8039);
nand U11125 (N_11125,N_8133,N_8061);
nand U11126 (N_11126,N_6245,N_6155);
nor U11127 (N_11127,N_8643,N_7744);
nor U11128 (N_11128,N_6445,N_8411);
and U11129 (N_11129,N_7576,N_6922);
or U11130 (N_11130,N_8040,N_8064);
and U11131 (N_11131,N_8063,N_6970);
or U11132 (N_11132,N_8282,N_7142);
nor U11133 (N_11133,N_6642,N_6827);
nand U11134 (N_11134,N_7785,N_8283);
and U11135 (N_11135,N_6083,N_8359);
nand U11136 (N_11136,N_6602,N_6760);
and U11137 (N_11137,N_7575,N_7118);
or U11138 (N_11138,N_6014,N_7820);
and U11139 (N_11139,N_8774,N_7199);
xor U11140 (N_11140,N_8913,N_8795);
xor U11141 (N_11141,N_8388,N_8372);
nand U11142 (N_11142,N_7503,N_6074);
or U11143 (N_11143,N_8882,N_6807);
nand U11144 (N_11144,N_7266,N_7410);
and U11145 (N_11145,N_7767,N_7880);
and U11146 (N_11146,N_8007,N_7712);
nand U11147 (N_11147,N_7553,N_7107);
and U11148 (N_11148,N_8281,N_8627);
and U11149 (N_11149,N_6763,N_7504);
xnor U11150 (N_11150,N_8937,N_8927);
and U11151 (N_11151,N_8977,N_6446);
or U11152 (N_11152,N_8673,N_6880);
or U11153 (N_11153,N_7174,N_7150);
or U11154 (N_11154,N_8689,N_6887);
xnor U11155 (N_11155,N_7999,N_6596);
nor U11156 (N_11156,N_8182,N_7040);
nor U11157 (N_11157,N_6979,N_8374);
xnor U11158 (N_11158,N_7992,N_8436);
nor U11159 (N_11159,N_8443,N_6015);
and U11160 (N_11160,N_8033,N_6467);
and U11161 (N_11161,N_7997,N_7991);
or U11162 (N_11162,N_8589,N_6693);
nand U11163 (N_11163,N_7626,N_7269);
nand U11164 (N_11164,N_6432,N_8588);
nand U11165 (N_11165,N_8735,N_7109);
and U11166 (N_11166,N_8221,N_7647);
and U11167 (N_11167,N_8205,N_8441);
nand U11168 (N_11168,N_8053,N_6580);
and U11169 (N_11169,N_6139,N_6746);
nor U11170 (N_11170,N_7535,N_8320);
and U11171 (N_11171,N_6294,N_8043);
nand U11172 (N_11172,N_8621,N_7089);
xnor U11173 (N_11173,N_6104,N_6046);
xor U11174 (N_11174,N_7076,N_8231);
and U11175 (N_11175,N_7578,N_8817);
and U11176 (N_11176,N_7310,N_8330);
nand U11177 (N_11177,N_7651,N_6911);
and U11178 (N_11178,N_7165,N_6929);
or U11179 (N_11179,N_8323,N_7670);
and U11180 (N_11180,N_6622,N_6078);
nor U11181 (N_11181,N_8462,N_6080);
or U11182 (N_11182,N_8068,N_8833);
or U11183 (N_11183,N_8342,N_8196);
xnor U11184 (N_11184,N_8719,N_8785);
nand U11185 (N_11185,N_6528,N_8601);
xor U11186 (N_11186,N_7261,N_8827);
and U11187 (N_11187,N_7666,N_8249);
and U11188 (N_11188,N_6994,N_6070);
or U11189 (N_11189,N_6307,N_8542);
nor U11190 (N_11190,N_7051,N_6519);
nor U11191 (N_11191,N_6512,N_8347);
nand U11192 (N_11192,N_6448,N_8497);
or U11193 (N_11193,N_8433,N_6671);
or U11194 (N_11194,N_8761,N_6386);
and U11195 (N_11195,N_8431,N_6084);
and U11196 (N_11196,N_6584,N_8593);
nor U11197 (N_11197,N_7239,N_7295);
or U11198 (N_11198,N_6698,N_8714);
nor U11199 (N_11199,N_6723,N_8016);
nand U11200 (N_11200,N_6806,N_6130);
xor U11201 (N_11201,N_6858,N_6806);
and U11202 (N_11202,N_6947,N_7767);
or U11203 (N_11203,N_8454,N_7087);
nand U11204 (N_11204,N_6673,N_7385);
and U11205 (N_11205,N_6645,N_8233);
and U11206 (N_11206,N_6023,N_8926);
and U11207 (N_11207,N_8639,N_6817);
or U11208 (N_11208,N_8633,N_6220);
nand U11209 (N_11209,N_8900,N_7634);
xnor U11210 (N_11210,N_6668,N_7382);
nor U11211 (N_11211,N_6878,N_7732);
and U11212 (N_11212,N_7919,N_7692);
nor U11213 (N_11213,N_7130,N_8884);
or U11214 (N_11214,N_6273,N_7451);
nand U11215 (N_11215,N_8358,N_7686);
or U11216 (N_11216,N_6396,N_6151);
or U11217 (N_11217,N_6928,N_6330);
nand U11218 (N_11218,N_8711,N_6580);
nor U11219 (N_11219,N_6835,N_6229);
and U11220 (N_11220,N_7127,N_8739);
or U11221 (N_11221,N_6478,N_8496);
nor U11222 (N_11222,N_8722,N_7436);
xnor U11223 (N_11223,N_7100,N_7682);
nor U11224 (N_11224,N_7852,N_8991);
or U11225 (N_11225,N_8379,N_6292);
or U11226 (N_11226,N_7822,N_6625);
or U11227 (N_11227,N_7101,N_7286);
and U11228 (N_11228,N_8399,N_6628);
nand U11229 (N_11229,N_7412,N_7073);
and U11230 (N_11230,N_7194,N_7663);
nor U11231 (N_11231,N_7336,N_8925);
nand U11232 (N_11232,N_7476,N_8126);
nand U11233 (N_11233,N_6709,N_8634);
and U11234 (N_11234,N_6485,N_6578);
and U11235 (N_11235,N_8303,N_8971);
nand U11236 (N_11236,N_8168,N_8703);
or U11237 (N_11237,N_7776,N_7138);
or U11238 (N_11238,N_8581,N_8249);
nand U11239 (N_11239,N_8860,N_6829);
nand U11240 (N_11240,N_8485,N_8956);
nor U11241 (N_11241,N_7766,N_7243);
and U11242 (N_11242,N_6679,N_8844);
and U11243 (N_11243,N_7500,N_7677);
nand U11244 (N_11244,N_7639,N_7813);
xnor U11245 (N_11245,N_8100,N_8531);
nand U11246 (N_11246,N_7542,N_8579);
nand U11247 (N_11247,N_6828,N_6536);
or U11248 (N_11248,N_7184,N_8593);
xor U11249 (N_11249,N_7026,N_7199);
nand U11250 (N_11250,N_8999,N_6298);
and U11251 (N_11251,N_7202,N_7930);
or U11252 (N_11252,N_8485,N_7244);
nor U11253 (N_11253,N_6503,N_8556);
and U11254 (N_11254,N_6327,N_6239);
nand U11255 (N_11255,N_6497,N_7590);
nor U11256 (N_11256,N_8547,N_7017);
nand U11257 (N_11257,N_6315,N_7638);
nor U11258 (N_11258,N_6541,N_7367);
nor U11259 (N_11259,N_7752,N_8424);
nand U11260 (N_11260,N_7366,N_6387);
or U11261 (N_11261,N_8666,N_8500);
nand U11262 (N_11262,N_7354,N_8320);
or U11263 (N_11263,N_8433,N_8311);
and U11264 (N_11264,N_7343,N_8163);
and U11265 (N_11265,N_8541,N_7826);
nor U11266 (N_11266,N_8331,N_7284);
or U11267 (N_11267,N_6303,N_7161);
and U11268 (N_11268,N_7562,N_8170);
nor U11269 (N_11269,N_7118,N_6115);
or U11270 (N_11270,N_6137,N_6482);
nand U11271 (N_11271,N_6364,N_8310);
nand U11272 (N_11272,N_7854,N_7451);
or U11273 (N_11273,N_8716,N_8365);
nand U11274 (N_11274,N_6188,N_8141);
or U11275 (N_11275,N_6888,N_7154);
xnor U11276 (N_11276,N_8890,N_8124);
or U11277 (N_11277,N_7217,N_8511);
or U11278 (N_11278,N_8272,N_6252);
nor U11279 (N_11279,N_7564,N_7373);
and U11280 (N_11280,N_6751,N_6793);
or U11281 (N_11281,N_8615,N_7132);
or U11282 (N_11282,N_7678,N_7217);
nor U11283 (N_11283,N_7897,N_8750);
or U11284 (N_11284,N_8465,N_6954);
nand U11285 (N_11285,N_6941,N_7781);
xnor U11286 (N_11286,N_8713,N_7800);
nand U11287 (N_11287,N_8821,N_6551);
or U11288 (N_11288,N_8393,N_7053);
or U11289 (N_11289,N_6922,N_7111);
nand U11290 (N_11290,N_7554,N_7114);
or U11291 (N_11291,N_8762,N_7543);
nand U11292 (N_11292,N_6485,N_7242);
or U11293 (N_11293,N_8402,N_6379);
xnor U11294 (N_11294,N_8516,N_8858);
nand U11295 (N_11295,N_7261,N_8243);
nand U11296 (N_11296,N_7124,N_6957);
or U11297 (N_11297,N_7838,N_6886);
nor U11298 (N_11298,N_6077,N_8717);
nand U11299 (N_11299,N_6609,N_7454);
nand U11300 (N_11300,N_6789,N_8662);
nor U11301 (N_11301,N_7629,N_6306);
nor U11302 (N_11302,N_8882,N_6272);
xnor U11303 (N_11303,N_6146,N_8197);
and U11304 (N_11304,N_8469,N_7604);
and U11305 (N_11305,N_6379,N_6889);
nand U11306 (N_11306,N_7351,N_7251);
nand U11307 (N_11307,N_7114,N_7856);
nor U11308 (N_11308,N_8212,N_6592);
or U11309 (N_11309,N_6569,N_7894);
or U11310 (N_11310,N_6478,N_8882);
and U11311 (N_11311,N_6817,N_6638);
nand U11312 (N_11312,N_7489,N_7701);
nor U11313 (N_11313,N_7783,N_8312);
nor U11314 (N_11314,N_8500,N_7385);
nor U11315 (N_11315,N_6240,N_7035);
nor U11316 (N_11316,N_8289,N_8812);
nand U11317 (N_11317,N_8248,N_6868);
or U11318 (N_11318,N_6360,N_8979);
nand U11319 (N_11319,N_7057,N_7029);
and U11320 (N_11320,N_8490,N_8198);
or U11321 (N_11321,N_8518,N_8363);
xnor U11322 (N_11322,N_6033,N_7357);
nor U11323 (N_11323,N_6523,N_7601);
and U11324 (N_11324,N_6436,N_8085);
nor U11325 (N_11325,N_7178,N_7212);
and U11326 (N_11326,N_6550,N_7309);
or U11327 (N_11327,N_7260,N_6342);
or U11328 (N_11328,N_6664,N_8213);
nor U11329 (N_11329,N_7920,N_7803);
nand U11330 (N_11330,N_8125,N_6730);
nand U11331 (N_11331,N_7579,N_6729);
or U11332 (N_11332,N_6522,N_8134);
nor U11333 (N_11333,N_6813,N_8111);
and U11334 (N_11334,N_8186,N_8088);
and U11335 (N_11335,N_7974,N_6690);
and U11336 (N_11336,N_7419,N_8412);
nor U11337 (N_11337,N_7378,N_6777);
nor U11338 (N_11338,N_8315,N_6961);
xor U11339 (N_11339,N_6563,N_6065);
nand U11340 (N_11340,N_6379,N_7772);
or U11341 (N_11341,N_8464,N_7787);
xnor U11342 (N_11342,N_8495,N_6237);
nand U11343 (N_11343,N_8389,N_8708);
or U11344 (N_11344,N_6615,N_6237);
nand U11345 (N_11345,N_7396,N_7631);
and U11346 (N_11346,N_6232,N_6707);
or U11347 (N_11347,N_8852,N_7393);
nand U11348 (N_11348,N_6904,N_8192);
xnor U11349 (N_11349,N_6285,N_8590);
nor U11350 (N_11350,N_7112,N_8415);
nand U11351 (N_11351,N_7950,N_7463);
nand U11352 (N_11352,N_8660,N_7083);
or U11353 (N_11353,N_6558,N_8463);
nor U11354 (N_11354,N_6684,N_7236);
or U11355 (N_11355,N_7683,N_7932);
or U11356 (N_11356,N_6194,N_7998);
nor U11357 (N_11357,N_8179,N_6895);
xor U11358 (N_11358,N_6184,N_7148);
nand U11359 (N_11359,N_6175,N_8611);
and U11360 (N_11360,N_7471,N_6537);
nor U11361 (N_11361,N_7874,N_7448);
nor U11362 (N_11362,N_6808,N_6287);
xor U11363 (N_11363,N_7360,N_6423);
nand U11364 (N_11364,N_7321,N_7820);
or U11365 (N_11365,N_6488,N_8188);
nor U11366 (N_11366,N_8980,N_7911);
or U11367 (N_11367,N_6479,N_7091);
nand U11368 (N_11368,N_6445,N_8658);
nand U11369 (N_11369,N_7106,N_8109);
or U11370 (N_11370,N_8774,N_6305);
nand U11371 (N_11371,N_7558,N_7304);
or U11372 (N_11372,N_7265,N_7350);
xor U11373 (N_11373,N_7303,N_7842);
nor U11374 (N_11374,N_7688,N_6473);
and U11375 (N_11375,N_6099,N_8802);
nand U11376 (N_11376,N_7964,N_8841);
nor U11377 (N_11377,N_8492,N_7536);
and U11378 (N_11378,N_8817,N_6466);
nor U11379 (N_11379,N_8295,N_8952);
nand U11380 (N_11380,N_8556,N_6448);
and U11381 (N_11381,N_7355,N_7897);
nand U11382 (N_11382,N_6994,N_7038);
nand U11383 (N_11383,N_6272,N_6805);
nor U11384 (N_11384,N_6911,N_7443);
nand U11385 (N_11385,N_8694,N_7047);
or U11386 (N_11386,N_8134,N_7805);
nand U11387 (N_11387,N_8437,N_6308);
and U11388 (N_11388,N_7685,N_6671);
and U11389 (N_11389,N_8064,N_8379);
nand U11390 (N_11390,N_6494,N_8366);
nand U11391 (N_11391,N_7631,N_6416);
nand U11392 (N_11392,N_8457,N_7613);
nor U11393 (N_11393,N_6869,N_7820);
xnor U11394 (N_11394,N_6362,N_8727);
xor U11395 (N_11395,N_7834,N_8280);
and U11396 (N_11396,N_8646,N_6630);
or U11397 (N_11397,N_6857,N_7739);
or U11398 (N_11398,N_8063,N_7922);
and U11399 (N_11399,N_6060,N_7110);
nor U11400 (N_11400,N_7323,N_6385);
nand U11401 (N_11401,N_8838,N_8483);
nor U11402 (N_11402,N_7277,N_6422);
nand U11403 (N_11403,N_8163,N_8144);
and U11404 (N_11404,N_6395,N_8352);
nand U11405 (N_11405,N_8139,N_6186);
nor U11406 (N_11406,N_8181,N_8362);
nor U11407 (N_11407,N_6278,N_8779);
nor U11408 (N_11408,N_7556,N_7873);
nor U11409 (N_11409,N_7783,N_7353);
or U11410 (N_11410,N_6407,N_8819);
and U11411 (N_11411,N_6640,N_6732);
nor U11412 (N_11412,N_7148,N_6730);
nand U11413 (N_11413,N_6173,N_8723);
nand U11414 (N_11414,N_8777,N_8577);
nand U11415 (N_11415,N_8991,N_8796);
or U11416 (N_11416,N_6200,N_8719);
nor U11417 (N_11417,N_7457,N_8796);
xnor U11418 (N_11418,N_7538,N_7724);
and U11419 (N_11419,N_7589,N_6383);
xnor U11420 (N_11420,N_8720,N_6127);
nand U11421 (N_11421,N_6392,N_7050);
or U11422 (N_11422,N_8033,N_8402);
nor U11423 (N_11423,N_6129,N_8201);
nor U11424 (N_11424,N_7625,N_8129);
or U11425 (N_11425,N_7593,N_7992);
or U11426 (N_11426,N_8528,N_6339);
xnor U11427 (N_11427,N_7751,N_7303);
nand U11428 (N_11428,N_6771,N_7972);
or U11429 (N_11429,N_8390,N_6607);
nand U11430 (N_11430,N_8947,N_6812);
or U11431 (N_11431,N_8300,N_6446);
xnor U11432 (N_11432,N_7875,N_7123);
nor U11433 (N_11433,N_8413,N_8220);
nor U11434 (N_11434,N_6854,N_8262);
nand U11435 (N_11435,N_7916,N_6126);
or U11436 (N_11436,N_7059,N_7468);
nand U11437 (N_11437,N_8376,N_8975);
nand U11438 (N_11438,N_8997,N_8563);
or U11439 (N_11439,N_7351,N_8119);
nor U11440 (N_11440,N_6350,N_8789);
nand U11441 (N_11441,N_7659,N_7490);
nor U11442 (N_11442,N_6664,N_6661);
or U11443 (N_11443,N_6334,N_6562);
nor U11444 (N_11444,N_8670,N_7252);
xnor U11445 (N_11445,N_8242,N_7452);
nand U11446 (N_11446,N_8757,N_8800);
and U11447 (N_11447,N_7278,N_8966);
or U11448 (N_11448,N_8361,N_7079);
and U11449 (N_11449,N_6440,N_7292);
or U11450 (N_11450,N_6471,N_8482);
or U11451 (N_11451,N_8779,N_8099);
or U11452 (N_11452,N_7562,N_6173);
or U11453 (N_11453,N_6125,N_8011);
nand U11454 (N_11454,N_8848,N_8350);
nand U11455 (N_11455,N_6211,N_8001);
or U11456 (N_11456,N_7978,N_6077);
and U11457 (N_11457,N_8439,N_8829);
and U11458 (N_11458,N_6617,N_6142);
xnor U11459 (N_11459,N_8110,N_6588);
nor U11460 (N_11460,N_7130,N_6858);
nand U11461 (N_11461,N_7387,N_6616);
or U11462 (N_11462,N_8562,N_8057);
nor U11463 (N_11463,N_6036,N_8392);
or U11464 (N_11464,N_8830,N_6365);
and U11465 (N_11465,N_7348,N_6007);
and U11466 (N_11466,N_6723,N_6007);
nand U11467 (N_11467,N_8933,N_6768);
nor U11468 (N_11468,N_6536,N_8510);
nor U11469 (N_11469,N_8721,N_7614);
nor U11470 (N_11470,N_7172,N_6012);
nand U11471 (N_11471,N_6993,N_6647);
and U11472 (N_11472,N_8592,N_8460);
xnor U11473 (N_11473,N_8303,N_6686);
xnor U11474 (N_11474,N_7032,N_8632);
nor U11475 (N_11475,N_7153,N_6256);
and U11476 (N_11476,N_7025,N_6946);
nor U11477 (N_11477,N_7848,N_6313);
and U11478 (N_11478,N_7631,N_8785);
or U11479 (N_11479,N_7835,N_7941);
or U11480 (N_11480,N_7508,N_6536);
or U11481 (N_11481,N_7788,N_8477);
or U11482 (N_11482,N_7268,N_7929);
nor U11483 (N_11483,N_7551,N_6415);
nor U11484 (N_11484,N_6673,N_8154);
xnor U11485 (N_11485,N_8582,N_8532);
and U11486 (N_11486,N_6914,N_7752);
nand U11487 (N_11487,N_6201,N_6849);
or U11488 (N_11488,N_6444,N_6480);
or U11489 (N_11489,N_7767,N_7895);
and U11490 (N_11490,N_8153,N_6928);
and U11491 (N_11491,N_6345,N_6312);
or U11492 (N_11492,N_8410,N_7820);
nor U11493 (N_11493,N_7924,N_8453);
or U11494 (N_11494,N_8975,N_8791);
and U11495 (N_11495,N_7775,N_6134);
xnor U11496 (N_11496,N_6968,N_6705);
or U11497 (N_11497,N_8929,N_6739);
nand U11498 (N_11498,N_6390,N_8656);
nor U11499 (N_11499,N_7963,N_6551);
nor U11500 (N_11500,N_6086,N_8243);
nand U11501 (N_11501,N_6093,N_7309);
or U11502 (N_11502,N_8274,N_6143);
or U11503 (N_11503,N_8441,N_8562);
nand U11504 (N_11504,N_7485,N_7888);
and U11505 (N_11505,N_6862,N_8235);
nor U11506 (N_11506,N_8826,N_7224);
or U11507 (N_11507,N_6593,N_7371);
or U11508 (N_11508,N_8400,N_7254);
nand U11509 (N_11509,N_7108,N_8129);
and U11510 (N_11510,N_7585,N_7250);
nor U11511 (N_11511,N_8433,N_6954);
or U11512 (N_11512,N_8211,N_8665);
or U11513 (N_11513,N_8951,N_6427);
nor U11514 (N_11514,N_6597,N_7114);
nand U11515 (N_11515,N_7186,N_7925);
and U11516 (N_11516,N_8316,N_6972);
nor U11517 (N_11517,N_6020,N_6355);
nor U11518 (N_11518,N_8182,N_6310);
xor U11519 (N_11519,N_7977,N_8050);
xor U11520 (N_11520,N_6447,N_6675);
nand U11521 (N_11521,N_8070,N_7801);
xor U11522 (N_11522,N_8150,N_6973);
or U11523 (N_11523,N_8593,N_8772);
nand U11524 (N_11524,N_7454,N_8331);
or U11525 (N_11525,N_6700,N_7318);
nor U11526 (N_11526,N_6148,N_6972);
and U11527 (N_11527,N_7804,N_7367);
nor U11528 (N_11528,N_7959,N_6201);
nand U11529 (N_11529,N_8953,N_8656);
nand U11530 (N_11530,N_7216,N_6243);
or U11531 (N_11531,N_6069,N_7660);
nor U11532 (N_11532,N_8715,N_6945);
nor U11533 (N_11533,N_8412,N_6695);
and U11534 (N_11534,N_6109,N_6008);
nor U11535 (N_11535,N_6725,N_8420);
or U11536 (N_11536,N_6216,N_8048);
nor U11537 (N_11537,N_7770,N_8418);
and U11538 (N_11538,N_8717,N_6898);
xor U11539 (N_11539,N_7568,N_7307);
nor U11540 (N_11540,N_7944,N_6817);
nand U11541 (N_11541,N_8782,N_6699);
nand U11542 (N_11542,N_6497,N_8558);
and U11543 (N_11543,N_7073,N_6030);
nand U11544 (N_11544,N_6923,N_7267);
nand U11545 (N_11545,N_6435,N_7609);
nor U11546 (N_11546,N_8856,N_7582);
nand U11547 (N_11547,N_7627,N_8253);
or U11548 (N_11548,N_7090,N_6612);
and U11549 (N_11549,N_6701,N_8955);
nand U11550 (N_11550,N_7485,N_8357);
or U11551 (N_11551,N_6869,N_8314);
nand U11552 (N_11552,N_6606,N_6882);
or U11553 (N_11553,N_8548,N_7205);
nand U11554 (N_11554,N_6350,N_7497);
xnor U11555 (N_11555,N_7331,N_8858);
and U11556 (N_11556,N_7934,N_8766);
nor U11557 (N_11557,N_8535,N_7809);
nor U11558 (N_11558,N_8623,N_6013);
nand U11559 (N_11559,N_6953,N_8848);
or U11560 (N_11560,N_6484,N_7999);
nand U11561 (N_11561,N_8201,N_7980);
or U11562 (N_11562,N_6945,N_8271);
and U11563 (N_11563,N_8990,N_8862);
or U11564 (N_11564,N_7488,N_6720);
xnor U11565 (N_11565,N_6924,N_8969);
or U11566 (N_11566,N_7682,N_7589);
nand U11567 (N_11567,N_6046,N_8998);
or U11568 (N_11568,N_7823,N_7467);
or U11569 (N_11569,N_7170,N_7331);
nor U11570 (N_11570,N_7897,N_8912);
or U11571 (N_11571,N_8133,N_6957);
nor U11572 (N_11572,N_7874,N_7196);
or U11573 (N_11573,N_7180,N_6402);
or U11574 (N_11574,N_8565,N_8111);
or U11575 (N_11575,N_7982,N_8103);
or U11576 (N_11576,N_6660,N_8097);
nand U11577 (N_11577,N_6017,N_8439);
nand U11578 (N_11578,N_7174,N_7814);
nor U11579 (N_11579,N_6144,N_8773);
nor U11580 (N_11580,N_7809,N_6571);
and U11581 (N_11581,N_8223,N_6163);
or U11582 (N_11582,N_8572,N_8691);
nand U11583 (N_11583,N_8118,N_7911);
xor U11584 (N_11584,N_7239,N_6690);
or U11585 (N_11585,N_7407,N_6772);
and U11586 (N_11586,N_7062,N_8005);
and U11587 (N_11587,N_7199,N_8586);
nor U11588 (N_11588,N_6145,N_8965);
nand U11589 (N_11589,N_8788,N_7525);
or U11590 (N_11590,N_8446,N_6432);
xor U11591 (N_11591,N_6373,N_7426);
or U11592 (N_11592,N_8404,N_6688);
or U11593 (N_11593,N_8451,N_6210);
nand U11594 (N_11594,N_6393,N_7395);
and U11595 (N_11595,N_6213,N_6061);
and U11596 (N_11596,N_8508,N_7278);
nor U11597 (N_11597,N_7917,N_6032);
and U11598 (N_11598,N_8581,N_7095);
or U11599 (N_11599,N_7143,N_7725);
nand U11600 (N_11600,N_7224,N_8637);
or U11601 (N_11601,N_7121,N_7616);
or U11602 (N_11602,N_8758,N_6494);
nor U11603 (N_11603,N_6909,N_6168);
nand U11604 (N_11604,N_8621,N_6168);
nor U11605 (N_11605,N_6989,N_7302);
or U11606 (N_11606,N_8390,N_6535);
nor U11607 (N_11607,N_7468,N_7623);
or U11608 (N_11608,N_7317,N_6874);
nand U11609 (N_11609,N_8164,N_8436);
nand U11610 (N_11610,N_8464,N_7984);
nand U11611 (N_11611,N_7538,N_8353);
nor U11612 (N_11612,N_8352,N_8201);
and U11613 (N_11613,N_8858,N_7732);
or U11614 (N_11614,N_7754,N_8194);
and U11615 (N_11615,N_7464,N_8531);
and U11616 (N_11616,N_6895,N_8051);
and U11617 (N_11617,N_7870,N_6338);
and U11618 (N_11618,N_7729,N_7004);
or U11619 (N_11619,N_8849,N_7978);
and U11620 (N_11620,N_6338,N_7727);
and U11621 (N_11621,N_7186,N_7762);
nand U11622 (N_11622,N_7125,N_6730);
nor U11623 (N_11623,N_8483,N_8160);
nand U11624 (N_11624,N_7677,N_8674);
nand U11625 (N_11625,N_8687,N_7097);
nand U11626 (N_11626,N_7735,N_8223);
and U11627 (N_11627,N_7379,N_7123);
nand U11628 (N_11628,N_7823,N_6874);
nand U11629 (N_11629,N_8084,N_8055);
or U11630 (N_11630,N_7036,N_6016);
nand U11631 (N_11631,N_8025,N_8530);
nor U11632 (N_11632,N_7543,N_8179);
or U11633 (N_11633,N_7828,N_7879);
or U11634 (N_11634,N_7094,N_8269);
nand U11635 (N_11635,N_8000,N_7126);
or U11636 (N_11636,N_6015,N_8949);
nor U11637 (N_11637,N_6236,N_7548);
xor U11638 (N_11638,N_7749,N_7627);
nor U11639 (N_11639,N_6364,N_6856);
nor U11640 (N_11640,N_7557,N_8281);
nand U11641 (N_11641,N_8680,N_6832);
nand U11642 (N_11642,N_8986,N_6874);
nor U11643 (N_11643,N_8897,N_6490);
nor U11644 (N_11644,N_8914,N_8832);
nor U11645 (N_11645,N_8428,N_6314);
nor U11646 (N_11646,N_6912,N_6468);
and U11647 (N_11647,N_7266,N_8344);
or U11648 (N_11648,N_7498,N_8747);
and U11649 (N_11649,N_8559,N_8640);
nand U11650 (N_11650,N_6963,N_8932);
or U11651 (N_11651,N_7480,N_8001);
nor U11652 (N_11652,N_6991,N_6772);
nor U11653 (N_11653,N_6574,N_8498);
or U11654 (N_11654,N_6854,N_8744);
nor U11655 (N_11655,N_8881,N_7255);
and U11656 (N_11656,N_8415,N_7037);
nand U11657 (N_11657,N_8095,N_6880);
nand U11658 (N_11658,N_6718,N_8204);
or U11659 (N_11659,N_7883,N_8191);
nor U11660 (N_11660,N_6427,N_7424);
nand U11661 (N_11661,N_8560,N_8879);
and U11662 (N_11662,N_7283,N_6614);
and U11663 (N_11663,N_6183,N_6577);
nand U11664 (N_11664,N_8006,N_8702);
and U11665 (N_11665,N_7159,N_7707);
nor U11666 (N_11666,N_6190,N_6865);
nand U11667 (N_11667,N_6944,N_8240);
nand U11668 (N_11668,N_6153,N_7811);
nor U11669 (N_11669,N_6977,N_8150);
or U11670 (N_11670,N_6843,N_6500);
or U11671 (N_11671,N_8844,N_7637);
and U11672 (N_11672,N_8880,N_8838);
nand U11673 (N_11673,N_6704,N_8224);
nand U11674 (N_11674,N_8133,N_6253);
and U11675 (N_11675,N_6750,N_7161);
nor U11676 (N_11676,N_6146,N_8423);
or U11677 (N_11677,N_7155,N_8289);
and U11678 (N_11678,N_7615,N_7898);
and U11679 (N_11679,N_7037,N_6942);
and U11680 (N_11680,N_7006,N_7901);
and U11681 (N_11681,N_8828,N_8275);
nand U11682 (N_11682,N_8169,N_7966);
nand U11683 (N_11683,N_7460,N_7909);
xnor U11684 (N_11684,N_8902,N_8686);
or U11685 (N_11685,N_6468,N_7030);
or U11686 (N_11686,N_7884,N_8823);
nor U11687 (N_11687,N_7384,N_8150);
nand U11688 (N_11688,N_7517,N_6456);
and U11689 (N_11689,N_6144,N_6170);
nor U11690 (N_11690,N_7298,N_7421);
nand U11691 (N_11691,N_7306,N_8163);
nand U11692 (N_11692,N_6699,N_8244);
nor U11693 (N_11693,N_8048,N_6540);
nand U11694 (N_11694,N_6892,N_8242);
nor U11695 (N_11695,N_6687,N_8062);
and U11696 (N_11696,N_6353,N_6032);
or U11697 (N_11697,N_6877,N_8087);
nand U11698 (N_11698,N_7040,N_7823);
or U11699 (N_11699,N_6970,N_7964);
nor U11700 (N_11700,N_7977,N_6842);
nor U11701 (N_11701,N_6590,N_8895);
nor U11702 (N_11702,N_6408,N_6854);
and U11703 (N_11703,N_7279,N_6955);
and U11704 (N_11704,N_7457,N_6930);
nor U11705 (N_11705,N_6239,N_6051);
xnor U11706 (N_11706,N_6046,N_7863);
xor U11707 (N_11707,N_8761,N_7670);
nand U11708 (N_11708,N_6526,N_7480);
or U11709 (N_11709,N_7617,N_8548);
nor U11710 (N_11710,N_6920,N_6081);
nand U11711 (N_11711,N_8307,N_8220);
nor U11712 (N_11712,N_8566,N_7214);
nor U11713 (N_11713,N_7085,N_6337);
nor U11714 (N_11714,N_6026,N_7218);
or U11715 (N_11715,N_6604,N_7897);
nor U11716 (N_11716,N_6457,N_8022);
and U11717 (N_11717,N_6722,N_6202);
nand U11718 (N_11718,N_7880,N_6060);
nand U11719 (N_11719,N_7182,N_6893);
or U11720 (N_11720,N_8197,N_6121);
and U11721 (N_11721,N_6923,N_7561);
or U11722 (N_11722,N_6905,N_6174);
and U11723 (N_11723,N_8339,N_7497);
nor U11724 (N_11724,N_6456,N_7658);
or U11725 (N_11725,N_8527,N_7328);
or U11726 (N_11726,N_8729,N_6304);
or U11727 (N_11727,N_6878,N_6488);
nor U11728 (N_11728,N_8518,N_7333);
or U11729 (N_11729,N_6977,N_6651);
and U11730 (N_11730,N_6448,N_7691);
and U11731 (N_11731,N_7754,N_8385);
nand U11732 (N_11732,N_8989,N_6842);
or U11733 (N_11733,N_8778,N_6351);
nor U11734 (N_11734,N_8746,N_8071);
nor U11735 (N_11735,N_8546,N_6455);
xor U11736 (N_11736,N_7567,N_8719);
nor U11737 (N_11737,N_6641,N_7571);
and U11738 (N_11738,N_7298,N_7381);
nand U11739 (N_11739,N_6082,N_8618);
or U11740 (N_11740,N_8724,N_7486);
nand U11741 (N_11741,N_6416,N_8364);
and U11742 (N_11742,N_6895,N_8843);
or U11743 (N_11743,N_7703,N_7735);
nor U11744 (N_11744,N_7802,N_6385);
nand U11745 (N_11745,N_6155,N_6635);
nor U11746 (N_11746,N_7839,N_6526);
nor U11747 (N_11747,N_6507,N_7435);
nand U11748 (N_11748,N_6001,N_6639);
and U11749 (N_11749,N_6659,N_7675);
nand U11750 (N_11750,N_8029,N_6410);
nand U11751 (N_11751,N_7146,N_8621);
nor U11752 (N_11752,N_7219,N_8755);
nor U11753 (N_11753,N_6130,N_8845);
nand U11754 (N_11754,N_7292,N_8859);
nand U11755 (N_11755,N_7127,N_8113);
or U11756 (N_11756,N_6319,N_6771);
and U11757 (N_11757,N_7251,N_7421);
and U11758 (N_11758,N_8300,N_6138);
and U11759 (N_11759,N_6718,N_6438);
nor U11760 (N_11760,N_7796,N_8377);
nor U11761 (N_11761,N_8626,N_8321);
nor U11762 (N_11762,N_7650,N_8986);
and U11763 (N_11763,N_8149,N_6793);
nor U11764 (N_11764,N_8268,N_7632);
nor U11765 (N_11765,N_8435,N_6400);
nand U11766 (N_11766,N_6072,N_7816);
or U11767 (N_11767,N_8918,N_7128);
xnor U11768 (N_11768,N_7990,N_6688);
and U11769 (N_11769,N_7735,N_8958);
and U11770 (N_11770,N_7246,N_6194);
or U11771 (N_11771,N_8812,N_7327);
or U11772 (N_11772,N_7126,N_8475);
nor U11773 (N_11773,N_6784,N_7868);
or U11774 (N_11774,N_6736,N_6573);
and U11775 (N_11775,N_6689,N_7396);
or U11776 (N_11776,N_7545,N_7619);
and U11777 (N_11777,N_7496,N_6420);
nor U11778 (N_11778,N_8916,N_7306);
nand U11779 (N_11779,N_7976,N_7261);
or U11780 (N_11780,N_7280,N_6130);
nand U11781 (N_11781,N_6756,N_6761);
nor U11782 (N_11782,N_6008,N_6943);
or U11783 (N_11783,N_7343,N_6608);
nand U11784 (N_11784,N_8178,N_6162);
nor U11785 (N_11785,N_7000,N_6088);
xnor U11786 (N_11786,N_8825,N_7343);
nor U11787 (N_11787,N_7314,N_7176);
nor U11788 (N_11788,N_7097,N_7539);
nor U11789 (N_11789,N_7114,N_8673);
and U11790 (N_11790,N_7012,N_6712);
or U11791 (N_11791,N_6656,N_6660);
nand U11792 (N_11792,N_7764,N_8187);
or U11793 (N_11793,N_8919,N_7733);
or U11794 (N_11794,N_8695,N_8002);
nor U11795 (N_11795,N_8462,N_7017);
nand U11796 (N_11796,N_6121,N_7352);
nand U11797 (N_11797,N_8128,N_7749);
xnor U11798 (N_11798,N_7438,N_8643);
nor U11799 (N_11799,N_7399,N_8596);
nor U11800 (N_11800,N_7605,N_6623);
or U11801 (N_11801,N_6612,N_8809);
nand U11802 (N_11802,N_8010,N_7691);
xnor U11803 (N_11803,N_8120,N_6133);
nand U11804 (N_11804,N_7382,N_8812);
or U11805 (N_11805,N_8587,N_7083);
nand U11806 (N_11806,N_8183,N_7433);
and U11807 (N_11807,N_6573,N_8436);
and U11808 (N_11808,N_6863,N_7495);
and U11809 (N_11809,N_6128,N_8976);
nor U11810 (N_11810,N_6165,N_7110);
and U11811 (N_11811,N_7505,N_6391);
and U11812 (N_11812,N_8443,N_8077);
or U11813 (N_11813,N_6540,N_8567);
and U11814 (N_11814,N_7978,N_7995);
and U11815 (N_11815,N_8166,N_6232);
or U11816 (N_11816,N_7156,N_8941);
nand U11817 (N_11817,N_7539,N_7442);
nor U11818 (N_11818,N_8164,N_6143);
and U11819 (N_11819,N_6461,N_8114);
nor U11820 (N_11820,N_6955,N_6491);
and U11821 (N_11821,N_8768,N_6262);
nor U11822 (N_11822,N_8572,N_6056);
nor U11823 (N_11823,N_6154,N_6171);
nand U11824 (N_11824,N_7139,N_8813);
or U11825 (N_11825,N_8728,N_6793);
nand U11826 (N_11826,N_6931,N_6993);
xnor U11827 (N_11827,N_7148,N_6372);
and U11828 (N_11828,N_8839,N_8428);
or U11829 (N_11829,N_7703,N_6814);
or U11830 (N_11830,N_6475,N_8658);
xor U11831 (N_11831,N_8226,N_8754);
nor U11832 (N_11832,N_6524,N_6899);
or U11833 (N_11833,N_8005,N_8521);
or U11834 (N_11834,N_6319,N_6121);
and U11835 (N_11835,N_8937,N_7300);
nor U11836 (N_11836,N_8389,N_7709);
or U11837 (N_11837,N_8958,N_7996);
and U11838 (N_11838,N_6909,N_7887);
or U11839 (N_11839,N_6292,N_7275);
or U11840 (N_11840,N_7999,N_7674);
and U11841 (N_11841,N_8761,N_8864);
nand U11842 (N_11842,N_6847,N_8824);
nand U11843 (N_11843,N_6265,N_6348);
and U11844 (N_11844,N_6041,N_7014);
nor U11845 (N_11845,N_7670,N_8662);
nand U11846 (N_11846,N_8044,N_7476);
xor U11847 (N_11847,N_8267,N_6424);
and U11848 (N_11848,N_7148,N_6449);
or U11849 (N_11849,N_6202,N_8130);
and U11850 (N_11850,N_7513,N_6021);
and U11851 (N_11851,N_6541,N_7586);
or U11852 (N_11852,N_7518,N_8855);
xnor U11853 (N_11853,N_8048,N_8559);
or U11854 (N_11854,N_8050,N_8236);
nor U11855 (N_11855,N_8018,N_8151);
and U11856 (N_11856,N_8868,N_8741);
or U11857 (N_11857,N_8921,N_6458);
and U11858 (N_11858,N_8806,N_6021);
or U11859 (N_11859,N_8343,N_7864);
and U11860 (N_11860,N_8510,N_8079);
or U11861 (N_11861,N_6138,N_6056);
nor U11862 (N_11862,N_6743,N_8088);
xnor U11863 (N_11863,N_6989,N_8268);
nor U11864 (N_11864,N_7549,N_6731);
and U11865 (N_11865,N_6678,N_7444);
nand U11866 (N_11866,N_8517,N_7457);
and U11867 (N_11867,N_6759,N_6671);
and U11868 (N_11868,N_7495,N_8659);
or U11869 (N_11869,N_8191,N_6900);
xor U11870 (N_11870,N_6573,N_7431);
nand U11871 (N_11871,N_6638,N_8459);
xor U11872 (N_11872,N_8713,N_7410);
and U11873 (N_11873,N_8151,N_7174);
nor U11874 (N_11874,N_7237,N_7016);
nor U11875 (N_11875,N_8436,N_6839);
and U11876 (N_11876,N_6788,N_6078);
and U11877 (N_11877,N_6183,N_8424);
nor U11878 (N_11878,N_7733,N_6166);
or U11879 (N_11879,N_7597,N_6460);
or U11880 (N_11880,N_7425,N_8199);
nor U11881 (N_11881,N_7567,N_6932);
and U11882 (N_11882,N_6404,N_7308);
nor U11883 (N_11883,N_8760,N_6594);
nor U11884 (N_11884,N_6151,N_6891);
nor U11885 (N_11885,N_7776,N_6849);
and U11886 (N_11886,N_6024,N_6938);
nor U11887 (N_11887,N_8621,N_7104);
nand U11888 (N_11888,N_8017,N_7507);
nand U11889 (N_11889,N_8272,N_7879);
and U11890 (N_11890,N_6164,N_8573);
nor U11891 (N_11891,N_8152,N_7731);
and U11892 (N_11892,N_7441,N_8384);
and U11893 (N_11893,N_6616,N_8130);
nand U11894 (N_11894,N_6165,N_7238);
and U11895 (N_11895,N_6759,N_7816);
or U11896 (N_11896,N_6170,N_7373);
nand U11897 (N_11897,N_6681,N_7041);
or U11898 (N_11898,N_7349,N_8198);
and U11899 (N_11899,N_8975,N_6055);
or U11900 (N_11900,N_6156,N_6938);
xnor U11901 (N_11901,N_7689,N_8524);
and U11902 (N_11902,N_7997,N_8042);
xor U11903 (N_11903,N_7697,N_8061);
nor U11904 (N_11904,N_8065,N_6469);
nand U11905 (N_11905,N_7506,N_7835);
nor U11906 (N_11906,N_6341,N_6534);
nor U11907 (N_11907,N_6518,N_8590);
or U11908 (N_11908,N_7200,N_8105);
nor U11909 (N_11909,N_7478,N_8462);
nor U11910 (N_11910,N_6641,N_7040);
nand U11911 (N_11911,N_8935,N_8530);
xnor U11912 (N_11912,N_8840,N_8389);
or U11913 (N_11913,N_7851,N_8168);
or U11914 (N_11914,N_7089,N_7327);
or U11915 (N_11915,N_8541,N_7899);
or U11916 (N_11916,N_6874,N_8684);
nor U11917 (N_11917,N_8067,N_8651);
or U11918 (N_11918,N_6203,N_6925);
nor U11919 (N_11919,N_6745,N_8873);
xor U11920 (N_11920,N_7138,N_8810);
nor U11921 (N_11921,N_6232,N_7705);
or U11922 (N_11922,N_7918,N_8485);
or U11923 (N_11923,N_7305,N_6989);
nor U11924 (N_11924,N_8251,N_7576);
and U11925 (N_11925,N_8155,N_7502);
nand U11926 (N_11926,N_8013,N_8091);
xnor U11927 (N_11927,N_8834,N_8699);
nor U11928 (N_11928,N_8409,N_6298);
nor U11929 (N_11929,N_6562,N_8443);
nand U11930 (N_11930,N_7465,N_6810);
nor U11931 (N_11931,N_7610,N_6268);
or U11932 (N_11932,N_7862,N_8898);
nand U11933 (N_11933,N_6878,N_6083);
and U11934 (N_11934,N_8916,N_8576);
nor U11935 (N_11935,N_6023,N_6969);
and U11936 (N_11936,N_7954,N_8421);
or U11937 (N_11937,N_8435,N_7198);
and U11938 (N_11938,N_8296,N_8747);
nor U11939 (N_11939,N_7330,N_8793);
and U11940 (N_11940,N_7837,N_8431);
nor U11941 (N_11941,N_6465,N_7039);
nand U11942 (N_11942,N_8793,N_6320);
nor U11943 (N_11943,N_8393,N_8733);
and U11944 (N_11944,N_8946,N_8461);
or U11945 (N_11945,N_8351,N_6738);
and U11946 (N_11946,N_6445,N_7506);
and U11947 (N_11947,N_8948,N_7885);
xnor U11948 (N_11948,N_8777,N_7588);
or U11949 (N_11949,N_8713,N_6620);
and U11950 (N_11950,N_7205,N_8933);
xnor U11951 (N_11951,N_8224,N_6365);
nor U11952 (N_11952,N_6669,N_7707);
nand U11953 (N_11953,N_6357,N_6399);
and U11954 (N_11954,N_6679,N_7624);
nand U11955 (N_11955,N_8986,N_8366);
xor U11956 (N_11956,N_8358,N_7149);
nor U11957 (N_11957,N_6783,N_7240);
and U11958 (N_11958,N_6190,N_7030);
nor U11959 (N_11959,N_8869,N_8703);
nand U11960 (N_11960,N_7041,N_8169);
and U11961 (N_11961,N_8829,N_8443);
and U11962 (N_11962,N_6824,N_8522);
and U11963 (N_11963,N_6863,N_6281);
or U11964 (N_11964,N_6678,N_8894);
and U11965 (N_11965,N_8053,N_6002);
and U11966 (N_11966,N_6321,N_7491);
nand U11967 (N_11967,N_7247,N_8381);
and U11968 (N_11968,N_8970,N_6655);
nor U11969 (N_11969,N_8954,N_6377);
xnor U11970 (N_11970,N_6227,N_8046);
and U11971 (N_11971,N_7621,N_6831);
nor U11972 (N_11972,N_7275,N_6988);
xnor U11973 (N_11973,N_6231,N_7034);
nand U11974 (N_11974,N_8521,N_7695);
and U11975 (N_11975,N_6270,N_8101);
and U11976 (N_11976,N_8977,N_7066);
or U11977 (N_11977,N_7853,N_7518);
nand U11978 (N_11978,N_6952,N_6290);
or U11979 (N_11979,N_7328,N_7552);
and U11980 (N_11980,N_7830,N_7641);
or U11981 (N_11981,N_6358,N_7160);
and U11982 (N_11982,N_7563,N_6243);
nor U11983 (N_11983,N_8981,N_7015);
nor U11984 (N_11984,N_8340,N_7551);
nor U11985 (N_11985,N_6361,N_6964);
nor U11986 (N_11986,N_7966,N_7169);
nand U11987 (N_11987,N_6099,N_6690);
nor U11988 (N_11988,N_6852,N_8354);
or U11989 (N_11989,N_6505,N_6692);
xnor U11990 (N_11990,N_8620,N_6019);
nor U11991 (N_11991,N_7054,N_7370);
xnor U11992 (N_11992,N_7882,N_8441);
xor U11993 (N_11993,N_8786,N_8627);
nor U11994 (N_11994,N_8455,N_8412);
nor U11995 (N_11995,N_6488,N_8736);
and U11996 (N_11996,N_7138,N_6270);
xor U11997 (N_11997,N_7611,N_7672);
xnor U11998 (N_11998,N_7028,N_6872);
and U11999 (N_11999,N_8683,N_6552);
or U12000 (N_12000,N_11557,N_10239);
and U12001 (N_12001,N_10599,N_10864);
or U12002 (N_12002,N_11204,N_11176);
nand U12003 (N_12003,N_11921,N_10028);
nor U12004 (N_12004,N_11784,N_11883);
xor U12005 (N_12005,N_11905,N_11459);
nand U12006 (N_12006,N_10308,N_9107);
and U12007 (N_12007,N_9158,N_9860);
xor U12008 (N_12008,N_9822,N_10684);
nor U12009 (N_12009,N_11214,N_11353);
xnor U12010 (N_12010,N_9144,N_11997);
or U12011 (N_12011,N_9913,N_11275);
and U12012 (N_12012,N_11162,N_11229);
nand U12013 (N_12013,N_11568,N_11213);
nor U12014 (N_12014,N_9093,N_10530);
xor U12015 (N_12015,N_9876,N_11485);
and U12016 (N_12016,N_11645,N_11281);
nor U12017 (N_12017,N_10162,N_11516);
nor U12018 (N_12018,N_11634,N_9960);
nand U12019 (N_12019,N_11196,N_11564);
or U12020 (N_12020,N_9234,N_10708);
and U12021 (N_12021,N_10742,N_9492);
and U12022 (N_12022,N_10422,N_11335);
and U12023 (N_12023,N_11394,N_9317);
xor U12024 (N_12024,N_10492,N_11963);
nor U12025 (N_12025,N_10836,N_11683);
and U12026 (N_12026,N_9374,N_9590);
nand U12027 (N_12027,N_11741,N_11014);
and U12028 (N_12028,N_10786,N_10469);
nor U12029 (N_12029,N_9662,N_11679);
nand U12030 (N_12030,N_11492,N_9136);
nor U12031 (N_12031,N_11413,N_9568);
nand U12032 (N_12032,N_11999,N_11414);
or U12033 (N_12033,N_11234,N_11606);
nor U12034 (N_12034,N_10484,N_10704);
nand U12035 (N_12035,N_9165,N_10342);
nor U12036 (N_12036,N_11582,N_10848);
nand U12037 (N_12037,N_9983,N_10459);
nor U12038 (N_12038,N_10040,N_9402);
nand U12039 (N_12039,N_10041,N_11276);
nor U12040 (N_12040,N_10688,N_9365);
or U12041 (N_12041,N_10080,N_11280);
nor U12042 (N_12042,N_9918,N_10971);
and U12043 (N_12043,N_11677,N_9303);
nor U12044 (N_12044,N_11870,N_9294);
or U12045 (N_12045,N_9438,N_11748);
or U12046 (N_12046,N_10754,N_10750);
nor U12047 (N_12047,N_11903,N_10557);
or U12048 (N_12048,N_11308,N_9609);
or U12049 (N_12049,N_11722,N_11168);
or U12050 (N_12050,N_11576,N_9362);
nand U12051 (N_12051,N_9541,N_11293);
nor U12052 (N_12052,N_9270,N_11800);
xnor U12053 (N_12053,N_11114,N_10715);
nand U12054 (N_12054,N_10532,N_10771);
nor U12055 (N_12055,N_11099,N_11198);
or U12056 (N_12056,N_10358,N_11296);
nor U12057 (N_12057,N_11989,N_9092);
nor U12058 (N_12058,N_10978,N_11478);
or U12059 (N_12059,N_9195,N_9847);
nand U12060 (N_12060,N_9368,N_10156);
nand U12061 (N_12061,N_11826,N_10416);
xnor U12062 (N_12062,N_10632,N_11809);
or U12063 (N_12063,N_11828,N_11090);
and U12064 (N_12064,N_9618,N_11332);
nor U12065 (N_12065,N_9321,N_10697);
nand U12066 (N_12066,N_10101,N_10999);
xor U12067 (N_12067,N_11687,N_9117);
nor U12068 (N_12068,N_11235,N_10252);
nand U12069 (N_12069,N_10986,N_9785);
nor U12070 (N_12070,N_10602,N_9420);
nor U12071 (N_12071,N_10478,N_9780);
and U12072 (N_12072,N_10776,N_11104);
nor U12073 (N_12073,N_10914,N_9258);
xnor U12074 (N_12074,N_9166,N_10558);
and U12075 (N_12075,N_11618,N_11794);
and U12076 (N_12076,N_11141,N_11001);
nor U12077 (N_12077,N_9941,N_9608);
and U12078 (N_12078,N_9613,N_9663);
or U12079 (N_12079,N_10507,N_10471);
nand U12080 (N_12080,N_10816,N_11314);
nor U12081 (N_12081,N_9298,N_9703);
nor U12082 (N_12082,N_9939,N_11372);
and U12083 (N_12083,N_9472,N_11547);
or U12084 (N_12084,N_9480,N_10493);
nand U12085 (N_12085,N_10293,N_10220);
and U12086 (N_12086,N_9306,N_9723);
nor U12087 (N_12087,N_9831,N_9288);
xor U12088 (N_12088,N_10344,N_10887);
or U12089 (N_12089,N_10994,N_11065);
nor U12090 (N_12090,N_9873,N_10721);
or U12091 (N_12091,N_9226,N_9796);
or U12092 (N_12092,N_10212,N_9393);
and U12093 (N_12093,N_9058,N_9494);
nor U12094 (N_12094,N_10906,N_11920);
nor U12095 (N_12095,N_9877,N_11540);
nor U12096 (N_12096,N_10032,N_10320);
nand U12097 (N_12097,N_11191,N_11644);
or U12098 (N_12098,N_9328,N_9192);
nand U12099 (N_12099,N_11475,N_10995);
nor U12100 (N_12100,N_11451,N_10681);
nand U12101 (N_12101,N_10727,N_9081);
xor U12102 (N_12102,N_11325,N_11123);
nand U12103 (N_12103,N_11672,N_10762);
and U12104 (N_12104,N_9084,N_10354);
xor U12105 (N_12105,N_11087,N_10908);
and U12106 (N_12106,N_9361,N_9152);
and U12107 (N_12107,N_10611,N_10938);
and U12108 (N_12108,N_9826,N_10907);
nor U12109 (N_12109,N_11048,N_9811);
or U12110 (N_12110,N_10965,N_9196);
or U12111 (N_12111,N_9187,N_11597);
nand U12112 (N_12112,N_11703,N_11089);
nand U12113 (N_12113,N_10335,N_10133);
or U12114 (N_12114,N_9764,N_10172);
nor U12115 (N_12115,N_9712,N_11390);
or U12116 (N_12116,N_9341,N_9171);
and U12117 (N_12117,N_10426,N_10858);
nand U12118 (N_12118,N_9399,N_10741);
and U12119 (N_12119,N_10548,N_11039);
and U12120 (N_12120,N_11236,N_11689);
and U12121 (N_12121,N_10967,N_11094);
nand U12122 (N_12122,N_10137,N_9370);
nand U12123 (N_12123,N_11831,N_9799);
or U12124 (N_12124,N_9202,N_9211);
nor U12125 (N_12125,N_10187,N_11955);
or U12126 (N_12126,N_9732,N_9366);
xor U12127 (N_12127,N_10264,N_10305);
or U12128 (N_12128,N_9934,N_11237);
xnor U12129 (N_12129,N_11712,N_11768);
nor U12130 (N_12130,N_9520,N_11355);
nor U12131 (N_12131,N_10165,N_9631);
and U12132 (N_12132,N_10545,N_11719);
or U12133 (N_12133,N_10045,N_9350);
and U12134 (N_12134,N_11248,N_9583);
nand U12135 (N_12135,N_9903,N_10217);
nand U12136 (N_12136,N_9175,N_11134);
nand U12137 (N_12137,N_11560,N_9616);
nand U12138 (N_12138,N_10109,N_9997);
nor U12139 (N_12139,N_10631,N_11145);
and U12140 (N_12140,N_11043,N_9035);
xnor U12141 (N_12141,N_10279,N_10328);
and U12142 (N_12142,N_11944,N_10977);
and U12143 (N_12143,N_11652,N_11643);
and U12144 (N_12144,N_9032,N_10788);
nand U12145 (N_12145,N_9463,N_9238);
nand U12146 (N_12146,N_10433,N_11249);
nand U12147 (N_12147,N_10755,N_11889);
nor U12148 (N_12148,N_9881,N_11493);
and U12149 (N_12149,N_11185,N_10227);
nand U12150 (N_12150,N_9369,N_10090);
nor U12151 (N_12151,N_10573,N_11482);
nand U12152 (N_12152,N_9129,N_9809);
nand U12153 (N_12153,N_11812,N_11780);
nor U12154 (N_12154,N_10757,N_10539);
or U12155 (N_12155,N_9228,N_9911);
nand U12156 (N_12156,N_11421,N_9676);
and U12157 (N_12157,N_11461,N_11667);
nor U12158 (N_12158,N_10654,N_9853);
and U12159 (N_12159,N_10694,N_11639);
or U12160 (N_12160,N_10853,N_9557);
nand U12161 (N_12161,N_10719,N_9888);
nand U12162 (N_12162,N_11840,N_11476);
nor U12163 (N_12163,N_11961,N_11170);
or U12164 (N_12164,N_11795,N_9561);
and U12165 (N_12165,N_10331,N_10141);
nor U12166 (N_12166,N_11893,N_9473);
nand U12167 (N_12167,N_11154,N_9006);
or U12168 (N_12168,N_11327,N_11630);
and U12169 (N_12169,N_11147,N_9830);
nor U12170 (N_12170,N_10517,N_9720);
nand U12171 (N_12171,N_11849,N_10083);
and U12172 (N_12172,N_11337,N_10520);
or U12173 (N_12173,N_11788,N_10278);
xor U12174 (N_12174,N_11698,N_11379);
nor U12175 (N_12175,N_11468,N_10093);
and U12176 (N_12176,N_11585,N_11344);
nor U12177 (N_12177,N_11616,N_10854);
nor U12178 (N_12178,N_11439,N_10726);
nand U12179 (N_12179,N_9680,N_9257);
nand U12180 (N_12180,N_9617,N_11601);
nand U12181 (N_12181,N_10556,N_10650);
and U12182 (N_12182,N_9336,N_9833);
nor U12183 (N_12183,N_11910,N_11024);
nor U12184 (N_12184,N_10325,N_9542);
nor U12185 (N_12185,N_9169,N_10889);
or U12186 (N_12186,N_11947,N_11077);
or U12187 (N_12187,N_11085,N_10886);
or U12188 (N_12188,N_9414,N_9668);
nand U12189 (N_12189,N_11657,N_11956);
nor U12190 (N_12190,N_11031,N_10525);
and U12191 (N_12191,N_11251,N_9545);
xor U12192 (N_12192,N_10379,N_11362);
xor U12193 (N_12193,N_11142,N_9926);
or U12194 (N_12194,N_9223,N_11388);
and U12195 (N_12195,N_9669,N_9790);
nand U12196 (N_12196,N_11462,N_9020);
or U12197 (N_12197,N_10114,N_9709);
nor U12198 (N_12198,N_9858,N_11874);
or U12199 (N_12199,N_11149,N_9586);
nand U12200 (N_12200,N_9064,N_11965);
nand U12201 (N_12201,N_10249,N_9610);
nor U12202 (N_12202,N_11161,N_10054);
nor U12203 (N_12203,N_9793,N_11226);
nand U12204 (N_12204,N_10929,N_10300);
and U12205 (N_12205,N_11017,N_9897);
nor U12206 (N_12206,N_11858,N_10782);
or U12207 (N_12207,N_11628,N_10541);
and U12208 (N_12208,N_9572,N_11307);
xnor U12209 (N_12209,N_10457,N_10559);
and U12210 (N_12210,N_9424,N_10489);
nand U12211 (N_12211,N_11726,N_9003);
nand U12212 (N_12212,N_9466,N_9379);
or U12213 (N_12213,N_11025,N_10255);
xnor U12214 (N_12214,N_10138,N_10823);
and U12215 (N_12215,N_10871,N_9971);
or U12216 (N_12216,N_9671,N_11897);
and U12217 (N_12217,N_11931,N_11431);
and U12218 (N_12218,N_9803,N_11028);
and U12219 (N_12219,N_9046,N_11864);
nand U12220 (N_12220,N_11533,N_10961);
or U12221 (N_12221,N_9124,N_10553);
or U12222 (N_12222,N_9415,N_10928);
nand U12223 (N_12223,N_11650,N_11815);
xnor U12224 (N_12224,N_11736,N_11009);
and U12225 (N_12225,N_10505,N_11295);
nand U12226 (N_12226,N_11756,N_10496);
nor U12227 (N_12227,N_10304,N_10461);
nand U12228 (N_12228,N_10732,N_10794);
nor U12229 (N_12229,N_11448,N_10449);
and U12230 (N_12230,N_10913,N_10501);
or U12231 (N_12231,N_10926,N_10306);
or U12232 (N_12232,N_11347,N_10572);
or U12233 (N_12233,N_10565,N_10261);
nor U12234 (N_12234,N_11358,N_10506);
nor U12235 (N_12235,N_9677,N_9318);
and U12236 (N_12236,N_10462,N_9885);
and U12237 (N_12237,N_10295,N_9607);
nand U12238 (N_12238,N_11323,N_10890);
and U12239 (N_12239,N_9157,N_9286);
nor U12240 (N_12240,N_11410,N_9025);
nand U12241 (N_12241,N_9797,N_10659);
nand U12242 (N_12242,N_9731,N_10529);
nor U12243 (N_12243,N_11240,N_9951);
xnor U12244 (N_12244,N_11040,N_10567);
nand U12245 (N_12245,N_10134,N_11823);
nor U12246 (N_12246,N_10594,N_11329);
nor U12247 (N_12247,N_11357,N_10185);
and U12248 (N_12248,N_9711,N_9183);
or U12249 (N_12249,N_11591,N_11139);
and U12250 (N_12250,N_11239,N_11341);
nand U12251 (N_12251,N_9437,N_10330);
nand U12252 (N_12252,N_9821,N_9390);
nand U12253 (N_12253,N_10096,N_10934);
nor U12254 (N_12254,N_10065,N_11749);
or U12255 (N_12255,N_9267,N_10235);
and U12256 (N_12256,N_11203,N_11289);
xnor U12257 (N_12257,N_10383,N_11488);
or U12258 (N_12258,N_10515,N_10346);
and U12259 (N_12259,N_11682,N_10375);
or U12260 (N_12260,N_9241,N_9577);
or U12261 (N_12261,N_11019,N_11381);
or U12262 (N_12262,N_10476,N_10680);
or U12263 (N_12263,N_10604,N_11232);
nor U12264 (N_12264,N_10148,N_10877);
nor U12265 (N_12265,N_9304,N_9315);
or U12266 (N_12266,N_10174,N_11817);
or U12267 (N_12267,N_10991,N_11531);
or U12268 (N_12268,N_11896,N_11924);
nand U12269 (N_12269,N_9217,N_9330);
or U12270 (N_12270,N_9180,N_9639);
nand U12271 (N_12271,N_11177,N_11589);
xnor U12272 (N_12272,N_10244,N_11465);
nor U12273 (N_12273,N_11003,N_11036);
nor U12274 (N_12274,N_11503,N_11411);
xnor U12275 (N_12275,N_10523,N_10297);
or U12276 (N_12276,N_11467,N_10152);
nand U12277 (N_12277,N_9846,N_11284);
xnor U12278 (N_12278,N_10960,N_10372);
nor U12279 (N_12279,N_11975,N_10368);
nand U12280 (N_12280,N_10531,N_10921);
and U12281 (N_12281,N_11026,N_9491);
nand U12282 (N_12282,N_11497,N_9173);
nor U12283 (N_12283,N_10899,N_9702);
or U12284 (N_12284,N_10091,N_11885);
nor U12285 (N_12285,N_10625,N_11157);
nor U12286 (N_12286,N_9271,N_9701);
and U12287 (N_12287,N_11258,N_10147);
xor U12288 (N_12288,N_9445,N_9102);
nand U12289 (N_12289,N_10840,N_11769);
nand U12290 (N_12290,N_10648,N_10466);
or U12291 (N_12291,N_9573,N_11098);
nand U12292 (N_12292,N_11522,N_10497);
nand U12293 (N_12293,N_11030,N_10922);
nor U12294 (N_12294,N_11244,N_11304);
nor U12295 (N_12295,N_9518,N_9292);
and U12296 (N_12296,N_11539,N_9194);
or U12297 (N_12297,N_9584,N_10470);
and U12298 (N_12298,N_10287,N_9347);
xnor U12299 (N_12299,N_11988,N_9506);
and U12300 (N_12300,N_11750,N_9970);
or U12301 (N_12301,N_10561,N_11396);
and U12302 (N_12302,N_10009,N_11612);
nor U12303 (N_12303,N_9485,N_11869);
nand U12304 (N_12304,N_11061,N_9028);
nor U12305 (N_12305,N_11755,N_11778);
or U12306 (N_12306,N_11427,N_10740);
xor U12307 (N_12307,N_11441,N_11658);
nand U12308 (N_12308,N_9387,N_11434);
xor U12309 (N_12309,N_11480,N_11268);
or U12310 (N_12310,N_11369,N_11838);
nand U12311 (N_12311,N_11211,N_9932);
and U12312 (N_12312,N_10294,N_10714);
nand U12313 (N_12313,N_9052,N_9191);
or U12314 (N_12314,N_11015,N_10224);
or U12315 (N_12315,N_11895,N_9981);
nor U12316 (N_12316,N_11888,N_10369);
and U12317 (N_12317,N_9508,N_11338);
and U12318 (N_12318,N_11603,N_10809);
or U12319 (N_12319,N_11510,N_9080);
nand U12320 (N_12320,N_10870,N_10046);
or U12321 (N_12321,N_11799,N_10425);
or U12322 (N_12322,N_10350,N_11352);
nand U12323 (N_12323,N_9276,N_10064);
nor U12324 (N_12324,N_11514,N_10464);
nand U12325 (N_12325,N_11620,N_9458);
nand U12326 (N_12326,N_9496,N_9637);
and U12327 (N_12327,N_9013,N_9956);
or U12328 (N_12328,N_10535,N_10958);
nor U12329 (N_12329,N_10215,N_10073);
or U12330 (N_12330,N_10381,N_9523);
or U12331 (N_12331,N_10730,N_10323);
or U12332 (N_12332,N_10711,N_9045);
nand U12333 (N_12333,N_10199,N_10316);
nor U12334 (N_12334,N_10108,N_9786);
nor U12335 (N_12335,N_10208,N_10500);
and U12336 (N_12336,N_10736,N_9229);
nand U12337 (N_12337,N_10966,N_11286);
and U12338 (N_12338,N_11534,N_10670);
and U12339 (N_12339,N_10514,N_10789);
nor U12340 (N_12340,N_10831,N_10124);
nand U12341 (N_12341,N_11136,N_10665);
or U12342 (N_12342,N_9487,N_10445);
or U12343 (N_12343,N_9788,N_10472);
or U12344 (N_12344,N_9957,N_9733);
or U12345 (N_12345,N_9478,N_10393);
nand U12346 (N_12346,N_10980,N_11773);
and U12347 (N_12347,N_10078,N_10098);
or U12348 (N_12348,N_10498,N_9208);
nand U12349 (N_12349,N_10709,N_9820);
or U12350 (N_12350,N_9209,N_11970);
nor U12351 (N_12351,N_9834,N_9116);
and U12352 (N_12352,N_9683,N_11671);
nand U12353 (N_12353,N_11285,N_10544);
nand U12354 (N_12354,N_10062,N_10382);
or U12355 (N_12355,N_10568,N_10438);
nor U12356 (N_12356,N_10336,N_9367);
nand U12357 (N_12357,N_11222,N_10403);
nand U12358 (N_12358,N_11876,N_9470);
nor U12359 (N_12359,N_10251,N_9930);
xnor U12360 (N_12360,N_9296,N_10319);
nand U12361 (N_12361,N_11695,N_10280);
nor U12362 (N_12362,N_11260,N_11595);
or U12363 (N_12363,N_11496,N_11886);
or U12364 (N_12364,N_10605,N_9299);
nand U12365 (N_12365,N_10432,N_11538);
or U12366 (N_12366,N_9823,N_10552);
xnor U12367 (N_12367,N_11267,N_10821);
nand U12368 (N_12368,N_11117,N_11761);
nor U12369 (N_12369,N_9356,N_11706);
and U12370 (N_12370,N_11453,N_10662);
or U12371 (N_12371,N_11571,N_9378);
nor U12372 (N_12372,N_10089,N_9091);
xnor U12373 (N_12373,N_11899,N_9908);
nor U12374 (N_12374,N_9757,N_10164);
nand U12375 (N_12375,N_9040,N_10576);
and U12376 (N_12376,N_10269,N_10677);
and U12377 (N_12377,N_10190,N_11545);
nand U12378 (N_12378,N_9449,N_9978);
xnor U12379 (N_12379,N_9079,N_11452);
and U12380 (N_12380,N_11743,N_11629);
and U12381 (N_12381,N_11941,N_9138);
or U12382 (N_12382,N_9581,N_9314);
nand U12383 (N_12383,N_10895,N_10233);
nand U12384 (N_12384,N_11623,N_10790);
and U12385 (N_12385,N_11716,N_11680);
xnor U12386 (N_12386,N_9504,N_11300);
nor U12387 (N_12387,N_11807,N_11673);
and U12388 (N_12388,N_9495,N_11816);
nand U12389 (N_12389,N_9685,N_11604);
or U12390 (N_12390,N_11907,N_11298);
xnor U12391 (N_12391,N_10214,N_9556);
nand U12392 (N_12392,N_11766,N_9986);
xor U12393 (N_12393,N_11076,N_10849);
or U12394 (N_12394,N_9570,N_10198);
nor U12395 (N_12395,N_10852,N_11386);
or U12396 (N_12396,N_9620,N_11106);
nand U12397 (N_12397,N_11062,N_9710);
nor U12398 (N_12398,N_10982,N_11103);
or U12399 (N_12399,N_10104,N_10006);
nand U12400 (N_12400,N_10935,N_9900);
nand U12401 (N_12401,N_9651,N_10522);
nor U12402 (N_12402,N_10981,N_10752);
nand U12403 (N_12403,N_11072,N_9687);
nor U12404 (N_12404,N_10226,N_11608);
and U12405 (N_12405,N_9975,N_10247);
nand U12406 (N_12406,N_10389,N_11501);
or U12407 (N_12407,N_11813,N_9384);
nand U12408 (N_12408,N_9312,N_9513);
nand U12409 (N_12409,N_9522,N_9598);
and U12410 (N_12410,N_11884,N_9658);
or U12411 (N_12411,N_10160,N_11209);
nand U12412 (N_12412,N_11745,N_9098);
nor U12413 (N_12413,N_11909,N_11105);
and U12414 (N_12414,N_11206,N_9634);
nor U12415 (N_12415,N_11050,N_11567);
or U12416 (N_12416,N_10878,N_10271);
or U12417 (N_12417,N_10942,N_9746);
nand U12418 (N_12418,N_9666,N_10924);
nand U12419 (N_12419,N_9022,N_10893);
and U12420 (N_12420,N_10804,N_9726);
nor U12421 (N_12421,N_11617,N_11697);
nand U12422 (N_12422,N_10598,N_9805);
nor U12423 (N_12423,N_9579,N_9139);
or U12424 (N_12424,N_11368,N_11977);
nand U12425 (N_12425,N_10024,N_10661);
or U12426 (N_12426,N_9898,N_10972);
and U12427 (N_12427,N_10050,N_10276);
nor U12428 (N_12428,N_11356,N_10392);
or U12429 (N_12429,N_11744,N_11517);
nor U12430 (N_12430,N_10990,N_9212);
nand U12431 (N_12431,N_9319,N_10092);
and U12432 (N_12432,N_9467,N_11912);
and U12433 (N_12433,N_9931,N_10792);
nand U12434 (N_12434,N_11887,N_10467);
nand U12435 (N_12435,N_10097,N_9146);
nor U12436 (N_12436,N_11423,N_11197);
xor U12437 (N_12437,N_9812,N_10491);
nor U12438 (N_12438,N_9429,N_10210);
nand U12439 (N_12439,N_11445,N_9235);
nand U12440 (N_12440,N_10760,N_11696);
nand U12441 (N_12441,N_9452,N_11607);
nand U12442 (N_12442,N_11187,N_10408);
nand U12443 (N_12443,N_10808,N_10314);
or U12444 (N_12444,N_10191,N_9255);
or U12445 (N_12445,N_11231,N_11966);
nor U12446 (N_12446,N_10728,N_9088);
nand U12447 (N_12447,N_9887,N_9309);
or U12448 (N_12448,N_10970,N_11638);
and U12449 (N_12449,N_11500,N_9612);
and U12450 (N_12450,N_11688,N_10613);
nand U12451 (N_12451,N_11370,N_11982);
or U12452 (N_12452,N_10746,N_10458);
and U12453 (N_12453,N_9263,N_10894);
or U12454 (N_12454,N_9679,N_9546);
xnor U12455 (N_12455,N_11569,N_9442);
and U12456 (N_12456,N_9451,N_9069);
nand U12457 (N_12457,N_10371,N_11536);
and U12458 (N_12458,N_11395,N_10820);
or U12459 (N_12459,N_9653,N_11186);
nor U12460 (N_12460,N_10504,N_9737);
nor U12461 (N_12461,N_9724,N_10299);
xor U12462 (N_12462,N_9543,N_11714);
nor U12463 (N_12463,N_10463,N_9027);
and U12464 (N_12464,N_10061,N_10434);
nor U12465 (N_12465,N_10429,N_10891);
or U12466 (N_12466,N_11430,N_11287);
or U12467 (N_12467,N_10150,N_10881);
and U12468 (N_12468,N_11986,N_9264);
or U12469 (N_12469,N_11302,N_11605);
nor U12470 (N_12470,N_10231,N_9179);
nand U12471 (N_12471,N_10581,N_10333);
nor U12472 (N_12472,N_9394,N_10232);
xnor U12473 (N_12473,N_9562,N_9596);
nand U12474 (N_12474,N_11233,N_11751);
and U12475 (N_12475,N_11692,N_9946);
nor U12476 (N_12476,N_10259,N_9441);
xor U12477 (N_12477,N_9422,N_10976);
and U12478 (N_12478,N_11526,N_10321);
nand U12479 (N_12479,N_10574,N_11096);
nand U12480 (N_12480,N_10340,N_11055);
and U12481 (N_12481,N_9991,N_9053);
nand U12482 (N_12482,N_10118,N_11400);
or U12483 (N_12483,N_11913,N_9973);
nand U12484 (N_12484,N_10855,N_11575);
and U12485 (N_12485,N_10571,N_11389);
xor U12486 (N_12486,N_9961,N_11270);
and U12487 (N_12487,N_9874,N_11363);
xor U12488 (N_12488,N_10518,N_11179);
or U12489 (N_12489,N_9435,N_9029);
xnor U12490 (N_12490,N_10710,N_9459);
nor U12491 (N_12491,N_9085,N_9632);
and U12492 (N_12492,N_11262,N_10699);
and U12493 (N_12493,N_9086,N_9159);
or U12494 (N_12494,N_11727,N_10813);
nor U12495 (N_12495,N_11006,N_11406);
nor U12496 (N_12496,N_10242,N_9210);
nor U12497 (N_12497,N_11360,N_9963);
and U12498 (N_12498,N_10339,N_10052);
and U12499 (N_12499,N_11731,N_10483);
nor U12500 (N_12500,N_9331,N_9260);
nand U12501 (N_12501,N_10737,N_9057);
nor U12502 (N_12502,N_9996,N_11700);
nor U12503 (N_12503,N_9642,N_10860);
xnor U12504 (N_12504,N_9924,N_11306);
and U12505 (N_12505,N_9625,N_11660);
or U12506 (N_12506,N_11715,N_11340);
or U12507 (N_12507,N_9503,N_10801);
nand U12508 (N_12508,N_11824,N_11960);
nand U12509 (N_12509,N_9528,N_10044);
nor U12510 (N_12510,N_10051,N_11980);
and U12511 (N_12511,N_10384,N_9411);
nand U12512 (N_12512,N_9386,N_9167);
nand U12513 (N_12513,N_11917,N_11776);
nor U12514 (N_12514,N_10872,N_11967);
and U12515 (N_12515,N_10386,N_10984);
nor U12516 (N_12516,N_10812,N_11188);
and U12517 (N_12517,N_10034,N_9240);
nor U12518 (N_12518,N_10550,N_11053);
nand U12519 (N_12519,N_10674,N_9363);
and U12520 (N_12520,N_9601,N_9061);
nor U12521 (N_12521,N_9033,N_11163);
and U12522 (N_12522,N_9421,N_10189);
and U12523 (N_12523,N_9216,N_10705);
or U12524 (N_12524,N_9933,N_10769);
nand U12525 (N_12525,N_9443,N_9962);
xnor U12526 (N_12526,N_11738,N_9706);
nand U12527 (N_12527,N_9048,N_10480);
xnor U12528 (N_12528,N_10207,N_9814);
or U12529 (N_12529,N_11927,N_11730);
xnor U12530 (N_12530,N_10621,N_9010);
or U12531 (N_12531,N_11541,N_9071);
and U12532 (N_12532,N_9501,N_11092);
nor U12533 (N_12533,N_10318,N_10646);
or U12534 (N_12534,N_11278,N_9070);
xor U12535 (N_12535,N_10658,N_9870);
nand U12536 (N_12536,N_9126,N_11290);
nand U12537 (N_12537,N_11084,N_10919);
nor U12538 (N_12538,N_11635,N_10793);
nor U12539 (N_12539,N_11733,N_11227);
or U12540 (N_12540,N_9089,N_11119);
nand U12541 (N_12541,N_9324,N_11580);
nor U12542 (N_12542,N_9714,N_11212);
nor U12543 (N_12543,N_10007,N_9310);
xnor U12544 (N_12544,N_9334,N_9246);
xnor U12545 (N_12545,N_9431,N_11704);
nand U12546 (N_12546,N_9657,N_9385);
and U12547 (N_12547,N_10842,N_11494);
or U12548 (N_12548,N_9564,N_9742);
and U12549 (N_12549,N_10363,N_9254);
and U12550 (N_12550,N_11848,N_11221);
and U12551 (N_12551,N_9966,N_10647);
or U12552 (N_12552,N_9498,N_11747);
nand U12553 (N_12553,N_10312,N_9725);
or U12554 (N_12554,N_9974,N_10365);
nand U12555 (N_12555,N_9947,N_9927);
nand U12556 (N_12556,N_9377,N_10651);
nor U12557 (N_12557,N_11821,N_9912);
and U12558 (N_12558,N_9787,N_9575);
nor U12559 (N_12559,N_11521,N_9252);
or U12560 (N_12560,N_9882,N_9130);
nand U12561 (N_12561,N_9624,N_9824);
or U12562 (N_12562,N_10263,N_11959);
or U12563 (N_12563,N_9836,N_10357);
xor U12564 (N_12564,N_11862,N_11064);
and U12565 (N_12565,N_10376,N_9450);
and U12566 (N_12566,N_11190,N_11587);
or U12567 (N_12567,N_10015,N_10690);
xor U12568 (N_12568,N_10839,N_9699);
nand U12569 (N_12569,N_9261,N_11929);
nor U12570 (N_12570,N_9177,N_9340);
nor U12571 (N_12571,N_10370,N_11277);
or U12572 (N_12572,N_10707,N_11984);
nand U12573 (N_12573,N_10502,N_11490);
xnor U12574 (N_12574,N_10112,N_10837);
and U12575 (N_12575,N_11107,N_11225);
nand U12576 (N_12576,N_9705,N_11842);
nor U12577 (N_12577,N_10620,N_9308);
xor U12578 (N_12578,N_10201,N_9433);
nand U12579 (N_12579,N_9397,N_10008);
nor U12580 (N_12580,N_10402,N_9511);
nand U12581 (N_12581,N_11444,N_10237);
nor U12582 (N_12582,N_10380,N_10968);
nand U12583 (N_12583,N_10026,N_9256);
or U12584 (N_12584,N_11169,N_9067);
and U12585 (N_12585,N_10560,N_11419);
and U12586 (N_12586,N_9794,N_9244);
nor U12587 (N_12587,N_9410,N_10268);
nand U12588 (N_12588,N_11495,N_10784);
xnor U12589 (N_12589,N_9735,N_10927);
xor U12590 (N_12590,N_11511,N_11563);
nand U12591 (N_12591,N_11566,N_10937);
nor U12592 (N_12592,N_9313,N_10687);
nand U12593 (N_12593,N_9675,N_9630);
and U12594 (N_12594,N_11837,N_10166);
and U12595 (N_12595,N_11872,N_9510);
nand U12596 (N_12596,N_10920,N_9342);
or U12597 (N_12597,N_10626,N_9000);
nor U12598 (N_12598,N_10592,N_9585);
and U12599 (N_12599,N_10151,N_10103);
and U12600 (N_12600,N_11063,N_11998);
xor U12601 (N_12601,N_9749,N_11269);
or U12602 (N_12602,N_10192,N_9358);
or U12603 (N_12603,N_9619,N_9859);
nand U12604 (N_12604,N_9905,N_9206);
and U12605 (N_12605,N_9615,N_9481);
nand U12606 (N_12606,N_10667,N_11305);
nor U12607 (N_12607,N_9552,N_9896);
xnor U12608 (N_12608,N_10685,N_11825);
nor U12609 (N_12609,N_9643,N_11112);
and U12610 (N_12610,N_10448,N_9444);
and U12611 (N_12611,N_9305,N_11487);
xor U12612 (N_12612,N_11655,N_9999);
and U12613 (N_12613,N_10406,N_9479);
nand U12614 (N_12614,N_11075,N_9036);
nor U12615 (N_12615,N_11246,N_9760);
and U12616 (N_12616,N_11380,N_9417);
nor U12617 (N_12617,N_11250,N_11456);
and U12618 (N_12618,N_9977,N_10218);
nand U12619 (N_12619,N_11904,N_11611);
nand U12620 (N_12620,N_9739,N_11969);
nor U12621 (N_12621,N_11259,N_9333);
or U12622 (N_12622,N_9134,N_11382);
and U12623 (N_12623,N_10394,N_11130);
nor U12624 (N_12624,N_11771,N_11868);
xor U12625 (N_12625,N_9646,N_9004);
nor U12626 (N_12626,N_9916,N_11489);
nand U12627 (N_12627,N_10186,N_11523);
and U12628 (N_12628,N_11402,N_11619);
nand U12629 (N_12629,N_11691,N_9761);
and U12630 (N_12630,N_9059,N_10035);
nor U12631 (N_12631,N_11707,N_10791);
nand U12632 (N_12632,N_9555,N_10623);
nor U12633 (N_12633,N_10575,N_10143);
or U12634 (N_12634,N_10364,N_9548);
nor U12635 (N_12635,N_9227,N_9178);
or U12636 (N_12636,N_11027,N_11156);
or U12637 (N_12637,N_9734,N_9863);
and U12638 (N_12638,N_11255,N_10723);
and U12639 (N_12639,N_10807,N_11202);
or U12640 (N_12640,N_9284,N_11850);
or U12641 (N_12641,N_10175,N_10817);
and U12642 (N_12642,N_10443,N_10485);
or U12643 (N_12643,N_9549,N_10596);
nand U12644 (N_12644,N_10374,N_11785);
nor U12645 (N_12645,N_9536,N_9477);
nand U12646 (N_12646,N_9490,N_10033);
nand U12647 (N_12647,N_9147,N_10136);
nor U12648 (N_12648,N_11624,N_9185);
nor U12649 (N_12649,N_11449,N_9594);
or U12650 (N_12650,N_10417,N_11220);
nand U12651 (N_12651,N_11046,N_9582);
nand U12652 (N_12652,N_9408,N_11670);
or U12653 (N_12653,N_10473,N_11832);
nand U12654 (N_12654,N_9728,N_9835);
or U12655 (N_12655,N_9722,N_9297);
or U12656 (N_12656,N_10985,N_10952);
nand U12657 (N_12657,N_10660,N_9274);
nand U12658 (N_12658,N_10859,N_11012);
nand U12659 (N_12659,N_11625,N_10818);
nand U12660 (N_12660,N_11365,N_10917);
nand U12661 (N_12661,N_9242,N_10939);
nand U12662 (N_12662,N_11574,N_9985);
xnor U12663 (N_12663,N_11873,N_9563);
xnor U12664 (N_12664,N_10633,N_9289);
nor U12665 (N_12665,N_10954,N_10437);
nor U12666 (N_12666,N_9285,N_9024);
or U12667 (N_12667,N_11317,N_11935);
nand U12668 (N_12668,N_10989,N_11765);
or U12669 (N_12669,N_10284,N_10144);
and U12670 (N_12670,N_9182,N_11925);
xnor U12671 (N_12671,N_11757,N_11649);
and U12672 (N_12672,N_10686,N_11000);
and U12673 (N_12673,N_9681,N_11189);
or U12674 (N_12674,N_9248,N_9694);
and U12675 (N_12675,N_11180,N_9649);
xor U12676 (N_12676,N_9295,N_10885);
nand U12677 (N_12677,N_11086,N_11708);
nor U12678 (N_12678,N_10282,N_9143);
nand U12679 (N_12679,N_10799,N_10456);
nor U12680 (N_12680,N_10861,N_11529);
nor U12681 (N_12681,N_11109,N_9137);
nand U12682 (N_12682,N_11772,N_11590);
nor U12683 (N_12683,N_9695,N_10486);
xor U12684 (N_12684,N_10749,N_10524);
and U12685 (N_12685,N_10689,N_9660);
nor U12686 (N_12686,N_11647,N_9259);
nor U12687 (N_12687,N_9489,N_9214);
and U12688 (N_12688,N_10618,N_10963);
nand U12689 (N_12689,N_9762,N_10196);
nor U12690 (N_12690,N_9453,N_10814);
or U12691 (N_12691,N_11763,N_11843);
nand U12692 (N_12692,N_11181,N_11095);
nand U12693 (N_12693,N_11551,N_11299);
and U12694 (N_12694,N_9635,N_9120);
xor U12695 (N_12695,N_9364,N_9770);
nor U12696 (N_12696,N_11173,N_10542);
nand U12697 (N_12697,N_11309,N_9837);
nand U12698 (N_12698,N_11860,N_11732);
nand U12699 (N_12699,N_9987,N_10225);
or U12700 (N_12700,N_10428,N_10634);
or U12701 (N_12701,N_10036,N_11646);
or U12702 (N_12702,N_11922,N_11120);
nand U12703 (N_12703,N_11052,N_10367);
nand U12704 (N_12704,N_11686,N_10716);
nor U12705 (N_12705,N_10349,N_9266);
and U12706 (N_12706,N_10987,N_9193);
nor U12707 (N_12707,N_9633,N_11640);
nand U12708 (N_12708,N_10058,N_11957);
or U12709 (N_12709,N_10758,N_11132);
nand U12710 (N_12710,N_9592,N_10761);
or U12711 (N_12711,N_9281,N_11991);
and U12712 (N_12712,N_11535,N_9696);
or U12713 (N_12713,N_10135,N_11822);
nand U12714 (N_12714,N_10583,N_11199);
nand U12715 (N_12715,N_9108,N_10020);
or U12716 (N_12716,N_9854,N_11010);
nor U12717 (N_12717,N_10759,N_10586);
and U12718 (N_12718,N_10311,N_10768);
or U12719 (N_12719,N_10802,N_10281);
nor U12720 (N_12720,N_10447,N_9409);
nor U12721 (N_12721,N_11178,N_9034);
and U12722 (N_12722,N_11542,N_10998);
or U12723 (N_12723,N_10351,N_9959);
nand U12724 (N_12724,N_10979,N_10643);
or U12725 (N_12725,N_10796,N_9533);
xnor U12726 (N_12726,N_11932,N_9428);
nor U12727 (N_12727,N_10943,N_11845);
and U12728 (N_12728,N_10892,N_9993);
nand U12729 (N_12729,N_10722,N_11515);
nand U12730 (N_12730,N_11952,N_11737);
xor U12731 (N_12731,N_11626,N_11328);
nor U12732 (N_12732,N_11948,N_9776);
and U12733 (N_12733,N_9090,N_9909);
nand U12734 (N_12734,N_10785,N_9919);
and U12735 (N_12735,N_9754,N_11930);
nor U12736 (N_12736,N_9647,N_10642);
xnor U12737 (N_12737,N_11364,N_10847);
and U12738 (N_12738,N_10203,N_11463);
and U12739 (N_12739,N_11979,N_10862);
or U12740 (N_12740,N_11792,N_11324);
nor U12741 (N_12741,N_9106,N_10780);
and U12742 (N_12742,N_11167,N_10037);
or U12743 (N_12743,N_9576,N_9636);
and U12744 (N_12744,N_11405,N_10366);
nand U12745 (N_12745,N_9516,N_9767);
and U12746 (N_12746,N_11808,N_9894);
nor U12747 (N_12747,N_9448,N_9174);
nor U12748 (N_12748,N_9895,N_10413);
or U12749 (N_12749,N_9950,N_9645);
xor U12750 (N_12750,N_11034,N_9163);
and U12751 (N_12751,N_11228,N_11450);
nand U12752 (N_12752,N_10100,N_9332);
nand U12753 (N_12753,N_9804,N_11333);
and U12754 (N_12754,N_10857,N_11676);
nand U12755 (N_12755,N_11224,N_10733);
nor U12756 (N_12756,N_9872,N_11990);
nand U12757 (N_12757,N_9818,N_11252);
nor U12758 (N_12758,N_9560,N_11584);
or U12759 (N_12759,N_11088,N_10549);
nor U12760 (N_12760,N_10031,N_9031);
nand U12761 (N_12761,N_11108,N_10419);
xnor U12762 (N_12762,N_9829,N_10213);
nor U12763 (N_12763,N_11118,N_9886);
nand U12764 (N_12764,N_10409,N_9160);
nor U12765 (N_12765,N_10418,N_9078);
nand U12766 (N_12766,N_10778,N_11319);
or U12767 (N_12767,N_10543,N_10822);
nand U12768 (N_12768,N_11637,N_9407);
nor U12769 (N_12769,N_9967,N_11469);
or U12770 (N_12770,N_11022,N_10718);
and U12771 (N_12771,N_11477,N_10649);
and U12772 (N_12772,N_11158,N_10027);
or U12773 (N_12773,N_10452,N_11742);
and U12774 (N_12774,N_9775,N_9502);
nand U12775 (N_12775,N_10657,N_11294);
xnor U12776 (N_12776,N_10307,N_9401);
or U12777 (N_12777,N_10534,N_11415);
xor U12778 (N_12778,N_10074,N_10038);
or U12779 (N_12779,N_10444,N_9692);
nand U12780 (N_12780,N_11263,N_9468);
nand U12781 (N_12781,N_10183,N_9396);
and U12782 (N_12782,N_11192,N_10002);
nor U12783 (N_12783,N_10302,N_9938);
or U12784 (N_12784,N_11457,N_11393);
and U12785 (N_12785,N_11651,N_9540);
or U12786 (N_12786,N_11656,N_11210);
and U12787 (N_12787,N_10725,N_11124);
xnor U12788 (N_12788,N_10125,N_9097);
nor U12789 (N_12789,N_11717,N_11777);
or U12790 (N_12790,N_11532,N_11424);
or U12791 (N_12791,N_11753,N_11350);
and U12792 (N_12792,N_9599,N_10608);
nand U12793 (N_12793,N_10763,N_10117);
xnor U12794 (N_12794,N_10513,N_10411);
nand U12795 (N_12795,N_9083,N_10169);
and U12796 (N_12796,N_9525,N_11033);
and U12797 (N_12797,N_11374,N_9906);
xor U12798 (N_12798,N_9604,N_9741);
nor U12799 (N_12799,N_10115,N_10579);
or U12800 (N_12800,N_9672,N_10744);
nor U12801 (N_12801,N_11746,N_9375);
nand U12802 (N_12802,N_11900,N_9861);
or U12803 (N_12803,N_9145,N_11974);
and U12804 (N_12804,N_11016,N_9247);
nand U12805 (N_12805,N_11416,N_9716);
or U12806 (N_12806,N_11499,N_10806);
and U12807 (N_12807,N_9151,N_11811);
or U12808 (N_12808,N_9606,N_9382);
nand U12809 (N_12809,N_10679,N_9883);
or U12810 (N_12810,N_11455,N_11829);
nand U12811 (N_12811,N_9515,N_10729);
or U12812 (N_12812,N_11041,N_9005);
nor U12813 (N_12813,N_9447,N_10077);
nand U12814 (N_12814,N_11506,N_9795);
nand U12815 (N_12815,N_11537,N_9641);
and U12816 (N_12816,N_11091,N_9935);
xnor U12817 (N_12817,N_11890,N_9611);
nor U12818 (N_12818,N_9427,N_9800);
nand U12819 (N_12819,N_10155,N_11417);
and U12820 (N_12820,N_11425,N_9654);
nor U12821 (N_12821,N_11383,N_11351);
nand U12822 (N_12822,N_11678,N_11371);
nor U12823 (N_12823,N_10149,N_9103);
and U12824 (N_12824,N_10094,N_11473);
and U12825 (N_12825,N_9250,N_11339);
and U12826 (N_12826,N_10167,N_10084);
nand U12827 (N_12827,N_11083,N_10863);
or U12828 (N_12828,N_11122,N_11852);
nand U12829 (N_12829,N_10315,N_10014);
and U12830 (N_12830,N_9075,N_11994);
and U12831 (N_12831,N_9042,N_10829);
nand U12832 (N_12832,N_9355,N_11614);
nand U12833 (N_12833,N_11943,N_9721);
nand U12834 (N_12834,N_10180,N_10329);
nand U12835 (N_12835,N_10833,N_9073);
and U12836 (N_12836,N_11830,N_10775);
or U12837 (N_12837,N_10347,N_11786);
xnor U12838 (N_12838,N_10345,N_10337);
nand U12839 (N_12839,N_10326,N_10378);
nand U12840 (N_12840,N_9110,N_9162);
nand U12841 (N_12841,N_10277,N_11121);
xor U12842 (N_12842,N_11038,N_10257);
nor U12843 (N_12843,N_11291,N_9980);
nor U12844 (N_12844,N_10404,N_10069);
xnor U12845 (N_12845,N_10488,N_11818);
nor U12846 (N_12846,N_9100,N_9943);
and U12847 (N_12847,N_10262,N_9290);
and U12848 (N_12848,N_9142,N_10835);
nor U12849 (N_12849,N_9287,N_11833);
nand U12850 (N_12850,N_10421,N_9026);
nand U12851 (N_12851,N_9469,N_11435);
and U12852 (N_12852,N_10359,N_9852);
xnor U12853 (N_12853,N_10011,N_11437);
nor U12854 (N_12854,N_10388,N_10825);
or U12855 (N_12855,N_9713,N_9253);
and U12856 (N_12856,N_10322,N_11681);
nand U12857 (N_12857,N_11583,N_10962);
or U12858 (N_12858,N_10400,N_10540);
or U12859 (N_12859,N_11546,N_9150);
nand U12860 (N_12860,N_10765,N_10446);
or U12861 (N_12861,N_10909,N_10170);
nand U12862 (N_12862,N_11964,N_9815);
nor U12863 (N_12863,N_11550,N_11343);
nand U12864 (N_12864,N_9530,N_9659);
nor U12865 (N_12865,N_11422,N_11641);
nand U12866 (N_12866,N_11021,N_10010);
xor U12867 (N_12867,N_10587,N_11555);
nand U12868 (N_12868,N_11728,N_10195);
nand U12869 (N_12869,N_10260,N_9153);
nand U12870 (N_12870,N_10200,N_9914);
or U12871 (N_12871,N_9307,N_9763);
or U12872 (N_12872,N_9249,N_10675);
nand U12873 (N_12873,N_10916,N_9360);
and U12874 (N_12874,N_10075,N_9664);
nor U12875 (N_12875,N_10479,N_11216);
and U12876 (N_12876,N_11946,N_9380);
nor U12877 (N_12877,N_10883,N_9021);
or U12878 (N_12878,N_10272,N_9603);
and U12879 (N_12879,N_11675,N_10795);
or U12880 (N_12880,N_10590,N_9779);
or U12881 (N_12881,N_9055,N_10275);
nor U12882 (N_12882,N_9844,N_10387);
and U12883 (N_12883,N_11805,N_9689);
nor U12884 (N_12884,N_11253,N_9337);
xnor U12885 (N_12885,N_10188,N_9500);
nand U12886 (N_12886,N_11796,N_11334);
or U12887 (N_12887,N_10918,N_11512);
nor U12888 (N_12888,N_11330,N_9627);
or U12889 (N_12889,N_11438,N_9940);
nor U12890 (N_12890,N_9050,N_10431);
nand U12891 (N_12891,N_10865,N_9395);
xor U12892 (N_12892,N_11155,N_9148);
xnor U12893 (N_12893,N_9707,N_10787);
or U12894 (N_12894,N_11429,N_11586);
nor U12895 (N_12895,N_10230,N_11354);
nand U12896 (N_12896,N_11049,N_11839);
nand U12897 (N_12897,N_9758,N_10205);
or U12898 (N_12898,N_10246,N_10441);
nand U12899 (N_12899,N_11940,N_9047);
nor U12900 (N_12900,N_10298,N_10874);
or U12901 (N_12901,N_10105,N_11472);
xnor U12902 (N_12902,N_11312,N_11505);
nor U12903 (N_12903,N_9708,N_11578);
or U12904 (N_12904,N_10176,N_9684);
and U12905 (N_12905,N_11404,N_9928);
xor U12906 (N_12906,N_10941,N_11793);
nor U12907 (N_12907,N_10250,N_11376);
nand U12908 (N_12908,N_11767,N_11195);
or U12909 (N_12909,N_10600,N_11648);
nor U12910 (N_12910,N_9686,N_11942);
nor U12911 (N_12911,N_9231,N_9899);
and U12912 (N_12912,N_11320,N_11553);
nor U12913 (N_12913,N_11789,N_11498);
or U12914 (N_12914,N_11659,N_10016);
nand U12915 (N_12915,N_10739,N_10682);
and U12916 (N_12916,N_9936,N_10171);
and U12917 (N_12917,N_9729,N_9283);
xor U12918 (N_12918,N_9845,N_9802);
or U12919 (N_12919,N_9769,N_11693);
nor U12920 (N_12920,N_10490,N_10332);
and U12921 (N_12921,N_11070,N_10401);
or U12922 (N_12922,N_10173,N_11067);
or U12923 (N_12923,N_10288,N_10265);
or U12924 (N_12924,N_11528,N_11856);
or U12925 (N_12925,N_9065,N_10102);
or U12926 (N_12926,N_10361,N_11292);
and U12927 (N_12927,N_9205,N_9526);
and U12928 (N_12928,N_10353,N_9547);
nand U12929 (N_12929,N_11348,N_11995);
nand U12930 (N_12930,N_9131,N_10450);
nor U12931 (N_12931,N_10267,N_10751);
nand U12932 (N_12932,N_11622,N_10897);
and U12933 (N_12933,N_11908,N_9109);
nor U12934 (N_12934,N_10310,N_11201);
nand U12935 (N_12935,N_9920,N_11243);
nand U12936 (N_12936,N_9121,N_9168);
nand U12937 (N_12937,N_11937,N_10876);
or U12938 (N_12938,N_9189,N_11549);
and U12939 (N_12939,N_10291,N_9648);
and U12940 (N_12940,N_9752,N_11479);
xor U12941 (N_12941,N_9915,N_9891);
nand U12942 (N_12942,N_10617,N_10211);
nand U12943 (N_12943,N_10121,N_9218);
or U12944 (N_12944,N_9738,N_9204);
xor U12945 (N_12945,N_9186,N_11592);
or U12946 (N_12946,N_9600,N_9224);
nand U12947 (N_12947,N_11847,N_11057);
or U12948 (N_12948,N_9864,N_9509);
nand U12949 (N_12949,N_10653,N_11011);
and U12950 (N_12950,N_9806,N_11316);
nand U12951 (N_12951,N_11519,N_9371);
xor U12952 (N_12952,N_9041,N_11739);
and U12953 (N_12953,N_11894,N_9406);
nor U12954 (N_12954,N_9391,N_10274);
nand U12955 (N_12955,N_11433,N_10229);
nand U12956 (N_12956,N_9866,N_11774);
nand U12957 (N_12957,N_9984,N_10029);
and U12958 (N_12958,N_9357,N_10944);
and U12959 (N_12959,N_11674,N_11562);
nor U12960 (N_12960,N_10546,N_10766);
nand U12961 (N_12961,N_9316,N_11257);
and U12962 (N_12962,N_11140,N_9718);
nor U12963 (N_12963,N_10012,N_11058);
or U12964 (N_12964,N_10700,N_10615);
and U12965 (N_12965,N_9461,N_9269);
nor U12966 (N_12966,N_10712,N_10066);
or U12967 (N_12967,N_11878,N_10948);
or U12968 (N_12968,N_11458,N_9965);
or U12969 (N_12969,N_9392,N_10683);
nand U12970 (N_12970,N_10803,N_11266);
or U12971 (N_12971,N_9122,N_10499);
and U12972 (N_12972,N_10236,N_10503);
or U12973 (N_12973,N_11841,N_9992);
xnor U12974 (N_12974,N_9587,N_10140);
or U12975 (N_12975,N_11137,N_11401);
nor U12976 (N_12976,N_10695,N_11906);
and U12977 (N_12977,N_10734,N_10720);
nor U12978 (N_12978,N_9416,N_9118);
or U12979 (N_12979,N_9038,N_10436);
and U12980 (N_12980,N_10202,N_11861);
and U12981 (N_12981,N_9161,N_9621);
or U12982 (N_12982,N_10373,N_11759);
nor U12983 (N_12983,N_11301,N_10256);
and U12984 (N_12984,N_11790,N_11976);
and U12985 (N_12985,N_11342,N_11440);
or U12986 (N_12986,N_11880,N_11310);
nand U12987 (N_12987,N_11171,N_11916);
nor U12988 (N_12988,N_11615,N_9383);
or U12989 (N_12989,N_9789,N_10904);
and U12990 (N_12990,N_10113,N_9475);
and U12991 (N_12991,N_10338,N_9850);
xor U12992 (N_12992,N_10969,N_11735);
nand U12993 (N_12993,N_9972,N_11200);
or U12994 (N_12994,N_9771,N_11770);
xnor U12995 (N_12995,N_9880,N_9051);
and U12996 (N_12996,N_10258,N_10678);
and U12997 (N_12997,N_11518,N_10474);
nand U12998 (N_12998,N_9792,N_11524);
nand U12999 (N_12999,N_9623,N_10888);
nor U13000 (N_13000,N_10399,N_9750);
nor U13001 (N_13001,N_10912,N_9871);
and U13002 (N_13002,N_11978,N_9719);
xor U13003 (N_13003,N_11004,N_11791);
nor U13004 (N_13004,N_10494,N_10774);
and U13005 (N_13005,N_9807,N_10194);
and U13006 (N_13006,N_10868,N_11346);
or U13007 (N_13007,N_10693,N_10828);
nand U13008 (N_13008,N_11915,N_9614);
and U13009 (N_13009,N_10879,N_9200);
xnor U13010 (N_13010,N_11509,N_11871);
and U13011 (N_13011,N_10869,N_10973);
nor U13012 (N_13012,N_10902,N_10666);
and U13013 (N_13013,N_9744,N_9531);
nor U13014 (N_13014,N_10698,N_10724);
nand U13015 (N_13015,N_9236,N_9565);
nor U13016 (N_13016,N_9551,N_9781);
or U13017 (N_13017,N_9434,N_10088);
nand U13018 (N_13018,N_11855,N_11366);
or U13019 (N_13019,N_10110,N_11664);
nand U13020 (N_13020,N_9039,N_9373);
nor U13021 (N_13021,N_10898,N_9432);
xor U13022 (N_13022,N_9688,N_9589);
or U13023 (N_13023,N_11245,N_11846);
nor U13024 (N_13024,N_9095,N_11175);
or U13025 (N_13025,N_10341,N_10783);
nand U13026 (N_13026,N_9893,N_11126);
nand U13027 (N_13027,N_9460,N_10933);
or U13028 (N_13028,N_10640,N_11668);
or U13029 (N_13029,N_9953,N_11527);
and U13030 (N_13030,N_10953,N_10245);
or U13031 (N_13031,N_9436,N_11901);
nand U13032 (N_13032,N_11556,N_10048);
and U13033 (N_13033,N_11446,N_10841);
and U13034 (N_13034,N_9203,N_11711);
and U13035 (N_13035,N_11762,N_9778);
and U13036 (N_13036,N_11798,N_9398);
nand U13037 (N_13037,N_10671,N_10844);
or U13038 (N_13038,N_10395,N_10204);
nor U13039 (N_13039,N_11074,N_9990);
nand U13040 (N_13040,N_9917,N_9343);
nand U13041 (N_13041,N_9389,N_11853);
nor U13042 (N_13042,N_9338,N_9094);
or U13043 (N_13043,N_11653,N_10770);
and U13044 (N_13044,N_11882,N_11408);
or U13045 (N_13045,N_10120,N_11143);
or U13046 (N_13046,N_9519,N_11045);
xnor U13047 (N_13047,N_11428,N_10435);
nand U13048 (N_13048,N_10779,N_9273);
or U13049 (N_13049,N_9323,N_10508);
nor U13050 (N_13050,N_11854,N_11020);
xnor U13051 (N_13051,N_9982,N_11525);
nand U13052 (N_13052,N_10830,N_9665);
nor U13053 (N_13053,N_10691,N_10222);
nand U13054 (N_13054,N_9597,N_9798);
or U13055 (N_13055,N_9230,N_9638);
nor U13056 (N_13056,N_11097,N_11460);
nor U13057 (N_13057,N_10936,N_9949);
xor U13058 (N_13058,N_9457,N_9629);
nor U13059 (N_13059,N_10635,N_11230);
and U13060 (N_13060,N_10781,N_9008);
xnor U13061 (N_13061,N_9497,N_9076);
nor U13062 (N_13062,N_10564,N_11164);
or U13063 (N_13063,N_9268,N_11632);
nand U13064 (N_13064,N_9400,N_11359);
nand U13065 (N_13065,N_11116,N_11205);
xor U13066 (N_13066,N_10398,N_9745);
xnor U13067 (N_13067,N_10811,N_9925);
and U13068 (N_13068,N_9537,N_11669);
nand U13069 (N_13069,N_10424,N_10911);
and U13070 (N_13070,N_11420,N_11548);
or U13071 (N_13071,N_11261,N_11082);
and U13072 (N_13072,N_11148,N_9403);
and U13073 (N_13073,N_9527,N_9777);
or U13074 (N_13074,N_11127,N_9149);
or U13075 (N_13075,N_10735,N_10614);
and U13076 (N_13076,N_10362,N_10158);
nor U13077 (N_13077,N_11923,N_11378);
and U13078 (N_13078,N_10289,N_11008);
nor U13079 (N_13079,N_11144,N_10005);
nor U13080 (N_13080,N_11005,N_10946);
nand U13081 (N_13081,N_10956,N_10551);
or U13082 (N_13082,N_9412,N_11051);
nor U13083 (N_13083,N_11442,N_10059);
or U13084 (N_13084,N_9439,N_11047);
or U13085 (N_13085,N_11573,N_11981);
and U13086 (N_13086,N_9320,N_10901);
or U13087 (N_13087,N_10241,N_9344);
and U13088 (N_13088,N_11705,N_10747);
and U13089 (N_13089,N_9507,N_10959);
and U13090 (N_13090,N_9311,N_11699);
nor U13091 (N_13091,N_11621,N_10360);
nand U13092 (N_13092,N_11552,N_10767);
nand U13093 (N_13093,N_11802,N_11131);
nor U13094 (N_13094,N_10673,N_11834);
and U13095 (N_13095,N_9825,N_11879);
and U13096 (N_13096,N_10085,N_11412);
nand U13097 (N_13097,N_11013,N_10079);
or U13098 (N_13098,N_9605,N_10055);
nand U13099 (N_13099,N_10652,N_9857);
or U13100 (N_13100,N_9774,N_10286);
nor U13101 (N_13101,N_11779,N_9215);
nand U13102 (N_13102,N_10554,N_10582);
nand U13103 (N_13103,N_9554,N_11265);
or U13104 (N_13104,N_11071,N_9535);
nand U13105 (N_13105,N_11023,N_9213);
nor U13106 (N_13106,N_10900,N_9462);
or U13107 (N_13107,N_10106,N_10127);
nand U13108 (N_13108,N_11863,N_9569);
xor U13109 (N_13109,N_10945,N_10177);
or U13110 (N_13110,N_11572,N_10248);
and U13111 (N_13111,N_10128,N_10528);
or U13112 (N_13112,N_11782,N_11223);
nand U13113 (N_13113,N_10629,N_11559);
nor U13114 (N_13114,N_9979,N_9232);
or U13115 (N_13115,N_11996,N_10427);
or U13116 (N_13116,N_9484,N_9910);
or U13117 (N_13117,N_10578,N_10451);
nor U13118 (N_13118,N_11939,N_9302);
and U13119 (N_13119,N_10056,N_9524);
and U13120 (N_13120,N_10595,N_9784);
nor U13121 (N_13121,N_11914,N_10593);
and U13122 (N_13122,N_11297,N_11110);
or U13123 (N_13123,N_9819,N_11464);
and U13124 (N_13124,N_10181,N_9736);
nor U13125 (N_13125,N_9354,N_9082);
xnor U13126 (N_13126,N_11724,N_11636);
nor U13127 (N_13127,N_9700,N_9958);
nand U13128 (N_13128,N_10023,N_11579);
or U13129 (N_13129,N_11018,N_11331);
and U13130 (N_13130,N_11066,N_10182);
nand U13131 (N_13131,N_10290,N_11764);
nand U13132 (N_13132,N_10412,N_9471);
nand U13133 (N_13133,N_10253,N_9486);
nand U13134 (N_13134,N_9464,N_9381);
nor U13135 (N_13135,N_11056,N_11483);
and U13136 (N_13136,N_9023,N_11182);
nor U13137 (N_13137,N_9740,N_10296);
and U13138 (N_13138,N_9759,N_9278);
and U13139 (N_13139,N_10606,N_11138);
nor U13140 (N_13140,N_9404,N_9682);
or U13141 (N_13141,N_11600,N_9335);
nand U13142 (N_13142,N_10301,N_9019);
or U13143 (N_13143,N_10193,N_9851);
or U13144 (N_13144,N_11665,N_11803);
or U13145 (N_13145,N_10420,N_11530);
nand U13146 (N_13146,N_10951,N_11810);
nand U13147 (N_13147,N_11407,N_11694);
and U13148 (N_13148,N_10159,N_11663);
xnor U13149 (N_13149,N_11044,N_9591);
and U13150 (N_13150,N_10619,N_9074);
nand U13151 (N_13151,N_10465,N_10731);
or U13152 (N_13152,N_10087,N_11115);
nor U13153 (N_13153,N_9650,N_10254);
and U13154 (N_13154,N_10993,N_9810);
nor U13155 (N_13155,N_9376,N_10585);
and U13156 (N_13156,N_10000,N_10013);
nor U13157 (N_13157,N_11718,N_11073);
or U13158 (N_13158,N_11159,N_10216);
nor U13159 (N_13159,N_9066,N_11602);
and U13160 (N_13160,N_9125,N_10132);
nand U13161 (N_13161,N_9184,N_9225);
nor U13162 (N_13162,N_11042,N_10070);
nand U13163 (N_13163,N_9839,N_10068);
xnor U13164 (N_13164,N_11554,N_10630);
and U13165 (N_13165,N_9222,N_9593);
nor U13166 (N_13166,N_9282,N_9521);
xor U13167 (N_13167,N_11313,N_9644);
and U13168 (N_13168,N_9923,N_11054);
xnor U13169 (N_13169,N_9674,N_9969);
nor U13170 (N_13170,N_11471,N_10334);
nand U13171 (N_13171,N_9446,N_10355);
nor U13172 (N_13172,N_9105,N_10396);
or U13173 (N_13173,N_11384,N_11035);
nand U13174 (N_13174,N_9944,N_9529);
nor U13175 (N_13175,N_9327,N_10627);
and U13176 (N_13176,N_10566,N_11409);
and U13177 (N_13177,N_10798,N_9456);
xor U13178 (N_13178,N_9077,N_9123);
nand U13179 (N_13179,N_9030,N_10974);
and U13180 (N_13180,N_9454,N_9862);
and U13181 (N_13181,N_9727,N_11193);
and U13182 (N_13182,N_9207,N_9164);
nor U13183 (N_13183,N_11661,N_10832);
nand U13184 (N_13184,N_10930,N_11710);
or U13185 (N_13185,N_10772,N_10764);
and U13186 (N_13186,N_9219,N_11814);
nand U13187 (N_13187,N_11254,N_9512);
and U13188 (N_13188,N_10702,N_11507);
nor U13189 (N_13189,N_11194,N_9233);
and U13190 (N_13190,N_10243,N_9514);
nand U13191 (N_13191,N_10021,N_10179);
nand U13192 (N_13192,N_10607,N_10570);
and U13193 (N_13193,N_11502,N_10875);
nand U13194 (N_13194,N_11690,N_11160);
and U13195 (N_13195,N_11336,N_9156);
and U13196 (N_13196,N_9889,N_11926);
nor U13197 (N_13197,N_9730,N_9715);
nand U13198 (N_13198,N_9348,N_9251);
and U13199 (N_13199,N_10234,N_9670);
nand U13200 (N_13200,N_9104,N_10950);
nand U13201 (N_13201,N_11113,N_9221);
or U13202 (N_13202,N_9220,N_11153);
nor U13203 (N_13203,N_11345,N_10664);
nand U13204 (N_13204,N_10588,N_9652);
nor U13205 (N_13205,N_11238,N_9007);
or U13206 (N_13206,N_9868,N_10527);
and U13207 (N_13207,N_10317,N_11432);
nor U13208 (N_13208,N_10957,N_9190);
nand U13209 (N_13209,N_11215,N_10824);
or U13210 (N_13210,N_11593,N_11311);
or U13211 (N_13211,N_9329,N_11135);
or U13212 (N_13212,N_10468,N_10385);
and U13213 (N_13213,N_9801,N_10512);
xor U13214 (N_13214,N_9816,N_11361);
nand U13215 (N_13215,N_9423,N_9656);
nor U13216 (N_13216,N_9602,N_10303);
xnor U13217 (N_13217,N_11271,N_11958);
nand U13218 (N_13218,N_11247,N_10209);
nand U13219 (N_13219,N_10107,N_11418);
or U13220 (N_13220,N_9198,N_9995);
nor U13221 (N_13221,N_11558,N_10915);
nor U13222 (N_13222,N_10636,N_11403);
nor U13223 (N_13223,N_11387,N_11283);
or U13224 (N_13224,N_10639,N_11125);
nor U13225 (N_13225,N_9011,N_9280);
nand U13226 (N_13226,N_11218,N_10838);
and U13227 (N_13227,N_10348,N_10309);
nand U13228 (N_13228,N_9002,N_9132);
or U13229 (N_13229,N_10516,N_11543);
nor U13230 (N_13230,N_10555,N_9553);
and U13231 (N_13231,N_10738,N_9346);
and U13232 (N_13232,N_9751,N_10597);
and U13233 (N_13233,N_9848,N_9856);
nand U13234 (N_13234,N_9698,N_11588);
nand U13235 (N_13235,N_9277,N_11797);
or U13236 (N_13236,N_10703,N_9351);
nand U13237 (N_13237,N_10624,N_10454);
xor U13238 (N_13238,N_11100,N_10057);
nand U13239 (N_13239,N_11398,N_10851);
nor U13240 (N_13240,N_10577,N_9968);
nor U13241 (N_13241,N_11596,N_10988);
xnor U13242 (N_13242,N_11151,N_9017);
xnor U13243 (N_13243,N_11486,N_11783);
and U13244 (N_13244,N_9640,N_10157);
or U13245 (N_13245,N_11068,N_11654);
nand U13246 (N_13246,N_9838,N_9755);
nor U13247 (N_13247,N_11752,N_10562);
or U13248 (N_13248,N_9907,N_9339);
nor U13249 (N_13249,N_10495,N_11836);
and U13250 (N_13250,N_11713,N_10071);
and U13251 (N_13251,N_9783,N_9904);
xor U13252 (N_13252,N_11581,N_11633);
or U13253 (N_13253,N_9952,N_10949);
xor U13254 (N_13254,N_10845,N_10086);
nor U13255 (N_13255,N_11397,N_11443);
nor U13256 (N_13256,N_9349,N_11972);
or U13257 (N_13257,N_10638,N_10641);
and U13258 (N_13258,N_10356,N_9176);
and U13259 (N_13259,N_10324,N_11720);
nand U13260 (N_13260,N_9655,N_11484);
and U13261 (N_13261,N_11303,N_11174);
nand U13262 (N_13262,N_10696,N_9060);
nand U13263 (N_13263,N_10460,N_9588);
xnor U13264 (N_13264,N_11470,N_10081);
nand U13265 (N_13265,N_10487,N_9976);
xor U13266 (N_13266,N_10672,N_11349);
nor U13267 (N_13267,N_10049,N_10139);
nor U13268 (N_13268,N_11504,N_11513);
and U13269 (N_13269,N_9115,N_10283);
nor U13270 (N_13270,N_11758,N_9291);
xnor U13271 (N_13271,N_10414,N_10019);
and U13272 (N_13272,N_9243,N_10644);
xnor U13273 (N_13273,N_10923,N_10430);
or U13274 (N_13274,N_11133,N_11642);
nor U13275 (N_13275,N_11709,N_11129);
and U13276 (N_13276,N_9016,N_9056);
nor U13277 (N_13277,N_10663,N_10082);
or U13278 (N_13278,N_10228,N_9114);
or U13279 (N_13279,N_11911,N_10580);
or U13280 (N_13280,N_9474,N_11399);
and U13281 (N_13281,N_11865,N_9068);
or U13282 (N_13282,N_9018,N_9772);
or U13283 (N_13283,N_10511,N_11288);
and U13284 (N_13284,N_10442,N_11322);
and U13285 (N_13285,N_9488,N_9012);
and U13286 (N_13286,N_11985,N_10701);
nor U13287 (N_13287,N_10910,N_10453);
nor U13288 (N_13288,N_10126,N_10880);
and U13289 (N_13289,N_10519,N_11721);
nand U13290 (N_13290,N_10391,N_11953);
nor U13291 (N_13291,N_9272,N_10153);
xnor U13292 (N_13292,N_9239,N_9580);
nor U13293 (N_13293,N_11069,N_10099);
or U13294 (N_13294,N_10238,N_11491);
nor U13295 (N_13295,N_10142,N_10067);
nand U13296 (N_13296,N_9559,N_11684);
and U13297 (N_13297,N_11949,N_9154);
nor U13298 (N_13298,N_10996,N_10905);
and U13299 (N_13299,N_9828,N_9827);
xor U13300 (N_13300,N_11101,N_11938);
xor U13301 (N_13301,N_9628,N_11326);
nand U13302 (N_13302,N_10975,N_10439);
and U13303 (N_13303,N_10997,N_11241);
nand U13304 (N_13304,N_11598,N_11219);
nor U13305 (N_13305,N_11936,N_11844);
xnor U13306 (N_13306,N_10285,N_9418);
nor U13307 (N_13307,N_10273,N_10676);
or U13308 (N_13308,N_11274,N_10992);
and U13309 (N_13309,N_9054,N_10521);
and U13310 (N_13310,N_10612,N_9072);
or U13311 (N_13311,N_11918,N_10645);
and U13312 (N_13312,N_9465,N_11060);
or U13313 (N_13313,N_9199,N_10628);
and U13314 (N_13314,N_10390,N_9756);
or U13315 (N_13315,N_11951,N_11150);
nor U13316 (N_13316,N_11385,N_11367);
nor U13317 (N_13317,N_9044,N_10983);
or U13318 (N_13318,N_10668,N_10717);
nand U13319 (N_13319,N_10047,N_9101);
nand U13320 (N_13320,N_9493,N_9326);
nand U13321 (N_13321,N_10292,N_11891);
nor U13322 (N_13322,N_11666,N_9879);
and U13323 (N_13323,N_11740,N_9279);
xor U13324 (N_13324,N_10777,N_10352);
or U13325 (N_13325,N_9043,N_10873);
nand U13326 (N_13326,N_11859,N_9141);
and U13327 (N_13327,N_9419,N_11804);
xnor U13328 (N_13328,N_11426,N_9955);
nand U13329 (N_13329,N_9197,N_10270);
or U13330 (N_13330,N_9843,N_10122);
xor U13331 (N_13331,N_11725,N_11835);
or U13332 (N_13332,N_10313,N_10538);
and U13333 (N_13333,N_9813,N_9099);
nor U13334 (N_13334,N_9994,N_11701);
nor U13335 (N_13335,N_9353,N_10810);
or U13336 (N_13336,N_11481,N_9201);
and U13337 (N_13337,N_9921,N_10206);
or U13338 (N_13338,N_11992,N_9595);
nand U13339 (N_13339,N_10656,N_11172);
or U13340 (N_13340,N_9661,N_11987);
xnor U13341 (N_13341,N_9929,N_11508);
xor U13342 (N_13342,N_9405,N_10745);
nand U13343 (N_13343,N_11892,N_11945);
or U13344 (N_13344,N_10004,N_10131);
nor U13345 (N_13345,N_11933,N_11820);
or U13346 (N_13346,N_11867,N_9372);
and U13347 (N_13347,N_10931,N_10343);
or U13348 (N_13348,N_11081,N_9622);
nor U13349 (N_13349,N_11029,N_11282);
and U13350 (N_13350,N_10017,N_9747);
nand U13351 (N_13351,N_9001,N_11080);
nor U13352 (N_13352,N_10223,N_10397);
and U13353 (N_13353,N_11971,N_10655);
and U13354 (N_13354,N_11279,N_10063);
and U13355 (N_13355,N_10455,N_10116);
or U13356 (N_13356,N_10060,N_11111);
nor U13357 (N_13357,N_11032,N_9817);
nor U13358 (N_13358,N_10591,N_9922);
or U13359 (N_13359,N_9170,N_11662);
nor U13360 (N_13360,N_11613,N_9942);
nor U13361 (N_13361,N_11577,N_10903);
nand U13362 (N_13362,N_10111,N_10168);
or U13363 (N_13363,N_10537,N_11775);
xor U13364 (N_13364,N_9690,N_9037);
nand U13365 (N_13365,N_9768,N_9534);
nor U13366 (N_13366,N_10955,N_11968);
and U13367 (N_13367,N_11610,N_9188);
xor U13368 (N_13368,N_9571,N_10753);
and U13369 (N_13369,N_9869,N_10896);
or U13370 (N_13370,N_11801,N_10533);
and U13371 (N_13371,N_10800,N_9748);
and U13372 (N_13372,N_10815,N_11242);
nor U13373 (N_13373,N_10526,N_10266);
nor U13374 (N_13374,N_9517,N_11875);
nand U13375 (N_13375,N_11866,N_9135);
nor U13376 (N_13376,N_11207,N_10163);
nor U13377 (N_13377,N_10856,N_9062);
and U13378 (N_13378,N_9626,N_11183);
or U13379 (N_13379,N_11685,N_10589);
or U13380 (N_13380,N_10477,N_10940);
and U13381 (N_13381,N_11093,N_9765);
nand U13382 (N_13382,N_10601,N_10440);
or U13383 (N_13383,N_10947,N_9678);
nor U13384 (N_13384,N_11561,N_10603);
nor U13385 (N_13385,N_11079,N_9140);
xnor U13386 (N_13386,N_10547,N_10866);
and U13387 (N_13387,N_9133,N_9476);
nand U13388 (N_13388,N_10622,N_11734);
nor U13389 (N_13389,N_9539,N_9842);
nor U13390 (N_13390,N_10053,N_11166);
nor U13391 (N_13391,N_10178,N_9937);
nor U13392 (N_13392,N_9691,N_11321);
and U13393 (N_13393,N_10129,N_10609);
nand U13394 (N_13394,N_10221,N_11787);
or U13395 (N_13395,N_11819,N_10637);
or U13396 (N_13396,N_11919,N_10748);
and U13397 (N_13397,N_10743,N_11377);
and U13398 (N_13398,N_10003,N_9265);
or U13399 (N_13399,N_10001,N_11631);
and U13400 (N_13400,N_11002,N_9717);
or U13401 (N_13401,N_9119,N_10145);
and U13402 (N_13402,N_9782,N_11544);
nor U13403 (N_13403,N_11881,N_9015);
nor U13404 (N_13404,N_11208,N_11599);
or U13405 (N_13405,N_9275,N_9884);
nand U13406 (N_13406,N_9841,N_10184);
xor U13407 (N_13407,N_9014,N_9954);
nand U13408 (N_13408,N_11217,N_11928);
or U13409 (N_13409,N_9875,N_10616);
nor U13410 (N_13410,N_10018,N_11037);
nand U13411 (N_13411,N_11272,N_10146);
and U13412 (N_13412,N_11520,N_11447);
and U13413 (N_13413,N_11315,N_11078);
and U13414 (N_13414,N_11973,N_9413);
or U13415 (N_13415,N_9892,N_9753);
or U13416 (N_13416,N_11474,N_10827);
xor U13417 (N_13417,N_9322,N_11184);
nand U13418 (N_13418,N_9181,N_9505);
nand U13419 (N_13419,N_11993,N_9172);
nor U13420 (N_13420,N_9791,N_10713);
or U13421 (N_13421,N_9988,N_9878);
and U13422 (N_13422,N_10569,N_10536);
and U13423 (N_13423,N_9867,N_9049);
xor U13424 (N_13424,N_10610,N_9087);
or U13425 (N_13425,N_10669,N_10039);
nand U13426 (N_13426,N_11950,N_10072);
or U13427 (N_13427,N_11851,N_9155);
and U13428 (N_13428,N_10797,N_10219);
or U13429 (N_13429,N_10076,N_10119);
or U13430 (N_13430,N_11391,N_9558);
nor U13431 (N_13431,N_10584,N_11152);
or U13432 (N_13432,N_9113,N_11594);
and U13433 (N_13433,N_9567,N_10130);
and U13434 (N_13434,N_10095,N_10563);
nor U13435 (N_13435,N_9544,N_9550);
or U13436 (N_13436,N_9890,N_10197);
or U13437 (N_13437,N_9532,N_10826);
or U13438 (N_13438,N_11954,N_11877);
nand U13439 (N_13439,N_10510,N_9352);
nand U13440 (N_13440,N_9697,N_11007);
or U13441 (N_13441,N_9855,N_10410);
nor U13442 (N_13442,N_9112,N_10481);
or U13443 (N_13443,N_9293,N_9359);
nor U13444 (N_13444,N_9111,N_9865);
and U13445 (N_13445,N_9574,N_11760);
or U13446 (N_13446,N_9483,N_9673);
or U13447 (N_13447,N_10377,N_10482);
and U13448 (N_13448,N_9237,N_11702);
xnor U13449 (N_13449,N_10692,N_9667);
nor U13450 (N_13450,N_10407,N_10819);
or U13451 (N_13451,N_9455,N_11256);
nand U13452 (N_13452,N_9440,N_10415);
or U13453 (N_13453,N_9832,N_11962);
nand U13454 (N_13454,N_11264,N_9430);
nand U13455 (N_13455,N_11373,N_9482);
and U13456 (N_13456,N_9704,N_9426);
or U13457 (N_13457,N_10846,N_9945);
and U13458 (N_13458,N_10154,N_9566);
or U13459 (N_13459,N_9096,N_11570);
or U13460 (N_13460,N_9127,N_10405);
or U13461 (N_13461,N_11754,N_9773);
nor U13462 (N_13462,N_11273,N_11827);
nor U13463 (N_13463,N_11983,N_9989);
nand U13464 (N_13464,N_11729,N_11375);
and U13465 (N_13465,N_9499,N_9300);
nor U13466 (N_13466,N_9693,N_9766);
nand U13467 (N_13467,N_11318,N_9425);
and U13468 (N_13468,N_11059,N_10867);
nor U13469 (N_13469,N_9325,N_9840);
nor U13470 (N_13470,N_9388,N_10240);
nor U13471 (N_13471,N_10161,N_9948);
or U13472 (N_13472,N_9849,N_10932);
and U13473 (N_13473,N_9301,N_11454);
nor U13474 (N_13474,N_11781,N_9901);
nor U13475 (N_13475,N_11436,N_11466);
and U13476 (N_13476,N_10834,N_10025);
nand U13477 (N_13477,N_11898,N_10042);
and U13478 (N_13478,N_10706,N_10043);
nor U13479 (N_13479,N_10123,N_11392);
nor U13480 (N_13480,N_11565,N_10756);
and U13481 (N_13481,N_10423,N_10022);
or U13482 (N_13482,N_11627,N_9538);
nor U13483 (N_13483,N_10805,N_11857);
nor U13484 (N_13484,N_10882,N_10475);
nor U13485 (N_13485,N_9063,N_9998);
nor U13486 (N_13486,N_11902,N_11102);
nor U13487 (N_13487,N_9964,N_9262);
nor U13488 (N_13488,N_10843,N_9345);
nor U13489 (N_13489,N_9578,N_9128);
nand U13490 (N_13490,N_11723,N_9009);
and U13491 (N_13491,N_10327,N_10964);
and U13492 (N_13492,N_11165,N_10030);
or U13493 (N_13493,N_11146,N_11128);
nand U13494 (N_13494,N_9808,N_9245);
and U13495 (N_13495,N_9902,N_10509);
and U13496 (N_13496,N_9743,N_10925);
and U13497 (N_13497,N_11934,N_11609);
or U13498 (N_13498,N_10850,N_10884);
nand U13499 (N_13499,N_10773,N_11806);
nand U13500 (N_13500,N_10595,N_9970);
nand U13501 (N_13501,N_11144,N_10420);
or U13502 (N_13502,N_11253,N_11338);
or U13503 (N_13503,N_11352,N_11310);
or U13504 (N_13504,N_9942,N_11302);
nand U13505 (N_13505,N_9113,N_10101);
xnor U13506 (N_13506,N_10047,N_10474);
and U13507 (N_13507,N_10126,N_11117);
xnor U13508 (N_13508,N_11324,N_10460);
or U13509 (N_13509,N_10684,N_9407);
nand U13510 (N_13510,N_9872,N_9833);
and U13511 (N_13511,N_11865,N_9371);
nand U13512 (N_13512,N_11668,N_11369);
nand U13513 (N_13513,N_11385,N_11338);
and U13514 (N_13514,N_10758,N_9042);
or U13515 (N_13515,N_10066,N_10533);
or U13516 (N_13516,N_11095,N_10626);
or U13517 (N_13517,N_9728,N_10732);
or U13518 (N_13518,N_11715,N_11307);
and U13519 (N_13519,N_9397,N_9586);
nor U13520 (N_13520,N_10496,N_11083);
nand U13521 (N_13521,N_11615,N_9504);
nand U13522 (N_13522,N_10444,N_11512);
nand U13523 (N_13523,N_11126,N_9142);
or U13524 (N_13524,N_9666,N_9451);
and U13525 (N_13525,N_10935,N_9673);
and U13526 (N_13526,N_10055,N_9912);
nand U13527 (N_13527,N_9760,N_11989);
and U13528 (N_13528,N_11619,N_10326);
nand U13529 (N_13529,N_11929,N_10961);
nor U13530 (N_13530,N_10554,N_10962);
xor U13531 (N_13531,N_11284,N_11296);
nor U13532 (N_13532,N_9385,N_10994);
nor U13533 (N_13533,N_11112,N_11201);
and U13534 (N_13534,N_11529,N_10787);
or U13535 (N_13535,N_11435,N_11931);
nand U13536 (N_13536,N_10914,N_9910);
or U13537 (N_13537,N_9624,N_9446);
or U13538 (N_13538,N_10463,N_10630);
nor U13539 (N_13539,N_9166,N_10642);
nand U13540 (N_13540,N_10612,N_9546);
or U13541 (N_13541,N_11570,N_9242);
or U13542 (N_13542,N_9261,N_11345);
xor U13543 (N_13543,N_10983,N_9620);
and U13544 (N_13544,N_11515,N_10880);
nand U13545 (N_13545,N_10530,N_9660);
nor U13546 (N_13546,N_9673,N_9080);
nor U13547 (N_13547,N_9096,N_9743);
nor U13548 (N_13548,N_10486,N_10756);
and U13549 (N_13549,N_10738,N_9118);
nand U13550 (N_13550,N_11367,N_10080);
and U13551 (N_13551,N_10060,N_11918);
or U13552 (N_13552,N_11263,N_10696);
or U13553 (N_13553,N_11016,N_11980);
nand U13554 (N_13554,N_11487,N_9754);
and U13555 (N_13555,N_10485,N_9469);
and U13556 (N_13556,N_11610,N_11567);
nand U13557 (N_13557,N_9577,N_9674);
nor U13558 (N_13558,N_10141,N_11296);
and U13559 (N_13559,N_11851,N_9328);
nand U13560 (N_13560,N_11888,N_11045);
and U13561 (N_13561,N_10152,N_10301);
and U13562 (N_13562,N_11034,N_9874);
and U13563 (N_13563,N_10079,N_11679);
nor U13564 (N_13564,N_10403,N_10197);
and U13565 (N_13565,N_11875,N_10359);
or U13566 (N_13566,N_10242,N_11129);
or U13567 (N_13567,N_10984,N_10310);
and U13568 (N_13568,N_11143,N_9817);
nor U13569 (N_13569,N_9823,N_11534);
nor U13570 (N_13570,N_9924,N_10630);
xnor U13571 (N_13571,N_10886,N_10599);
nor U13572 (N_13572,N_10469,N_9345);
and U13573 (N_13573,N_9999,N_9431);
xor U13574 (N_13574,N_9200,N_10859);
nor U13575 (N_13575,N_9323,N_11679);
or U13576 (N_13576,N_10408,N_11681);
xnor U13577 (N_13577,N_9081,N_11868);
and U13578 (N_13578,N_10528,N_9698);
or U13579 (N_13579,N_10560,N_10185);
nor U13580 (N_13580,N_11251,N_11408);
nand U13581 (N_13581,N_9320,N_9001);
and U13582 (N_13582,N_10788,N_9368);
nor U13583 (N_13583,N_9771,N_11948);
and U13584 (N_13584,N_9943,N_9676);
and U13585 (N_13585,N_11314,N_11605);
nor U13586 (N_13586,N_10882,N_10074);
nor U13587 (N_13587,N_10336,N_9894);
nor U13588 (N_13588,N_11080,N_9022);
nor U13589 (N_13589,N_10539,N_11892);
or U13590 (N_13590,N_10365,N_9610);
nand U13591 (N_13591,N_9377,N_10546);
and U13592 (N_13592,N_11996,N_9867);
or U13593 (N_13593,N_9797,N_10033);
or U13594 (N_13594,N_9790,N_11846);
nand U13595 (N_13595,N_11298,N_11984);
or U13596 (N_13596,N_10446,N_9970);
nand U13597 (N_13597,N_10160,N_9335);
nand U13598 (N_13598,N_11760,N_9254);
nand U13599 (N_13599,N_9459,N_11587);
nor U13600 (N_13600,N_9463,N_10349);
nand U13601 (N_13601,N_10005,N_10090);
nand U13602 (N_13602,N_11712,N_9289);
nand U13603 (N_13603,N_11577,N_10501);
xnor U13604 (N_13604,N_9567,N_9231);
nor U13605 (N_13605,N_11172,N_11176);
or U13606 (N_13606,N_9355,N_10025);
nand U13607 (N_13607,N_10031,N_11595);
nor U13608 (N_13608,N_10942,N_10106);
xor U13609 (N_13609,N_9665,N_10544);
or U13610 (N_13610,N_11375,N_10995);
nand U13611 (N_13611,N_10004,N_11644);
nand U13612 (N_13612,N_9086,N_9282);
nand U13613 (N_13613,N_10402,N_9269);
or U13614 (N_13614,N_11040,N_11865);
or U13615 (N_13615,N_9242,N_11295);
nor U13616 (N_13616,N_10887,N_10953);
or U13617 (N_13617,N_10504,N_9845);
and U13618 (N_13618,N_9537,N_9150);
nor U13619 (N_13619,N_9013,N_10129);
or U13620 (N_13620,N_11109,N_9784);
or U13621 (N_13621,N_10396,N_9736);
nand U13622 (N_13622,N_10098,N_10430);
or U13623 (N_13623,N_9982,N_10595);
nor U13624 (N_13624,N_11301,N_11308);
and U13625 (N_13625,N_10250,N_11853);
and U13626 (N_13626,N_9930,N_9333);
nor U13627 (N_13627,N_9005,N_10777);
and U13628 (N_13628,N_11561,N_11116);
nand U13629 (N_13629,N_11167,N_9701);
xor U13630 (N_13630,N_11386,N_10833);
nor U13631 (N_13631,N_10363,N_11667);
xnor U13632 (N_13632,N_11464,N_11502);
and U13633 (N_13633,N_9519,N_11308);
nand U13634 (N_13634,N_9793,N_9839);
nor U13635 (N_13635,N_9707,N_10609);
nand U13636 (N_13636,N_11767,N_10850);
nor U13637 (N_13637,N_10481,N_11926);
or U13638 (N_13638,N_11222,N_11682);
and U13639 (N_13639,N_10891,N_10943);
nand U13640 (N_13640,N_11872,N_11109);
or U13641 (N_13641,N_9585,N_10893);
nor U13642 (N_13642,N_11131,N_9174);
and U13643 (N_13643,N_10266,N_10831);
or U13644 (N_13644,N_10938,N_9119);
and U13645 (N_13645,N_11412,N_11034);
xnor U13646 (N_13646,N_10540,N_9729);
nand U13647 (N_13647,N_9784,N_11912);
xnor U13648 (N_13648,N_10990,N_10690);
or U13649 (N_13649,N_10521,N_10201);
xor U13650 (N_13650,N_9180,N_9675);
and U13651 (N_13651,N_10671,N_9444);
and U13652 (N_13652,N_11587,N_11320);
and U13653 (N_13653,N_10337,N_10658);
and U13654 (N_13654,N_10889,N_10719);
nor U13655 (N_13655,N_9561,N_11894);
or U13656 (N_13656,N_10876,N_10299);
or U13657 (N_13657,N_10888,N_9421);
nand U13658 (N_13658,N_9543,N_11422);
or U13659 (N_13659,N_11161,N_10051);
nor U13660 (N_13660,N_10077,N_9444);
nor U13661 (N_13661,N_10254,N_9830);
and U13662 (N_13662,N_11524,N_10411);
nand U13663 (N_13663,N_11827,N_9891);
nand U13664 (N_13664,N_9216,N_11009);
nor U13665 (N_13665,N_10457,N_10850);
nor U13666 (N_13666,N_10064,N_9642);
or U13667 (N_13667,N_9725,N_10467);
and U13668 (N_13668,N_11169,N_11522);
nor U13669 (N_13669,N_9556,N_11951);
nor U13670 (N_13670,N_9578,N_10702);
or U13671 (N_13671,N_9542,N_11360);
nand U13672 (N_13672,N_11670,N_11198);
nor U13673 (N_13673,N_9578,N_11537);
and U13674 (N_13674,N_10731,N_9133);
nor U13675 (N_13675,N_11131,N_9267);
and U13676 (N_13676,N_9928,N_11202);
nand U13677 (N_13677,N_10623,N_11170);
and U13678 (N_13678,N_10369,N_10752);
nand U13679 (N_13679,N_11327,N_9774);
nand U13680 (N_13680,N_11965,N_9396);
nor U13681 (N_13681,N_10118,N_11832);
nor U13682 (N_13682,N_9866,N_9544);
nor U13683 (N_13683,N_10456,N_11024);
nor U13684 (N_13684,N_11863,N_9699);
nand U13685 (N_13685,N_10555,N_10523);
or U13686 (N_13686,N_9537,N_11117);
or U13687 (N_13687,N_10267,N_11533);
nand U13688 (N_13688,N_9862,N_10520);
xnor U13689 (N_13689,N_10238,N_10170);
and U13690 (N_13690,N_10971,N_11259);
or U13691 (N_13691,N_11712,N_10799);
or U13692 (N_13692,N_10342,N_11306);
nand U13693 (N_13693,N_10982,N_9516);
and U13694 (N_13694,N_9250,N_11719);
or U13695 (N_13695,N_10130,N_11381);
nor U13696 (N_13696,N_11699,N_10823);
and U13697 (N_13697,N_11877,N_11727);
nand U13698 (N_13698,N_9778,N_9723);
nor U13699 (N_13699,N_10844,N_9457);
nand U13700 (N_13700,N_11818,N_10090);
nand U13701 (N_13701,N_10824,N_9452);
xnor U13702 (N_13702,N_10910,N_9148);
or U13703 (N_13703,N_9454,N_11592);
or U13704 (N_13704,N_10250,N_10500);
and U13705 (N_13705,N_9095,N_9221);
nand U13706 (N_13706,N_10217,N_11428);
and U13707 (N_13707,N_10993,N_9384);
and U13708 (N_13708,N_10791,N_11928);
nand U13709 (N_13709,N_9694,N_10390);
and U13710 (N_13710,N_10250,N_11387);
nand U13711 (N_13711,N_10442,N_10050);
nand U13712 (N_13712,N_9580,N_11902);
or U13713 (N_13713,N_11952,N_9997);
nand U13714 (N_13714,N_11119,N_10022);
and U13715 (N_13715,N_11078,N_10025);
nand U13716 (N_13716,N_9387,N_11905);
nand U13717 (N_13717,N_10654,N_10818);
or U13718 (N_13718,N_9186,N_10343);
and U13719 (N_13719,N_10250,N_10568);
nand U13720 (N_13720,N_9367,N_10242);
xor U13721 (N_13721,N_10077,N_11447);
xnor U13722 (N_13722,N_11424,N_9448);
nand U13723 (N_13723,N_11963,N_9804);
or U13724 (N_13724,N_11127,N_9769);
and U13725 (N_13725,N_9094,N_10112);
nor U13726 (N_13726,N_10289,N_9787);
or U13727 (N_13727,N_10146,N_11818);
or U13728 (N_13728,N_9483,N_11998);
and U13729 (N_13729,N_9852,N_11725);
nor U13730 (N_13730,N_9430,N_9088);
or U13731 (N_13731,N_11658,N_10053);
xor U13732 (N_13732,N_9359,N_9086);
nand U13733 (N_13733,N_10143,N_9653);
nor U13734 (N_13734,N_9857,N_10182);
nand U13735 (N_13735,N_11477,N_11411);
and U13736 (N_13736,N_11400,N_9190);
or U13737 (N_13737,N_11176,N_10080);
nand U13738 (N_13738,N_11853,N_11229);
or U13739 (N_13739,N_9796,N_11344);
nand U13740 (N_13740,N_9483,N_11454);
xor U13741 (N_13741,N_9450,N_11155);
or U13742 (N_13742,N_10147,N_9778);
nor U13743 (N_13743,N_10906,N_10453);
and U13744 (N_13744,N_10521,N_9279);
xor U13745 (N_13745,N_10363,N_10594);
nand U13746 (N_13746,N_10996,N_11698);
and U13747 (N_13747,N_10929,N_11236);
and U13748 (N_13748,N_10281,N_10734);
or U13749 (N_13749,N_9282,N_9401);
nand U13750 (N_13750,N_11021,N_9282);
nor U13751 (N_13751,N_9896,N_9971);
nor U13752 (N_13752,N_9673,N_10559);
or U13753 (N_13753,N_11564,N_11284);
nand U13754 (N_13754,N_11367,N_9741);
xnor U13755 (N_13755,N_10609,N_11017);
or U13756 (N_13756,N_10919,N_11360);
nand U13757 (N_13757,N_10951,N_10807);
and U13758 (N_13758,N_10624,N_10488);
or U13759 (N_13759,N_11845,N_11533);
or U13760 (N_13760,N_10674,N_9580);
or U13761 (N_13761,N_9422,N_11558);
or U13762 (N_13762,N_10342,N_10798);
or U13763 (N_13763,N_9154,N_9725);
nand U13764 (N_13764,N_10797,N_10102);
and U13765 (N_13765,N_10084,N_10780);
nor U13766 (N_13766,N_10768,N_10671);
nand U13767 (N_13767,N_10636,N_11892);
xnor U13768 (N_13768,N_9285,N_10590);
nand U13769 (N_13769,N_11002,N_9632);
nand U13770 (N_13770,N_11127,N_10218);
or U13771 (N_13771,N_9681,N_10167);
and U13772 (N_13772,N_10257,N_11695);
nand U13773 (N_13773,N_9259,N_9968);
nand U13774 (N_13774,N_10690,N_11886);
nor U13775 (N_13775,N_11756,N_11561);
nor U13776 (N_13776,N_11507,N_10173);
nor U13777 (N_13777,N_9068,N_9555);
nand U13778 (N_13778,N_10858,N_11408);
nor U13779 (N_13779,N_9351,N_10437);
and U13780 (N_13780,N_11408,N_9031);
nor U13781 (N_13781,N_9334,N_9738);
and U13782 (N_13782,N_11771,N_10115);
nor U13783 (N_13783,N_10056,N_10917);
nand U13784 (N_13784,N_9203,N_10198);
and U13785 (N_13785,N_11236,N_11922);
and U13786 (N_13786,N_9824,N_10522);
and U13787 (N_13787,N_11172,N_9561);
and U13788 (N_13788,N_10429,N_9653);
and U13789 (N_13789,N_9614,N_9059);
nor U13790 (N_13790,N_11524,N_9424);
or U13791 (N_13791,N_9795,N_10544);
or U13792 (N_13792,N_10131,N_11853);
nand U13793 (N_13793,N_10806,N_10953);
or U13794 (N_13794,N_11591,N_10683);
nand U13795 (N_13795,N_9649,N_11253);
or U13796 (N_13796,N_10952,N_10685);
and U13797 (N_13797,N_11316,N_11251);
or U13798 (N_13798,N_11517,N_11748);
nor U13799 (N_13799,N_11290,N_10448);
or U13800 (N_13800,N_11077,N_11571);
and U13801 (N_13801,N_11596,N_10229);
or U13802 (N_13802,N_11909,N_9139);
nor U13803 (N_13803,N_9497,N_10285);
and U13804 (N_13804,N_9561,N_9978);
or U13805 (N_13805,N_9448,N_9835);
xnor U13806 (N_13806,N_9478,N_10500);
nor U13807 (N_13807,N_9371,N_9380);
and U13808 (N_13808,N_10403,N_11275);
xor U13809 (N_13809,N_10491,N_10350);
nor U13810 (N_13810,N_9050,N_11025);
nand U13811 (N_13811,N_9292,N_10346);
nand U13812 (N_13812,N_9390,N_9509);
and U13813 (N_13813,N_10546,N_10182);
nand U13814 (N_13814,N_11306,N_11428);
nand U13815 (N_13815,N_11564,N_9903);
and U13816 (N_13816,N_9446,N_10432);
and U13817 (N_13817,N_11806,N_9358);
and U13818 (N_13818,N_9422,N_10862);
nand U13819 (N_13819,N_9858,N_11193);
nor U13820 (N_13820,N_10852,N_10342);
nor U13821 (N_13821,N_9574,N_10255);
and U13822 (N_13822,N_11279,N_9257);
or U13823 (N_13823,N_9079,N_11811);
and U13824 (N_13824,N_11740,N_11625);
or U13825 (N_13825,N_11855,N_9737);
nor U13826 (N_13826,N_9258,N_11824);
or U13827 (N_13827,N_10258,N_11803);
or U13828 (N_13828,N_9992,N_11779);
and U13829 (N_13829,N_11520,N_11656);
or U13830 (N_13830,N_9424,N_10577);
and U13831 (N_13831,N_9689,N_9283);
and U13832 (N_13832,N_10821,N_10125);
or U13833 (N_13833,N_10068,N_9336);
and U13834 (N_13834,N_11267,N_10220);
xor U13835 (N_13835,N_10129,N_10196);
and U13836 (N_13836,N_10682,N_11912);
nand U13837 (N_13837,N_10578,N_10585);
and U13838 (N_13838,N_9366,N_10076);
nor U13839 (N_13839,N_11093,N_9188);
nor U13840 (N_13840,N_10626,N_9938);
and U13841 (N_13841,N_11963,N_11548);
or U13842 (N_13842,N_9163,N_10095);
or U13843 (N_13843,N_10340,N_11917);
or U13844 (N_13844,N_9125,N_10426);
nor U13845 (N_13845,N_10964,N_9195);
or U13846 (N_13846,N_10373,N_11766);
or U13847 (N_13847,N_9744,N_9826);
nand U13848 (N_13848,N_11474,N_10510);
nand U13849 (N_13849,N_9352,N_9235);
nor U13850 (N_13850,N_11969,N_10015);
xor U13851 (N_13851,N_10294,N_10366);
nor U13852 (N_13852,N_11772,N_10805);
nand U13853 (N_13853,N_11642,N_11606);
or U13854 (N_13854,N_10181,N_10488);
xnor U13855 (N_13855,N_10070,N_11264);
and U13856 (N_13856,N_9415,N_10995);
and U13857 (N_13857,N_11884,N_9485);
nor U13858 (N_13858,N_9379,N_9305);
nor U13859 (N_13859,N_11788,N_10441);
nand U13860 (N_13860,N_10990,N_9229);
or U13861 (N_13861,N_11496,N_9043);
and U13862 (N_13862,N_9914,N_9991);
xnor U13863 (N_13863,N_10268,N_9884);
or U13864 (N_13864,N_9484,N_10460);
and U13865 (N_13865,N_11885,N_9115);
or U13866 (N_13866,N_10591,N_10123);
or U13867 (N_13867,N_9657,N_10322);
nor U13868 (N_13868,N_9421,N_10278);
nor U13869 (N_13869,N_10955,N_11562);
xnor U13870 (N_13870,N_9030,N_9919);
nor U13871 (N_13871,N_9495,N_11396);
or U13872 (N_13872,N_9593,N_11979);
or U13873 (N_13873,N_11936,N_9045);
or U13874 (N_13874,N_9215,N_11774);
nand U13875 (N_13875,N_10366,N_10900);
and U13876 (N_13876,N_11403,N_9644);
nand U13877 (N_13877,N_10907,N_9081);
nor U13878 (N_13878,N_9666,N_11713);
nand U13879 (N_13879,N_10026,N_9311);
nor U13880 (N_13880,N_9326,N_11674);
and U13881 (N_13881,N_9050,N_9928);
or U13882 (N_13882,N_9049,N_11160);
xor U13883 (N_13883,N_9177,N_10129);
or U13884 (N_13884,N_9224,N_11869);
nand U13885 (N_13885,N_10557,N_9266);
nand U13886 (N_13886,N_11365,N_11723);
nand U13887 (N_13887,N_9432,N_10251);
and U13888 (N_13888,N_9428,N_10021);
nand U13889 (N_13889,N_11124,N_11749);
and U13890 (N_13890,N_10536,N_11671);
or U13891 (N_13891,N_11167,N_11422);
or U13892 (N_13892,N_9061,N_11839);
nand U13893 (N_13893,N_9236,N_11416);
or U13894 (N_13894,N_11836,N_11899);
or U13895 (N_13895,N_10292,N_10300);
nor U13896 (N_13896,N_9205,N_9228);
or U13897 (N_13897,N_9331,N_9493);
nor U13898 (N_13898,N_11848,N_9322);
nand U13899 (N_13899,N_9958,N_9509);
xor U13900 (N_13900,N_10631,N_11464);
nand U13901 (N_13901,N_11437,N_9146);
nor U13902 (N_13902,N_11606,N_11883);
and U13903 (N_13903,N_10141,N_10839);
nand U13904 (N_13904,N_10869,N_11715);
nand U13905 (N_13905,N_10621,N_9604);
or U13906 (N_13906,N_10663,N_11046);
or U13907 (N_13907,N_10028,N_9333);
nor U13908 (N_13908,N_9114,N_9189);
nor U13909 (N_13909,N_11754,N_10784);
nor U13910 (N_13910,N_11588,N_10212);
xnor U13911 (N_13911,N_11096,N_9027);
or U13912 (N_13912,N_9886,N_10594);
nand U13913 (N_13913,N_10324,N_10429);
and U13914 (N_13914,N_10368,N_11517);
or U13915 (N_13915,N_11135,N_11056);
nand U13916 (N_13916,N_11200,N_9275);
xnor U13917 (N_13917,N_9632,N_10528);
xor U13918 (N_13918,N_10003,N_11341);
nand U13919 (N_13919,N_10266,N_9307);
or U13920 (N_13920,N_9166,N_9397);
nor U13921 (N_13921,N_9372,N_9178);
nor U13922 (N_13922,N_9305,N_9132);
and U13923 (N_13923,N_11128,N_10272);
xnor U13924 (N_13924,N_10226,N_10190);
and U13925 (N_13925,N_11737,N_10520);
xor U13926 (N_13926,N_9972,N_10201);
nor U13927 (N_13927,N_11195,N_11756);
nand U13928 (N_13928,N_11921,N_10578);
and U13929 (N_13929,N_11524,N_10916);
nor U13930 (N_13930,N_11229,N_11474);
and U13931 (N_13931,N_10007,N_9913);
nand U13932 (N_13932,N_11464,N_9594);
nor U13933 (N_13933,N_10203,N_9689);
nand U13934 (N_13934,N_9954,N_9136);
xor U13935 (N_13935,N_11294,N_10422);
nand U13936 (N_13936,N_11345,N_10064);
nand U13937 (N_13937,N_10123,N_9904);
and U13938 (N_13938,N_10981,N_10533);
and U13939 (N_13939,N_10913,N_9770);
or U13940 (N_13940,N_10692,N_9882);
or U13941 (N_13941,N_9437,N_11825);
nor U13942 (N_13942,N_10410,N_11612);
nand U13943 (N_13943,N_9446,N_9027);
and U13944 (N_13944,N_9683,N_10931);
nand U13945 (N_13945,N_11189,N_11370);
or U13946 (N_13946,N_11007,N_9748);
xor U13947 (N_13947,N_11514,N_9264);
and U13948 (N_13948,N_9447,N_10025);
nand U13949 (N_13949,N_9900,N_10189);
nand U13950 (N_13950,N_11661,N_9402);
nand U13951 (N_13951,N_9593,N_9442);
xor U13952 (N_13952,N_11661,N_9067);
or U13953 (N_13953,N_9836,N_10411);
nand U13954 (N_13954,N_10031,N_11160);
nor U13955 (N_13955,N_10911,N_9493);
nand U13956 (N_13956,N_10637,N_11611);
nor U13957 (N_13957,N_11731,N_11292);
and U13958 (N_13958,N_9119,N_11131);
nor U13959 (N_13959,N_9692,N_10612);
and U13960 (N_13960,N_10908,N_11171);
nor U13961 (N_13961,N_11580,N_11689);
nand U13962 (N_13962,N_11642,N_9368);
and U13963 (N_13963,N_10566,N_10630);
nand U13964 (N_13964,N_11714,N_9686);
nand U13965 (N_13965,N_11074,N_9250);
or U13966 (N_13966,N_11772,N_9131);
or U13967 (N_13967,N_9836,N_10047);
or U13968 (N_13968,N_10972,N_10684);
and U13969 (N_13969,N_11759,N_10785);
or U13970 (N_13970,N_11440,N_9134);
nand U13971 (N_13971,N_10825,N_9809);
nand U13972 (N_13972,N_11916,N_11812);
or U13973 (N_13973,N_9997,N_11351);
nor U13974 (N_13974,N_11805,N_9186);
xor U13975 (N_13975,N_9726,N_10750);
or U13976 (N_13976,N_9933,N_9668);
or U13977 (N_13977,N_11255,N_9554);
and U13978 (N_13978,N_9805,N_10231);
nand U13979 (N_13979,N_9492,N_10796);
and U13980 (N_13980,N_10817,N_11695);
and U13981 (N_13981,N_11878,N_11558);
or U13982 (N_13982,N_9411,N_11956);
and U13983 (N_13983,N_11697,N_9866);
nand U13984 (N_13984,N_11944,N_10928);
nor U13985 (N_13985,N_9567,N_10839);
or U13986 (N_13986,N_10491,N_10564);
and U13987 (N_13987,N_9530,N_11119);
and U13988 (N_13988,N_11826,N_9448);
nor U13989 (N_13989,N_10646,N_10279);
or U13990 (N_13990,N_10094,N_10769);
or U13991 (N_13991,N_10648,N_10089);
or U13992 (N_13992,N_11343,N_9669);
xnor U13993 (N_13993,N_10615,N_10089);
and U13994 (N_13994,N_10852,N_11032);
nor U13995 (N_13995,N_11769,N_10142);
and U13996 (N_13996,N_11348,N_9171);
nand U13997 (N_13997,N_11966,N_11642);
or U13998 (N_13998,N_11761,N_9213);
or U13999 (N_13999,N_10938,N_9984);
and U14000 (N_14000,N_11168,N_9682);
nor U14001 (N_14001,N_10907,N_10379);
or U14002 (N_14002,N_10473,N_10701);
or U14003 (N_14003,N_11172,N_11099);
nand U14004 (N_14004,N_10407,N_10736);
or U14005 (N_14005,N_11197,N_11451);
and U14006 (N_14006,N_10521,N_9166);
or U14007 (N_14007,N_9762,N_10634);
nor U14008 (N_14008,N_11862,N_10982);
nand U14009 (N_14009,N_9462,N_11637);
or U14010 (N_14010,N_10293,N_11334);
xor U14011 (N_14011,N_11204,N_10459);
nor U14012 (N_14012,N_10224,N_11256);
xor U14013 (N_14013,N_10924,N_10361);
and U14014 (N_14014,N_10734,N_10130);
nand U14015 (N_14015,N_11795,N_11019);
nand U14016 (N_14016,N_10812,N_11901);
nor U14017 (N_14017,N_9008,N_9596);
nand U14018 (N_14018,N_11033,N_10683);
nand U14019 (N_14019,N_10546,N_11183);
and U14020 (N_14020,N_9520,N_9731);
nand U14021 (N_14021,N_11140,N_9308);
and U14022 (N_14022,N_9596,N_9363);
nor U14023 (N_14023,N_9255,N_10833);
nand U14024 (N_14024,N_11314,N_9016);
nand U14025 (N_14025,N_10149,N_10379);
nand U14026 (N_14026,N_10078,N_11166);
and U14027 (N_14027,N_11599,N_11334);
nor U14028 (N_14028,N_10691,N_10034);
nor U14029 (N_14029,N_11578,N_9546);
or U14030 (N_14030,N_11759,N_9198);
xnor U14031 (N_14031,N_11070,N_10624);
xnor U14032 (N_14032,N_9442,N_11040);
nor U14033 (N_14033,N_10906,N_9020);
or U14034 (N_14034,N_10137,N_11270);
or U14035 (N_14035,N_10600,N_9373);
nor U14036 (N_14036,N_10716,N_9235);
nor U14037 (N_14037,N_11664,N_11075);
xnor U14038 (N_14038,N_10799,N_11855);
nor U14039 (N_14039,N_11079,N_9375);
or U14040 (N_14040,N_10246,N_9646);
and U14041 (N_14041,N_11452,N_10559);
nand U14042 (N_14042,N_11781,N_9981);
nor U14043 (N_14043,N_10873,N_10360);
nand U14044 (N_14044,N_9530,N_9586);
nor U14045 (N_14045,N_10795,N_9725);
or U14046 (N_14046,N_10767,N_11620);
and U14047 (N_14047,N_9555,N_10554);
and U14048 (N_14048,N_9400,N_9207);
nor U14049 (N_14049,N_11325,N_11636);
and U14050 (N_14050,N_11235,N_9119);
or U14051 (N_14051,N_9333,N_9951);
or U14052 (N_14052,N_9892,N_11075);
and U14053 (N_14053,N_10344,N_9860);
nand U14054 (N_14054,N_9136,N_9928);
nand U14055 (N_14055,N_9627,N_11510);
or U14056 (N_14056,N_9737,N_9764);
and U14057 (N_14057,N_9414,N_9975);
or U14058 (N_14058,N_9265,N_10526);
xnor U14059 (N_14059,N_9864,N_10940);
nor U14060 (N_14060,N_11476,N_9611);
nand U14061 (N_14061,N_10184,N_10960);
or U14062 (N_14062,N_9169,N_11547);
nor U14063 (N_14063,N_10760,N_9600);
nor U14064 (N_14064,N_11725,N_10726);
nand U14065 (N_14065,N_10064,N_10390);
nand U14066 (N_14066,N_11379,N_11747);
and U14067 (N_14067,N_11885,N_9624);
or U14068 (N_14068,N_9249,N_9046);
nand U14069 (N_14069,N_9759,N_9341);
nor U14070 (N_14070,N_10582,N_11496);
and U14071 (N_14071,N_10560,N_10289);
and U14072 (N_14072,N_11953,N_10461);
xnor U14073 (N_14073,N_11276,N_11986);
or U14074 (N_14074,N_10013,N_9944);
xor U14075 (N_14075,N_9613,N_10009);
and U14076 (N_14076,N_11944,N_11418);
and U14077 (N_14077,N_10611,N_9101);
xor U14078 (N_14078,N_9824,N_9807);
nand U14079 (N_14079,N_11868,N_11965);
xor U14080 (N_14080,N_10437,N_10074);
nand U14081 (N_14081,N_9387,N_11484);
xor U14082 (N_14082,N_9445,N_10223);
and U14083 (N_14083,N_10355,N_9696);
nand U14084 (N_14084,N_10874,N_9963);
and U14085 (N_14085,N_11065,N_11369);
or U14086 (N_14086,N_11106,N_9195);
nor U14087 (N_14087,N_9280,N_10959);
nor U14088 (N_14088,N_9334,N_9336);
nand U14089 (N_14089,N_10704,N_9355);
or U14090 (N_14090,N_9909,N_10438);
nand U14091 (N_14091,N_11265,N_9092);
nand U14092 (N_14092,N_11595,N_9657);
nor U14093 (N_14093,N_10010,N_10476);
or U14094 (N_14094,N_10610,N_9714);
nand U14095 (N_14095,N_9559,N_11436);
and U14096 (N_14096,N_11891,N_10659);
nor U14097 (N_14097,N_11672,N_11973);
and U14098 (N_14098,N_11030,N_10484);
and U14099 (N_14099,N_11918,N_9556);
xnor U14100 (N_14100,N_9623,N_10793);
and U14101 (N_14101,N_11787,N_11829);
and U14102 (N_14102,N_10132,N_10825);
or U14103 (N_14103,N_11816,N_10274);
and U14104 (N_14104,N_11913,N_9468);
or U14105 (N_14105,N_10279,N_11870);
nand U14106 (N_14106,N_9468,N_11079);
nor U14107 (N_14107,N_10473,N_10851);
xor U14108 (N_14108,N_9203,N_9567);
nand U14109 (N_14109,N_11762,N_10142);
or U14110 (N_14110,N_11053,N_9127);
or U14111 (N_14111,N_9948,N_10853);
and U14112 (N_14112,N_10577,N_10294);
or U14113 (N_14113,N_9975,N_11871);
or U14114 (N_14114,N_10451,N_11639);
or U14115 (N_14115,N_11188,N_10113);
nand U14116 (N_14116,N_11063,N_9474);
and U14117 (N_14117,N_9721,N_9042);
xnor U14118 (N_14118,N_9904,N_9122);
and U14119 (N_14119,N_10830,N_9900);
or U14120 (N_14120,N_10497,N_10352);
or U14121 (N_14121,N_11057,N_10170);
or U14122 (N_14122,N_11930,N_11518);
and U14123 (N_14123,N_11583,N_11059);
or U14124 (N_14124,N_9214,N_9992);
nand U14125 (N_14125,N_10760,N_11835);
or U14126 (N_14126,N_9965,N_11978);
and U14127 (N_14127,N_9121,N_10114);
nand U14128 (N_14128,N_9630,N_10044);
nand U14129 (N_14129,N_9169,N_10536);
nor U14130 (N_14130,N_11867,N_11413);
and U14131 (N_14131,N_9717,N_10968);
or U14132 (N_14132,N_9041,N_11496);
or U14133 (N_14133,N_10389,N_11143);
or U14134 (N_14134,N_11956,N_9442);
and U14135 (N_14135,N_9074,N_11596);
nor U14136 (N_14136,N_10343,N_10291);
nand U14137 (N_14137,N_10619,N_10716);
xor U14138 (N_14138,N_10003,N_9618);
or U14139 (N_14139,N_9745,N_10591);
nand U14140 (N_14140,N_10795,N_9359);
and U14141 (N_14141,N_10876,N_9549);
nand U14142 (N_14142,N_10284,N_11702);
or U14143 (N_14143,N_10577,N_10339);
and U14144 (N_14144,N_9640,N_10983);
or U14145 (N_14145,N_11387,N_11167);
or U14146 (N_14146,N_10920,N_11638);
nand U14147 (N_14147,N_11166,N_11921);
nor U14148 (N_14148,N_11498,N_10325);
or U14149 (N_14149,N_9234,N_9321);
or U14150 (N_14150,N_9264,N_9643);
or U14151 (N_14151,N_11065,N_10286);
and U14152 (N_14152,N_9563,N_10238);
nand U14153 (N_14153,N_10160,N_11567);
nor U14154 (N_14154,N_9816,N_11412);
nand U14155 (N_14155,N_11025,N_9083);
or U14156 (N_14156,N_10579,N_9359);
nor U14157 (N_14157,N_11558,N_11399);
xor U14158 (N_14158,N_10214,N_11538);
nor U14159 (N_14159,N_9722,N_9325);
nand U14160 (N_14160,N_10764,N_9611);
and U14161 (N_14161,N_10652,N_9384);
nand U14162 (N_14162,N_11798,N_10340);
nor U14163 (N_14163,N_11179,N_11294);
nand U14164 (N_14164,N_9583,N_9193);
and U14165 (N_14165,N_9825,N_11445);
nand U14166 (N_14166,N_9460,N_11906);
nor U14167 (N_14167,N_11416,N_10477);
or U14168 (N_14168,N_11953,N_11329);
nand U14169 (N_14169,N_11520,N_10418);
nand U14170 (N_14170,N_9407,N_9330);
or U14171 (N_14171,N_11828,N_10968);
and U14172 (N_14172,N_10389,N_11222);
and U14173 (N_14173,N_9232,N_10901);
nor U14174 (N_14174,N_11135,N_10996);
nor U14175 (N_14175,N_10606,N_11790);
and U14176 (N_14176,N_9347,N_11495);
or U14177 (N_14177,N_11955,N_11157);
or U14178 (N_14178,N_11982,N_11589);
nand U14179 (N_14179,N_9659,N_10557);
nand U14180 (N_14180,N_11686,N_9082);
xor U14181 (N_14181,N_10317,N_9928);
xor U14182 (N_14182,N_10545,N_11858);
and U14183 (N_14183,N_9623,N_11884);
nor U14184 (N_14184,N_11109,N_10368);
nand U14185 (N_14185,N_11609,N_9471);
or U14186 (N_14186,N_10258,N_9059);
and U14187 (N_14187,N_11632,N_9005);
nor U14188 (N_14188,N_9154,N_11327);
and U14189 (N_14189,N_9351,N_10179);
nor U14190 (N_14190,N_10293,N_9283);
and U14191 (N_14191,N_10121,N_9861);
or U14192 (N_14192,N_10163,N_10857);
nand U14193 (N_14193,N_9861,N_9572);
xnor U14194 (N_14194,N_9269,N_9989);
xnor U14195 (N_14195,N_9856,N_10492);
nand U14196 (N_14196,N_10024,N_10722);
or U14197 (N_14197,N_10576,N_9319);
or U14198 (N_14198,N_9746,N_11353);
nor U14199 (N_14199,N_10430,N_10957);
xor U14200 (N_14200,N_11281,N_9966);
and U14201 (N_14201,N_11012,N_11807);
and U14202 (N_14202,N_11627,N_10806);
and U14203 (N_14203,N_10685,N_9143);
or U14204 (N_14204,N_10138,N_10260);
and U14205 (N_14205,N_11682,N_11546);
nor U14206 (N_14206,N_9589,N_9216);
nand U14207 (N_14207,N_11957,N_10532);
or U14208 (N_14208,N_10501,N_9651);
or U14209 (N_14209,N_10224,N_10945);
nand U14210 (N_14210,N_9680,N_9401);
xor U14211 (N_14211,N_9201,N_11247);
or U14212 (N_14212,N_10787,N_11723);
xnor U14213 (N_14213,N_9274,N_9407);
nand U14214 (N_14214,N_9955,N_10866);
xor U14215 (N_14215,N_11284,N_11734);
and U14216 (N_14216,N_11007,N_10088);
and U14217 (N_14217,N_9279,N_9719);
or U14218 (N_14218,N_10098,N_9634);
nand U14219 (N_14219,N_10773,N_9210);
nor U14220 (N_14220,N_10357,N_9123);
nand U14221 (N_14221,N_11952,N_10403);
or U14222 (N_14222,N_9640,N_9745);
and U14223 (N_14223,N_10640,N_9906);
or U14224 (N_14224,N_9129,N_11644);
or U14225 (N_14225,N_10980,N_10011);
or U14226 (N_14226,N_10968,N_11969);
or U14227 (N_14227,N_9798,N_9818);
xnor U14228 (N_14228,N_10496,N_11635);
xor U14229 (N_14229,N_10579,N_11865);
and U14230 (N_14230,N_11225,N_10447);
and U14231 (N_14231,N_9167,N_11005);
nor U14232 (N_14232,N_11663,N_9298);
nor U14233 (N_14233,N_11071,N_9368);
nor U14234 (N_14234,N_11606,N_10778);
or U14235 (N_14235,N_10654,N_10140);
or U14236 (N_14236,N_9980,N_11893);
or U14237 (N_14237,N_10454,N_10230);
or U14238 (N_14238,N_10088,N_9648);
and U14239 (N_14239,N_11021,N_9552);
or U14240 (N_14240,N_11210,N_11477);
nor U14241 (N_14241,N_11056,N_10417);
or U14242 (N_14242,N_9756,N_9730);
nand U14243 (N_14243,N_10762,N_11819);
nor U14244 (N_14244,N_10171,N_11968);
nor U14245 (N_14245,N_9388,N_11972);
nor U14246 (N_14246,N_10655,N_9895);
nand U14247 (N_14247,N_9617,N_9985);
or U14248 (N_14248,N_11129,N_11180);
nand U14249 (N_14249,N_10096,N_9852);
and U14250 (N_14250,N_9199,N_11503);
nand U14251 (N_14251,N_11737,N_11258);
nand U14252 (N_14252,N_10971,N_10807);
nor U14253 (N_14253,N_9274,N_11465);
and U14254 (N_14254,N_9573,N_10834);
xnor U14255 (N_14255,N_9278,N_9548);
and U14256 (N_14256,N_9778,N_11683);
nor U14257 (N_14257,N_9894,N_11820);
and U14258 (N_14258,N_10814,N_10799);
or U14259 (N_14259,N_11140,N_10656);
and U14260 (N_14260,N_11617,N_9593);
nor U14261 (N_14261,N_10050,N_10045);
or U14262 (N_14262,N_11654,N_9086);
nand U14263 (N_14263,N_10559,N_11310);
and U14264 (N_14264,N_11881,N_11397);
nor U14265 (N_14265,N_10487,N_11566);
or U14266 (N_14266,N_10541,N_11431);
or U14267 (N_14267,N_11909,N_11631);
nand U14268 (N_14268,N_11406,N_11850);
and U14269 (N_14269,N_11320,N_10038);
or U14270 (N_14270,N_9587,N_10408);
and U14271 (N_14271,N_10214,N_9609);
or U14272 (N_14272,N_11854,N_10135);
xor U14273 (N_14273,N_10693,N_9887);
nand U14274 (N_14274,N_9869,N_9957);
or U14275 (N_14275,N_9811,N_10247);
nor U14276 (N_14276,N_11440,N_10880);
or U14277 (N_14277,N_11719,N_10840);
or U14278 (N_14278,N_11291,N_9741);
and U14279 (N_14279,N_11448,N_10273);
nor U14280 (N_14280,N_11185,N_11144);
xor U14281 (N_14281,N_9283,N_9125);
or U14282 (N_14282,N_10214,N_11138);
xnor U14283 (N_14283,N_10630,N_10655);
nor U14284 (N_14284,N_9841,N_9901);
nand U14285 (N_14285,N_9200,N_11041);
nand U14286 (N_14286,N_11661,N_9695);
and U14287 (N_14287,N_11493,N_11145);
and U14288 (N_14288,N_11711,N_11535);
nand U14289 (N_14289,N_9571,N_9802);
and U14290 (N_14290,N_10376,N_9868);
or U14291 (N_14291,N_11316,N_11399);
xor U14292 (N_14292,N_10430,N_9920);
and U14293 (N_14293,N_9359,N_10006);
nand U14294 (N_14294,N_11168,N_9786);
and U14295 (N_14295,N_11125,N_9093);
nand U14296 (N_14296,N_9630,N_11980);
nand U14297 (N_14297,N_10192,N_10718);
or U14298 (N_14298,N_9780,N_11295);
nor U14299 (N_14299,N_11112,N_9371);
nor U14300 (N_14300,N_11554,N_11265);
and U14301 (N_14301,N_9930,N_9699);
nand U14302 (N_14302,N_11964,N_11815);
nor U14303 (N_14303,N_11805,N_10235);
or U14304 (N_14304,N_10641,N_9202);
and U14305 (N_14305,N_9446,N_10265);
nand U14306 (N_14306,N_11149,N_9002);
or U14307 (N_14307,N_11817,N_11158);
xor U14308 (N_14308,N_10978,N_9302);
xor U14309 (N_14309,N_10486,N_9582);
xnor U14310 (N_14310,N_10577,N_11780);
nor U14311 (N_14311,N_9073,N_9572);
nand U14312 (N_14312,N_11027,N_11598);
or U14313 (N_14313,N_11318,N_10183);
and U14314 (N_14314,N_9705,N_10133);
nor U14315 (N_14315,N_10372,N_10195);
xnor U14316 (N_14316,N_9423,N_9138);
and U14317 (N_14317,N_9853,N_10251);
and U14318 (N_14318,N_10401,N_11826);
nor U14319 (N_14319,N_9005,N_10955);
xor U14320 (N_14320,N_11991,N_11436);
and U14321 (N_14321,N_10838,N_11832);
xnor U14322 (N_14322,N_11643,N_9598);
xnor U14323 (N_14323,N_9364,N_11473);
and U14324 (N_14324,N_10659,N_10430);
xor U14325 (N_14325,N_9730,N_10286);
nor U14326 (N_14326,N_11986,N_9470);
nand U14327 (N_14327,N_9115,N_11480);
and U14328 (N_14328,N_10127,N_10129);
nor U14329 (N_14329,N_11561,N_9500);
nand U14330 (N_14330,N_10109,N_9297);
nand U14331 (N_14331,N_9583,N_9399);
or U14332 (N_14332,N_10559,N_10476);
or U14333 (N_14333,N_9257,N_10965);
nor U14334 (N_14334,N_9892,N_10679);
nor U14335 (N_14335,N_11941,N_11099);
xnor U14336 (N_14336,N_9128,N_10847);
or U14337 (N_14337,N_11997,N_9268);
nand U14338 (N_14338,N_11953,N_11236);
nand U14339 (N_14339,N_10039,N_9745);
and U14340 (N_14340,N_10967,N_11586);
or U14341 (N_14341,N_10301,N_11678);
nand U14342 (N_14342,N_9366,N_9268);
and U14343 (N_14343,N_11494,N_9443);
nand U14344 (N_14344,N_11050,N_10901);
nand U14345 (N_14345,N_11499,N_9719);
nand U14346 (N_14346,N_9782,N_10094);
nand U14347 (N_14347,N_10250,N_10319);
nand U14348 (N_14348,N_9563,N_9047);
nor U14349 (N_14349,N_9643,N_11295);
nand U14350 (N_14350,N_11518,N_9416);
nor U14351 (N_14351,N_10326,N_10087);
and U14352 (N_14352,N_9706,N_11301);
nand U14353 (N_14353,N_9014,N_11993);
or U14354 (N_14354,N_11007,N_10394);
nor U14355 (N_14355,N_11464,N_9719);
and U14356 (N_14356,N_11434,N_10376);
and U14357 (N_14357,N_11306,N_11525);
and U14358 (N_14358,N_10871,N_10768);
xnor U14359 (N_14359,N_10941,N_11330);
nand U14360 (N_14360,N_11787,N_9494);
nor U14361 (N_14361,N_9746,N_11807);
nor U14362 (N_14362,N_9883,N_10014);
nor U14363 (N_14363,N_11398,N_11479);
nor U14364 (N_14364,N_10004,N_11161);
or U14365 (N_14365,N_9454,N_11951);
nor U14366 (N_14366,N_11691,N_11167);
nor U14367 (N_14367,N_9642,N_9917);
nor U14368 (N_14368,N_11541,N_11495);
nand U14369 (N_14369,N_9628,N_11218);
nor U14370 (N_14370,N_10966,N_11859);
nor U14371 (N_14371,N_11159,N_9661);
or U14372 (N_14372,N_10866,N_9647);
and U14373 (N_14373,N_9944,N_10634);
nor U14374 (N_14374,N_10629,N_10018);
nor U14375 (N_14375,N_11741,N_11573);
or U14376 (N_14376,N_9132,N_10772);
nor U14377 (N_14377,N_11941,N_11799);
or U14378 (N_14378,N_9448,N_10951);
nor U14379 (N_14379,N_10030,N_11965);
nor U14380 (N_14380,N_10674,N_11898);
nor U14381 (N_14381,N_9774,N_10061);
nand U14382 (N_14382,N_9520,N_11330);
and U14383 (N_14383,N_11001,N_11923);
or U14384 (N_14384,N_9421,N_11297);
or U14385 (N_14385,N_10564,N_10770);
nand U14386 (N_14386,N_11853,N_11637);
nand U14387 (N_14387,N_9876,N_9869);
nand U14388 (N_14388,N_9696,N_11971);
and U14389 (N_14389,N_10359,N_10561);
nor U14390 (N_14390,N_11061,N_11603);
nor U14391 (N_14391,N_10991,N_11946);
nand U14392 (N_14392,N_9264,N_10740);
or U14393 (N_14393,N_10150,N_9586);
nand U14394 (N_14394,N_11800,N_10365);
or U14395 (N_14395,N_10669,N_10659);
nor U14396 (N_14396,N_9734,N_9621);
nor U14397 (N_14397,N_10133,N_9146);
nor U14398 (N_14398,N_9825,N_10835);
nor U14399 (N_14399,N_11760,N_9624);
nor U14400 (N_14400,N_10721,N_11320);
or U14401 (N_14401,N_9864,N_10827);
and U14402 (N_14402,N_9495,N_10151);
or U14403 (N_14403,N_11922,N_10829);
nor U14404 (N_14404,N_9048,N_11011);
nand U14405 (N_14405,N_10958,N_11548);
nor U14406 (N_14406,N_11389,N_10968);
or U14407 (N_14407,N_11763,N_10374);
nand U14408 (N_14408,N_10673,N_9712);
nand U14409 (N_14409,N_9810,N_9571);
nor U14410 (N_14410,N_9941,N_9488);
nand U14411 (N_14411,N_9368,N_9638);
or U14412 (N_14412,N_9165,N_11888);
or U14413 (N_14413,N_9857,N_10896);
and U14414 (N_14414,N_9784,N_9307);
or U14415 (N_14415,N_10444,N_11119);
nand U14416 (N_14416,N_9994,N_11704);
or U14417 (N_14417,N_10298,N_11661);
nor U14418 (N_14418,N_9786,N_9472);
or U14419 (N_14419,N_9365,N_9139);
nor U14420 (N_14420,N_11745,N_10466);
nor U14421 (N_14421,N_11098,N_10772);
and U14422 (N_14422,N_9788,N_11544);
or U14423 (N_14423,N_11307,N_11144);
or U14424 (N_14424,N_10275,N_9312);
nand U14425 (N_14425,N_9088,N_10469);
xor U14426 (N_14426,N_9291,N_9120);
and U14427 (N_14427,N_9276,N_10233);
nor U14428 (N_14428,N_10402,N_9238);
nand U14429 (N_14429,N_11839,N_9338);
and U14430 (N_14430,N_9092,N_10169);
nand U14431 (N_14431,N_10864,N_11945);
and U14432 (N_14432,N_10241,N_11093);
or U14433 (N_14433,N_10347,N_10448);
and U14434 (N_14434,N_10354,N_9664);
xnor U14435 (N_14435,N_11847,N_11131);
and U14436 (N_14436,N_10549,N_11404);
or U14437 (N_14437,N_10839,N_11448);
nor U14438 (N_14438,N_9313,N_11830);
nor U14439 (N_14439,N_11840,N_10004);
nand U14440 (N_14440,N_9776,N_10338);
nor U14441 (N_14441,N_11878,N_11345);
and U14442 (N_14442,N_9918,N_11019);
or U14443 (N_14443,N_11001,N_10206);
xor U14444 (N_14444,N_9812,N_11702);
nor U14445 (N_14445,N_11004,N_10977);
nor U14446 (N_14446,N_11427,N_9009);
or U14447 (N_14447,N_11231,N_10289);
or U14448 (N_14448,N_11478,N_11551);
or U14449 (N_14449,N_10005,N_11337);
and U14450 (N_14450,N_9904,N_9230);
or U14451 (N_14451,N_9177,N_10871);
nand U14452 (N_14452,N_10925,N_11743);
or U14453 (N_14453,N_10603,N_9803);
and U14454 (N_14454,N_9644,N_9759);
nor U14455 (N_14455,N_11122,N_11178);
nand U14456 (N_14456,N_9347,N_10215);
xor U14457 (N_14457,N_11340,N_9846);
nor U14458 (N_14458,N_9859,N_11803);
or U14459 (N_14459,N_9657,N_9333);
nor U14460 (N_14460,N_11735,N_11211);
nor U14461 (N_14461,N_11098,N_9904);
and U14462 (N_14462,N_10099,N_10447);
and U14463 (N_14463,N_11411,N_9026);
and U14464 (N_14464,N_11816,N_9275);
and U14465 (N_14465,N_10710,N_9810);
nand U14466 (N_14466,N_9240,N_11391);
and U14467 (N_14467,N_11064,N_11107);
and U14468 (N_14468,N_10510,N_11283);
nor U14469 (N_14469,N_10088,N_10820);
or U14470 (N_14470,N_10237,N_9142);
nor U14471 (N_14471,N_9789,N_9124);
or U14472 (N_14472,N_10458,N_10511);
xnor U14473 (N_14473,N_10818,N_9031);
and U14474 (N_14474,N_10724,N_11940);
nor U14475 (N_14475,N_11926,N_9035);
or U14476 (N_14476,N_9090,N_9253);
nand U14477 (N_14477,N_11164,N_11445);
and U14478 (N_14478,N_9062,N_11244);
and U14479 (N_14479,N_10351,N_11850);
nand U14480 (N_14480,N_9833,N_11303);
nand U14481 (N_14481,N_11076,N_11147);
nor U14482 (N_14482,N_9796,N_10089);
nor U14483 (N_14483,N_10219,N_10736);
nor U14484 (N_14484,N_9744,N_9097);
nand U14485 (N_14485,N_10085,N_9640);
nand U14486 (N_14486,N_11082,N_10770);
or U14487 (N_14487,N_10075,N_9245);
nand U14488 (N_14488,N_10993,N_11042);
xnor U14489 (N_14489,N_9837,N_10734);
nor U14490 (N_14490,N_10676,N_10922);
or U14491 (N_14491,N_10047,N_9069);
or U14492 (N_14492,N_10421,N_9006);
or U14493 (N_14493,N_9606,N_10754);
or U14494 (N_14494,N_11230,N_9942);
or U14495 (N_14495,N_9221,N_11336);
and U14496 (N_14496,N_10199,N_11246);
or U14497 (N_14497,N_11083,N_9192);
or U14498 (N_14498,N_10790,N_9932);
nor U14499 (N_14499,N_10949,N_10330);
nor U14500 (N_14500,N_11019,N_11940);
nand U14501 (N_14501,N_10804,N_9944);
or U14502 (N_14502,N_9098,N_9859);
nand U14503 (N_14503,N_9001,N_10739);
or U14504 (N_14504,N_11080,N_10973);
nand U14505 (N_14505,N_9799,N_9148);
and U14506 (N_14506,N_9685,N_10348);
nand U14507 (N_14507,N_9074,N_10293);
or U14508 (N_14508,N_10080,N_11852);
nor U14509 (N_14509,N_9807,N_10556);
nand U14510 (N_14510,N_9217,N_9332);
or U14511 (N_14511,N_9058,N_9991);
nor U14512 (N_14512,N_9024,N_10694);
or U14513 (N_14513,N_11132,N_9403);
nor U14514 (N_14514,N_10179,N_11991);
nand U14515 (N_14515,N_11546,N_9903);
nor U14516 (N_14516,N_11265,N_10580);
xnor U14517 (N_14517,N_9196,N_10110);
xnor U14518 (N_14518,N_9310,N_11866);
nand U14519 (N_14519,N_10297,N_11350);
and U14520 (N_14520,N_9803,N_10738);
and U14521 (N_14521,N_10844,N_9210);
nor U14522 (N_14522,N_9183,N_9560);
or U14523 (N_14523,N_9783,N_11630);
nand U14524 (N_14524,N_9732,N_9130);
nor U14525 (N_14525,N_9913,N_10427);
nor U14526 (N_14526,N_10210,N_10425);
nor U14527 (N_14527,N_9153,N_11001);
nand U14528 (N_14528,N_11971,N_10844);
or U14529 (N_14529,N_10268,N_9114);
or U14530 (N_14530,N_9102,N_11720);
and U14531 (N_14531,N_9296,N_10152);
or U14532 (N_14532,N_9161,N_11957);
or U14533 (N_14533,N_10448,N_9946);
nor U14534 (N_14534,N_10536,N_10680);
nor U14535 (N_14535,N_10655,N_10573);
nor U14536 (N_14536,N_10663,N_9040);
nor U14537 (N_14537,N_11591,N_11424);
or U14538 (N_14538,N_9272,N_11798);
and U14539 (N_14539,N_9323,N_11586);
and U14540 (N_14540,N_11024,N_10801);
nand U14541 (N_14541,N_10128,N_10889);
nor U14542 (N_14542,N_10704,N_9767);
and U14543 (N_14543,N_9258,N_10166);
nor U14544 (N_14544,N_10874,N_9677);
or U14545 (N_14545,N_9086,N_10186);
or U14546 (N_14546,N_11133,N_10257);
xnor U14547 (N_14547,N_10549,N_11522);
and U14548 (N_14548,N_9375,N_9170);
xor U14549 (N_14549,N_11440,N_9123);
or U14550 (N_14550,N_10289,N_11085);
and U14551 (N_14551,N_10920,N_10557);
xnor U14552 (N_14552,N_9240,N_11891);
nor U14553 (N_14553,N_9422,N_11232);
nand U14554 (N_14554,N_9459,N_9480);
xnor U14555 (N_14555,N_10592,N_10202);
nand U14556 (N_14556,N_11715,N_9713);
nand U14557 (N_14557,N_11818,N_10445);
nor U14558 (N_14558,N_9403,N_10662);
nand U14559 (N_14559,N_10612,N_11982);
or U14560 (N_14560,N_10834,N_11685);
xor U14561 (N_14561,N_11670,N_9041);
nor U14562 (N_14562,N_9148,N_10057);
nand U14563 (N_14563,N_10646,N_9194);
nor U14564 (N_14564,N_11033,N_9081);
nand U14565 (N_14565,N_11562,N_10085);
nand U14566 (N_14566,N_9443,N_9725);
nor U14567 (N_14567,N_11809,N_11007);
nand U14568 (N_14568,N_10957,N_9866);
xor U14569 (N_14569,N_9995,N_9941);
and U14570 (N_14570,N_9927,N_9058);
nor U14571 (N_14571,N_10593,N_9985);
and U14572 (N_14572,N_9609,N_11168);
and U14573 (N_14573,N_10663,N_10774);
and U14574 (N_14574,N_11155,N_11510);
nand U14575 (N_14575,N_9058,N_9973);
nand U14576 (N_14576,N_9033,N_11042);
or U14577 (N_14577,N_9287,N_11145);
or U14578 (N_14578,N_11660,N_10178);
nor U14579 (N_14579,N_11322,N_10592);
nor U14580 (N_14580,N_11121,N_11830);
or U14581 (N_14581,N_9677,N_11636);
and U14582 (N_14582,N_10986,N_11747);
nand U14583 (N_14583,N_9988,N_11643);
nand U14584 (N_14584,N_10207,N_11005);
nand U14585 (N_14585,N_9914,N_11917);
nand U14586 (N_14586,N_11971,N_10384);
nand U14587 (N_14587,N_11099,N_10449);
and U14588 (N_14588,N_9091,N_11767);
and U14589 (N_14589,N_10169,N_9060);
or U14590 (N_14590,N_10716,N_10615);
nand U14591 (N_14591,N_10581,N_11190);
nand U14592 (N_14592,N_10085,N_11524);
nor U14593 (N_14593,N_10461,N_11813);
or U14594 (N_14594,N_9255,N_10575);
and U14595 (N_14595,N_11716,N_9799);
or U14596 (N_14596,N_9060,N_9258);
nand U14597 (N_14597,N_10631,N_11741);
nand U14598 (N_14598,N_10796,N_11583);
or U14599 (N_14599,N_11101,N_11492);
and U14600 (N_14600,N_9333,N_9133);
and U14601 (N_14601,N_10405,N_10410);
and U14602 (N_14602,N_11985,N_9511);
xor U14603 (N_14603,N_11681,N_9074);
nand U14604 (N_14604,N_9232,N_10572);
and U14605 (N_14605,N_9373,N_9889);
and U14606 (N_14606,N_10710,N_9635);
nor U14607 (N_14607,N_10596,N_11997);
nand U14608 (N_14608,N_10019,N_11119);
and U14609 (N_14609,N_9654,N_10856);
or U14610 (N_14610,N_10429,N_11506);
nand U14611 (N_14611,N_11567,N_11723);
or U14612 (N_14612,N_10448,N_9254);
nor U14613 (N_14613,N_10263,N_10252);
nand U14614 (N_14614,N_9249,N_11965);
or U14615 (N_14615,N_11397,N_9026);
nor U14616 (N_14616,N_11540,N_10386);
or U14617 (N_14617,N_10814,N_11824);
nor U14618 (N_14618,N_9829,N_9861);
xnor U14619 (N_14619,N_9024,N_9044);
or U14620 (N_14620,N_9703,N_11421);
nor U14621 (N_14621,N_11251,N_10224);
nor U14622 (N_14622,N_10847,N_10103);
nand U14623 (N_14623,N_10175,N_9603);
nand U14624 (N_14624,N_9961,N_11211);
and U14625 (N_14625,N_9489,N_10352);
and U14626 (N_14626,N_9247,N_10817);
and U14627 (N_14627,N_9055,N_9391);
or U14628 (N_14628,N_11577,N_10423);
nand U14629 (N_14629,N_9987,N_11480);
or U14630 (N_14630,N_10141,N_9125);
nand U14631 (N_14631,N_11129,N_11605);
nor U14632 (N_14632,N_9937,N_9497);
xnor U14633 (N_14633,N_9095,N_9233);
and U14634 (N_14634,N_11250,N_11140);
nor U14635 (N_14635,N_11712,N_10869);
nand U14636 (N_14636,N_9493,N_10868);
or U14637 (N_14637,N_9913,N_9326);
and U14638 (N_14638,N_9835,N_10377);
nor U14639 (N_14639,N_9721,N_9519);
nand U14640 (N_14640,N_9025,N_10035);
xnor U14641 (N_14641,N_9425,N_9071);
nand U14642 (N_14642,N_9190,N_9857);
nor U14643 (N_14643,N_10868,N_11438);
nor U14644 (N_14644,N_11381,N_10458);
xnor U14645 (N_14645,N_11108,N_11457);
and U14646 (N_14646,N_9369,N_11108);
and U14647 (N_14647,N_10385,N_9939);
nand U14648 (N_14648,N_9451,N_9408);
or U14649 (N_14649,N_10932,N_10357);
and U14650 (N_14650,N_9224,N_11325);
nor U14651 (N_14651,N_11389,N_10939);
nand U14652 (N_14652,N_9707,N_10877);
nand U14653 (N_14653,N_11491,N_9273);
or U14654 (N_14654,N_9038,N_11121);
nor U14655 (N_14655,N_9190,N_11626);
and U14656 (N_14656,N_11786,N_11204);
nand U14657 (N_14657,N_11801,N_11433);
or U14658 (N_14658,N_9500,N_11351);
nand U14659 (N_14659,N_10471,N_11773);
nor U14660 (N_14660,N_10824,N_9664);
or U14661 (N_14661,N_10663,N_10757);
nor U14662 (N_14662,N_11293,N_9232);
xnor U14663 (N_14663,N_11435,N_9942);
or U14664 (N_14664,N_11111,N_11159);
or U14665 (N_14665,N_10007,N_10777);
nor U14666 (N_14666,N_9799,N_9511);
nand U14667 (N_14667,N_9223,N_11685);
nand U14668 (N_14668,N_9456,N_11241);
or U14669 (N_14669,N_9089,N_11947);
nor U14670 (N_14670,N_11855,N_10033);
xor U14671 (N_14671,N_11646,N_11476);
and U14672 (N_14672,N_9823,N_9387);
xnor U14673 (N_14673,N_10467,N_11078);
or U14674 (N_14674,N_10491,N_10653);
nor U14675 (N_14675,N_9889,N_10998);
and U14676 (N_14676,N_9391,N_9768);
nor U14677 (N_14677,N_9871,N_11595);
and U14678 (N_14678,N_10016,N_9213);
nor U14679 (N_14679,N_9247,N_9058);
nand U14680 (N_14680,N_11512,N_9103);
and U14681 (N_14681,N_9530,N_11057);
nor U14682 (N_14682,N_9296,N_10798);
nand U14683 (N_14683,N_11626,N_9273);
and U14684 (N_14684,N_11053,N_9064);
or U14685 (N_14685,N_9137,N_10784);
or U14686 (N_14686,N_9202,N_11814);
nor U14687 (N_14687,N_9672,N_9813);
xnor U14688 (N_14688,N_9954,N_11553);
nor U14689 (N_14689,N_10032,N_10881);
nor U14690 (N_14690,N_10667,N_10974);
or U14691 (N_14691,N_10706,N_10751);
or U14692 (N_14692,N_10048,N_10132);
nand U14693 (N_14693,N_11223,N_10743);
nor U14694 (N_14694,N_11917,N_10780);
nor U14695 (N_14695,N_9465,N_11761);
nand U14696 (N_14696,N_10808,N_11980);
or U14697 (N_14697,N_9182,N_9321);
and U14698 (N_14698,N_9288,N_10839);
or U14699 (N_14699,N_9120,N_10920);
and U14700 (N_14700,N_9537,N_11505);
nand U14701 (N_14701,N_11418,N_9135);
or U14702 (N_14702,N_10737,N_9262);
xnor U14703 (N_14703,N_9296,N_10274);
nand U14704 (N_14704,N_10032,N_11412);
nand U14705 (N_14705,N_10655,N_9060);
xor U14706 (N_14706,N_10516,N_9626);
nand U14707 (N_14707,N_10777,N_10264);
nand U14708 (N_14708,N_10092,N_9390);
or U14709 (N_14709,N_9366,N_10909);
xor U14710 (N_14710,N_11789,N_10690);
or U14711 (N_14711,N_11386,N_11262);
and U14712 (N_14712,N_11518,N_10977);
nor U14713 (N_14713,N_10299,N_11818);
or U14714 (N_14714,N_11410,N_10765);
nor U14715 (N_14715,N_9977,N_11217);
or U14716 (N_14716,N_11917,N_11962);
nand U14717 (N_14717,N_11037,N_10828);
nand U14718 (N_14718,N_9456,N_10149);
nand U14719 (N_14719,N_11023,N_9014);
nand U14720 (N_14720,N_11964,N_10738);
and U14721 (N_14721,N_9921,N_9207);
and U14722 (N_14722,N_11230,N_9034);
xor U14723 (N_14723,N_10560,N_10210);
xor U14724 (N_14724,N_9018,N_11232);
nor U14725 (N_14725,N_10673,N_9869);
nand U14726 (N_14726,N_10279,N_9055);
xnor U14727 (N_14727,N_11682,N_11044);
or U14728 (N_14728,N_11812,N_10647);
nand U14729 (N_14729,N_10432,N_11540);
and U14730 (N_14730,N_10114,N_9151);
nor U14731 (N_14731,N_10289,N_9260);
nor U14732 (N_14732,N_11580,N_10530);
nor U14733 (N_14733,N_11537,N_9415);
nand U14734 (N_14734,N_11500,N_9105);
or U14735 (N_14735,N_10721,N_11972);
and U14736 (N_14736,N_9438,N_9255);
and U14737 (N_14737,N_9050,N_9912);
nor U14738 (N_14738,N_10126,N_11556);
or U14739 (N_14739,N_10333,N_10954);
or U14740 (N_14740,N_11924,N_9370);
nand U14741 (N_14741,N_10992,N_11969);
or U14742 (N_14742,N_11348,N_10262);
nor U14743 (N_14743,N_10788,N_9064);
nor U14744 (N_14744,N_10589,N_10105);
nand U14745 (N_14745,N_9325,N_10350);
nand U14746 (N_14746,N_11251,N_9189);
nor U14747 (N_14747,N_10992,N_10030);
xnor U14748 (N_14748,N_9413,N_9033);
or U14749 (N_14749,N_9408,N_10713);
nand U14750 (N_14750,N_10348,N_9022);
xnor U14751 (N_14751,N_9292,N_9483);
nand U14752 (N_14752,N_9555,N_9851);
and U14753 (N_14753,N_10456,N_11180);
or U14754 (N_14754,N_11869,N_9374);
and U14755 (N_14755,N_9474,N_11364);
nor U14756 (N_14756,N_11640,N_10474);
and U14757 (N_14757,N_11463,N_10907);
and U14758 (N_14758,N_11212,N_10627);
nand U14759 (N_14759,N_9053,N_11501);
or U14760 (N_14760,N_11054,N_9704);
nand U14761 (N_14761,N_9048,N_11256);
nand U14762 (N_14762,N_11936,N_9019);
nand U14763 (N_14763,N_9915,N_10188);
and U14764 (N_14764,N_9262,N_9619);
or U14765 (N_14765,N_10107,N_11711);
nor U14766 (N_14766,N_9708,N_10658);
nor U14767 (N_14767,N_10557,N_10732);
and U14768 (N_14768,N_9137,N_10711);
nor U14769 (N_14769,N_9225,N_9967);
nand U14770 (N_14770,N_9841,N_11277);
xnor U14771 (N_14771,N_11852,N_9430);
or U14772 (N_14772,N_9600,N_9999);
nand U14773 (N_14773,N_11587,N_11406);
or U14774 (N_14774,N_11744,N_9393);
and U14775 (N_14775,N_11463,N_10375);
and U14776 (N_14776,N_10442,N_10221);
xnor U14777 (N_14777,N_11501,N_10868);
and U14778 (N_14778,N_9384,N_11416);
and U14779 (N_14779,N_10659,N_9875);
nand U14780 (N_14780,N_11043,N_11896);
nor U14781 (N_14781,N_11479,N_10872);
nor U14782 (N_14782,N_11045,N_9772);
or U14783 (N_14783,N_9725,N_11612);
or U14784 (N_14784,N_9338,N_9623);
or U14785 (N_14785,N_11839,N_9904);
nand U14786 (N_14786,N_9900,N_11502);
nor U14787 (N_14787,N_9283,N_11831);
and U14788 (N_14788,N_9363,N_10943);
nor U14789 (N_14789,N_9336,N_10199);
or U14790 (N_14790,N_10596,N_9687);
xor U14791 (N_14791,N_9701,N_9308);
or U14792 (N_14792,N_9096,N_11719);
nand U14793 (N_14793,N_11302,N_9977);
and U14794 (N_14794,N_10269,N_11177);
nand U14795 (N_14795,N_10945,N_9051);
nand U14796 (N_14796,N_10692,N_9433);
nand U14797 (N_14797,N_10733,N_9706);
nor U14798 (N_14798,N_11667,N_9641);
and U14799 (N_14799,N_11326,N_10981);
nor U14800 (N_14800,N_11211,N_11149);
xnor U14801 (N_14801,N_10402,N_9536);
nand U14802 (N_14802,N_9728,N_10922);
and U14803 (N_14803,N_10182,N_11549);
xnor U14804 (N_14804,N_10683,N_9934);
and U14805 (N_14805,N_11258,N_9185);
and U14806 (N_14806,N_11405,N_10816);
xnor U14807 (N_14807,N_9606,N_11975);
or U14808 (N_14808,N_11273,N_11824);
xor U14809 (N_14809,N_11777,N_9672);
xor U14810 (N_14810,N_11512,N_10701);
and U14811 (N_14811,N_11985,N_10054);
and U14812 (N_14812,N_11584,N_11136);
nand U14813 (N_14813,N_10130,N_10225);
xnor U14814 (N_14814,N_10109,N_10012);
and U14815 (N_14815,N_11592,N_9537);
or U14816 (N_14816,N_11625,N_9885);
nand U14817 (N_14817,N_9971,N_11922);
and U14818 (N_14818,N_10017,N_10061);
and U14819 (N_14819,N_11732,N_9342);
and U14820 (N_14820,N_10270,N_11021);
and U14821 (N_14821,N_9589,N_9546);
nor U14822 (N_14822,N_11774,N_10109);
xor U14823 (N_14823,N_10404,N_11124);
and U14824 (N_14824,N_9058,N_9745);
or U14825 (N_14825,N_11992,N_10231);
nor U14826 (N_14826,N_11131,N_10932);
or U14827 (N_14827,N_9799,N_11495);
and U14828 (N_14828,N_9581,N_9141);
nand U14829 (N_14829,N_9920,N_10411);
nand U14830 (N_14830,N_11695,N_10922);
nor U14831 (N_14831,N_10265,N_11015);
xnor U14832 (N_14832,N_10172,N_11837);
or U14833 (N_14833,N_10095,N_10416);
xor U14834 (N_14834,N_11657,N_9256);
nand U14835 (N_14835,N_9150,N_9314);
nand U14836 (N_14836,N_11137,N_10424);
or U14837 (N_14837,N_9446,N_10483);
nor U14838 (N_14838,N_10140,N_11358);
nand U14839 (N_14839,N_10618,N_10762);
nand U14840 (N_14840,N_9127,N_9935);
and U14841 (N_14841,N_9591,N_10156);
nor U14842 (N_14842,N_10253,N_11113);
or U14843 (N_14843,N_11797,N_9535);
nand U14844 (N_14844,N_11150,N_10144);
nor U14845 (N_14845,N_10055,N_11659);
or U14846 (N_14846,N_10807,N_11119);
nor U14847 (N_14847,N_11015,N_9668);
and U14848 (N_14848,N_9993,N_11970);
nor U14849 (N_14849,N_11292,N_10670);
or U14850 (N_14850,N_9334,N_9019);
xor U14851 (N_14851,N_10641,N_10138);
nand U14852 (N_14852,N_10611,N_11324);
nor U14853 (N_14853,N_10427,N_9251);
nand U14854 (N_14854,N_9324,N_11359);
and U14855 (N_14855,N_10253,N_10027);
xnor U14856 (N_14856,N_11484,N_9146);
nor U14857 (N_14857,N_9816,N_11011);
nor U14858 (N_14858,N_10542,N_10583);
xor U14859 (N_14859,N_9364,N_9168);
nor U14860 (N_14860,N_9086,N_9195);
nand U14861 (N_14861,N_9710,N_11538);
or U14862 (N_14862,N_11197,N_11012);
nor U14863 (N_14863,N_9540,N_9679);
and U14864 (N_14864,N_11163,N_11182);
and U14865 (N_14865,N_9977,N_9493);
or U14866 (N_14866,N_10680,N_11587);
nand U14867 (N_14867,N_10366,N_9946);
nand U14868 (N_14868,N_10821,N_11633);
xnor U14869 (N_14869,N_9290,N_10200);
nand U14870 (N_14870,N_11832,N_10875);
or U14871 (N_14871,N_10317,N_11356);
or U14872 (N_14872,N_9281,N_9822);
or U14873 (N_14873,N_11569,N_10575);
or U14874 (N_14874,N_9742,N_9194);
xor U14875 (N_14875,N_10903,N_10522);
nor U14876 (N_14876,N_10505,N_9098);
nand U14877 (N_14877,N_10642,N_11467);
nand U14878 (N_14878,N_9860,N_10964);
nor U14879 (N_14879,N_10185,N_10452);
xor U14880 (N_14880,N_11222,N_9931);
or U14881 (N_14881,N_9352,N_10389);
nand U14882 (N_14882,N_10025,N_10276);
nand U14883 (N_14883,N_11388,N_9152);
and U14884 (N_14884,N_9275,N_10063);
xnor U14885 (N_14885,N_9022,N_10879);
nor U14886 (N_14886,N_9013,N_11980);
or U14887 (N_14887,N_11693,N_10455);
xnor U14888 (N_14888,N_9426,N_10571);
nor U14889 (N_14889,N_11312,N_9666);
nand U14890 (N_14890,N_11478,N_11956);
and U14891 (N_14891,N_9560,N_9380);
xnor U14892 (N_14892,N_11024,N_10393);
and U14893 (N_14893,N_10481,N_10526);
nand U14894 (N_14894,N_11961,N_11745);
nor U14895 (N_14895,N_9128,N_10649);
nand U14896 (N_14896,N_11004,N_9790);
nand U14897 (N_14897,N_9877,N_10518);
nor U14898 (N_14898,N_9465,N_11654);
nor U14899 (N_14899,N_10906,N_10813);
and U14900 (N_14900,N_10985,N_11524);
or U14901 (N_14901,N_9526,N_9987);
and U14902 (N_14902,N_9368,N_11550);
and U14903 (N_14903,N_10145,N_11069);
and U14904 (N_14904,N_11433,N_10021);
or U14905 (N_14905,N_11287,N_10281);
and U14906 (N_14906,N_9531,N_10538);
nand U14907 (N_14907,N_10549,N_9224);
nand U14908 (N_14908,N_10406,N_11678);
and U14909 (N_14909,N_9917,N_10887);
and U14910 (N_14910,N_9830,N_10173);
or U14911 (N_14911,N_9034,N_10962);
or U14912 (N_14912,N_10704,N_10051);
and U14913 (N_14913,N_10167,N_11046);
nand U14914 (N_14914,N_10224,N_9870);
nor U14915 (N_14915,N_9200,N_10974);
nand U14916 (N_14916,N_11953,N_9820);
nand U14917 (N_14917,N_9552,N_10505);
xnor U14918 (N_14918,N_11215,N_9371);
nand U14919 (N_14919,N_10541,N_9198);
or U14920 (N_14920,N_9869,N_11208);
nor U14921 (N_14921,N_11220,N_9184);
xnor U14922 (N_14922,N_11235,N_10608);
or U14923 (N_14923,N_9039,N_10889);
nand U14924 (N_14924,N_10623,N_9157);
nand U14925 (N_14925,N_11892,N_9060);
nand U14926 (N_14926,N_10573,N_11051);
nor U14927 (N_14927,N_9598,N_9708);
nand U14928 (N_14928,N_10397,N_9112);
or U14929 (N_14929,N_9934,N_9894);
xnor U14930 (N_14930,N_11386,N_11443);
and U14931 (N_14931,N_10982,N_9383);
nand U14932 (N_14932,N_11599,N_10412);
nor U14933 (N_14933,N_9719,N_11074);
and U14934 (N_14934,N_11096,N_9251);
and U14935 (N_14935,N_11713,N_9549);
or U14936 (N_14936,N_11282,N_11200);
or U14937 (N_14937,N_11266,N_11850);
nand U14938 (N_14938,N_10338,N_10748);
and U14939 (N_14939,N_11202,N_11141);
and U14940 (N_14940,N_10992,N_11324);
nand U14941 (N_14941,N_11755,N_11959);
nand U14942 (N_14942,N_9579,N_9323);
nor U14943 (N_14943,N_10590,N_10316);
and U14944 (N_14944,N_9502,N_9185);
nor U14945 (N_14945,N_10885,N_10541);
nand U14946 (N_14946,N_9416,N_11329);
and U14947 (N_14947,N_11560,N_10328);
xnor U14948 (N_14948,N_11544,N_10222);
nor U14949 (N_14949,N_11999,N_11852);
nor U14950 (N_14950,N_11352,N_9654);
and U14951 (N_14951,N_9088,N_10778);
or U14952 (N_14952,N_9175,N_11149);
xnor U14953 (N_14953,N_11379,N_10033);
nand U14954 (N_14954,N_10795,N_10627);
nor U14955 (N_14955,N_9033,N_11718);
or U14956 (N_14956,N_9091,N_9234);
and U14957 (N_14957,N_11448,N_11595);
nor U14958 (N_14958,N_10427,N_11900);
nand U14959 (N_14959,N_10572,N_11262);
xor U14960 (N_14960,N_9654,N_11756);
nand U14961 (N_14961,N_9659,N_11316);
nor U14962 (N_14962,N_11980,N_9439);
or U14963 (N_14963,N_10574,N_11381);
and U14964 (N_14964,N_10950,N_11918);
or U14965 (N_14965,N_10382,N_10485);
nor U14966 (N_14966,N_10308,N_10393);
or U14967 (N_14967,N_9628,N_10472);
nor U14968 (N_14968,N_9787,N_9906);
xnor U14969 (N_14969,N_9666,N_9574);
xnor U14970 (N_14970,N_11344,N_9473);
and U14971 (N_14971,N_11850,N_9548);
nor U14972 (N_14972,N_11903,N_10520);
and U14973 (N_14973,N_11996,N_9885);
or U14974 (N_14974,N_9620,N_10770);
nand U14975 (N_14975,N_9570,N_10531);
nand U14976 (N_14976,N_11452,N_9427);
and U14977 (N_14977,N_10126,N_11573);
nor U14978 (N_14978,N_11818,N_9271);
or U14979 (N_14979,N_10199,N_9613);
nand U14980 (N_14980,N_9752,N_10927);
or U14981 (N_14981,N_10634,N_9042);
and U14982 (N_14982,N_9766,N_9159);
and U14983 (N_14983,N_9323,N_10647);
or U14984 (N_14984,N_11893,N_11612);
nor U14985 (N_14985,N_10860,N_11937);
xnor U14986 (N_14986,N_11904,N_11254);
nand U14987 (N_14987,N_11536,N_9200);
and U14988 (N_14988,N_10069,N_10154);
nand U14989 (N_14989,N_9344,N_11384);
and U14990 (N_14990,N_9248,N_9855);
and U14991 (N_14991,N_9896,N_11729);
nand U14992 (N_14992,N_10546,N_9976);
xnor U14993 (N_14993,N_11707,N_10331);
nor U14994 (N_14994,N_11371,N_9583);
or U14995 (N_14995,N_9489,N_10608);
nand U14996 (N_14996,N_9302,N_11638);
nor U14997 (N_14997,N_10672,N_11411);
nand U14998 (N_14998,N_9655,N_11269);
or U14999 (N_14999,N_10511,N_11718);
xor UO_0 (O_0,N_12950,N_13385);
and UO_1 (O_1,N_14569,N_14365);
xor UO_2 (O_2,N_13153,N_12496);
nor UO_3 (O_3,N_13361,N_14710);
and UO_4 (O_4,N_13339,N_14017);
and UO_5 (O_5,N_13424,N_14721);
and UO_6 (O_6,N_14012,N_14744);
and UO_7 (O_7,N_14810,N_12275);
or UO_8 (O_8,N_14548,N_12256);
and UO_9 (O_9,N_12291,N_12387);
nand UO_10 (O_10,N_14795,N_14013);
nor UO_11 (O_11,N_12126,N_12145);
nor UO_12 (O_12,N_14902,N_12238);
nor UO_13 (O_13,N_14245,N_13287);
nand UO_14 (O_14,N_12909,N_14919);
nand UO_15 (O_15,N_13299,N_12357);
xor UO_16 (O_16,N_12107,N_14426);
or UO_17 (O_17,N_13636,N_14461);
or UO_18 (O_18,N_12494,N_12712);
nand UO_19 (O_19,N_14262,N_14661);
or UO_20 (O_20,N_14082,N_12098);
nand UO_21 (O_21,N_12472,N_13133);
or UO_22 (O_22,N_14400,N_12285);
xor UO_23 (O_23,N_13386,N_13030);
or UO_24 (O_24,N_12622,N_13043);
xnor UO_25 (O_25,N_14553,N_12991);
nand UO_26 (O_26,N_14490,N_12488);
or UO_27 (O_27,N_13231,N_14189);
nand UO_28 (O_28,N_13208,N_13304);
or UO_29 (O_29,N_13931,N_12922);
nand UO_30 (O_30,N_12742,N_14059);
nand UO_31 (O_31,N_12842,N_12913);
or UO_32 (O_32,N_12438,N_14107);
nand UO_33 (O_33,N_14255,N_13176);
or UO_34 (O_34,N_12758,N_13178);
or UO_35 (O_35,N_12867,N_12644);
nor UO_36 (O_36,N_12914,N_14971);
nand UO_37 (O_37,N_14544,N_12430);
xor UO_38 (O_38,N_12433,N_13880);
or UO_39 (O_39,N_14364,N_13877);
xnor UO_40 (O_40,N_13051,N_13653);
xnor UO_41 (O_41,N_13130,N_13204);
nor UO_42 (O_42,N_13732,N_13134);
xnor UO_43 (O_43,N_13785,N_13066);
and UO_44 (O_44,N_14417,N_13210);
nand UO_45 (O_45,N_14608,N_13371);
nand UO_46 (O_46,N_13852,N_14446);
or UO_47 (O_47,N_13556,N_13567);
or UO_48 (O_48,N_14429,N_14595);
xnor UO_49 (O_49,N_12590,N_13121);
and UO_50 (O_50,N_13725,N_12095);
and UO_51 (O_51,N_14924,N_14628);
or UO_52 (O_52,N_13892,N_13464);
and UO_53 (O_53,N_12329,N_13158);
nor UO_54 (O_54,N_14979,N_12563);
or UO_55 (O_55,N_12785,N_13702);
and UO_56 (O_56,N_12169,N_13778);
nand UO_57 (O_57,N_12232,N_14787);
nor UO_58 (O_58,N_14805,N_12201);
or UO_59 (O_59,N_13159,N_12760);
xor UO_60 (O_60,N_13705,N_13952);
nor UO_61 (O_61,N_14881,N_13094);
xor UO_62 (O_62,N_14875,N_14237);
nand UO_63 (O_63,N_13920,N_12578);
and UO_64 (O_64,N_13677,N_12980);
and UO_65 (O_65,N_14503,N_14954);
nand UO_66 (O_66,N_13598,N_13316);
or UO_67 (O_67,N_12153,N_12694);
and UO_68 (O_68,N_14662,N_13715);
or UO_69 (O_69,N_14823,N_13274);
nand UO_70 (O_70,N_13654,N_14404);
nor UO_71 (O_71,N_13194,N_12230);
nor UO_72 (O_72,N_12748,N_14127);
and UO_73 (O_73,N_14571,N_14943);
nand UO_74 (O_74,N_13536,N_13675);
nand UO_75 (O_75,N_14444,N_12709);
nand UO_76 (O_76,N_12820,N_13533);
nand UO_77 (O_77,N_13724,N_14858);
or UO_78 (O_78,N_14501,N_14874);
or UO_79 (O_79,N_14181,N_14125);
or UO_80 (O_80,N_13528,N_14148);
and UO_81 (O_81,N_13340,N_13930);
nor UO_82 (O_82,N_13330,N_13729);
nor UO_83 (O_83,N_13844,N_13777);
nand UO_84 (O_84,N_13363,N_13638);
and UO_85 (O_85,N_14754,N_12701);
or UO_86 (O_86,N_14260,N_12612);
nand UO_87 (O_87,N_13879,N_14990);
or UO_88 (O_88,N_12025,N_12405);
nand UO_89 (O_89,N_14287,N_13200);
and UO_90 (O_90,N_12257,N_13649);
nor UO_91 (O_91,N_12354,N_12983);
or UO_92 (O_92,N_14049,N_12425);
nand UO_93 (O_93,N_14132,N_12523);
nand UO_94 (O_94,N_12199,N_14887);
nor UO_95 (O_95,N_13048,N_13755);
or UO_96 (O_96,N_14341,N_14645);
xnor UO_97 (O_97,N_13792,N_13356);
or UO_98 (O_98,N_12152,N_13017);
and UO_99 (O_99,N_14855,N_12575);
nand UO_100 (O_100,N_12930,N_14879);
and UO_101 (O_101,N_14334,N_12318);
or UO_102 (O_102,N_12834,N_13303);
nand UO_103 (O_103,N_14793,N_14817);
nand UO_104 (O_104,N_13397,N_12277);
and UO_105 (O_105,N_12055,N_14983);
nand UO_106 (O_106,N_14032,N_14992);
or UO_107 (O_107,N_12378,N_13587);
nand UO_108 (O_108,N_12455,N_12640);
nor UO_109 (O_109,N_13849,N_13914);
and UO_110 (O_110,N_13375,N_12428);
nand UO_111 (O_111,N_14144,N_13993);
nor UO_112 (O_112,N_13314,N_12822);
nand UO_113 (O_113,N_14796,N_12423);
and UO_114 (O_114,N_13630,N_14854);
or UO_115 (O_115,N_12300,N_12416);
nor UO_116 (O_116,N_12988,N_14438);
nand UO_117 (O_117,N_12131,N_14183);
nor UO_118 (O_118,N_12008,N_13581);
nor UO_119 (O_119,N_14547,N_12422);
xnor UO_120 (O_120,N_14730,N_13582);
and UO_121 (O_121,N_13148,N_12402);
xnor UO_122 (O_122,N_14379,N_12944);
and UO_123 (O_123,N_14213,N_13486);
and UO_124 (O_124,N_12133,N_14207);
nor UO_125 (O_125,N_13593,N_14699);
nand UO_126 (O_126,N_13874,N_12541);
nand UO_127 (O_127,N_14938,N_13881);
nor UO_128 (O_128,N_13129,N_14228);
or UO_129 (O_129,N_14939,N_12332);
nor UO_130 (O_130,N_12029,N_12629);
and UO_131 (O_131,N_13980,N_14118);
or UO_132 (O_132,N_13222,N_12193);
nand UO_133 (O_133,N_12091,N_13747);
nand UO_134 (O_134,N_12485,N_12280);
or UO_135 (O_135,N_14828,N_13232);
and UO_136 (O_136,N_13911,N_13083);
or UO_137 (O_137,N_14169,N_13112);
nor UO_138 (O_138,N_12048,N_12086);
xnor UO_139 (O_139,N_13662,N_13292);
or UO_140 (O_140,N_14358,N_13678);
xnor UO_141 (O_141,N_14980,N_14372);
nand UO_142 (O_142,N_12219,N_14928);
or UO_143 (O_143,N_12030,N_13322);
xnor UO_144 (O_144,N_12075,N_13994);
xor UO_145 (O_145,N_12375,N_12879);
nor UO_146 (O_146,N_12961,N_14987);
or UO_147 (O_147,N_12617,N_13501);
and UO_148 (O_148,N_14981,N_14057);
and UO_149 (O_149,N_12418,N_13012);
nor UO_150 (O_150,N_13984,N_14290);
and UO_151 (O_151,N_12157,N_13191);
nor UO_152 (O_152,N_13426,N_13922);
nand UO_153 (O_153,N_14840,N_13529);
nand UO_154 (O_154,N_13313,N_13864);
or UO_155 (O_155,N_12123,N_14020);
nand UO_156 (O_156,N_13916,N_14582);
or UO_157 (O_157,N_12828,N_14398);
or UO_158 (O_158,N_14425,N_12755);
nand UO_159 (O_159,N_12887,N_13166);
and UO_160 (O_160,N_14653,N_13698);
nand UO_161 (O_161,N_12047,N_13047);
or UO_162 (O_162,N_14682,N_14143);
or UO_163 (O_163,N_13933,N_14532);
nor UO_164 (O_164,N_13589,N_12945);
nor UO_165 (O_165,N_13201,N_12937);
nand UO_166 (O_166,N_14128,N_12090);
nor UO_167 (O_167,N_12396,N_13364);
nor UO_168 (O_168,N_13487,N_14665);
nand UO_169 (O_169,N_14578,N_13910);
nand UO_170 (O_170,N_14014,N_12076);
or UO_171 (O_171,N_13506,N_13218);
and UO_172 (O_172,N_13890,N_14593);
xor UO_173 (O_173,N_13497,N_14027);
or UO_174 (O_174,N_14849,N_13895);
nor UO_175 (O_175,N_14937,N_13409);
or UO_176 (O_176,N_13633,N_12217);
and UO_177 (O_177,N_12907,N_14324);
nand UO_178 (O_178,N_14709,N_14588);
xnor UO_179 (O_179,N_14575,N_12186);
and UO_180 (O_180,N_12643,N_14751);
nand UO_181 (O_181,N_13046,N_13646);
xor UO_182 (O_182,N_14205,N_13077);
and UO_183 (O_183,N_13008,N_12373);
nand UO_184 (O_184,N_12417,N_14918);
nor UO_185 (O_185,N_14089,N_13449);
xor UO_186 (O_186,N_14623,N_13887);
nand UO_187 (O_187,N_12847,N_12733);
nand UO_188 (O_188,N_13557,N_13513);
nand UO_189 (O_189,N_14355,N_13246);
and UO_190 (O_190,N_14516,N_12502);
and UO_191 (O_191,N_12268,N_14515);
or UO_192 (O_192,N_13059,N_12014);
and UO_193 (O_193,N_13642,N_12593);
or UO_194 (O_194,N_14909,N_12018);
nand UO_195 (O_195,N_12779,N_12013);
nand UO_196 (O_196,N_13320,N_12279);
nand UO_197 (O_197,N_12841,N_12895);
and UO_198 (O_198,N_12498,N_12208);
and UO_199 (O_199,N_13087,N_13180);
and UO_200 (O_200,N_13751,N_13522);
xnor UO_201 (O_201,N_13171,N_13081);
and UO_202 (O_202,N_13157,N_14149);
and UO_203 (O_203,N_14440,N_12977);
or UO_204 (O_204,N_13147,N_13885);
nand UO_205 (O_205,N_14244,N_13866);
or UO_206 (O_206,N_14023,N_14778);
xnor UO_207 (O_207,N_12110,N_14815);
xor UO_208 (O_208,N_13762,N_13643);
nand UO_209 (O_209,N_13639,N_14176);
and UO_210 (O_210,N_13305,N_12264);
or UO_211 (O_211,N_13045,N_13746);
xnor UO_212 (O_212,N_12866,N_12549);
and UO_213 (O_213,N_12936,N_13515);
nand UO_214 (O_214,N_12518,N_14996);
and UO_215 (O_215,N_13277,N_13106);
nand UO_216 (O_216,N_12151,N_14455);
or UO_217 (O_217,N_13031,N_13179);
xnor UO_218 (O_218,N_12299,N_12624);
and UO_219 (O_219,N_14413,N_13668);
and UO_220 (O_220,N_12883,N_13987);
nand UO_221 (O_221,N_14742,N_12283);
or UO_222 (O_222,N_12715,N_14015);
nor UO_223 (O_223,N_12311,N_12171);
nor UO_224 (O_224,N_13118,N_12298);
or UO_225 (O_225,N_13215,N_13569);
and UO_226 (O_226,N_12235,N_12835);
or UO_227 (O_227,N_13597,N_12376);
and UO_228 (O_228,N_12960,N_12184);
nand UO_229 (O_229,N_14872,N_14208);
nand UO_230 (O_230,N_13769,N_12105);
xnor UO_231 (O_231,N_13764,N_13604);
nor UO_232 (O_232,N_14008,N_13007);
and UO_233 (O_233,N_13658,N_13050);
nand UO_234 (O_234,N_12522,N_12223);
nor UO_235 (O_235,N_13685,N_12707);
nand UO_236 (O_236,N_13447,N_14789);
nand UO_237 (O_237,N_13056,N_13360);
and UO_238 (O_238,N_13413,N_14367);
or UO_239 (O_239,N_12811,N_14982);
nand UO_240 (O_240,N_14129,N_12435);
or UO_241 (O_241,N_14740,N_14388);
nor UO_242 (O_242,N_13982,N_14408);
nand UO_243 (O_243,N_13956,N_13713);
and UO_244 (O_244,N_14018,N_13467);
and UO_245 (O_245,N_12140,N_13188);
nor UO_246 (O_246,N_14476,N_12252);
nand UO_247 (O_247,N_14399,N_13518);
and UO_248 (O_248,N_14878,N_14487);
or UO_249 (O_249,N_12974,N_12161);
nand UO_250 (O_250,N_12807,N_12539);
and UO_251 (O_251,N_14783,N_12411);
and UO_252 (O_252,N_12984,N_13953);
or UO_253 (O_253,N_14791,N_12971);
nand UO_254 (O_254,N_13635,N_13973);
nor UO_255 (O_255,N_14138,N_14974);
and UO_256 (O_256,N_12069,N_13508);
or UO_257 (O_257,N_12713,N_14322);
or UO_258 (O_258,N_14994,N_14328);
xor UO_259 (O_259,N_13839,N_13527);
nand UO_260 (O_260,N_13794,N_12917);
xnor UO_261 (O_261,N_12393,N_13504);
nor UO_262 (O_262,N_12920,N_14777);
nand UO_263 (O_263,N_13144,N_13369);
or UO_264 (O_264,N_13768,N_12985);
or UO_265 (O_265,N_14812,N_13009);
nor UO_266 (O_266,N_14147,N_12456);
and UO_267 (O_267,N_14293,N_13560);
nand UO_268 (O_268,N_12697,N_12177);
and UO_269 (O_269,N_13122,N_12767);
nand UO_270 (O_270,N_12011,N_12412);
and UO_271 (O_271,N_13950,N_12838);
and UO_272 (O_272,N_13706,N_13132);
nand UO_273 (O_273,N_14093,N_13483);
xnor UO_274 (O_274,N_14901,N_12761);
xnor UO_275 (O_275,N_13760,N_12625);
nor UO_276 (O_276,N_14759,N_12750);
or UO_277 (O_277,N_14882,N_12855);
and UO_278 (O_278,N_12413,N_14256);
nand UO_279 (O_279,N_14660,N_14150);
xor UO_280 (O_280,N_13070,N_12849);
nand UO_281 (O_281,N_12832,N_12964);
nor UO_282 (O_282,N_12739,N_12222);
nand UO_283 (O_283,N_14242,N_13381);
or UO_284 (O_284,N_13152,N_12249);
or UO_285 (O_285,N_14302,N_12946);
and UO_286 (O_286,N_13185,N_13860);
nand UO_287 (O_287,N_13281,N_14312);
or UO_288 (O_288,N_12893,N_14718);
nor UO_289 (O_289,N_14058,N_13544);
or UO_290 (O_290,N_13594,N_14458);
or UO_291 (O_291,N_14473,N_14335);
nand UO_292 (O_292,N_13869,N_14510);
nand UO_293 (O_293,N_13553,N_12108);
nand UO_294 (O_294,N_13595,N_13261);
nor UO_295 (O_295,N_12245,N_12792);
nand UO_296 (O_296,N_12179,N_14268);
nand UO_297 (O_297,N_12253,N_13173);
and UO_298 (O_298,N_14270,N_14507);
or UO_299 (O_299,N_13583,N_14329);
or UO_300 (O_300,N_13970,N_14055);
and UO_301 (O_301,N_13290,N_12554);
and UO_302 (O_302,N_12001,N_13960);
xnor UO_303 (O_303,N_14349,N_14196);
xnor UO_304 (O_304,N_13310,N_12797);
or UO_305 (O_305,N_12512,N_13472);
nand UO_306 (O_306,N_14641,N_12061);
xnor UO_307 (O_307,N_13831,N_14694);
nand UO_308 (O_308,N_13396,N_12198);
nor UO_309 (O_309,N_12328,N_14862);
nor UO_310 (O_310,N_13296,N_12419);
nand UO_311 (O_311,N_12799,N_14463);
nand UO_312 (O_312,N_13688,N_14366);
nor UO_313 (O_313,N_14570,N_14401);
nand UO_314 (O_314,N_13606,N_14637);
and UO_315 (O_315,N_12657,N_14936);
nand UO_316 (O_316,N_12084,N_12642);
nand UO_317 (O_317,N_13298,N_14765);
or UO_318 (O_318,N_14484,N_13532);
nor UO_319 (O_319,N_13523,N_13624);
nand UO_320 (O_320,N_13736,N_12732);
and UO_321 (O_321,N_14871,N_14326);
nand UO_322 (O_322,N_12437,N_12610);
nand UO_323 (O_323,N_13475,N_13207);
or UO_324 (O_324,N_13840,N_14842);
nand UO_325 (O_325,N_12781,N_13610);
and UO_326 (O_326,N_13378,N_13942);
nand UO_327 (O_327,N_14217,N_12060);
nor UO_328 (O_328,N_14827,N_14566);
nor UO_329 (O_329,N_12929,N_14844);
or UO_330 (O_330,N_13803,N_13203);
and UO_331 (O_331,N_12233,N_12440);
nand UO_332 (O_332,N_13875,N_12115);
and UO_333 (O_333,N_14384,N_14542);
nand UO_334 (O_334,N_12756,N_14469);
or UO_335 (O_335,N_12192,N_12035);
and UO_336 (O_336,N_13548,N_14175);
nand UO_337 (O_337,N_13740,N_14738);
nor UO_338 (O_338,N_14830,N_13405);
xnor UO_339 (O_339,N_13433,N_13758);
and UO_340 (O_340,N_13326,N_14346);
and UO_341 (O_341,N_14609,N_14241);
nor UO_342 (O_342,N_12764,N_14917);
nor UO_343 (O_343,N_12730,N_14199);
and UO_344 (O_344,N_13791,N_12475);
nand UO_345 (O_345,N_12336,N_14638);
nor UO_346 (O_346,N_13665,N_14003);
and UO_347 (O_347,N_12821,N_14371);
nand UO_348 (O_348,N_14154,N_13438);
nor UO_349 (O_349,N_12211,N_14177);
or UO_350 (O_350,N_12740,N_14596);
or UO_351 (O_351,N_14382,N_13411);
and UO_352 (O_352,N_12802,N_12400);
xor UO_353 (O_353,N_14838,N_14482);
or UO_354 (O_354,N_12596,N_14356);
and UO_355 (O_355,N_12053,N_12665);
or UO_356 (O_356,N_14927,N_14412);
nor UO_357 (O_357,N_12150,N_14890);
and UO_358 (O_358,N_13871,N_12863);
nor UO_359 (O_359,N_13350,N_12019);
nor UO_360 (O_360,N_12528,N_12609);
xor UO_361 (O_361,N_12774,N_14550);
or UO_362 (O_362,N_13968,N_13941);
nor UO_363 (O_363,N_14377,N_12274);
or UO_364 (O_364,N_14806,N_12386);
and UO_365 (O_365,N_12452,N_14198);
and UO_366 (O_366,N_13079,N_13068);
or UO_367 (O_367,N_14519,N_14449);
nor UO_368 (O_368,N_13123,N_14774);
nand UO_369 (O_369,N_14479,N_12514);
and UO_370 (O_370,N_12087,N_14697);
xnor UO_371 (O_371,N_14215,N_13919);
and UO_372 (O_372,N_12225,N_14826);
and UO_373 (O_373,N_13086,N_12190);
or UO_374 (O_374,N_12228,N_12754);
xor UO_375 (O_375,N_14965,N_13470);
nor UO_376 (O_376,N_13796,N_13223);
or UO_377 (O_377,N_14707,N_12490);
nand UO_378 (O_378,N_13093,N_14362);
xor UO_379 (O_379,N_12982,N_14168);
or UO_380 (O_380,N_13855,N_14693);
and UO_381 (O_381,N_12260,N_12651);
xnor UO_382 (O_382,N_13812,N_12818);
and UO_383 (O_383,N_12202,N_12672);
nor UO_384 (O_384,N_12941,N_13451);
and UO_385 (O_385,N_13141,N_13435);
xnor UO_386 (O_386,N_14145,N_12796);
nor UO_387 (O_387,N_13311,N_12762);
nand UO_388 (O_388,N_14253,N_14866);
nand UO_389 (O_389,N_12766,N_13641);
nor UO_390 (O_390,N_14407,N_13670);
or UO_391 (O_391,N_12517,N_13868);
nor UO_392 (O_392,N_14952,N_12641);
nor UO_393 (O_393,N_13924,N_12689);
nor UO_394 (O_394,N_13393,N_13496);
nor UO_395 (O_395,N_13212,N_13985);
and UO_396 (O_396,N_14822,N_12896);
or UO_397 (O_397,N_13562,N_12392);
and UO_398 (O_398,N_14581,N_13695);
nand UO_399 (O_399,N_13004,N_13739);
nor UO_400 (O_400,N_13285,N_14420);
and UO_401 (O_401,N_12436,N_13731);
nand UO_402 (O_402,N_13591,N_14852);
and UO_403 (O_403,N_13932,N_13437);
or UO_404 (O_404,N_12269,N_13347);
nand UO_405 (O_405,N_13830,N_13734);
or UO_406 (O_406,N_14785,N_12874);
or UO_407 (O_407,N_12585,N_12408);
and UO_408 (O_408,N_13495,N_13154);
or UO_409 (O_409,N_13111,N_13810);
or UO_410 (O_410,N_12505,N_13749);
nand UO_411 (O_411,N_13779,N_13790);
xor UO_412 (O_412,N_12829,N_14000);
nor UO_413 (O_413,N_13935,N_14305);
xnor UO_414 (O_414,N_12331,N_12571);
nand UO_415 (O_415,N_12031,N_14528);
and UO_416 (O_416,N_14026,N_13388);
nor UO_417 (O_417,N_12815,N_14171);
and UO_418 (O_418,N_13632,N_12159);
and UO_419 (O_419,N_12071,N_13319);
and UO_420 (O_420,N_14886,N_13485);
nor UO_421 (O_421,N_12652,N_13867);
nand UO_422 (O_422,N_14223,N_13091);
nand UO_423 (O_423,N_12121,N_12286);
nor UO_424 (O_424,N_14500,N_13843);
and UO_425 (O_425,N_12484,N_12282);
nor UO_426 (O_426,N_13691,N_12906);
or UO_427 (O_427,N_12924,N_12457);
or UO_428 (O_428,N_12825,N_13140);
or UO_429 (O_429,N_14997,N_12716);
or UO_430 (O_430,N_13998,N_12663);
nor UO_431 (O_431,N_14700,N_14834);
or UO_432 (O_432,N_13186,N_13482);
and UO_433 (O_433,N_12586,N_12788);
nor UO_434 (O_434,N_13846,N_12165);
nor UO_435 (O_435,N_14478,N_14843);
or UO_436 (O_436,N_12858,N_13711);
nand UO_437 (O_437,N_12236,N_14188);
nand UO_438 (O_438,N_13989,N_14383);
and UO_439 (O_439,N_12717,N_13344);
nor UO_440 (O_440,N_12749,N_14746);
or UO_441 (O_441,N_14360,N_12784);
nor UO_442 (O_442,N_12602,N_13484);
xnor UO_443 (O_443,N_14466,N_14761);
or UO_444 (O_444,N_13795,N_13255);
and UO_445 (O_445,N_13681,N_14483);
nand UO_446 (O_446,N_13019,N_12744);
nor UO_447 (O_447,N_12827,N_13064);
and UO_448 (O_448,N_14337,N_14405);
xnor UO_449 (O_449,N_14706,N_14678);
and UO_450 (O_450,N_14576,N_14666);
or UO_451 (O_451,N_13833,N_14243);
nor UO_452 (O_452,N_12789,N_12656);
xor UO_453 (O_453,N_14338,N_14941);
xor UO_454 (O_454,N_14319,N_13227);
and UO_455 (O_455,N_14643,N_12662);
nor UO_456 (O_456,N_13219,N_14597);
nor UO_457 (O_457,N_12359,N_14948);
nor UO_458 (O_458,N_12931,N_14279);
xor UO_459 (O_459,N_12857,N_12068);
or UO_460 (O_460,N_12923,N_14495);
nor UO_461 (O_461,N_13052,N_13631);
or UO_462 (O_462,N_13089,N_12466);
nand UO_463 (O_463,N_14139,N_13502);
and UO_464 (O_464,N_12003,N_13494);
or UO_465 (O_465,N_12630,N_13837);
or UO_466 (O_466,N_12989,N_12038);
and UO_467 (O_467,N_14092,N_13826);
nand UO_468 (O_468,N_13707,N_14523);
xor UO_469 (O_469,N_14233,N_13620);
nor UO_470 (O_470,N_14635,N_13139);
and UO_471 (O_471,N_13936,N_13242);
or UO_472 (O_472,N_13683,N_12606);
and UO_473 (O_473,N_14323,N_13689);
xnor UO_474 (O_474,N_14353,N_14736);
nor UO_475 (O_475,N_14191,N_14594);
nor UO_476 (O_476,N_12097,N_14922);
and UO_477 (O_477,N_12458,N_12546);
xnor UO_478 (O_478,N_13854,N_14561);
xnor UO_479 (O_479,N_12246,N_13872);
or UO_480 (O_480,N_13859,N_12163);
and UO_481 (O_481,N_14658,N_12478);
xnor UO_482 (O_482,N_14266,N_12894);
and UO_483 (O_483,N_14031,N_12308);
nor UO_484 (O_484,N_14613,N_12556);
and UO_485 (O_485,N_12022,N_13616);
nand UO_486 (O_486,N_14178,N_12024);
xor UO_487 (O_487,N_12237,N_12362);
or UO_488 (O_488,N_12465,N_14598);
nand UO_489 (O_489,N_14433,N_14564);
or UO_490 (O_490,N_14111,N_12627);
nand UO_491 (O_491,N_13323,N_14048);
nand UO_492 (O_492,N_13126,N_14116);
or UO_493 (O_493,N_13991,N_14640);
nand UO_494 (O_494,N_12925,N_14633);
and UO_495 (O_495,N_13710,N_14010);
nor UO_496 (O_496,N_13808,N_14186);
nor UO_497 (O_497,N_14568,N_12798);
nor UO_498 (O_498,N_13596,N_14527);
nor UO_499 (O_499,N_13551,N_13006);
or UO_500 (O_500,N_13534,N_13542);
and UO_501 (O_501,N_12693,N_14807);
or UO_502 (O_502,N_13835,N_14164);
nand UO_503 (O_503,N_14674,N_14393);
xor UO_504 (O_504,N_13478,N_14257);
and UO_505 (O_505,N_12495,N_12284);
xor UO_506 (O_506,N_12695,N_12614);
or UO_507 (O_507,N_12959,N_13170);
and UO_508 (O_508,N_14540,N_13716);
and UO_509 (O_509,N_12187,N_12875);
xor UO_510 (O_510,N_12322,N_13554);
xnor UO_511 (O_511,N_12613,N_12979);
and UO_512 (O_512,N_14300,N_14766);
nor UO_513 (O_513,N_12720,N_13058);
nand UO_514 (O_514,N_14146,N_14916);
xor UO_515 (O_515,N_13603,N_12853);
xnor UO_516 (O_516,N_12962,N_13499);
or UO_517 (O_517,N_12659,N_12587);
and UO_518 (O_518,N_14447,N_12935);
and UO_519 (O_519,N_14745,N_14976);
or UO_520 (O_520,N_12580,N_14342);
nand UO_521 (O_521,N_12294,N_13380);
or UO_522 (O_522,N_14583,N_12410);
or UO_523 (O_523,N_14261,N_13590);
and UO_524 (O_524,N_12948,N_13213);
and UO_525 (O_525,N_13098,N_13481);
nor UO_526 (O_526,N_13442,N_14239);
nand UO_527 (O_527,N_14820,N_12684);
and UO_528 (O_528,N_13816,N_12653);
and UO_529 (O_529,N_12812,N_12530);
nor UO_530 (O_530,N_14716,N_14359);
nand UO_531 (O_531,N_14663,N_14573);
nand UO_532 (O_532,N_14590,N_13062);
or UO_533 (O_533,N_14068,N_13927);
and UO_534 (O_534,N_14508,N_13726);
nand UO_535 (O_535,N_14786,N_13694);
nor UO_536 (O_536,N_12859,N_13318);
and UO_537 (O_537,N_12787,N_12467);
xnor UO_538 (O_538,N_12940,N_13423);
nor UO_539 (O_539,N_14910,N_12244);
and UO_540 (O_540,N_13545,N_12303);
nor UO_541 (O_541,N_12751,N_12675);
or UO_542 (O_542,N_12350,N_14236);
nand UO_543 (O_543,N_13730,N_13018);
nand UO_544 (O_544,N_12356,N_14967);
nor UO_545 (O_545,N_14309,N_12844);
nor UO_546 (O_546,N_14675,N_14900);
nand UO_547 (O_547,N_14836,N_14950);
or UO_548 (O_548,N_14411,N_12527);
nor UO_549 (O_549,N_12889,N_13561);
or UO_550 (O_550,N_12723,N_12840);
nor UO_551 (O_551,N_13609,N_13269);
nor UO_552 (O_552,N_14727,N_14600);
xnor UO_553 (O_553,N_13468,N_12746);
and UO_554 (O_554,N_14543,N_12584);
nand UO_555 (O_555,N_12506,N_12317);
xnor UO_556 (O_556,N_12234,N_12409);
or UO_557 (O_557,N_13814,N_12453);
and UO_558 (O_558,N_14225,N_14883);
or UO_559 (O_559,N_13002,N_12164);
xnor UO_560 (O_560,N_12080,N_13053);
and UO_561 (O_561,N_12623,N_12852);
nor UO_562 (O_562,N_13799,N_13617);
or UO_563 (O_563,N_13954,N_12065);
nand UO_564 (O_564,N_12667,N_12521);
nor UO_565 (O_565,N_13205,N_14671);
or UO_566 (O_566,N_13366,N_14318);
nand UO_567 (O_567,N_12561,N_13902);
nor UO_568 (O_568,N_14956,N_13955);
and UO_569 (O_569,N_14235,N_13964);
nor UO_570 (O_570,N_14681,N_13801);
or UO_571 (O_571,N_13748,N_12358);
nand UO_572 (O_572,N_13415,N_12015);
and UO_573 (O_573,N_13150,N_12477);
or UO_574 (O_574,N_13977,N_14340);
or UO_575 (O_575,N_13460,N_14285);
nand UO_576 (O_576,N_12990,N_12491);
and UO_577 (O_577,N_14664,N_12391);
nor UO_578 (O_578,N_12388,N_12544);
and UO_579 (O_579,N_13718,N_12010);
xnor UO_580 (O_580,N_13408,N_13028);
and UO_581 (O_581,N_12195,N_12678);
and UO_582 (O_582,N_12891,N_12573);
nor UO_583 (O_583,N_12239,N_12611);
xnor UO_584 (O_584,N_13061,N_14289);
nand UO_585 (O_585,N_14086,N_14354);
nand UO_586 (O_586,N_12509,N_14443);
or UO_587 (O_587,N_13510,N_14465);
or UO_588 (O_588,N_13817,N_13906);
or UO_589 (O_589,N_13085,N_13648);
or UO_590 (O_590,N_12647,N_12324);
nand UO_591 (O_591,N_13605,N_12769);
or UO_592 (O_592,N_13457,N_12231);
or UO_593 (O_593,N_13549,N_14846);
and UO_594 (O_594,N_14480,N_13682);
or UO_595 (O_595,N_14770,N_12724);
or UO_596 (O_596,N_13842,N_12486);
or UO_597 (O_597,N_12101,N_12542);
nand UO_598 (O_598,N_12566,N_14833);
xor UO_599 (O_599,N_13184,N_12594);
or UO_600 (O_600,N_12646,N_12532);
nand UO_601 (O_601,N_13135,N_14656);
nand UO_602 (O_602,N_14995,N_12892);
xnor UO_603 (O_603,N_12515,N_14069);
nor UO_604 (O_604,N_14076,N_14703);
xnor UO_605 (O_605,N_14741,N_14194);
nand UO_606 (O_606,N_12052,N_14567);
and UO_607 (O_607,N_14603,N_13181);
or UO_608 (O_608,N_13332,N_13757);
or UO_609 (O_609,N_13741,N_12531);
xor UO_610 (O_610,N_14102,N_14753);
and UO_611 (O_611,N_14525,N_13573);
and UO_612 (O_612,N_12081,N_14247);
and UO_613 (O_613,N_14333,N_13623);
nand UO_614 (O_614,N_13848,N_13588);
nor UO_615 (O_615,N_13252,N_14368);
nor UO_616 (O_616,N_14115,N_13402);
or UO_617 (O_617,N_13983,N_13996);
and UO_618 (O_618,N_12567,N_14387);
nor UO_619 (O_619,N_12125,N_13637);
or UO_620 (O_620,N_12803,N_13249);
or UO_621 (O_621,N_12999,N_14007);
nor UO_622 (O_622,N_12178,N_12130);
nand UO_623 (O_623,N_14546,N_12598);
or UO_624 (O_624,N_13674,N_13142);
nand UO_625 (O_625,N_12172,N_14839);
nand UO_626 (O_626,N_12552,N_13032);
nor UO_627 (O_627,N_13951,N_14867);
xor UO_628 (O_628,N_14180,N_13579);
or UO_629 (O_629,N_14680,N_14868);
nand UO_630 (O_630,N_14580,N_12993);
and UO_631 (O_631,N_13217,N_14043);
nand UO_632 (O_632,N_14961,N_14712);
and UO_633 (O_633,N_13789,N_12686);
nand UO_634 (O_634,N_12088,N_12942);
nand UO_635 (O_635,N_12188,N_12032);
nand UO_636 (O_636,N_14374,N_12743);
or UO_637 (O_637,N_13090,N_13492);
nor UO_638 (O_638,N_13107,N_12447);
and UO_639 (O_639,N_12072,N_14797);
xnor UO_640 (O_640,N_14348,N_14514);
and UO_641 (O_641,N_14397,N_14631);
nor UO_642 (O_642,N_13315,N_14668);
nand UO_643 (O_643,N_12679,N_13782);
nor UO_644 (O_644,N_12954,N_12139);
or UO_645 (O_645,N_14698,N_12209);
nand UO_646 (O_646,N_14726,N_12353);
or UO_647 (O_647,N_14657,N_14903);
or UO_648 (O_648,N_14897,N_12809);
nand UO_649 (O_649,N_12559,N_12189);
nor UO_650 (O_650,N_12004,N_12017);
nand UO_651 (O_651,N_13809,N_14504);
nand UO_652 (O_652,N_13618,N_13976);
nor UO_653 (O_653,N_12213,N_14166);
or UO_654 (O_654,N_12295,N_14870);
nor UO_655 (O_655,N_14945,N_13520);
nand UO_656 (O_656,N_13673,N_12267);
nand UO_657 (O_657,N_13325,N_14914);
or UO_658 (O_658,N_14911,N_14179);
nor UO_659 (O_659,N_12155,N_14065);
nand UO_660 (O_660,N_13990,N_12676);
nand UO_661 (O_661,N_13918,N_14275);
or UO_662 (O_662,N_12046,N_12278);
or UO_663 (O_663,N_12607,N_14280);
or UO_664 (O_664,N_13550,N_12703);
and UO_665 (O_665,N_14112,N_14152);
nor UO_666 (O_666,N_14436,N_14029);
nand UO_667 (O_667,N_12290,N_12103);
and UO_668 (O_668,N_13585,N_13165);
or UO_669 (O_669,N_14467,N_14652);
or UO_670 (O_670,N_13334,N_13256);
xor UO_671 (O_671,N_14067,N_14141);
and UO_672 (O_672,N_12568,N_13209);
or UO_673 (O_673,N_13264,N_12261);
nand UO_674 (O_674,N_14230,N_12479);
nor UO_675 (O_675,N_12638,N_12364);
or UO_676 (O_676,N_14930,N_14607);
nor UO_677 (O_677,N_12579,N_12868);
nand UO_678 (O_678,N_14281,N_14402);
nor UO_679 (O_679,N_13407,N_13063);
or UO_680 (O_680,N_12041,N_13049);
nand UO_681 (O_681,N_14428,N_14422);
or UO_682 (O_682,N_13276,N_14978);
and UO_683 (O_683,N_12067,N_12346);
nor UO_684 (O_684,N_14224,N_13893);
nor UO_685 (O_685,N_13392,N_12560);
or UO_686 (O_686,N_12116,N_14824);
and UO_687 (O_687,N_12250,N_12658);
nor UO_688 (O_688,N_13700,N_14299);
and UO_689 (O_689,N_14489,N_12039);
nand UO_690 (O_690,N_12735,N_12281);
nor UO_691 (O_691,N_13979,N_12902);
nand UO_692 (O_692,N_14054,N_13257);
nor UO_693 (O_693,N_13278,N_12036);
nand UO_694 (O_694,N_14441,N_14265);
and UO_695 (O_695,N_13221,N_12673);
or UO_696 (O_696,N_14612,N_14792);
or UO_697 (O_697,N_12768,N_14975);
nor UO_698 (O_698,N_13444,N_14506);
nor UO_699 (O_699,N_14782,N_12726);
or UO_700 (O_700,N_14124,N_13680);
nor UO_701 (O_701,N_12897,N_14913);
or UO_702 (O_702,N_14185,N_12564);
nand UO_703 (O_703,N_14123,N_13055);
or UO_704 (O_704,N_12526,N_14959);
nor UO_705 (O_705,N_14034,N_14905);
and UO_706 (O_706,N_12503,N_12548);
xnor UO_707 (O_707,N_13650,N_12320);
nor UO_708 (O_708,N_12848,N_13896);
nand UO_709 (O_709,N_13805,N_12727);
or UO_710 (O_710,N_12943,N_14853);
and UO_711 (O_711,N_13733,N_12463);
nor UO_712 (O_712,N_14851,N_13717);
or UO_713 (O_713,N_14380,N_13915);
or UO_714 (O_714,N_14320,N_12381);
nand UO_715 (O_715,N_13679,N_13412);
nand UO_716 (O_716,N_12109,N_14819);
nor UO_717 (O_717,N_12780,N_12776);
nor UO_718 (O_718,N_12454,N_13563);
nor UO_719 (O_719,N_14555,N_12273);
nor UO_720 (O_720,N_12138,N_12460);
nor UO_721 (O_721,N_12132,N_14001);
nor UO_722 (O_722,N_13802,N_12407);
nand UO_723 (O_723,N_12207,N_12698);
xnor UO_724 (O_724,N_13949,N_12682);
nor UO_725 (O_725,N_13825,N_12368);
or UO_726 (O_726,N_14773,N_12414);
xor UO_727 (O_727,N_12448,N_13823);
or UO_728 (O_728,N_14021,N_13343);
xor UO_729 (O_729,N_12009,N_14998);
nor UO_730 (O_730,N_12191,N_14297);
or UO_731 (O_731,N_13559,N_13417);
or UO_732 (O_732,N_13832,N_12243);
nor UO_733 (O_733,N_12953,N_13466);
or UO_734 (O_734,N_13907,N_14369);
nand UO_735 (O_735,N_13145,N_12367);
and UO_736 (O_736,N_14760,N_13182);
xor UO_737 (O_737,N_12204,N_13162);
nand UO_738 (O_738,N_13268,N_12898);
nor UO_739 (O_739,N_14811,N_12581);
nand UO_740 (O_740,N_13301,N_13414);
xor UO_741 (O_741,N_13329,N_13195);
nor UO_742 (O_742,N_12688,N_13167);
or UO_743 (O_743,N_13113,N_14232);
or UO_744 (O_744,N_12648,N_14639);
or UO_745 (O_745,N_14051,N_12933);
nand UO_746 (O_746,N_12881,N_13897);
nor UO_747 (O_747,N_14769,N_13286);
and UO_748 (O_748,N_12379,N_13820);
and UO_749 (O_749,N_12714,N_13509);
nand UO_750 (O_750,N_14908,N_13765);
and UO_751 (O_751,N_14585,N_14162);
nor UO_752 (O_752,N_13168,N_13686);
nand UO_753 (O_753,N_12939,N_13822);
nand UO_754 (O_754,N_13797,N_14557);
and UO_755 (O_755,N_13177,N_14481);
nand UO_756 (O_756,N_14193,N_12771);
nand UO_757 (O_757,N_14160,N_13420);
nand UO_758 (O_758,N_14227,N_14216);
and UO_759 (O_759,N_14258,N_13939);
or UO_760 (O_760,N_13657,N_12321);
nand UO_761 (O_761,N_13307,N_13440);
or UO_762 (O_762,N_13240,N_12543);
nand UO_763 (O_763,N_14776,N_13013);
or UO_764 (O_764,N_14263,N_12973);
or UO_765 (O_765,N_14539,N_13622);
nand UO_766 (O_766,N_12504,N_13889);
nand UO_767 (O_767,N_14562,N_13541);
xor UO_768 (O_768,N_12813,N_13333);
or UO_769 (O_769,N_12621,N_13462);
or UO_770 (O_770,N_12000,N_13988);
nand UO_771 (O_771,N_12185,N_14629);
xor UO_772 (O_772,N_14800,N_14904);
nor UO_773 (O_773,N_14316,N_12508);
xor UO_774 (O_774,N_12555,N_14611);
or UO_775 (O_775,N_12302,N_12865);
or UO_776 (O_776,N_14317,N_14448);
nor UO_777 (O_777,N_13275,N_13355);
xnor UO_778 (O_778,N_14373,N_14526);
nor UO_779 (O_779,N_14472,N_13265);
nor UO_780 (O_780,N_13401,N_12326);
xor UO_781 (O_781,N_13387,N_14869);
nor UO_782 (O_782,N_12664,N_13999);
or UO_783 (O_783,N_12077,N_14192);
or UO_784 (O_784,N_12102,N_14108);
nor UO_785 (O_785,N_13404,N_14331);
nand UO_786 (O_786,N_12520,N_12910);
nor UO_787 (O_787,N_12777,N_14551);
or UO_788 (O_788,N_14857,N_14784);
nor UO_789 (O_789,N_14161,N_12770);
nor UO_790 (O_790,N_13225,N_13723);
or UO_791 (O_791,N_14762,N_13608);
nand UO_792 (O_792,N_14231,N_13943);
nor UO_793 (O_793,N_13306,N_14130);
and UO_794 (O_794,N_14061,N_14865);
and UO_795 (O_795,N_12649,N_14432);
or UO_796 (O_796,N_13377,N_14589);
xor UO_797 (O_797,N_13033,N_12226);
and UO_798 (O_798,N_13080,N_14025);
nor UO_799 (O_799,N_13202,N_14642);
nand UO_800 (O_800,N_14378,N_14002);
and UO_801 (O_801,N_13384,N_14418);
and UO_802 (O_802,N_13845,N_13946);
nand UO_803 (O_803,N_13163,N_13042);
and UO_804 (O_804,N_14311,N_13291);
nand UO_805 (O_805,N_14376,N_13701);
or UO_806 (O_806,N_12057,N_14779);
nor UO_807 (O_807,N_13969,N_14211);
xnor UO_808 (O_808,N_13505,N_14101);
nand UO_809 (O_809,N_14758,N_13312);
nand UO_810 (O_810,N_14957,N_13000);
nor UO_811 (O_811,N_12995,N_12808);
or UO_812 (O_812,N_13570,N_12183);
or UO_813 (O_813,N_12882,N_12372);
and UO_814 (O_814,N_14040,N_13521);
and UO_815 (O_815,N_13214,N_12142);
nand UO_816 (O_816,N_13190,N_13925);
nor UO_817 (O_817,N_12499,N_14841);
nand UO_818 (O_818,N_13834,N_13295);
xnor UO_819 (O_819,N_13088,N_12021);
and UO_820 (O_820,N_14644,N_12801);
nand UO_821 (O_821,N_13100,N_14204);
or UO_822 (O_822,N_14735,N_14172);
nor UO_823 (O_823,N_12168,N_12670);
nor UO_824 (O_824,N_13647,N_14264);
nor UO_825 (O_825,N_14053,N_12343);
or UO_826 (O_826,N_13263,N_14273);
nand UO_827 (O_827,N_14419,N_14679);
and UO_828 (O_828,N_13525,N_13489);
nor UO_829 (O_829,N_14617,N_12374);
nand UO_830 (O_830,N_13742,N_14327);
nor UO_831 (O_831,N_14106,N_12572);
and UO_832 (O_832,N_12007,N_14649);
nor UO_833 (O_833,N_13317,N_13908);
or UO_834 (O_834,N_12242,N_13421);
or UO_835 (O_835,N_12156,N_13516);
nand UO_836 (O_836,N_13273,N_12160);
xnor UO_837 (O_837,N_14837,N_14719);
and UO_838 (O_838,N_12836,N_14696);
nor UO_839 (O_839,N_14790,N_13357);
nand UO_840 (O_840,N_14277,N_13965);
nor UO_841 (O_841,N_12137,N_13719);
nor UO_842 (O_842,N_14511,N_14920);
nor UO_843 (O_843,N_14931,N_13704);
nor UO_844 (O_844,N_14684,N_14655);
nand UO_845 (O_845,N_13967,N_14494);
nor UO_846 (O_846,N_12175,N_14803);
or UO_847 (O_847,N_13863,N_14906);
nand UO_848 (O_848,N_14298,N_14536);
or UO_849 (O_849,N_14396,N_12383);
nor UO_850 (O_850,N_13841,N_13069);
or UO_851 (O_851,N_14861,N_14743);
nor UO_852 (O_852,N_14768,N_14505);
xnor UO_853 (O_853,N_12592,N_14016);
xor UO_854 (O_854,N_14410,N_14734);
and UO_855 (O_855,N_12804,N_12553);
nor UO_856 (O_856,N_14451,N_13469);
nor UO_857 (O_857,N_14343,N_14541);
xnor UO_858 (O_858,N_12604,N_13010);
or UO_859 (O_859,N_14220,N_14537);
nor UO_860 (O_860,N_14958,N_12791);
nor UO_861 (O_861,N_14748,N_14295);
nand UO_862 (O_862,N_13308,N_13894);
or UO_863 (O_863,N_12918,N_12537);
nor UO_864 (O_864,N_14153,N_12341);
nand UO_865 (O_865,N_12947,N_14064);
or UO_866 (O_866,N_12128,N_14799);
nand UO_867 (O_867,N_12976,N_14454);
and UO_868 (O_868,N_13075,N_12443);
nor UO_869 (O_869,N_14066,N_12958);
nor UO_870 (O_870,N_12843,N_13025);
and UO_871 (O_871,N_14592,N_13020);
nand UO_872 (O_872,N_12558,N_14513);
and UO_873 (O_873,N_14431,N_13829);
nor UO_874 (O_874,N_12292,N_14685);
nor UO_875 (O_875,N_13040,N_13601);
and UO_876 (O_876,N_14182,N_14794);
nand UO_877 (O_877,N_12489,N_13226);
and UO_878 (O_878,N_13016,N_12846);
xnor UO_879 (O_879,N_14084,N_13786);
or UO_880 (O_880,N_14151,N_12297);
nand UO_881 (O_881,N_13676,N_13199);
and UO_882 (O_882,N_13477,N_13944);
and UO_883 (O_883,N_12487,N_14174);
nand UO_884 (O_884,N_14896,N_12884);
and UO_885 (O_885,N_14019,N_12911);
and UO_886 (O_886,N_13883,N_13699);
and UO_887 (O_887,N_14050,N_12721);
nand UO_888 (O_888,N_13672,N_13260);
xnor UO_889 (O_889,N_14876,N_13110);
nand UO_890 (O_890,N_14452,N_13455);
or UO_891 (O_891,N_14091,N_12965);
nand UO_892 (O_892,N_14955,N_13904);
and UO_893 (O_893,N_14813,N_13787);
and UO_894 (O_894,N_14414,N_14352);
or UO_895 (O_895,N_14294,N_13798);
nor UO_896 (O_896,N_13728,N_12919);
nor UO_897 (O_897,N_13015,N_13961);
nand UO_898 (O_898,N_13458,N_13909);
nand UO_899 (O_899,N_13888,N_14415);
or UO_900 (O_900,N_13399,N_12634);
and UO_901 (O_901,N_13367,N_13037);
nand UO_902 (O_902,N_13538,N_14672);
nor UO_903 (O_903,N_13856,N_12626);
xnor UO_904 (O_904,N_14764,N_14884);
or UO_905 (O_905,N_14695,N_12143);
or UO_906 (O_906,N_13021,N_12775);
or UO_907 (O_907,N_13600,N_14163);
nor UO_908 (O_908,N_12023,N_13586);
and UO_909 (O_909,N_12671,N_13948);
nand UO_910 (O_910,N_14140,N_14530);
xnor UO_911 (O_911,N_14816,N_13767);
nor UO_912 (O_912,N_12337,N_12117);
or UO_913 (O_913,N_12669,N_12681);
or UO_914 (O_914,N_13697,N_12241);
nor UO_915 (O_915,N_14942,N_14989);
and UO_916 (O_916,N_14646,N_14276);
nor UO_917 (O_917,N_12141,N_14403);
and UO_918 (O_918,N_14308,N_12483);
nand UO_919 (O_919,N_12352,N_12205);
nor UO_920 (O_920,N_12981,N_13857);
nand UO_921 (O_921,N_13480,N_12304);
and UO_922 (O_922,N_13828,N_14891);
or UO_923 (O_923,N_13398,N_13712);
nand UO_924 (O_924,N_12439,N_12705);
nor UO_925 (O_925,N_13836,N_14973);
and UO_926 (O_926,N_12704,N_14885);
or UO_927 (O_927,N_13400,N_12361);
or UO_928 (O_928,N_14103,N_12200);
nor UO_929 (O_929,N_12955,N_12229);
nand UO_930 (O_930,N_14863,N_13374);
nor UO_931 (O_931,N_13611,N_12180);
nand UO_932 (O_932,N_14259,N_12366);
nand UO_933 (O_933,N_14781,N_14708);
nor UO_934 (O_934,N_12618,N_12569);
or UO_935 (O_935,N_12497,N_12608);
or UO_936 (O_936,N_13602,N_14804);
nor UO_937 (O_937,N_12601,N_13373);
and UO_938 (O_938,N_14687,N_14714);
or UO_939 (O_939,N_12538,N_14272);
and UO_940 (O_940,N_13708,N_12870);
or UO_941 (O_941,N_14286,N_14889);
nand UO_942 (O_942,N_13614,N_14385);
or UO_943 (O_943,N_12872,N_12339);
nand UO_944 (O_944,N_13917,N_12677);
nand UO_945 (O_945,N_14798,N_14267);
or UO_946 (O_946,N_14968,N_12500);
and UO_947 (O_947,N_12270,N_14070);
and UO_948 (O_948,N_14621,N_13995);
and UO_949 (O_949,N_13078,N_14351);
nor UO_950 (O_950,N_14552,N_12655);
nor UO_951 (O_951,N_12830,N_13488);
or UO_952 (O_952,N_14190,N_12741);
and UO_953 (O_953,N_12680,N_14296);
xor UO_954 (O_954,N_14301,N_14599);
nor UO_955 (O_955,N_12135,N_13327);
nor UO_956 (O_956,N_14389,N_14072);
nand UO_957 (O_957,N_12406,N_14339);
nor UO_958 (O_958,N_12176,N_14689);
nor UO_959 (O_959,N_14572,N_13821);
nand UO_960 (O_960,N_13229,N_13690);
nor UO_961 (O_961,N_13448,N_13773);
or UO_962 (O_962,N_14090,N_14757);
nand UO_963 (O_963,N_12683,N_14085);
nand UO_964 (O_964,N_14471,N_13572);
nand UO_965 (O_965,N_14676,N_12028);
nor UO_966 (O_966,N_13471,N_14893);
nand UO_967 (O_967,N_14690,N_13432);
or UO_968 (O_968,N_13770,N_13428);
nand UO_969 (O_969,N_14202,N_12079);
and UO_970 (O_970,N_14485,N_13628);
xnor UO_971 (O_971,N_13788,N_13427);
and UO_972 (O_972,N_14705,N_12173);
nor UO_973 (O_973,N_12773,N_12382);
nand UO_974 (O_974,N_14563,N_13727);
or UO_975 (O_975,N_13975,N_14713);
or UO_976 (O_976,N_13491,N_13766);
and UO_977 (O_977,N_13743,N_12986);
and UO_978 (O_978,N_13714,N_12431);
and UO_979 (O_979,N_12377,N_13666);
and UO_980 (O_980,N_12149,N_12752);
nand UO_981 (O_981,N_14391,N_12535);
nand UO_982 (O_982,N_14964,N_12728);
or UO_983 (O_983,N_14970,N_13230);
nor UO_984 (O_984,N_13436,N_13379);
nor UO_985 (O_985,N_12794,N_12873);
nand UO_986 (O_986,N_13138,N_12146);
or UO_987 (O_987,N_12059,N_12826);
xnor UO_988 (O_988,N_14347,N_13824);
or UO_989 (O_989,N_14771,N_13160);
or UO_990 (O_990,N_14701,N_12915);
and UO_991 (O_991,N_12576,N_14963);
or UO_992 (O_992,N_13337,N_12795);
nor UO_993 (O_993,N_13101,N_14724);
nor UO_994 (O_994,N_13060,N_12660);
or UO_995 (O_995,N_12861,N_12220);
nand UO_996 (O_996,N_13754,N_14720);
xor UO_997 (O_997,N_12476,N_14558);
or UO_998 (O_998,N_13349,N_13783);
or UO_999 (O_999,N_12119,N_13116);
nand UO_1000 (O_1000,N_12114,N_14497);
nor UO_1001 (O_1001,N_13870,N_14895);
and UO_1002 (O_1002,N_14052,N_14470);
nor UO_1003 (O_1003,N_12468,N_13804);
nor UO_1004 (O_1004,N_13253,N_12360);
nand UO_1005 (O_1005,N_12736,N_12819);
and UO_1006 (O_1006,N_14991,N_12111);
and UO_1007 (O_1007,N_14845,N_14898);
nand UO_1008 (O_1008,N_14739,N_12969);
nand UO_1009 (O_1009,N_13041,N_14099);
xnor UO_1010 (O_1010,N_14499,N_14126);
nor UO_1011 (O_1011,N_14098,N_13640);
nor UO_1012 (O_1012,N_14219,N_12871);
and UO_1013 (O_1013,N_12951,N_14203);
nand UO_1014 (O_1014,N_14915,N_13071);
or UO_1015 (O_1015,N_13038,N_13359);
xnor UO_1016 (O_1016,N_12711,N_14271);
and UO_1017 (O_1017,N_12154,N_12247);
and UO_1018 (O_1018,N_13878,N_12196);
nor UO_1019 (O_1019,N_12384,N_12070);
nand UO_1020 (O_1020,N_13986,N_12210);
and UO_1021 (O_1021,N_13612,N_14310);
and UO_1022 (O_1022,N_14767,N_14829);
and UO_1023 (O_1023,N_12315,N_12927);
nor UO_1024 (O_1024,N_14605,N_14114);
nor UO_1025 (O_1025,N_12349,N_14173);
and UO_1026 (O_1026,N_12221,N_13267);
nor UO_1027 (O_1027,N_14729,N_14434);
nor UO_1028 (O_1028,N_14814,N_12158);
nor UO_1029 (O_1029,N_12533,N_12112);
or UO_1030 (O_1030,N_14269,N_14370);
nand UO_1031 (O_1031,N_14856,N_12370);
nand UO_1032 (O_1032,N_14363,N_12557);
or UO_1033 (O_1033,N_12314,N_12551);
xor UO_1034 (O_1034,N_13321,N_12492);
or UO_1035 (O_1035,N_14392,N_12970);
nor UO_1036 (O_1036,N_13282,N_12020);
nand UO_1037 (O_1037,N_14110,N_14860);
nand UO_1038 (O_1038,N_13763,N_12330);
and UO_1039 (O_1039,N_14088,N_13196);
nand UO_1040 (O_1040,N_13780,N_12042);
or UO_1041 (O_1041,N_12967,N_12254);
or UO_1042 (O_1042,N_14864,N_13124);
or UO_1043 (O_1043,N_12968,N_12975);
or UO_1044 (O_1044,N_14274,N_13389);
nand UO_1045 (O_1045,N_12334,N_13811);
nor UO_1046 (O_1046,N_14907,N_14459);
or UO_1047 (O_1047,N_14077,N_13737);
xor UO_1048 (O_1048,N_12272,N_13599);
and UO_1049 (O_1049,N_14238,N_14226);
nor UO_1050 (O_1050,N_12888,N_12570);
and UO_1051 (O_1051,N_12251,N_12194);
or UO_1052 (O_1052,N_13390,N_13696);
nand UO_1053 (O_1053,N_12545,N_12258);
or UO_1054 (O_1054,N_13011,N_14969);
or UO_1055 (O_1055,N_12805,N_12074);
nand UO_1056 (O_1056,N_13234,N_14946);
nor UO_1057 (O_1057,N_12903,N_12389);
nor UO_1058 (O_1058,N_12363,N_14406);
nand UO_1059 (O_1059,N_13109,N_13807);
and UO_1060 (O_1060,N_14252,N_12574);
and UO_1061 (O_1061,N_14491,N_12166);
or UO_1062 (O_1062,N_12833,N_12063);
nand UO_1063 (O_1063,N_13254,N_13358);
nand UO_1064 (O_1064,N_13815,N_13886);
and UO_1065 (O_1065,N_14538,N_14078);
and UO_1066 (O_1066,N_13280,N_12708);
nand UO_1067 (O_1067,N_12510,N_12900);
nor UO_1068 (O_1068,N_14579,N_12424);
or UO_1069 (O_1069,N_12262,N_14894);
and UO_1070 (O_1070,N_14079,N_14498);
and UO_1071 (O_1071,N_12073,N_14278);
nand UO_1072 (O_1072,N_12170,N_13395);
nand UO_1073 (O_1073,N_13873,N_14627);
nor UO_1074 (O_1074,N_13095,N_13416);
or UO_1075 (O_1075,N_13220,N_12619);
and UO_1076 (O_1076,N_12860,N_14306);
xnor UO_1077 (O_1077,N_12026,N_12347);
nand UO_1078 (O_1078,N_14520,N_14809);
and UO_1079 (O_1079,N_14953,N_12404);
nor UO_1080 (O_1080,N_12082,N_13865);
nor UO_1081 (O_1081,N_14993,N_12921);
nand UO_1082 (O_1082,N_12470,N_14006);
or UO_1083 (O_1083,N_13187,N_13459);
or UO_1084 (O_1084,N_13500,N_14669);
nand UO_1085 (O_1085,N_13761,N_14313);
xnor UO_1086 (O_1086,N_14250,N_14113);
nand UO_1087 (O_1087,N_12850,N_12605);
and UO_1088 (O_1088,N_14601,N_12403);
nor UO_1089 (O_1089,N_14584,N_12862);
or UO_1090 (O_1090,N_14131,N_12118);
or UO_1091 (O_1091,N_14283,N_14212);
and UO_1092 (O_1092,N_12307,N_12690);
or UO_1093 (O_1093,N_13391,N_12216);
nor UO_1094 (O_1094,N_14756,N_13687);
nor UO_1095 (O_1095,N_12122,N_12912);
or UO_1096 (O_1096,N_14554,N_12511);
nor UO_1097 (O_1097,N_13035,N_12027);
and UO_1098 (O_1098,N_13014,N_14096);
nor UO_1099 (O_1099,N_13882,N_12591);
or UO_1100 (O_1100,N_12427,N_13383);
and UO_1101 (O_1101,N_13446,N_12583);
nand UO_1102 (O_1102,N_13003,N_13819);
or UO_1103 (O_1103,N_14187,N_13335);
nand UO_1104 (O_1104,N_14046,N_14780);
nor UO_1105 (O_1105,N_14209,N_12636);
and UO_1106 (O_1106,N_14120,N_14142);
nand UO_1107 (O_1107,N_13443,N_14105);
and UO_1108 (O_1108,N_12395,N_13241);
nand UO_1109 (O_1109,N_14626,N_14011);
and UO_1110 (O_1110,N_13336,N_13667);
xor UO_1111 (O_1111,N_14197,N_12399);
nand UO_1112 (O_1112,N_12949,N_13250);
and UO_1113 (O_1113,N_14960,N_12916);
and UO_1114 (O_1114,N_12507,N_14725);
nand UO_1115 (O_1115,N_13288,N_13537);
or UO_1116 (O_1116,N_13099,N_13974);
nor UO_1117 (O_1117,N_13901,N_14632);
nor UO_1118 (O_1118,N_12397,N_14755);
or UO_1119 (O_1119,N_14512,N_13193);
nor UO_1120 (O_1120,N_13945,N_13328);
and UO_1121 (O_1121,N_13669,N_12654);
nor UO_1122 (O_1122,N_13236,N_12786);
or UO_1123 (O_1123,N_13626,N_13198);
or UO_1124 (O_1124,N_14934,N_12313);
nand UO_1125 (O_1125,N_14122,N_13445);
and UO_1126 (O_1126,N_12817,N_13452);
and UO_1127 (O_1127,N_12631,N_12316);
nor UO_1128 (O_1128,N_12089,N_13565);
xor UO_1129 (O_1129,N_12037,N_13753);
nor UO_1130 (O_1130,N_13514,N_14045);
nor UO_1131 (O_1131,N_12469,N_14614);
or UO_1132 (O_1132,N_14445,N_13558);
nand UO_1133 (O_1133,N_14925,N_12099);
or UO_1134 (O_1134,N_14686,N_13450);
nor UO_1135 (O_1135,N_14683,N_12371);
nand UO_1136 (O_1136,N_12524,N_13029);
and UO_1137 (O_1137,N_13362,N_14659);
or UO_1138 (O_1138,N_14314,N_12351);
nor UO_1139 (O_1139,N_13905,N_13108);
nand UO_1140 (O_1140,N_13005,N_12637);
or UO_1141 (O_1141,N_12096,N_14818);
nor UO_1142 (O_1142,N_12806,N_12928);
nand UO_1143 (O_1143,N_13621,N_13057);
xnor UO_1144 (O_1144,N_12957,N_14604);
or UO_1145 (O_1145,N_13963,N_13898);
xor UO_1146 (O_1146,N_14521,N_13074);
and UO_1147 (O_1147,N_13940,N_13136);
nand UO_1148 (O_1148,N_13197,N_12577);
or UO_1149 (O_1149,N_14453,N_12932);
or UO_1150 (O_1150,N_14651,N_14456);
nand UO_1151 (O_1151,N_12092,N_14292);
or UO_1152 (O_1152,N_13781,N_12259);
nor UO_1153 (O_1153,N_12255,N_12136);
xnor UO_1154 (O_1154,N_12540,N_12854);
or UO_1155 (O_1155,N_14288,N_14888);
xor UO_1156 (O_1156,N_12218,N_13463);
nor UO_1157 (O_1157,N_14984,N_14524);
and UO_1158 (O_1158,N_12734,N_12783);
nand UO_1159 (O_1159,N_14075,N_13243);
nor UO_1160 (O_1160,N_12224,N_14097);
or UO_1161 (O_1161,N_13394,N_13735);
and UO_1162 (O_1162,N_14095,N_12696);
xor UO_1163 (O_1163,N_12426,N_13044);
nand UO_1164 (O_1164,N_13248,N_13512);
or UO_1165 (O_1165,N_12934,N_14972);
nand UO_1166 (O_1166,N_13526,N_13211);
and UO_1167 (O_1167,N_13535,N_12214);
and UO_1168 (O_1168,N_14474,N_13921);
nand UO_1169 (O_1169,N_14457,N_13297);
nor UO_1170 (O_1170,N_13174,N_13039);
xnor UO_1171 (O_1171,N_13228,N_14715);
and UO_1172 (O_1172,N_14648,N_14409);
nor UO_1173 (O_1173,N_13302,N_14951);
and UO_1174 (O_1174,N_12271,N_13410);
or UO_1175 (O_1175,N_14117,N_13659);
and UO_1176 (O_1176,N_13259,N_14825);
nand UO_1177 (O_1177,N_13431,N_13279);
xnor UO_1178 (O_1178,N_13912,N_14531);
xnor UO_1179 (O_1179,N_13530,N_12051);
or UO_1180 (O_1180,N_14940,N_14832);
xnor UO_1181 (O_1181,N_14464,N_13114);
nand UO_1182 (O_1182,N_14028,N_14248);
nand UO_1183 (O_1183,N_14315,N_14625);
and UO_1184 (O_1184,N_13957,N_13619);
and UO_1185 (O_1185,N_13105,N_12148);
or UO_1186 (O_1186,N_13756,N_13793);
and UO_1187 (O_1187,N_12113,N_12441);
or UO_1188 (O_1188,N_13119,N_12589);
nor UO_1189 (O_1189,N_14121,N_12415);
nor UO_1190 (O_1190,N_14024,N_12129);
and UO_1191 (O_1191,N_14394,N_13838);
nand UO_1192 (O_1192,N_13251,N_12702);
xnor UO_1193 (O_1193,N_13937,N_13092);
nand UO_1194 (O_1194,N_13345,N_13172);
nor UO_1195 (O_1195,N_13775,N_14850);
nor UO_1196 (O_1196,N_12480,N_13224);
nand UO_1197 (O_1197,N_12869,N_12369);
or UO_1198 (O_1198,N_12661,N_13574);
or UO_1199 (O_1199,N_14158,N_14988);
nor UO_1200 (O_1200,N_12582,N_14847);
or UO_1201 (O_1201,N_13294,N_14545);
nor UO_1202 (O_1202,N_13926,N_14039);
xnor UO_1203 (O_1203,N_13370,N_14439);
or UO_1204 (O_1204,N_13645,N_13072);
nand UO_1205 (O_1205,N_12106,N_14667);
nor UO_1206 (O_1206,N_14200,N_12342);
and UO_1207 (O_1207,N_12310,N_13938);
nor UO_1208 (O_1208,N_13784,N_14345);
and UO_1209 (O_1209,N_12450,N_13175);
or UO_1210 (O_1210,N_12380,N_14157);
or UO_1211 (O_1211,N_12445,N_12248);
or UO_1212 (O_1212,N_13233,N_12886);
nand UO_1213 (O_1213,N_12722,N_14336);
nor UO_1214 (O_1214,N_12996,N_12731);
nor UO_1215 (O_1215,N_12513,N_14935);
or UO_1216 (O_1216,N_12765,N_13903);
or UO_1217 (O_1217,N_12814,N_13022);
nand UO_1218 (O_1218,N_12182,N_12877);
xor UO_1219 (O_1219,N_13161,N_13564);
or UO_1220 (O_1220,N_13546,N_12174);
nand UO_1221 (O_1221,N_12212,N_13997);
or UO_1222 (O_1222,N_12049,N_13576);
or UO_1223 (O_1223,N_14234,N_13959);
and UO_1224 (O_1224,N_14775,N_12782);
nand UO_1225 (O_1225,N_12325,N_13192);
nor UO_1226 (O_1226,N_12385,N_14304);
nor UO_1227 (O_1227,N_12348,N_14430);
nand UO_1228 (O_1228,N_13036,N_13660);
nand UO_1229 (O_1229,N_13664,N_14677);
and UO_1230 (O_1230,N_13237,N_12167);
and UO_1231 (O_1231,N_13104,N_14022);
nand UO_1232 (O_1232,N_14670,N_13403);
and UO_1233 (O_1233,N_12880,N_13978);
or UO_1234 (O_1234,N_12978,N_14421);
nor UO_1235 (O_1235,N_12666,N_12956);
or UO_1236 (O_1236,N_14210,N_13507);
nand UO_1237 (O_1237,N_14692,N_14037);
nor UO_1238 (O_1238,N_13577,N_13117);
or UO_1239 (O_1239,N_12301,N_13958);
nand UO_1240 (O_1240,N_13076,N_13456);
or UO_1241 (O_1241,N_14587,N_13352);
nand UO_1242 (O_1242,N_12597,N_12926);
or UO_1243 (O_1243,N_13552,N_12562);
nand UO_1244 (O_1244,N_12446,N_14165);
and UO_1245 (O_1245,N_14923,N_12266);
xnor UO_1246 (O_1246,N_12473,N_14386);
nand UO_1247 (O_1247,N_13692,N_14184);
or UO_1248 (O_1248,N_12005,N_13584);
or UO_1249 (O_1249,N_14731,N_14462);
and UO_1250 (O_1250,N_12451,N_13353);
nor UO_1251 (O_1251,N_14080,N_13981);
or UO_1252 (O_1252,N_14159,N_14577);
xnor UO_1253 (O_1253,N_13547,N_12908);
xor UO_1254 (O_1254,N_14565,N_12823);
nor UO_1255 (O_1255,N_12420,N_13884);
and UO_1256 (O_1256,N_12333,N_13309);
and UO_1257 (O_1257,N_14688,N_12529);
and UO_1258 (O_1258,N_12952,N_14460);
and UO_1259 (O_1259,N_12824,N_13923);
and UO_1260 (O_1260,N_12344,N_12481);
or UO_1261 (O_1261,N_13962,N_13847);
and UO_1262 (O_1262,N_13722,N_12085);
nand UO_1263 (O_1263,N_12104,N_13853);
nand UO_1264 (O_1264,N_14529,N_13850);
and UO_1265 (O_1265,N_12296,N_12120);
nand UO_1266 (O_1266,N_13661,N_12394);
and UO_1267 (O_1267,N_14835,N_14620);
nand UO_1268 (O_1268,N_12100,N_12044);
and UO_1269 (O_1269,N_14517,N_14586);
nand UO_1270 (O_1270,N_13434,N_14999);
or UO_1271 (O_1271,N_12856,N_12633);
or UO_1272 (O_1272,N_13644,N_14229);
nor UO_1273 (O_1273,N_13149,N_12206);
and UO_1274 (O_1274,N_13615,N_14390);
and UO_1275 (O_1275,N_13425,N_14477);
or UO_1276 (O_1276,N_12078,N_14249);
xnor UO_1277 (O_1277,N_13663,N_13891);
and UO_1278 (O_1278,N_12197,N_14330);
nor UO_1279 (O_1279,N_12839,N_14831);
nor UO_1280 (O_1280,N_13474,N_14606);
and UO_1281 (O_1281,N_14650,N_13703);
xnor UO_1282 (O_1282,N_14475,N_12588);
nor UO_1283 (O_1283,N_14518,N_14624);
or UO_1284 (O_1284,N_13806,N_14647);
or UO_1285 (O_1285,N_13258,N_13137);
xor UO_1286 (O_1286,N_12434,N_14654);
xnor UO_1287 (O_1287,N_13519,N_12288);
and UO_1288 (O_1288,N_14350,N_14622);
and UO_1289 (O_1289,N_13709,N_12800);
nor UO_1290 (O_1290,N_13324,N_13498);
nor UO_1291 (O_1291,N_13262,N_12994);
and UO_1292 (O_1292,N_13244,N_13913);
nand UO_1293 (O_1293,N_13235,N_12963);
and UO_1294 (O_1294,N_14133,N_12338);
and UO_1295 (O_1295,N_14488,N_14030);
xor UO_1296 (O_1296,N_14221,N_14509);
nand UO_1297 (O_1297,N_13024,N_12547);
and UO_1298 (O_1298,N_14877,N_13341);
nand UO_1299 (O_1299,N_13655,N_14732);
nor UO_1300 (O_1300,N_13155,N_14630);
xnor UO_1301 (O_1301,N_14005,N_12700);
or UO_1302 (O_1302,N_13862,N_12534);
nor UO_1303 (O_1303,N_12340,N_13183);
nor UO_1304 (O_1304,N_13771,N_12904);
xor UO_1305 (O_1305,N_12147,N_14083);
or UO_1306 (O_1306,N_12054,N_13143);
and UO_1307 (O_1307,N_13592,N_12401);
xnor UO_1308 (O_1308,N_14284,N_14450);
and UO_1309 (O_1309,N_14071,N_14170);
xor UO_1310 (O_1310,N_14880,N_14109);
or UO_1311 (O_1311,N_14044,N_12747);
nor UO_1312 (O_1312,N_13652,N_12265);
nor UO_1313 (O_1313,N_12525,N_12421);
xnor UO_1314 (O_1314,N_12066,N_14321);
and UO_1315 (O_1315,N_12687,N_12668);
or UO_1316 (O_1316,N_14437,N_13131);
nor UO_1317 (O_1317,N_13473,N_12006);
nand UO_1318 (O_1318,N_13365,N_14591);
or UO_1319 (O_1319,N_14137,N_14004);
nor UO_1320 (O_1320,N_13097,N_14673);
nand UO_1321 (O_1321,N_14357,N_14772);
nor UO_1322 (O_1322,N_13992,N_12058);
nand UO_1323 (O_1323,N_14763,N_12289);
xnor UO_1324 (O_1324,N_14691,N_12215);
or UO_1325 (O_1325,N_13026,N_14063);
and UO_1326 (O_1326,N_13289,N_14424);
or UO_1327 (O_1327,N_13627,N_12639);
xnor UO_1328 (O_1328,N_12276,N_12482);
nand UO_1329 (O_1329,N_14933,N_14251);
or UO_1330 (O_1330,N_14549,N_14041);
nor UO_1331 (O_1331,N_12293,N_12845);
nand UO_1332 (O_1332,N_13429,N_14962);
nor UO_1333 (O_1333,N_13543,N_13772);
or UO_1334 (O_1334,N_12181,N_12345);
nor UO_1335 (O_1335,N_13115,N_12550);
or UO_1336 (O_1336,N_13752,N_13465);
and UO_1337 (O_1337,N_14427,N_14081);
and UO_1338 (O_1338,N_13776,N_13156);
xor UO_1339 (O_1339,N_13971,N_13517);
nor UO_1340 (O_1340,N_14788,N_14156);
nand UO_1341 (O_1341,N_12603,N_13247);
xor UO_1342 (O_1342,N_12323,N_14533);
or UO_1343 (O_1343,N_13580,N_14802);
nand UO_1344 (O_1344,N_14912,N_12729);
nand UO_1345 (O_1345,N_13774,N_12083);
or UO_1346 (O_1346,N_12365,N_13245);
xor UO_1347 (O_1347,N_14214,N_13745);
nand UO_1348 (O_1348,N_13800,N_12710);
and UO_1349 (O_1349,N_12240,N_14704);
nor UO_1350 (O_1350,N_13738,N_14167);
xor UO_1351 (O_1351,N_14502,N_14074);
nand UO_1352 (O_1352,N_14749,N_14332);
nor UO_1353 (O_1353,N_13001,N_14047);
xnor UO_1354 (O_1354,N_13270,N_13493);
or UO_1355 (O_1355,N_12309,N_14750);
or UO_1356 (O_1356,N_14094,N_12635);
or UO_1357 (O_1357,N_13430,N_14848);
nand UO_1358 (O_1358,N_13972,N_14702);
nor UO_1359 (O_1359,N_14560,N_13406);
nor UO_1360 (O_1360,N_12616,N_12442);
and UO_1361 (O_1361,N_12464,N_14206);
nor UO_1362 (O_1362,N_12094,N_12691);
and UO_1363 (O_1363,N_13206,N_12519);
nor UO_1364 (O_1364,N_13607,N_13629);
nand UO_1365 (O_1365,N_13346,N_13750);
xor UO_1366 (O_1366,N_12203,N_14062);
nor UO_1367 (O_1367,N_13490,N_12628);
and UO_1368 (O_1368,N_13555,N_12034);
nand UO_1369 (O_1369,N_12319,N_13966);
nor UO_1370 (O_1370,N_14395,N_12012);
nor UO_1371 (O_1371,N_12692,N_14136);
nand UO_1372 (O_1372,N_14636,N_12093);
or UO_1373 (O_1373,N_14038,N_14119);
nand UO_1374 (O_1374,N_12398,N_13348);
nand UO_1375 (O_1375,N_12461,N_13338);
or UO_1376 (O_1376,N_13067,N_13065);
or UO_1377 (O_1377,N_14291,N_14344);
nor UO_1378 (O_1378,N_14486,N_14616);
nor UO_1379 (O_1379,N_13947,N_12685);
and UO_1380 (O_1380,N_12992,N_13461);
nand UO_1381 (O_1381,N_14134,N_12124);
and UO_1382 (O_1382,N_13120,N_13813);
nor UO_1383 (O_1383,N_14752,N_13272);
nor UO_1384 (O_1384,N_12899,N_12763);
nor UO_1385 (O_1385,N_14808,N_14737);
nand UO_1386 (O_1386,N_14728,N_14722);
nand UO_1387 (O_1387,N_13876,N_14104);
xor UO_1388 (O_1388,N_13568,N_14246);
and UO_1389 (O_1389,N_12738,N_13827);
or UO_1390 (O_1390,N_13720,N_12753);
nand UO_1391 (O_1391,N_13671,N_12471);
nor UO_1392 (O_1392,N_12227,N_14723);
or UO_1393 (O_1393,N_13454,N_14135);
nand UO_1394 (O_1394,N_12355,N_14921);
xnor UO_1395 (O_1395,N_14944,N_12501);
and UO_1396 (O_1396,N_12002,N_13331);
or UO_1397 (O_1397,N_13342,N_12905);
nor UO_1398 (O_1398,N_12718,N_12033);
xnor UO_1399 (O_1399,N_13934,N_14493);
or UO_1400 (O_1400,N_14442,N_14892);
and UO_1401 (O_1401,N_13900,N_13164);
xor UO_1402 (O_1402,N_13571,N_12016);
or UO_1403 (O_1403,N_14926,N_12759);
or UO_1404 (O_1404,N_14375,N_14717);
nor UO_1405 (O_1405,N_13419,N_14060);
and UO_1406 (O_1406,N_12831,N_14201);
or UO_1407 (O_1407,N_12459,N_12162);
nand UO_1408 (O_1408,N_12615,N_12810);
nand UO_1409 (O_1409,N_13418,N_12287);
and UO_1410 (O_1410,N_13479,N_12040);
nand UO_1411 (O_1411,N_13693,N_14073);
nand UO_1412 (O_1412,N_14042,N_12816);
and UO_1413 (O_1413,N_13503,N_12462);
nand UO_1414 (O_1414,N_14747,N_14610);
nand UO_1415 (O_1415,N_12474,N_14873);
and UO_1416 (O_1416,N_14535,N_14325);
nor UO_1417 (O_1417,N_13239,N_12056);
and UO_1418 (O_1418,N_12737,N_13054);
xor UO_1419 (O_1419,N_12127,N_13082);
nor UO_1420 (O_1420,N_12757,N_13511);
or UO_1421 (O_1421,N_14033,N_13929);
nor UO_1422 (O_1422,N_12987,N_12998);
nor UO_1423 (O_1423,N_13084,N_12144);
or UO_1424 (O_1424,N_13566,N_12885);
or UO_1425 (O_1425,N_12327,N_14634);
nand UO_1426 (O_1426,N_13300,N_14801);
xor UO_1427 (O_1427,N_14522,N_13293);
and UO_1428 (O_1428,N_14966,N_13073);
or UO_1429 (O_1429,N_14574,N_12390);
nand UO_1430 (O_1430,N_14929,N_14615);
nor UO_1431 (O_1431,N_12312,N_14468);
nand UO_1432 (O_1432,N_12997,N_14056);
xor UO_1433 (O_1433,N_12045,N_13216);
xor UO_1434 (O_1434,N_13422,N_14496);
or UO_1435 (O_1435,N_14240,N_14307);
nand UO_1436 (O_1436,N_12043,N_12595);
and UO_1437 (O_1437,N_13354,N_14361);
nand UO_1438 (O_1438,N_12429,N_14947);
xor UO_1439 (O_1439,N_12890,N_13382);
xor UO_1440 (O_1440,N_12650,N_13238);
xnor UO_1441 (O_1441,N_12719,N_13858);
nor UO_1442 (O_1442,N_13851,N_14381);
or UO_1443 (O_1443,N_13439,N_14303);
nor UO_1444 (O_1444,N_14009,N_12778);
or UO_1445 (O_1445,N_13266,N_13899);
nor UO_1446 (O_1446,N_14559,N_13531);
nor UO_1447 (O_1447,N_13453,N_14986);
nor UO_1448 (O_1448,N_12600,N_13102);
nand UO_1449 (O_1449,N_13861,N_12972);
xor UO_1450 (O_1450,N_12516,N_14899);
nand UO_1451 (O_1451,N_14218,N_12725);
or UO_1452 (O_1452,N_13540,N_14949);
nand UO_1453 (O_1453,N_13684,N_13625);
nor UO_1454 (O_1454,N_13613,N_12620);
nand UO_1455 (O_1455,N_12793,N_13027);
and UO_1456 (O_1456,N_12632,N_14087);
or UO_1457 (O_1457,N_12536,N_12966);
or UO_1458 (O_1458,N_13441,N_12064);
nand UO_1459 (O_1459,N_12674,N_12134);
nand UO_1460 (O_1460,N_13928,N_14035);
or UO_1461 (O_1461,N_14618,N_14435);
nor UO_1462 (O_1462,N_13376,N_13034);
and UO_1463 (O_1463,N_13524,N_12864);
nor UO_1464 (O_1464,N_14602,N_12938);
xor UO_1465 (O_1465,N_14985,N_12706);
and UO_1466 (O_1466,N_13578,N_12062);
or UO_1467 (O_1467,N_14619,N_14859);
nor UO_1468 (O_1468,N_12306,N_13721);
nor UO_1469 (O_1469,N_12335,N_13189);
xnor UO_1470 (O_1470,N_12901,N_13656);
or UO_1471 (O_1471,N_13127,N_14416);
or UO_1472 (O_1472,N_12790,N_14556);
and UO_1473 (O_1473,N_13759,N_12699);
nand UO_1474 (O_1474,N_14733,N_12876);
nor UO_1475 (O_1475,N_14932,N_13151);
or UO_1476 (O_1476,N_14711,N_13128);
and UO_1477 (O_1477,N_12599,N_13103);
nand UO_1478 (O_1478,N_13744,N_12745);
and UO_1479 (O_1479,N_12432,N_14222);
nor UO_1480 (O_1480,N_12565,N_12851);
and UO_1481 (O_1481,N_14821,N_14282);
nor UO_1482 (O_1482,N_14195,N_12050);
and UO_1483 (O_1483,N_14100,N_14155);
nor UO_1484 (O_1484,N_14423,N_12493);
and UO_1485 (O_1485,N_13271,N_13539);
nand UO_1486 (O_1486,N_13023,N_12449);
or UO_1487 (O_1487,N_13169,N_14977);
and UO_1488 (O_1488,N_12444,N_12878);
or UO_1489 (O_1489,N_12837,N_13146);
xor UO_1490 (O_1490,N_13351,N_13368);
and UO_1491 (O_1491,N_12772,N_14036);
nor UO_1492 (O_1492,N_12305,N_14254);
nand UO_1493 (O_1493,N_14492,N_13651);
or UO_1494 (O_1494,N_13575,N_13818);
nand UO_1495 (O_1495,N_14534,N_13096);
and UO_1496 (O_1496,N_13476,N_13125);
nor UO_1497 (O_1497,N_12645,N_13283);
nand UO_1498 (O_1498,N_13372,N_13634);
and UO_1499 (O_1499,N_13284,N_12263);
and UO_1500 (O_1500,N_12660,N_13324);
or UO_1501 (O_1501,N_12927,N_12510);
or UO_1502 (O_1502,N_14894,N_12526);
nor UO_1503 (O_1503,N_13701,N_14689);
or UO_1504 (O_1504,N_14300,N_13543);
and UO_1505 (O_1505,N_14231,N_12480);
nor UO_1506 (O_1506,N_14891,N_12229);
or UO_1507 (O_1507,N_12549,N_12073);
nor UO_1508 (O_1508,N_13773,N_12977);
or UO_1509 (O_1509,N_14215,N_13713);
or UO_1510 (O_1510,N_13409,N_14536);
nand UO_1511 (O_1511,N_14904,N_12292);
and UO_1512 (O_1512,N_13713,N_14037);
xor UO_1513 (O_1513,N_12093,N_13982);
xor UO_1514 (O_1514,N_14213,N_12949);
nand UO_1515 (O_1515,N_14017,N_13416);
xor UO_1516 (O_1516,N_13221,N_12488);
nand UO_1517 (O_1517,N_12941,N_12496);
nand UO_1518 (O_1518,N_12396,N_12515);
and UO_1519 (O_1519,N_13048,N_12438);
nand UO_1520 (O_1520,N_13540,N_12019);
and UO_1521 (O_1521,N_13403,N_12048);
and UO_1522 (O_1522,N_13651,N_12352);
and UO_1523 (O_1523,N_14628,N_14923);
and UO_1524 (O_1524,N_14781,N_13106);
nand UO_1525 (O_1525,N_12270,N_14898);
nor UO_1526 (O_1526,N_13340,N_14571);
nand UO_1527 (O_1527,N_12921,N_12722);
xor UO_1528 (O_1528,N_12967,N_13168);
or UO_1529 (O_1529,N_14614,N_14915);
or UO_1530 (O_1530,N_13540,N_13574);
and UO_1531 (O_1531,N_12621,N_12094);
nand UO_1532 (O_1532,N_13182,N_12079);
or UO_1533 (O_1533,N_13416,N_14299);
nor UO_1534 (O_1534,N_12125,N_13402);
nand UO_1535 (O_1535,N_12719,N_14650);
and UO_1536 (O_1536,N_12055,N_13091);
xnor UO_1537 (O_1537,N_12316,N_14442);
nand UO_1538 (O_1538,N_12166,N_13117);
nand UO_1539 (O_1539,N_12092,N_13016);
nor UO_1540 (O_1540,N_13742,N_13012);
and UO_1541 (O_1541,N_14823,N_12445);
or UO_1542 (O_1542,N_13177,N_12334);
nand UO_1543 (O_1543,N_13060,N_12116);
and UO_1544 (O_1544,N_13938,N_13744);
xor UO_1545 (O_1545,N_13556,N_12958);
nand UO_1546 (O_1546,N_12931,N_12897);
or UO_1547 (O_1547,N_14205,N_13325);
nand UO_1548 (O_1548,N_14745,N_14494);
nand UO_1549 (O_1549,N_13942,N_13604);
nor UO_1550 (O_1550,N_14842,N_12663);
nor UO_1551 (O_1551,N_12578,N_13510);
nor UO_1552 (O_1552,N_14797,N_14480);
nor UO_1553 (O_1553,N_14239,N_14794);
nand UO_1554 (O_1554,N_13659,N_14928);
and UO_1555 (O_1555,N_14347,N_13339);
nor UO_1556 (O_1556,N_14497,N_13233);
or UO_1557 (O_1557,N_14328,N_13399);
or UO_1558 (O_1558,N_13997,N_13915);
nand UO_1559 (O_1559,N_13102,N_12382);
nand UO_1560 (O_1560,N_13984,N_14518);
and UO_1561 (O_1561,N_12012,N_12583);
xor UO_1562 (O_1562,N_13261,N_14739);
nand UO_1563 (O_1563,N_12104,N_14038);
or UO_1564 (O_1564,N_13210,N_14977);
or UO_1565 (O_1565,N_13342,N_12343);
and UO_1566 (O_1566,N_14820,N_14500);
or UO_1567 (O_1567,N_12862,N_12570);
xor UO_1568 (O_1568,N_13716,N_12255);
or UO_1569 (O_1569,N_14181,N_14541);
or UO_1570 (O_1570,N_14911,N_12381);
nand UO_1571 (O_1571,N_12335,N_14801);
or UO_1572 (O_1572,N_13310,N_13720);
and UO_1573 (O_1573,N_12283,N_12542);
xor UO_1574 (O_1574,N_14394,N_14492);
and UO_1575 (O_1575,N_13916,N_12531);
and UO_1576 (O_1576,N_12506,N_14093);
nand UO_1577 (O_1577,N_14238,N_13089);
nand UO_1578 (O_1578,N_14460,N_14420);
nor UO_1579 (O_1579,N_13936,N_13441);
xor UO_1580 (O_1580,N_12568,N_13627);
xnor UO_1581 (O_1581,N_13415,N_12882);
or UO_1582 (O_1582,N_13860,N_12181);
and UO_1583 (O_1583,N_12670,N_13361);
nand UO_1584 (O_1584,N_14221,N_13787);
nor UO_1585 (O_1585,N_13564,N_13358);
nor UO_1586 (O_1586,N_12636,N_12035);
nor UO_1587 (O_1587,N_12588,N_12631);
and UO_1588 (O_1588,N_12736,N_13279);
and UO_1589 (O_1589,N_14447,N_12073);
and UO_1590 (O_1590,N_13005,N_13836);
nor UO_1591 (O_1591,N_14071,N_13264);
nand UO_1592 (O_1592,N_12647,N_12506);
nand UO_1593 (O_1593,N_13255,N_12926);
nor UO_1594 (O_1594,N_12811,N_14723);
and UO_1595 (O_1595,N_13507,N_14216);
nand UO_1596 (O_1596,N_12629,N_12635);
or UO_1597 (O_1597,N_13616,N_12819);
xnor UO_1598 (O_1598,N_13329,N_14608);
xor UO_1599 (O_1599,N_13027,N_14114);
xnor UO_1600 (O_1600,N_13705,N_12529);
or UO_1601 (O_1601,N_12251,N_12548);
xnor UO_1602 (O_1602,N_14579,N_13998);
and UO_1603 (O_1603,N_14796,N_13098);
and UO_1604 (O_1604,N_14584,N_12614);
xor UO_1605 (O_1605,N_12101,N_12288);
and UO_1606 (O_1606,N_12430,N_12969);
nor UO_1607 (O_1607,N_12650,N_14021);
nand UO_1608 (O_1608,N_14217,N_13857);
nand UO_1609 (O_1609,N_13072,N_13326);
and UO_1610 (O_1610,N_12305,N_13691);
or UO_1611 (O_1611,N_13148,N_13556);
or UO_1612 (O_1612,N_14901,N_12047);
and UO_1613 (O_1613,N_14008,N_14711);
or UO_1614 (O_1614,N_14404,N_12778);
and UO_1615 (O_1615,N_14349,N_13516);
and UO_1616 (O_1616,N_14216,N_12908);
nor UO_1617 (O_1617,N_14392,N_13008);
nor UO_1618 (O_1618,N_14949,N_12720);
xor UO_1619 (O_1619,N_14704,N_12380);
nand UO_1620 (O_1620,N_13139,N_14445);
nand UO_1621 (O_1621,N_12518,N_13584);
and UO_1622 (O_1622,N_13805,N_14049);
nand UO_1623 (O_1623,N_12692,N_13436);
nand UO_1624 (O_1624,N_13367,N_14457);
or UO_1625 (O_1625,N_13839,N_12642);
and UO_1626 (O_1626,N_13764,N_12167);
and UO_1627 (O_1627,N_12600,N_12566);
xor UO_1628 (O_1628,N_13346,N_12826);
xnor UO_1629 (O_1629,N_13737,N_13914);
nand UO_1630 (O_1630,N_13127,N_13078);
or UO_1631 (O_1631,N_12857,N_13205);
nand UO_1632 (O_1632,N_12002,N_12130);
nor UO_1633 (O_1633,N_13395,N_13418);
nand UO_1634 (O_1634,N_14125,N_13425);
nand UO_1635 (O_1635,N_13834,N_12444);
or UO_1636 (O_1636,N_14075,N_12614);
nor UO_1637 (O_1637,N_14299,N_14367);
or UO_1638 (O_1638,N_14866,N_12552);
or UO_1639 (O_1639,N_14096,N_14434);
and UO_1640 (O_1640,N_14675,N_13005);
or UO_1641 (O_1641,N_13334,N_13498);
nand UO_1642 (O_1642,N_13402,N_14984);
or UO_1643 (O_1643,N_13015,N_12132);
nor UO_1644 (O_1644,N_13494,N_13362);
nand UO_1645 (O_1645,N_13014,N_14794);
nand UO_1646 (O_1646,N_13848,N_13351);
nor UO_1647 (O_1647,N_12346,N_12774);
and UO_1648 (O_1648,N_12401,N_13259);
or UO_1649 (O_1649,N_14717,N_12846);
nor UO_1650 (O_1650,N_13777,N_14085);
and UO_1651 (O_1651,N_13000,N_13316);
nor UO_1652 (O_1652,N_13284,N_12902);
or UO_1653 (O_1653,N_14702,N_12638);
or UO_1654 (O_1654,N_13681,N_13087);
nor UO_1655 (O_1655,N_14947,N_13847);
nand UO_1656 (O_1656,N_13293,N_13443);
nor UO_1657 (O_1657,N_12028,N_13620);
or UO_1658 (O_1658,N_13274,N_12206);
nand UO_1659 (O_1659,N_12501,N_12373);
nand UO_1660 (O_1660,N_12273,N_12254);
nor UO_1661 (O_1661,N_14280,N_12699);
nand UO_1662 (O_1662,N_14870,N_12440);
or UO_1663 (O_1663,N_14048,N_13468);
and UO_1664 (O_1664,N_14043,N_14912);
xnor UO_1665 (O_1665,N_13231,N_14949);
nand UO_1666 (O_1666,N_12817,N_14824);
and UO_1667 (O_1667,N_14802,N_14819);
nand UO_1668 (O_1668,N_13167,N_13409);
nor UO_1669 (O_1669,N_13249,N_14718);
xnor UO_1670 (O_1670,N_12277,N_12932);
xor UO_1671 (O_1671,N_13840,N_12231);
or UO_1672 (O_1672,N_12154,N_13188);
nand UO_1673 (O_1673,N_12740,N_14543);
and UO_1674 (O_1674,N_14243,N_12226);
xor UO_1675 (O_1675,N_14565,N_14517);
nor UO_1676 (O_1676,N_13152,N_14052);
xor UO_1677 (O_1677,N_13683,N_13497);
nand UO_1678 (O_1678,N_12845,N_14963);
and UO_1679 (O_1679,N_12572,N_12219);
nand UO_1680 (O_1680,N_13381,N_12543);
nor UO_1681 (O_1681,N_12406,N_14271);
nand UO_1682 (O_1682,N_12405,N_12922);
or UO_1683 (O_1683,N_14428,N_14580);
or UO_1684 (O_1684,N_12108,N_12429);
nor UO_1685 (O_1685,N_12203,N_14480);
and UO_1686 (O_1686,N_13646,N_13724);
nand UO_1687 (O_1687,N_13582,N_13414);
and UO_1688 (O_1688,N_13252,N_14256);
and UO_1689 (O_1689,N_13562,N_13162);
nor UO_1690 (O_1690,N_12714,N_13583);
or UO_1691 (O_1691,N_12104,N_12751);
nand UO_1692 (O_1692,N_14311,N_14070);
nand UO_1693 (O_1693,N_14839,N_13329);
and UO_1694 (O_1694,N_14985,N_13356);
nor UO_1695 (O_1695,N_12665,N_13908);
nor UO_1696 (O_1696,N_13714,N_13101);
nand UO_1697 (O_1697,N_12440,N_12567);
and UO_1698 (O_1698,N_14194,N_12500);
nand UO_1699 (O_1699,N_12698,N_13810);
or UO_1700 (O_1700,N_12004,N_13054);
nor UO_1701 (O_1701,N_12213,N_14872);
nand UO_1702 (O_1702,N_14191,N_13551);
and UO_1703 (O_1703,N_13793,N_14327);
or UO_1704 (O_1704,N_14407,N_13250);
nor UO_1705 (O_1705,N_13778,N_12724);
nand UO_1706 (O_1706,N_12209,N_12624);
nor UO_1707 (O_1707,N_13925,N_14973);
nor UO_1708 (O_1708,N_14990,N_13814);
or UO_1709 (O_1709,N_12707,N_14656);
xor UO_1710 (O_1710,N_14157,N_14463);
and UO_1711 (O_1711,N_13142,N_12213);
nand UO_1712 (O_1712,N_12055,N_14748);
nand UO_1713 (O_1713,N_14731,N_12587);
xnor UO_1714 (O_1714,N_13492,N_12699);
or UO_1715 (O_1715,N_13495,N_14358);
nand UO_1716 (O_1716,N_12041,N_12611);
nand UO_1717 (O_1717,N_14478,N_14304);
nor UO_1718 (O_1718,N_12832,N_12033);
or UO_1719 (O_1719,N_14778,N_14044);
nand UO_1720 (O_1720,N_12485,N_14623);
or UO_1721 (O_1721,N_13756,N_13281);
nand UO_1722 (O_1722,N_12150,N_12978);
and UO_1723 (O_1723,N_12137,N_13115);
nand UO_1724 (O_1724,N_14021,N_13027);
nor UO_1725 (O_1725,N_12904,N_14690);
nor UO_1726 (O_1726,N_12641,N_13951);
or UO_1727 (O_1727,N_13146,N_12149);
or UO_1728 (O_1728,N_12448,N_14327);
nand UO_1729 (O_1729,N_14501,N_14603);
nor UO_1730 (O_1730,N_14556,N_14791);
and UO_1731 (O_1731,N_13263,N_13464);
nor UO_1732 (O_1732,N_12019,N_12593);
nand UO_1733 (O_1733,N_14568,N_12223);
nor UO_1734 (O_1734,N_14569,N_14433);
nand UO_1735 (O_1735,N_13259,N_12301);
nand UO_1736 (O_1736,N_13125,N_12586);
nor UO_1737 (O_1737,N_13770,N_13426);
nor UO_1738 (O_1738,N_14753,N_12176);
nor UO_1739 (O_1739,N_13696,N_12874);
xnor UO_1740 (O_1740,N_12022,N_13027);
nor UO_1741 (O_1741,N_12958,N_14229);
and UO_1742 (O_1742,N_13151,N_14156);
nor UO_1743 (O_1743,N_14103,N_14819);
nand UO_1744 (O_1744,N_12671,N_13350);
xor UO_1745 (O_1745,N_12593,N_12830);
or UO_1746 (O_1746,N_12492,N_13852);
nor UO_1747 (O_1747,N_13128,N_14485);
or UO_1748 (O_1748,N_14099,N_13644);
nor UO_1749 (O_1749,N_13931,N_13399);
and UO_1750 (O_1750,N_12332,N_13427);
and UO_1751 (O_1751,N_12505,N_12087);
nor UO_1752 (O_1752,N_13982,N_12503);
nor UO_1753 (O_1753,N_12685,N_12322);
and UO_1754 (O_1754,N_12462,N_12871);
nand UO_1755 (O_1755,N_14282,N_14543);
and UO_1756 (O_1756,N_14486,N_13394);
and UO_1757 (O_1757,N_12273,N_14496);
and UO_1758 (O_1758,N_13842,N_13538);
nand UO_1759 (O_1759,N_12775,N_12987);
nand UO_1760 (O_1760,N_13473,N_13275);
and UO_1761 (O_1761,N_13757,N_14330);
nand UO_1762 (O_1762,N_14641,N_12973);
nand UO_1763 (O_1763,N_14694,N_13434);
and UO_1764 (O_1764,N_14123,N_14817);
and UO_1765 (O_1765,N_14720,N_13079);
nor UO_1766 (O_1766,N_12473,N_14161);
nor UO_1767 (O_1767,N_14138,N_14507);
nor UO_1768 (O_1768,N_14648,N_12358);
and UO_1769 (O_1769,N_14973,N_12532);
nand UO_1770 (O_1770,N_14373,N_12216);
nor UO_1771 (O_1771,N_13641,N_13959);
and UO_1772 (O_1772,N_12058,N_12412);
nor UO_1773 (O_1773,N_12085,N_13266);
nand UO_1774 (O_1774,N_14269,N_13441);
or UO_1775 (O_1775,N_12927,N_13284);
xnor UO_1776 (O_1776,N_14736,N_13230);
or UO_1777 (O_1777,N_12243,N_14290);
xnor UO_1778 (O_1778,N_13137,N_13938);
or UO_1779 (O_1779,N_14892,N_14671);
nor UO_1780 (O_1780,N_14940,N_13798);
xor UO_1781 (O_1781,N_12109,N_13906);
nand UO_1782 (O_1782,N_12167,N_14879);
nor UO_1783 (O_1783,N_13478,N_13431);
nand UO_1784 (O_1784,N_12184,N_12510);
xor UO_1785 (O_1785,N_14558,N_14043);
and UO_1786 (O_1786,N_13657,N_13610);
or UO_1787 (O_1787,N_13854,N_13251);
and UO_1788 (O_1788,N_12584,N_13968);
or UO_1789 (O_1789,N_14393,N_14137);
xnor UO_1790 (O_1790,N_13145,N_12958);
nand UO_1791 (O_1791,N_12389,N_13735);
and UO_1792 (O_1792,N_12125,N_14556);
and UO_1793 (O_1793,N_13575,N_12160);
nor UO_1794 (O_1794,N_12089,N_14441);
and UO_1795 (O_1795,N_14193,N_12563);
and UO_1796 (O_1796,N_13452,N_12481);
and UO_1797 (O_1797,N_14636,N_14361);
and UO_1798 (O_1798,N_14980,N_12142);
nand UO_1799 (O_1799,N_12913,N_13533);
nand UO_1800 (O_1800,N_12257,N_14550);
or UO_1801 (O_1801,N_13507,N_12691);
xnor UO_1802 (O_1802,N_12465,N_13743);
nor UO_1803 (O_1803,N_12685,N_13914);
or UO_1804 (O_1804,N_12516,N_12215);
and UO_1805 (O_1805,N_14756,N_14035);
and UO_1806 (O_1806,N_14812,N_12322);
and UO_1807 (O_1807,N_13302,N_12373);
nand UO_1808 (O_1808,N_12587,N_12926);
and UO_1809 (O_1809,N_13433,N_12273);
xor UO_1810 (O_1810,N_12480,N_13271);
and UO_1811 (O_1811,N_14254,N_12171);
nor UO_1812 (O_1812,N_13290,N_14851);
nand UO_1813 (O_1813,N_12329,N_12007);
nand UO_1814 (O_1814,N_13009,N_12329);
nand UO_1815 (O_1815,N_13748,N_13078);
and UO_1816 (O_1816,N_14628,N_12990);
and UO_1817 (O_1817,N_13818,N_12803);
nor UO_1818 (O_1818,N_12522,N_12177);
nor UO_1819 (O_1819,N_13646,N_12905);
nor UO_1820 (O_1820,N_13123,N_14164);
and UO_1821 (O_1821,N_12444,N_12409);
xor UO_1822 (O_1822,N_14210,N_13548);
nor UO_1823 (O_1823,N_12752,N_12879);
and UO_1824 (O_1824,N_13030,N_12403);
nor UO_1825 (O_1825,N_12766,N_14370);
and UO_1826 (O_1826,N_12926,N_13286);
or UO_1827 (O_1827,N_14006,N_14984);
xnor UO_1828 (O_1828,N_14490,N_14067);
and UO_1829 (O_1829,N_13515,N_13323);
nor UO_1830 (O_1830,N_12767,N_13121);
nor UO_1831 (O_1831,N_13136,N_13998);
nor UO_1832 (O_1832,N_14015,N_13788);
and UO_1833 (O_1833,N_14592,N_13754);
xnor UO_1834 (O_1834,N_13226,N_13329);
and UO_1835 (O_1835,N_13635,N_13023);
nand UO_1836 (O_1836,N_12551,N_14291);
nor UO_1837 (O_1837,N_12833,N_14207);
nand UO_1838 (O_1838,N_12808,N_13137);
and UO_1839 (O_1839,N_14948,N_13490);
nor UO_1840 (O_1840,N_14597,N_12176);
and UO_1841 (O_1841,N_12274,N_13625);
and UO_1842 (O_1842,N_12611,N_14289);
nand UO_1843 (O_1843,N_13467,N_14096);
nand UO_1844 (O_1844,N_12482,N_14102);
and UO_1845 (O_1845,N_13730,N_12907);
nor UO_1846 (O_1846,N_12052,N_13325);
or UO_1847 (O_1847,N_14210,N_12944);
nor UO_1848 (O_1848,N_12384,N_12373);
nand UO_1849 (O_1849,N_13144,N_12603);
and UO_1850 (O_1850,N_12108,N_13377);
and UO_1851 (O_1851,N_14520,N_13027);
nor UO_1852 (O_1852,N_12970,N_14082);
nand UO_1853 (O_1853,N_14266,N_12842);
or UO_1854 (O_1854,N_12476,N_13298);
xnor UO_1855 (O_1855,N_14617,N_14109);
nand UO_1856 (O_1856,N_12391,N_12241);
xor UO_1857 (O_1857,N_13131,N_13127);
or UO_1858 (O_1858,N_14578,N_13220);
nand UO_1859 (O_1859,N_12975,N_12195);
or UO_1860 (O_1860,N_14228,N_13242);
nor UO_1861 (O_1861,N_13135,N_13064);
nand UO_1862 (O_1862,N_13555,N_13711);
nand UO_1863 (O_1863,N_13581,N_14420);
nand UO_1864 (O_1864,N_12162,N_13077);
and UO_1865 (O_1865,N_14332,N_13825);
or UO_1866 (O_1866,N_14644,N_14582);
and UO_1867 (O_1867,N_13399,N_12011);
nand UO_1868 (O_1868,N_13677,N_12202);
nand UO_1869 (O_1869,N_13408,N_12267);
and UO_1870 (O_1870,N_12025,N_13047);
and UO_1871 (O_1871,N_13228,N_14319);
or UO_1872 (O_1872,N_13066,N_13973);
and UO_1873 (O_1873,N_12368,N_14535);
and UO_1874 (O_1874,N_14570,N_13260);
nand UO_1875 (O_1875,N_12592,N_12086);
nor UO_1876 (O_1876,N_12370,N_12028);
nand UO_1877 (O_1877,N_14349,N_12669);
nand UO_1878 (O_1878,N_12784,N_13993);
and UO_1879 (O_1879,N_12967,N_14887);
nand UO_1880 (O_1880,N_13579,N_12225);
nor UO_1881 (O_1881,N_14661,N_12526);
nor UO_1882 (O_1882,N_14869,N_14868);
nor UO_1883 (O_1883,N_12781,N_12855);
or UO_1884 (O_1884,N_13177,N_12229);
and UO_1885 (O_1885,N_13421,N_13534);
nand UO_1886 (O_1886,N_12376,N_13461);
nor UO_1887 (O_1887,N_13272,N_13317);
xor UO_1888 (O_1888,N_12474,N_13648);
nor UO_1889 (O_1889,N_12602,N_14166);
or UO_1890 (O_1890,N_12996,N_12220);
nor UO_1891 (O_1891,N_13614,N_13065);
and UO_1892 (O_1892,N_14291,N_13316);
or UO_1893 (O_1893,N_13018,N_13589);
xnor UO_1894 (O_1894,N_13860,N_12707);
nand UO_1895 (O_1895,N_12371,N_13427);
xor UO_1896 (O_1896,N_14106,N_14827);
or UO_1897 (O_1897,N_13523,N_14847);
nor UO_1898 (O_1898,N_14886,N_12594);
or UO_1899 (O_1899,N_13900,N_13248);
or UO_1900 (O_1900,N_14696,N_12774);
nand UO_1901 (O_1901,N_14516,N_13883);
nor UO_1902 (O_1902,N_14718,N_12076);
nor UO_1903 (O_1903,N_13528,N_13786);
or UO_1904 (O_1904,N_12709,N_13846);
and UO_1905 (O_1905,N_14592,N_14708);
and UO_1906 (O_1906,N_14832,N_13578);
nand UO_1907 (O_1907,N_12890,N_14608);
nand UO_1908 (O_1908,N_12553,N_13364);
nor UO_1909 (O_1909,N_13394,N_13823);
or UO_1910 (O_1910,N_14428,N_12355);
nor UO_1911 (O_1911,N_14555,N_14851);
or UO_1912 (O_1912,N_13762,N_12144);
nand UO_1913 (O_1913,N_12670,N_13967);
or UO_1914 (O_1914,N_14399,N_12073);
and UO_1915 (O_1915,N_14014,N_14641);
or UO_1916 (O_1916,N_12585,N_14106);
and UO_1917 (O_1917,N_13209,N_12412);
and UO_1918 (O_1918,N_13391,N_12266);
and UO_1919 (O_1919,N_14092,N_13572);
xnor UO_1920 (O_1920,N_14846,N_14901);
nand UO_1921 (O_1921,N_14332,N_12105);
and UO_1922 (O_1922,N_14283,N_13612);
nand UO_1923 (O_1923,N_13522,N_14444);
or UO_1924 (O_1924,N_13819,N_13674);
or UO_1925 (O_1925,N_13368,N_14208);
nor UO_1926 (O_1926,N_13569,N_12568);
and UO_1927 (O_1927,N_14655,N_12404);
nor UO_1928 (O_1928,N_14555,N_14994);
nor UO_1929 (O_1929,N_13883,N_13034);
and UO_1930 (O_1930,N_13052,N_12627);
and UO_1931 (O_1931,N_13161,N_13502);
xnor UO_1932 (O_1932,N_13234,N_12984);
and UO_1933 (O_1933,N_13393,N_12024);
nor UO_1934 (O_1934,N_12649,N_12940);
nand UO_1935 (O_1935,N_13102,N_12383);
nor UO_1936 (O_1936,N_12732,N_14686);
xor UO_1937 (O_1937,N_14371,N_12219);
nand UO_1938 (O_1938,N_12025,N_12546);
or UO_1939 (O_1939,N_13460,N_14496);
or UO_1940 (O_1940,N_14887,N_12859);
or UO_1941 (O_1941,N_14138,N_13547);
or UO_1942 (O_1942,N_13179,N_14544);
nor UO_1943 (O_1943,N_12828,N_14174);
nand UO_1944 (O_1944,N_13508,N_14551);
nor UO_1945 (O_1945,N_13396,N_12067);
and UO_1946 (O_1946,N_14835,N_12755);
nor UO_1947 (O_1947,N_13141,N_12174);
nand UO_1948 (O_1948,N_13983,N_13836);
and UO_1949 (O_1949,N_14445,N_13467);
nand UO_1950 (O_1950,N_12535,N_13448);
nor UO_1951 (O_1951,N_13944,N_13661);
and UO_1952 (O_1952,N_14433,N_13641);
and UO_1953 (O_1953,N_12505,N_12409);
and UO_1954 (O_1954,N_14109,N_13370);
and UO_1955 (O_1955,N_12628,N_13420);
nor UO_1956 (O_1956,N_12084,N_13892);
nand UO_1957 (O_1957,N_12235,N_14026);
nand UO_1958 (O_1958,N_13623,N_14713);
and UO_1959 (O_1959,N_13386,N_13395);
nand UO_1960 (O_1960,N_14457,N_14142);
nor UO_1961 (O_1961,N_13443,N_14708);
or UO_1962 (O_1962,N_13984,N_13124);
nor UO_1963 (O_1963,N_13055,N_14701);
and UO_1964 (O_1964,N_13146,N_14097);
nand UO_1965 (O_1965,N_13397,N_14168);
nor UO_1966 (O_1966,N_13354,N_12435);
or UO_1967 (O_1967,N_14576,N_14116);
and UO_1968 (O_1968,N_12361,N_13138);
and UO_1969 (O_1969,N_14982,N_12810);
or UO_1970 (O_1970,N_13831,N_13901);
or UO_1971 (O_1971,N_14321,N_12582);
or UO_1972 (O_1972,N_14210,N_14495);
or UO_1973 (O_1973,N_14593,N_14125);
or UO_1974 (O_1974,N_12358,N_14206);
or UO_1975 (O_1975,N_12796,N_13537);
nor UO_1976 (O_1976,N_14001,N_12054);
or UO_1977 (O_1977,N_13682,N_14646);
or UO_1978 (O_1978,N_12730,N_14585);
and UO_1979 (O_1979,N_13340,N_14498);
nand UO_1980 (O_1980,N_13581,N_12857);
nand UO_1981 (O_1981,N_14692,N_13712);
or UO_1982 (O_1982,N_14279,N_13650);
and UO_1983 (O_1983,N_13126,N_14624);
or UO_1984 (O_1984,N_14142,N_12333);
xnor UO_1985 (O_1985,N_14326,N_12929);
or UO_1986 (O_1986,N_12884,N_13919);
nor UO_1987 (O_1987,N_12020,N_12519);
or UO_1988 (O_1988,N_13974,N_13415);
or UO_1989 (O_1989,N_14471,N_12198);
xnor UO_1990 (O_1990,N_12426,N_12747);
xnor UO_1991 (O_1991,N_14355,N_14424);
nor UO_1992 (O_1992,N_13730,N_14297);
and UO_1993 (O_1993,N_13517,N_14663);
nand UO_1994 (O_1994,N_13251,N_13292);
nor UO_1995 (O_1995,N_14968,N_12807);
nand UO_1996 (O_1996,N_12045,N_14729);
and UO_1997 (O_1997,N_13300,N_13624);
xor UO_1998 (O_1998,N_12463,N_12455);
and UO_1999 (O_1999,N_13164,N_14922);
endmodule