module basic_3000_30000_3500_50_levels_5xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,In_2500,In_2501,In_2502,In_2503,In_2504,In_2505,In_2506,In_2507,In_2508,In_2509,In_2510,In_2511,In_2512,In_2513,In_2514,In_2515,In_2516,In_2517,In_2518,In_2519,In_2520,In_2521,In_2522,In_2523,In_2524,In_2525,In_2526,In_2527,In_2528,In_2529,In_2530,In_2531,In_2532,In_2533,In_2534,In_2535,In_2536,In_2537,In_2538,In_2539,In_2540,In_2541,In_2542,In_2543,In_2544,In_2545,In_2546,In_2547,In_2548,In_2549,In_2550,In_2551,In_2552,In_2553,In_2554,In_2555,In_2556,In_2557,In_2558,In_2559,In_2560,In_2561,In_2562,In_2563,In_2564,In_2565,In_2566,In_2567,In_2568,In_2569,In_2570,In_2571,In_2572,In_2573,In_2574,In_2575,In_2576,In_2577,In_2578,In_2579,In_2580,In_2581,In_2582,In_2583,In_2584,In_2585,In_2586,In_2587,In_2588,In_2589,In_2590,In_2591,In_2592,In_2593,In_2594,In_2595,In_2596,In_2597,In_2598,In_2599,In_2600,In_2601,In_2602,In_2603,In_2604,In_2605,In_2606,In_2607,In_2608,In_2609,In_2610,In_2611,In_2612,In_2613,In_2614,In_2615,In_2616,In_2617,In_2618,In_2619,In_2620,In_2621,In_2622,In_2623,In_2624,In_2625,In_2626,In_2627,In_2628,In_2629,In_2630,In_2631,In_2632,In_2633,In_2634,In_2635,In_2636,In_2637,In_2638,In_2639,In_2640,In_2641,In_2642,In_2643,In_2644,In_2645,In_2646,In_2647,In_2648,In_2649,In_2650,In_2651,In_2652,In_2653,In_2654,In_2655,In_2656,In_2657,In_2658,In_2659,In_2660,In_2661,In_2662,In_2663,In_2664,In_2665,In_2666,In_2667,In_2668,In_2669,In_2670,In_2671,In_2672,In_2673,In_2674,In_2675,In_2676,In_2677,In_2678,In_2679,In_2680,In_2681,In_2682,In_2683,In_2684,In_2685,In_2686,In_2687,In_2688,In_2689,In_2690,In_2691,In_2692,In_2693,In_2694,In_2695,In_2696,In_2697,In_2698,In_2699,In_2700,In_2701,In_2702,In_2703,In_2704,In_2705,In_2706,In_2707,In_2708,In_2709,In_2710,In_2711,In_2712,In_2713,In_2714,In_2715,In_2716,In_2717,In_2718,In_2719,In_2720,In_2721,In_2722,In_2723,In_2724,In_2725,In_2726,In_2727,In_2728,In_2729,In_2730,In_2731,In_2732,In_2733,In_2734,In_2735,In_2736,In_2737,In_2738,In_2739,In_2740,In_2741,In_2742,In_2743,In_2744,In_2745,In_2746,In_2747,In_2748,In_2749,In_2750,In_2751,In_2752,In_2753,In_2754,In_2755,In_2756,In_2757,In_2758,In_2759,In_2760,In_2761,In_2762,In_2763,In_2764,In_2765,In_2766,In_2767,In_2768,In_2769,In_2770,In_2771,In_2772,In_2773,In_2774,In_2775,In_2776,In_2777,In_2778,In_2779,In_2780,In_2781,In_2782,In_2783,In_2784,In_2785,In_2786,In_2787,In_2788,In_2789,In_2790,In_2791,In_2792,In_2793,In_2794,In_2795,In_2796,In_2797,In_2798,In_2799,In_2800,In_2801,In_2802,In_2803,In_2804,In_2805,In_2806,In_2807,In_2808,In_2809,In_2810,In_2811,In_2812,In_2813,In_2814,In_2815,In_2816,In_2817,In_2818,In_2819,In_2820,In_2821,In_2822,In_2823,In_2824,In_2825,In_2826,In_2827,In_2828,In_2829,In_2830,In_2831,In_2832,In_2833,In_2834,In_2835,In_2836,In_2837,In_2838,In_2839,In_2840,In_2841,In_2842,In_2843,In_2844,In_2845,In_2846,In_2847,In_2848,In_2849,In_2850,In_2851,In_2852,In_2853,In_2854,In_2855,In_2856,In_2857,In_2858,In_2859,In_2860,In_2861,In_2862,In_2863,In_2864,In_2865,In_2866,In_2867,In_2868,In_2869,In_2870,In_2871,In_2872,In_2873,In_2874,In_2875,In_2876,In_2877,In_2878,In_2879,In_2880,In_2881,In_2882,In_2883,In_2884,In_2885,In_2886,In_2887,In_2888,In_2889,In_2890,In_2891,In_2892,In_2893,In_2894,In_2895,In_2896,In_2897,In_2898,In_2899,In_2900,In_2901,In_2902,In_2903,In_2904,In_2905,In_2906,In_2907,In_2908,In_2909,In_2910,In_2911,In_2912,In_2913,In_2914,In_2915,In_2916,In_2917,In_2918,In_2919,In_2920,In_2921,In_2922,In_2923,In_2924,In_2925,In_2926,In_2927,In_2928,In_2929,In_2930,In_2931,In_2932,In_2933,In_2934,In_2935,In_2936,In_2937,In_2938,In_2939,In_2940,In_2941,In_2942,In_2943,In_2944,In_2945,In_2946,In_2947,In_2948,In_2949,In_2950,In_2951,In_2952,In_2953,In_2954,In_2955,In_2956,In_2957,In_2958,In_2959,In_2960,In_2961,In_2962,In_2963,In_2964,In_2965,In_2966,In_2967,In_2968,In_2969,In_2970,In_2971,In_2972,In_2973,In_2974,In_2975,In_2976,In_2977,In_2978,In_2979,In_2980,In_2981,In_2982,In_2983,In_2984,In_2985,In_2986,In_2987,In_2988,In_2989,In_2990,In_2991,In_2992,In_2993,In_2994,In_2995,In_2996,In_2997,In_2998,In_2999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999,O_3000,O_3001,O_3002,O_3003,O_3004,O_3005,O_3006,O_3007,O_3008,O_3009,O_3010,O_3011,O_3012,O_3013,O_3014,O_3015,O_3016,O_3017,O_3018,O_3019,O_3020,O_3021,O_3022,O_3023,O_3024,O_3025,O_3026,O_3027,O_3028,O_3029,O_3030,O_3031,O_3032,O_3033,O_3034,O_3035,O_3036,O_3037,O_3038,O_3039,O_3040,O_3041,O_3042,O_3043,O_3044,O_3045,O_3046,O_3047,O_3048,O_3049,O_3050,O_3051,O_3052,O_3053,O_3054,O_3055,O_3056,O_3057,O_3058,O_3059,O_3060,O_3061,O_3062,O_3063,O_3064,O_3065,O_3066,O_3067,O_3068,O_3069,O_3070,O_3071,O_3072,O_3073,O_3074,O_3075,O_3076,O_3077,O_3078,O_3079,O_3080,O_3081,O_3082,O_3083,O_3084,O_3085,O_3086,O_3087,O_3088,O_3089,O_3090,O_3091,O_3092,O_3093,O_3094,O_3095,O_3096,O_3097,O_3098,O_3099,O_3100,O_3101,O_3102,O_3103,O_3104,O_3105,O_3106,O_3107,O_3108,O_3109,O_3110,O_3111,O_3112,O_3113,O_3114,O_3115,O_3116,O_3117,O_3118,O_3119,O_3120,O_3121,O_3122,O_3123,O_3124,O_3125,O_3126,O_3127,O_3128,O_3129,O_3130,O_3131,O_3132,O_3133,O_3134,O_3135,O_3136,O_3137,O_3138,O_3139,O_3140,O_3141,O_3142,O_3143,O_3144,O_3145,O_3146,O_3147,O_3148,O_3149,O_3150,O_3151,O_3152,O_3153,O_3154,O_3155,O_3156,O_3157,O_3158,O_3159,O_3160,O_3161,O_3162,O_3163,O_3164,O_3165,O_3166,O_3167,O_3168,O_3169,O_3170,O_3171,O_3172,O_3173,O_3174,O_3175,O_3176,O_3177,O_3178,O_3179,O_3180,O_3181,O_3182,O_3183,O_3184,O_3185,O_3186,O_3187,O_3188,O_3189,O_3190,O_3191,O_3192,O_3193,O_3194,O_3195,O_3196,O_3197,O_3198,O_3199,O_3200,O_3201,O_3202,O_3203,O_3204,O_3205,O_3206,O_3207,O_3208,O_3209,O_3210,O_3211,O_3212,O_3213,O_3214,O_3215,O_3216,O_3217,O_3218,O_3219,O_3220,O_3221,O_3222,O_3223,O_3224,O_3225,O_3226,O_3227,O_3228,O_3229,O_3230,O_3231,O_3232,O_3233,O_3234,O_3235,O_3236,O_3237,O_3238,O_3239,O_3240,O_3241,O_3242,O_3243,O_3244,O_3245,O_3246,O_3247,O_3248,O_3249,O_3250,O_3251,O_3252,O_3253,O_3254,O_3255,O_3256,O_3257,O_3258,O_3259,O_3260,O_3261,O_3262,O_3263,O_3264,O_3265,O_3266,O_3267,O_3268,O_3269,O_3270,O_3271,O_3272,O_3273,O_3274,O_3275,O_3276,O_3277,O_3278,O_3279,O_3280,O_3281,O_3282,O_3283,O_3284,O_3285,O_3286,O_3287,O_3288,O_3289,O_3290,O_3291,O_3292,O_3293,O_3294,O_3295,O_3296,O_3297,O_3298,O_3299,O_3300,O_3301,O_3302,O_3303,O_3304,O_3305,O_3306,O_3307,O_3308,O_3309,O_3310,O_3311,O_3312,O_3313,O_3314,O_3315,O_3316,O_3317,O_3318,O_3319,O_3320,O_3321,O_3322,O_3323,O_3324,O_3325,O_3326,O_3327,O_3328,O_3329,O_3330,O_3331,O_3332,O_3333,O_3334,O_3335,O_3336,O_3337,O_3338,O_3339,O_3340,O_3341,O_3342,O_3343,O_3344,O_3345,O_3346,O_3347,O_3348,O_3349,O_3350,O_3351,O_3352,O_3353,O_3354,O_3355,O_3356,O_3357,O_3358,O_3359,O_3360,O_3361,O_3362,O_3363,O_3364,O_3365,O_3366,O_3367,O_3368,O_3369,O_3370,O_3371,O_3372,O_3373,O_3374,O_3375,O_3376,O_3377,O_3378,O_3379,O_3380,O_3381,O_3382,O_3383,O_3384,O_3385,O_3386,O_3387,O_3388,O_3389,O_3390,O_3391,O_3392,O_3393,O_3394,O_3395,O_3396,O_3397,O_3398,O_3399,O_3400,O_3401,O_3402,O_3403,O_3404,O_3405,O_3406,O_3407,O_3408,O_3409,O_3410,O_3411,O_3412,O_3413,O_3414,O_3415,O_3416,O_3417,O_3418,O_3419,O_3420,O_3421,O_3422,O_3423,O_3424,O_3425,O_3426,O_3427,O_3428,O_3429,O_3430,O_3431,O_3432,O_3433,O_3434,O_3435,O_3436,O_3437,O_3438,O_3439,O_3440,O_3441,O_3442,O_3443,O_3444,O_3445,O_3446,O_3447,O_3448,O_3449,O_3450,O_3451,O_3452,O_3453,O_3454,O_3455,O_3456,O_3457,O_3458,O_3459,O_3460,O_3461,O_3462,O_3463,O_3464,O_3465,O_3466,O_3467,O_3468,O_3469,O_3470,O_3471,O_3472,O_3473,O_3474,O_3475,O_3476,O_3477,O_3478,O_3479,O_3480,O_3481,O_3482,O_3483,O_3484,O_3485,O_3486,O_3487,O_3488,O_3489,O_3490,O_3491,O_3492,O_3493,O_3494,O_3495,O_3496,O_3497,O_3498,O_3499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999,N_25000,N_25001,N_25002,N_25003,N_25004,N_25005,N_25006,N_25007,N_25008,N_25009,N_25010,N_25011,N_25012,N_25013,N_25014,N_25015,N_25016,N_25017,N_25018,N_25019,N_25020,N_25021,N_25022,N_25023,N_25024,N_25025,N_25026,N_25027,N_25028,N_25029,N_25030,N_25031,N_25032,N_25033,N_25034,N_25035,N_25036,N_25037,N_25038,N_25039,N_25040,N_25041,N_25042,N_25043,N_25044,N_25045,N_25046,N_25047,N_25048,N_25049,N_25050,N_25051,N_25052,N_25053,N_25054,N_25055,N_25056,N_25057,N_25058,N_25059,N_25060,N_25061,N_25062,N_25063,N_25064,N_25065,N_25066,N_25067,N_25068,N_25069,N_25070,N_25071,N_25072,N_25073,N_25074,N_25075,N_25076,N_25077,N_25078,N_25079,N_25080,N_25081,N_25082,N_25083,N_25084,N_25085,N_25086,N_25087,N_25088,N_25089,N_25090,N_25091,N_25092,N_25093,N_25094,N_25095,N_25096,N_25097,N_25098,N_25099,N_25100,N_25101,N_25102,N_25103,N_25104,N_25105,N_25106,N_25107,N_25108,N_25109,N_25110,N_25111,N_25112,N_25113,N_25114,N_25115,N_25116,N_25117,N_25118,N_25119,N_25120,N_25121,N_25122,N_25123,N_25124,N_25125,N_25126,N_25127,N_25128,N_25129,N_25130,N_25131,N_25132,N_25133,N_25134,N_25135,N_25136,N_25137,N_25138,N_25139,N_25140,N_25141,N_25142,N_25143,N_25144,N_25145,N_25146,N_25147,N_25148,N_25149,N_25150,N_25151,N_25152,N_25153,N_25154,N_25155,N_25156,N_25157,N_25158,N_25159,N_25160,N_25161,N_25162,N_25163,N_25164,N_25165,N_25166,N_25167,N_25168,N_25169,N_25170,N_25171,N_25172,N_25173,N_25174,N_25175,N_25176,N_25177,N_25178,N_25179,N_25180,N_25181,N_25182,N_25183,N_25184,N_25185,N_25186,N_25187,N_25188,N_25189,N_25190,N_25191,N_25192,N_25193,N_25194,N_25195,N_25196,N_25197,N_25198,N_25199,N_25200,N_25201,N_25202,N_25203,N_25204,N_25205,N_25206,N_25207,N_25208,N_25209,N_25210,N_25211,N_25212,N_25213,N_25214,N_25215,N_25216,N_25217,N_25218,N_25219,N_25220,N_25221,N_25222,N_25223,N_25224,N_25225,N_25226,N_25227,N_25228,N_25229,N_25230,N_25231,N_25232,N_25233,N_25234,N_25235,N_25236,N_25237,N_25238,N_25239,N_25240,N_25241,N_25242,N_25243,N_25244,N_25245,N_25246,N_25247,N_25248,N_25249,N_25250,N_25251,N_25252,N_25253,N_25254,N_25255,N_25256,N_25257,N_25258,N_25259,N_25260,N_25261,N_25262,N_25263,N_25264,N_25265,N_25266,N_25267,N_25268,N_25269,N_25270,N_25271,N_25272,N_25273,N_25274,N_25275,N_25276,N_25277,N_25278,N_25279,N_25280,N_25281,N_25282,N_25283,N_25284,N_25285,N_25286,N_25287,N_25288,N_25289,N_25290,N_25291,N_25292,N_25293,N_25294,N_25295,N_25296,N_25297,N_25298,N_25299,N_25300,N_25301,N_25302,N_25303,N_25304,N_25305,N_25306,N_25307,N_25308,N_25309,N_25310,N_25311,N_25312,N_25313,N_25314,N_25315,N_25316,N_25317,N_25318,N_25319,N_25320,N_25321,N_25322,N_25323,N_25324,N_25325,N_25326,N_25327,N_25328,N_25329,N_25330,N_25331,N_25332,N_25333,N_25334,N_25335,N_25336,N_25337,N_25338,N_25339,N_25340,N_25341,N_25342,N_25343,N_25344,N_25345,N_25346,N_25347,N_25348,N_25349,N_25350,N_25351,N_25352,N_25353,N_25354,N_25355,N_25356,N_25357,N_25358,N_25359,N_25360,N_25361,N_25362,N_25363,N_25364,N_25365,N_25366,N_25367,N_25368,N_25369,N_25370,N_25371,N_25372,N_25373,N_25374,N_25375,N_25376,N_25377,N_25378,N_25379,N_25380,N_25381,N_25382,N_25383,N_25384,N_25385,N_25386,N_25387,N_25388,N_25389,N_25390,N_25391,N_25392,N_25393,N_25394,N_25395,N_25396,N_25397,N_25398,N_25399,N_25400,N_25401,N_25402,N_25403,N_25404,N_25405,N_25406,N_25407,N_25408,N_25409,N_25410,N_25411,N_25412,N_25413,N_25414,N_25415,N_25416,N_25417,N_25418,N_25419,N_25420,N_25421,N_25422,N_25423,N_25424,N_25425,N_25426,N_25427,N_25428,N_25429,N_25430,N_25431,N_25432,N_25433,N_25434,N_25435,N_25436,N_25437,N_25438,N_25439,N_25440,N_25441,N_25442,N_25443,N_25444,N_25445,N_25446,N_25447,N_25448,N_25449,N_25450,N_25451,N_25452,N_25453,N_25454,N_25455,N_25456,N_25457,N_25458,N_25459,N_25460,N_25461,N_25462,N_25463,N_25464,N_25465,N_25466,N_25467,N_25468,N_25469,N_25470,N_25471,N_25472,N_25473,N_25474,N_25475,N_25476,N_25477,N_25478,N_25479,N_25480,N_25481,N_25482,N_25483,N_25484,N_25485,N_25486,N_25487,N_25488,N_25489,N_25490,N_25491,N_25492,N_25493,N_25494,N_25495,N_25496,N_25497,N_25498,N_25499,N_25500,N_25501,N_25502,N_25503,N_25504,N_25505,N_25506,N_25507,N_25508,N_25509,N_25510,N_25511,N_25512,N_25513,N_25514,N_25515,N_25516,N_25517,N_25518,N_25519,N_25520,N_25521,N_25522,N_25523,N_25524,N_25525,N_25526,N_25527,N_25528,N_25529,N_25530,N_25531,N_25532,N_25533,N_25534,N_25535,N_25536,N_25537,N_25538,N_25539,N_25540,N_25541,N_25542,N_25543,N_25544,N_25545,N_25546,N_25547,N_25548,N_25549,N_25550,N_25551,N_25552,N_25553,N_25554,N_25555,N_25556,N_25557,N_25558,N_25559,N_25560,N_25561,N_25562,N_25563,N_25564,N_25565,N_25566,N_25567,N_25568,N_25569,N_25570,N_25571,N_25572,N_25573,N_25574,N_25575,N_25576,N_25577,N_25578,N_25579,N_25580,N_25581,N_25582,N_25583,N_25584,N_25585,N_25586,N_25587,N_25588,N_25589,N_25590,N_25591,N_25592,N_25593,N_25594,N_25595,N_25596,N_25597,N_25598,N_25599,N_25600,N_25601,N_25602,N_25603,N_25604,N_25605,N_25606,N_25607,N_25608,N_25609,N_25610,N_25611,N_25612,N_25613,N_25614,N_25615,N_25616,N_25617,N_25618,N_25619,N_25620,N_25621,N_25622,N_25623,N_25624,N_25625,N_25626,N_25627,N_25628,N_25629,N_25630,N_25631,N_25632,N_25633,N_25634,N_25635,N_25636,N_25637,N_25638,N_25639,N_25640,N_25641,N_25642,N_25643,N_25644,N_25645,N_25646,N_25647,N_25648,N_25649,N_25650,N_25651,N_25652,N_25653,N_25654,N_25655,N_25656,N_25657,N_25658,N_25659,N_25660,N_25661,N_25662,N_25663,N_25664,N_25665,N_25666,N_25667,N_25668,N_25669,N_25670,N_25671,N_25672,N_25673,N_25674,N_25675,N_25676,N_25677,N_25678,N_25679,N_25680,N_25681,N_25682,N_25683,N_25684,N_25685,N_25686,N_25687,N_25688,N_25689,N_25690,N_25691,N_25692,N_25693,N_25694,N_25695,N_25696,N_25697,N_25698,N_25699,N_25700,N_25701,N_25702,N_25703,N_25704,N_25705,N_25706,N_25707,N_25708,N_25709,N_25710,N_25711,N_25712,N_25713,N_25714,N_25715,N_25716,N_25717,N_25718,N_25719,N_25720,N_25721,N_25722,N_25723,N_25724,N_25725,N_25726,N_25727,N_25728,N_25729,N_25730,N_25731,N_25732,N_25733,N_25734,N_25735,N_25736,N_25737,N_25738,N_25739,N_25740,N_25741,N_25742,N_25743,N_25744,N_25745,N_25746,N_25747,N_25748,N_25749,N_25750,N_25751,N_25752,N_25753,N_25754,N_25755,N_25756,N_25757,N_25758,N_25759,N_25760,N_25761,N_25762,N_25763,N_25764,N_25765,N_25766,N_25767,N_25768,N_25769,N_25770,N_25771,N_25772,N_25773,N_25774,N_25775,N_25776,N_25777,N_25778,N_25779,N_25780,N_25781,N_25782,N_25783,N_25784,N_25785,N_25786,N_25787,N_25788,N_25789,N_25790,N_25791,N_25792,N_25793,N_25794,N_25795,N_25796,N_25797,N_25798,N_25799,N_25800,N_25801,N_25802,N_25803,N_25804,N_25805,N_25806,N_25807,N_25808,N_25809,N_25810,N_25811,N_25812,N_25813,N_25814,N_25815,N_25816,N_25817,N_25818,N_25819,N_25820,N_25821,N_25822,N_25823,N_25824,N_25825,N_25826,N_25827,N_25828,N_25829,N_25830,N_25831,N_25832,N_25833,N_25834,N_25835,N_25836,N_25837,N_25838,N_25839,N_25840,N_25841,N_25842,N_25843,N_25844,N_25845,N_25846,N_25847,N_25848,N_25849,N_25850,N_25851,N_25852,N_25853,N_25854,N_25855,N_25856,N_25857,N_25858,N_25859,N_25860,N_25861,N_25862,N_25863,N_25864,N_25865,N_25866,N_25867,N_25868,N_25869,N_25870,N_25871,N_25872,N_25873,N_25874,N_25875,N_25876,N_25877,N_25878,N_25879,N_25880,N_25881,N_25882,N_25883,N_25884,N_25885,N_25886,N_25887,N_25888,N_25889,N_25890,N_25891,N_25892,N_25893,N_25894,N_25895,N_25896,N_25897,N_25898,N_25899,N_25900,N_25901,N_25902,N_25903,N_25904,N_25905,N_25906,N_25907,N_25908,N_25909,N_25910,N_25911,N_25912,N_25913,N_25914,N_25915,N_25916,N_25917,N_25918,N_25919,N_25920,N_25921,N_25922,N_25923,N_25924,N_25925,N_25926,N_25927,N_25928,N_25929,N_25930,N_25931,N_25932,N_25933,N_25934,N_25935,N_25936,N_25937,N_25938,N_25939,N_25940,N_25941,N_25942,N_25943,N_25944,N_25945,N_25946,N_25947,N_25948,N_25949,N_25950,N_25951,N_25952,N_25953,N_25954,N_25955,N_25956,N_25957,N_25958,N_25959,N_25960,N_25961,N_25962,N_25963,N_25964,N_25965,N_25966,N_25967,N_25968,N_25969,N_25970,N_25971,N_25972,N_25973,N_25974,N_25975,N_25976,N_25977,N_25978,N_25979,N_25980,N_25981,N_25982,N_25983,N_25984,N_25985,N_25986,N_25987,N_25988,N_25989,N_25990,N_25991,N_25992,N_25993,N_25994,N_25995,N_25996,N_25997,N_25998,N_25999,N_26000,N_26001,N_26002,N_26003,N_26004,N_26005,N_26006,N_26007,N_26008,N_26009,N_26010,N_26011,N_26012,N_26013,N_26014,N_26015,N_26016,N_26017,N_26018,N_26019,N_26020,N_26021,N_26022,N_26023,N_26024,N_26025,N_26026,N_26027,N_26028,N_26029,N_26030,N_26031,N_26032,N_26033,N_26034,N_26035,N_26036,N_26037,N_26038,N_26039,N_26040,N_26041,N_26042,N_26043,N_26044,N_26045,N_26046,N_26047,N_26048,N_26049,N_26050,N_26051,N_26052,N_26053,N_26054,N_26055,N_26056,N_26057,N_26058,N_26059,N_26060,N_26061,N_26062,N_26063,N_26064,N_26065,N_26066,N_26067,N_26068,N_26069,N_26070,N_26071,N_26072,N_26073,N_26074,N_26075,N_26076,N_26077,N_26078,N_26079,N_26080,N_26081,N_26082,N_26083,N_26084,N_26085,N_26086,N_26087,N_26088,N_26089,N_26090,N_26091,N_26092,N_26093,N_26094,N_26095,N_26096,N_26097,N_26098,N_26099,N_26100,N_26101,N_26102,N_26103,N_26104,N_26105,N_26106,N_26107,N_26108,N_26109,N_26110,N_26111,N_26112,N_26113,N_26114,N_26115,N_26116,N_26117,N_26118,N_26119,N_26120,N_26121,N_26122,N_26123,N_26124,N_26125,N_26126,N_26127,N_26128,N_26129,N_26130,N_26131,N_26132,N_26133,N_26134,N_26135,N_26136,N_26137,N_26138,N_26139,N_26140,N_26141,N_26142,N_26143,N_26144,N_26145,N_26146,N_26147,N_26148,N_26149,N_26150,N_26151,N_26152,N_26153,N_26154,N_26155,N_26156,N_26157,N_26158,N_26159,N_26160,N_26161,N_26162,N_26163,N_26164,N_26165,N_26166,N_26167,N_26168,N_26169,N_26170,N_26171,N_26172,N_26173,N_26174,N_26175,N_26176,N_26177,N_26178,N_26179,N_26180,N_26181,N_26182,N_26183,N_26184,N_26185,N_26186,N_26187,N_26188,N_26189,N_26190,N_26191,N_26192,N_26193,N_26194,N_26195,N_26196,N_26197,N_26198,N_26199,N_26200,N_26201,N_26202,N_26203,N_26204,N_26205,N_26206,N_26207,N_26208,N_26209,N_26210,N_26211,N_26212,N_26213,N_26214,N_26215,N_26216,N_26217,N_26218,N_26219,N_26220,N_26221,N_26222,N_26223,N_26224,N_26225,N_26226,N_26227,N_26228,N_26229,N_26230,N_26231,N_26232,N_26233,N_26234,N_26235,N_26236,N_26237,N_26238,N_26239,N_26240,N_26241,N_26242,N_26243,N_26244,N_26245,N_26246,N_26247,N_26248,N_26249,N_26250,N_26251,N_26252,N_26253,N_26254,N_26255,N_26256,N_26257,N_26258,N_26259,N_26260,N_26261,N_26262,N_26263,N_26264,N_26265,N_26266,N_26267,N_26268,N_26269,N_26270,N_26271,N_26272,N_26273,N_26274,N_26275,N_26276,N_26277,N_26278,N_26279,N_26280,N_26281,N_26282,N_26283,N_26284,N_26285,N_26286,N_26287,N_26288,N_26289,N_26290,N_26291,N_26292,N_26293,N_26294,N_26295,N_26296,N_26297,N_26298,N_26299,N_26300,N_26301,N_26302,N_26303,N_26304,N_26305,N_26306,N_26307,N_26308,N_26309,N_26310,N_26311,N_26312,N_26313,N_26314,N_26315,N_26316,N_26317,N_26318,N_26319,N_26320,N_26321,N_26322,N_26323,N_26324,N_26325,N_26326,N_26327,N_26328,N_26329,N_26330,N_26331,N_26332,N_26333,N_26334,N_26335,N_26336,N_26337,N_26338,N_26339,N_26340,N_26341,N_26342,N_26343,N_26344,N_26345,N_26346,N_26347,N_26348,N_26349,N_26350,N_26351,N_26352,N_26353,N_26354,N_26355,N_26356,N_26357,N_26358,N_26359,N_26360,N_26361,N_26362,N_26363,N_26364,N_26365,N_26366,N_26367,N_26368,N_26369,N_26370,N_26371,N_26372,N_26373,N_26374,N_26375,N_26376,N_26377,N_26378,N_26379,N_26380,N_26381,N_26382,N_26383,N_26384,N_26385,N_26386,N_26387,N_26388,N_26389,N_26390,N_26391,N_26392,N_26393,N_26394,N_26395,N_26396,N_26397,N_26398,N_26399,N_26400,N_26401,N_26402,N_26403,N_26404,N_26405,N_26406,N_26407,N_26408,N_26409,N_26410,N_26411,N_26412,N_26413,N_26414,N_26415,N_26416,N_26417,N_26418,N_26419,N_26420,N_26421,N_26422,N_26423,N_26424,N_26425,N_26426,N_26427,N_26428,N_26429,N_26430,N_26431,N_26432,N_26433,N_26434,N_26435,N_26436,N_26437,N_26438,N_26439,N_26440,N_26441,N_26442,N_26443,N_26444,N_26445,N_26446,N_26447,N_26448,N_26449,N_26450,N_26451,N_26452,N_26453,N_26454,N_26455,N_26456,N_26457,N_26458,N_26459,N_26460,N_26461,N_26462,N_26463,N_26464,N_26465,N_26466,N_26467,N_26468,N_26469,N_26470,N_26471,N_26472,N_26473,N_26474,N_26475,N_26476,N_26477,N_26478,N_26479,N_26480,N_26481,N_26482,N_26483,N_26484,N_26485,N_26486,N_26487,N_26488,N_26489,N_26490,N_26491,N_26492,N_26493,N_26494,N_26495,N_26496,N_26497,N_26498,N_26499,N_26500,N_26501,N_26502,N_26503,N_26504,N_26505,N_26506,N_26507,N_26508,N_26509,N_26510,N_26511,N_26512,N_26513,N_26514,N_26515,N_26516,N_26517,N_26518,N_26519,N_26520,N_26521,N_26522,N_26523,N_26524,N_26525,N_26526,N_26527,N_26528,N_26529,N_26530,N_26531,N_26532,N_26533,N_26534,N_26535,N_26536,N_26537,N_26538,N_26539,N_26540,N_26541,N_26542,N_26543,N_26544,N_26545,N_26546,N_26547,N_26548,N_26549,N_26550,N_26551,N_26552,N_26553,N_26554,N_26555,N_26556,N_26557,N_26558,N_26559,N_26560,N_26561,N_26562,N_26563,N_26564,N_26565,N_26566,N_26567,N_26568,N_26569,N_26570,N_26571,N_26572,N_26573,N_26574,N_26575,N_26576,N_26577,N_26578,N_26579,N_26580,N_26581,N_26582,N_26583,N_26584,N_26585,N_26586,N_26587,N_26588,N_26589,N_26590,N_26591,N_26592,N_26593,N_26594,N_26595,N_26596,N_26597,N_26598,N_26599,N_26600,N_26601,N_26602,N_26603,N_26604,N_26605,N_26606,N_26607,N_26608,N_26609,N_26610,N_26611,N_26612,N_26613,N_26614,N_26615,N_26616,N_26617,N_26618,N_26619,N_26620,N_26621,N_26622,N_26623,N_26624,N_26625,N_26626,N_26627,N_26628,N_26629,N_26630,N_26631,N_26632,N_26633,N_26634,N_26635,N_26636,N_26637,N_26638,N_26639,N_26640,N_26641,N_26642,N_26643,N_26644,N_26645,N_26646,N_26647,N_26648,N_26649,N_26650,N_26651,N_26652,N_26653,N_26654,N_26655,N_26656,N_26657,N_26658,N_26659,N_26660,N_26661,N_26662,N_26663,N_26664,N_26665,N_26666,N_26667,N_26668,N_26669,N_26670,N_26671,N_26672,N_26673,N_26674,N_26675,N_26676,N_26677,N_26678,N_26679,N_26680,N_26681,N_26682,N_26683,N_26684,N_26685,N_26686,N_26687,N_26688,N_26689,N_26690,N_26691,N_26692,N_26693,N_26694,N_26695,N_26696,N_26697,N_26698,N_26699,N_26700,N_26701,N_26702,N_26703,N_26704,N_26705,N_26706,N_26707,N_26708,N_26709,N_26710,N_26711,N_26712,N_26713,N_26714,N_26715,N_26716,N_26717,N_26718,N_26719,N_26720,N_26721,N_26722,N_26723,N_26724,N_26725,N_26726,N_26727,N_26728,N_26729,N_26730,N_26731,N_26732,N_26733,N_26734,N_26735,N_26736,N_26737,N_26738,N_26739,N_26740,N_26741,N_26742,N_26743,N_26744,N_26745,N_26746,N_26747,N_26748,N_26749,N_26750,N_26751,N_26752,N_26753,N_26754,N_26755,N_26756,N_26757,N_26758,N_26759,N_26760,N_26761,N_26762,N_26763,N_26764,N_26765,N_26766,N_26767,N_26768,N_26769,N_26770,N_26771,N_26772,N_26773,N_26774,N_26775,N_26776,N_26777,N_26778,N_26779,N_26780,N_26781,N_26782,N_26783,N_26784,N_26785,N_26786,N_26787,N_26788,N_26789,N_26790,N_26791,N_26792,N_26793,N_26794,N_26795,N_26796,N_26797,N_26798,N_26799,N_26800,N_26801,N_26802,N_26803,N_26804,N_26805,N_26806,N_26807,N_26808,N_26809,N_26810,N_26811,N_26812,N_26813,N_26814,N_26815,N_26816,N_26817,N_26818,N_26819,N_26820,N_26821,N_26822,N_26823,N_26824,N_26825,N_26826,N_26827,N_26828,N_26829,N_26830,N_26831,N_26832,N_26833,N_26834,N_26835,N_26836,N_26837,N_26838,N_26839,N_26840,N_26841,N_26842,N_26843,N_26844,N_26845,N_26846,N_26847,N_26848,N_26849,N_26850,N_26851,N_26852,N_26853,N_26854,N_26855,N_26856,N_26857,N_26858,N_26859,N_26860,N_26861,N_26862,N_26863,N_26864,N_26865,N_26866,N_26867,N_26868,N_26869,N_26870,N_26871,N_26872,N_26873,N_26874,N_26875,N_26876,N_26877,N_26878,N_26879,N_26880,N_26881,N_26882,N_26883,N_26884,N_26885,N_26886,N_26887,N_26888,N_26889,N_26890,N_26891,N_26892,N_26893,N_26894,N_26895,N_26896,N_26897,N_26898,N_26899,N_26900,N_26901,N_26902,N_26903,N_26904,N_26905,N_26906,N_26907,N_26908,N_26909,N_26910,N_26911,N_26912,N_26913,N_26914,N_26915,N_26916,N_26917,N_26918,N_26919,N_26920,N_26921,N_26922,N_26923,N_26924,N_26925,N_26926,N_26927,N_26928,N_26929,N_26930,N_26931,N_26932,N_26933,N_26934,N_26935,N_26936,N_26937,N_26938,N_26939,N_26940,N_26941,N_26942,N_26943,N_26944,N_26945,N_26946,N_26947,N_26948,N_26949,N_26950,N_26951,N_26952,N_26953,N_26954,N_26955,N_26956,N_26957,N_26958,N_26959,N_26960,N_26961,N_26962,N_26963,N_26964,N_26965,N_26966,N_26967,N_26968,N_26969,N_26970,N_26971,N_26972,N_26973,N_26974,N_26975,N_26976,N_26977,N_26978,N_26979,N_26980,N_26981,N_26982,N_26983,N_26984,N_26985,N_26986,N_26987,N_26988,N_26989,N_26990,N_26991,N_26992,N_26993,N_26994,N_26995,N_26996,N_26997,N_26998,N_26999,N_27000,N_27001,N_27002,N_27003,N_27004,N_27005,N_27006,N_27007,N_27008,N_27009,N_27010,N_27011,N_27012,N_27013,N_27014,N_27015,N_27016,N_27017,N_27018,N_27019,N_27020,N_27021,N_27022,N_27023,N_27024,N_27025,N_27026,N_27027,N_27028,N_27029,N_27030,N_27031,N_27032,N_27033,N_27034,N_27035,N_27036,N_27037,N_27038,N_27039,N_27040,N_27041,N_27042,N_27043,N_27044,N_27045,N_27046,N_27047,N_27048,N_27049,N_27050,N_27051,N_27052,N_27053,N_27054,N_27055,N_27056,N_27057,N_27058,N_27059,N_27060,N_27061,N_27062,N_27063,N_27064,N_27065,N_27066,N_27067,N_27068,N_27069,N_27070,N_27071,N_27072,N_27073,N_27074,N_27075,N_27076,N_27077,N_27078,N_27079,N_27080,N_27081,N_27082,N_27083,N_27084,N_27085,N_27086,N_27087,N_27088,N_27089,N_27090,N_27091,N_27092,N_27093,N_27094,N_27095,N_27096,N_27097,N_27098,N_27099,N_27100,N_27101,N_27102,N_27103,N_27104,N_27105,N_27106,N_27107,N_27108,N_27109,N_27110,N_27111,N_27112,N_27113,N_27114,N_27115,N_27116,N_27117,N_27118,N_27119,N_27120,N_27121,N_27122,N_27123,N_27124,N_27125,N_27126,N_27127,N_27128,N_27129,N_27130,N_27131,N_27132,N_27133,N_27134,N_27135,N_27136,N_27137,N_27138,N_27139,N_27140,N_27141,N_27142,N_27143,N_27144,N_27145,N_27146,N_27147,N_27148,N_27149,N_27150,N_27151,N_27152,N_27153,N_27154,N_27155,N_27156,N_27157,N_27158,N_27159,N_27160,N_27161,N_27162,N_27163,N_27164,N_27165,N_27166,N_27167,N_27168,N_27169,N_27170,N_27171,N_27172,N_27173,N_27174,N_27175,N_27176,N_27177,N_27178,N_27179,N_27180,N_27181,N_27182,N_27183,N_27184,N_27185,N_27186,N_27187,N_27188,N_27189,N_27190,N_27191,N_27192,N_27193,N_27194,N_27195,N_27196,N_27197,N_27198,N_27199,N_27200,N_27201,N_27202,N_27203,N_27204,N_27205,N_27206,N_27207,N_27208,N_27209,N_27210,N_27211,N_27212,N_27213,N_27214,N_27215,N_27216,N_27217,N_27218,N_27219,N_27220,N_27221,N_27222,N_27223,N_27224,N_27225,N_27226,N_27227,N_27228,N_27229,N_27230,N_27231,N_27232,N_27233,N_27234,N_27235,N_27236,N_27237,N_27238,N_27239,N_27240,N_27241,N_27242,N_27243,N_27244,N_27245,N_27246,N_27247,N_27248,N_27249,N_27250,N_27251,N_27252,N_27253,N_27254,N_27255,N_27256,N_27257,N_27258,N_27259,N_27260,N_27261,N_27262,N_27263,N_27264,N_27265,N_27266,N_27267,N_27268,N_27269,N_27270,N_27271,N_27272,N_27273,N_27274,N_27275,N_27276,N_27277,N_27278,N_27279,N_27280,N_27281,N_27282,N_27283,N_27284,N_27285,N_27286,N_27287,N_27288,N_27289,N_27290,N_27291,N_27292,N_27293,N_27294,N_27295,N_27296,N_27297,N_27298,N_27299,N_27300,N_27301,N_27302,N_27303,N_27304,N_27305,N_27306,N_27307,N_27308,N_27309,N_27310,N_27311,N_27312,N_27313,N_27314,N_27315,N_27316,N_27317,N_27318,N_27319,N_27320,N_27321,N_27322,N_27323,N_27324,N_27325,N_27326,N_27327,N_27328,N_27329,N_27330,N_27331,N_27332,N_27333,N_27334,N_27335,N_27336,N_27337,N_27338,N_27339,N_27340,N_27341,N_27342,N_27343,N_27344,N_27345,N_27346,N_27347,N_27348,N_27349,N_27350,N_27351,N_27352,N_27353,N_27354,N_27355,N_27356,N_27357,N_27358,N_27359,N_27360,N_27361,N_27362,N_27363,N_27364,N_27365,N_27366,N_27367,N_27368,N_27369,N_27370,N_27371,N_27372,N_27373,N_27374,N_27375,N_27376,N_27377,N_27378,N_27379,N_27380,N_27381,N_27382,N_27383,N_27384,N_27385,N_27386,N_27387,N_27388,N_27389,N_27390,N_27391,N_27392,N_27393,N_27394,N_27395,N_27396,N_27397,N_27398,N_27399,N_27400,N_27401,N_27402,N_27403,N_27404,N_27405,N_27406,N_27407,N_27408,N_27409,N_27410,N_27411,N_27412,N_27413,N_27414,N_27415,N_27416,N_27417,N_27418,N_27419,N_27420,N_27421,N_27422,N_27423,N_27424,N_27425,N_27426,N_27427,N_27428,N_27429,N_27430,N_27431,N_27432,N_27433,N_27434,N_27435,N_27436,N_27437,N_27438,N_27439,N_27440,N_27441,N_27442,N_27443,N_27444,N_27445,N_27446,N_27447,N_27448,N_27449,N_27450,N_27451,N_27452,N_27453,N_27454,N_27455,N_27456,N_27457,N_27458,N_27459,N_27460,N_27461,N_27462,N_27463,N_27464,N_27465,N_27466,N_27467,N_27468,N_27469,N_27470,N_27471,N_27472,N_27473,N_27474,N_27475,N_27476,N_27477,N_27478,N_27479,N_27480,N_27481,N_27482,N_27483,N_27484,N_27485,N_27486,N_27487,N_27488,N_27489,N_27490,N_27491,N_27492,N_27493,N_27494,N_27495,N_27496,N_27497,N_27498,N_27499,N_27500,N_27501,N_27502,N_27503,N_27504,N_27505,N_27506,N_27507,N_27508,N_27509,N_27510,N_27511,N_27512,N_27513,N_27514,N_27515,N_27516,N_27517,N_27518,N_27519,N_27520,N_27521,N_27522,N_27523,N_27524,N_27525,N_27526,N_27527,N_27528,N_27529,N_27530,N_27531,N_27532,N_27533,N_27534,N_27535,N_27536,N_27537,N_27538,N_27539,N_27540,N_27541,N_27542,N_27543,N_27544,N_27545,N_27546,N_27547,N_27548,N_27549,N_27550,N_27551,N_27552,N_27553,N_27554,N_27555,N_27556,N_27557,N_27558,N_27559,N_27560,N_27561,N_27562,N_27563,N_27564,N_27565,N_27566,N_27567,N_27568,N_27569,N_27570,N_27571,N_27572,N_27573,N_27574,N_27575,N_27576,N_27577,N_27578,N_27579,N_27580,N_27581,N_27582,N_27583,N_27584,N_27585,N_27586,N_27587,N_27588,N_27589,N_27590,N_27591,N_27592,N_27593,N_27594,N_27595,N_27596,N_27597,N_27598,N_27599,N_27600,N_27601,N_27602,N_27603,N_27604,N_27605,N_27606,N_27607,N_27608,N_27609,N_27610,N_27611,N_27612,N_27613,N_27614,N_27615,N_27616,N_27617,N_27618,N_27619,N_27620,N_27621,N_27622,N_27623,N_27624,N_27625,N_27626,N_27627,N_27628,N_27629,N_27630,N_27631,N_27632,N_27633,N_27634,N_27635,N_27636,N_27637,N_27638,N_27639,N_27640,N_27641,N_27642,N_27643,N_27644,N_27645,N_27646,N_27647,N_27648,N_27649,N_27650,N_27651,N_27652,N_27653,N_27654,N_27655,N_27656,N_27657,N_27658,N_27659,N_27660,N_27661,N_27662,N_27663,N_27664,N_27665,N_27666,N_27667,N_27668,N_27669,N_27670,N_27671,N_27672,N_27673,N_27674,N_27675,N_27676,N_27677,N_27678,N_27679,N_27680,N_27681,N_27682,N_27683,N_27684,N_27685,N_27686,N_27687,N_27688,N_27689,N_27690,N_27691,N_27692,N_27693,N_27694,N_27695,N_27696,N_27697,N_27698,N_27699,N_27700,N_27701,N_27702,N_27703,N_27704,N_27705,N_27706,N_27707,N_27708,N_27709,N_27710,N_27711,N_27712,N_27713,N_27714,N_27715,N_27716,N_27717,N_27718,N_27719,N_27720,N_27721,N_27722,N_27723,N_27724,N_27725,N_27726,N_27727,N_27728,N_27729,N_27730,N_27731,N_27732,N_27733,N_27734,N_27735,N_27736,N_27737,N_27738,N_27739,N_27740,N_27741,N_27742,N_27743,N_27744,N_27745,N_27746,N_27747,N_27748,N_27749,N_27750,N_27751,N_27752,N_27753,N_27754,N_27755,N_27756,N_27757,N_27758,N_27759,N_27760,N_27761,N_27762,N_27763,N_27764,N_27765,N_27766,N_27767,N_27768,N_27769,N_27770,N_27771,N_27772,N_27773,N_27774,N_27775,N_27776,N_27777,N_27778,N_27779,N_27780,N_27781,N_27782,N_27783,N_27784,N_27785,N_27786,N_27787,N_27788,N_27789,N_27790,N_27791,N_27792,N_27793,N_27794,N_27795,N_27796,N_27797,N_27798,N_27799,N_27800,N_27801,N_27802,N_27803,N_27804,N_27805,N_27806,N_27807,N_27808,N_27809,N_27810,N_27811,N_27812,N_27813,N_27814,N_27815,N_27816,N_27817,N_27818,N_27819,N_27820,N_27821,N_27822,N_27823,N_27824,N_27825,N_27826,N_27827,N_27828,N_27829,N_27830,N_27831,N_27832,N_27833,N_27834,N_27835,N_27836,N_27837,N_27838,N_27839,N_27840,N_27841,N_27842,N_27843,N_27844,N_27845,N_27846,N_27847,N_27848,N_27849,N_27850,N_27851,N_27852,N_27853,N_27854,N_27855,N_27856,N_27857,N_27858,N_27859,N_27860,N_27861,N_27862,N_27863,N_27864,N_27865,N_27866,N_27867,N_27868,N_27869,N_27870,N_27871,N_27872,N_27873,N_27874,N_27875,N_27876,N_27877,N_27878,N_27879,N_27880,N_27881,N_27882,N_27883,N_27884,N_27885,N_27886,N_27887,N_27888,N_27889,N_27890,N_27891,N_27892,N_27893,N_27894,N_27895,N_27896,N_27897,N_27898,N_27899,N_27900,N_27901,N_27902,N_27903,N_27904,N_27905,N_27906,N_27907,N_27908,N_27909,N_27910,N_27911,N_27912,N_27913,N_27914,N_27915,N_27916,N_27917,N_27918,N_27919,N_27920,N_27921,N_27922,N_27923,N_27924,N_27925,N_27926,N_27927,N_27928,N_27929,N_27930,N_27931,N_27932,N_27933,N_27934,N_27935,N_27936,N_27937,N_27938,N_27939,N_27940,N_27941,N_27942,N_27943,N_27944,N_27945,N_27946,N_27947,N_27948,N_27949,N_27950,N_27951,N_27952,N_27953,N_27954,N_27955,N_27956,N_27957,N_27958,N_27959,N_27960,N_27961,N_27962,N_27963,N_27964,N_27965,N_27966,N_27967,N_27968,N_27969,N_27970,N_27971,N_27972,N_27973,N_27974,N_27975,N_27976,N_27977,N_27978,N_27979,N_27980,N_27981,N_27982,N_27983,N_27984,N_27985,N_27986,N_27987,N_27988,N_27989,N_27990,N_27991,N_27992,N_27993,N_27994,N_27995,N_27996,N_27997,N_27998,N_27999,N_28000,N_28001,N_28002,N_28003,N_28004,N_28005,N_28006,N_28007,N_28008,N_28009,N_28010,N_28011,N_28012,N_28013,N_28014,N_28015,N_28016,N_28017,N_28018,N_28019,N_28020,N_28021,N_28022,N_28023,N_28024,N_28025,N_28026,N_28027,N_28028,N_28029,N_28030,N_28031,N_28032,N_28033,N_28034,N_28035,N_28036,N_28037,N_28038,N_28039,N_28040,N_28041,N_28042,N_28043,N_28044,N_28045,N_28046,N_28047,N_28048,N_28049,N_28050,N_28051,N_28052,N_28053,N_28054,N_28055,N_28056,N_28057,N_28058,N_28059,N_28060,N_28061,N_28062,N_28063,N_28064,N_28065,N_28066,N_28067,N_28068,N_28069,N_28070,N_28071,N_28072,N_28073,N_28074,N_28075,N_28076,N_28077,N_28078,N_28079,N_28080,N_28081,N_28082,N_28083,N_28084,N_28085,N_28086,N_28087,N_28088,N_28089,N_28090,N_28091,N_28092,N_28093,N_28094,N_28095,N_28096,N_28097,N_28098,N_28099,N_28100,N_28101,N_28102,N_28103,N_28104,N_28105,N_28106,N_28107,N_28108,N_28109,N_28110,N_28111,N_28112,N_28113,N_28114,N_28115,N_28116,N_28117,N_28118,N_28119,N_28120,N_28121,N_28122,N_28123,N_28124,N_28125,N_28126,N_28127,N_28128,N_28129,N_28130,N_28131,N_28132,N_28133,N_28134,N_28135,N_28136,N_28137,N_28138,N_28139,N_28140,N_28141,N_28142,N_28143,N_28144,N_28145,N_28146,N_28147,N_28148,N_28149,N_28150,N_28151,N_28152,N_28153,N_28154,N_28155,N_28156,N_28157,N_28158,N_28159,N_28160,N_28161,N_28162,N_28163,N_28164,N_28165,N_28166,N_28167,N_28168,N_28169,N_28170,N_28171,N_28172,N_28173,N_28174,N_28175,N_28176,N_28177,N_28178,N_28179,N_28180,N_28181,N_28182,N_28183,N_28184,N_28185,N_28186,N_28187,N_28188,N_28189,N_28190,N_28191,N_28192,N_28193,N_28194,N_28195,N_28196,N_28197,N_28198,N_28199,N_28200,N_28201,N_28202,N_28203,N_28204,N_28205,N_28206,N_28207,N_28208,N_28209,N_28210,N_28211,N_28212,N_28213,N_28214,N_28215,N_28216,N_28217,N_28218,N_28219,N_28220,N_28221,N_28222,N_28223,N_28224,N_28225,N_28226,N_28227,N_28228,N_28229,N_28230,N_28231,N_28232,N_28233,N_28234,N_28235,N_28236,N_28237,N_28238,N_28239,N_28240,N_28241,N_28242,N_28243,N_28244,N_28245,N_28246,N_28247,N_28248,N_28249,N_28250,N_28251,N_28252,N_28253,N_28254,N_28255,N_28256,N_28257,N_28258,N_28259,N_28260,N_28261,N_28262,N_28263,N_28264,N_28265,N_28266,N_28267,N_28268,N_28269,N_28270,N_28271,N_28272,N_28273,N_28274,N_28275,N_28276,N_28277,N_28278,N_28279,N_28280,N_28281,N_28282,N_28283,N_28284,N_28285,N_28286,N_28287,N_28288,N_28289,N_28290,N_28291,N_28292,N_28293,N_28294,N_28295,N_28296,N_28297,N_28298,N_28299,N_28300,N_28301,N_28302,N_28303,N_28304,N_28305,N_28306,N_28307,N_28308,N_28309,N_28310,N_28311,N_28312,N_28313,N_28314,N_28315,N_28316,N_28317,N_28318,N_28319,N_28320,N_28321,N_28322,N_28323,N_28324,N_28325,N_28326,N_28327,N_28328,N_28329,N_28330,N_28331,N_28332,N_28333,N_28334,N_28335,N_28336,N_28337,N_28338,N_28339,N_28340,N_28341,N_28342,N_28343,N_28344,N_28345,N_28346,N_28347,N_28348,N_28349,N_28350,N_28351,N_28352,N_28353,N_28354,N_28355,N_28356,N_28357,N_28358,N_28359,N_28360,N_28361,N_28362,N_28363,N_28364,N_28365,N_28366,N_28367,N_28368,N_28369,N_28370,N_28371,N_28372,N_28373,N_28374,N_28375,N_28376,N_28377,N_28378,N_28379,N_28380,N_28381,N_28382,N_28383,N_28384,N_28385,N_28386,N_28387,N_28388,N_28389,N_28390,N_28391,N_28392,N_28393,N_28394,N_28395,N_28396,N_28397,N_28398,N_28399,N_28400,N_28401,N_28402,N_28403,N_28404,N_28405,N_28406,N_28407,N_28408,N_28409,N_28410,N_28411,N_28412,N_28413,N_28414,N_28415,N_28416,N_28417,N_28418,N_28419,N_28420,N_28421,N_28422,N_28423,N_28424,N_28425,N_28426,N_28427,N_28428,N_28429,N_28430,N_28431,N_28432,N_28433,N_28434,N_28435,N_28436,N_28437,N_28438,N_28439,N_28440,N_28441,N_28442,N_28443,N_28444,N_28445,N_28446,N_28447,N_28448,N_28449,N_28450,N_28451,N_28452,N_28453,N_28454,N_28455,N_28456,N_28457,N_28458,N_28459,N_28460,N_28461,N_28462,N_28463,N_28464,N_28465,N_28466,N_28467,N_28468,N_28469,N_28470,N_28471,N_28472,N_28473,N_28474,N_28475,N_28476,N_28477,N_28478,N_28479,N_28480,N_28481,N_28482,N_28483,N_28484,N_28485,N_28486,N_28487,N_28488,N_28489,N_28490,N_28491,N_28492,N_28493,N_28494,N_28495,N_28496,N_28497,N_28498,N_28499,N_28500,N_28501,N_28502,N_28503,N_28504,N_28505,N_28506,N_28507,N_28508,N_28509,N_28510,N_28511,N_28512,N_28513,N_28514,N_28515,N_28516,N_28517,N_28518,N_28519,N_28520,N_28521,N_28522,N_28523,N_28524,N_28525,N_28526,N_28527,N_28528,N_28529,N_28530,N_28531,N_28532,N_28533,N_28534,N_28535,N_28536,N_28537,N_28538,N_28539,N_28540,N_28541,N_28542,N_28543,N_28544,N_28545,N_28546,N_28547,N_28548,N_28549,N_28550,N_28551,N_28552,N_28553,N_28554,N_28555,N_28556,N_28557,N_28558,N_28559,N_28560,N_28561,N_28562,N_28563,N_28564,N_28565,N_28566,N_28567,N_28568,N_28569,N_28570,N_28571,N_28572,N_28573,N_28574,N_28575,N_28576,N_28577,N_28578,N_28579,N_28580,N_28581,N_28582,N_28583,N_28584,N_28585,N_28586,N_28587,N_28588,N_28589,N_28590,N_28591,N_28592,N_28593,N_28594,N_28595,N_28596,N_28597,N_28598,N_28599,N_28600,N_28601,N_28602,N_28603,N_28604,N_28605,N_28606,N_28607,N_28608,N_28609,N_28610,N_28611,N_28612,N_28613,N_28614,N_28615,N_28616,N_28617,N_28618,N_28619,N_28620,N_28621,N_28622,N_28623,N_28624,N_28625,N_28626,N_28627,N_28628,N_28629,N_28630,N_28631,N_28632,N_28633,N_28634,N_28635,N_28636,N_28637,N_28638,N_28639,N_28640,N_28641,N_28642,N_28643,N_28644,N_28645,N_28646,N_28647,N_28648,N_28649,N_28650,N_28651,N_28652,N_28653,N_28654,N_28655,N_28656,N_28657,N_28658,N_28659,N_28660,N_28661,N_28662,N_28663,N_28664,N_28665,N_28666,N_28667,N_28668,N_28669,N_28670,N_28671,N_28672,N_28673,N_28674,N_28675,N_28676,N_28677,N_28678,N_28679,N_28680,N_28681,N_28682,N_28683,N_28684,N_28685,N_28686,N_28687,N_28688,N_28689,N_28690,N_28691,N_28692,N_28693,N_28694,N_28695,N_28696,N_28697,N_28698,N_28699,N_28700,N_28701,N_28702,N_28703,N_28704,N_28705,N_28706,N_28707,N_28708,N_28709,N_28710,N_28711,N_28712,N_28713,N_28714,N_28715,N_28716,N_28717,N_28718,N_28719,N_28720,N_28721,N_28722,N_28723,N_28724,N_28725,N_28726,N_28727,N_28728,N_28729,N_28730,N_28731,N_28732,N_28733,N_28734,N_28735,N_28736,N_28737,N_28738,N_28739,N_28740,N_28741,N_28742,N_28743,N_28744,N_28745,N_28746,N_28747,N_28748,N_28749,N_28750,N_28751,N_28752,N_28753,N_28754,N_28755,N_28756,N_28757,N_28758,N_28759,N_28760,N_28761,N_28762,N_28763,N_28764,N_28765,N_28766,N_28767,N_28768,N_28769,N_28770,N_28771,N_28772,N_28773,N_28774,N_28775,N_28776,N_28777,N_28778,N_28779,N_28780,N_28781,N_28782,N_28783,N_28784,N_28785,N_28786,N_28787,N_28788,N_28789,N_28790,N_28791,N_28792,N_28793,N_28794,N_28795,N_28796,N_28797,N_28798,N_28799,N_28800,N_28801,N_28802,N_28803,N_28804,N_28805,N_28806,N_28807,N_28808,N_28809,N_28810,N_28811,N_28812,N_28813,N_28814,N_28815,N_28816,N_28817,N_28818,N_28819,N_28820,N_28821,N_28822,N_28823,N_28824,N_28825,N_28826,N_28827,N_28828,N_28829,N_28830,N_28831,N_28832,N_28833,N_28834,N_28835,N_28836,N_28837,N_28838,N_28839,N_28840,N_28841,N_28842,N_28843,N_28844,N_28845,N_28846,N_28847,N_28848,N_28849,N_28850,N_28851,N_28852,N_28853,N_28854,N_28855,N_28856,N_28857,N_28858,N_28859,N_28860,N_28861,N_28862,N_28863,N_28864,N_28865,N_28866,N_28867,N_28868,N_28869,N_28870,N_28871,N_28872,N_28873,N_28874,N_28875,N_28876,N_28877,N_28878,N_28879,N_28880,N_28881,N_28882,N_28883,N_28884,N_28885,N_28886,N_28887,N_28888,N_28889,N_28890,N_28891,N_28892,N_28893,N_28894,N_28895,N_28896,N_28897,N_28898,N_28899,N_28900,N_28901,N_28902,N_28903,N_28904,N_28905,N_28906,N_28907,N_28908,N_28909,N_28910,N_28911,N_28912,N_28913,N_28914,N_28915,N_28916,N_28917,N_28918,N_28919,N_28920,N_28921,N_28922,N_28923,N_28924,N_28925,N_28926,N_28927,N_28928,N_28929,N_28930,N_28931,N_28932,N_28933,N_28934,N_28935,N_28936,N_28937,N_28938,N_28939,N_28940,N_28941,N_28942,N_28943,N_28944,N_28945,N_28946,N_28947,N_28948,N_28949,N_28950,N_28951,N_28952,N_28953,N_28954,N_28955,N_28956,N_28957,N_28958,N_28959,N_28960,N_28961,N_28962,N_28963,N_28964,N_28965,N_28966,N_28967,N_28968,N_28969,N_28970,N_28971,N_28972,N_28973,N_28974,N_28975,N_28976,N_28977,N_28978,N_28979,N_28980,N_28981,N_28982,N_28983,N_28984,N_28985,N_28986,N_28987,N_28988,N_28989,N_28990,N_28991,N_28992,N_28993,N_28994,N_28995,N_28996,N_28997,N_28998,N_28999,N_29000,N_29001,N_29002,N_29003,N_29004,N_29005,N_29006,N_29007,N_29008,N_29009,N_29010,N_29011,N_29012,N_29013,N_29014,N_29015,N_29016,N_29017,N_29018,N_29019,N_29020,N_29021,N_29022,N_29023,N_29024,N_29025,N_29026,N_29027,N_29028,N_29029,N_29030,N_29031,N_29032,N_29033,N_29034,N_29035,N_29036,N_29037,N_29038,N_29039,N_29040,N_29041,N_29042,N_29043,N_29044,N_29045,N_29046,N_29047,N_29048,N_29049,N_29050,N_29051,N_29052,N_29053,N_29054,N_29055,N_29056,N_29057,N_29058,N_29059,N_29060,N_29061,N_29062,N_29063,N_29064,N_29065,N_29066,N_29067,N_29068,N_29069,N_29070,N_29071,N_29072,N_29073,N_29074,N_29075,N_29076,N_29077,N_29078,N_29079,N_29080,N_29081,N_29082,N_29083,N_29084,N_29085,N_29086,N_29087,N_29088,N_29089,N_29090,N_29091,N_29092,N_29093,N_29094,N_29095,N_29096,N_29097,N_29098,N_29099,N_29100,N_29101,N_29102,N_29103,N_29104,N_29105,N_29106,N_29107,N_29108,N_29109,N_29110,N_29111,N_29112,N_29113,N_29114,N_29115,N_29116,N_29117,N_29118,N_29119,N_29120,N_29121,N_29122,N_29123,N_29124,N_29125,N_29126,N_29127,N_29128,N_29129,N_29130,N_29131,N_29132,N_29133,N_29134,N_29135,N_29136,N_29137,N_29138,N_29139,N_29140,N_29141,N_29142,N_29143,N_29144,N_29145,N_29146,N_29147,N_29148,N_29149,N_29150,N_29151,N_29152,N_29153,N_29154,N_29155,N_29156,N_29157,N_29158,N_29159,N_29160,N_29161,N_29162,N_29163,N_29164,N_29165,N_29166,N_29167,N_29168,N_29169,N_29170,N_29171,N_29172,N_29173,N_29174,N_29175,N_29176,N_29177,N_29178,N_29179,N_29180,N_29181,N_29182,N_29183,N_29184,N_29185,N_29186,N_29187,N_29188,N_29189,N_29190,N_29191,N_29192,N_29193,N_29194,N_29195,N_29196,N_29197,N_29198,N_29199,N_29200,N_29201,N_29202,N_29203,N_29204,N_29205,N_29206,N_29207,N_29208,N_29209,N_29210,N_29211,N_29212,N_29213,N_29214,N_29215,N_29216,N_29217,N_29218,N_29219,N_29220,N_29221,N_29222,N_29223,N_29224,N_29225,N_29226,N_29227,N_29228,N_29229,N_29230,N_29231,N_29232,N_29233,N_29234,N_29235,N_29236,N_29237,N_29238,N_29239,N_29240,N_29241,N_29242,N_29243,N_29244,N_29245,N_29246,N_29247,N_29248,N_29249,N_29250,N_29251,N_29252,N_29253,N_29254,N_29255,N_29256,N_29257,N_29258,N_29259,N_29260,N_29261,N_29262,N_29263,N_29264,N_29265,N_29266,N_29267,N_29268,N_29269,N_29270,N_29271,N_29272,N_29273,N_29274,N_29275,N_29276,N_29277,N_29278,N_29279,N_29280,N_29281,N_29282,N_29283,N_29284,N_29285,N_29286,N_29287,N_29288,N_29289,N_29290,N_29291,N_29292,N_29293,N_29294,N_29295,N_29296,N_29297,N_29298,N_29299,N_29300,N_29301,N_29302,N_29303,N_29304,N_29305,N_29306,N_29307,N_29308,N_29309,N_29310,N_29311,N_29312,N_29313,N_29314,N_29315,N_29316,N_29317,N_29318,N_29319,N_29320,N_29321,N_29322,N_29323,N_29324,N_29325,N_29326,N_29327,N_29328,N_29329,N_29330,N_29331,N_29332,N_29333,N_29334,N_29335,N_29336,N_29337,N_29338,N_29339,N_29340,N_29341,N_29342,N_29343,N_29344,N_29345,N_29346,N_29347,N_29348,N_29349,N_29350,N_29351,N_29352,N_29353,N_29354,N_29355,N_29356,N_29357,N_29358,N_29359,N_29360,N_29361,N_29362,N_29363,N_29364,N_29365,N_29366,N_29367,N_29368,N_29369,N_29370,N_29371,N_29372,N_29373,N_29374,N_29375,N_29376,N_29377,N_29378,N_29379,N_29380,N_29381,N_29382,N_29383,N_29384,N_29385,N_29386,N_29387,N_29388,N_29389,N_29390,N_29391,N_29392,N_29393,N_29394,N_29395,N_29396,N_29397,N_29398,N_29399,N_29400,N_29401,N_29402,N_29403,N_29404,N_29405,N_29406,N_29407,N_29408,N_29409,N_29410,N_29411,N_29412,N_29413,N_29414,N_29415,N_29416,N_29417,N_29418,N_29419,N_29420,N_29421,N_29422,N_29423,N_29424,N_29425,N_29426,N_29427,N_29428,N_29429,N_29430,N_29431,N_29432,N_29433,N_29434,N_29435,N_29436,N_29437,N_29438,N_29439,N_29440,N_29441,N_29442,N_29443,N_29444,N_29445,N_29446,N_29447,N_29448,N_29449,N_29450,N_29451,N_29452,N_29453,N_29454,N_29455,N_29456,N_29457,N_29458,N_29459,N_29460,N_29461,N_29462,N_29463,N_29464,N_29465,N_29466,N_29467,N_29468,N_29469,N_29470,N_29471,N_29472,N_29473,N_29474,N_29475,N_29476,N_29477,N_29478,N_29479,N_29480,N_29481,N_29482,N_29483,N_29484,N_29485,N_29486,N_29487,N_29488,N_29489,N_29490,N_29491,N_29492,N_29493,N_29494,N_29495,N_29496,N_29497,N_29498,N_29499,N_29500,N_29501,N_29502,N_29503,N_29504,N_29505,N_29506,N_29507,N_29508,N_29509,N_29510,N_29511,N_29512,N_29513,N_29514,N_29515,N_29516,N_29517,N_29518,N_29519,N_29520,N_29521,N_29522,N_29523,N_29524,N_29525,N_29526,N_29527,N_29528,N_29529,N_29530,N_29531,N_29532,N_29533,N_29534,N_29535,N_29536,N_29537,N_29538,N_29539,N_29540,N_29541,N_29542,N_29543,N_29544,N_29545,N_29546,N_29547,N_29548,N_29549,N_29550,N_29551,N_29552,N_29553,N_29554,N_29555,N_29556,N_29557,N_29558,N_29559,N_29560,N_29561,N_29562,N_29563,N_29564,N_29565,N_29566,N_29567,N_29568,N_29569,N_29570,N_29571,N_29572,N_29573,N_29574,N_29575,N_29576,N_29577,N_29578,N_29579,N_29580,N_29581,N_29582,N_29583,N_29584,N_29585,N_29586,N_29587,N_29588,N_29589,N_29590,N_29591,N_29592,N_29593,N_29594,N_29595,N_29596,N_29597,N_29598,N_29599,N_29600,N_29601,N_29602,N_29603,N_29604,N_29605,N_29606,N_29607,N_29608,N_29609,N_29610,N_29611,N_29612,N_29613,N_29614,N_29615,N_29616,N_29617,N_29618,N_29619,N_29620,N_29621,N_29622,N_29623,N_29624,N_29625,N_29626,N_29627,N_29628,N_29629,N_29630,N_29631,N_29632,N_29633,N_29634,N_29635,N_29636,N_29637,N_29638,N_29639,N_29640,N_29641,N_29642,N_29643,N_29644,N_29645,N_29646,N_29647,N_29648,N_29649,N_29650,N_29651,N_29652,N_29653,N_29654,N_29655,N_29656,N_29657,N_29658,N_29659,N_29660,N_29661,N_29662,N_29663,N_29664,N_29665,N_29666,N_29667,N_29668,N_29669,N_29670,N_29671,N_29672,N_29673,N_29674,N_29675,N_29676,N_29677,N_29678,N_29679,N_29680,N_29681,N_29682,N_29683,N_29684,N_29685,N_29686,N_29687,N_29688,N_29689,N_29690,N_29691,N_29692,N_29693,N_29694,N_29695,N_29696,N_29697,N_29698,N_29699,N_29700,N_29701,N_29702,N_29703,N_29704,N_29705,N_29706,N_29707,N_29708,N_29709,N_29710,N_29711,N_29712,N_29713,N_29714,N_29715,N_29716,N_29717,N_29718,N_29719,N_29720,N_29721,N_29722,N_29723,N_29724,N_29725,N_29726,N_29727,N_29728,N_29729,N_29730,N_29731,N_29732,N_29733,N_29734,N_29735,N_29736,N_29737,N_29738,N_29739,N_29740,N_29741,N_29742,N_29743,N_29744,N_29745,N_29746,N_29747,N_29748,N_29749,N_29750,N_29751,N_29752,N_29753,N_29754,N_29755,N_29756,N_29757,N_29758,N_29759,N_29760,N_29761,N_29762,N_29763,N_29764,N_29765,N_29766,N_29767,N_29768,N_29769,N_29770,N_29771,N_29772,N_29773,N_29774,N_29775,N_29776,N_29777,N_29778,N_29779,N_29780,N_29781,N_29782,N_29783,N_29784,N_29785,N_29786,N_29787,N_29788,N_29789,N_29790,N_29791,N_29792,N_29793,N_29794,N_29795,N_29796,N_29797,N_29798,N_29799,N_29800,N_29801,N_29802,N_29803,N_29804,N_29805,N_29806,N_29807,N_29808,N_29809,N_29810,N_29811,N_29812,N_29813,N_29814,N_29815,N_29816,N_29817,N_29818,N_29819,N_29820,N_29821,N_29822,N_29823,N_29824,N_29825,N_29826,N_29827,N_29828,N_29829,N_29830,N_29831,N_29832,N_29833,N_29834,N_29835,N_29836,N_29837,N_29838,N_29839,N_29840,N_29841,N_29842,N_29843,N_29844,N_29845,N_29846,N_29847,N_29848,N_29849,N_29850,N_29851,N_29852,N_29853,N_29854,N_29855,N_29856,N_29857,N_29858,N_29859,N_29860,N_29861,N_29862,N_29863,N_29864,N_29865,N_29866,N_29867,N_29868,N_29869,N_29870,N_29871,N_29872,N_29873,N_29874,N_29875,N_29876,N_29877,N_29878,N_29879,N_29880,N_29881,N_29882,N_29883,N_29884,N_29885,N_29886,N_29887,N_29888,N_29889,N_29890,N_29891,N_29892,N_29893,N_29894,N_29895,N_29896,N_29897,N_29898,N_29899,N_29900,N_29901,N_29902,N_29903,N_29904,N_29905,N_29906,N_29907,N_29908,N_29909,N_29910,N_29911,N_29912,N_29913,N_29914,N_29915,N_29916,N_29917,N_29918,N_29919,N_29920,N_29921,N_29922,N_29923,N_29924,N_29925,N_29926,N_29927,N_29928,N_29929,N_29930,N_29931,N_29932,N_29933,N_29934,N_29935,N_29936,N_29937,N_29938,N_29939,N_29940,N_29941,N_29942,N_29943,N_29944,N_29945,N_29946,N_29947,N_29948,N_29949,N_29950,N_29951,N_29952,N_29953,N_29954,N_29955,N_29956,N_29957,N_29958,N_29959,N_29960,N_29961,N_29962,N_29963,N_29964,N_29965,N_29966,N_29967,N_29968,N_29969,N_29970,N_29971,N_29972,N_29973,N_29974,N_29975,N_29976,N_29977,N_29978,N_29979,N_29980,N_29981,N_29982,N_29983,N_29984,N_29985,N_29986,N_29987,N_29988,N_29989,N_29990,N_29991,N_29992,N_29993,N_29994,N_29995,N_29996,N_29997,N_29998,N_29999;
nand U0 (N_0,In_2538,In_636);
nand U1 (N_1,In_2510,In_1922);
nand U2 (N_2,In_1698,In_2294);
nand U3 (N_3,In_1444,In_517);
nand U4 (N_4,In_2689,In_358);
or U5 (N_5,In_304,In_2898);
nor U6 (N_6,In_2785,In_1527);
or U7 (N_7,In_1531,In_738);
or U8 (N_8,In_2399,In_2152);
nand U9 (N_9,In_364,In_1462);
or U10 (N_10,In_2605,In_1009);
or U11 (N_11,In_331,In_2729);
nand U12 (N_12,In_2226,In_1979);
and U13 (N_13,In_1608,In_2723);
nand U14 (N_14,In_203,In_491);
nand U15 (N_15,In_2883,In_2179);
and U16 (N_16,In_2449,In_693);
nor U17 (N_17,In_2156,In_2951);
and U18 (N_18,In_2186,In_702);
nor U19 (N_19,In_1692,In_819);
nand U20 (N_20,In_1162,In_2523);
nor U21 (N_21,In_2329,In_1606);
xnor U22 (N_22,In_2699,In_1533);
or U23 (N_23,In_1559,In_1025);
nand U24 (N_24,In_804,In_589);
and U25 (N_25,In_412,In_809);
xor U26 (N_26,In_2344,In_882);
xor U27 (N_27,In_1006,In_1223);
and U28 (N_28,In_110,In_284);
or U29 (N_29,In_2199,In_330);
or U30 (N_30,In_1784,In_236);
nand U31 (N_31,In_0,In_1643);
or U32 (N_32,In_265,In_934);
and U33 (N_33,In_2066,In_2210);
nor U34 (N_34,In_211,In_274);
nand U35 (N_35,In_313,In_1656);
and U36 (N_36,In_896,In_1385);
nand U37 (N_37,In_2998,In_82);
and U38 (N_38,In_1196,In_1911);
and U39 (N_39,In_878,In_642);
nand U40 (N_40,In_891,In_2583);
and U41 (N_41,In_2021,In_272);
nand U42 (N_42,In_1891,In_1779);
or U43 (N_43,In_724,In_2823);
or U44 (N_44,In_1284,In_2556);
nor U45 (N_45,In_1239,In_1429);
nor U46 (N_46,In_2459,In_250);
and U47 (N_47,In_1893,In_2901);
and U48 (N_48,In_2767,In_1279);
or U49 (N_49,In_2805,In_2351);
and U50 (N_50,In_670,In_575);
xor U51 (N_51,In_437,In_1603);
and U52 (N_52,In_200,In_1085);
or U53 (N_53,In_239,In_1122);
or U54 (N_54,In_1616,In_2920);
nand U55 (N_55,In_2558,In_2637);
and U56 (N_56,In_1637,In_1056);
or U57 (N_57,In_1282,In_661);
and U58 (N_58,In_205,In_1325);
or U59 (N_59,In_1872,In_801);
or U60 (N_60,In_1370,In_2600);
or U61 (N_61,In_2890,In_2650);
nor U62 (N_62,In_1959,In_944);
nor U63 (N_63,In_8,In_548);
nor U64 (N_64,In_1316,In_768);
nor U65 (N_65,In_2803,In_1622);
nor U66 (N_66,In_543,In_1428);
nand U67 (N_67,In_1189,In_1881);
and U68 (N_68,In_1151,In_2345);
nand U69 (N_69,In_1393,In_354);
nor U70 (N_70,In_753,In_2029);
and U71 (N_71,In_1408,In_116);
and U72 (N_72,In_2830,In_1463);
or U73 (N_73,In_2277,In_2441);
nand U74 (N_74,In_7,In_654);
nor U75 (N_75,In_1921,In_1053);
xnor U76 (N_76,In_1237,In_521);
nand U77 (N_77,In_1937,In_1803);
or U78 (N_78,In_182,In_2978);
nand U79 (N_79,In_2014,In_1542);
and U80 (N_80,In_632,In_230);
nor U81 (N_81,In_1360,In_2771);
xor U82 (N_82,In_1406,In_903);
and U83 (N_83,In_184,In_2279);
and U84 (N_84,In_2621,In_2239);
or U85 (N_85,In_2589,In_2299);
nand U86 (N_86,In_705,In_1846);
and U87 (N_87,In_2322,In_1773);
nor U88 (N_88,In_1347,In_2659);
and U89 (N_89,In_2057,In_1045);
or U90 (N_90,In_2293,In_1657);
xor U91 (N_91,In_1743,In_1210);
and U92 (N_92,In_1432,In_746);
xor U93 (N_93,In_513,In_1211);
xor U94 (N_94,In_401,In_953);
nor U95 (N_95,In_817,In_410);
and U96 (N_96,In_2712,In_1330);
nand U97 (N_97,In_2011,In_504);
nor U98 (N_98,In_2457,In_2560);
and U99 (N_99,In_319,In_2458);
and U100 (N_100,In_2751,In_2874);
xnor U101 (N_101,In_138,In_1700);
nor U102 (N_102,In_2974,In_2539);
and U103 (N_103,In_2573,In_1195);
nand U104 (N_104,In_2330,In_2599);
or U105 (N_105,In_2914,In_787);
and U106 (N_106,In_2675,In_292);
nor U107 (N_107,In_2969,In_1276);
or U108 (N_108,In_733,In_2015);
or U109 (N_109,In_1250,In_835);
or U110 (N_110,In_2073,In_1248);
and U111 (N_111,In_385,In_811);
and U112 (N_112,In_1716,In_902);
or U113 (N_113,In_2832,In_1016);
or U114 (N_114,In_949,In_1246);
or U115 (N_115,In_1477,In_641);
or U116 (N_116,In_1355,In_1371);
and U117 (N_117,In_41,In_2690);
or U118 (N_118,In_129,In_372);
nand U119 (N_119,In_2224,In_140);
nand U120 (N_120,In_2948,In_2648);
or U121 (N_121,In_1687,In_604);
and U122 (N_122,In_554,In_2582);
nand U123 (N_123,In_1887,In_21);
or U124 (N_124,In_849,In_792);
or U125 (N_125,In_1680,In_1183);
nor U126 (N_126,In_72,In_937);
and U127 (N_127,In_1520,In_101);
or U128 (N_128,In_2045,In_1361);
and U129 (N_129,In_1058,In_1618);
nor U130 (N_130,In_1468,In_537);
nor U131 (N_131,In_1352,In_463);
xnor U132 (N_132,In_681,In_1066);
or U133 (N_133,In_2262,In_659);
nand U134 (N_134,In_244,In_2090);
and U135 (N_135,In_195,In_1132);
nor U136 (N_136,In_2320,In_545);
xnor U137 (N_137,In_2982,In_1503);
nor U138 (N_138,In_1288,In_523);
or U139 (N_139,In_749,In_2182);
and U140 (N_140,In_1178,In_2514);
or U141 (N_141,In_2851,In_1351);
and U142 (N_142,In_2203,In_1677);
or U143 (N_143,In_1167,In_1142);
nand U144 (N_144,In_452,In_2072);
and U145 (N_145,In_223,In_925);
and U146 (N_146,In_1696,In_2384);
or U147 (N_147,In_2632,In_2524);
and U148 (N_148,In_1127,In_473);
nor U149 (N_149,In_1544,In_1599);
nor U150 (N_150,In_38,In_2761);
and U151 (N_151,In_732,In_97);
and U152 (N_152,In_1720,In_1746);
or U153 (N_153,In_1648,In_422);
and U154 (N_154,In_2835,In_39);
nand U155 (N_155,In_2040,In_1731);
nor U156 (N_156,In_327,In_1146);
nor U157 (N_157,In_2430,In_119);
or U158 (N_158,In_14,In_969);
nor U159 (N_159,In_2041,In_2815);
and U160 (N_160,In_1069,In_1835);
nand U161 (N_161,In_1051,In_580);
nand U162 (N_162,In_1427,In_2779);
nor U163 (N_163,In_1868,In_566);
and U164 (N_164,In_1577,In_496);
nor U165 (N_165,In_210,In_2083);
and U166 (N_166,In_1430,In_1668);
nand U167 (N_167,In_1386,In_2472);
nand U168 (N_168,In_2502,In_451);
nand U169 (N_169,In_959,In_55);
and U170 (N_170,In_2929,In_719);
nor U171 (N_171,In_569,In_409);
nand U172 (N_172,In_2587,In_2735);
or U173 (N_173,In_1526,In_2343);
nand U174 (N_174,In_2939,In_1034);
and U175 (N_175,In_2122,In_427);
or U176 (N_176,In_865,In_1421);
and U177 (N_177,In_901,In_294);
or U178 (N_178,In_434,In_215);
or U179 (N_179,In_89,In_508);
nand U180 (N_180,In_666,In_1448);
or U181 (N_181,In_597,In_391);
and U182 (N_182,In_1861,In_2380);
nor U183 (N_183,In_947,In_2244);
nor U184 (N_184,In_1073,In_2933);
nor U185 (N_185,In_912,In_1392);
and U186 (N_186,In_181,In_1889);
nor U187 (N_187,In_593,In_83);
xnor U188 (N_188,In_1359,In_966);
or U189 (N_189,In_2130,In_759);
or U190 (N_190,In_2402,In_881);
nor U191 (N_191,In_723,In_22);
nand U192 (N_192,In_336,In_2542);
and U193 (N_193,In_850,In_1925);
nand U194 (N_194,In_216,In_2398);
nand U195 (N_195,In_1435,In_544);
nor U196 (N_196,In_2216,In_439);
xnor U197 (N_197,In_1120,In_2953);
nor U198 (N_198,In_2572,In_2428);
and U199 (N_199,In_2099,In_2371);
or U200 (N_200,In_591,In_799);
or U201 (N_201,In_1244,In_1561);
or U202 (N_202,In_2337,In_687);
nand U203 (N_203,In_596,In_2498);
xor U204 (N_204,In_2652,In_2112);
or U205 (N_205,In_1280,In_2264);
nor U206 (N_206,In_1528,In_1763);
xor U207 (N_207,In_1332,In_2468);
xnor U208 (N_208,In_1164,In_2944);
or U209 (N_209,In_1585,In_1666);
nor U210 (N_210,In_2527,In_2217);
nor U211 (N_211,In_2943,In_1032);
nand U212 (N_212,In_1958,In_567);
and U213 (N_213,In_291,In_1710);
nand U214 (N_214,In_1469,In_810);
or U215 (N_215,In_1290,In_1281);
nand U216 (N_216,In_2697,In_989);
nor U217 (N_217,In_1970,In_1856);
nand U218 (N_218,In_1240,In_1465);
nor U219 (N_219,In_2684,In_2067);
or U220 (N_220,In_2005,In_2229);
nor U221 (N_221,In_286,In_196);
and U222 (N_222,In_2742,In_1083);
and U223 (N_223,In_1335,In_188);
nand U224 (N_224,In_2155,In_2149);
and U225 (N_225,In_5,In_2038);
nor U226 (N_226,In_2205,In_1764);
xnor U227 (N_227,In_1150,In_2984);
nor U228 (N_228,In_1673,In_1342);
and U229 (N_229,In_635,In_647);
and U230 (N_230,In_1619,In_688);
xnor U231 (N_231,In_2976,In_1800);
or U232 (N_232,In_2454,In_1339);
nand U233 (N_233,In_1641,In_1317);
or U234 (N_234,In_948,In_255);
or U235 (N_235,In_2598,In_2418);
nand U236 (N_236,In_467,In_431);
and U237 (N_237,In_352,In_563);
and U238 (N_238,In_1809,In_1452);
nor U239 (N_239,In_1109,In_1285);
nand U240 (N_240,In_1836,In_2750);
nand U241 (N_241,In_1088,In_770);
or U242 (N_242,In_796,In_1484);
and U243 (N_243,In_2204,In_2999);
nand U244 (N_244,In_271,In_2247);
nand U245 (N_245,In_2195,In_2850);
nand U246 (N_246,In_1137,In_2053);
xor U247 (N_247,In_2241,In_1046);
and U248 (N_248,In_2055,In_1512);
nand U249 (N_249,In_2574,In_154);
and U250 (N_250,In_2054,In_2036);
nand U251 (N_251,In_275,In_1261);
or U252 (N_252,In_2911,In_2460);
or U253 (N_253,In_2051,In_2476);
nand U254 (N_254,In_1133,In_1569);
and U255 (N_255,In_2645,In_2717);
nand U256 (N_256,In_701,In_2087);
or U257 (N_257,In_797,In_1778);
nor U258 (N_258,In_1967,In_1909);
or U259 (N_259,In_1888,In_1047);
xnor U260 (N_260,In_2989,In_697);
and U261 (N_261,In_617,In_1214);
nand U262 (N_262,In_1838,In_213);
nor U263 (N_263,In_1257,In_1005);
and U264 (N_264,In_1262,In_333);
nor U265 (N_265,In_2421,In_1156);
nor U266 (N_266,In_2385,In_201);
nand U267 (N_267,In_1023,In_2482);
and U268 (N_268,In_1556,In_2635);
or U269 (N_269,In_24,In_1268);
and U270 (N_270,In_25,In_757);
nand U271 (N_271,In_1505,In_1108);
or U272 (N_272,In_1942,In_886);
or U273 (N_273,In_2480,In_469);
and U274 (N_274,In_2190,In_2081);
xor U275 (N_275,In_1082,In_67);
or U276 (N_276,In_1049,In_321);
and U277 (N_277,In_2,In_1830);
nor U278 (N_278,In_1334,In_374);
nand U279 (N_279,In_2870,In_2392);
nand U280 (N_280,In_1530,In_542);
or U281 (N_281,In_2726,In_2658);
or U282 (N_282,In_2420,In_2923);
and U283 (N_283,In_289,In_156);
nor U284 (N_284,In_2396,In_1772);
or U285 (N_285,In_1434,In_529);
nor U286 (N_286,In_2386,In_1617);
nand U287 (N_287,In_1078,In_587);
or U288 (N_288,In_1372,In_1848);
xnor U289 (N_289,In_2634,In_2234);
nand U290 (N_290,In_561,In_531);
xnor U291 (N_291,In_2786,In_1594);
or U292 (N_292,In_2909,In_2076);
or U293 (N_293,In_2888,In_2465);
nor U294 (N_294,In_1695,In_967);
xnor U295 (N_295,In_51,In_1795);
nand U296 (N_296,In_908,In_1808);
and U297 (N_297,In_1587,In_462);
and U298 (N_298,In_1601,In_440);
or U299 (N_299,In_1158,In_1766);
and U300 (N_300,In_836,In_2533);
xnor U301 (N_301,In_386,In_731);
and U302 (N_302,In_1501,In_1327);
nand U303 (N_303,In_955,In_803);
or U304 (N_304,In_994,In_546);
nor U305 (N_305,In_1343,In_1532);
nor U306 (N_306,In_446,In_127);
and U307 (N_307,In_2875,In_1417);
nand U308 (N_308,In_772,In_1684);
nand U309 (N_309,In_44,In_958);
and U310 (N_310,In_306,In_873);
and U311 (N_311,In_574,In_1013);
nand U312 (N_312,In_2483,In_2569);
nor U313 (N_313,In_520,In_1715);
and U314 (N_314,In_943,In_1173);
nand U315 (N_315,In_480,In_2431);
and U316 (N_316,In_2283,In_2721);
nor U317 (N_317,In_1283,In_1265);
or U318 (N_318,In_2694,In_1907);
nand U319 (N_319,In_242,In_2938);
and U320 (N_320,In_2327,In_1018);
xnor U321 (N_321,In_2397,In_2448);
and U322 (N_322,In_2926,In_2113);
or U323 (N_323,In_833,In_1381);
or U324 (N_324,In_2529,In_2893);
and U325 (N_325,In_863,In_146);
nor U326 (N_326,In_1769,In_455);
or U327 (N_327,In_1033,In_2025);
xnor U328 (N_328,In_2052,In_2173);
nand U329 (N_329,In_2764,In_2987);
and U330 (N_330,In_823,In_2627);
nor U331 (N_331,In_305,In_1117);
nor U332 (N_332,In_1377,In_1090);
nor U333 (N_333,In_2378,In_1445);
nand U334 (N_334,In_2983,In_279);
nor U335 (N_335,In_1124,In_2221);
xnor U336 (N_336,In_465,In_2592);
nand U337 (N_337,In_2143,In_2284);
or U338 (N_338,In_615,In_754);
and U339 (N_339,In_2810,In_458);
nor U340 (N_340,In_468,In_2641);
xnor U341 (N_341,In_880,In_1969);
or U342 (N_342,In_1642,In_143);
nor U343 (N_343,In_285,In_1256);
xnor U344 (N_344,In_2991,In_1638);
and U345 (N_345,In_2075,In_490);
nor U346 (N_346,In_1035,In_104);
nand U347 (N_347,In_1039,In_2278);
and U348 (N_348,In_672,In_59);
xnor U349 (N_349,In_1757,In_30);
nor U350 (N_350,In_1551,In_494);
xnor U351 (N_351,In_813,In_2417);
and U352 (N_352,In_1380,In_472);
or U353 (N_353,In_756,In_322);
xor U354 (N_354,In_2732,In_1274);
nor U355 (N_355,In_1554,In_805);
nand U356 (N_356,In_2961,In_109);
nor U357 (N_357,In_1135,In_194);
xnor U358 (N_358,In_1067,In_1492);
nand U359 (N_359,In_618,In_894);
nor U360 (N_360,In_831,In_1884);
and U361 (N_361,In_481,In_332);
nand U362 (N_362,In_640,In_2248);
nor U363 (N_363,In_235,In_560);
and U364 (N_364,In_2595,In_423);
nand U365 (N_365,In_1983,In_1115);
or U366 (N_366,In_1095,In_1971);
or U367 (N_367,In_946,In_1052);
nor U368 (N_368,In_2887,In_1728);
and U369 (N_369,In_1539,In_2528);
nand U370 (N_370,In_1043,In_1216);
nor U371 (N_371,In_1676,In_2654);
nor U372 (N_372,In_2309,In_1449);
nand U373 (N_373,In_176,In_1988);
nor U374 (N_374,In_1699,In_2114);
or U375 (N_375,In_318,In_198);
or U376 (N_376,In_1876,In_978);
xor U377 (N_377,In_2633,In_457);
and U378 (N_378,In_739,In_1304);
nor U379 (N_379,In_2972,In_1894);
xnor U380 (N_380,In_2246,In_1933);
nor U381 (N_381,In_2791,In_1790);
and U382 (N_382,In_2686,In_1770);
nand U383 (N_383,In_827,In_2968);
and U384 (N_384,In_15,In_2710);
nor U385 (N_385,In_2030,In_2773);
nand U386 (N_386,In_982,In_2936);
or U387 (N_387,In_2930,In_1995);
nor U388 (N_388,In_2058,In_820);
or U389 (N_389,In_2331,In_1549);
nand U390 (N_390,In_1962,In_2607);
nor U391 (N_391,In_565,In_2032);
nand U392 (N_392,In_2432,In_1948);
and U393 (N_393,In_362,In_1704);
or U394 (N_394,In_2367,In_2841);
nor U395 (N_395,In_418,In_920);
and U396 (N_396,In_1583,In_2154);
nor U397 (N_397,In_2222,In_17);
nand U398 (N_398,In_2346,In_2450);
xor U399 (N_399,In_2734,In_1956);
and U400 (N_400,In_161,In_2281);
xnor U401 (N_401,In_1524,In_1134);
nand U402 (N_402,In_550,In_838);
nand U403 (N_403,In_2842,In_2174);
nor U404 (N_404,In_2985,In_1661);
nor U405 (N_405,In_717,In_945);
and U406 (N_406,In_2146,In_264);
nor U407 (N_407,In_855,In_668);
nor U408 (N_408,In_611,In_2282);
xor U409 (N_409,In_1096,In_1071);
nand U410 (N_410,In_1537,In_1940);
nor U411 (N_411,In_2243,In_2877);
nand U412 (N_412,In_342,In_939);
nor U413 (N_413,In_1759,In_2772);
nand U414 (N_414,In_1788,In_2640);
nor U415 (N_415,In_940,In_35);
or U416 (N_416,In_1507,In_1890);
and U417 (N_417,In_1148,In_1785);
or U418 (N_418,In_2892,In_656);
or U419 (N_419,In_2197,In_2097);
or U420 (N_420,In_1689,In_1738);
or U421 (N_421,In_784,In_2638);
nor U422 (N_422,In_299,In_471);
nor U423 (N_423,In_2504,In_2352);
nand U424 (N_424,In_380,In_2956);
or U425 (N_425,In_2963,In_28);
or U426 (N_426,In_2389,In_445);
xor U427 (N_427,In_1841,In_1300);
and U428 (N_428,In_1,In_996);
nand U429 (N_429,In_2251,In_2446);
and U430 (N_430,In_2519,In_2618);
xor U431 (N_431,In_180,In_1560);
or U432 (N_432,In_1263,In_2272);
nor U433 (N_433,In_1411,In_2880);
nand U434 (N_434,In_33,In_229);
nor U435 (N_435,In_1225,In_2374);
nand U436 (N_436,In_1185,In_31);
nand U437 (N_437,In_2715,In_1792);
or U438 (N_438,In_2844,In_77);
or U439 (N_439,In_1076,In_1902);
or U440 (N_440,In_1114,In_1609);
nor U441 (N_441,In_2549,In_1374);
or U442 (N_442,In_2960,In_85);
and U443 (N_443,In_2702,In_157);
nor U444 (N_444,In_405,In_1513);
nand U445 (N_445,In_1605,In_2409);
nand U446 (N_446,In_1973,In_2501);
and U447 (N_447,In_64,In_2491);
and U448 (N_448,In_428,In_2092);
xnor U449 (N_449,In_1050,In_2579);
and U450 (N_450,In_2235,In_482);
and U451 (N_451,In_1141,In_2861);
nand U452 (N_452,In_136,In_1929);
nor U453 (N_453,In_432,In_1663);
and U454 (N_454,In_2670,In_2828);
or U455 (N_455,In_649,In_1777);
nand U456 (N_456,In_2082,In_875);
and U457 (N_457,In_628,In_1447);
or U458 (N_458,In_483,In_2980);
and U459 (N_459,In_56,In_2427);
nand U460 (N_460,In_2608,In_2731);
or U461 (N_461,In_413,In_2796);
and U462 (N_462,In_2564,In_2037);
and U463 (N_463,In_1844,In_144);
and U464 (N_464,In_231,In_1188);
or U465 (N_465,In_1624,In_918);
nor U466 (N_466,In_1831,In_557);
nand U467 (N_467,In_2394,In_1946);
nand U468 (N_468,In_81,In_991);
and U469 (N_469,In_1315,In_2847);
and U470 (N_470,In_479,In_1705);
or U471 (N_471,In_2077,In_1485);
nor U472 (N_472,In_303,In_500);
and U473 (N_473,In_2680,In_2230);
xnor U474 (N_474,In_2897,In_2419);
xnor U475 (N_475,In_631,In_1003);
or U476 (N_476,In_1719,In_1259);
or U477 (N_477,In_1296,In_1901);
nor U478 (N_478,In_1842,In_2370);
nor U479 (N_479,In_1102,In_2683);
nand U480 (N_480,In_478,In_2535);
and U481 (N_481,In_276,In_2471);
nand U482 (N_482,In_2907,In_2825);
or U483 (N_483,In_2563,In_2286);
or U484 (N_484,In_466,In_1388);
and U485 (N_485,In_2138,In_2981);
or U486 (N_486,In_658,In_2100);
and U487 (N_487,In_602,In_1328);
and U488 (N_488,In_526,In_1194);
nand U489 (N_489,In_206,In_745);
nor U490 (N_490,In_95,In_1002);
and U491 (N_491,In_1707,In_2121);
or U492 (N_492,In_2342,In_495);
nand U493 (N_493,In_131,In_348);
nor U494 (N_494,In_1238,In_2878);
nor U495 (N_495,In_2616,In_1936);
nor U496 (N_496,In_1456,In_842);
or U497 (N_497,In_2383,In_87);
and U498 (N_498,In_2191,In_1021);
nand U499 (N_499,In_1612,In_1660);
or U500 (N_500,In_2060,In_2140);
nand U501 (N_501,In_2782,In_2903);
nand U502 (N_502,In_2442,In_2590);
nor U503 (N_503,In_2954,In_343);
or U504 (N_504,In_2778,In_2496);
nand U505 (N_505,In_2056,In_2740);
xor U506 (N_506,In_460,In_212);
or U507 (N_507,In_1475,In_1904);
or U508 (N_508,In_191,In_1206);
or U509 (N_509,In_844,In_2148);
nor U510 (N_510,In_541,In_1235);
or U511 (N_511,In_2860,In_1479);
nand U512 (N_512,In_1140,In_2671);
or U513 (N_513,In_2361,In_1786);
and U514 (N_514,In_916,In_2720);
and U515 (N_515,In_96,In_660);
or U516 (N_516,In_2799,In_1105);
nand U517 (N_517,In_1204,In_425);
nor U518 (N_518,In_2006,In_1312);
or U519 (N_519,In_442,In_2228);
xnor U520 (N_520,In_1019,In_390);
or U521 (N_521,In_1113,In_917);
and U522 (N_522,In_287,In_2912);
xor U523 (N_523,In_1659,In_2365);
and U524 (N_524,In_2382,In_1038);
or U525 (N_525,In_990,In_629);
and U526 (N_526,In_2407,In_2678);
nor U527 (N_527,In_789,In_2376);
nor U528 (N_528,In_1991,In_1845);
and U529 (N_529,In_74,In_1678);
and U530 (N_530,In_92,In_2125);
xnor U531 (N_531,In_1251,In_2485);
xor U532 (N_532,In_1340,In_346);
or U533 (N_533,In_1324,In_2261);
or U534 (N_534,In_616,In_2128);
nand U535 (N_535,In_378,In_1546);
nand U536 (N_536,In_2604,In_2176);
xnor U537 (N_537,In_682,In_1059);
and U538 (N_538,In_2393,In_1147);
or U539 (N_539,In_760,In_1832);
nand U540 (N_540,In_2555,In_121);
or U541 (N_541,In_1871,In_115);
nand U542 (N_542,In_450,In_1100);
nor U543 (N_543,In_734,In_1801);
xor U544 (N_544,In_2922,In_2511);
nand U545 (N_545,In_1190,In_341);
or U546 (N_546,In_1927,In_10);
or U547 (N_547,In_2068,In_2647);
nand U548 (N_548,In_780,In_369);
xnor U549 (N_549,In_1226,In_2473);
xor U550 (N_550,In_869,In_2798);
or U551 (N_551,In_1636,In_726);
nand U552 (N_552,In_954,In_1664);
nand U553 (N_553,In_52,In_111);
or U554 (N_554,In_2770,In_2044);
nand U555 (N_555,In_2411,In_1741);
nand U556 (N_556,In_1266,In_159);
nand U557 (N_557,In_309,In_1511);
or U558 (N_558,In_281,In_262);
and U559 (N_559,In_1509,In_1875);
and U560 (N_560,In_2207,In_153);
nor U561 (N_561,In_2354,In_2840);
and U562 (N_562,In_2879,In_1490);
and U563 (N_563,In_1847,In_2273);
nor U564 (N_564,In_2967,In_2802);
nor U565 (N_565,In_2335,In_748);
nor U566 (N_566,In_411,In_2245);
nand U567 (N_567,In_2395,In_808);
nand U568 (N_568,In_1589,In_1683);
and U569 (N_569,In_727,In_2208);
nand U570 (N_570,In_2255,In_2001);
nand U571 (N_571,In_347,In_417);
and U572 (N_572,In_1582,In_376);
nor U573 (N_573,In_2063,In_1271);
or U574 (N_574,In_2775,In_1953);
xnor U575 (N_575,In_1717,In_2947);
nor U576 (N_576,In_1614,In_2096);
nand U577 (N_577,In_997,In_1153);
nand U578 (N_578,In_627,In_2406);
nand U579 (N_579,In_308,In_1443);
and U580 (N_580,In_2602,In_1155);
and U581 (N_581,In_1128,In_2256);
nor U582 (N_582,In_1758,In_527);
nand U583 (N_583,In_927,In_2444);
nor U584 (N_584,In_2797,In_1389);
and U585 (N_585,In_2324,In_2626);
nand U586 (N_586,In_325,In_2308);
nor U587 (N_587,In_2748,In_1394);
or U588 (N_588,In_988,In_1482);
nor U589 (N_589,In_2910,In_2267);
or U590 (N_590,In_1552,In_1525);
or U591 (N_591,In_453,In_791);
xor U592 (N_592,In_2258,In_2387);
nor U593 (N_593,In_2003,In_570);
and U594 (N_594,In_73,In_1961);
nor U595 (N_595,In_2788,In_923);
nand U596 (N_596,In_1396,In_2813);
nand U597 (N_597,In_2614,In_578);
or U598 (N_598,In_1472,In_254);
xor U599 (N_599,In_2202,In_1849);
nand U600 (N_600,In_2628,In_572);
nor U601 (N_601,N_175,In_2578);
nor U602 (N_602,In_1048,In_1807);
or U603 (N_603,In_2467,In_70);
nor U604 (N_604,In_1125,N_59);
nor U605 (N_605,In_1087,In_2749);
or U606 (N_606,In_251,In_1917);
or U607 (N_607,In_1097,In_2970);
nor U608 (N_608,N_369,N_452);
or U609 (N_609,In_2571,N_120);
or U610 (N_610,In_497,In_1375);
and U611 (N_611,N_372,In_61);
and U612 (N_612,N_385,In_365);
nor U613 (N_613,In_2091,In_665);
nand U614 (N_614,In_2843,In_2129);
and U615 (N_615,N_215,In_2804);
nand U616 (N_616,In_19,In_762);
nor U617 (N_617,In_202,In_2856);
or U618 (N_618,N_1,N_129);
nor U619 (N_619,In_2470,In_2094);
xor U620 (N_620,In_2137,In_1119);
or U621 (N_621,In_1877,N_325);
nor U622 (N_622,In_1913,In_853);
xnor U623 (N_623,In_503,In_334);
and U624 (N_624,In_1649,In_2168);
nand U625 (N_625,In_1850,In_1419);
nor U626 (N_626,In_2462,In_363);
nand U627 (N_627,N_253,In_876);
and U628 (N_628,In_1647,In_2007);
nor U629 (N_629,N_22,In_60);
nand U630 (N_630,In_1028,In_1213);
and U631 (N_631,N_92,N_183);
and U632 (N_632,In_2415,N_336);
and U633 (N_633,In_1063,In_58);
and U634 (N_634,N_460,In_783);
xnor U635 (N_635,N_159,N_445);
nor U636 (N_636,In_895,In_1821);
or U637 (N_637,In_1767,In_485);
nand U638 (N_638,In_714,In_1091);
nand U639 (N_639,In_2776,In_2611);
nor U640 (N_640,In_1960,In_1584);
nor U641 (N_641,N_164,N_565);
and U642 (N_642,In_2934,In_1407);
nor U643 (N_643,N_20,In_765);
nor U644 (N_644,N_24,In_2517);
or U645 (N_645,N_473,In_1433);
xor U646 (N_646,N_586,In_2757);
nand U647 (N_647,N_111,In_151);
xor U648 (N_648,In_1514,In_1191);
nand U649 (N_649,In_712,In_2317);
nand U650 (N_650,In_1812,N_469);
and U651 (N_651,In_169,N_553);
nor U652 (N_652,In_2362,In_634);
nor U653 (N_653,In_856,In_930);
nor U654 (N_654,In_852,In_377);
xnor U655 (N_655,In_877,N_399);
nand U656 (N_656,In_2979,In_1422);
xnor U657 (N_657,In_238,In_168);
and U658 (N_658,N_308,In_1797);
or U659 (N_659,In_1567,In_883);
and U660 (N_660,In_2711,In_2534);
and U661 (N_661,In_1177,N_515);
and U662 (N_662,N_133,In_470);
or U663 (N_663,In_2925,N_543);
and U664 (N_664,In_1476,N_488);
nor U665 (N_665,N_307,In_1234);
or U666 (N_666,In_269,In_1851);
and U667 (N_667,N_468,In_2673);
and U668 (N_668,In_2429,In_1943);
nand U669 (N_669,In_415,In_2837);
nor U670 (N_670,In_2042,In_1756);
nand U671 (N_671,In_1130,In_766);
nand U672 (N_672,In_2784,N_541);
nand U673 (N_673,N_593,In_2639);
nor U674 (N_674,N_174,In_232);
or U675 (N_675,In_1457,In_1878);
or U676 (N_676,In_2606,In_108);
or U677 (N_677,In_2185,N_427);
nand U678 (N_678,N_115,In_1968);
nor U679 (N_679,In_2369,In_2225);
or U680 (N_680,In_847,In_1706);
xor U681 (N_681,In_233,In_1358);
and U682 (N_682,In_2692,In_2755);
nor U683 (N_683,In_1761,In_2035);
nor U684 (N_684,In_691,In_2593);
nand U685 (N_685,N_118,In_2214);
nand U686 (N_686,In_737,N_52);
and U687 (N_687,In_904,In_1935);
nor U688 (N_688,In_355,In_178);
nor U689 (N_689,N_114,In_488);
nor U690 (N_690,In_1510,N_499);
nor U691 (N_691,In_1441,In_2009);
nor U692 (N_692,In_2706,In_547);
and U693 (N_693,N_524,In_1138);
nand U694 (N_694,In_2086,In_1879);
or U695 (N_695,In_2492,In_1752);
nor U696 (N_696,N_82,In_1897);
nor U697 (N_697,N_205,In_1287);
or U698 (N_698,In_2488,In_900);
nand U699 (N_699,In_1873,N_391);
and U700 (N_700,In_404,N_31);
and U701 (N_701,In_1278,In_1308);
nand U702 (N_702,In_559,In_914);
nand U703 (N_703,In_1712,N_126);
and U704 (N_704,N_132,In_1089);
nor U705 (N_705,In_135,N_416);
or U706 (N_706,In_2973,In_1912);
nand U707 (N_707,In_2777,In_773);
xor U708 (N_708,In_449,In_1610);
nand U709 (N_709,N_589,In_1024);
nand U710 (N_710,In_2158,In_2737);
or U711 (N_711,In_588,In_100);
nor U712 (N_712,In_802,In_806);
or U713 (N_713,N_513,In_1976);
or U714 (N_714,In_2131,N_122);
or U715 (N_715,In_326,N_362);
or U716 (N_716,In_1833,In_1273);
nor U717 (N_717,N_458,N_590);
and U718 (N_718,In_23,In_266);
xor U719 (N_719,In_2636,In_2059);
and U720 (N_720,In_1632,In_711);
nor U721 (N_721,In_2849,In_2661);
and U722 (N_722,In_1722,N_453);
and U723 (N_723,In_1202,In_76);
nand U724 (N_724,In_43,N_23);
nor U725 (N_725,N_236,In_57);
nand U726 (N_726,In_1607,N_10);
nand U727 (N_727,In_837,In_986);
and U728 (N_728,In_2808,In_614);
nor U729 (N_729,N_279,In_256);
or U730 (N_730,In_368,In_1802);
or U731 (N_731,N_148,In_2872);
nor U732 (N_732,In_2900,N_123);
nor U733 (N_733,In_2744,In_270);
and U734 (N_734,In_935,In_2789);
or U735 (N_735,In_1667,In_2048);
and U736 (N_736,In_828,N_125);
nor U737 (N_737,In_86,In_1571);
or U738 (N_738,In_47,In_1245);
nand U739 (N_739,In_1346,In_1523);
xor U740 (N_740,In_1305,In_2110);
and U741 (N_741,N_395,In_2400);
and U742 (N_742,In_2292,In_2852);
or U743 (N_743,N_267,N_491);
or U744 (N_744,In_843,In_2964);
or U745 (N_745,In_1197,In_539);
and U746 (N_746,In_2730,In_2913);
and U747 (N_747,In_2359,In_2466);
or U748 (N_748,In_2725,N_591);
nor U749 (N_749,N_80,In_2794);
or U750 (N_750,In_1121,In_2145);
nand U751 (N_751,In_1180,In_353);
and U752 (N_752,In_921,In_2236);
xor U753 (N_753,In_752,N_397);
and U754 (N_754,In_793,N_270);
xnor U755 (N_755,In_2642,In_938);
or U756 (N_756,In_718,In_2904);
nor U757 (N_757,In_2657,In_208);
or U758 (N_758,In_1254,In_516);
and U759 (N_759,N_273,N_562);
nor U760 (N_760,In_2372,In_535);
nor U761 (N_761,In_1776,In_1748);
nand U762 (N_762,In_394,N_190);
nand U763 (N_763,In_1502,In_1080);
xnor U764 (N_764,In_769,In_1212);
or U765 (N_765,In_2487,In_1941);
nor U766 (N_766,N_383,In_357);
and U767 (N_767,N_57,In_1401);
nand U768 (N_768,In_311,N_285);
or U769 (N_769,In_1437,In_1272);
nor U770 (N_770,In_259,N_480);
xnor U771 (N_771,In_1154,N_418);
nand U772 (N_772,N_76,N_442);
or U773 (N_773,N_360,N_559);
xnor U774 (N_774,In_2275,In_2147);
nand U775 (N_775,N_229,In_1219);
and U776 (N_776,In_2955,In_2685);
or U777 (N_777,N_45,N_588);
or U778 (N_778,N_220,N_404);
nand U779 (N_779,In_2567,In_263);
or U780 (N_780,In_320,In_2811);
or U781 (N_781,In_1857,In_2596);
or U782 (N_782,In_2624,In_2945);
and U783 (N_783,In_214,N_298);
xor U784 (N_784,In_1635,In_562);
nand U785 (N_785,In_741,In_963);
and U786 (N_786,In_2232,In_1885);
nand U787 (N_787,N_37,N_247);
and U788 (N_788,In_475,In_1275);
and U789 (N_789,In_2610,N_492);
nor U790 (N_790,In_248,In_1563);
or U791 (N_791,In_777,N_153);
and U792 (N_792,In_1628,N_545);
and U793 (N_793,In_2824,N_119);
and U794 (N_794,In_1218,In_130);
nand U795 (N_795,In_1558,In_2134);
nand U796 (N_796,In_684,In_2377);
or U797 (N_797,In_2288,N_547);
and U798 (N_798,In_2196,In_32);
nor U799 (N_799,In_370,N_531);
xor U800 (N_800,In_49,In_1198);
nand U801 (N_801,N_527,N_293);
xor U802 (N_802,In_393,In_2591);
nor U803 (N_803,In_2136,N_27);
nand U804 (N_804,N_17,In_2434);
and U805 (N_805,In_2340,In_1898);
and U806 (N_806,In_2161,N_340);
or U807 (N_807,In_1144,In_1319);
or U808 (N_808,In_1703,In_2357);
or U809 (N_809,In_2486,In_2941);
or U810 (N_810,In_273,N_314);
and U811 (N_811,N_276,In_199);
and U812 (N_812,N_415,In_858);
xor U813 (N_813,In_1007,N_328);
or U814 (N_814,In_1466,N_60);
or U815 (N_815,In_1416,In_582);
or U816 (N_816,In_932,N_333);
and U817 (N_817,In_735,N_331);
or U818 (N_818,In_794,N_529);
and U819 (N_819,In_1733,In_1924);
nand U820 (N_820,In_2391,In_1209);
and U821 (N_821,In_179,In_6);
nand U822 (N_822,In_700,In_1950);
xor U823 (N_823,In_598,In_2708);
xor U824 (N_824,In_1399,In_68);
and U825 (N_825,In_1813,In_592);
xnor U826 (N_826,In_1163,N_390);
nand U827 (N_827,In_1674,In_2806);
and U828 (N_828,In_48,In_1747);
and U829 (N_829,In_1027,N_484);
or U830 (N_830,N_568,In_2338);
nor U831 (N_831,In_209,N_112);
nor U832 (N_832,In_722,In_2325);
nor U833 (N_833,N_514,In_1574);
nor U834 (N_834,In_2756,In_2516);
xnor U835 (N_835,In_2439,In_2265);
and U836 (N_836,N_2,In_2070);
and U837 (N_837,In_1729,In_1481);
nor U838 (N_838,N_65,N_546);
nand U839 (N_839,In_1152,In_301);
nand U840 (N_840,In_1363,In_2801);
or U841 (N_841,In_771,N_187);
nor U842 (N_842,N_566,In_2000);
nand U843 (N_843,N_393,In_298);
and U844 (N_844,In_2049,In_2594);
nor U845 (N_845,In_34,In_525);
xor U846 (N_846,In_1438,In_1883);
nand U847 (N_847,In_1760,N_425);
nor U848 (N_848,In_461,In_105);
nand U849 (N_849,In_102,N_209);
nand U850 (N_850,N_58,In_980);
nand U851 (N_851,In_2445,In_859);
nand U852 (N_852,In_1103,In_1458);
or U853 (N_853,N_38,N_15);
nand U854 (N_854,In_2752,In_664);
xnor U855 (N_855,In_88,In_2839);
and U856 (N_856,N_91,N_97);
or U857 (N_857,In_1365,In_1892);
xor U858 (N_858,In_112,In_2997);
nand U859 (N_859,In_2117,In_1072);
or U860 (N_860,In_1690,In_147);
and U861 (N_861,In_190,N_292);
and U862 (N_862,In_1496,In_2028);
xnor U863 (N_863,N_444,N_475);
nand U864 (N_864,In_1611,N_160);
nand U865 (N_865,N_146,In_942);
and U866 (N_866,N_501,In_1553);
xor U867 (N_867,In_1822,N_224);
nand U868 (N_868,N_186,In_464);
or U869 (N_869,In_2169,N_343);
nor U870 (N_870,N_461,In_2151);
nand U871 (N_871,N_238,N_281);
nor U872 (N_872,In_1789,In_708);
nand U873 (N_873,In_1774,In_1299);
and U874 (N_874,In_2410,In_118);
or U875 (N_875,In_1331,In_761);
nand U876 (N_876,N_447,In_1323);
nor U877 (N_877,In_915,In_680);
or U878 (N_878,In_2551,In_2280);
nand U879 (N_879,In_359,N_34);
nor U880 (N_880,In_2304,In_1997);
nand U881 (N_881,In_122,In_976);
or U882 (N_882,In_220,In_2436);
or U883 (N_883,In_2495,In_964);
or U884 (N_884,N_231,In_774);
or U885 (N_885,In_1436,In_1734);
xnor U886 (N_886,N_556,In_444);
and U887 (N_887,In_1538,N_596);
nor U888 (N_888,In_1806,In_2623);
and U889 (N_889,In_992,In_2211);
nand U890 (N_890,N_200,In_2727);
xor U891 (N_891,In_1409,In_1990);
xnor U892 (N_892,In_2565,In_800);
nor U893 (N_893,In_1562,In_703);
nor U894 (N_894,In_382,N_335);
or U895 (N_895,N_179,In_845);
nor U896 (N_896,In_2333,In_2506);
and U897 (N_897,In_2753,In_145);
nor U898 (N_898,In_65,In_2762);
nand U899 (N_899,In_1828,N_213);
nand U900 (N_900,N_67,In_2026);
nand U901 (N_901,N_509,In_2163);
xnor U902 (N_902,In_2975,In_2559);
or U903 (N_903,In_2166,N_261);
nand U904 (N_904,N_466,In_781);
or U905 (N_905,N_216,In_2422);
or U906 (N_906,In_2719,In_345);
nor U907 (N_907,In_2868,In_968);
and U908 (N_908,In_657,In_438);
or U909 (N_909,In_63,N_235);
nand U910 (N_910,In_2831,In_2935);
or U911 (N_911,In_1298,In_2184);
nand U912 (N_912,N_454,In_568);
nand U913 (N_913,In_2339,In_1908);
xor U914 (N_914,In_2453,N_311);
nor U915 (N_915,N_46,In_2132);
or U916 (N_916,In_2027,In_814);
nor U917 (N_917,In_1978,In_1597);
nand U918 (N_918,N_438,In_207);
or U919 (N_919,In_107,In_2713);
nor U920 (N_920,In_2977,N_256);
and U921 (N_921,In_1008,In_2433);
or U922 (N_922,In_1231,N_479);
nand U923 (N_923,N_344,In_1491);
and U924 (N_924,N_486,N_137);
or U925 (N_925,N_505,In_829);
xor U926 (N_926,N_278,In_2693);
nand U927 (N_927,In_815,In_501);
nand U928 (N_928,In_2769,In_2557);
nand U929 (N_929,In_1745,In_1397);
nor U930 (N_930,In_1623,In_1403);
nand U931 (N_931,N_7,In_571);
nand U932 (N_932,N_203,In_1870);
nor U933 (N_933,N_240,In_951);
or U934 (N_934,In_249,In_1309);
or U935 (N_935,In_2062,In_1011);
or U936 (N_936,In_2946,In_366);
nand U937 (N_937,In_2754,In_606);
nor U938 (N_938,In_2093,In_1765);
or U939 (N_939,N_464,In_2665);
or U940 (N_940,In_2957,In_1054);
nor U941 (N_941,In_258,In_2401);
and U942 (N_942,In_1489,N_436);
and U943 (N_943,In_1735,In_2213);
nand U944 (N_944,In_375,N_287);
and U945 (N_945,N_365,N_379);
xnor U946 (N_946,N_140,N_577);
nor U947 (N_947,In_192,In_1860);
xnor U948 (N_948,In_1600,In_20);
and U949 (N_949,In_1253,N_30);
nor U950 (N_950,In_2537,In_1593);
or U951 (N_951,In_1157,N_208);
and U952 (N_952,In_1853,N_482);
and U953 (N_953,In_1791,In_899);
and U954 (N_954,In_414,In_884);
xnor U955 (N_955,In_2084,In_158);
and U956 (N_956,In_183,In_1998);
xnor U957 (N_957,N_502,N_306);
or U958 (N_958,In_1965,In_1161);
xor U959 (N_959,In_477,In_713);
and U960 (N_960,In_2002,N_167);
nor U961 (N_961,N_232,In_2915);
or U962 (N_962,N_585,In_240);
and U963 (N_963,In_2253,In_929);
and U964 (N_964,N_446,In_1464);
nand U965 (N_965,In_2829,N_440);
xnor U966 (N_966,N_594,In_128);
nand U967 (N_967,In_2118,In_257);
nand U968 (N_968,In_1233,In_134);
or U969 (N_969,In_910,In_2845);
and U970 (N_970,N_56,In_226);
and U971 (N_971,In_1473,In_360);
nand U972 (N_972,In_1843,In_45);
nor U973 (N_973,In_1175,In_671);
or U974 (N_974,N_230,In_1367);
or U975 (N_975,In_1737,In_1781);
or U976 (N_976,In_907,N_41);
and U977 (N_977,In_2489,In_2625);
nand U978 (N_978,In_798,In_124);
and U979 (N_979,N_419,In_2390);
nand U980 (N_980,In_2215,In_1650);
or U981 (N_981,In_2503,In_486);
nand U982 (N_982,N_171,In_1170);
nor U983 (N_983,In_2817,N_580);
nand U984 (N_984,N_8,In_141);
nand U985 (N_985,In_860,In_822);
xnor U986 (N_986,In_812,N_581);
nand U987 (N_987,In_1136,N_206);
nor U988 (N_988,N_266,N_595);
nor U989 (N_989,N_376,N_66);
nor U990 (N_990,N_326,N_172);
or U991 (N_991,In_826,In_2050);
or U992 (N_992,In_2584,In_2321);
nor U993 (N_993,In_2886,N_495);
xor U994 (N_994,In_2869,N_42);
nand U995 (N_995,In_519,In_1564);
or U996 (N_996,In_1499,N_389);
nor U997 (N_997,N_432,In_1269);
and U998 (N_998,In_2619,In_1366);
nand U999 (N_999,N_189,N_338);
nor U1000 (N_1000,In_788,In_2509);
nand U1001 (N_1001,In_1101,N_373);
nand U1002 (N_1002,In_53,In_1951);
nor U1003 (N_1003,N_145,In_2966);
or U1004 (N_1004,In_1930,In_1545);
and U1005 (N_1005,In_2836,In_507);
nand U1006 (N_1006,N_144,In_2240);
nand U1007 (N_1007,In_1333,In_1487);
nor U1008 (N_1008,N_506,In_1920);
nor U1009 (N_1009,In_499,In_1986);
nand U1010 (N_1010,In_514,In_505);
xnor U1011 (N_1011,In_1320,In_2080);
nor U1012 (N_1012,N_459,In_2774);
nor U1013 (N_1013,In_2995,In_906);
and U1014 (N_1014,In_2681,In_2233);
or U1015 (N_1015,In_2477,In_2919);
and U1016 (N_1016,In_534,In_2663);
and U1017 (N_1017,In_2104,In_2709);
nand U1018 (N_1018,In_1260,N_194);
nand U1019 (N_1019,In_767,N_341);
and U1020 (N_1020,N_456,N_400);
nor U1021 (N_1021,N_241,In_854);
nand U1022 (N_1022,In_1750,N_380);
nand U1023 (N_1023,In_241,N_269);
or U1024 (N_1024,In_166,In_1384);
nor U1025 (N_1025,In_1579,In_36);
nor U1026 (N_1026,N_321,In_956);
nor U1027 (N_1027,In_2065,In_1205);
nand U1028 (N_1028,N_158,N_142);
nor U1029 (N_1029,In_1768,In_402);
nor U1030 (N_1030,N_29,In_1548);
nor U1031 (N_1031,In_2274,In_2178);
and U1032 (N_1032,N_346,In_252);
and U1033 (N_1033,N_170,N_567);
or U1034 (N_1034,In_1726,In_2889);
nor U1035 (N_1035,In_476,In_620);
and U1036 (N_1036,N_420,In_2119);
nor U1037 (N_1037,In_2162,In_2297);
nand U1038 (N_1038,In_398,In_747);
or U1039 (N_1039,In_698,In_2175);
nand U1040 (N_1040,N_470,In_1215);
and U1041 (N_1041,In_1425,In_2451);
and U1042 (N_1042,In_2061,In_779);
xnor U1043 (N_1043,N_537,In_2871);
or U1044 (N_1044,N_0,In_506);
and U1045 (N_1045,In_1744,In_1555);
nand U1046 (N_1046,In_317,In_2728);
and U1047 (N_1047,In_2033,In_484);
nor U1048 (N_1048,In_79,In_1926);
and U1049 (N_1049,In_692,In_2017);
xnor U1050 (N_1050,In_1814,N_557);
xnor U1051 (N_1051,In_1017,In_2268);
or U1052 (N_1052,In_2546,In_2716);
nand U1053 (N_1053,In_2674,N_493);
or U1054 (N_1054,N_388,N_355);
nor U1055 (N_1055,In_1798,In_1753);
and U1056 (N_1056,N_40,In_1297);
nand U1057 (N_1057,In_1839,N_467);
nor U1058 (N_1058,In_1702,In_2687);
nor U1059 (N_1059,N_43,In_310);
nor U1060 (N_1060,In_1910,In_1424);
nand U1061 (N_1061,N_508,In_1344);
nor U1062 (N_1062,In_662,In_2423);
or U1063 (N_1063,In_893,In_46);
nand U1064 (N_1064,In_1000,In_1996);
nand U1065 (N_1065,In_2996,In_426);
nand U1066 (N_1066,In_511,N_157);
xor U1067 (N_1067,In_928,In_1686);
nand U1068 (N_1068,In_2668,N_242);
and U1069 (N_1069,In_1508,N_197);
nor U1070 (N_1070,In_2356,N_465);
nand U1071 (N_1071,In_1732,N_571);
nor U1072 (N_1072,N_462,In_2242);
nand U1073 (N_1073,N_472,In_2768);
and U1074 (N_1074,In_1529,In_351);
xor U1075 (N_1075,In_177,In_113);
nor U1076 (N_1076,In_1015,N_69);
or U1077 (N_1077,N_526,In_117);
nor U1078 (N_1078,In_674,In_75);
nor U1079 (N_1079,In_1029,N_579);
nor U1080 (N_1080,In_758,In_1823);
nor U1081 (N_1081,N_163,In_2008);
and U1082 (N_1082,N_9,In_2669);
and U1083 (N_1083,In_2918,N_572);
or U1084 (N_1084,N_342,In_2617);
nand U1085 (N_1085,In_1708,In_2820);
nand U1086 (N_1086,In_839,In_751);
nand U1087 (N_1087,In_1829,In_1118);
or U1088 (N_1088,In_510,In_474);
nor U1089 (N_1089,In_1566,N_345);
nor U1090 (N_1090,In_1725,N_127);
nand U1091 (N_1091,In_612,In_1460);
or U1092 (N_1092,In_2004,N_147);
and U1093 (N_1093,In_174,N_525);
or U1094 (N_1094,In_2662,In_599);
and U1095 (N_1095,N_471,N_166);
xnor U1096 (N_1096,In_54,In_667);
and U1097 (N_1097,In_1519,In_933);
nand U1098 (N_1098,In_1338,In_1478);
nor U1099 (N_1099,In_2109,In_871);
nor U1100 (N_1100,In_1947,In_1169);
nor U1101 (N_1101,In_2566,In_221);
xnor U1102 (N_1102,In_1852,In_695);
or U1103 (N_1103,In_1654,In_93);
nand U1104 (N_1104,In_2653,N_421);
or U1105 (N_1105,In_2353,In_998);
and U1106 (N_1106,N_139,In_2882);
and U1107 (N_1107,In_1258,In_1264);
and U1108 (N_1108,In_2105,In_2314);
and U1109 (N_1109,N_316,In_2722);
nand U1110 (N_1110,N_496,In_1688);
or U1111 (N_1111,In_626,In_2010);
or U1112 (N_1112,In_581,N_12);
and U1113 (N_1113,In_2311,In_296);
and U1114 (N_1114,In_583,In_2937);
nor U1115 (N_1115,In_721,N_599);
nor U1116 (N_1116,In_245,N_431);
xnor U1117 (N_1117,In_300,In_2303);
and U1118 (N_1118,In_1376,In_197);
xor U1119 (N_1119,N_201,In_2494);
or U1120 (N_1120,In_448,N_521);
and U1121 (N_1121,In_1931,In_2707);
or U1122 (N_1122,In_268,In_2127);
nor U1123 (N_1123,In_139,In_2181);
and U1124 (N_1124,In_643,N_53);
or U1125 (N_1125,In_2765,N_225);
nor U1126 (N_1126,N_563,N_255);
nand U1127 (N_1127,In_2200,In_558);
nor U1128 (N_1128,In_1578,In_1486);
and U1129 (N_1129,In_1867,N_555);
or U1130 (N_1130,In_619,In_78);
nand U1131 (N_1131,N_211,In_1518);
or U1132 (N_1132,N_251,In_669);
nand U1133 (N_1133,N_350,In_1222);
nor U1134 (N_1134,In_1952,In_1440);
or U1135 (N_1135,In_646,In_2787);
nor U1136 (N_1136,N_417,In_816);
nor U1137 (N_1137,N_149,N_485);
nand U1138 (N_1138,In_1291,In_1311);
and U1139 (N_1139,In_148,In_1739);
nand U1140 (N_1140,In_1179,N_339);
and U1141 (N_1141,In_1357,In_1055);
nand U1142 (N_1142,In_1303,N_219);
nor U1143 (N_1143,In_2994,In_1426);
xor U1144 (N_1144,N_500,In_2561);
nor U1145 (N_1145,In_2826,In_2865);
or U1146 (N_1146,N_182,In_2780);
or U1147 (N_1147,N_212,In_2758);
nand U1148 (N_1148,In_1306,In_2676);
and U1149 (N_1149,N_130,In_1662);
nor U1150 (N_1150,In_2257,In_2474);
or U1151 (N_1151,In_655,In_1228);
or U1152 (N_1152,In_1022,In_807);
or U1153 (N_1153,In_2289,In_2677);
and U1154 (N_1154,N_551,N_569);
nor U1155 (N_1155,In_2069,In_1862);
and U1156 (N_1156,N_398,In_282);
nand U1157 (N_1157,N_18,In_2167);
nor U1158 (N_1158,In_1985,In_1938);
and U1159 (N_1159,N_303,N_512);
and U1160 (N_1160,In_862,In_2368);
nand U1161 (N_1161,In_328,In_2023);
nand U1162 (N_1162,In_2545,In_2440);
and U1163 (N_1163,N_560,N_154);
nor U1164 (N_1164,In_970,In_2347);
nand U1165 (N_1165,In_1896,In_103);
or U1166 (N_1166,In_725,In_2554);
or U1167 (N_1167,In_297,In_487);
nor U1168 (N_1168,In_1536,N_239);
nor U1169 (N_1169,N_561,In_1252);
and U1170 (N_1170,In_3,In_1899);
and U1171 (N_1171,N_426,N_21);
nand U1172 (N_1172,N_327,In_979);
nand U1173 (N_1173,In_1455,In_608);
or U1174 (N_1174,N_117,In_2157);
and U1175 (N_1175,N_392,In_98);
nor U1176 (N_1176,In_2315,In_2783);
and U1177 (N_1177,N_548,In_2993);
nand U1178 (N_1178,In_2612,In_1353);
or U1179 (N_1179,In_2102,In_2536);
xnor U1180 (N_1180,In_2139,In_167);
and U1181 (N_1181,In_2747,N_150);
xnor U1182 (N_1182,In_2313,N_455);
nor U1183 (N_1183,In_2585,In_2106);
nand U1184 (N_1184,In_1236,In_699);
or U1185 (N_1185,N_94,N_504);
nand U1186 (N_1186,In_492,In_926);
and U1187 (N_1187,In_2085,N_250);
or U1188 (N_1188,In_1672,In_2876);
nor U1189 (N_1189,N_244,N_487);
nor U1190 (N_1190,In_2609,In_729);
nor U1191 (N_1191,In_237,In_1691);
nand U1192 (N_1192,In_2300,In_2522);
nand U1193 (N_1193,In_1714,In_1497);
nand U1194 (N_1194,In_898,In_1337);
or U1195 (N_1195,In_1804,N_70);
or U1196 (N_1196,In_2481,In_972);
nand U1197 (N_1197,In_218,In_2540);
or U1198 (N_1198,N_227,In_1014);
xnor U1199 (N_1199,N_450,In_728);
and U1200 (N_1200,N_814,In_2746);
and U1201 (N_1201,In_1854,N_1066);
xnor U1202 (N_1202,In_1031,N_891);
nor U1203 (N_1203,N_625,In_2490);
nor U1204 (N_1204,N_188,In_2701);
nor U1205 (N_1205,In_1192,In_94);
nor U1206 (N_1206,N_859,N_651);
and U1207 (N_1207,In_2098,In_2846);
or U1208 (N_1208,In_2630,In_950);
and U1209 (N_1209,N_717,In_1718);
or U1210 (N_1210,In_931,N_284);
nand U1211 (N_1211,In_152,N_533);
nand U1212 (N_1212,N_847,In_2249);
nand U1213 (N_1213,N_807,In_71);
xor U1214 (N_1214,In_302,N_1080);
nand U1215 (N_1215,In_2940,N_789);
nor U1216 (N_1216,N_896,N_246);
nor U1217 (N_1217,In_555,In_1945);
and U1218 (N_1218,In_1919,In_498);
and U1219 (N_1219,N_1041,N_297);
and U1220 (N_1220,N_1185,N_1171);
nand U1221 (N_1221,In_1863,N_1142);
xor U1222 (N_1222,N_583,In_515);
and U1223 (N_1223,N_518,In_840);
nand U1224 (N_1224,In_1207,In_651);
nand U1225 (N_1225,In_2827,In_834);
and U1226 (N_1226,N_574,N_805);
or U1227 (N_1227,N_178,N_414);
nand U1228 (N_1228,N_874,N_620);
or U1229 (N_1229,N_746,N_890);
nand U1230 (N_1230,In_2414,N_820);
nand U1231 (N_1231,N_836,In_253);
and U1232 (N_1232,N_1162,N_940);
nand U1233 (N_1233,N_73,In_2123);
and U1234 (N_1234,In_1568,N_295);
nand U1235 (N_1235,N_249,N_353);
nor U1236 (N_1236,In_2656,N_723);
and U1237 (N_1237,N_1064,N_877);
xor U1238 (N_1238,In_1439,In_706);
nand U1239 (N_1239,N_610,N_334);
nand U1240 (N_1240,N_99,N_102);
nor U1241 (N_1241,In_2499,N_520);
nand U1242 (N_1242,In_985,N_730);
nand U1243 (N_1243,In_1354,N_196);
nor U1244 (N_1244,N_680,In_2416);
nand U1245 (N_1245,N_113,In_2688);
xor U1246 (N_1246,In_2323,N_435);
nor U1247 (N_1247,N_1107,In_2615);
nand U1248 (N_1248,In_1914,N_1070);
and U1249 (N_1249,N_636,In_1165);
or U1250 (N_1250,N_962,N_1146);
nand U1251 (N_1251,In_160,N_1172);
nand U1252 (N_1252,N_234,In_1713);
and U1253 (N_1253,N_952,In_164);
and U1254 (N_1254,In_1186,In_316);
and U1255 (N_1255,In_1498,N_430);
or U1256 (N_1256,In_1094,In_2478);
and U1257 (N_1257,N_908,In_280);
nand U1258 (N_1258,N_498,N_1174);
nand U1259 (N_1259,N_619,In_2220);
nand U1260 (N_1260,In_1387,N_775);
or U1261 (N_1261,In_388,In_2016);
nand U1262 (N_1262,In_2150,N_101);
nand U1263 (N_1263,In_1453,N_834);
or U1264 (N_1264,In_890,N_1094);
and U1265 (N_1265,N_386,In_1591);
nor U1266 (N_1266,N_84,N_1059);
xnor U1267 (N_1267,In_2464,In_2862);
nand U1268 (N_1268,In_530,N_356);
xor U1269 (N_1269,N_1166,N_192);
and U1270 (N_1270,N_1121,In_1415);
nor U1271 (N_1271,In_512,In_1974);
xor U1272 (N_1272,In_80,N_116);
nand U1273 (N_1273,In_295,N_288);
nand U1274 (N_1274,In_62,In_1104);
xnor U1275 (N_1275,In_1977,N_669);
xnor U1276 (N_1276,N_1143,N_745);
nor U1277 (N_1277,In_247,N_690);
or U1278 (N_1278,N_424,N_1084);
and U1279 (N_1279,N_1024,In_2895);
nor U1280 (N_1280,N_494,N_771);
and U1281 (N_1281,In_2500,In_785);
nor U1282 (N_1282,In_1573,In_1572);
xor U1283 (N_1283,In_1655,In_288);
xnor U1284 (N_1284,N_756,In_2550);
or U1285 (N_1285,N_1036,In_848);
nand U1286 (N_1286,In_540,N_5);
or U1287 (N_1287,In_995,N_999);
and U1288 (N_1288,In_984,In_889);
or U1289 (N_1289,In_905,In_435);
nor U1290 (N_1290,N_128,In_1736);
and U1291 (N_1291,In_2575,In_1506);
nand U1292 (N_1292,N_352,In_420);
and U1293 (N_1293,In_2816,In_424);
nand U1294 (N_1294,N_62,In_2298);
nand U1295 (N_1295,N_758,In_2124);
nor U1296 (N_1296,In_960,N_1160);
nand U1297 (N_1297,N_744,N_13);
or U1298 (N_1298,N_1087,N_1089);
nor U1299 (N_1299,In_2046,In_2463);
nand U1300 (N_1300,In_1289,N_738);
xnor U1301 (N_1301,N_374,In_1782);
or U1302 (N_1302,N_882,In_2206);
nand U1303 (N_1303,N_934,In_694);
or U1304 (N_1304,N_930,In_818);
or U1305 (N_1305,N_1114,In_2194);
and U1306 (N_1306,N_274,N_1043);
nor U1307 (N_1307,In_4,In_106);
or U1308 (N_1308,In_778,In_2959);
nor U1309 (N_1309,In_821,N_381);
or U1310 (N_1310,N_645,N_185);
nand U1311 (N_1311,N_1175,N_1039);
nand U1312 (N_1312,N_603,N_946);
and U1313 (N_1313,N_779,N_784);
nand U1314 (N_1314,N_841,N_710);
and U1315 (N_1315,N_676,In_2660);
nor U1316 (N_1316,In_91,N_448);
or U1317 (N_1317,In_2521,N_697);
nor U1318 (N_1318,In_2336,N_840);
or U1319 (N_1319,In_2548,In_663);
nand U1320 (N_1320,In_125,In_204);
nor U1321 (N_1321,In_763,In_879);
xnor U1322 (N_1322,In_400,N_1136);
xnor U1323 (N_1323,In_1454,In_1993);
or U1324 (N_1324,N_904,N_702);
nor U1325 (N_1325,N_720,N_793);
nand U1326 (N_1326,N_827,N_1168);
and U1327 (N_1327,N_319,N_931);
nor U1328 (N_1328,N_968,In_2238);
and U1329 (N_1329,In_2254,N_866);
or U1330 (N_1330,N_977,In_1697);
or U1331 (N_1331,N_1187,N_835);
nor U1332 (N_1332,In_1645,In_1107);
xor U1333 (N_1333,N_918,N_1192);
or U1334 (N_1334,N_312,N_731);
or U1335 (N_1335,In_1866,N_89);
xor U1336 (N_1336,In_1516,N_79);
or U1337 (N_1337,In_2107,In_1595);
nor U1338 (N_1338,In_1145,In_2990);
and U1339 (N_1339,N_1061,N_262);
xor U1340 (N_1340,N_265,In_392);
nand U1341 (N_1341,N_1088,In_2812);
nand U1342 (N_1342,N_752,N_1179);
xor U1343 (N_1343,In_1057,In_2360);
nand U1344 (N_1344,In_2334,N_1027);
or U1345 (N_1345,In_1515,In_2928);
nor U1346 (N_1346,N_644,N_68);
nand U1347 (N_1347,In_2022,In_1326);
and U1348 (N_1348,N_674,In_2095);
nor U1349 (N_1349,In_892,N_61);
nand U1350 (N_1350,In_1362,N_1191);
or U1351 (N_1351,In_2885,In_2260);
and U1352 (N_1352,In_1450,N_1047);
or U1353 (N_1353,In_1220,In_909);
or U1354 (N_1354,In_1820,N_83);
or U1355 (N_1355,In_1895,N_323);
nor U1356 (N_1356,In_1391,In_1026);
nor U1357 (N_1357,N_1152,N_162);
nand U1358 (N_1358,N_1009,N_1078);
nand U1359 (N_1359,In_1181,N_1026);
nand U1360 (N_1360,In_2855,In_18);
and U1361 (N_1361,N_156,N_879);
or U1362 (N_1362,In_716,In_246);
and U1363 (N_1363,N_876,N_131);
or U1364 (N_1364,In_126,N_1091);
nand U1365 (N_1365,N_510,In_419);
nor U1366 (N_1366,In_90,N_1038);
nand U1367 (N_1367,In_2296,N_617);
and U1368 (N_1368,In_2679,N_135);
or U1369 (N_1369,N_503,N_587);
nor U1370 (N_1370,In_2646,N_785);
nor U1371 (N_1371,N_913,In_2859);
or U1372 (N_1372,N_252,In_2425);
nor U1373 (N_1373,In_977,In_2413);
nor U1374 (N_1374,N_957,In_585);
nor U1375 (N_1375,N_919,N_821);
or U1376 (N_1376,N_704,N_592);
or U1377 (N_1377,In_1535,In_2553);
nand U1378 (N_1378,In_2733,N_949);
xnor U1379 (N_1379,In_952,N_886);
nand U1380 (N_1380,N_1013,In_957);
nand U1381 (N_1381,In_120,In_1982);
nand U1382 (N_1382,In_2183,N_722);
or U1383 (N_1383,N_575,In_742);
and U1384 (N_1384,N_169,N_633);
nand U1385 (N_1385,In_2745,In_260);
and U1386 (N_1386,N_1072,In_1984);
or U1387 (N_1387,N_1032,In_2475);
nand U1388 (N_1388,N_614,N_707);
or U1389 (N_1389,In_1805,In_2949);
nor U1390 (N_1390,N_396,N_924);
xnor U1391 (N_1391,In_339,In_1675);
nand U1392 (N_1392,N_1181,N_993);
nand U1393 (N_1393,In_2695,N_50);
and U1394 (N_1394,N_910,N_1060);
nor U1395 (N_1395,N_367,In_2714);
and U1396 (N_1396,In_2833,N_695);
nand U1397 (N_1397,In_720,In_1794);
or U1398 (N_1398,N_622,In_395);
and U1399 (N_1399,N_1120,In_613);
nor U1400 (N_1400,In_2921,In_408);
and U1401 (N_1401,N_109,N_181);
and U1402 (N_1402,N_661,In_2629);
xnor U1403 (N_1403,N_976,N_221);
xnor U1404 (N_1404,N_933,In_2800);
or U1405 (N_1405,N_844,In_2819);
or U1406 (N_1406,N_736,In_1129);
nor U1407 (N_1407,N_842,In_2461);
and U1408 (N_1408,In_1471,In_1176);
and U1409 (N_1409,N_737,In_2724);
xnor U1410 (N_1410,In_678,N_302);
xor U1411 (N_1411,In_2089,In_2366);
or U1412 (N_1412,In_2942,N_843);
nand U1413 (N_1413,N_6,In_2219);
nor U1414 (N_1414,In_1092,N_632);
and U1415 (N_1415,In_2103,In_2363);
or U1416 (N_1416,N_77,In_1412);
nand U1417 (N_1417,In_2115,In_1633);
and U1418 (N_1418,N_943,N_540);
or U1419 (N_1419,N_248,N_1074);
nor U1420 (N_1420,In_1916,In_1627);
or U1421 (N_1421,N_264,N_199);
and U1422 (N_1422,In_1815,N_698);
or U1423 (N_1423,In_26,N_1197);
or U1424 (N_1424,In_1061,N_693);
or U1425 (N_1425,In_1442,In_1799);
and U1426 (N_1426,In_2736,N_916);
and U1427 (N_1427,In_1626,In_2672);
and U1428 (N_1428,In_2586,In_1630);
or U1429 (N_1429,N_729,In_1493);
nand U1430 (N_1430,In_27,N_640);
or U1431 (N_1431,In_1470,In_2790);
nand U1432 (N_1432,In_1550,In_344);
nand U1433 (N_1433,N_451,N_996);
or U1434 (N_1434,N_751,N_1104);
or U1435 (N_1435,In_2927,N_497);
xor U1436 (N_1436,In_1004,N_838);
or U1437 (N_1437,N_315,In_193);
and U1438 (N_1438,N_687,N_490);
nand U1439 (N_1439,In_509,In_1928);
nand U1440 (N_1440,In_1932,In_2741);
or U1441 (N_1441,N_1093,In_1064);
and U1442 (N_1442,N_1167,In_1787);
nor U1443 (N_1443,In_2291,In_2520);
xnor U1444 (N_1444,In_603,N_822);
and U1445 (N_1445,N_180,N_780);
and U1446 (N_1446,N_11,In_1200);
nand U1447 (N_1447,N_1010,N_792);
and U1448 (N_1448,N_357,In_2854);
nor U1449 (N_1449,N_35,N_39);
nand U1450 (N_1450,N_865,In_607);
nor U1451 (N_1451,In_1826,In_1682);
and U1452 (N_1452,N_337,In_1270);
nand U1453 (N_1453,In_1754,In_2350);
nor U1454 (N_1454,In_2493,In_407);
nor U1455 (N_1455,N_1030,N_14);
nand U1456 (N_1456,N_743,N_198);
nor U1457 (N_1457,N_26,In_1495);
or U1458 (N_1458,N_826,N_726);
nand U1459 (N_1459,In_638,In_1740);
and U1460 (N_1460,N_1022,In_459);
and U1461 (N_1461,N_942,In_312);
or U1462 (N_1462,In_277,N_449);
nor U1463 (N_1463,In_2601,N_377);
and U1464 (N_1464,In_149,N_1025);
or U1465 (N_1465,In_851,In_2570);
and U1466 (N_1466,N_1052,N_405);
and U1467 (N_1467,In_776,In_493);
nand U1468 (N_1468,In_685,N_1170);
nor U1469 (N_1469,N_966,N_1173);
nor U1470 (N_1470,N_382,N_871);
xnor U1471 (N_1471,N_954,In_172);
nand U1472 (N_1472,N_228,N_606);
nor U1473 (N_1473,In_1949,In_1681);
nand U1474 (N_1474,N_903,N_925);
nand U1475 (N_1475,N_81,In_1547);
and U1476 (N_1476,N_88,In_1855);
or U1477 (N_1477,N_898,In_2108);
nand U1478 (N_1478,N_641,In_1652);
xor U1479 (N_1479,N_55,In_2187);
nand U1480 (N_1480,N_519,In_2576);
nor U1481 (N_1481,In_40,In_1994);
and U1482 (N_1482,In_744,In_1229);
or U1483 (N_1483,In_162,N_476);
nand U1484 (N_1484,In_846,In_2443);
or U1485 (N_1485,N_463,In_227);
xnor U1486 (N_1486,N_741,N_709);
nor U1487 (N_1487,In_443,N_1029);
or U1488 (N_1488,N_864,In_1644);
nor U1489 (N_1489,N_917,In_1329);
nor U1490 (N_1490,N_1099,N_971);
and U1491 (N_1491,In_114,N_612);
nor U1492 (N_1492,N_778,In_1395);
nor U1493 (N_1493,N_554,In_2906);
or U1494 (N_1494,N_1195,In_790);
nor U1495 (N_1495,In_609,In_1201);
nor U1496 (N_1496,N_921,N_243);
nand U1497 (N_1497,In_2698,In_2766);
xor U1498 (N_1498,N_837,In_69);
nor U1499 (N_1499,N_788,In_887);
and U1500 (N_1500,In_1241,In_403);
or U1501 (N_1501,In_454,In_2899);
or U1502 (N_1502,In_2437,N_670);
xnor U1503 (N_1503,In_707,N_706);
and U1504 (N_1504,N_1155,In_1160);
and U1505 (N_1505,N_928,In_329);
nand U1506 (N_1506,N_786,N_796);
and U1507 (N_1507,In_350,In_1540);
nand U1508 (N_1508,In_2101,In_1957);
or U1509 (N_1509,In_2703,In_885);
and U1510 (N_1510,N_912,N_1086);
and U1511 (N_1511,N_1006,N_897);
or U1512 (N_1512,N_666,N_668);
and U1513 (N_1513,N_1063,In_1413);
or U1514 (N_1514,N_535,In_573);
nand U1515 (N_1515,N_685,In_379);
nand U1516 (N_1516,N_210,In_1307);
or U1517 (N_1517,In_222,N_530);
or U1518 (N_1518,In_2541,In_1864);
nor U1519 (N_1519,In_1110,N_714);
or U1520 (N_1520,N_364,N_1046);
or U1521 (N_1521,N_1067,In_1062);
or U1522 (N_1522,N_1102,N_1117);
and U1523 (N_1523,In_1596,N_601);
or U1524 (N_1524,In_1203,In_1398);
and U1525 (N_1525,In_962,N_653);
and U1526 (N_1526,N_892,In_2896);
and U1527 (N_1527,N_361,N_825);
and U1528 (N_1528,In_919,In_857);
nand U1529 (N_1529,In_2447,N_375);
or U1530 (N_1530,In_2088,N_662);
and U1531 (N_1531,In_1541,In_2328);
nand U1532 (N_1532,In_1249,N_951);
and U1533 (N_1533,In_2484,N_1165);
and U1534 (N_1534,In_2530,In_2231);
nor U1535 (N_1535,N_665,In_689);
or U1536 (N_1536,N_1068,In_1042);
or U1537 (N_1537,N_973,In_170);
nand U1538 (N_1538,N_772,In_2905);
xor U1539 (N_1539,In_888,In_696);
xor U1540 (N_1540,N_1129,In_2424);
nor U1541 (N_1541,In_2917,N_1008);
nand U1542 (N_1542,N_72,In_2469);
or U1543 (N_1543,N_1126,N_770);
nor U1544 (N_1544,N_739,N_516);
nor U1545 (N_1545,N_1018,In_577);
xnor U1546 (N_1546,In_1126,N_795);
and U1547 (N_1547,N_291,N_1071);
or U1548 (N_1548,In_150,In_361);
nor U1549 (N_1549,In_335,In_1602);
and U1550 (N_1550,In_2822,N_1033);
nor U1551 (N_1551,N_1019,N_855);
nor U1552 (N_1552,N_721,In_941);
and U1553 (N_1553,N_656,N_223);
xnor U1554 (N_1554,N_1077,In_1060);
nor U1555 (N_1555,In_1972,In_1369);
and U1556 (N_1556,In_1159,In_1727);
nand U1557 (N_1557,N_347,N_108);
and U1558 (N_1558,In_1255,In_290);
nand U1559 (N_1559,N_78,In_2212);
xor U1560 (N_1560,N_608,N_1076);
nand U1561 (N_1561,N_618,N_104);
nand U1562 (N_1562,N_411,In_2620);
and U1563 (N_1563,N_970,In_1400);
and U1564 (N_1564,In_2198,N_204);
nand U1565 (N_1565,N_749,N_378);
nand U1566 (N_1566,N_412,In_549);
nand U1567 (N_1567,In_1410,In_2031);
nor U1568 (N_1568,In_1634,N_136);
nor U1569 (N_1569,N_1182,In_2682);
or U1570 (N_1570,In_186,In_2141);
nand U1571 (N_1571,N_652,In_396);
xnor U1572 (N_1572,In_1586,N_936);
and U1573 (N_1573,In_2218,N_988);
and U1574 (N_1574,N_1058,In_2305);
and U1575 (N_1575,N_387,N_929);
xnor U1576 (N_1576,In_2452,N_740);
nor U1577 (N_1577,N_961,In_743);
or U1578 (N_1578,N_1113,N_564);
and U1579 (N_1579,N_686,In_132);
nand U1580 (N_1580,In_2332,N_1014);
xor U1581 (N_1581,In_1243,In_2358);
xnor U1582 (N_1582,N_791,In_16);
xor U1583 (N_1583,N_600,N_408);
or U1584 (N_1584,In_1480,N_800);
and U1585 (N_1585,N_332,N_578);
nand U1586 (N_1586,In_1081,N_1125);
or U1587 (N_1587,In_755,In_622);
nand U1588 (N_1588,In_1084,N_1183);
or U1589 (N_1589,N_1054,In_1693);
nand U1590 (N_1590,In_1099,In_2079);
nor U1591 (N_1591,In_2894,In_2603);
and U1592 (N_1592,In_2631,N_768);
nor U1593 (N_1593,N_409,In_1390);
or U1594 (N_1594,In_1923,N_885);
and U1595 (N_1595,N_900,N_922);
or U1596 (N_1596,N_90,In_1827);
or U1597 (N_1597,N_647,In_2580);
and U1598 (N_1598,N_1176,In_1112);
nand U1599 (N_1599,N_428,N_1180);
nand U1600 (N_1600,N_1157,N_833);
nor U1601 (N_1601,N_613,In_433);
or U1602 (N_1602,N_700,N_760);
or U1603 (N_1603,In_1336,In_1166);
nor U1604 (N_1604,N_899,N_1015);
nand U1605 (N_1605,In_870,In_2988);
xor U1606 (N_1606,N_1012,N_967);
nor U1607 (N_1607,N_926,In_594);
nor U1608 (N_1608,N_869,In_1037);
and U1609 (N_1609,In_2866,N_724);
xor U1610 (N_1610,In_983,In_1402);
or U1611 (N_1611,In_2507,N_689);
nor U1612 (N_1612,In_679,In_2992);
and U1613 (N_1613,In_1886,N_634);
nand U1614 (N_1614,N_995,N_517);
and U1615 (N_1615,N_1016,N_433);
nand U1616 (N_1616,N_701,In_2931);
nand U1617 (N_1617,In_1030,In_1780);
or U1618 (N_1618,In_1824,N_177);
and U1619 (N_1619,In_387,In_293);
or U1620 (N_1620,N_1169,In_1903);
or U1621 (N_1621,N_1132,In_1685);
and U1622 (N_1622,N_534,N_831);
and U1623 (N_1623,In_2188,N_280);
nand U1624 (N_1624,In_2515,N_747);
nor U1625 (N_1625,N_275,N_1190);
nor U1626 (N_1626,In_2691,N_932);
or U1627 (N_1627,N_1044,N_47);
and U1628 (N_1628,N_1053,N_1199);
xor U1629 (N_1629,N_682,In_2718);
or U1630 (N_1630,In_2848,N_963);
and U1631 (N_1631,In_1356,N_1079);
nor U1632 (N_1632,In_1483,N_777);
nor U1633 (N_1633,N_32,In_1817);
nor U1634 (N_1634,In_1640,N_1164);
nor U1635 (N_1635,In_2408,In_2252);
nand U1636 (N_1636,N_732,In_399);
or U1637 (N_1637,In_782,In_551);
nand U1638 (N_1638,In_2020,In_2018);
nor U1639 (N_1639,N_868,N_1144);
nor U1640 (N_1640,N_296,In_552);
xor U1641 (N_1641,In_1651,N_1073);
nand U1642 (N_1642,In_338,In_874);
and U1643 (N_1643,In_2426,N_773);
nand U1644 (N_1644,In_1065,In_2455);
or U1645 (N_1645,In_2135,In_29);
nand U1646 (N_1646,In_913,In_1658);
nor U1647 (N_1647,In_528,N_542);
and U1648 (N_1648,In_2544,N_1138);
nor U1649 (N_1649,N_237,N_829);
or U1650 (N_1650,N_1151,In_1840);
xor U1651 (N_1651,In_1580,In_1810);
and U1652 (N_1652,In_595,N_654);
nand U1653 (N_1653,In_2120,In_1944);
nor U1654 (N_1654,In_1474,N_407);
and U1655 (N_1655,N_371,In_228);
nand U1656 (N_1656,N_1178,In_2547);
and U1657 (N_1657,In_686,N_624);
nor U1658 (N_1658,In_2958,In_2552);
and U1659 (N_1659,N_909,N_849);
nand U1660 (N_1660,In_2276,In_2209);
or U1661 (N_1661,N_161,In_1348);
or U1662 (N_1662,N_1196,N_1108);
and U1663 (N_1663,In_2891,In_13);
xnor U1664 (N_1664,N_401,In_1858);
xor U1665 (N_1665,In_2562,N_678);
and U1666 (N_1666,In_2807,N_64);
nor U1667 (N_1667,In_133,In_637);
nor U1668 (N_1668,In_1451,N_511);
and U1669 (N_1669,In_2064,In_2153);
nor U1670 (N_1670,N_550,In_2189);
and U1671 (N_1671,N_658,In_2965);
or U1672 (N_1672,N_318,In_710);
and U1673 (N_1673,In_1629,N_984);
nor U1674 (N_1674,N_684,In_2047);
xor U1675 (N_1675,N_1194,N_478);
and U1676 (N_1676,N_1148,In_1631);
or U1677 (N_1677,N_1150,In_1086);
xnor U1678 (N_1678,N_733,In_1869);
nor U1679 (N_1679,In_1368,N_615);
nand U1680 (N_1680,N_71,In_1041);
xor U1681 (N_1681,N_798,In_653);
or U1682 (N_1682,In_2864,In_1825);
and U1683 (N_1683,In_2952,N_173);
or U1684 (N_1684,In_1149,N_1111);
xnor U1685 (N_1685,N_366,In_922);
nand U1686 (N_1686,N_1141,N_742);
nor U1687 (N_1687,In_2739,In_2142);
and U1688 (N_1688,N_539,N_1154);
nand U1689 (N_1689,In_1625,N_1123);
or U1690 (N_1690,In_337,In_2039);
nor U1691 (N_1691,In_981,In_832);
or U1692 (N_1692,N_168,N_895);
nand U1693 (N_1693,N_889,In_2814);
nor U1694 (N_1694,In_225,In_2597);
or U1695 (N_1695,In_1459,N_958);
nor U1696 (N_1696,N_832,In_1915);
and U1697 (N_1697,N_304,N_44);
nor U1698 (N_1698,In_1217,In_841);
and U1699 (N_1699,In_1723,N_969);
or U1700 (N_1700,N_1092,In_2531);
and U1701 (N_1701,N_790,In_2177);
nor U1702 (N_1702,In_2341,N_1119);
nor U1703 (N_1703,N_597,In_1834);
xnor U1704 (N_1704,In_1711,In_2649);
nor U1705 (N_1705,In_2853,N_121);
xor U1706 (N_1706,In_2237,N_907);
nand U1707 (N_1707,N_631,N_1003);
or U1708 (N_1708,In_2266,In_1966);
or U1709 (N_1709,In_1079,In_2193);
and U1710 (N_1710,In_1934,In_2666);
nand U1711 (N_1711,N_1184,N_990);
and U1712 (N_1712,In_489,N_948);
nor U1713 (N_1713,N_25,In_2622);
and U1714 (N_1714,N_853,In_185);
or U1715 (N_1715,N_878,N_716);
nand U1716 (N_1716,In_2223,In_1796);
nand U1717 (N_1717,In_1504,N_1007);
or U1718 (N_1718,N_1002,In_2078);
xor U1719 (N_1719,In_553,N_604);
xnor U1720 (N_1720,N_1147,N_794);
nor U1721 (N_1721,N_49,In_911);
and U1722 (N_1722,N_1097,In_730);
xor U1723 (N_1723,In_1701,In_397);
xor U1724 (N_1724,In_66,In_2588);
xnor U1725 (N_1725,In_1819,In_2643);
nand U1726 (N_1726,In_2667,In_1771);
nand U1727 (N_1727,N_884,In_456);
and U1728 (N_1728,In_2932,In_2456);
nor U1729 (N_1729,N_1153,N_875);
or U1730 (N_1730,In_234,N_854);
and U1731 (N_1731,In_1020,N_781);
or U1732 (N_1732,N_638,N_98);
or U1733 (N_1733,N_358,N_719);
and U1734 (N_1734,In_861,In_2250);
nand U1735 (N_1735,N_850,In_1557);
nor U1736 (N_1736,In_2319,N_329);
or U1737 (N_1737,In_1837,N_1011);
nand U1738 (N_1738,N_573,In_1168);
nand U1739 (N_1739,N_1037,N_635);
nand U1740 (N_1740,In_736,In_367);
and U1741 (N_1741,N_1133,In_2364);
nor U1742 (N_1742,In_650,N_902);
nand U1743 (N_1743,N_1156,N_776);
and U1744 (N_1744,N_1105,In_2508);
nand U1745 (N_1745,In_2704,In_1859);
nand U1746 (N_1746,N_305,In_2479);
xor U1747 (N_1747,In_137,In_1906);
or U1748 (N_1748,N_1051,N_923);
nand U1749 (N_1749,N_299,N_828);
nor U1750 (N_1750,In_1187,N_410);
and U1751 (N_1751,N_422,In_704);
and U1752 (N_1752,N_429,In_1364);
nand U1753 (N_1753,In_163,N_1085);
xnor U1754 (N_1754,N_728,In_536);
nand U1755 (N_1755,N_217,In_1267);
or U1756 (N_1756,In_189,In_1992);
nor U1757 (N_1757,In_2759,N_994);
nor U1758 (N_1758,N_1083,In_406);
or U1759 (N_1759,In_2705,N_439);
and U1760 (N_1760,In_2170,In_2924);
or U1761 (N_1761,N_887,In_1313);
and U1762 (N_1762,N_880,N_787);
xor U1763 (N_1763,In_1131,N_85);
and U1764 (N_1764,In_1581,In_576);
and U1765 (N_1765,N_705,N_911);
and U1766 (N_1766,In_2307,N_1193);
and U1767 (N_1767,In_2285,In_1182);
nor U1768 (N_1768,In_2497,In_37);
nor U1769 (N_1769,In_2405,In_961);
or U1770 (N_1770,N_474,In_556);
xor U1771 (N_1771,In_1423,N_819);
or U1772 (N_1772,In_1074,In_2165);
and U1773 (N_1773,N_1122,N_955);
or U1774 (N_1774,N_522,N_960);
nor U1775 (N_1775,In_1488,N_810);
xnor U1776 (N_1776,N_1139,In_2971);
and U1777 (N_1777,In_830,N_576);
nor U1778 (N_1778,N_901,N_1075);
nor U1779 (N_1779,N_605,N_1000);
nor U1780 (N_1780,N_523,In_1174);
and U1781 (N_1781,N_1048,N_1127);
and U1782 (N_1782,In_2867,In_1292);
nand U1783 (N_1783,N_856,In_1001);
xor U1784 (N_1784,In_315,N_715);
or U1785 (N_1785,N_852,In_1314);
and U1786 (N_1786,N_1055,In_2381);
and U1787 (N_1787,In_1543,N_642);
or U1788 (N_1788,In_2763,N_106);
nand U1789 (N_1789,N_1177,In_12);
or U1790 (N_1790,N_322,N_1096);
nor U1791 (N_1791,N_406,N_975);
nor U1792 (N_1792,In_1143,In_1588);
nand U1793 (N_1793,In_1724,In_1010);
nor U1794 (N_1794,N_1069,N_991);
or U1795 (N_1795,N_986,In_2795);
nand U1796 (N_1796,In_673,In_2301);
and U1797 (N_1797,N_93,In_2435);
or U1798 (N_1798,In_1874,In_715);
nand U1799 (N_1799,N_324,N_860);
and U1800 (N_1800,N_1569,N_1362);
and U1801 (N_1801,N_667,N_808);
nor U1802 (N_1802,N_972,N_1649);
or U1803 (N_1803,N_1638,N_1364);
and U1804 (N_1804,N_1360,N_1109);
nor U1805 (N_1805,N_1130,N_384);
nor U1806 (N_1806,N_1752,N_1585);
nand U1807 (N_1807,In_2512,N_1632);
nor U1808 (N_1808,N_1241,N_1527);
and U1809 (N_1809,N_1627,In_868);
or U1810 (N_1810,N_1737,N_725);
and U1811 (N_1811,N_155,N_621);
nor U1812 (N_1812,N_195,N_1749);
or U1813 (N_1813,N_1355,N_1219);
and U1814 (N_1814,N_1686,N_607);
nor U1815 (N_1815,N_1441,In_356);
and U1816 (N_1816,In_648,N_1418);
and U1817 (N_1817,In_1590,N_1534);
or U1818 (N_1818,N_1348,In_1379);
nor U1819 (N_1819,N_107,N_1466);
and U1820 (N_1820,N_1320,In_42);
nand U1821 (N_1821,N_1384,N_1528);
and U1822 (N_1822,N_1381,N_1584);
nor U1823 (N_1823,In_2171,N_1688);
xnor U1824 (N_1824,N_1442,N_1504);
nor U1825 (N_1825,N_1616,N_368);
nor U1826 (N_1826,N_294,N_54);
xor U1827 (N_1827,In_1694,In_2270);
nor U1828 (N_1828,N_1578,N_1318);
xor U1829 (N_1829,N_1586,N_1407);
or U1830 (N_1830,In_123,N_423);
or U1831 (N_1831,In_2577,N_992);
nand U1832 (N_1832,N_1427,N_691);
nor U1833 (N_1833,In_1199,N_1495);
or U1834 (N_1834,N_1660,In_633);
nand U1835 (N_1835,N_1572,N_271);
or U1836 (N_1836,N_1602,N_207);
and U1837 (N_1837,N_1748,N_659);
and U1838 (N_1838,In_1345,N_1789);
nand U1839 (N_1839,N_1394,In_187);
or U1840 (N_1840,N_245,N_165);
nor U1841 (N_1841,N_184,N_1550);
nand U1842 (N_1842,In_1570,N_1304);
and U1843 (N_1843,N_1343,In_1980);
or U1844 (N_1844,In_2581,N_1598);
xnor U1845 (N_1845,N_1573,N_639);
or U1846 (N_1846,In_2738,N_1716);
nor U1847 (N_1847,In_1446,N_1392);
nor U1848 (N_1848,N_1425,N_1005);
or U1849 (N_1849,N_549,N_348);
and U1850 (N_1850,N_1396,N_1506);
or U1851 (N_1851,In_1431,N_483);
xnor U1852 (N_1852,N_1476,N_1536);
or U1853 (N_1853,N_1450,N_218);
or U1854 (N_1854,N_1189,N_1634);
nand U1855 (N_1855,N_1349,N_1551);
and U1856 (N_1856,N_1731,N_1494);
xnor U1857 (N_1857,N_317,N_1735);
and U1858 (N_1858,In_864,N_1582);
nand U1859 (N_1859,N_1736,N_1723);
nand U1860 (N_1860,N_1116,N_1780);
and U1861 (N_1861,N_1714,N_1332);
or U1862 (N_1862,N_1763,N_671);
and U1863 (N_1863,N_1258,In_381);
nand U1864 (N_1864,N_906,N_1298);
and U1865 (N_1865,N_1408,In_1077);
or U1866 (N_1866,N_1677,N_1758);
nand U1867 (N_1867,N_679,In_349);
and U1868 (N_1868,N_1276,In_307);
and U1869 (N_1869,N_1095,N_1422);
nand U1870 (N_1870,In_1565,N_1514);
or U1871 (N_1871,N_1614,N_1438);
nor U1872 (N_1872,N_1786,N_394);
or U1873 (N_1873,N_1788,N_1545);
and U1874 (N_1874,N_443,In_532);
or U1875 (N_1875,N_1727,N_1775);
xnor U1876 (N_1876,N_1511,N_1245);
nor U1877 (N_1877,N_437,N_1202);
nand U1878 (N_1878,In_173,N_1200);
nand U1879 (N_1879,N_1698,N_1031);
or U1880 (N_1880,N_1314,N_1574);
nor U1881 (N_1881,N_1215,N_1591);
nand U1882 (N_1882,In_1575,N_1553);
nand U1883 (N_1883,N_363,N_1315);
nand U1884 (N_1884,In_1613,N_1712);
or U1885 (N_1885,N_434,In_524);
nand U1886 (N_1886,N_1691,In_1075);
nor U1887 (N_1887,N_1718,N_1730);
or U1888 (N_1888,In_764,N_1299);
nand U1889 (N_1889,N_703,N_1242);
nor U1890 (N_1890,N_1657,N_1503);
xnor U1891 (N_1891,N_1244,N_1567);
nand U1892 (N_1892,N_812,In_283);
or U1893 (N_1893,N_1268,N_1352);
and U1894 (N_1894,N_870,N_1681);
and U1895 (N_1895,In_2373,N_1717);
and U1896 (N_1896,In_1783,N_1741);
and U1897 (N_1897,N_1414,N_1216);
xor U1898 (N_1898,N_1020,N_1254);
xor U1899 (N_1899,In_2781,N_1502);
or U1900 (N_1900,N_1629,N_883);
nor U1901 (N_1901,N_1546,In_1322);
nor U1902 (N_1902,N_301,N_1222);
xor U1903 (N_1903,N_1112,N_650);
or U1904 (N_1904,N_1001,N_143);
nand U1905 (N_1905,N_1376,N_1556);
nand U1906 (N_1906,N_51,N_489);
nand U1907 (N_1907,N_1531,N_1600);
or U1908 (N_1908,N_1778,In_2192);
or U1909 (N_1909,N_570,N_3);
xor U1910 (N_1910,N_558,In_2164);
nor U1911 (N_1911,N_1239,N_1785);
or U1912 (N_1912,N_978,In_645);
nand U1913 (N_1913,N_754,N_1519);
and U1914 (N_1914,N_1101,In_1882);
and U1915 (N_1915,N_1238,N_1410);
and U1916 (N_1916,In_1671,N_1365);
and U1917 (N_1917,N_1501,N_1554);
nor U1918 (N_1918,N_657,In_975);
xor U1919 (N_1919,N_759,In_219);
nor U1920 (N_1920,N_1322,N_1278);
and U1921 (N_1921,N_1398,N_1768);
or U1922 (N_1922,N_1443,N_1754);
or U1923 (N_1923,N_1473,N_1766);
and U1924 (N_1924,N_1188,N_1255);
or U1925 (N_1925,N_1333,N_1577);
and U1926 (N_1926,In_324,In_1709);
and U1927 (N_1927,In_1964,N_1272);
nand U1928 (N_1928,N_96,N_677);
nand U1929 (N_1929,N_1761,N_905);
nor U1930 (N_1930,N_260,N_1608);
and U1931 (N_1931,N_1237,N_1225);
or U1932 (N_1932,N_441,In_795);
and U1933 (N_1933,N_1491,N_648);
nand U1934 (N_1934,N_134,N_1706);
nor U1935 (N_1935,In_1227,N_1377);
or U1936 (N_1936,N_1635,N_1500);
nor U1937 (N_1937,N_1659,In_1230);
nor U1938 (N_1938,N_965,N_1583);
nand U1939 (N_1939,N_1652,N_1799);
and U1940 (N_1940,N_1415,In_786);
nor U1941 (N_1941,In_1981,In_683);
xor U1942 (N_1942,N_1439,N_1389);
or U1943 (N_1943,In_2568,N_359);
and U1944 (N_1944,N_1436,N_1021);
and U1945 (N_1945,N_1680,N_532);
nor U1946 (N_1946,N_1339,In_2793);
nor U1947 (N_1947,N_1779,N_1689);
and U1948 (N_1948,N_1416,In_155);
or U1949 (N_1949,N_152,N_1571);
and U1950 (N_1950,In_897,N_1430);
or U1951 (N_1951,N_1581,N_893);
or U1952 (N_1952,N_1651,N_1482);
or U1953 (N_1953,N_1312,In_600);
nor U1954 (N_1954,N_1746,N_1284);
and U1955 (N_1955,In_2159,N_1198);
nor U1956 (N_1956,N_1363,N_1767);
xor U1957 (N_1957,N_1004,N_1693);
and U1958 (N_1958,N_1687,In_1639);
xnor U1959 (N_1959,N_1391,N_110);
and U1960 (N_1960,N_1560,In_1811);
nand U1961 (N_1961,N_1461,In_2126);
nand U1962 (N_1962,In_639,N_1300);
nor U1963 (N_1963,In_1040,In_2525);
xor U1964 (N_1964,In_1420,N_672);
and U1965 (N_1965,N_851,N_1106);
nor U1966 (N_1966,N_1224,N_974);
and U1967 (N_1967,In_421,In_2379);
and U1968 (N_1968,N_1448,In_2613);
nand U1969 (N_1969,In_2074,N_1295);
xnor U1970 (N_1970,In_9,N_1429);
and U1971 (N_1971,N_1508,N_1711);
xor U1972 (N_1972,N_1379,N_873);
and U1973 (N_1973,N_1475,In_2144);
or U1974 (N_1974,In_1500,N_1543);
nor U1975 (N_1975,N_1499,In_872);
or U1976 (N_1976,N_664,N_1353);
nand U1977 (N_1977,N_1675,N_1601);
or U1978 (N_1978,In_2349,In_99);
nand U1979 (N_1979,N_1062,N_1633);
and U1980 (N_1980,N_1411,In_601);
and U1981 (N_1981,In_2012,N_1794);
and U1982 (N_1982,N_1751,N_1462);
or U1983 (N_1983,In_924,N_1366);
nor U1984 (N_1984,In_2962,N_1424);
nand U1985 (N_1985,N_1724,N_945);
nand U1986 (N_1986,In_1295,N_1537);
xnor U1987 (N_1987,N_1158,In_971);
and U1988 (N_1988,N_1286,N_1217);
and U1989 (N_1989,N_290,In_447);
nor U1990 (N_1990,N_1742,N_1640);
or U1991 (N_1991,N_1517,N_1399);
nor U1992 (N_1992,In_610,N_1274);
nand U1993 (N_1993,N_987,N_1690);
and U1994 (N_1994,N_1262,N_857);
and U1995 (N_1995,In_323,In_2526);
and U1996 (N_1996,In_243,In_1044);
nand U1997 (N_1997,N_699,N_1368);
or U1998 (N_1998,N_1309,N_1787);
or U1999 (N_1999,N_1606,N_755);
or U2000 (N_2000,N_1404,N_1679);
nand U2001 (N_2001,N_1228,In_2518);
and U2002 (N_2002,N_867,N_1760);
nor U2003 (N_2003,N_649,In_429);
nor U2004 (N_2004,N_1658,N_1646);
nor U2005 (N_2005,In_1171,N_1434);
nor U2006 (N_2006,N_1694,In_1653);
and U2007 (N_2007,N_1294,In_1286);
xor U2008 (N_2008,N_753,N_1292);
and U2009 (N_2009,N_1326,N_1486);
and U2010 (N_2010,N_818,N_1421);
nor U2011 (N_2011,N_1103,N_1340);
nand U2012 (N_2012,N_402,In_340);
nand U2013 (N_2013,N_1720,In_1404);
or U2014 (N_2014,N_75,In_624);
or U2015 (N_2015,N_1269,In_2019);
and U2016 (N_2016,In_1534,N_1469);
or U2017 (N_2017,N_1753,N_1209);
nand U2018 (N_2018,N_1647,N_797);
or U2019 (N_2019,In_1106,N_927);
nand U2020 (N_2020,In_2302,N_1615);
nand U2021 (N_2021,N_1465,N_1636);
nor U2022 (N_2022,N_584,N_1544);
nand U2023 (N_2023,N_257,N_816);
nand U2024 (N_2024,In_538,In_1111);
and U2025 (N_2025,N_1208,In_1620);
and U2026 (N_2026,N_259,N_263);
or U2027 (N_2027,N_1603,N_1100);
nor U2028 (N_2028,N_1493,In_2644);
nand U2029 (N_2029,In_586,In_1975);
nor U2030 (N_2030,In_2513,N_1163);
nor U2031 (N_2031,In_2310,In_1730);
and U2032 (N_2032,N_681,N_1373);
and U2033 (N_2033,N_1734,N_655);
or U2034 (N_2034,In_973,In_1193);
nand U2035 (N_2035,N_258,N_1701);
or U2036 (N_2036,N_1496,N_1678);
or U2037 (N_2037,N_1065,N_1774);
or U2038 (N_2038,In_2412,N_1385);
and U2039 (N_2039,N_1207,N_1257);
nor U2040 (N_2040,N_1260,N_1468);
nor U2041 (N_2041,In_1012,N_981);
and U2042 (N_2042,N_947,In_621);
nand U2043 (N_2043,N_1604,In_590);
xor U2044 (N_2044,N_1057,In_2071);
and U2045 (N_2045,N_1729,In_676);
nand U2046 (N_2046,In_1093,In_1139);
and U2047 (N_2047,N_801,In_522);
nand U2048 (N_2048,N_815,In_2227);
nor U2049 (N_2049,N_1524,N_1497);
and U2050 (N_2050,N_1642,In_2881);
and U2051 (N_2051,N_1618,In_314);
nand U2052 (N_2052,N_1612,N_86);
nand U2053 (N_2053,N_1489,N_1211);
xnor U2054 (N_2054,N_1699,N_727);
or U2055 (N_2055,N_1732,N_538);
nor U2056 (N_2056,N_1256,N_1484);
and U2057 (N_2057,N_959,N_950);
nor U2058 (N_2058,In_1669,N_1263);
nor U2059 (N_2059,In_1098,N_1575);
nor U2060 (N_2060,N_1700,N_1243);
nor U2061 (N_2061,N_626,In_278);
nand U2062 (N_2062,N_1128,N_1645);
and U2063 (N_2063,N_914,N_1204);
nor U2064 (N_2064,N_1131,In_2375);
xor U2065 (N_2065,N_1655,N_1464);
or U2066 (N_2066,N_1371,In_690);
nand U2067 (N_2067,N_214,N_1719);
and U2068 (N_2068,In_2172,N_1764);
nand U2069 (N_2069,N_1049,N_1336);
and U2070 (N_2070,In_1621,N_1676);
or U2071 (N_2071,In_1742,In_1302);
nor U2072 (N_2072,N_1374,N_1498);
or U2073 (N_2073,N_1552,In_171);
or U2074 (N_2074,In_1294,N_1725);
nand U2075 (N_2075,N_1722,N_939);
and U2076 (N_2076,N_1710,N_63);
or U2077 (N_2077,N_1643,N_1684);
or U2078 (N_2078,In_1184,N_802);
or U2079 (N_2079,In_2133,In_2259);
nor U2080 (N_2080,N_1588,In_1592);
xor U2081 (N_2081,N_48,N_1653);
nand U2082 (N_2082,N_1650,N_1610);
nor U2083 (N_2083,N_277,N_1017);
nor U2084 (N_2084,N_1311,N_1301);
nand U2085 (N_2085,In_630,N_1370);
or U2086 (N_2086,N_1291,In_652);
and U2087 (N_2087,N_313,In_1598);
and U2088 (N_2088,In_2655,N_1338);
or U2089 (N_2089,N_1685,N_881);
and U2090 (N_2090,N_1715,In_2295);
nor U2091 (N_2091,In_2857,N_507);
or U2092 (N_2092,N_694,N_1437);
and U2093 (N_2093,N_997,N_1666);
and U2094 (N_2094,In_2902,N_1492);
nand U2095 (N_2095,In_1749,N_1221);
nor U2096 (N_2096,N_370,N_330);
nor U2097 (N_2097,N_1265,N_1798);
nor U2098 (N_2098,N_1235,In_1517);
and U2099 (N_2099,In_1905,N_823);
xor U2100 (N_2100,N_1530,N_915);
or U2101 (N_2101,N_1525,In_677);
nand U2102 (N_2102,N_1509,N_1206);
or U2103 (N_2103,N_1283,In_1989);
and U2104 (N_2104,N_1288,In_2287);
or U2105 (N_2105,N_1784,N_1406);
or U2106 (N_2106,N_1232,N_1034);
nand U2107 (N_2107,In_2043,N_1328);
nand U2108 (N_2108,N_861,In_1762);
nor U2109 (N_2109,In_2696,N_1297);
and U2110 (N_2110,In_436,N_95);
or U2111 (N_2111,N_528,N_1617);
xnor U2112 (N_2112,N_1605,In_1954);
or U2113 (N_2113,N_1478,In_2884);
or U2114 (N_2114,N_782,In_1900);
nor U2115 (N_2115,N_1665,N_1446);
nor U2116 (N_2116,In_1310,N_1557);
nand U2117 (N_2117,In_2700,N_799);
xnor U2118 (N_2118,N_1744,N_980);
nand U2119 (N_2119,N_1713,In_384);
or U2120 (N_2120,N_1579,N_1792);
nor U2121 (N_2121,N_1401,N_1743);
nand U2122 (N_2122,N_1229,In_1461);
nand U2123 (N_2123,N_985,N_1673);
nand U2124 (N_2124,N_1565,N_1212);
nand U2125 (N_2125,N_1419,N_1487);
and U2126 (N_2126,In_1963,N_1772);
nand U2127 (N_2127,N_1186,In_2388);
nor U2128 (N_2128,In_2180,N_1334);
or U2129 (N_2129,In_416,N_1644);
nand U2130 (N_2130,N_1704,N_1387);
nor U2131 (N_2131,N_1327,N_1261);
nand U2132 (N_2132,N_1628,N_1342);
or U2133 (N_2133,N_609,N_983);
and U2134 (N_2134,N_1372,In_2318);
and U2135 (N_2135,N_16,In_84);
or U2136 (N_2136,N_1769,N_1279);
nand U2137 (N_2137,In_11,In_2326);
nand U2138 (N_2138,N_1115,N_1426);
nand U2139 (N_2139,N_1323,In_1999);
or U2140 (N_2140,N_202,N_1367);
nor U2141 (N_2141,N_1369,In_2908);
nor U2142 (N_2142,N_536,N_1040);
nand U2143 (N_2143,In_644,N_1563);
nor U2144 (N_2144,N_1435,In_430);
nor U2145 (N_2145,N_1431,In_1293);
and U2146 (N_2146,N_1757,N_1576);
nor U2147 (N_2147,In_1232,N_1630);
nor U2148 (N_2148,N_1739,N_1782);
nand U2149 (N_2149,N_1383,In_2858);
or U2150 (N_2150,N_1518,N_457);
and U2151 (N_2151,N_1354,N_1762);
nand U2152 (N_2152,N_1303,N_1287);
xor U2153 (N_2153,In_2404,N_1459);
or U2154 (N_2154,In_1208,N_1662);
or U2155 (N_2155,N_349,In_564);
or U2156 (N_2156,In_965,N_646);
nand U2157 (N_2157,In_2201,N_1449);
or U2158 (N_2158,N_1683,N_1388);
nor U2159 (N_2159,N_1559,In_974);
or U2160 (N_2160,In_1224,N_1444);
and U2161 (N_2161,N_1510,N_863);
xnor U2162 (N_2162,N_1654,N_1479);
xnor U2163 (N_2163,N_1361,N_1231);
or U2164 (N_2164,N_1471,N_403);
xor U2165 (N_2165,In_1522,N_1620);
nor U2166 (N_2166,N_1275,N_763);
nor U2167 (N_2167,N_1619,In_1987);
or U2168 (N_2168,N_1214,In_2986);
and U2169 (N_2169,N_1035,N_1280);
and U2170 (N_2170,In_2809,N_1624);
nand U2171 (N_2171,N_1535,N_806);
nand U2172 (N_2172,N_1266,N_1023);
or U2173 (N_2173,In_2269,N_1317);
nor U2174 (N_2174,N_1134,N_1795);
or U2175 (N_2175,N_1522,N_1682);
nand U2176 (N_2176,N_683,N_1721);
nor U2177 (N_2177,N_1777,In_623);
nand U2178 (N_2178,In_373,N_1313);
and U2179 (N_2179,N_552,In_2034);
nor U2180 (N_2180,N_1447,In_2348);
nor U2181 (N_2181,N_1203,N_1771);
nand U2182 (N_2182,N_105,N_1135);
and U2183 (N_2183,N_1289,N_1667);
or U2184 (N_2184,N_1733,N_1454);
or U2185 (N_2185,In_389,N_138);
or U2186 (N_2186,N_1490,N_1648);
or U2187 (N_2187,N_1293,N_226);
xor U2188 (N_2188,N_848,N_1580);
xnor U2189 (N_2189,In_2821,N_1270);
nand U2190 (N_2190,N_354,N_830);
and U2191 (N_2191,N_1595,N_1759);
nor U2192 (N_2192,N_1705,N_1773);
nand U2193 (N_2193,N_1335,N_1250);
and U2194 (N_2194,In_1070,N_1310);
and U2195 (N_2195,N_1252,In_267);
nand U2196 (N_2196,In_2873,N_711);
or U2197 (N_2197,N_286,In_142);
and U2198 (N_2198,N_956,N_627);
or U2199 (N_2199,N_1596,N_87);
nor U2200 (N_2200,In_1247,N_283);
and U2201 (N_2201,N_1307,N_1347);
or U2202 (N_2202,N_1562,In_1350);
nor U2203 (N_2203,N_282,N_1783);
and U2204 (N_2204,In_1378,N_1597);
nor U2205 (N_2205,In_1939,N_811);
and U2206 (N_2206,N_1098,In_824);
nand U2207 (N_2207,In_2950,N_1248);
nand U2208 (N_2208,In_775,N_1282);
nand U2209 (N_2209,N_1456,N_1521);
nand U2210 (N_2210,N_1671,N_1590);
and U2211 (N_2211,N_1341,N_1382);
nor U2212 (N_2212,In_1172,N_1045);
nand U2213 (N_2213,N_1621,N_1613);
xor U2214 (N_2214,In_224,N_1453);
nor U2215 (N_2215,N_1296,N_1668);
or U2216 (N_2216,In_1341,N_1285);
nand U2217 (N_2217,N_481,In_2760);
and U2218 (N_2218,In_1604,N_477);
nand U2219 (N_2219,N_1477,N_1290);
and U2220 (N_2220,N_1692,N_1393);
nand U2221 (N_2221,N_817,N_735);
nor U2222 (N_2222,N_1674,N_1337);
and U2223 (N_2223,N_1483,In_2271);
and U2224 (N_2224,In_1955,N_765);
nand U2225 (N_2225,N_1413,N_1423);
or U2226 (N_2226,N_191,N_1082);
nor U2227 (N_2227,N_413,N_1670);
nand U2228 (N_2228,N_1555,N_1118);
nand U2229 (N_2229,N_762,N_998);
nor U2230 (N_2230,In_987,N_1319);
or U2231 (N_2231,In_1221,N_1709);
nor U2232 (N_2232,N_1375,N_1227);
and U2233 (N_2233,N_1755,N_351);
nand U2234 (N_2234,N_1223,In_1373);
nand U2235 (N_2235,N_151,N_1481);
or U2236 (N_2236,N_1050,N_757);
nand U2237 (N_2237,N_1790,N_944);
xor U2238 (N_2238,In_165,In_2306);
or U2239 (N_2239,N_1747,N_1708);
nand U2240 (N_2240,N_839,N_708);
or U2241 (N_2241,N_1472,N_1233);
and U2242 (N_2242,N_1386,In_2290);
and U2243 (N_2243,In_625,In_1467);
or U2244 (N_2244,N_1697,N_1538);
and U2245 (N_2245,In_2013,N_1344);
nor U2246 (N_2246,N_1594,In_2792);
nor U2247 (N_2247,N_1641,N_1230);
or U2248 (N_2248,N_1351,N_1081);
or U2249 (N_2249,N_1623,N_1558);
and U2250 (N_2250,N_1234,In_1576);
or U2251 (N_2251,N_1432,N_1420);
or U2252 (N_2252,N_1205,N_1793);
nor U2253 (N_2253,N_1137,In_1721);
xor U2254 (N_2254,N_629,N_872);
nor U2255 (N_2255,N_1474,N_4);
and U2256 (N_2256,In_1793,In_2532);
or U2257 (N_2257,N_692,N_1259);
nor U2258 (N_2258,N_1599,N_1316);
nor U2259 (N_2259,In_441,In_579);
or U2260 (N_2260,N_982,N_783);
nand U2261 (N_2261,N_813,N_1548);
and U2262 (N_2262,N_289,In_2116);
nor U2263 (N_2263,N_1568,N_1467);
or U2264 (N_2264,In_2863,In_584);
and U2265 (N_2265,N_1251,N_1329);
nand U2266 (N_2266,N_1330,N_320);
and U2267 (N_2267,N_193,N_1397);
nand U2268 (N_2268,N_1346,N_1161);
nand U2269 (N_2269,N_1587,In_2312);
nand U2270 (N_2270,N_1428,N_1308);
nand U2271 (N_2271,In_1615,N_1145);
or U2272 (N_2272,N_935,N_1592);
and U2273 (N_2273,N_637,N_19);
or U2274 (N_2274,N_673,N_1264);
nand U2275 (N_2275,N_1412,In_1665);
xnor U2276 (N_2276,N_1350,N_804);
nand U2277 (N_2277,In_175,N_809);
and U2278 (N_2278,In_1818,N_1570);
or U2279 (N_2279,N_1218,N_1505);
and U2280 (N_2280,N_1380,N_300);
xnor U2281 (N_2281,N_764,N_1523);
or U2282 (N_2282,In_2160,In_1918);
and U2283 (N_2283,N_696,N_1589);
xnor U2284 (N_2284,N_920,In_217);
xor U2285 (N_2285,In_518,N_1470);
nand U2286 (N_2286,N_1541,N_33);
and U2287 (N_2287,N_1539,N_103);
and U2288 (N_2288,N_1305,N_1090);
nand U2289 (N_2289,In_709,N_712);
and U2290 (N_2290,In_1418,N_1140);
nor U2291 (N_2291,N_1253,N_1695);
nand U2292 (N_2292,N_1042,N_1325);
or U2293 (N_2293,N_611,N_1797);
nand U2294 (N_2294,N_1547,In_533);
xnor U2295 (N_2295,N_1281,N_616);
or U2296 (N_2296,N_1460,N_846);
or U2297 (N_2297,N_1656,N_222);
and U2298 (N_2298,N_1669,N_1331);
or U2299 (N_2299,N_1356,N_254);
nand U2300 (N_2300,N_1540,N_28);
nor U2301 (N_2301,N_1028,N_1417);
nand U2302 (N_2302,N_660,In_1301);
or U2303 (N_2303,In_2024,N_1765);
and U2304 (N_2304,In_2838,N_675);
and U2305 (N_2305,N_1542,In_2664);
and U2306 (N_2306,In_675,In_1123);
and U2307 (N_2307,In_750,In_1277);
xnor U2308 (N_2308,N_1756,In_1414);
and U2309 (N_2309,N_953,In_1775);
nand U2310 (N_2310,N_1631,N_1516);
or U2311 (N_2311,N_1726,N_1452);
nand U2312 (N_2312,In_2263,N_858);
nor U2313 (N_2313,N_718,N_582);
or U2314 (N_2314,N_1776,N_1738);
nand U2315 (N_2315,N_1564,N_1213);
or U2316 (N_2316,In_2316,N_1321);
nand U2317 (N_2317,N_1267,N_1740);
and U2318 (N_2318,N_1791,N_1626);
nand U2319 (N_2319,N_1220,N_1745);
nor U2320 (N_2320,In_1242,N_1770);
and U2321 (N_2321,In_1318,In_1679);
nor U2322 (N_2322,N_1395,N_964);
xnor U2323 (N_2323,N_1390,In_1521);
and U2324 (N_2324,N_713,In_50);
and U2325 (N_2325,N_1513,N_1663);
and U2326 (N_2326,N_628,N_767);
xor U2327 (N_2327,In_1865,N_1403);
and U2328 (N_2328,N_1661,N_663);
nor U2329 (N_2329,N_1622,In_1646);
xnor U2330 (N_2330,N_766,N_862);
nand U2331 (N_2331,In_1880,In_1116);
nand U2332 (N_2332,N_1110,In_605);
or U2333 (N_2333,In_2818,N_1702);
and U2334 (N_2334,N_176,N_1358);
nand U2335 (N_2335,In_1816,N_941);
or U2336 (N_2336,N_36,N_1520);
nor U2337 (N_2337,N_1703,N_1781);
or U2338 (N_2338,N_1485,In_2505);
nand U2339 (N_2339,N_1409,In_1068);
and U2340 (N_2340,In_1755,N_623);
or U2341 (N_2341,In_1405,N_774);
and U2342 (N_2342,In_261,N_938);
or U2343 (N_2343,N_1526,N_824);
and U2344 (N_2344,N_309,N_1149);
xnor U2345 (N_2345,N_141,N_1359);
and U2346 (N_2346,N_1345,N_1609);
nor U2347 (N_2347,N_1639,In_1494);
xor U2348 (N_2348,N_100,In_1751);
nor U2349 (N_2349,N_761,N_1402);
nor U2350 (N_2350,N_1433,In_1036);
nor U2351 (N_2351,N_1728,N_937);
nor U2352 (N_2352,In_2834,N_1611);
and U2353 (N_2353,N_1159,In_2916);
or U2354 (N_2354,N_1458,N_688);
nand U2355 (N_2355,N_1463,N_1566);
or U2356 (N_2356,N_602,N_1480);
and U2357 (N_2357,N_1696,N_1277);
nand U2358 (N_2358,N_1455,N_1247);
or U2359 (N_2359,In_867,N_1357);
nor U2360 (N_2360,In_999,In_1382);
nand U2361 (N_2361,N_1707,In_2355);
and U2362 (N_2362,N_1672,In_825);
or U2363 (N_2363,N_1302,N_803);
nand U2364 (N_2364,In_993,N_750);
nand U2365 (N_2365,N_1515,N_1457);
or U2366 (N_2366,In_1383,N_1532);
xnor U2367 (N_2367,N_1378,N_1271);
nor U2368 (N_2368,N_1561,In_371);
nand U2369 (N_2369,In_740,In_2743);
nand U2370 (N_2370,N_1249,In_502);
and U2371 (N_2371,N_1210,N_1625);
nor U2372 (N_2372,N_1488,N_1549);
nor U2373 (N_2373,In_383,N_1512);
nor U2374 (N_2374,In_2403,N_1507);
nor U2375 (N_2375,In_1670,N_310);
nand U2376 (N_2376,N_1533,N_1056);
or U2377 (N_2377,N_1607,N_1246);
nand U2378 (N_2378,In_2651,N_1400);
or U2379 (N_2379,In_2543,N_233);
or U2380 (N_2380,N_894,N_598);
or U2381 (N_2381,N_630,In_866);
or U2382 (N_2382,In_2438,N_1124);
xnor U2383 (N_2383,N_1273,N_544);
xnor U2384 (N_2384,N_1440,N_989);
or U2385 (N_2385,N_124,N_888);
xor U2386 (N_2386,N_1240,N_1529);
nand U2387 (N_2387,N_1593,In_2111);
nand U2388 (N_2388,N_1445,N_1796);
xnor U2389 (N_2389,N_1236,N_1637);
nand U2390 (N_2390,N_1226,N_748);
nor U2391 (N_2391,In_936,N_268);
xnor U2392 (N_2392,N_1405,N_1664);
xnor U2393 (N_2393,N_1324,In_1349);
or U2394 (N_2394,N_1451,N_845);
or U2395 (N_2395,N_74,In_1321);
nor U2396 (N_2396,N_643,N_734);
or U2397 (N_2397,N_272,N_769);
or U2398 (N_2398,N_1306,N_1750);
nand U2399 (N_2399,N_979,N_1201);
or U2400 (N_2400,N_2213,N_2012);
nor U2401 (N_2401,N_2269,N_1972);
xnor U2402 (N_2402,N_2302,N_2310);
xor U2403 (N_2403,N_2284,N_2134);
or U2404 (N_2404,N_2055,N_2068);
nor U2405 (N_2405,N_2201,N_2285);
or U2406 (N_2406,N_2325,N_2211);
and U2407 (N_2407,N_1960,N_1835);
nand U2408 (N_2408,N_2014,N_1858);
nand U2409 (N_2409,N_2172,N_2305);
xnor U2410 (N_2410,N_2150,N_1973);
and U2411 (N_2411,N_2176,N_2322);
and U2412 (N_2412,N_2094,N_2330);
and U2413 (N_2413,N_2158,N_1864);
nand U2414 (N_2414,N_1970,N_2279);
xnor U2415 (N_2415,N_2359,N_1892);
nand U2416 (N_2416,N_2171,N_1860);
nand U2417 (N_2417,N_2178,N_1980);
or U2418 (N_2418,N_2214,N_1852);
and U2419 (N_2419,N_1935,N_1933);
xnor U2420 (N_2420,N_2126,N_2292);
and U2421 (N_2421,N_2095,N_1913);
nor U2422 (N_2422,N_2028,N_2326);
nand U2423 (N_2423,N_2358,N_1848);
and U2424 (N_2424,N_2362,N_2147);
and U2425 (N_2425,N_2007,N_2145);
nor U2426 (N_2426,N_1899,N_2392);
nor U2427 (N_2427,N_2100,N_2329);
and U2428 (N_2428,N_2005,N_1807);
and U2429 (N_2429,N_2203,N_2179);
and U2430 (N_2430,N_2127,N_2166);
and U2431 (N_2431,N_1982,N_1841);
or U2432 (N_2432,N_1989,N_1901);
nand U2433 (N_2433,N_2066,N_2076);
xnor U2434 (N_2434,N_1884,N_1920);
xor U2435 (N_2435,N_1906,N_2016);
or U2436 (N_2436,N_2118,N_2009);
xor U2437 (N_2437,N_2064,N_2247);
nand U2438 (N_2438,N_2257,N_2311);
or U2439 (N_2439,N_2289,N_2104);
or U2440 (N_2440,N_2236,N_2349);
and U2441 (N_2441,N_1844,N_1806);
or U2442 (N_2442,N_2031,N_2390);
and U2443 (N_2443,N_2061,N_1838);
nor U2444 (N_2444,N_2306,N_2137);
nand U2445 (N_2445,N_2174,N_1905);
and U2446 (N_2446,N_2393,N_1976);
xor U2447 (N_2447,N_2320,N_2338);
xor U2448 (N_2448,N_1925,N_2309);
and U2449 (N_2449,N_2394,N_2177);
nand U2450 (N_2450,N_2042,N_1804);
nor U2451 (N_2451,N_2190,N_2114);
nand U2452 (N_2452,N_1996,N_2092);
xor U2453 (N_2453,N_2221,N_1827);
xnor U2454 (N_2454,N_1910,N_2164);
or U2455 (N_2455,N_2207,N_1801);
xnor U2456 (N_2456,N_2335,N_1891);
and U2457 (N_2457,N_1867,N_2002);
nor U2458 (N_2458,N_2381,N_1893);
nor U2459 (N_2459,N_2004,N_2024);
or U2460 (N_2460,N_2108,N_2079);
nand U2461 (N_2461,N_1947,N_2008);
xnor U2462 (N_2462,N_1829,N_2270);
nor U2463 (N_2463,N_1942,N_1941);
and U2464 (N_2464,N_1992,N_1926);
or U2465 (N_2465,N_1997,N_1832);
xor U2466 (N_2466,N_2165,N_2384);
nand U2467 (N_2467,N_2057,N_2345);
or U2468 (N_2468,N_2139,N_2181);
xnor U2469 (N_2469,N_1831,N_2003);
xnor U2470 (N_2470,N_1971,N_2208);
nand U2471 (N_2471,N_2183,N_2136);
and U2472 (N_2472,N_1874,N_2169);
nor U2473 (N_2473,N_2202,N_2367);
nor U2474 (N_2474,N_2343,N_1887);
nand U2475 (N_2475,N_1963,N_1930);
or U2476 (N_2476,N_2131,N_2132);
and U2477 (N_2477,N_1950,N_2280);
nand U2478 (N_2478,N_2121,N_2375);
xnor U2479 (N_2479,N_1965,N_2246);
nand U2480 (N_2480,N_2106,N_2277);
and U2481 (N_2481,N_1800,N_2383);
and U2482 (N_2482,N_2088,N_1911);
and U2483 (N_2483,N_2373,N_2288);
xnor U2484 (N_2484,N_1803,N_1914);
or U2485 (N_2485,N_2113,N_2060);
or U2486 (N_2486,N_2152,N_2017);
or U2487 (N_2487,N_2315,N_2111);
and U2488 (N_2488,N_2116,N_2225);
or U2489 (N_2489,N_1889,N_2380);
xnor U2490 (N_2490,N_1932,N_2205);
nor U2491 (N_2491,N_2197,N_2080);
and U2492 (N_2492,N_1951,N_1962);
or U2493 (N_2493,N_1882,N_2268);
nand U2494 (N_2494,N_2259,N_2049);
nor U2495 (N_2495,N_2010,N_1855);
and U2496 (N_2496,N_2232,N_2244);
and U2497 (N_2497,N_2078,N_2189);
nor U2498 (N_2498,N_2239,N_2101);
and U2499 (N_2499,N_1929,N_1819);
or U2500 (N_2500,N_2091,N_2308);
and U2501 (N_2501,N_2258,N_2307);
nor U2502 (N_2502,N_2097,N_1846);
xor U2503 (N_2503,N_1869,N_1938);
nand U2504 (N_2504,N_2245,N_2224);
or U2505 (N_2505,N_2048,N_1810);
and U2506 (N_2506,N_2160,N_2252);
xnor U2507 (N_2507,N_1902,N_2046);
nand U2508 (N_2508,N_2267,N_1999);
or U2509 (N_2509,N_1988,N_2355);
nand U2510 (N_2510,N_2196,N_2281);
nand U2511 (N_2511,N_2243,N_2102);
or U2512 (N_2512,N_2083,N_2368);
and U2513 (N_2513,N_2153,N_2036);
nor U2514 (N_2514,N_1948,N_1880);
and U2515 (N_2515,N_2276,N_2334);
or U2516 (N_2516,N_1866,N_2364);
or U2517 (N_2517,N_2220,N_1854);
or U2518 (N_2518,N_2229,N_2140);
and U2519 (N_2519,N_2303,N_2328);
nand U2520 (N_2520,N_2347,N_2282);
or U2521 (N_2521,N_2223,N_2143);
nor U2522 (N_2522,N_1824,N_1915);
nand U2523 (N_2523,N_1837,N_2234);
and U2524 (N_2524,N_1991,N_1818);
nand U2525 (N_2525,N_2059,N_2058);
or U2526 (N_2526,N_2301,N_1834);
or U2527 (N_2527,N_1817,N_2238);
nand U2528 (N_2528,N_2337,N_1978);
or U2529 (N_2529,N_2378,N_2099);
nor U2530 (N_2530,N_2209,N_2210);
and U2531 (N_2531,N_2021,N_2151);
or U2532 (N_2532,N_1944,N_2141);
and U2533 (N_2533,N_2093,N_2191);
nor U2534 (N_2534,N_1875,N_1968);
and U2535 (N_2535,N_1928,N_2045);
nand U2536 (N_2536,N_1850,N_2256);
nor U2537 (N_2537,N_2346,N_2212);
nor U2538 (N_2538,N_2129,N_1990);
nand U2539 (N_2539,N_2295,N_1871);
and U2540 (N_2540,N_1809,N_1853);
nand U2541 (N_2541,N_1987,N_1956);
xnor U2542 (N_2542,N_2228,N_2148);
nand U2543 (N_2543,N_1815,N_2299);
or U2544 (N_2544,N_1908,N_2149);
nand U2545 (N_2545,N_2231,N_2371);
nand U2546 (N_2546,N_2218,N_2376);
or U2547 (N_2547,N_1808,N_1878);
and U2548 (N_2548,N_2242,N_1862);
or U2549 (N_2549,N_2386,N_2037);
or U2550 (N_2550,N_1975,N_2233);
xnor U2551 (N_2551,N_1821,N_2157);
or U2552 (N_2552,N_2314,N_2366);
and U2553 (N_2553,N_2204,N_1895);
or U2554 (N_2554,N_2065,N_2318);
and U2555 (N_2555,N_2047,N_2348);
or U2556 (N_2556,N_2109,N_2173);
nand U2557 (N_2557,N_2250,N_2357);
or U2558 (N_2558,N_2027,N_1856);
or U2559 (N_2559,N_1903,N_1857);
or U2560 (N_2560,N_2087,N_2025);
nor U2561 (N_2561,N_1877,N_2133);
nor U2562 (N_2562,N_1885,N_2275);
nand U2563 (N_2563,N_2369,N_2274);
xor U2564 (N_2564,N_1812,N_2188);
or U2565 (N_2565,N_2029,N_1964);
nor U2566 (N_2566,N_1966,N_2331);
or U2567 (N_2567,N_1912,N_2217);
and U2568 (N_2568,N_2324,N_1974);
or U2569 (N_2569,N_2265,N_1890);
nor U2570 (N_2570,N_2241,N_2001);
and U2571 (N_2571,N_2070,N_2163);
nand U2572 (N_2572,N_1888,N_2353);
and U2573 (N_2573,N_2138,N_2071);
and U2574 (N_2574,N_2184,N_1825);
and U2575 (N_2575,N_1979,N_1943);
nand U2576 (N_2576,N_2119,N_1953);
nor U2577 (N_2577,N_1937,N_1945);
nor U2578 (N_2578,N_2086,N_2255);
nor U2579 (N_2579,N_2344,N_2056);
nand U2580 (N_2580,N_2170,N_1983);
xor U2581 (N_2581,N_1961,N_1816);
or U2582 (N_2582,N_2354,N_2273);
nand U2583 (N_2583,N_2293,N_2044);
and U2584 (N_2584,N_2222,N_2352);
nand U2585 (N_2585,N_1828,N_2041);
nand U2586 (N_2586,N_2248,N_1811);
nor U2587 (N_2587,N_2263,N_1886);
nand U2588 (N_2588,N_2193,N_1917);
nor U2589 (N_2589,N_2074,N_2240);
or U2590 (N_2590,N_1870,N_1986);
and U2591 (N_2591,N_1923,N_1826);
and U2592 (N_2592,N_2135,N_2105);
nand U2593 (N_2593,N_2006,N_2261);
nand U2594 (N_2594,N_1839,N_1805);
nor U2595 (N_2595,N_2385,N_1897);
nor U2596 (N_2596,N_1936,N_2327);
xnor U2597 (N_2597,N_1967,N_2249);
nand U2598 (N_2598,N_2374,N_2144);
nand U2599 (N_2599,N_1919,N_2198);
nor U2600 (N_2600,N_2332,N_1879);
nand U2601 (N_2601,N_2199,N_2351);
nand U2602 (N_2602,N_1952,N_2013);
nor U2603 (N_2603,N_2278,N_2339);
nor U2604 (N_2604,N_1836,N_2216);
xnor U2605 (N_2605,N_1849,N_2391);
nand U2606 (N_2606,N_2067,N_2283);
nand U2607 (N_2607,N_2082,N_2363);
and U2608 (N_2608,N_2075,N_1940);
and U2609 (N_2609,N_2341,N_2266);
nand U2610 (N_2610,N_2388,N_2312);
and U2611 (N_2611,N_1916,N_2396);
xor U2612 (N_2612,N_2186,N_1939);
nand U2613 (N_2613,N_2015,N_1830);
nor U2614 (N_2614,N_1840,N_2297);
or U2615 (N_2615,N_2206,N_2018);
nand U2616 (N_2616,N_2096,N_2146);
nand U2617 (N_2617,N_2040,N_2395);
and U2618 (N_2618,N_2124,N_2286);
nor U2619 (N_2619,N_1959,N_1949);
and U2620 (N_2620,N_2185,N_2054);
nor U2621 (N_2621,N_1865,N_1981);
and U2622 (N_2622,N_2072,N_1847);
nor U2623 (N_2623,N_2272,N_2077);
or U2624 (N_2624,N_2382,N_1843);
and U2625 (N_2625,N_2291,N_1863);
or U2626 (N_2626,N_1995,N_1924);
nand U2627 (N_2627,N_1909,N_2115);
or U2628 (N_2628,N_2317,N_1993);
and U2629 (N_2629,N_2154,N_2237);
nor U2630 (N_2630,N_2084,N_2398);
nor U2631 (N_2631,N_2032,N_1907);
nor U2632 (N_2632,N_2063,N_2011);
or U2633 (N_2633,N_2187,N_2200);
xnor U2634 (N_2634,N_1896,N_2107);
nor U2635 (N_2635,N_1984,N_2264);
nand U2636 (N_2636,N_2030,N_2377);
and U2637 (N_2637,N_2313,N_2123);
nand U2638 (N_2638,N_1823,N_1845);
xnor U2639 (N_2639,N_2321,N_1898);
or U2640 (N_2640,N_2038,N_2182);
nand U2641 (N_2641,N_2142,N_1894);
xnor U2642 (N_2642,N_1820,N_1969);
nor U2643 (N_2643,N_2022,N_1873);
nand U2644 (N_2644,N_2298,N_1883);
nor U2645 (N_2645,N_2035,N_2175);
or U2646 (N_2646,N_2336,N_2120);
or U2647 (N_2647,N_2370,N_2168);
nand U2648 (N_2648,N_1922,N_2167);
xor U2649 (N_2649,N_1861,N_2069);
and U2650 (N_2650,N_2287,N_2156);
or U2651 (N_2651,N_2110,N_1994);
and U2652 (N_2652,N_2379,N_2340);
or U2653 (N_2653,N_1822,N_2254);
and U2654 (N_2654,N_2260,N_2062);
and U2655 (N_2655,N_1955,N_2050);
and U2656 (N_2656,N_2180,N_2161);
nor U2657 (N_2657,N_1931,N_2389);
nand U2658 (N_2658,N_2235,N_2034);
and U2659 (N_2659,N_2033,N_1904);
xor U2660 (N_2660,N_2300,N_1918);
xor U2661 (N_2661,N_2262,N_1957);
nor U2662 (N_2662,N_2051,N_2130);
xor U2663 (N_2663,N_2271,N_2304);
and U2664 (N_2664,N_2226,N_1985);
or U2665 (N_2665,N_2192,N_1859);
xnor U2666 (N_2666,N_2019,N_1872);
nor U2667 (N_2667,N_2215,N_1900);
nand U2668 (N_2668,N_2361,N_2290);
nor U2669 (N_2669,N_2365,N_2053);
and U2670 (N_2670,N_1842,N_1868);
and U2671 (N_2671,N_1927,N_2194);
xor U2672 (N_2672,N_1977,N_1998);
nand U2673 (N_2673,N_2043,N_2103);
and U2674 (N_2674,N_2073,N_1954);
or U2675 (N_2675,N_2081,N_2397);
nand U2676 (N_2676,N_1813,N_2387);
xor U2677 (N_2677,N_2085,N_2342);
and U2678 (N_2678,N_2195,N_1958);
xnor U2679 (N_2679,N_2122,N_1876);
or U2680 (N_2680,N_2251,N_1934);
and U2681 (N_2681,N_2316,N_2333);
and U2682 (N_2682,N_1921,N_2020);
or U2683 (N_2683,N_2219,N_2000);
or U2684 (N_2684,N_2350,N_2356);
and U2685 (N_2685,N_2230,N_1946);
nor U2686 (N_2686,N_2125,N_2253);
or U2687 (N_2687,N_2112,N_2098);
nor U2688 (N_2688,N_2155,N_2360);
nor U2689 (N_2689,N_2323,N_2090);
nor U2690 (N_2690,N_1814,N_2159);
xor U2691 (N_2691,N_1881,N_2372);
or U2692 (N_2692,N_2023,N_2117);
nand U2693 (N_2693,N_1833,N_2296);
xor U2694 (N_2694,N_2227,N_2294);
nand U2695 (N_2695,N_2026,N_2162);
nor U2696 (N_2696,N_1802,N_1851);
or U2697 (N_2697,N_2128,N_2399);
nand U2698 (N_2698,N_2319,N_2089);
xor U2699 (N_2699,N_2039,N_2052);
nand U2700 (N_2700,N_2327,N_2221);
nand U2701 (N_2701,N_1893,N_1934);
nor U2702 (N_2702,N_2045,N_2191);
and U2703 (N_2703,N_1864,N_2353);
or U2704 (N_2704,N_2015,N_1942);
and U2705 (N_2705,N_2201,N_2011);
xnor U2706 (N_2706,N_2346,N_2144);
or U2707 (N_2707,N_1917,N_2008);
nand U2708 (N_2708,N_2120,N_1954);
or U2709 (N_2709,N_2386,N_1829);
nand U2710 (N_2710,N_2021,N_1934);
and U2711 (N_2711,N_1938,N_1889);
nand U2712 (N_2712,N_2118,N_1815);
xor U2713 (N_2713,N_1855,N_2160);
nand U2714 (N_2714,N_1974,N_2056);
nand U2715 (N_2715,N_1814,N_1958);
nand U2716 (N_2716,N_2340,N_2203);
and U2717 (N_2717,N_2147,N_2281);
nand U2718 (N_2718,N_2203,N_2247);
and U2719 (N_2719,N_1947,N_2134);
nor U2720 (N_2720,N_2076,N_2033);
or U2721 (N_2721,N_2123,N_2334);
nand U2722 (N_2722,N_2392,N_1987);
nand U2723 (N_2723,N_1934,N_2258);
or U2724 (N_2724,N_2106,N_2373);
or U2725 (N_2725,N_2092,N_1901);
or U2726 (N_2726,N_2155,N_1936);
or U2727 (N_2727,N_2129,N_2364);
or U2728 (N_2728,N_2306,N_2212);
nand U2729 (N_2729,N_2271,N_2189);
nor U2730 (N_2730,N_2049,N_2124);
nor U2731 (N_2731,N_2254,N_2120);
xnor U2732 (N_2732,N_2057,N_2259);
nand U2733 (N_2733,N_2377,N_2038);
nor U2734 (N_2734,N_2204,N_2147);
nor U2735 (N_2735,N_1964,N_1855);
nand U2736 (N_2736,N_2324,N_2292);
nor U2737 (N_2737,N_2376,N_1839);
and U2738 (N_2738,N_2327,N_2066);
or U2739 (N_2739,N_2210,N_1988);
and U2740 (N_2740,N_1987,N_2204);
or U2741 (N_2741,N_2327,N_2277);
nand U2742 (N_2742,N_2191,N_2079);
xor U2743 (N_2743,N_1824,N_1935);
xor U2744 (N_2744,N_2155,N_1989);
and U2745 (N_2745,N_1911,N_2023);
xor U2746 (N_2746,N_2235,N_2329);
nor U2747 (N_2747,N_1801,N_2368);
xnor U2748 (N_2748,N_2392,N_2176);
nor U2749 (N_2749,N_1868,N_2009);
nand U2750 (N_2750,N_1926,N_2160);
and U2751 (N_2751,N_2370,N_2285);
xor U2752 (N_2752,N_1968,N_1815);
and U2753 (N_2753,N_1808,N_1890);
or U2754 (N_2754,N_2088,N_1945);
nor U2755 (N_2755,N_2078,N_1906);
nand U2756 (N_2756,N_2031,N_2342);
and U2757 (N_2757,N_2098,N_2177);
and U2758 (N_2758,N_2011,N_1900);
nand U2759 (N_2759,N_2053,N_1862);
nand U2760 (N_2760,N_1825,N_1890);
or U2761 (N_2761,N_2366,N_1908);
or U2762 (N_2762,N_1968,N_1891);
or U2763 (N_2763,N_2169,N_2162);
and U2764 (N_2764,N_2113,N_1895);
and U2765 (N_2765,N_2126,N_2282);
and U2766 (N_2766,N_2236,N_1908);
or U2767 (N_2767,N_1894,N_2296);
or U2768 (N_2768,N_2097,N_2326);
and U2769 (N_2769,N_1891,N_2148);
nand U2770 (N_2770,N_2335,N_2073);
and U2771 (N_2771,N_2089,N_2271);
nand U2772 (N_2772,N_2327,N_1884);
nor U2773 (N_2773,N_2178,N_1954);
nor U2774 (N_2774,N_2338,N_2021);
or U2775 (N_2775,N_2313,N_1899);
nor U2776 (N_2776,N_2040,N_2079);
or U2777 (N_2777,N_2099,N_2278);
nor U2778 (N_2778,N_1869,N_2165);
or U2779 (N_2779,N_2240,N_2393);
and U2780 (N_2780,N_2050,N_2342);
or U2781 (N_2781,N_2212,N_1904);
and U2782 (N_2782,N_2186,N_2201);
and U2783 (N_2783,N_2210,N_2126);
and U2784 (N_2784,N_2320,N_2364);
nor U2785 (N_2785,N_2018,N_1938);
and U2786 (N_2786,N_2021,N_1825);
nor U2787 (N_2787,N_2005,N_2321);
or U2788 (N_2788,N_2340,N_2361);
or U2789 (N_2789,N_1853,N_2087);
nor U2790 (N_2790,N_1824,N_2351);
or U2791 (N_2791,N_1949,N_2197);
nor U2792 (N_2792,N_1943,N_1946);
or U2793 (N_2793,N_2001,N_2119);
nor U2794 (N_2794,N_2050,N_2352);
nand U2795 (N_2795,N_2041,N_2042);
and U2796 (N_2796,N_2265,N_2391);
xnor U2797 (N_2797,N_2104,N_2218);
xor U2798 (N_2798,N_1843,N_1956);
or U2799 (N_2799,N_2083,N_2158);
nand U2800 (N_2800,N_2280,N_1968);
or U2801 (N_2801,N_2383,N_2352);
xnor U2802 (N_2802,N_2390,N_2361);
xnor U2803 (N_2803,N_2253,N_2224);
and U2804 (N_2804,N_1823,N_1938);
xnor U2805 (N_2805,N_2063,N_2089);
nand U2806 (N_2806,N_1908,N_2075);
nor U2807 (N_2807,N_1869,N_2359);
and U2808 (N_2808,N_2365,N_1871);
nor U2809 (N_2809,N_2067,N_1864);
nand U2810 (N_2810,N_1942,N_2345);
xor U2811 (N_2811,N_2209,N_2132);
nor U2812 (N_2812,N_1948,N_2195);
nand U2813 (N_2813,N_1897,N_2257);
nand U2814 (N_2814,N_2022,N_2358);
and U2815 (N_2815,N_1835,N_2233);
or U2816 (N_2816,N_2151,N_1959);
nor U2817 (N_2817,N_2317,N_2116);
nand U2818 (N_2818,N_1852,N_2234);
or U2819 (N_2819,N_2041,N_2373);
nor U2820 (N_2820,N_1900,N_2306);
or U2821 (N_2821,N_1915,N_2113);
nand U2822 (N_2822,N_1958,N_1875);
nand U2823 (N_2823,N_2170,N_2084);
or U2824 (N_2824,N_2383,N_1884);
nor U2825 (N_2825,N_1944,N_2118);
and U2826 (N_2826,N_2200,N_2192);
and U2827 (N_2827,N_1854,N_1943);
or U2828 (N_2828,N_2263,N_1976);
nand U2829 (N_2829,N_1913,N_1910);
xor U2830 (N_2830,N_1825,N_2016);
nand U2831 (N_2831,N_2380,N_2350);
nor U2832 (N_2832,N_2277,N_1828);
and U2833 (N_2833,N_1846,N_2315);
nor U2834 (N_2834,N_1969,N_1946);
nand U2835 (N_2835,N_1872,N_2172);
and U2836 (N_2836,N_1922,N_1982);
nor U2837 (N_2837,N_2168,N_2349);
xnor U2838 (N_2838,N_2149,N_2239);
nor U2839 (N_2839,N_2012,N_2383);
nand U2840 (N_2840,N_2134,N_2140);
and U2841 (N_2841,N_2141,N_2254);
xor U2842 (N_2842,N_1935,N_2032);
nand U2843 (N_2843,N_2319,N_2206);
or U2844 (N_2844,N_1805,N_2237);
and U2845 (N_2845,N_2238,N_1978);
xor U2846 (N_2846,N_1826,N_2023);
nand U2847 (N_2847,N_2282,N_2199);
nand U2848 (N_2848,N_1832,N_1929);
nand U2849 (N_2849,N_1958,N_1941);
nor U2850 (N_2850,N_2073,N_2091);
and U2851 (N_2851,N_2242,N_1999);
and U2852 (N_2852,N_2002,N_1960);
nand U2853 (N_2853,N_2327,N_2231);
nand U2854 (N_2854,N_1885,N_1830);
nor U2855 (N_2855,N_2217,N_2102);
nor U2856 (N_2856,N_2176,N_1959);
or U2857 (N_2857,N_2295,N_1961);
nor U2858 (N_2858,N_2097,N_2183);
or U2859 (N_2859,N_1812,N_1980);
nand U2860 (N_2860,N_2326,N_2045);
or U2861 (N_2861,N_2284,N_2366);
and U2862 (N_2862,N_2247,N_1821);
and U2863 (N_2863,N_2399,N_1978);
nand U2864 (N_2864,N_2353,N_1945);
or U2865 (N_2865,N_2197,N_2318);
or U2866 (N_2866,N_2118,N_2256);
and U2867 (N_2867,N_1960,N_2088);
and U2868 (N_2868,N_2246,N_2285);
nand U2869 (N_2869,N_1924,N_2200);
or U2870 (N_2870,N_1857,N_2192);
and U2871 (N_2871,N_2171,N_2097);
nand U2872 (N_2872,N_2347,N_2085);
nor U2873 (N_2873,N_1808,N_1955);
or U2874 (N_2874,N_1806,N_2335);
nor U2875 (N_2875,N_2127,N_2251);
and U2876 (N_2876,N_2338,N_1827);
and U2877 (N_2877,N_2377,N_1932);
nor U2878 (N_2878,N_2132,N_1971);
and U2879 (N_2879,N_1927,N_2016);
and U2880 (N_2880,N_1843,N_2249);
nor U2881 (N_2881,N_2203,N_2284);
or U2882 (N_2882,N_1917,N_1889);
nand U2883 (N_2883,N_2323,N_1963);
nand U2884 (N_2884,N_2226,N_2277);
and U2885 (N_2885,N_2333,N_1850);
nand U2886 (N_2886,N_2302,N_2094);
nand U2887 (N_2887,N_1827,N_1949);
nor U2888 (N_2888,N_2040,N_1890);
nand U2889 (N_2889,N_2338,N_2059);
nor U2890 (N_2890,N_2018,N_2042);
nor U2891 (N_2891,N_1928,N_2067);
nor U2892 (N_2892,N_1874,N_1897);
and U2893 (N_2893,N_1951,N_2271);
and U2894 (N_2894,N_1996,N_1951);
or U2895 (N_2895,N_2365,N_2346);
or U2896 (N_2896,N_2245,N_1919);
nor U2897 (N_2897,N_2057,N_2014);
and U2898 (N_2898,N_1876,N_2366);
and U2899 (N_2899,N_2317,N_2324);
and U2900 (N_2900,N_1846,N_2060);
or U2901 (N_2901,N_1995,N_2227);
nand U2902 (N_2902,N_1979,N_1807);
and U2903 (N_2903,N_1934,N_1846);
nor U2904 (N_2904,N_2086,N_2023);
or U2905 (N_2905,N_1992,N_2104);
xor U2906 (N_2906,N_2047,N_1838);
and U2907 (N_2907,N_2154,N_1971);
or U2908 (N_2908,N_1870,N_2056);
and U2909 (N_2909,N_2303,N_2358);
nand U2910 (N_2910,N_2226,N_2122);
nor U2911 (N_2911,N_1819,N_2276);
nor U2912 (N_2912,N_2349,N_1815);
and U2913 (N_2913,N_2112,N_1843);
nand U2914 (N_2914,N_2322,N_2396);
or U2915 (N_2915,N_2190,N_1989);
nand U2916 (N_2916,N_2142,N_1899);
or U2917 (N_2917,N_1909,N_2108);
or U2918 (N_2918,N_2109,N_2304);
nand U2919 (N_2919,N_1868,N_2140);
nand U2920 (N_2920,N_2008,N_2221);
nor U2921 (N_2921,N_1922,N_2368);
nand U2922 (N_2922,N_1945,N_2038);
nor U2923 (N_2923,N_2054,N_1964);
or U2924 (N_2924,N_2256,N_1938);
and U2925 (N_2925,N_1989,N_2177);
nand U2926 (N_2926,N_2396,N_1997);
nand U2927 (N_2927,N_2299,N_2249);
nor U2928 (N_2928,N_1953,N_2096);
nand U2929 (N_2929,N_2221,N_2114);
and U2930 (N_2930,N_2163,N_2260);
nand U2931 (N_2931,N_2334,N_2140);
nor U2932 (N_2932,N_2336,N_1833);
xor U2933 (N_2933,N_2138,N_2204);
nand U2934 (N_2934,N_2315,N_2150);
xor U2935 (N_2935,N_2247,N_2276);
nand U2936 (N_2936,N_1984,N_1931);
nor U2937 (N_2937,N_2186,N_2034);
nand U2938 (N_2938,N_2300,N_2064);
nand U2939 (N_2939,N_1981,N_2273);
or U2940 (N_2940,N_2132,N_1957);
nand U2941 (N_2941,N_2080,N_1842);
and U2942 (N_2942,N_2162,N_2237);
nor U2943 (N_2943,N_1863,N_2272);
or U2944 (N_2944,N_2318,N_1873);
nand U2945 (N_2945,N_2018,N_2225);
nor U2946 (N_2946,N_2395,N_1987);
and U2947 (N_2947,N_1858,N_1833);
or U2948 (N_2948,N_2206,N_1889);
nor U2949 (N_2949,N_2397,N_2237);
nor U2950 (N_2950,N_2109,N_2341);
nor U2951 (N_2951,N_1846,N_2026);
or U2952 (N_2952,N_2009,N_1922);
or U2953 (N_2953,N_2316,N_2266);
and U2954 (N_2954,N_2215,N_2038);
nor U2955 (N_2955,N_2102,N_2103);
nor U2956 (N_2956,N_2314,N_1831);
and U2957 (N_2957,N_2114,N_2162);
xnor U2958 (N_2958,N_1810,N_2294);
xor U2959 (N_2959,N_2156,N_2173);
and U2960 (N_2960,N_2292,N_2060);
and U2961 (N_2961,N_1819,N_2016);
or U2962 (N_2962,N_2354,N_1830);
and U2963 (N_2963,N_1997,N_1901);
and U2964 (N_2964,N_1946,N_2060);
and U2965 (N_2965,N_1998,N_2103);
or U2966 (N_2966,N_2216,N_2127);
nor U2967 (N_2967,N_2305,N_1996);
nor U2968 (N_2968,N_2058,N_1880);
nand U2969 (N_2969,N_2120,N_2156);
or U2970 (N_2970,N_1984,N_1800);
and U2971 (N_2971,N_2224,N_1981);
nor U2972 (N_2972,N_1930,N_2371);
or U2973 (N_2973,N_1876,N_2205);
nand U2974 (N_2974,N_2292,N_2005);
and U2975 (N_2975,N_2227,N_2257);
and U2976 (N_2976,N_2284,N_2224);
nor U2977 (N_2977,N_2284,N_2042);
or U2978 (N_2978,N_1979,N_1929);
and U2979 (N_2979,N_1818,N_1864);
and U2980 (N_2980,N_1877,N_2236);
nand U2981 (N_2981,N_2357,N_1817);
or U2982 (N_2982,N_2260,N_2223);
or U2983 (N_2983,N_2326,N_2276);
nor U2984 (N_2984,N_1844,N_2378);
and U2985 (N_2985,N_2066,N_2057);
or U2986 (N_2986,N_2127,N_1952);
nand U2987 (N_2987,N_2031,N_2049);
and U2988 (N_2988,N_2085,N_1893);
nor U2989 (N_2989,N_1919,N_1855);
xor U2990 (N_2990,N_1843,N_2149);
xor U2991 (N_2991,N_1826,N_2169);
or U2992 (N_2992,N_2070,N_2364);
or U2993 (N_2993,N_2118,N_1943);
nor U2994 (N_2994,N_1899,N_1903);
nand U2995 (N_2995,N_1898,N_1967);
or U2996 (N_2996,N_2220,N_2015);
nor U2997 (N_2997,N_2094,N_2081);
or U2998 (N_2998,N_2372,N_1946);
nand U2999 (N_2999,N_2142,N_2208);
nor U3000 (N_3000,N_2437,N_2893);
nor U3001 (N_3001,N_2837,N_2551);
nor U3002 (N_3002,N_2601,N_2883);
and U3003 (N_3003,N_2629,N_2713);
or U3004 (N_3004,N_2895,N_2412);
nor U3005 (N_3005,N_2990,N_2591);
or U3006 (N_3006,N_2825,N_2832);
nand U3007 (N_3007,N_2593,N_2946);
or U3008 (N_3008,N_2435,N_2670);
or U3009 (N_3009,N_2821,N_2633);
nor U3010 (N_3010,N_2902,N_2568);
nor U3011 (N_3011,N_2456,N_2449);
xor U3012 (N_3012,N_2698,N_2522);
or U3013 (N_3013,N_2903,N_2636);
or U3014 (N_3014,N_2779,N_2729);
or U3015 (N_3015,N_2726,N_2656);
nand U3016 (N_3016,N_2776,N_2661);
nor U3017 (N_3017,N_2637,N_2972);
or U3018 (N_3018,N_2938,N_2860);
nand U3019 (N_3019,N_2823,N_2847);
nor U3020 (N_3020,N_2735,N_2703);
nand U3021 (N_3021,N_2557,N_2662);
and U3022 (N_3022,N_2487,N_2442);
or U3023 (N_3023,N_2801,N_2748);
nor U3024 (N_3024,N_2686,N_2548);
nand U3025 (N_3025,N_2966,N_2813);
or U3026 (N_3026,N_2669,N_2410);
or U3027 (N_3027,N_2616,N_2898);
and U3028 (N_3028,N_2417,N_2798);
nand U3029 (N_3029,N_2599,N_2500);
nor U3030 (N_3030,N_2645,N_2411);
or U3031 (N_3031,N_2790,N_2434);
nand U3032 (N_3032,N_2960,N_2916);
or U3033 (N_3033,N_2414,N_2931);
and U3034 (N_3034,N_2588,N_2774);
xnor U3035 (N_3035,N_2885,N_2788);
and U3036 (N_3036,N_2524,N_2852);
or U3037 (N_3037,N_2759,N_2705);
nor U3038 (N_3038,N_2582,N_2905);
and U3039 (N_3039,N_2841,N_2419);
and U3040 (N_3040,N_2767,N_2867);
or U3041 (N_3041,N_2746,N_2976);
nand U3042 (N_3042,N_2514,N_2809);
nor U3043 (N_3043,N_2802,N_2477);
nor U3044 (N_3044,N_2440,N_2708);
nor U3045 (N_3045,N_2423,N_2653);
nand U3046 (N_3046,N_2448,N_2738);
nor U3047 (N_3047,N_2592,N_2888);
xor U3048 (N_3048,N_2935,N_2877);
or U3049 (N_3049,N_2838,N_2531);
and U3050 (N_3050,N_2534,N_2589);
nand U3051 (N_3051,N_2754,N_2875);
nand U3052 (N_3052,N_2554,N_2818);
nor U3053 (N_3053,N_2753,N_2536);
and U3054 (N_3054,N_2913,N_2612);
and U3055 (N_3055,N_2615,N_2929);
nor U3056 (N_3056,N_2547,N_2822);
and U3057 (N_3057,N_2780,N_2783);
nand U3058 (N_3058,N_2680,N_2855);
and U3059 (N_3059,N_2947,N_2701);
and U3060 (N_3060,N_2733,N_2720);
and U3061 (N_3061,N_2585,N_2829);
or U3062 (N_3062,N_2626,N_2652);
nor U3063 (N_3063,N_2850,N_2846);
or U3064 (N_3064,N_2493,N_2743);
xor U3065 (N_3065,N_2803,N_2925);
or U3066 (N_3066,N_2725,N_2486);
or U3067 (N_3067,N_2769,N_2559);
or U3068 (N_3068,N_2770,N_2807);
and U3069 (N_3069,N_2512,N_2498);
xor U3070 (N_3070,N_2576,N_2664);
nor U3071 (N_3071,N_2580,N_2900);
xnor U3072 (N_3072,N_2539,N_2438);
or U3073 (N_3073,N_2810,N_2861);
nor U3074 (N_3074,N_2622,N_2630);
nand U3075 (N_3075,N_2673,N_2899);
nor U3076 (N_3076,N_2518,N_2749);
nor U3077 (N_3077,N_2842,N_2492);
or U3078 (N_3078,N_2640,N_2918);
nor U3079 (N_3079,N_2692,N_2517);
and U3080 (N_3080,N_2716,N_2922);
nand U3081 (N_3081,N_2714,N_2556);
nor U3082 (N_3082,N_2892,N_2679);
nor U3083 (N_3083,N_2856,N_2942);
or U3084 (N_3084,N_2695,N_2975);
nor U3085 (N_3085,N_2526,N_2717);
and U3086 (N_3086,N_2934,N_2873);
nor U3087 (N_3087,N_2843,N_2808);
nor U3088 (N_3088,N_2660,N_2994);
and U3089 (N_3089,N_2933,N_2866);
nor U3090 (N_3090,N_2451,N_2572);
nand U3091 (N_3091,N_2455,N_2891);
nor U3092 (N_3092,N_2654,N_2468);
nor U3093 (N_3093,N_2608,N_2944);
and U3094 (N_3094,N_2422,N_2949);
or U3095 (N_3095,N_2583,N_2722);
nand U3096 (N_3096,N_2404,N_2605);
and U3097 (N_3097,N_2447,N_2416);
or U3098 (N_3098,N_2858,N_2687);
and U3099 (N_3099,N_2594,N_2503);
and U3100 (N_3100,N_2986,N_2804);
or U3101 (N_3101,N_2479,N_2621);
or U3102 (N_3102,N_2688,N_2550);
or U3103 (N_3103,N_2833,N_2967);
nor U3104 (N_3104,N_2870,N_2491);
nor U3105 (N_3105,N_2765,N_2740);
nand U3106 (N_3106,N_2771,N_2567);
nor U3107 (N_3107,N_2489,N_2955);
or U3108 (N_3108,N_2405,N_2509);
and U3109 (N_3109,N_2980,N_2979);
or U3110 (N_3110,N_2627,N_2655);
xor U3111 (N_3111,N_2865,N_2459);
xnor U3112 (N_3112,N_2785,N_2791);
or U3113 (N_3113,N_2834,N_2415);
and U3114 (N_3114,N_2964,N_2831);
nand U3115 (N_3115,N_2483,N_2881);
nand U3116 (N_3116,N_2816,N_2909);
nand U3117 (N_3117,N_2777,N_2401);
nor U3118 (N_3118,N_2794,N_2712);
nor U3119 (N_3119,N_2768,N_2425);
nor U3120 (N_3120,N_2677,N_2930);
nand U3121 (N_3121,N_2824,N_2982);
and U3122 (N_3122,N_2577,N_2667);
xnor U3123 (N_3123,N_2528,N_2869);
nor U3124 (N_3124,N_2786,N_2525);
nand U3125 (N_3125,N_2797,N_2619);
and U3126 (N_3126,N_2646,N_2886);
nor U3127 (N_3127,N_2689,N_2795);
nor U3128 (N_3128,N_2732,N_2436);
nand U3129 (N_3129,N_2443,N_2945);
or U3130 (N_3130,N_2812,N_2610);
xnor U3131 (N_3131,N_2475,N_2995);
and U3132 (N_3132,N_2672,N_2523);
nor U3133 (N_3133,N_2978,N_2623);
and U3134 (N_3134,N_2649,N_2723);
or U3135 (N_3135,N_2403,N_2991);
and U3136 (N_3136,N_2853,N_2527);
or U3137 (N_3137,N_2697,N_2839);
and U3138 (N_3138,N_2647,N_2541);
or U3139 (N_3139,N_2682,N_2474);
nand U3140 (N_3140,N_2683,N_2472);
or U3141 (N_3141,N_2710,N_2533);
or U3142 (N_3142,N_2755,N_2575);
nand U3143 (N_3143,N_2868,N_2745);
nor U3144 (N_3144,N_2537,N_2985);
nand U3145 (N_3145,N_2782,N_2956);
and U3146 (N_3146,N_2872,N_2932);
and U3147 (N_3147,N_2494,N_2439);
or U3148 (N_3148,N_2943,N_2917);
nor U3149 (N_3149,N_2773,N_2819);
or U3150 (N_3150,N_2502,N_2927);
or U3151 (N_3151,N_2634,N_2458);
nand U3152 (N_3152,N_2406,N_2958);
nor U3153 (N_3153,N_2566,N_2454);
nand U3154 (N_3154,N_2461,N_2507);
or U3155 (N_3155,N_2573,N_2457);
or U3156 (N_3156,N_2614,N_2618);
or U3157 (N_3157,N_2400,N_2959);
and U3158 (N_3158,N_2569,N_2988);
or U3159 (N_3159,N_2894,N_2989);
or U3160 (N_3160,N_2420,N_2815);
nand U3161 (N_3161,N_2999,N_2445);
or U3162 (N_3162,N_2481,N_2828);
nand U3163 (N_3163,N_2879,N_2515);
nand U3164 (N_3164,N_2957,N_2484);
nor U3165 (N_3165,N_2639,N_2665);
nor U3166 (N_3166,N_2793,N_2657);
and U3167 (N_3167,N_2620,N_2545);
and U3168 (N_3168,N_2981,N_2742);
and U3169 (N_3169,N_2826,N_2787);
or U3170 (N_3170,N_2625,N_2516);
nor U3171 (N_3171,N_2501,N_2952);
and U3172 (N_3172,N_2659,N_2542);
or U3173 (N_3173,N_2805,N_2650);
xnor U3174 (N_3174,N_2549,N_2921);
and U3175 (N_3175,N_2876,N_2467);
nor U3176 (N_3176,N_2889,N_2453);
nand U3177 (N_3177,N_2587,N_2799);
nand U3178 (N_3178,N_2737,N_2977);
or U3179 (N_3179,N_2408,N_2854);
or U3180 (N_3180,N_2444,N_2506);
or U3181 (N_3181,N_2996,N_2685);
and U3182 (N_3182,N_2983,N_2693);
nand U3183 (N_3183,N_2718,N_2878);
nor U3184 (N_3184,N_2520,N_2584);
nand U3185 (N_3185,N_2721,N_2750);
xnor U3186 (N_3186,N_2963,N_2544);
nand U3187 (N_3187,N_2849,N_2789);
xnor U3188 (N_3188,N_2702,N_2606);
and U3189 (N_3189,N_2497,N_2597);
or U3190 (N_3190,N_2904,N_2464);
and U3191 (N_3191,N_2914,N_2936);
or U3192 (N_3192,N_2574,N_2998);
nand U3193 (N_3193,N_2758,N_2845);
and U3194 (N_3194,N_2951,N_2954);
nor U3195 (N_3195,N_2603,N_2806);
or U3196 (N_3196,N_2736,N_2910);
xnor U3197 (N_3197,N_2560,N_2920);
nand U3198 (N_3198,N_2562,N_2864);
nand U3199 (N_3199,N_2632,N_2476);
nand U3200 (N_3200,N_2540,N_2744);
and U3201 (N_3201,N_2973,N_2643);
nand U3202 (N_3202,N_2923,N_2519);
nand U3203 (N_3203,N_2604,N_2613);
xor U3204 (N_3204,N_2496,N_2402);
and U3205 (N_3205,N_2666,N_2811);
and U3206 (N_3206,N_2432,N_2413);
nand U3207 (N_3207,N_2800,N_2752);
nand U3208 (N_3208,N_2836,N_2901);
nand U3209 (N_3209,N_2485,N_2939);
and U3210 (N_3210,N_2874,N_2747);
nand U3211 (N_3211,N_2535,N_2529);
nor U3212 (N_3212,N_2510,N_2764);
and U3213 (N_3213,N_2595,N_2792);
and U3214 (N_3214,N_2907,N_2546);
or U3215 (N_3215,N_2511,N_2678);
nand U3216 (N_3216,N_2579,N_2840);
and U3217 (N_3217,N_2429,N_2424);
and U3218 (N_3218,N_2694,N_2763);
nand U3219 (N_3219,N_2407,N_2696);
or U3220 (N_3220,N_2641,N_2699);
nor U3221 (N_3221,N_2863,N_2638);
nand U3222 (N_3222,N_2598,N_2658);
and U3223 (N_3223,N_2814,N_2882);
nand U3224 (N_3224,N_2897,N_2940);
or U3225 (N_3225,N_2928,N_2706);
or U3226 (N_3226,N_2426,N_2480);
or U3227 (N_3227,N_2428,N_2766);
nand U3228 (N_3228,N_2961,N_2478);
or U3229 (N_3229,N_2607,N_2441);
or U3230 (N_3230,N_2731,N_2887);
xnor U3231 (N_3231,N_2851,N_2611);
or U3232 (N_3232,N_2564,N_2926);
nor U3233 (N_3233,N_2908,N_2896);
xnor U3234 (N_3234,N_2704,N_2473);
nand U3235 (N_3235,N_2884,N_2796);
nor U3236 (N_3236,N_2993,N_2739);
xnor U3237 (N_3237,N_2675,N_2727);
nor U3238 (N_3238,N_2997,N_2602);
or U3239 (N_3239,N_2586,N_2471);
and U3240 (N_3240,N_2446,N_2499);
and U3241 (N_3241,N_2969,N_2470);
or U3242 (N_3242,N_2827,N_2561);
nor U3243 (N_3243,N_2962,N_2671);
or U3244 (N_3244,N_2430,N_2906);
or U3245 (N_3245,N_2674,N_2950);
nand U3246 (N_3246,N_2600,N_2642);
nand U3247 (N_3247,N_2970,N_2691);
nand U3248 (N_3248,N_2711,N_2609);
or U3249 (N_3249,N_2558,N_2684);
and U3250 (N_3250,N_2505,N_2450);
xor U3251 (N_3251,N_2715,N_2974);
nand U3252 (N_3252,N_2830,N_2543);
or U3253 (N_3253,N_2948,N_2761);
nand U3254 (N_3254,N_2760,N_2463);
nor U3255 (N_3255,N_2762,N_2775);
and U3256 (N_3256,N_2987,N_2552);
nor U3257 (N_3257,N_2427,N_2984);
and U3258 (N_3258,N_2668,N_2571);
and U3259 (N_3259,N_2912,N_2488);
or U3260 (N_3260,N_2521,N_2418);
nor U3261 (N_3261,N_2757,N_2971);
nor U3262 (N_3262,N_2663,N_2578);
nand U3263 (N_3263,N_2465,N_2469);
or U3264 (N_3264,N_2452,N_2532);
xnor U3265 (N_3265,N_2690,N_2538);
nor U3266 (N_3266,N_2915,N_2624);
nor U3267 (N_3267,N_2462,N_2857);
or U3268 (N_3268,N_2859,N_2992);
and U3269 (N_3269,N_2635,N_2756);
and U3270 (N_3270,N_2965,N_2741);
nand U3271 (N_3271,N_2504,N_2553);
nand U3272 (N_3272,N_2631,N_2707);
nor U3273 (N_3273,N_2482,N_2565);
and U3274 (N_3274,N_2937,N_2570);
or U3275 (N_3275,N_2772,N_2433);
or U3276 (N_3276,N_2719,N_2513);
and U3277 (N_3277,N_2644,N_2835);
or U3278 (N_3278,N_2941,N_2778);
and U3279 (N_3279,N_2890,N_2848);
and U3280 (N_3280,N_2490,N_2911);
or U3281 (N_3281,N_2862,N_2628);
nor U3282 (N_3282,N_2676,N_2880);
nor U3283 (N_3283,N_2953,N_2409);
nand U3284 (N_3284,N_2590,N_2555);
xor U3285 (N_3285,N_2700,N_2844);
or U3286 (N_3286,N_2781,N_2919);
nand U3287 (N_3287,N_2596,N_2495);
and U3288 (N_3288,N_2751,N_2421);
nor U3289 (N_3289,N_2460,N_2581);
and U3290 (N_3290,N_2681,N_2431);
nand U3291 (N_3291,N_2728,N_2648);
and U3292 (N_3292,N_2530,N_2709);
nand U3293 (N_3293,N_2820,N_2924);
nor U3294 (N_3294,N_2724,N_2784);
nand U3295 (N_3295,N_2871,N_2651);
or U3296 (N_3296,N_2817,N_2508);
and U3297 (N_3297,N_2563,N_2730);
and U3298 (N_3298,N_2617,N_2734);
and U3299 (N_3299,N_2466,N_2968);
or U3300 (N_3300,N_2982,N_2823);
and U3301 (N_3301,N_2687,N_2425);
and U3302 (N_3302,N_2956,N_2517);
or U3303 (N_3303,N_2781,N_2514);
xnor U3304 (N_3304,N_2807,N_2583);
nor U3305 (N_3305,N_2815,N_2964);
nor U3306 (N_3306,N_2887,N_2853);
and U3307 (N_3307,N_2518,N_2706);
nor U3308 (N_3308,N_2951,N_2871);
nor U3309 (N_3309,N_2935,N_2539);
nand U3310 (N_3310,N_2805,N_2926);
or U3311 (N_3311,N_2963,N_2436);
nand U3312 (N_3312,N_2736,N_2815);
or U3313 (N_3313,N_2482,N_2595);
nor U3314 (N_3314,N_2755,N_2693);
or U3315 (N_3315,N_2847,N_2876);
or U3316 (N_3316,N_2728,N_2581);
and U3317 (N_3317,N_2430,N_2805);
or U3318 (N_3318,N_2937,N_2406);
nand U3319 (N_3319,N_2697,N_2745);
or U3320 (N_3320,N_2890,N_2655);
and U3321 (N_3321,N_2943,N_2432);
nand U3322 (N_3322,N_2753,N_2960);
nand U3323 (N_3323,N_2531,N_2424);
nor U3324 (N_3324,N_2728,N_2789);
nor U3325 (N_3325,N_2448,N_2943);
or U3326 (N_3326,N_2796,N_2595);
nand U3327 (N_3327,N_2593,N_2834);
nor U3328 (N_3328,N_2755,N_2510);
or U3329 (N_3329,N_2955,N_2844);
and U3330 (N_3330,N_2710,N_2639);
xor U3331 (N_3331,N_2725,N_2850);
nand U3332 (N_3332,N_2501,N_2979);
and U3333 (N_3333,N_2655,N_2932);
nor U3334 (N_3334,N_2868,N_2448);
xor U3335 (N_3335,N_2598,N_2851);
or U3336 (N_3336,N_2464,N_2712);
or U3337 (N_3337,N_2578,N_2438);
and U3338 (N_3338,N_2977,N_2492);
or U3339 (N_3339,N_2594,N_2470);
or U3340 (N_3340,N_2513,N_2617);
and U3341 (N_3341,N_2497,N_2942);
nor U3342 (N_3342,N_2468,N_2756);
and U3343 (N_3343,N_2911,N_2882);
and U3344 (N_3344,N_2973,N_2478);
nor U3345 (N_3345,N_2913,N_2591);
or U3346 (N_3346,N_2809,N_2440);
nor U3347 (N_3347,N_2544,N_2907);
nor U3348 (N_3348,N_2483,N_2691);
or U3349 (N_3349,N_2750,N_2508);
nand U3350 (N_3350,N_2737,N_2658);
nand U3351 (N_3351,N_2424,N_2833);
nand U3352 (N_3352,N_2518,N_2583);
nand U3353 (N_3353,N_2894,N_2911);
xnor U3354 (N_3354,N_2917,N_2520);
xor U3355 (N_3355,N_2844,N_2428);
xor U3356 (N_3356,N_2425,N_2559);
or U3357 (N_3357,N_2447,N_2487);
nor U3358 (N_3358,N_2840,N_2542);
or U3359 (N_3359,N_2537,N_2445);
or U3360 (N_3360,N_2856,N_2844);
or U3361 (N_3361,N_2476,N_2747);
or U3362 (N_3362,N_2453,N_2839);
nor U3363 (N_3363,N_2545,N_2499);
nor U3364 (N_3364,N_2848,N_2952);
nand U3365 (N_3365,N_2970,N_2784);
and U3366 (N_3366,N_2892,N_2402);
or U3367 (N_3367,N_2561,N_2686);
nor U3368 (N_3368,N_2576,N_2428);
nand U3369 (N_3369,N_2894,N_2667);
xnor U3370 (N_3370,N_2485,N_2907);
xnor U3371 (N_3371,N_2549,N_2715);
and U3372 (N_3372,N_2634,N_2994);
nor U3373 (N_3373,N_2476,N_2448);
nor U3374 (N_3374,N_2985,N_2782);
nor U3375 (N_3375,N_2819,N_2829);
nand U3376 (N_3376,N_2962,N_2852);
nand U3377 (N_3377,N_2803,N_2574);
nor U3378 (N_3378,N_2718,N_2918);
nor U3379 (N_3379,N_2827,N_2612);
or U3380 (N_3380,N_2550,N_2572);
nand U3381 (N_3381,N_2645,N_2706);
or U3382 (N_3382,N_2952,N_2448);
nand U3383 (N_3383,N_2767,N_2737);
xor U3384 (N_3384,N_2717,N_2504);
xor U3385 (N_3385,N_2640,N_2509);
or U3386 (N_3386,N_2654,N_2819);
or U3387 (N_3387,N_2461,N_2457);
nand U3388 (N_3388,N_2780,N_2952);
and U3389 (N_3389,N_2682,N_2405);
nand U3390 (N_3390,N_2661,N_2612);
nand U3391 (N_3391,N_2692,N_2998);
and U3392 (N_3392,N_2627,N_2794);
and U3393 (N_3393,N_2442,N_2577);
or U3394 (N_3394,N_2918,N_2584);
nor U3395 (N_3395,N_2919,N_2701);
nor U3396 (N_3396,N_2755,N_2934);
or U3397 (N_3397,N_2959,N_2922);
nand U3398 (N_3398,N_2590,N_2912);
and U3399 (N_3399,N_2715,N_2812);
nand U3400 (N_3400,N_2987,N_2685);
xnor U3401 (N_3401,N_2962,N_2846);
and U3402 (N_3402,N_2541,N_2457);
nor U3403 (N_3403,N_2810,N_2719);
nand U3404 (N_3404,N_2578,N_2636);
nand U3405 (N_3405,N_2752,N_2433);
xor U3406 (N_3406,N_2914,N_2748);
nor U3407 (N_3407,N_2842,N_2713);
nand U3408 (N_3408,N_2447,N_2525);
nand U3409 (N_3409,N_2536,N_2632);
and U3410 (N_3410,N_2597,N_2650);
and U3411 (N_3411,N_2581,N_2992);
and U3412 (N_3412,N_2737,N_2773);
and U3413 (N_3413,N_2543,N_2982);
nor U3414 (N_3414,N_2762,N_2709);
and U3415 (N_3415,N_2918,N_2962);
and U3416 (N_3416,N_2786,N_2841);
or U3417 (N_3417,N_2964,N_2892);
xnor U3418 (N_3418,N_2770,N_2733);
nor U3419 (N_3419,N_2879,N_2756);
or U3420 (N_3420,N_2848,N_2911);
and U3421 (N_3421,N_2497,N_2825);
nand U3422 (N_3422,N_2413,N_2509);
nand U3423 (N_3423,N_2993,N_2990);
nor U3424 (N_3424,N_2634,N_2954);
and U3425 (N_3425,N_2753,N_2761);
nand U3426 (N_3426,N_2631,N_2734);
and U3427 (N_3427,N_2756,N_2434);
or U3428 (N_3428,N_2828,N_2408);
and U3429 (N_3429,N_2723,N_2909);
nand U3430 (N_3430,N_2852,N_2973);
nor U3431 (N_3431,N_2976,N_2979);
or U3432 (N_3432,N_2969,N_2895);
or U3433 (N_3433,N_2568,N_2912);
and U3434 (N_3434,N_2982,N_2531);
or U3435 (N_3435,N_2632,N_2498);
and U3436 (N_3436,N_2633,N_2917);
or U3437 (N_3437,N_2431,N_2723);
and U3438 (N_3438,N_2411,N_2806);
or U3439 (N_3439,N_2739,N_2792);
and U3440 (N_3440,N_2963,N_2872);
nand U3441 (N_3441,N_2802,N_2686);
nor U3442 (N_3442,N_2590,N_2596);
and U3443 (N_3443,N_2753,N_2500);
or U3444 (N_3444,N_2575,N_2808);
nand U3445 (N_3445,N_2820,N_2886);
xor U3446 (N_3446,N_2835,N_2906);
nand U3447 (N_3447,N_2883,N_2698);
and U3448 (N_3448,N_2615,N_2644);
nor U3449 (N_3449,N_2527,N_2966);
or U3450 (N_3450,N_2751,N_2499);
nand U3451 (N_3451,N_2678,N_2418);
and U3452 (N_3452,N_2957,N_2969);
and U3453 (N_3453,N_2979,N_2426);
and U3454 (N_3454,N_2432,N_2810);
or U3455 (N_3455,N_2551,N_2405);
nand U3456 (N_3456,N_2945,N_2984);
nand U3457 (N_3457,N_2415,N_2663);
xnor U3458 (N_3458,N_2585,N_2522);
nor U3459 (N_3459,N_2584,N_2940);
nand U3460 (N_3460,N_2807,N_2494);
or U3461 (N_3461,N_2526,N_2708);
nand U3462 (N_3462,N_2532,N_2688);
nand U3463 (N_3463,N_2825,N_2968);
nor U3464 (N_3464,N_2550,N_2902);
and U3465 (N_3465,N_2787,N_2588);
nor U3466 (N_3466,N_2734,N_2771);
nand U3467 (N_3467,N_2520,N_2958);
nand U3468 (N_3468,N_2715,N_2941);
nor U3469 (N_3469,N_2886,N_2813);
or U3470 (N_3470,N_2887,N_2695);
nand U3471 (N_3471,N_2468,N_2747);
or U3472 (N_3472,N_2753,N_2999);
and U3473 (N_3473,N_2527,N_2631);
and U3474 (N_3474,N_2818,N_2463);
nand U3475 (N_3475,N_2540,N_2940);
nand U3476 (N_3476,N_2698,N_2995);
or U3477 (N_3477,N_2860,N_2482);
nor U3478 (N_3478,N_2984,N_2493);
nor U3479 (N_3479,N_2768,N_2758);
and U3480 (N_3480,N_2939,N_2804);
nor U3481 (N_3481,N_2749,N_2733);
or U3482 (N_3482,N_2847,N_2685);
nor U3483 (N_3483,N_2419,N_2822);
xnor U3484 (N_3484,N_2945,N_2839);
and U3485 (N_3485,N_2886,N_2756);
and U3486 (N_3486,N_2756,N_2690);
or U3487 (N_3487,N_2932,N_2968);
nand U3488 (N_3488,N_2819,N_2810);
or U3489 (N_3489,N_2678,N_2504);
xor U3490 (N_3490,N_2525,N_2421);
nand U3491 (N_3491,N_2482,N_2666);
nor U3492 (N_3492,N_2808,N_2448);
and U3493 (N_3493,N_2883,N_2514);
or U3494 (N_3494,N_2499,N_2869);
nor U3495 (N_3495,N_2489,N_2427);
or U3496 (N_3496,N_2808,N_2785);
xor U3497 (N_3497,N_2588,N_2616);
and U3498 (N_3498,N_2531,N_2536);
or U3499 (N_3499,N_2590,N_2469);
nor U3500 (N_3500,N_2674,N_2851);
nand U3501 (N_3501,N_2937,N_2740);
and U3502 (N_3502,N_2454,N_2955);
and U3503 (N_3503,N_2978,N_2488);
or U3504 (N_3504,N_2564,N_2773);
nor U3505 (N_3505,N_2611,N_2919);
nand U3506 (N_3506,N_2675,N_2833);
and U3507 (N_3507,N_2418,N_2570);
nor U3508 (N_3508,N_2987,N_2768);
nor U3509 (N_3509,N_2655,N_2521);
nand U3510 (N_3510,N_2985,N_2792);
xnor U3511 (N_3511,N_2637,N_2570);
and U3512 (N_3512,N_2792,N_2879);
nand U3513 (N_3513,N_2796,N_2660);
and U3514 (N_3514,N_2975,N_2607);
and U3515 (N_3515,N_2404,N_2490);
nor U3516 (N_3516,N_2578,N_2715);
nand U3517 (N_3517,N_2400,N_2800);
and U3518 (N_3518,N_2788,N_2418);
and U3519 (N_3519,N_2695,N_2413);
nand U3520 (N_3520,N_2462,N_2756);
nor U3521 (N_3521,N_2884,N_2442);
and U3522 (N_3522,N_2441,N_2700);
and U3523 (N_3523,N_2845,N_2449);
nand U3524 (N_3524,N_2589,N_2505);
and U3525 (N_3525,N_2841,N_2740);
nor U3526 (N_3526,N_2402,N_2540);
or U3527 (N_3527,N_2784,N_2697);
nand U3528 (N_3528,N_2624,N_2473);
or U3529 (N_3529,N_2431,N_2874);
nand U3530 (N_3530,N_2561,N_2639);
and U3531 (N_3531,N_2621,N_2750);
nor U3532 (N_3532,N_2758,N_2963);
nand U3533 (N_3533,N_2810,N_2456);
or U3534 (N_3534,N_2523,N_2916);
nor U3535 (N_3535,N_2930,N_2991);
nor U3536 (N_3536,N_2814,N_2930);
xor U3537 (N_3537,N_2593,N_2794);
xor U3538 (N_3538,N_2927,N_2735);
and U3539 (N_3539,N_2675,N_2514);
nand U3540 (N_3540,N_2859,N_2616);
or U3541 (N_3541,N_2562,N_2837);
and U3542 (N_3542,N_2677,N_2593);
nand U3543 (N_3543,N_2762,N_2848);
nor U3544 (N_3544,N_2782,N_2640);
or U3545 (N_3545,N_2451,N_2579);
nand U3546 (N_3546,N_2554,N_2942);
xor U3547 (N_3547,N_2430,N_2846);
or U3548 (N_3548,N_2848,N_2826);
or U3549 (N_3549,N_2428,N_2618);
nand U3550 (N_3550,N_2532,N_2557);
or U3551 (N_3551,N_2763,N_2757);
nand U3552 (N_3552,N_2573,N_2477);
or U3553 (N_3553,N_2608,N_2986);
nand U3554 (N_3554,N_2412,N_2696);
or U3555 (N_3555,N_2984,N_2469);
nand U3556 (N_3556,N_2793,N_2976);
or U3557 (N_3557,N_2955,N_2526);
nor U3558 (N_3558,N_2954,N_2882);
nor U3559 (N_3559,N_2854,N_2791);
nor U3560 (N_3560,N_2461,N_2449);
nor U3561 (N_3561,N_2968,N_2775);
and U3562 (N_3562,N_2424,N_2953);
and U3563 (N_3563,N_2715,N_2845);
nor U3564 (N_3564,N_2503,N_2786);
and U3565 (N_3565,N_2803,N_2898);
nor U3566 (N_3566,N_2492,N_2703);
nand U3567 (N_3567,N_2723,N_2896);
nand U3568 (N_3568,N_2785,N_2741);
and U3569 (N_3569,N_2627,N_2791);
xnor U3570 (N_3570,N_2457,N_2425);
or U3571 (N_3571,N_2703,N_2555);
nor U3572 (N_3572,N_2591,N_2713);
or U3573 (N_3573,N_2532,N_2591);
or U3574 (N_3574,N_2947,N_2786);
and U3575 (N_3575,N_2799,N_2666);
and U3576 (N_3576,N_2568,N_2745);
and U3577 (N_3577,N_2494,N_2932);
nor U3578 (N_3578,N_2481,N_2980);
or U3579 (N_3579,N_2819,N_2590);
or U3580 (N_3580,N_2828,N_2927);
and U3581 (N_3581,N_2755,N_2569);
nor U3582 (N_3582,N_2643,N_2495);
xor U3583 (N_3583,N_2835,N_2572);
nor U3584 (N_3584,N_2458,N_2705);
nor U3585 (N_3585,N_2905,N_2451);
and U3586 (N_3586,N_2736,N_2792);
or U3587 (N_3587,N_2976,N_2694);
nand U3588 (N_3588,N_2581,N_2539);
nand U3589 (N_3589,N_2423,N_2794);
nor U3590 (N_3590,N_2558,N_2744);
or U3591 (N_3591,N_2766,N_2828);
or U3592 (N_3592,N_2583,N_2754);
or U3593 (N_3593,N_2854,N_2825);
xnor U3594 (N_3594,N_2427,N_2636);
and U3595 (N_3595,N_2488,N_2781);
or U3596 (N_3596,N_2693,N_2536);
nor U3597 (N_3597,N_2726,N_2985);
nand U3598 (N_3598,N_2564,N_2963);
nand U3599 (N_3599,N_2691,N_2745);
and U3600 (N_3600,N_3432,N_3398);
xnor U3601 (N_3601,N_3422,N_3329);
and U3602 (N_3602,N_3449,N_3479);
nor U3603 (N_3603,N_3150,N_3180);
nand U3604 (N_3604,N_3099,N_3297);
or U3605 (N_3605,N_3222,N_3084);
or U3606 (N_3606,N_3541,N_3106);
and U3607 (N_3607,N_3536,N_3247);
and U3608 (N_3608,N_3585,N_3320);
xor U3609 (N_3609,N_3548,N_3416);
nand U3610 (N_3610,N_3053,N_3396);
and U3611 (N_3611,N_3064,N_3273);
nand U3612 (N_3612,N_3505,N_3547);
xnor U3613 (N_3613,N_3108,N_3095);
nand U3614 (N_3614,N_3510,N_3278);
nor U3615 (N_3615,N_3216,N_3277);
nor U3616 (N_3616,N_3201,N_3267);
or U3617 (N_3617,N_3447,N_3306);
nand U3618 (N_3618,N_3014,N_3395);
and U3619 (N_3619,N_3575,N_3072);
nor U3620 (N_3620,N_3132,N_3570);
nand U3621 (N_3621,N_3070,N_3076);
or U3622 (N_3622,N_3562,N_3442);
nand U3623 (N_3623,N_3255,N_3250);
nand U3624 (N_3624,N_3314,N_3593);
and U3625 (N_3625,N_3451,N_3266);
or U3626 (N_3626,N_3098,N_3013);
nand U3627 (N_3627,N_3419,N_3433);
and U3628 (N_3628,N_3135,N_3022);
or U3629 (N_3629,N_3597,N_3217);
nand U3630 (N_3630,N_3345,N_3166);
or U3631 (N_3631,N_3424,N_3181);
nand U3632 (N_3632,N_3225,N_3293);
nand U3633 (N_3633,N_3435,N_3240);
and U3634 (N_3634,N_3552,N_3058);
nand U3635 (N_3635,N_3199,N_3592);
xor U3636 (N_3636,N_3349,N_3382);
or U3637 (N_3637,N_3056,N_3459);
and U3638 (N_3638,N_3391,N_3004);
nor U3639 (N_3639,N_3521,N_3326);
nor U3640 (N_3640,N_3378,N_3475);
nand U3641 (N_3641,N_3373,N_3558);
and U3642 (N_3642,N_3403,N_3178);
nor U3643 (N_3643,N_3185,N_3028);
and U3644 (N_3644,N_3439,N_3026);
xnor U3645 (N_3645,N_3532,N_3235);
and U3646 (N_3646,N_3500,N_3468);
nor U3647 (N_3647,N_3526,N_3389);
and U3648 (N_3648,N_3352,N_3173);
or U3649 (N_3649,N_3044,N_3342);
xor U3650 (N_3650,N_3138,N_3128);
or U3651 (N_3651,N_3234,N_3042);
nand U3652 (N_3652,N_3177,N_3126);
or U3653 (N_3653,N_3012,N_3259);
or U3654 (N_3654,N_3100,N_3289);
and U3655 (N_3655,N_3092,N_3283);
nand U3656 (N_3656,N_3244,N_3364);
or U3657 (N_3657,N_3290,N_3426);
and U3658 (N_3658,N_3107,N_3474);
nor U3659 (N_3659,N_3501,N_3233);
or U3660 (N_3660,N_3366,N_3334);
xor U3661 (N_3661,N_3415,N_3462);
and U3662 (N_3662,N_3469,N_3365);
nand U3663 (N_3663,N_3370,N_3425);
or U3664 (N_3664,N_3109,N_3412);
nand U3665 (N_3665,N_3402,N_3008);
nor U3666 (N_3666,N_3243,N_3060);
or U3667 (N_3667,N_3583,N_3379);
or U3668 (N_3668,N_3354,N_3112);
nor U3669 (N_3669,N_3404,N_3495);
and U3670 (N_3670,N_3227,N_3139);
and U3671 (N_3671,N_3172,N_3577);
xor U3672 (N_3672,N_3579,N_3035);
xor U3673 (N_3673,N_3492,N_3193);
or U3674 (N_3674,N_3551,N_3351);
nor U3675 (N_3675,N_3472,N_3061);
nand U3676 (N_3676,N_3586,N_3337);
nand U3677 (N_3677,N_3446,N_3321);
nand U3678 (N_3678,N_3184,N_3335);
nand U3679 (N_3679,N_3487,N_3027);
nand U3680 (N_3680,N_3163,N_3186);
or U3681 (N_3681,N_3068,N_3448);
nor U3682 (N_3682,N_3528,N_3271);
and U3683 (N_3683,N_3175,N_3343);
or U3684 (N_3684,N_3274,N_3197);
or U3685 (N_3685,N_3176,N_3527);
or U3686 (N_3686,N_3145,N_3587);
xnor U3687 (N_3687,N_3518,N_3405);
nand U3688 (N_3688,N_3434,N_3312);
or U3689 (N_3689,N_3350,N_3101);
xor U3690 (N_3690,N_3540,N_3553);
and U3691 (N_3691,N_3077,N_3050);
xnor U3692 (N_3692,N_3513,N_3021);
nand U3693 (N_3693,N_3386,N_3567);
nand U3694 (N_3694,N_3245,N_3102);
nor U3695 (N_3695,N_3535,N_3237);
and U3696 (N_3696,N_3104,N_3323);
nand U3697 (N_3697,N_3231,N_3230);
or U3698 (N_3698,N_3212,N_3117);
xor U3699 (N_3699,N_3168,N_3534);
nand U3700 (N_3700,N_3074,N_3158);
or U3701 (N_3701,N_3340,N_3143);
or U3702 (N_3702,N_3355,N_3020);
nor U3703 (N_3703,N_3006,N_3307);
and U3704 (N_3704,N_3576,N_3203);
or U3705 (N_3705,N_3480,N_3516);
and U3706 (N_3706,N_3580,N_3322);
and U3707 (N_3707,N_3530,N_3588);
nand U3708 (N_3708,N_3563,N_3221);
nor U3709 (N_3709,N_3003,N_3254);
and U3710 (N_3710,N_3589,N_3443);
nor U3711 (N_3711,N_3301,N_3377);
or U3712 (N_3712,N_3111,N_3493);
and U3713 (N_3713,N_3578,N_3187);
nor U3714 (N_3714,N_3327,N_3037);
nand U3715 (N_3715,N_3408,N_3401);
nor U3716 (N_3716,N_3292,N_3573);
nor U3717 (N_3717,N_3457,N_3539);
and U3718 (N_3718,N_3001,N_3188);
xnor U3719 (N_3719,N_3167,N_3287);
nor U3720 (N_3720,N_3206,N_3131);
nand U3721 (N_3721,N_3091,N_3236);
nor U3722 (N_3722,N_3110,N_3149);
nor U3723 (N_3723,N_3363,N_3204);
or U3724 (N_3724,N_3229,N_3399);
nor U3725 (N_3725,N_3394,N_3146);
and U3726 (N_3726,N_3114,N_3078);
xor U3727 (N_3727,N_3465,N_3062);
and U3728 (N_3728,N_3280,N_3407);
xnor U3729 (N_3729,N_3317,N_3452);
or U3730 (N_3730,N_3560,N_3262);
nor U3731 (N_3731,N_3392,N_3445);
nor U3732 (N_3732,N_3113,N_3136);
nor U3733 (N_3733,N_3137,N_3458);
nor U3734 (N_3734,N_3569,N_3380);
xor U3735 (N_3735,N_3319,N_3333);
or U3736 (N_3736,N_3599,N_3023);
or U3737 (N_3737,N_3444,N_3441);
or U3738 (N_3738,N_3356,N_3315);
nor U3739 (N_3739,N_3344,N_3454);
nor U3740 (N_3740,N_3367,N_3249);
or U3741 (N_3741,N_3466,N_3071);
nand U3742 (N_3742,N_3257,N_3502);
nor U3743 (N_3743,N_3121,N_3226);
or U3744 (N_3744,N_3397,N_3120);
and U3745 (N_3745,N_3471,N_3192);
nand U3746 (N_3746,N_3284,N_3122);
nor U3747 (N_3747,N_3515,N_3304);
or U3748 (N_3748,N_3461,N_3276);
nand U3749 (N_3749,N_3279,N_3088);
nor U3750 (N_3750,N_3118,N_3507);
or U3751 (N_3751,N_3134,N_3130);
nand U3752 (N_3752,N_3195,N_3160);
and U3753 (N_3753,N_3239,N_3253);
nand U3754 (N_3754,N_3223,N_3411);
nand U3755 (N_3755,N_3248,N_3269);
nor U3756 (N_3756,N_3010,N_3594);
or U3757 (N_3757,N_3478,N_3385);
nor U3758 (N_3758,N_3499,N_3059);
nand U3759 (N_3759,N_3034,N_3209);
nand U3760 (N_3760,N_3572,N_3511);
xnor U3761 (N_3761,N_3202,N_3311);
nand U3762 (N_3762,N_3543,N_3094);
nand U3763 (N_3763,N_3361,N_3305);
xnor U3764 (N_3764,N_3538,N_3413);
or U3765 (N_3765,N_3085,N_3232);
and U3766 (N_3766,N_3119,N_3252);
nor U3767 (N_3767,N_3557,N_3215);
nor U3768 (N_3768,N_3219,N_3238);
nand U3769 (N_3769,N_3453,N_3414);
and U3770 (N_3770,N_3241,N_3200);
nand U3771 (N_3771,N_3598,N_3295);
nor U3772 (N_3772,N_3481,N_3360);
nand U3773 (N_3773,N_3251,N_3224);
nand U3774 (N_3774,N_3048,N_3152);
nor U3775 (N_3775,N_3147,N_3484);
xor U3776 (N_3776,N_3332,N_3455);
nor U3777 (N_3777,N_3420,N_3325);
or U3778 (N_3778,N_3550,N_3596);
and U3779 (N_3779,N_3549,N_3330);
and U3780 (N_3780,N_3191,N_3038);
nor U3781 (N_3781,N_3018,N_3522);
and U3782 (N_3782,N_3073,N_3299);
and U3783 (N_3783,N_3517,N_3375);
nor U3784 (N_3784,N_3318,N_3463);
nand U3785 (N_3785,N_3157,N_3069);
nor U3786 (N_3786,N_3316,N_3116);
or U3787 (N_3787,N_3584,N_3151);
nand U3788 (N_3788,N_3440,N_3270);
or U3789 (N_3789,N_3007,N_3063);
nor U3790 (N_3790,N_3506,N_3488);
or U3791 (N_3791,N_3546,N_3542);
or U3792 (N_3792,N_3336,N_3179);
nor U3793 (N_3793,N_3388,N_3418);
nand U3794 (N_3794,N_3554,N_3368);
nor U3795 (N_3795,N_3519,N_3220);
and U3796 (N_3796,N_3002,N_3450);
nor U3797 (N_3797,N_3310,N_3156);
nor U3798 (N_3798,N_3384,N_3141);
and U3799 (N_3799,N_3300,N_3043);
or U3800 (N_3800,N_3347,N_3093);
or U3801 (N_3801,N_3508,N_3000);
and U3802 (N_3802,N_3524,N_3303);
or U3803 (N_3803,N_3559,N_3127);
or U3804 (N_3804,N_3490,N_3066);
nor U3805 (N_3805,N_3486,N_3437);
nor U3806 (N_3806,N_3090,N_3189);
or U3807 (N_3807,N_3590,N_3207);
nand U3808 (N_3808,N_3359,N_3574);
and U3809 (N_3809,N_3228,N_3369);
and U3810 (N_3810,N_3075,N_3242);
or U3811 (N_3811,N_3125,N_3258);
and U3812 (N_3812,N_3049,N_3467);
nor U3813 (N_3813,N_3282,N_3346);
and U3814 (N_3814,N_3039,N_3009);
xnor U3815 (N_3815,N_3464,N_3214);
or U3816 (N_3816,N_3086,N_3423);
or U3817 (N_3817,N_3040,N_3256);
nor U3818 (N_3818,N_3210,N_3371);
nand U3819 (N_3819,N_3264,N_3555);
xor U3820 (N_3820,N_3154,N_3159);
and U3821 (N_3821,N_3313,N_3483);
nor U3822 (N_3822,N_3011,N_3218);
and U3823 (N_3823,N_3065,N_3161);
nor U3824 (N_3824,N_3196,N_3328);
nand U3825 (N_3825,N_3436,N_3124);
or U3826 (N_3826,N_3041,N_3162);
nor U3827 (N_3827,N_3083,N_3308);
or U3828 (N_3828,N_3353,N_3531);
nand U3829 (N_3829,N_3190,N_3281);
nand U3830 (N_3830,N_3498,N_3571);
nand U3831 (N_3831,N_3097,N_3174);
nor U3832 (N_3832,N_3406,N_3144);
or U3833 (N_3833,N_3031,N_3261);
and U3834 (N_3834,N_3429,N_3182);
nor U3835 (N_3835,N_3080,N_3400);
and U3836 (N_3836,N_3544,N_3339);
nand U3837 (N_3837,N_3171,N_3194);
nand U3838 (N_3838,N_3067,N_3082);
nor U3839 (N_3839,N_3081,N_3268);
xnor U3840 (N_3840,N_3087,N_3105);
and U3841 (N_3841,N_3079,N_3142);
or U3842 (N_3842,N_3129,N_3165);
and U3843 (N_3843,N_3566,N_3438);
or U3844 (N_3844,N_3372,N_3005);
nor U3845 (N_3845,N_3123,N_3054);
and U3846 (N_3846,N_3512,N_3030);
nand U3847 (N_3847,N_3046,N_3476);
and U3848 (N_3848,N_3383,N_3497);
xor U3849 (N_3849,N_3430,N_3265);
nor U3850 (N_3850,N_3381,N_3051);
or U3851 (N_3851,N_3591,N_3148);
or U3852 (N_3852,N_3491,N_3409);
nand U3853 (N_3853,N_3545,N_3291);
nand U3854 (N_3854,N_3489,N_3155);
xnor U3855 (N_3855,N_3564,N_3561);
nor U3856 (N_3856,N_3032,N_3052);
or U3857 (N_3857,N_3015,N_3460);
xor U3858 (N_3858,N_3324,N_3431);
nor U3859 (N_3859,N_3523,N_3529);
or U3860 (N_3860,N_3568,N_3025);
nor U3861 (N_3861,N_3169,N_3211);
nand U3862 (N_3862,N_3427,N_3348);
xnor U3863 (N_3863,N_3358,N_3205);
or U3864 (N_3864,N_3362,N_3470);
and U3865 (N_3865,N_3341,N_3024);
or U3866 (N_3866,N_3374,N_3260);
nand U3867 (N_3867,N_3309,N_3033);
or U3868 (N_3868,N_3298,N_3417);
xnor U3869 (N_3869,N_3514,N_3164);
nand U3870 (N_3870,N_3055,N_3272);
or U3871 (N_3871,N_3477,N_3482);
xnor U3872 (N_3872,N_3504,N_3565);
xor U3873 (N_3873,N_3581,N_3331);
and U3874 (N_3874,N_3246,N_3387);
or U3875 (N_3875,N_3096,N_3338);
or U3876 (N_3876,N_3285,N_3410);
nor U3877 (N_3877,N_3525,N_3036);
nand U3878 (N_3878,N_3421,N_3556);
nand U3879 (N_3879,N_3485,N_3473);
nor U3880 (N_3880,N_3133,N_3153);
and U3881 (N_3881,N_3520,N_3428);
and U3882 (N_3882,N_3017,N_3019);
nand U3883 (N_3883,N_3103,N_3496);
and U3884 (N_3884,N_3595,N_3275);
nand U3885 (N_3885,N_3213,N_3503);
nand U3886 (N_3886,N_3376,N_3582);
xnor U3887 (N_3887,N_3288,N_3089);
nand U3888 (N_3888,N_3296,N_3393);
or U3889 (N_3889,N_3045,N_3057);
or U3890 (N_3890,N_3183,N_3357);
nand U3891 (N_3891,N_3533,N_3537);
nand U3892 (N_3892,N_3509,N_3170);
or U3893 (N_3893,N_3302,N_3198);
nor U3894 (N_3894,N_3016,N_3286);
or U3895 (N_3895,N_3115,N_3456);
nand U3896 (N_3896,N_3263,N_3494);
nand U3897 (N_3897,N_3140,N_3390);
xor U3898 (N_3898,N_3208,N_3029);
nor U3899 (N_3899,N_3294,N_3047);
nor U3900 (N_3900,N_3177,N_3097);
or U3901 (N_3901,N_3272,N_3465);
nand U3902 (N_3902,N_3356,N_3303);
and U3903 (N_3903,N_3170,N_3499);
xor U3904 (N_3904,N_3187,N_3548);
nor U3905 (N_3905,N_3320,N_3360);
or U3906 (N_3906,N_3256,N_3283);
nand U3907 (N_3907,N_3088,N_3048);
nor U3908 (N_3908,N_3141,N_3329);
or U3909 (N_3909,N_3507,N_3245);
and U3910 (N_3910,N_3571,N_3175);
or U3911 (N_3911,N_3098,N_3417);
nand U3912 (N_3912,N_3147,N_3585);
nor U3913 (N_3913,N_3112,N_3269);
nor U3914 (N_3914,N_3563,N_3361);
and U3915 (N_3915,N_3160,N_3441);
nand U3916 (N_3916,N_3242,N_3574);
nor U3917 (N_3917,N_3325,N_3446);
and U3918 (N_3918,N_3545,N_3175);
nand U3919 (N_3919,N_3204,N_3457);
nor U3920 (N_3920,N_3349,N_3111);
xor U3921 (N_3921,N_3232,N_3047);
nand U3922 (N_3922,N_3573,N_3382);
or U3923 (N_3923,N_3483,N_3185);
nand U3924 (N_3924,N_3470,N_3528);
nor U3925 (N_3925,N_3383,N_3400);
or U3926 (N_3926,N_3365,N_3529);
nor U3927 (N_3927,N_3385,N_3264);
and U3928 (N_3928,N_3185,N_3016);
xnor U3929 (N_3929,N_3377,N_3467);
nand U3930 (N_3930,N_3459,N_3166);
nor U3931 (N_3931,N_3406,N_3264);
and U3932 (N_3932,N_3304,N_3260);
or U3933 (N_3933,N_3211,N_3582);
or U3934 (N_3934,N_3244,N_3306);
nor U3935 (N_3935,N_3293,N_3442);
nand U3936 (N_3936,N_3536,N_3516);
and U3937 (N_3937,N_3598,N_3590);
nor U3938 (N_3938,N_3188,N_3051);
and U3939 (N_3939,N_3108,N_3184);
nand U3940 (N_3940,N_3393,N_3141);
or U3941 (N_3941,N_3170,N_3442);
nand U3942 (N_3942,N_3443,N_3154);
or U3943 (N_3943,N_3373,N_3308);
nor U3944 (N_3944,N_3187,N_3435);
or U3945 (N_3945,N_3124,N_3395);
nand U3946 (N_3946,N_3278,N_3030);
and U3947 (N_3947,N_3124,N_3052);
and U3948 (N_3948,N_3568,N_3530);
or U3949 (N_3949,N_3028,N_3352);
nor U3950 (N_3950,N_3215,N_3510);
nand U3951 (N_3951,N_3319,N_3338);
or U3952 (N_3952,N_3567,N_3355);
nor U3953 (N_3953,N_3240,N_3433);
nand U3954 (N_3954,N_3478,N_3448);
nand U3955 (N_3955,N_3301,N_3597);
nand U3956 (N_3956,N_3524,N_3089);
and U3957 (N_3957,N_3173,N_3346);
nor U3958 (N_3958,N_3287,N_3464);
and U3959 (N_3959,N_3095,N_3488);
xor U3960 (N_3960,N_3281,N_3027);
or U3961 (N_3961,N_3003,N_3479);
nor U3962 (N_3962,N_3011,N_3521);
nand U3963 (N_3963,N_3464,N_3238);
or U3964 (N_3964,N_3148,N_3496);
or U3965 (N_3965,N_3171,N_3278);
and U3966 (N_3966,N_3289,N_3547);
nor U3967 (N_3967,N_3226,N_3094);
nor U3968 (N_3968,N_3487,N_3317);
nor U3969 (N_3969,N_3451,N_3398);
or U3970 (N_3970,N_3051,N_3168);
and U3971 (N_3971,N_3239,N_3252);
nand U3972 (N_3972,N_3294,N_3023);
nand U3973 (N_3973,N_3401,N_3100);
or U3974 (N_3974,N_3113,N_3328);
nor U3975 (N_3975,N_3296,N_3033);
nand U3976 (N_3976,N_3511,N_3349);
xor U3977 (N_3977,N_3457,N_3570);
xnor U3978 (N_3978,N_3251,N_3491);
and U3979 (N_3979,N_3214,N_3439);
xnor U3980 (N_3980,N_3010,N_3225);
and U3981 (N_3981,N_3326,N_3049);
and U3982 (N_3982,N_3184,N_3446);
nor U3983 (N_3983,N_3104,N_3394);
nand U3984 (N_3984,N_3464,N_3415);
nor U3985 (N_3985,N_3422,N_3254);
xor U3986 (N_3986,N_3495,N_3048);
or U3987 (N_3987,N_3175,N_3529);
nand U3988 (N_3988,N_3357,N_3002);
xnor U3989 (N_3989,N_3329,N_3401);
xor U3990 (N_3990,N_3542,N_3246);
nand U3991 (N_3991,N_3354,N_3322);
xor U3992 (N_3992,N_3344,N_3055);
and U3993 (N_3993,N_3348,N_3037);
and U3994 (N_3994,N_3351,N_3503);
nand U3995 (N_3995,N_3322,N_3269);
nor U3996 (N_3996,N_3223,N_3122);
nor U3997 (N_3997,N_3558,N_3196);
nand U3998 (N_3998,N_3561,N_3299);
or U3999 (N_3999,N_3395,N_3429);
xnor U4000 (N_4000,N_3560,N_3320);
nand U4001 (N_4001,N_3305,N_3360);
nand U4002 (N_4002,N_3431,N_3320);
nand U4003 (N_4003,N_3026,N_3574);
and U4004 (N_4004,N_3145,N_3340);
nand U4005 (N_4005,N_3117,N_3434);
nor U4006 (N_4006,N_3333,N_3074);
and U4007 (N_4007,N_3233,N_3156);
nor U4008 (N_4008,N_3504,N_3416);
nor U4009 (N_4009,N_3425,N_3595);
nor U4010 (N_4010,N_3093,N_3203);
or U4011 (N_4011,N_3006,N_3162);
nor U4012 (N_4012,N_3417,N_3515);
nor U4013 (N_4013,N_3275,N_3103);
nor U4014 (N_4014,N_3163,N_3521);
and U4015 (N_4015,N_3186,N_3513);
nand U4016 (N_4016,N_3356,N_3279);
or U4017 (N_4017,N_3246,N_3037);
or U4018 (N_4018,N_3335,N_3431);
or U4019 (N_4019,N_3542,N_3076);
nor U4020 (N_4020,N_3554,N_3528);
nand U4021 (N_4021,N_3193,N_3006);
and U4022 (N_4022,N_3564,N_3018);
nor U4023 (N_4023,N_3520,N_3559);
nor U4024 (N_4024,N_3498,N_3149);
nand U4025 (N_4025,N_3115,N_3411);
nand U4026 (N_4026,N_3029,N_3376);
or U4027 (N_4027,N_3472,N_3223);
nor U4028 (N_4028,N_3321,N_3478);
or U4029 (N_4029,N_3565,N_3220);
or U4030 (N_4030,N_3292,N_3127);
nand U4031 (N_4031,N_3172,N_3497);
nand U4032 (N_4032,N_3341,N_3124);
nor U4033 (N_4033,N_3074,N_3453);
nand U4034 (N_4034,N_3277,N_3330);
and U4035 (N_4035,N_3008,N_3267);
or U4036 (N_4036,N_3591,N_3551);
and U4037 (N_4037,N_3456,N_3335);
and U4038 (N_4038,N_3088,N_3330);
and U4039 (N_4039,N_3339,N_3499);
nor U4040 (N_4040,N_3535,N_3135);
and U4041 (N_4041,N_3289,N_3234);
and U4042 (N_4042,N_3465,N_3173);
nand U4043 (N_4043,N_3086,N_3085);
nor U4044 (N_4044,N_3531,N_3133);
and U4045 (N_4045,N_3322,N_3204);
or U4046 (N_4046,N_3392,N_3242);
or U4047 (N_4047,N_3285,N_3392);
or U4048 (N_4048,N_3130,N_3360);
nor U4049 (N_4049,N_3039,N_3263);
xnor U4050 (N_4050,N_3289,N_3494);
or U4051 (N_4051,N_3336,N_3430);
nor U4052 (N_4052,N_3077,N_3294);
and U4053 (N_4053,N_3431,N_3338);
and U4054 (N_4054,N_3183,N_3142);
nor U4055 (N_4055,N_3224,N_3019);
or U4056 (N_4056,N_3506,N_3339);
and U4057 (N_4057,N_3506,N_3186);
nand U4058 (N_4058,N_3189,N_3019);
and U4059 (N_4059,N_3251,N_3225);
and U4060 (N_4060,N_3075,N_3079);
and U4061 (N_4061,N_3488,N_3192);
xnor U4062 (N_4062,N_3215,N_3493);
nor U4063 (N_4063,N_3309,N_3522);
nand U4064 (N_4064,N_3038,N_3480);
or U4065 (N_4065,N_3510,N_3474);
or U4066 (N_4066,N_3266,N_3544);
and U4067 (N_4067,N_3599,N_3467);
nor U4068 (N_4068,N_3450,N_3301);
and U4069 (N_4069,N_3257,N_3022);
nand U4070 (N_4070,N_3377,N_3389);
xor U4071 (N_4071,N_3469,N_3311);
xor U4072 (N_4072,N_3080,N_3507);
nor U4073 (N_4073,N_3112,N_3411);
nand U4074 (N_4074,N_3470,N_3596);
and U4075 (N_4075,N_3053,N_3063);
or U4076 (N_4076,N_3398,N_3117);
nor U4077 (N_4077,N_3521,N_3107);
xor U4078 (N_4078,N_3538,N_3325);
and U4079 (N_4079,N_3061,N_3093);
or U4080 (N_4080,N_3438,N_3305);
nor U4081 (N_4081,N_3087,N_3316);
or U4082 (N_4082,N_3293,N_3132);
or U4083 (N_4083,N_3189,N_3451);
or U4084 (N_4084,N_3463,N_3338);
nand U4085 (N_4085,N_3277,N_3117);
and U4086 (N_4086,N_3290,N_3269);
nor U4087 (N_4087,N_3378,N_3114);
xor U4088 (N_4088,N_3477,N_3024);
xor U4089 (N_4089,N_3002,N_3421);
nor U4090 (N_4090,N_3391,N_3403);
nand U4091 (N_4091,N_3309,N_3404);
and U4092 (N_4092,N_3201,N_3331);
nand U4093 (N_4093,N_3063,N_3055);
xnor U4094 (N_4094,N_3116,N_3040);
or U4095 (N_4095,N_3080,N_3406);
nand U4096 (N_4096,N_3514,N_3471);
nor U4097 (N_4097,N_3348,N_3178);
nand U4098 (N_4098,N_3324,N_3358);
xor U4099 (N_4099,N_3108,N_3203);
or U4100 (N_4100,N_3349,N_3191);
nand U4101 (N_4101,N_3264,N_3309);
nand U4102 (N_4102,N_3578,N_3269);
nor U4103 (N_4103,N_3098,N_3220);
or U4104 (N_4104,N_3537,N_3191);
nor U4105 (N_4105,N_3512,N_3383);
nor U4106 (N_4106,N_3264,N_3245);
nor U4107 (N_4107,N_3359,N_3596);
or U4108 (N_4108,N_3155,N_3202);
or U4109 (N_4109,N_3557,N_3009);
or U4110 (N_4110,N_3512,N_3425);
nand U4111 (N_4111,N_3148,N_3215);
nor U4112 (N_4112,N_3490,N_3002);
and U4113 (N_4113,N_3528,N_3101);
nand U4114 (N_4114,N_3217,N_3296);
or U4115 (N_4115,N_3398,N_3464);
xor U4116 (N_4116,N_3197,N_3318);
and U4117 (N_4117,N_3494,N_3276);
and U4118 (N_4118,N_3075,N_3191);
or U4119 (N_4119,N_3326,N_3362);
xnor U4120 (N_4120,N_3025,N_3491);
xnor U4121 (N_4121,N_3335,N_3024);
and U4122 (N_4122,N_3059,N_3212);
xnor U4123 (N_4123,N_3593,N_3202);
nand U4124 (N_4124,N_3360,N_3077);
nand U4125 (N_4125,N_3407,N_3294);
and U4126 (N_4126,N_3211,N_3502);
xnor U4127 (N_4127,N_3500,N_3374);
or U4128 (N_4128,N_3386,N_3198);
and U4129 (N_4129,N_3422,N_3006);
xor U4130 (N_4130,N_3452,N_3320);
or U4131 (N_4131,N_3141,N_3519);
and U4132 (N_4132,N_3466,N_3488);
or U4133 (N_4133,N_3284,N_3268);
and U4134 (N_4134,N_3022,N_3304);
nor U4135 (N_4135,N_3000,N_3019);
nand U4136 (N_4136,N_3467,N_3297);
nor U4137 (N_4137,N_3057,N_3023);
nor U4138 (N_4138,N_3336,N_3531);
nand U4139 (N_4139,N_3247,N_3069);
xor U4140 (N_4140,N_3022,N_3435);
nand U4141 (N_4141,N_3464,N_3504);
nor U4142 (N_4142,N_3450,N_3298);
nor U4143 (N_4143,N_3029,N_3242);
and U4144 (N_4144,N_3254,N_3054);
nor U4145 (N_4145,N_3215,N_3155);
and U4146 (N_4146,N_3292,N_3368);
nand U4147 (N_4147,N_3379,N_3185);
and U4148 (N_4148,N_3491,N_3163);
or U4149 (N_4149,N_3250,N_3093);
nor U4150 (N_4150,N_3284,N_3351);
xor U4151 (N_4151,N_3118,N_3239);
or U4152 (N_4152,N_3509,N_3199);
and U4153 (N_4153,N_3036,N_3031);
and U4154 (N_4154,N_3537,N_3313);
and U4155 (N_4155,N_3026,N_3367);
nand U4156 (N_4156,N_3497,N_3229);
and U4157 (N_4157,N_3334,N_3383);
nor U4158 (N_4158,N_3533,N_3095);
or U4159 (N_4159,N_3448,N_3098);
and U4160 (N_4160,N_3173,N_3079);
nand U4161 (N_4161,N_3434,N_3116);
nor U4162 (N_4162,N_3183,N_3017);
nor U4163 (N_4163,N_3075,N_3413);
and U4164 (N_4164,N_3255,N_3052);
and U4165 (N_4165,N_3254,N_3593);
or U4166 (N_4166,N_3079,N_3475);
nor U4167 (N_4167,N_3579,N_3529);
xnor U4168 (N_4168,N_3595,N_3180);
nand U4169 (N_4169,N_3494,N_3193);
nand U4170 (N_4170,N_3539,N_3304);
xor U4171 (N_4171,N_3451,N_3072);
and U4172 (N_4172,N_3227,N_3216);
nand U4173 (N_4173,N_3501,N_3278);
or U4174 (N_4174,N_3328,N_3457);
or U4175 (N_4175,N_3509,N_3046);
or U4176 (N_4176,N_3296,N_3488);
and U4177 (N_4177,N_3589,N_3164);
and U4178 (N_4178,N_3141,N_3127);
xnor U4179 (N_4179,N_3216,N_3519);
and U4180 (N_4180,N_3344,N_3483);
xor U4181 (N_4181,N_3317,N_3283);
or U4182 (N_4182,N_3153,N_3129);
nand U4183 (N_4183,N_3071,N_3274);
and U4184 (N_4184,N_3444,N_3549);
or U4185 (N_4185,N_3449,N_3512);
and U4186 (N_4186,N_3107,N_3105);
or U4187 (N_4187,N_3402,N_3383);
nand U4188 (N_4188,N_3475,N_3473);
nor U4189 (N_4189,N_3414,N_3341);
and U4190 (N_4190,N_3565,N_3060);
nor U4191 (N_4191,N_3219,N_3382);
or U4192 (N_4192,N_3485,N_3137);
and U4193 (N_4193,N_3572,N_3120);
or U4194 (N_4194,N_3509,N_3361);
nor U4195 (N_4195,N_3559,N_3458);
xor U4196 (N_4196,N_3471,N_3161);
nor U4197 (N_4197,N_3525,N_3447);
nor U4198 (N_4198,N_3237,N_3363);
nor U4199 (N_4199,N_3544,N_3418);
or U4200 (N_4200,N_4166,N_3850);
nor U4201 (N_4201,N_3950,N_3659);
nor U4202 (N_4202,N_3867,N_3662);
xor U4203 (N_4203,N_4175,N_4184);
and U4204 (N_4204,N_4048,N_3692);
xor U4205 (N_4205,N_3828,N_3743);
and U4206 (N_4206,N_3674,N_4099);
or U4207 (N_4207,N_4155,N_3627);
and U4208 (N_4208,N_3824,N_3992);
nor U4209 (N_4209,N_4195,N_3952);
and U4210 (N_4210,N_4016,N_4032);
and U4211 (N_4211,N_3904,N_4100);
or U4212 (N_4212,N_3975,N_4127);
nand U4213 (N_4213,N_3782,N_4086);
and U4214 (N_4214,N_3637,N_3754);
or U4215 (N_4215,N_4033,N_4156);
nor U4216 (N_4216,N_3874,N_3780);
nand U4217 (N_4217,N_4000,N_3636);
nor U4218 (N_4218,N_4054,N_3806);
xnor U4219 (N_4219,N_4119,N_4006);
nand U4220 (N_4220,N_3956,N_3673);
or U4221 (N_4221,N_3919,N_3752);
nand U4222 (N_4222,N_3954,N_3978);
nand U4223 (N_4223,N_4046,N_3642);
and U4224 (N_4224,N_3779,N_3876);
and U4225 (N_4225,N_4051,N_3615);
and U4226 (N_4226,N_3766,N_3696);
nor U4227 (N_4227,N_3823,N_4049);
nand U4228 (N_4228,N_4029,N_3624);
or U4229 (N_4229,N_3971,N_4167);
or U4230 (N_4230,N_3611,N_3861);
or U4231 (N_4231,N_3713,N_4142);
nand U4232 (N_4232,N_3848,N_4196);
nand U4233 (N_4233,N_3750,N_3807);
nand U4234 (N_4234,N_3990,N_4063);
nor U4235 (N_4235,N_3645,N_3676);
or U4236 (N_4236,N_3833,N_4084);
xor U4237 (N_4237,N_3706,N_3755);
or U4238 (N_4238,N_3973,N_4023);
nand U4239 (N_4239,N_3654,N_3870);
nand U4240 (N_4240,N_3858,N_3701);
or U4241 (N_4241,N_3658,N_3810);
xor U4242 (N_4242,N_4133,N_4126);
xor U4243 (N_4243,N_3809,N_3891);
and U4244 (N_4244,N_3830,N_4069);
or U4245 (N_4245,N_4015,N_3834);
and U4246 (N_4246,N_3923,N_4134);
and U4247 (N_4247,N_4059,N_3839);
nand U4248 (N_4248,N_4178,N_3953);
xor U4249 (N_4249,N_4075,N_4136);
or U4250 (N_4250,N_4001,N_3970);
nand U4251 (N_4251,N_4194,N_4064);
or U4252 (N_4252,N_3880,N_3957);
and U4253 (N_4253,N_3749,N_3966);
and U4254 (N_4254,N_3770,N_3688);
nand U4255 (N_4255,N_3836,N_3693);
or U4256 (N_4256,N_4012,N_3663);
nor U4257 (N_4257,N_3753,N_4082);
or U4258 (N_4258,N_3831,N_4101);
and U4259 (N_4259,N_3922,N_4190);
nand U4260 (N_4260,N_4189,N_3771);
nand U4261 (N_4261,N_4191,N_4068);
or U4262 (N_4262,N_3913,N_4122);
nand U4263 (N_4263,N_3717,N_4039);
xor U4264 (N_4264,N_4135,N_3719);
or U4265 (N_4265,N_3786,N_3631);
nand U4266 (N_4266,N_4174,N_3925);
nand U4267 (N_4267,N_3918,N_3835);
xnor U4268 (N_4268,N_4114,N_4081);
nor U4269 (N_4269,N_3605,N_3949);
or U4270 (N_4270,N_3948,N_3849);
nor U4271 (N_4271,N_4171,N_4104);
nand U4272 (N_4272,N_3984,N_3804);
nand U4273 (N_4273,N_3764,N_3668);
xnor U4274 (N_4274,N_4094,N_3821);
and U4275 (N_4275,N_3960,N_3630);
nor U4276 (N_4276,N_3999,N_4123);
nor U4277 (N_4277,N_3873,N_3812);
nor U4278 (N_4278,N_3846,N_3687);
and U4279 (N_4279,N_3801,N_3623);
and U4280 (N_4280,N_3715,N_3774);
xor U4281 (N_4281,N_4037,N_4028);
or U4282 (N_4282,N_3863,N_4007);
nand U4283 (N_4283,N_3738,N_3938);
or U4284 (N_4284,N_4169,N_4067);
and U4285 (N_4285,N_3845,N_3656);
nor U4286 (N_4286,N_3837,N_3758);
nand U4287 (N_4287,N_3665,N_4145);
and U4288 (N_4288,N_4020,N_3798);
nor U4289 (N_4289,N_3689,N_3964);
nor U4290 (N_4290,N_3794,N_3748);
nor U4291 (N_4291,N_3629,N_3737);
nor U4292 (N_4292,N_3632,N_3878);
xnor U4293 (N_4293,N_3881,N_3756);
and U4294 (N_4294,N_4073,N_3745);
nor U4295 (N_4295,N_4077,N_4160);
xnor U4296 (N_4296,N_3819,N_3751);
or U4297 (N_4297,N_4090,N_3790);
nand U4298 (N_4298,N_3886,N_4088);
or U4299 (N_4299,N_3998,N_3778);
and U4300 (N_4300,N_3727,N_3931);
nor U4301 (N_4301,N_3893,N_4117);
nand U4302 (N_4302,N_3664,N_3784);
or U4303 (N_4303,N_4177,N_4153);
or U4304 (N_4304,N_4198,N_3736);
or U4305 (N_4305,N_4095,N_4110);
or U4306 (N_4306,N_4098,N_3657);
or U4307 (N_4307,N_4188,N_3910);
nand U4308 (N_4308,N_3983,N_3997);
or U4309 (N_4309,N_3768,N_4144);
nor U4310 (N_4310,N_3683,N_3734);
and U4311 (N_4311,N_4091,N_3995);
nor U4312 (N_4312,N_4080,N_4140);
nand U4313 (N_4313,N_3760,N_4158);
or U4314 (N_4314,N_3808,N_4102);
nor U4315 (N_4315,N_4004,N_3871);
and U4316 (N_4316,N_3901,N_4009);
or U4317 (N_4317,N_3729,N_4053);
or U4318 (N_4318,N_4010,N_3606);
nor U4319 (N_4319,N_3967,N_3661);
or U4320 (N_4320,N_3847,N_3777);
nand U4321 (N_4321,N_4002,N_3912);
xnor U4322 (N_4322,N_3838,N_3672);
or U4323 (N_4323,N_3829,N_4109);
nand U4324 (N_4324,N_3993,N_3982);
nor U4325 (N_4325,N_3996,N_3647);
xnor U4326 (N_4326,N_3909,N_3939);
or U4327 (N_4327,N_4139,N_3969);
and U4328 (N_4328,N_3872,N_4118);
or U4329 (N_4329,N_3827,N_3900);
xnor U4330 (N_4330,N_3889,N_3811);
xnor U4331 (N_4331,N_4013,N_3936);
or U4332 (N_4332,N_4093,N_3958);
and U4333 (N_4333,N_4113,N_4116);
nand U4334 (N_4334,N_3628,N_4040);
or U4335 (N_4335,N_4065,N_3868);
nand U4336 (N_4336,N_3942,N_4172);
or U4337 (N_4337,N_4030,N_4143);
or U4338 (N_4338,N_4193,N_3724);
nand U4339 (N_4339,N_3805,N_3620);
nand U4340 (N_4340,N_3894,N_3601);
and U4341 (N_4341,N_3788,N_4034);
and U4342 (N_4342,N_3869,N_3722);
nor U4343 (N_4343,N_3670,N_4072);
nand U4344 (N_4344,N_3616,N_3703);
or U4345 (N_4345,N_3712,N_3655);
xnor U4346 (N_4346,N_3879,N_3787);
nor U4347 (N_4347,N_3841,N_4192);
xor U4348 (N_4348,N_3600,N_3702);
nand U4349 (N_4349,N_3860,N_3895);
nand U4350 (N_4350,N_4022,N_4120);
or U4351 (N_4351,N_3666,N_3684);
nand U4352 (N_4352,N_3789,N_3609);
and U4353 (N_4353,N_3816,N_3796);
and U4354 (N_4354,N_3933,N_3854);
or U4355 (N_4355,N_4026,N_3832);
xor U4356 (N_4356,N_3723,N_4149);
nor U4357 (N_4357,N_3897,N_3648);
or U4358 (N_4358,N_4105,N_4163);
or U4359 (N_4359,N_4108,N_3866);
and U4360 (N_4360,N_3698,N_4042);
and U4361 (N_4361,N_4173,N_3720);
and U4362 (N_4362,N_4057,N_3604);
nor U4363 (N_4363,N_3644,N_3815);
or U4364 (N_4364,N_4181,N_3639);
and U4365 (N_4365,N_4078,N_4005);
nand U4366 (N_4366,N_3682,N_3767);
and U4367 (N_4367,N_3769,N_3709);
nand U4368 (N_4368,N_4031,N_4035);
nand U4369 (N_4369,N_3864,N_3959);
and U4370 (N_4370,N_3716,N_3691);
nand U4371 (N_4371,N_3680,N_4045);
or U4372 (N_4372,N_3646,N_3859);
nand U4373 (N_4373,N_3785,N_3744);
or U4374 (N_4374,N_4076,N_3622);
or U4375 (N_4375,N_3621,N_3865);
nor U4376 (N_4376,N_3899,N_3898);
or U4377 (N_4377,N_3707,N_3705);
or U4378 (N_4378,N_3793,N_4154);
xnor U4379 (N_4379,N_3714,N_4041);
nor U4380 (N_4380,N_3905,N_3822);
nand U4381 (N_4381,N_3928,N_3856);
nand U4382 (N_4382,N_4106,N_4050);
nor U4383 (N_4383,N_4021,N_4125);
nand U4384 (N_4384,N_4047,N_3989);
or U4385 (N_4385,N_3799,N_3944);
or U4386 (N_4386,N_3802,N_3825);
xnor U4387 (N_4387,N_3685,N_3740);
nor U4388 (N_4388,N_3844,N_3943);
nand U4389 (N_4389,N_3932,N_3625);
nor U4390 (N_4390,N_3776,N_3914);
xor U4391 (N_4391,N_3617,N_4147);
nand U4392 (N_4392,N_3988,N_3669);
nand U4393 (N_4393,N_3710,N_3730);
nor U4394 (N_4394,N_3660,N_4137);
and U4395 (N_4395,N_4079,N_4089);
and U4396 (N_4396,N_3686,N_3902);
nand U4397 (N_4397,N_4199,N_4038);
nand U4398 (N_4398,N_3610,N_4187);
and U4399 (N_4399,N_3739,N_3941);
nand U4400 (N_4400,N_4097,N_3962);
or U4401 (N_4401,N_4165,N_3842);
nand U4402 (N_4402,N_4103,N_3921);
or U4403 (N_4403,N_3733,N_3795);
nor U4404 (N_4404,N_3651,N_4066);
nand U4405 (N_4405,N_4085,N_3862);
or U4406 (N_4406,N_4130,N_3792);
nand U4407 (N_4407,N_4027,N_3757);
nand U4408 (N_4408,N_3852,N_3728);
nand U4409 (N_4409,N_3635,N_3884);
and U4410 (N_4410,N_4025,N_3742);
or U4411 (N_4411,N_3979,N_3908);
xor U4412 (N_4412,N_3641,N_4096);
nand U4413 (N_4413,N_3851,N_3697);
or U4414 (N_4414,N_3653,N_3695);
or U4415 (N_4415,N_3711,N_3607);
and U4416 (N_4416,N_3762,N_3907);
xor U4417 (N_4417,N_3675,N_4128);
nor U4418 (N_4418,N_3976,N_4003);
and U4419 (N_4419,N_3618,N_3887);
nor U4420 (N_4420,N_3614,N_4043);
nand U4421 (N_4421,N_3857,N_3855);
or U4422 (N_4422,N_3735,N_4052);
nor U4423 (N_4423,N_4132,N_3917);
xor U4424 (N_4424,N_3761,N_3699);
nor U4425 (N_4425,N_3980,N_3935);
nand U4426 (N_4426,N_3986,N_3602);
or U4427 (N_4427,N_3924,N_3826);
and U4428 (N_4428,N_3985,N_3817);
xnor U4429 (N_4429,N_3883,N_3747);
and U4430 (N_4430,N_4157,N_3882);
nand U4431 (N_4431,N_3678,N_4044);
and U4432 (N_4432,N_4182,N_3934);
and U4433 (N_4433,N_4168,N_3840);
nand U4434 (N_4434,N_4148,N_3853);
nand U4435 (N_4435,N_3963,N_3612);
or U4436 (N_4436,N_4138,N_4011);
or U4437 (N_4437,N_3892,N_3818);
and U4438 (N_4438,N_3690,N_4074);
and U4439 (N_4439,N_3803,N_4121);
nand U4440 (N_4440,N_4186,N_3773);
nand U4441 (N_4441,N_3791,N_3991);
or U4442 (N_4442,N_3667,N_3903);
or U4443 (N_4443,N_3732,N_3955);
or U4444 (N_4444,N_4062,N_3741);
nand U4445 (N_4445,N_4061,N_3888);
and U4446 (N_4446,N_4115,N_4185);
nand U4447 (N_4447,N_3911,N_3940);
nor U4448 (N_4448,N_3783,N_3731);
nand U4449 (N_4449,N_4058,N_4071);
nor U4450 (N_4450,N_3643,N_3926);
and U4451 (N_4451,N_3929,N_3974);
and U4452 (N_4452,N_3677,N_3820);
nor U4453 (N_4453,N_4159,N_3721);
nor U4454 (N_4454,N_3896,N_3640);
nor U4455 (N_4455,N_4055,N_4017);
nand U4456 (N_4456,N_3746,N_4161);
nor U4457 (N_4457,N_3994,N_3877);
or U4458 (N_4458,N_3937,N_3945);
xnor U4459 (N_4459,N_4131,N_3700);
xor U4460 (N_4460,N_3800,N_3972);
and U4461 (N_4461,N_3650,N_4197);
nor U4462 (N_4462,N_4087,N_3885);
xnor U4463 (N_4463,N_3649,N_4111);
or U4464 (N_4464,N_3772,N_3916);
nand U4465 (N_4465,N_4124,N_3968);
or U4466 (N_4466,N_4018,N_4152);
and U4467 (N_4467,N_4183,N_4092);
xnor U4468 (N_4468,N_3681,N_3765);
xnor U4469 (N_4469,N_3965,N_3951);
nor U4470 (N_4470,N_4060,N_4150);
xnor U4471 (N_4471,N_3613,N_4141);
nand U4472 (N_4472,N_3813,N_3633);
xnor U4473 (N_4473,N_3930,N_3726);
nor U4474 (N_4474,N_3987,N_4129);
xnor U4475 (N_4475,N_3626,N_3634);
nand U4476 (N_4476,N_4179,N_4164);
nand U4477 (N_4477,N_3763,N_3619);
nand U4478 (N_4478,N_3694,N_4170);
and U4479 (N_4479,N_3927,N_3920);
nand U4480 (N_4480,N_3704,N_3915);
nand U4481 (N_4481,N_3797,N_4036);
nor U4482 (N_4482,N_4008,N_4162);
or U4483 (N_4483,N_4083,N_3718);
or U4484 (N_4484,N_4146,N_3608);
and U4485 (N_4485,N_4056,N_3843);
or U4486 (N_4486,N_3725,N_3671);
nor U4487 (N_4487,N_4107,N_3977);
nand U4488 (N_4488,N_4014,N_3603);
nor U4489 (N_4489,N_4024,N_3981);
xnor U4490 (N_4490,N_3961,N_3781);
nand U4491 (N_4491,N_3638,N_3759);
xnor U4492 (N_4492,N_4112,N_3875);
or U4493 (N_4493,N_3946,N_3906);
and U4494 (N_4494,N_3708,N_3679);
and U4495 (N_4495,N_4019,N_4176);
and U4496 (N_4496,N_4151,N_3947);
nand U4497 (N_4497,N_4180,N_3814);
nand U4498 (N_4498,N_3652,N_3890);
nor U4499 (N_4499,N_4070,N_3775);
or U4500 (N_4500,N_3955,N_3761);
and U4501 (N_4501,N_3836,N_4069);
nand U4502 (N_4502,N_3921,N_4168);
nand U4503 (N_4503,N_3884,N_3719);
and U4504 (N_4504,N_4098,N_4069);
or U4505 (N_4505,N_4132,N_3612);
and U4506 (N_4506,N_3895,N_3630);
nand U4507 (N_4507,N_3698,N_3739);
nand U4508 (N_4508,N_3807,N_4112);
and U4509 (N_4509,N_3819,N_4089);
or U4510 (N_4510,N_3667,N_3922);
or U4511 (N_4511,N_3819,N_4070);
or U4512 (N_4512,N_3631,N_3688);
xnor U4513 (N_4513,N_3831,N_4180);
or U4514 (N_4514,N_3609,N_3690);
nor U4515 (N_4515,N_4153,N_3961);
and U4516 (N_4516,N_4063,N_3613);
nor U4517 (N_4517,N_3893,N_4035);
or U4518 (N_4518,N_3692,N_3881);
or U4519 (N_4519,N_3787,N_3812);
and U4520 (N_4520,N_3643,N_4136);
xnor U4521 (N_4521,N_3731,N_4098);
and U4522 (N_4522,N_4097,N_4053);
or U4523 (N_4523,N_4129,N_4096);
xnor U4524 (N_4524,N_3919,N_3854);
nor U4525 (N_4525,N_3778,N_3883);
nand U4526 (N_4526,N_3836,N_4134);
nand U4527 (N_4527,N_4088,N_3618);
and U4528 (N_4528,N_3603,N_4026);
nand U4529 (N_4529,N_3761,N_3808);
nor U4530 (N_4530,N_4114,N_4179);
and U4531 (N_4531,N_3989,N_3935);
nor U4532 (N_4532,N_4095,N_4173);
or U4533 (N_4533,N_4117,N_3986);
and U4534 (N_4534,N_3929,N_4055);
and U4535 (N_4535,N_3644,N_3697);
nor U4536 (N_4536,N_4091,N_4108);
nand U4537 (N_4537,N_3871,N_3990);
nor U4538 (N_4538,N_3659,N_4180);
nor U4539 (N_4539,N_3659,N_3885);
or U4540 (N_4540,N_3972,N_4172);
and U4541 (N_4541,N_3827,N_4062);
nand U4542 (N_4542,N_4127,N_3722);
or U4543 (N_4543,N_3647,N_3740);
and U4544 (N_4544,N_3772,N_3779);
nor U4545 (N_4545,N_3847,N_3923);
xor U4546 (N_4546,N_3602,N_4014);
or U4547 (N_4547,N_3991,N_3851);
or U4548 (N_4548,N_3745,N_4185);
or U4549 (N_4549,N_3738,N_3765);
nand U4550 (N_4550,N_4063,N_3926);
or U4551 (N_4551,N_4165,N_3991);
or U4552 (N_4552,N_3815,N_3713);
nand U4553 (N_4553,N_4026,N_3838);
nand U4554 (N_4554,N_4084,N_3648);
and U4555 (N_4555,N_3757,N_3939);
and U4556 (N_4556,N_3799,N_3824);
nand U4557 (N_4557,N_4072,N_4058);
and U4558 (N_4558,N_3975,N_4122);
or U4559 (N_4559,N_3787,N_4104);
nand U4560 (N_4560,N_3947,N_3735);
or U4561 (N_4561,N_4041,N_4150);
nand U4562 (N_4562,N_3654,N_4023);
nor U4563 (N_4563,N_4141,N_3896);
or U4564 (N_4564,N_4065,N_4077);
nor U4565 (N_4565,N_3720,N_3816);
nand U4566 (N_4566,N_3763,N_4164);
nand U4567 (N_4567,N_3767,N_4065);
or U4568 (N_4568,N_3825,N_4171);
nand U4569 (N_4569,N_3761,N_4049);
nor U4570 (N_4570,N_3951,N_3695);
and U4571 (N_4571,N_3801,N_3701);
nor U4572 (N_4572,N_3625,N_4013);
nand U4573 (N_4573,N_4021,N_4157);
nor U4574 (N_4574,N_4139,N_3885);
and U4575 (N_4575,N_3918,N_3753);
or U4576 (N_4576,N_4153,N_3759);
nand U4577 (N_4577,N_4011,N_3876);
xnor U4578 (N_4578,N_3612,N_3738);
nor U4579 (N_4579,N_4042,N_3644);
or U4580 (N_4580,N_3640,N_4101);
nand U4581 (N_4581,N_3947,N_4154);
nor U4582 (N_4582,N_4084,N_3619);
or U4583 (N_4583,N_3979,N_3868);
nand U4584 (N_4584,N_3991,N_3728);
nor U4585 (N_4585,N_4007,N_3920);
and U4586 (N_4586,N_4095,N_4168);
xnor U4587 (N_4587,N_4020,N_3716);
nand U4588 (N_4588,N_4085,N_3792);
nor U4589 (N_4589,N_3863,N_4044);
and U4590 (N_4590,N_3960,N_3665);
or U4591 (N_4591,N_3998,N_3770);
or U4592 (N_4592,N_4006,N_3884);
or U4593 (N_4593,N_3823,N_4080);
nor U4594 (N_4594,N_4098,N_4053);
and U4595 (N_4595,N_3604,N_4157);
nor U4596 (N_4596,N_3828,N_4170);
and U4597 (N_4597,N_3658,N_4031);
or U4598 (N_4598,N_3840,N_4180);
or U4599 (N_4599,N_3715,N_3712);
nand U4600 (N_4600,N_3878,N_4108);
or U4601 (N_4601,N_3760,N_3614);
or U4602 (N_4602,N_3967,N_4101);
nor U4603 (N_4603,N_3684,N_3921);
and U4604 (N_4604,N_3784,N_3853);
nor U4605 (N_4605,N_4185,N_3971);
nand U4606 (N_4606,N_4094,N_3620);
nand U4607 (N_4607,N_4045,N_3783);
or U4608 (N_4608,N_4121,N_3711);
nand U4609 (N_4609,N_4050,N_4185);
nand U4610 (N_4610,N_4045,N_4120);
and U4611 (N_4611,N_4102,N_4062);
and U4612 (N_4612,N_4090,N_3784);
nor U4613 (N_4613,N_4057,N_3754);
nand U4614 (N_4614,N_3751,N_3780);
nor U4615 (N_4615,N_4131,N_4017);
and U4616 (N_4616,N_4183,N_4189);
or U4617 (N_4617,N_3645,N_3769);
nand U4618 (N_4618,N_3918,N_3685);
nand U4619 (N_4619,N_3634,N_3753);
and U4620 (N_4620,N_3757,N_4190);
nand U4621 (N_4621,N_4088,N_3790);
or U4622 (N_4622,N_3683,N_3839);
and U4623 (N_4623,N_4077,N_3672);
nand U4624 (N_4624,N_3666,N_3619);
nor U4625 (N_4625,N_3664,N_4000);
and U4626 (N_4626,N_3601,N_3910);
and U4627 (N_4627,N_3811,N_3803);
or U4628 (N_4628,N_3799,N_3728);
nand U4629 (N_4629,N_3878,N_3941);
nor U4630 (N_4630,N_4119,N_3677);
nand U4631 (N_4631,N_4047,N_3714);
or U4632 (N_4632,N_4036,N_3835);
nor U4633 (N_4633,N_3796,N_3741);
nand U4634 (N_4634,N_3934,N_3620);
nor U4635 (N_4635,N_4112,N_4083);
nand U4636 (N_4636,N_3785,N_4001);
or U4637 (N_4637,N_3923,N_3694);
and U4638 (N_4638,N_3799,N_4023);
and U4639 (N_4639,N_3904,N_4028);
nor U4640 (N_4640,N_4133,N_4062);
and U4641 (N_4641,N_4102,N_3726);
and U4642 (N_4642,N_4104,N_4042);
and U4643 (N_4643,N_4029,N_3925);
nor U4644 (N_4644,N_3815,N_3985);
nand U4645 (N_4645,N_3759,N_4185);
and U4646 (N_4646,N_3877,N_3610);
nand U4647 (N_4647,N_3974,N_4157);
xor U4648 (N_4648,N_3827,N_3627);
nand U4649 (N_4649,N_4134,N_3990);
xor U4650 (N_4650,N_3822,N_3993);
or U4651 (N_4651,N_3938,N_3970);
and U4652 (N_4652,N_3954,N_4108);
nor U4653 (N_4653,N_4120,N_3696);
and U4654 (N_4654,N_3797,N_4033);
and U4655 (N_4655,N_4198,N_4066);
xor U4656 (N_4656,N_3649,N_4031);
and U4657 (N_4657,N_3746,N_4045);
nor U4658 (N_4658,N_3719,N_3745);
nor U4659 (N_4659,N_3996,N_3875);
nor U4660 (N_4660,N_3905,N_3650);
nor U4661 (N_4661,N_4121,N_3724);
nand U4662 (N_4662,N_3690,N_4195);
or U4663 (N_4663,N_4022,N_3700);
nand U4664 (N_4664,N_4120,N_3948);
and U4665 (N_4665,N_3767,N_3731);
nor U4666 (N_4666,N_3686,N_3774);
or U4667 (N_4667,N_3671,N_4185);
nand U4668 (N_4668,N_4039,N_3627);
or U4669 (N_4669,N_3801,N_3808);
nand U4670 (N_4670,N_4156,N_4053);
nand U4671 (N_4671,N_4097,N_4073);
nand U4672 (N_4672,N_3723,N_3876);
nor U4673 (N_4673,N_4008,N_3902);
xnor U4674 (N_4674,N_4196,N_3926);
and U4675 (N_4675,N_3994,N_4098);
nor U4676 (N_4676,N_3866,N_3793);
nand U4677 (N_4677,N_4062,N_3649);
nor U4678 (N_4678,N_3626,N_3623);
nor U4679 (N_4679,N_3904,N_3868);
nor U4680 (N_4680,N_3710,N_3987);
or U4681 (N_4681,N_3631,N_3977);
and U4682 (N_4682,N_3613,N_4102);
nand U4683 (N_4683,N_4091,N_3858);
and U4684 (N_4684,N_3670,N_3991);
or U4685 (N_4685,N_3707,N_4085);
or U4686 (N_4686,N_3905,N_3947);
nor U4687 (N_4687,N_3920,N_3706);
and U4688 (N_4688,N_3930,N_3947);
and U4689 (N_4689,N_3608,N_3720);
nand U4690 (N_4690,N_4164,N_3691);
nor U4691 (N_4691,N_3608,N_3960);
and U4692 (N_4692,N_3699,N_3800);
nor U4693 (N_4693,N_3783,N_4016);
and U4694 (N_4694,N_3980,N_4090);
and U4695 (N_4695,N_3631,N_3613);
xnor U4696 (N_4696,N_3669,N_3793);
nor U4697 (N_4697,N_3876,N_3609);
and U4698 (N_4698,N_3892,N_4019);
and U4699 (N_4699,N_3772,N_4171);
nor U4700 (N_4700,N_3668,N_4102);
or U4701 (N_4701,N_3862,N_3945);
nor U4702 (N_4702,N_3998,N_3864);
and U4703 (N_4703,N_3806,N_4145);
or U4704 (N_4704,N_3613,N_3973);
nor U4705 (N_4705,N_3859,N_3827);
xnor U4706 (N_4706,N_4007,N_4146);
and U4707 (N_4707,N_4137,N_4048);
or U4708 (N_4708,N_4101,N_4028);
and U4709 (N_4709,N_3756,N_4118);
nand U4710 (N_4710,N_3843,N_3638);
nor U4711 (N_4711,N_4014,N_4028);
or U4712 (N_4712,N_4043,N_3814);
nor U4713 (N_4713,N_3915,N_3803);
nor U4714 (N_4714,N_4098,N_3837);
nor U4715 (N_4715,N_4121,N_3890);
or U4716 (N_4716,N_3964,N_3815);
xnor U4717 (N_4717,N_3775,N_3869);
and U4718 (N_4718,N_4098,N_4073);
nor U4719 (N_4719,N_3861,N_3679);
xnor U4720 (N_4720,N_3951,N_3943);
and U4721 (N_4721,N_4090,N_3639);
nor U4722 (N_4722,N_3965,N_4060);
and U4723 (N_4723,N_3789,N_3856);
or U4724 (N_4724,N_4048,N_4080);
nand U4725 (N_4725,N_4122,N_4183);
nand U4726 (N_4726,N_4104,N_4088);
nand U4727 (N_4727,N_3946,N_3649);
or U4728 (N_4728,N_4047,N_3752);
nand U4729 (N_4729,N_4172,N_3759);
nor U4730 (N_4730,N_3680,N_3906);
nand U4731 (N_4731,N_3737,N_3713);
or U4732 (N_4732,N_4168,N_3768);
and U4733 (N_4733,N_3765,N_3689);
and U4734 (N_4734,N_3892,N_4064);
or U4735 (N_4735,N_3687,N_4139);
nor U4736 (N_4736,N_4059,N_4130);
or U4737 (N_4737,N_3961,N_4120);
or U4738 (N_4738,N_3973,N_3684);
nand U4739 (N_4739,N_3714,N_4010);
xor U4740 (N_4740,N_3873,N_3841);
nor U4741 (N_4741,N_3791,N_3914);
or U4742 (N_4742,N_3765,N_3670);
nand U4743 (N_4743,N_3768,N_3842);
xor U4744 (N_4744,N_3695,N_3922);
or U4745 (N_4745,N_3712,N_3882);
and U4746 (N_4746,N_3883,N_3824);
nand U4747 (N_4747,N_3949,N_3737);
or U4748 (N_4748,N_3636,N_3799);
xnor U4749 (N_4749,N_3721,N_4173);
and U4750 (N_4750,N_3764,N_4185);
or U4751 (N_4751,N_3652,N_4088);
or U4752 (N_4752,N_4058,N_3674);
and U4753 (N_4753,N_3789,N_3802);
or U4754 (N_4754,N_4161,N_3832);
or U4755 (N_4755,N_3622,N_3867);
nand U4756 (N_4756,N_3798,N_3653);
and U4757 (N_4757,N_3926,N_3996);
nand U4758 (N_4758,N_4027,N_3887);
nor U4759 (N_4759,N_3699,N_3917);
or U4760 (N_4760,N_4188,N_4108);
or U4761 (N_4761,N_3939,N_3993);
nand U4762 (N_4762,N_3798,N_3630);
and U4763 (N_4763,N_3969,N_4043);
nor U4764 (N_4764,N_3630,N_3679);
nand U4765 (N_4765,N_3956,N_3781);
nand U4766 (N_4766,N_4078,N_3728);
nor U4767 (N_4767,N_4144,N_4058);
and U4768 (N_4768,N_3896,N_3972);
nand U4769 (N_4769,N_4014,N_3644);
or U4770 (N_4770,N_4039,N_3952);
or U4771 (N_4771,N_3799,N_4055);
and U4772 (N_4772,N_3712,N_3700);
nor U4773 (N_4773,N_3677,N_3764);
or U4774 (N_4774,N_4054,N_4108);
xor U4775 (N_4775,N_3998,N_4106);
or U4776 (N_4776,N_3680,N_3741);
nand U4777 (N_4777,N_3716,N_3873);
nand U4778 (N_4778,N_3710,N_4132);
or U4779 (N_4779,N_3609,N_3638);
nand U4780 (N_4780,N_4122,N_4119);
and U4781 (N_4781,N_3816,N_3866);
nor U4782 (N_4782,N_3992,N_3778);
and U4783 (N_4783,N_4089,N_4077);
nor U4784 (N_4784,N_3784,N_3793);
nor U4785 (N_4785,N_3941,N_3742);
or U4786 (N_4786,N_3837,N_3971);
nor U4787 (N_4787,N_4198,N_3715);
and U4788 (N_4788,N_4157,N_3774);
nand U4789 (N_4789,N_4151,N_4024);
or U4790 (N_4790,N_4037,N_3640);
nor U4791 (N_4791,N_4172,N_3732);
nand U4792 (N_4792,N_3607,N_4067);
nor U4793 (N_4793,N_4063,N_4075);
and U4794 (N_4794,N_4181,N_4167);
nor U4795 (N_4795,N_3801,N_3636);
nand U4796 (N_4796,N_3931,N_4108);
or U4797 (N_4797,N_4105,N_4194);
nor U4798 (N_4798,N_3992,N_3868);
nand U4799 (N_4799,N_3613,N_3856);
and U4800 (N_4800,N_4411,N_4733);
nor U4801 (N_4801,N_4267,N_4544);
nor U4802 (N_4802,N_4752,N_4684);
nor U4803 (N_4803,N_4424,N_4616);
or U4804 (N_4804,N_4521,N_4649);
nor U4805 (N_4805,N_4201,N_4788);
nand U4806 (N_4806,N_4564,N_4542);
and U4807 (N_4807,N_4703,N_4552);
nor U4808 (N_4808,N_4461,N_4712);
nand U4809 (N_4809,N_4233,N_4459);
nor U4810 (N_4810,N_4567,N_4429);
nor U4811 (N_4811,N_4454,N_4337);
nor U4812 (N_4812,N_4695,N_4549);
and U4813 (N_4813,N_4288,N_4401);
nor U4814 (N_4814,N_4642,N_4658);
nor U4815 (N_4815,N_4431,N_4646);
or U4816 (N_4816,N_4223,N_4210);
xnor U4817 (N_4817,N_4462,N_4230);
and U4818 (N_4818,N_4781,N_4395);
nand U4819 (N_4819,N_4204,N_4344);
nor U4820 (N_4820,N_4487,N_4770);
and U4821 (N_4821,N_4745,N_4691);
nand U4822 (N_4822,N_4301,N_4726);
nor U4823 (N_4823,N_4440,N_4696);
nor U4824 (N_4824,N_4479,N_4347);
and U4825 (N_4825,N_4207,N_4690);
or U4826 (N_4826,N_4506,N_4612);
and U4827 (N_4827,N_4309,N_4403);
nor U4828 (N_4828,N_4252,N_4764);
nand U4829 (N_4829,N_4596,N_4687);
or U4830 (N_4830,N_4650,N_4592);
nor U4831 (N_4831,N_4379,N_4334);
nor U4832 (N_4832,N_4465,N_4534);
nor U4833 (N_4833,N_4724,N_4546);
or U4834 (N_4834,N_4318,N_4212);
and U4835 (N_4835,N_4785,N_4372);
or U4836 (N_4836,N_4352,N_4746);
nor U4837 (N_4837,N_4485,N_4771);
nor U4838 (N_4838,N_4434,N_4317);
or U4839 (N_4839,N_4342,N_4216);
or U4840 (N_4840,N_4714,N_4773);
or U4841 (N_4841,N_4607,N_4340);
nand U4842 (N_4842,N_4550,N_4441);
xor U4843 (N_4843,N_4525,N_4271);
nand U4844 (N_4844,N_4772,N_4258);
nor U4845 (N_4845,N_4407,N_4576);
nand U4846 (N_4846,N_4548,N_4702);
and U4847 (N_4847,N_4200,N_4662);
nand U4848 (N_4848,N_4614,N_4219);
and U4849 (N_4849,N_4322,N_4728);
nand U4850 (N_4850,N_4275,N_4330);
and U4851 (N_4851,N_4541,N_4553);
and U4852 (N_4852,N_4523,N_4313);
and U4853 (N_4853,N_4300,N_4727);
and U4854 (N_4854,N_4613,N_4689);
nand U4855 (N_4855,N_4315,N_4756);
nand U4856 (N_4856,N_4621,N_4535);
nand U4857 (N_4857,N_4538,N_4452);
nor U4858 (N_4858,N_4493,N_4492);
or U4859 (N_4859,N_4566,N_4311);
nand U4860 (N_4860,N_4491,N_4617);
nand U4861 (N_4861,N_4758,N_4512);
nor U4862 (N_4862,N_4246,N_4448);
xnor U4863 (N_4863,N_4654,N_4326);
or U4864 (N_4864,N_4356,N_4398);
or U4865 (N_4865,N_4729,N_4355);
nand U4866 (N_4866,N_4648,N_4499);
and U4867 (N_4867,N_4672,N_4704);
nor U4868 (N_4868,N_4530,N_4244);
xor U4869 (N_4869,N_4470,N_4370);
nor U4870 (N_4870,N_4637,N_4765);
or U4871 (N_4871,N_4211,N_4639);
nor U4872 (N_4872,N_4447,N_4264);
nand U4873 (N_4873,N_4777,N_4604);
or U4874 (N_4874,N_4721,N_4477);
or U4875 (N_4875,N_4478,N_4725);
nand U4876 (N_4876,N_4786,N_4641);
or U4877 (N_4877,N_4511,N_4522);
nor U4878 (N_4878,N_4218,N_4547);
and U4879 (N_4879,N_4438,N_4577);
or U4880 (N_4880,N_4480,N_4673);
nand U4881 (N_4881,N_4240,N_4494);
nor U4882 (N_4882,N_4208,N_4296);
nand U4883 (N_4883,N_4519,N_4629);
nor U4884 (N_4884,N_4446,N_4775);
nand U4885 (N_4885,N_4738,N_4363);
nand U4886 (N_4886,N_4291,N_4780);
nand U4887 (N_4887,N_4466,N_4423);
xnor U4888 (N_4888,N_4283,N_4677);
nand U4889 (N_4889,N_4561,N_4625);
or U4890 (N_4890,N_4705,N_4268);
nand U4891 (N_4891,N_4560,N_4327);
nand U4892 (N_4892,N_4513,N_4536);
nand U4893 (N_4893,N_4473,N_4253);
nor U4894 (N_4894,N_4369,N_4720);
nand U4895 (N_4895,N_4715,N_4681);
nor U4896 (N_4896,N_4783,N_4586);
or U4897 (N_4897,N_4497,N_4394);
and U4898 (N_4898,N_4308,N_4338);
nor U4899 (N_4899,N_4333,N_4796);
or U4900 (N_4900,N_4782,N_4251);
xnor U4901 (N_4901,N_4631,N_4353);
or U4902 (N_4902,N_4261,N_4305);
nor U4903 (N_4903,N_4209,N_4217);
nor U4904 (N_4904,N_4555,N_4682);
and U4905 (N_4905,N_4382,N_4237);
nand U4906 (N_4906,N_4442,N_4391);
xor U4907 (N_4907,N_4412,N_4594);
or U4908 (N_4908,N_4659,N_4314);
and U4909 (N_4909,N_4471,N_4557);
or U4910 (N_4910,N_4761,N_4630);
and U4911 (N_4911,N_4573,N_4505);
xnor U4912 (N_4912,N_4793,N_4388);
or U4913 (N_4913,N_4601,N_4242);
nand U4914 (N_4914,N_4213,N_4375);
nor U4915 (N_4915,N_4508,N_4286);
nor U4916 (N_4916,N_4202,N_4414);
nand U4917 (N_4917,N_4651,N_4708);
or U4918 (N_4918,N_4257,N_4743);
nand U4919 (N_4919,N_4799,N_4439);
or U4920 (N_4920,N_4335,N_4609);
nand U4921 (N_4921,N_4362,N_4711);
xor U4922 (N_4922,N_4496,N_4437);
nor U4923 (N_4923,N_4475,N_4565);
nor U4924 (N_4924,N_4569,N_4774);
nand U4925 (N_4925,N_4716,N_4464);
and U4926 (N_4926,N_4776,N_4399);
nand U4927 (N_4927,N_4732,N_4556);
nand U4928 (N_4928,N_4749,N_4595);
xnor U4929 (N_4929,N_4409,N_4256);
nor U4930 (N_4930,N_4376,N_4384);
nor U4931 (N_4931,N_4387,N_4328);
or U4932 (N_4932,N_4323,N_4532);
nand U4933 (N_4933,N_4406,N_4762);
nor U4934 (N_4934,N_4250,N_4769);
nor U4935 (N_4935,N_4685,N_4510);
nor U4936 (N_4936,N_4664,N_4784);
and U4937 (N_4937,N_4647,N_4638);
or U4938 (N_4938,N_4221,N_4518);
nand U4939 (N_4939,N_4236,N_4348);
nand U4940 (N_4940,N_4377,N_4626);
nand U4941 (N_4941,N_4415,N_4490);
or U4942 (N_4942,N_4263,N_4226);
or U4943 (N_4943,N_4310,N_4768);
nor U4944 (N_4944,N_4710,N_4731);
and U4945 (N_4945,N_4618,N_4736);
nor U4946 (N_4946,N_4422,N_4635);
xnor U4947 (N_4947,N_4590,N_4287);
nand U4948 (N_4948,N_4366,N_4298);
nor U4949 (N_4949,N_4292,N_4605);
or U4950 (N_4950,N_4660,N_4306);
nand U4951 (N_4951,N_4599,N_4543);
nor U4952 (N_4952,N_4312,N_4591);
nand U4953 (N_4953,N_4767,N_4718);
nor U4954 (N_4954,N_4540,N_4674);
xor U4955 (N_4955,N_4336,N_4324);
nand U4956 (N_4956,N_4249,N_4572);
nand U4957 (N_4957,N_4484,N_4683);
nor U4958 (N_4958,N_4699,N_4717);
nand U4959 (N_4959,N_4449,N_4488);
nand U4960 (N_4960,N_4307,N_4329);
nor U4961 (N_4961,N_4627,N_4744);
or U4962 (N_4962,N_4486,N_4425);
and U4963 (N_4963,N_4500,N_4203);
nor U4964 (N_4964,N_4587,N_4750);
xor U4965 (N_4965,N_4432,N_4402);
xor U4966 (N_4966,N_4634,N_4443);
xnor U4967 (N_4967,N_4260,N_4467);
nor U4968 (N_4968,N_4719,N_4632);
or U4969 (N_4969,N_4241,N_4787);
nor U4970 (N_4970,N_4644,N_4483);
xor U4971 (N_4971,N_4220,N_4455);
or U4972 (N_4972,N_4740,N_4751);
nand U4973 (N_4973,N_4254,N_4516);
or U4974 (N_4974,N_4734,N_4420);
nor U4975 (N_4975,N_4515,N_4603);
xnor U4976 (N_4976,N_4610,N_4405);
or U4977 (N_4977,N_4795,N_4367);
or U4978 (N_4978,N_4284,N_4504);
or U4979 (N_4979,N_4694,N_4680);
and U4980 (N_4980,N_4289,N_4722);
nand U4981 (N_4981,N_4624,N_4619);
or U4982 (N_4982,N_4345,N_4574);
or U4983 (N_4983,N_4789,N_4670);
or U4984 (N_4984,N_4701,N_4528);
and U4985 (N_4985,N_4700,N_4418);
nand U4986 (N_4986,N_4693,N_4593);
xor U4987 (N_4987,N_4514,N_4757);
nand U4988 (N_4988,N_4224,N_4435);
or U4989 (N_4989,N_4606,N_4332);
nor U4990 (N_4990,N_4747,N_4481);
or U4991 (N_4991,N_4374,N_4274);
nor U4992 (N_4992,N_4688,N_4281);
and U4993 (N_4993,N_4381,N_4474);
or U4994 (N_4994,N_4341,N_4723);
and U4995 (N_4995,N_4400,N_4645);
nand U4996 (N_4996,N_4225,N_4293);
or U4997 (N_4997,N_4797,N_4667);
nand U4998 (N_4998,N_4735,N_4545);
nor U4999 (N_4999,N_4349,N_4299);
and U5000 (N_5000,N_4248,N_4350);
nor U5001 (N_5001,N_4419,N_4472);
nor U5002 (N_5002,N_4469,N_4503);
or U5003 (N_5003,N_4368,N_4359);
nor U5004 (N_5004,N_4668,N_4657);
nor U5005 (N_5005,N_4457,N_4529);
nor U5006 (N_5006,N_4669,N_4739);
or U5007 (N_5007,N_4779,N_4389);
nand U5008 (N_5008,N_4303,N_4417);
or U5009 (N_5009,N_4357,N_4526);
xor U5010 (N_5010,N_4214,N_4262);
nand U5011 (N_5011,N_4509,N_4222);
nor U5012 (N_5012,N_4235,N_4285);
nand U5013 (N_5013,N_4652,N_4458);
nand U5014 (N_5014,N_4663,N_4766);
nor U5015 (N_5015,N_4339,N_4297);
nand U5016 (N_5016,N_4302,N_4371);
nor U5017 (N_5017,N_4436,N_4623);
and U5018 (N_5018,N_4270,N_4451);
nor U5019 (N_5019,N_4378,N_4231);
xnor U5020 (N_5020,N_4794,N_4571);
or U5021 (N_5021,N_4255,N_4445);
nand U5022 (N_5022,N_4247,N_4570);
nor U5023 (N_5023,N_4498,N_4760);
and U5024 (N_5024,N_4427,N_4737);
xor U5025 (N_5025,N_4206,N_4597);
nand U5026 (N_5026,N_4205,N_4551);
or U5027 (N_5027,N_4383,N_4562);
nor U5028 (N_5028,N_4239,N_4468);
xnor U5029 (N_5029,N_4580,N_4321);
and U5030 (N_5030,N_4354,N_4581);
or U5031 (N_5031,N_4489,N_4450);
nand U5032 (N_5032,N_4234,N_4527);
and U5033 (N_5033,N_4707,N_4759);
nand U5034 (N_5034,N_4568,N_4393);
and U5035 (N_5035,N_4533,N_4421);
or U5036 (N_5036,N_4265,N_4665);
nand U5037 (N_5037,N_4410,N_4628);
and U5038 (N_5038,N_4476,N_4495);
xor U5039 (N_5039,N_4404,N_4413);
nor U5040 (N_5040,N_4295,N_4748);
or U5041 (N_5041,N_4358,N_4396);
or U5042 (N_5042,N_4675,N_4578);
nor U5043 (N_5043,N_4697,N_4360);
or U5044 (N_5044,N_4280,N_4582);
nor U5045 (N_5045,N_4640,N_4228);
nand U5046 (N_5046,N_4790,N_4713);
or U5047 (N_5047,N_4331,N_4351);
nor U5048 (N_5048,N_4386,N_4430);
and U5049 (N_5049,N_4380,N_4277);
or U5050 (N_5050,N_4778,N_4755);
nor U5051 (N_5051,N_4463,N_4453);
and U5052 (N_5052,N_4502,N_4622);
nor U5053 (N_5053,N_4365,N_4742);
xnor U5054 (N_5054,N_4278,N_4537);
and U5055 (N_5055,N_4215,N_4686);
nand U5056 (N_5056,N_4584,N_4575);
or U5057 (N_5057,N_4245,N_4679);
and U5058 (N_5058,N_4276,N_4266);
nor U5059 (N_5059,N_4373,N_4279);
or U5060 (N_5060,N_4428,N_4539);
and U5061 (N_5061,N_4671,N_4554);
and U5062 (N_5062,N_4456,N_4583);
or U5063 (N_5063,N_4602,N_4730);
nand U5064 (N_5064,N_4433,N_4643);
nor U5065 (N_5065,N_4319,N_4408);
nand U5066 (N_5066,N_4692,N_4661);
or U5067 (N_5067,N_4589,N_4559);
or U5068 (N_5068,N_4608,N_4792);
nor U5069 (N_5069,N_4524,N_4259);
or U5070 (N_5070,N_4588,N_4709);
nand U5071 (N_5071,N_4392,N_4364);
or U5072 (N_5072,N_4232,N_4678);
nand U5073 (N_5073,N_4754,N_4282);
nor U5074 (N_5074,N_4753,N_4698);
nand U5075 (N_5075,N_4666,N_4227);
nand U5076 (N_5076,N_4294,N_4238);
nand U5077 (N_5077,N_4229,N_4763);
or U5078 (N_5078,N_4520,N_4390);
nor U5079 (N_5079,N_4653,N_4444);
or U5080 (N_5080,N_4517,N_4558);
and U5081 (N_5081,N_4304,N_4585);
and U5082 (N_5082,N_4273,N_4460);
nand U5083 (N_5083,N_4426,N_4385);
xnor U5084 (N_5084,N_4361,N_4290);
nor U5085 (N_5085,N_4791,N_4343);
xor U5086 (N_5086,N_4531,N_4706);
and U5087 (N_5087,N_4611,N_4316);
or U5088 (N_5088,N_4636,N_4579);
nand U5089 (N_5089,N_4243,N_4269);
nand U5090 (N_5090,N_4507,N_4563);
nor U5091 (N_5091,N_4416,N_4272);
and U5092 (N_5092,N_4633,N_4482);
nor U5093 (N_5093,N_4397,N_4656);
xor U5094 (N_5094,N_4798,N_4676);
and U5095 (N_5095,N_4615,N_4620);
or U5096 (N_5096,N_4325,N_4346);
nand U5097 (N_5097,N_4320,N_4501);
nor U5098 (N_5098,N_4655,N_4741);
and U5099 (N_5099,N_4598,N_4600);
xnor U5100 (N_5100,N_4641,N_4356);
nand U5101 (N_5101,N_4524,N_4449);
and U5102 (N_5102,N_4321,N_4483);
nor U5103 (N_5103,N_4745,N_4674);
or U5104 (N_5104,N_4657,N_4256);
or U5105 (N_5105,N_4442,N_4588);
and U5106 (N_5106,N_4664,N_4372);
xor U5107 (N_5107,N_4793,N_4286);
and U5108 (N_5108,N_4727,N_4389);
nand U5109 (N_5109,N_4284,N_4441);
or U5110 (N_5110,N_4202,N_4602);
and U5111 (N_5111,N_4574,N_4298);
nor U5112 (N_5112,N_4702,N_4266);
nor U5113 (N_5113,N_4583,N_4614);
nor U5114 (N_5114,N_4648,N_4682);
nand U5115 (N_5115,N_4297,N_4383);
nor U5116 (N_5116,N_4345,N_4755);
and U5117 (N_5117,N_4627,N_4593);
or U5118 (N_5118,N_4223,N_4442);
nand U5119 (N_5119,N_4310,N_4694);
or U5120 (N_5120,N_4263,N_4666);
xnor U5121 (N_5121,N_4233,N_4490);
nor U5122 (N_5122,N_4392,N_4214);
and U5123 (N_5123,N_4554,N_4326);
and U5124 (N_5124,N_4721,N_4295);
and U5125 (N_5125,N_4442,N_4200);
nand U5126 (N_5126,N_4345,N_4743);
xnor U5127 (N_5127,N_4449,N_4590);
nor U5128 (N_5128,N_4427,N_4591);
and U5129 (N_5129,N_4679,N_4422);
nor U5130 (N_5130,N_4512,N_4264);
xnor U5131 (N_5131,N_4458,N_4741);
nand U5132 (N_5132,N_4228,N_4557);
nor U5133 (N_5133,N_4208,N_4234);
nor U5134 (N_5134,N_4787,N_4478);
and U5135 (N_5135,N_4710,N_4528);
or U5136 (N_5136,N_4776,N_4537);
nor U5137 (N_5137,N_4254,N_4230);
nand U5138 (N_5138,N_4728,N_4581);
and U5139 (N_5139,N_4757,N_4538);
nand U5140 (N_5140,N_4762,N_4450);
xor U5141 (N_5141,N_4727,N_4465);
and U5142 (N_5142,N_4644,N_4229);
nand U5143 (N_5143,N_4684,N_4728);
or U5144 (N_5144,N_4662,N_4628);
nor U5145 (N_5145,N_4543,N_4445);
nand U5146 (N_5146,N_4453,N_4479);
xnor U5147 (N_5147,N_4245,N_4578);
nor U5148 (N_5148,N_4660,N_4799);
and U5149 (N_5149,N_4520,N_4752);
or U5150 (N_5150,N_4635,N_4627);
or U5151 (N_5151,N_4477,N_4717);
nor U5152 (N_5152,N_4260,N_4377);
or U5153 (N_5153,N_4437,N_4746);
nand U5154 (N_5154,N_4461,N_4424);
nand U5155 (N_5155,N_4681,N_4235);
and U5156 (N_5156,N_4434,N_4512);
or U5157 (N_5157,N_4514,N_4232);
and U5158 (N_5158,N_4252,N_4241);
and U5159 (N_5159,N_4562,N_4634);
or U5160 (N_5160,N_4769,N_4789);
nor U5161 (N_5161,N_4350,N_4234);
or U5162 (N_5162,N_4441,N_4641);
and U5163 (N_5163,N_4460,N_4568);
or U5164 (N_5164,N_4376,N_4370);
or U5165 (N_5165,N_4790,N_4510);
nor U5166 (N_5166,N_4625,N_4469);
nand U5167 (N_5167,N_4688,N_4341);
or U5168 (N_5168,N_4522,N_4692);
and U5169 (N_5169,N_4435,N_4568);
nand U5170 (N_5170,N_4749,N_4326);
or U5171 (N_5171,N_4626,N_4268);
or U5172 (N_5172,N_4277,N_4360);
and U5173 (N_5173,N_4723,N_4473);
nor U5174 (N_5174,N_4777,N_4499);
and U5175 (N_5175,N_4388,N_4465);
or U5176 (N_5176,N_4313,N_4276);
nand U5177 (N_5177,N_4564,N_4648);
and U5178 (N_5178,N_4559,N_4351);
and U5179 (N_5179,N_4604,N_4633);
or U5180 (N_5180,N_4627,N_4732);
or U5181 (N_5181,N_4350,N_4566);
or U5182 (N_5182,N_4523,N_4376);
or U5183 (N_5183,N_4210,N_4202);
or U5184 (N_5184,N_4397,N_4474);
and U5185 (N_5185,N_4349,N_4738);
nand U5186 (N_5186,N_4462,N_4297);
nor U5187 (N_5187,N_4355,N_4359);
and U5188 (N_5188,N_4291,N_4584);
or U5189 (N_5189,N_4592,N_4583);
or U5190 (N_5190,N_4541,N_4774);
and U5191 (N_5191,N_4691,N_4224);
or U5192 (N_5192,N_4715,N_4649);
or U5193 (N_5193,N_4797,N_4657);
nor U5194 (N_5194,N_4703,N_4433);
and U5195 (N_5195,N_4257,N_4494);
xnor U5196 (N_5196,N_4368,N_4403);
and U5197 (N_5197,N_4361,N_4253);
and U5198 (N_5198,N_4772,N_4519);
and U5199 (N_5199,N_4570,N_4753);
or U5200 (N_5200,N_4728,N_4485);
xnor U5201 (N_5201,N_4591,N_4500);
or U5202 (N_5202,N_4383,N_4766);
nand U5203 (N_5203,N_4344,N_4585);
nand U5204 (N_5204,N_4778,N_4788);
nor U5205 (N_5205,N_4405,N_4202);
and U5206 (N_5206,N_4593,N_4298);
and U5207 (N_5207,N_4204,N_4560);
or U5208 (N_5208,N_4507,N_4560);
and U5209 (N_5209,N_4315,N_4542);
nor U5210 (N_5210,N_4710,N_4277);
or U5211 (N_5211,N_4211,N_4201);
nand U5212 (N_5212,N_4479,N_4419);
or U5213 (N_5213,N_4470,N_4230);
nor U5214 (N_5214,N_4710,N_4306);
xnor U5215 (N_5215,N_4369,N_4463);
and U5216 (N_5216,N_4469,N_4690);
nand U5217 (N_5217,N_4482,N_4613);
nand U5218 (N_5218,N_4286,N_4732);
or U5219 (N_5219,N_4640,N_4777);
or U5220 (N_5220,N_4674,N_4205);
and U5221 (N_5221,N_4430,N_4717);
xor U5222 (N_5222,N_4751,N_4798);
or U5223 (N_5223,N_4319,N_4573);
or U5224 (N_5224,N_4415,N_4226);
nor U5225 (N_5225,N_4204,N_4799);
nand U5226 (N_5226,N_4424,N_4744);
nand U5227 (N_5227,N_4788,N_4572);
or U5228 (N_5228,N_4791,N_4434);
or U5229 (N_5229,N_4371,N_4560);
nand U5230 (N_5230,N_4387,N_4687);
nor U5231 (N_5231,N_4509,N_4475);
nor U5232 (N_5232,N_4515,N_4487);
nand U5233 (N_5233,N_4345,N_4520);
and U5234 (N_5234,N_4616,N_4306);
and U5235 (N_5235,N_4427,N_4446);
xnor U5236 (N_5236,N_4526,N_4510);
nor U5237 (N_5237,N_4764,N_4346);
and U5238 (N_5238,N_4313,N_4771);
nand U5239 (N_5239,N_4464,N_4266);
nor U5240 (N_5240,N_4317,N_4584);
nand U5241 (N_5241,N_4359,N_4707);
and U5242 (N_5242,N_4610,N_4742);
or U5243 (N_5243,N_4722,N_4386);
and U5244 (N_5244,N_4794,N_4405);
xor U5245 (N_5245,N_4636,N_4250);
or U5246 (N_5246,N_4423,N_4446);
xnor U5247 (N_5247,N_4531,N_4663);
nand U5248 (N_5248,N_4490,N_4643);
nand U5249 (N_5249,N_4696,N_4521);
and U5250 (N_5250,N_4471,N_4213);
nor U5251 (N_5251,N_4561,N_4667);
and U5252 (N_5252,N_4600,N_4230);
or U5253 (N_5253,N_4535,N_4644);
or U5254 (N_5254,N_4213,N_4301);
and U5255 (N_5255,N_4606,N_4207);
and U5256 (N_5256,N_4553,N_4510);
nand U5257 (N_5257,N_4239,N_4264);
and U5258 (N_5258,N_4612,N_4317);
and U5259 (N_5259,N_4420,N_4574);
xnor U5260 (N_5260,N_4646,N_4429);
xor U5261 (N_5261,N_4524,N_4342);
and U5262 (N_5262,N_4616,N_4566);
xor U5263 (N_5263,N_4304,N_4645);
nand U5264 (N_5264,N_4410,N_4512);
and U5265 (N_5265,N_4785,N_4333);
and U5266 (N_5266,N_4756,N_4730);
or U5267 (N_5267,N_4514,N_4654);
nand U5268 (N_5268,N_4439,N_4618);
or U5269 (N_5269,N_4683,N_4210);
and U5270 (N_5270,N_4773,N_4508);
or U5271 (N_5271,N_4527,N_4424);
nor U5272 (N_5272,N_4717,N_4457);
and U5273 (N_5273,N_4646,N_4208);
and U5274 (N_5274,N_4242,N_4636);
and U5275 (N_5275,N_4650,N_4523);
nor U5276 (N_5276,N_4666,N_4270);
nor U5277 (N_5277,N_4235,N_4267);
nand U5278 (N_5278,N_4440,N_4798);
and U5279 (N_5279,N_4363,N_4638);
and U5280 (N_5280,N_4560,N_4425);
nor U5281 (N_5281,N_4509,N_4250);
or U5282 (N_5282,N_4610,N_4659);
and U5283 (N_5283,N_4576,N_4276);
nand U5284 (N_5284,N_4254,N_4215);
nor U5285 (N_5285,N_4615,N_4206);
nand U5286 (N_5286,N_4622,N_4773);
nand U5287 (N_5287,N_4650,N_4212);
nor U5288 (N_5288,N_4620,N_4732);
nor U5289 (N_5289,N_4439,N_4250);
nand U5290 (N_5290,N_4792,N_4447);
nor U5291 (N_5291,N_4538,N_4214);
or U5292 (N_5292,N_4372,N_4211);
nor U5293 (N_5293,N_4400,N_4393);
or U5294 (N_5294,N_4749,N_4561);
nor U5295 (N_5295,N_4327,N_4500);
nor U5296 (N_5296,N_4434,N_4366);
and U5297 (N_5297,N_4712,N_4310);
xor U5298 (N_5298,N_4492,N_4697);
nand U5299 (N_5299,N_4281,N_4672);
or U5300 (N_5300,N_4219,N_4738);
or U5301 (N_5301,N_4231,N_4222);
nor U5302 (N_5302,N_4346,N_4581);
and U5303 (N_5303,N_4314,N_4449);
xnor U5304 (N_5304,N_4724,N_4621);
or U5305 (N_5305,N_4750,N_4766);
and U5306 (N_5306,N_4342,N_4719);
nor U5307 (N_5307,N_4443,N_4524);
and U5308 (N_5308,N_4318,N_4563);
or U5309 (N_5309,N_4651,N_4308);
and U5310 (N_5310,N_4605,N_4387);
xnor U5311 (N_5311,N_4692,N_4484);
nand U5312 (N_5312,N_4374,N_4265);
nor U5313 (N_5313,N_4442,N_4648);
nand U5314 (N_5314,N_4602,N_4366);
or U5315 (N_5315,N_4537,N_4683);
nor U5316 (N_5316,N_4492,N_4635);
or U5317 (N_5317,N_4460,N_4534);
nand U5318 (N_5318,N_4453,N_4327);
nor U5319 (N_5319,N_4633,N_4489);
or U5320 (N_5320,N_4287,N_4761);
nand U5321 (N_5321,N_4275,N_4484);
and U5322 (N_5322,N_4603,N_4697);
or U5323 (N_5323,N_4507,N_4282);
and U5324 (N_5324,N_4661,N_4335);
and U5325 (N_5325,N_4233,N_4537);
nand U5326 (N_5326,N_4511,N_4572);
or U5327 (N_5327,N_4205,N_4320);
nor U5328 (N_5328,N_4551,N_4420);
nor U5329 (N_5329,N_4719,N_4544);
or U5330 (N_5330,N_4758,N_4635);
or U5331 (N_5331,N_4602,N_4265);
xor U5332 (N_5332,N_4299,N_4233);
nand U5333 (N_5333,N_4463,N_4225);
and U5334 (N_5334,N_4554,N_4365);
and U5335 (N_5335,N_4482,N_4634);
and U5336 (N_5336,N_4329,N_4638);
nand U5337 (N_5337,N_4352,N_4564);
xor U5338 (N_5338,N_4552,N_4713);
or U5339 (N_5339,N_4337,N_4442);
nand U5340 (N_5340,N_4788,N_4620);
xnor U5341 (N_5341,N_4203,N_4424);
nor U5342 (N_5342,N_4733,N_4346);
or U5343 (N_5343,N_4434,N_4662);
and U5344 (N_5344,N_4534,N_4637);
nor U5345 (N_5345,N_4418,N_4555);
or U5346 (N_5346,N_4557,N_4277);
or U5347 (N_5347,N_4274,N_4723);
and U5348 (N_5348,N_4727,N_4555);
nand U5349 (N_5349,N_4567,N_4565);
nand U5350 (N_5350,N_4317,N_4742);
nor U5351 (N_5351,N_4505,N_4694);
and U5352 (N_5352,N_4680,N_4585);
nand U5353 (N_5353,N_4343,N_4651);
xor U5354 (N_5354,N_4422,N_4610);
nor U5355 (N_5355,N_4252,N_4269);
and U5356 (N_5356,N_4224,N_4307);
and U5357 (N_5357,N_4259,N_4420);
nor U5358 (N_5358,N_4524,N_4689);
nor U5359 (N_5359,N_4780,N_4262);
or U5360 (N_5360,N_4421,N_4333);
and U5361 (N_5361,N_4654,N_4269);
nand U5362 (N_5362,N_4389,N_4676);
or U5363 (N_5363,N_4517,N_4335);
or U5364 (N_5364,N_4598,N_4670);
or U5365 (N_5365,N_4705,N_4315);
nand U5366 (N_5366,N_4206,N_4443);
nor U5367 (N_5367,N_4563,N_4663);
nor U5368 (N_5368,N_4339,N_4251);
nor U5369 (N_5369,N_4611,N_4277);
xnor U5370 (N_5370,N_4684,N_4687);
or U5371 (N_5371,N_4269,N_4696);
and U5372 (N_5372,N_4273,N_4209);
or U5373 (N_5373,N_4565,N_4349);
nand U5374 (N_5374,N_4241,N_4465);
nor U5375 (N_5375,N_4634,N_4623);
nand U5376 (N_5376,N_4747,N_4416);
nor U5377 (N_5377,N_4295,N_4467);
nand U5378 (N_5378,N_4740,N_4257);
and U5379 (N_5379,N_4211,N_4745);
and U5380 (N_5380,N_4403,N_4686);
or U5381 (N_5381,N_4751,N_4544);
or U5382 (N_5382,N_4278,N_4684);
nand U5383 (N_5383,N_4284,N_4641);
nand U5384 (N_5384,N_4329,N_4293);
nor U5385 (N_5385,N_4337,N_4429);
xnor U5386 (N_5386,N_4459,N_4601);
or U5387 (N_5387,N_4353,N_4730);
nor U5388 (N_5388,N_4523,N_4292);
nand U5389 (N_5389,N_4243,N_4637);
nand U5390 (N_5390,N_4485,N_4572);
nand U5391 (N_5391,N_4551,N_4716);
or U5392 (N_5392,N_4205,N_4799);
and U5393 (N_5393,N_4457,N_4692);
nand U5394 (N_5394,N_4294,N_4268);
nand U5395 (N_5395,N_4228,N_4602);
nand U5396 (N_5396,N_4780,N_4517);
xor U5397 (N_5397,N_4493,N_4390);
nor U5398 (N_5398,N_4241,N_4614);
nor U5399 (N_5399,N_4397,N_4282);
nor U5400 (N_5400,N_5309,N_4949);
and U5401 (N_5401,N_5300,N_5042);
nand U5402 (N_5402,N_4865,N_5068);
nand U5403 (N_5403,N_5319,N_5054);
and U5404 (N_5404,N_5194,N_4805);
nor U5405 (N_5405,N_4807,N_5182);
and U5406 (N_5406,N_5165,N_4849);
xor U5407 (N_5407,N_5126,N_5388);
nor U5408 (N_5408,N_5225,N_4830);
nand U5409 (N_5409,N_5084,N_4932);
nor U5410 (N_5410,N_5318,N_5022);
or U5411 (N_5411,N_5185,N_5003);
nand U5412 (N_5412,N_4973,N_4961);
and U5413 (N_5413,N_5023,N_4861);
and U5414 (N_5414,N_5016,N_5017);
or U5415 (N_5415,N_5273,N_5202);
and U5416 (N_5416,N_5232,N_5020);
nor U5417 (N_5417,N_5210,N_5127);
nor U5418 (N_5418,N_5006,N_5349);
nand U5419 (N_5419,N_5274,N_4968);
nand U5420 (N_5420,N_4903,N_5242);
and U5421 (N_5421,N_4819,N_5290);
and U5422 (N_5422,N_5164,N_5154);
and U5423 (N_5423,N_4917,N_4928);
nand U5424 (N_5424,N_5222,N_5078);
nor U5425 (N_5425,N_5293,N_5332);
or U5426 (N_5426,N_4842,N_4919);
and U5427 (N_5427,N_5088,N_4889);
or U5428 (N_5428,N_5122,N_4895);
nor U5429 (N_5429,N_5052,N_4952);
or U5430 (N_5430,N_5097,N_5179);
nor U5431 (N_5431,N_4839,N_5348);
and U5432 (N_5432,N_4974,N_5373);
xnor U5433 (N_5433,N_5099,N_5163);
nor U5434 (N_5434,N_5195,N_5077);
or U5435 (N_5435,N_5105,N_4915);
nand U5436 (N_5436,N_5385,N_4984);
nor U5437 (N_5437,N_4902,N_4951);
xnor U5438 (N_5438,N_5188,N_5158);
and U5439 (N_5439,N_5066,N_4906);
nor U5440 (N_5440,N_5303,N_5144);
or U5441 (N_5441,N_4815,N_5116);
nor U5442 (N_5442,N_4965,N_5346);
nor U5443 (N_5443,N_5050,N_5364);
or U5444 (N_5444,N_5313,N_4986);
nor U5445 (N_5445,N_5262,N_4810);
nand U5446 (N_5446,N_4963,N_5229);
and U5447 (N_5447,N_5245,N_4901);
and U5448 (N_5448,N_4890,N_5033);
and U5449 (N_5449,N_4851,N_5167);
nor U5450 (N_5450,N_5329,N_5384);
nand U5451 (N_5451,N_4884,N_5286);
nor U5452 (N_5452,N_5369,N_5252);
nor U5453 (N_5453,N_4898,N_5360);
nand U5454 (N_5454,N_4988,N_5362);
nand U5455 (N_5455,N_5184,N_5111);
nor U5456 (N_5456,N_5123,N_5287);
xnor U5457 (N_5457,N_5150,N_5135);
and U5458 (N_5458,N_4991,N_4858);
or U5459 (N_5459,N_4853,N_4883);
nand U5460 (N_5460,N_5342,N_4875);
nand U5461 (N_5461,N_5014,N_5043);
and U5462 (N_5462,N_5231,N_4960);
nor U5463 (N_5463,N_4941,N_5353);
or U5464 (N_5464,N_4891,N_4833);
and U5465 (N_5465,N_5024,N_5272);
xor U5466 (N_5466,N_5377,N_5219);
nor U5467 (N_5467,N_5217,N_4897);
or U5468 (N_5468,N_5086,N_5170);
or U5469 (N_5469,N_5314,N_5083);
or U5470 (N_5470,N_5302,N_4876);
and U5471 (N_5471,N_5098,N_5255);
and U5472 (N_5472,N_4967,N_4801);
nand U5473 (N_5473,N_5117,N_4878);
nor U5474 (N_5474,N_5007,N_4940);
or U5475 (N_5475,N_5000,N_5338);
nor U5476 (N_5476,N_5398,N_5191);
nor U5477 (N_5477,N_5056,N_5264);
nor U5478 (N_5478,N_4863,N_5193);
or U5479 (N_5479,N_5204,N_5399);
nor U5480 (N_5480,N_5028,N_4935);
and U5481 (N_5481,N_4855,N_5258);
or U5482 (N_5482,N_5048,N_4934);
and U5483 (N_5483,N_5376,N_5331);
nand U5484 (N_5484,N_5240,N_4859);
nand U5485 (N_5485,N_5027,N_5207);
and U5486 (N_5486,N_5354,N_4920);
nand U5487 (N_5487,N_5323,N_5128);
or U5488 (N_5488,N_5206,N_5366);
and U5489 (N_5489,N_4848,N_5269);
and U5490 (N_5490,N_5280,N_4956);
or U5491 (N_5491,N_5008,N_5352);
and U5492 (N_5492,N_5254,N_4995);
nand U5493 (N_5493,N_4983,N_5213);
nor U5494 (N_5494,N_5397,N_5134);
nor U5495 (N_5495,N_4845,N_5211);
or U5496 (N_5496,N_4981,N_5396);
or U5497 (N_5497,N_5316,N_4814);
or U5498 (N_5498,N_4894,N_5291);
nand U5499 (N_5499,N_5257,N_5114);
nor U5500 (N_5500,N_5103,N_5201);
nor U5501 (N_5501,N_5070,N_5351);
nand U5502 (N_5502,N_4809,N_4955);
and U5503 (N_5503,N_5214,N_5104);
or U5504 (N_5504,N_5238,N_4930);
xnor U5505 (N_5505,N_4971,N_5013);
or U5506 (N_5506,N_5367,N_5198);
xor U5507 (N_5507,N_5282,N_4804);
nor U5508 (N_5508,N_5289,N_4931);
or U5509 (N_5509,N_4850,N_5251);
and U5510 (N_5510,N_5386,N_5228);
nor U5511 (N_5511,N_5159,N_5005);
nand U5512 (N_5512,N_4912,N_5002);
nand U5513 (N_5513,N_4877,N_5069);
nor U5514 (N_5514,N_5139,N_4905);
nand U5515 (N_5515,N_5141,N_5259);
nand U5516 (N_5516,N_4882,N_5230);
and U5517 (N_5517,N_5315,N_4926);
or U5518 (N_5518,N_5326,N_4909);
nand U5519 (N_5519,N_4892,N_5243);
nand U5520 (N_5520,N_5328,N_4862);
nor U5521 (N_5521,N_5079,N_4871);
nor U5522 (N_5522,N_4914,N_5196);
nand U5523 (N_5523,N_5391,N_4911);
and U5524 (N_5524,N_5040,N_5010);
nand U5525 (N_5525,N_5039,N_5037);
and U5526 (N_5526,N_4860,N_4840);
or U5527 (N_5527,N_5160,N_5320);
xor U5528 (N_5528,N_5368,N_5265);
nor U5529 (N_5529,N_4993,N_4852);
nor U5530 (N_5530,N_4990,N_4837);
and U5531 (N_5531,N_4831,N_5284);
or U5532 (N_5532,N_5345,N_5142);
or U5533 (N_5533,N_5235,N_4950);
nand U5534 (N_5534,N_5018,N_5044);
xnor U5535 (N_5535,N_4998,N_5085);
nand U5536 (N_5536,N_4899,N_5246);
or U5537 (N_5537,N_4966,N_4887);
and U5538 (N_5538,N_4856,N_4812);
nand U5539 (N_5539,N_4997,N_5118);
nor U5540 (N_5540,N_4969,N_4907);
nand U5541 (N_5541,N_5339,N_5394);
nand U5542 (N_5542,N_5094,N_5183);
nor U5543 (N_5543,N_4854,N_5370);
or U5544 (N_5544,N_5268,N_5059);
and U5545 (N_5545,N_5120,N_5046);
xnor U5546 (N_5546,N_5301,N_5026);
or U5547 (N_5547,N_5087,N_5296);
or U5548 (N_5548,N_5172,N_5299);
xnor U5549 (N_5549,N_5067,N_5168);
and U5550 (N_5550,N_4835,N_4885);
nor U5551 (N_5551,N_5381,N_4923);
nor U5552 (N_5552,N_5261,N_4948);
xor U5553 (N_5553,N_4953,N_5270);
nand U5554 (N_5554,N_5065,N_4944);
and U5555 (N_5555,N_5157,N_5186);
xnor U5556 (N_5556,N_5223,N_4936);
or U5557 (N_5557,N_5176,N_5108);
and U5558 (N_5558,N_5393,N_5322);
or U5559 (N_5559,N_4888,N_5390);
xnor U5560 (N_5560,N_4846,N_5171);
or U5561 (N_5561,N_4904,N_5119);
and U5562 (N_5562,N_5004,N_4975);
or U5563 (N_5563,N_5330,N_5174);
and U5564 (N_5564,N_5343,N_5060);
and U5565 (N_5565,N_5278,N_4821);
or U5566 (N_5566,N_5389,N_4945);
and U5567 (N_5567,N_5387,N_5107);
or U5568 (N_5568,N_5241,N_4985);
xnor U5569 (N_5569,N_5140,N_5130);
and U5570 (N_5570,N_5295,N_5138);
nand U5571 (N_5571,N_4868,N_4823);
or U5572 (N_5572,N_4843,N_5285);
and U5573 (N_5573,N_4922,N_4994);
or U5574 (N_5574,N_4881,N_4816);
and U5575 (N_5575,N_5277,N_5064);
nor U5576 (N_5576,N_5304,N_5036);
nand U5577 (N_5577,N_5101,N_5106);
nor U5578 (N_5578,N_5260,N_4822);
or U5579 (N_5579,N_5350,N_5035);
or U5580 (N_5580,N_5129,N_4828);
xnor U5581 (N_5581,N_4976,N_5321);
nand U5582 (N_5582,N_5110,N_5325);
nand U5583 (N_5583,N_4829,N_5244);
or U5584 (N_5584,N_5173,N_5152);
or U5585 (N_5585,N_5132,N_4939);
nand U5586 (N_5586,N_5038,N_5212);
or U5587 (N_5587,N_5218,N_5216);
nor U5588 (N_5588,N_4864,N_5041);
nand U5589 (N_5589,N_5359,N_5121);
nand U5590 (N_5590,N_5061,N_5057);
xor U5591 (N_5591,N_4872,N_5292);
nor U5592 (N_5592,N_5177,N_4879);
nand U5593 (N_5593,N_4937,N_5334);
or U5594 (N_5594,N_5169,N_5009);
nand U5595 (N_5595,N_5310,N_5197);
or U5596 (N_5596,N_5317,N_4808);
or U5597 (N_5597,N_4954,N_5091);
nor U5598 (N_5598,N_5047,N_4943);
and U5599 (N_5599,N_5363,N_4924);
nor U5600 (N_5600,N_5200,N_5131);
or U5601 (N_5601,N_4929,N_5308);
or U5602 (N_5602,N_5199,N_4825);
and U5603 (N_5603,N_4921,N_4918);
nor U5604 (N_5604,N_5203,N_5011);
or U5605 (N_5605,N_5155,N_5081);
or U5606 (N_5606,N_4996,N_5221);
nor U5607 (N_5607,N_4886,N_4992);
and U5608 (N_5608,N_5015,N_4838);
nand U5609 (N_5609,N_4857,N_5112);
nand U5610 (N_5610,N_5256,N_5080);
nor U5611 (N_5611,N_5133,N_5374);
and U5612 (N_5612,N_5187,N_5297);
or U5613 (N_5613,N_5075,N_5102);
nor U5614 (N_5614,N_5147,N_5072);
nand U5615 (N_5615,N_5178,N_4933);
xnor U5616 (N_5616,N_5021,N_5283);
nand U5617 (N_5617,N_4925,N_5148);
or U5618 (N_5618,N_4972,N_4896);
and U5619 (N_5619,N_4847,N_5375);
or U5620 (N_5620,N_5324,N_4946);
nand U5621 (N_5621,N_4880,N_5115);
and U5622 (N_5622,N_5298,N_5109);
nor U5623 (N_5623,N_5205,N_5045);
nor U5624 (N_5624,N_5100,N_5090);
nand U5625 (N_5625,N_5336,N_5032);
and U5626 (N_5626,N_5344,N_5340);
nand U5627 (N_5627,N_4874,N_5236);
or U5628 (N_5628,N_4893,N_5181);
and U5629 (N_5629,N_5149,N_5306);
nor U5630 (N_5630,N_4820,N_5337);
nand U5631 (N_5631,N_4962,N_5288);
and U5632 (N_5632,N_5113,N_5145);
xor U5633 (N_5633,N_4908,N_4958);
nor U5634 (N_5634,N_4824,N_5380);
xor U5635 (N_5635,N_5092,N_4980);
or U5636 (N_5636,N_5266,N_5071);
and U5637 (N_5637,N_4827,N_5249);
nand U5638 (N_5638,N_5189,N_4942);
nor U5639 (N_5639,N_5250,N_5237);
nand U5640 (N_5640,N_5275,N_4959);
nand U5641 (N_5641,N_4841,N_5279);
or U5642 (N_5642,N_4832,N_4800);
and U5643 (N_5643,N_4873,N_5358);
and U5644 (N_5644,N_5311,N_4802);
and U5645 (N_5645,N_5209,N_5180);
nor U5646 (N_5646,N_5049,N_4999);
or U5647 (N_5647,N_4818,N_4957);
and U5648 (N_5648,N_4947,N_5124);
xor U5649 (N_5649,N_4866,N_5382);
nor U5650 (N_5650,N_4987,N_4916);
nor U5651 (N_5651,N_5030,N_5095);
and U5652 (N_5652,N_5058,N_4826);
or U5653 (N_5653,N_5215,N_5347);
and U5654 (N_5654,N_4900,N_4938);
nand U5655 (N_5655,N_5253,N_4817);
or U5656 (N_5656,N_5271,N_5034);
and U5657 (N_5657,N_4913,N_4813);
and U5658 (N_5658,N_5234,N_5153);
nand U5659 (N_5659,N_4982,N_5365);
nor U5660 (N_5660,N_4867,N_5190);
nand U5661 (N_5661,N_5276,N_4978);
xor U5662 (N_5662,N_5151,N_5220);
nor U5663 (N_5663,N_5357,N_4869);
nor U5664 (N_5664,N_5161,N_5082);
xor U5665 (N_5665,N_5096,N_5233);
xor U5666 (N_5666,N_4979,N_5208);
xnor U5667 (N_5667,N_5162,N_5335);
nand U5668 (N_5668,N_5305,N_5247);
nand U5669 (N_5669,N_5175,N_5312);
nand U5670 (N_5670,N_4977,N_5263);
and U5671 (N_5671,N_5379,N_5051);
and U5672 (N_5672,N_5055,N_5146);
nor U5673 (N_5673,N_4811,N_5341);
xnor U5674 (N_5674,N_5192,N_5001);
nand U5675 (N_5675,N_5166,N_5062);
nor U5676 (N_5676,N_4970,N_5029);
or U5677 (N_5677,N_4844,N_5012);
nor U5678 (N_5678,N_4989,N_5383);
nor U5679 (N_5679,N_5063,N_5136);
or U5680 (N_5680,N_4834,N_5143);
nand U5681 (N_5681,N_4806,N_5156);
nor U5682 (N_5682,N_5137,N_5073);
nand U5683 (N_5683,N_5031,N_5239);
nand U5684 (N_5684,N_4803,N_5248);
nor U5685 (N_5685,N_5307,N_5074);
nor U5686 (N_5686,N_5227,N_5093);
or U5687 (N_5687,N_5019,N_4836);
nand U5688 (N_5688,N_5125,N_5356);
or U5689 (N_5689,N_5327,N_5378);
or U5690 (N_5690,N_5333,N_5392);
or U5691 (N_5691,N_4910,N_5294);
nor U5692 (N_5692,N_5267,N_4964);
nor U5693 (N_5693,N_4870,N_5372);
or U5694 (N_5694,N_5395,N_5361);
nand U5695 (N_5695,N_5281,N_5089);
and U5696 (N_5696,N_5076,N_5355);
nand U5697 (N_5697,N_5053,N_5226);
nor U5698 (N_5698,N_5025,N_5371);
or U5699 (N_5699,N_4927,N_5224);
nand U5700 (N_5700,N_4985,N_4804);
and U5701 (N_5701,N_4974,N_4928);
and U5702 (N_5702,N_4946,N_5034);
or U5703 (N_5703,N_5125,N_5023);
nand U5704 (N_5704,N_5138,N_4853);
nor U5705 (N_5705,N_5281,N_5090);
nor U5706 (N_5706,N_5273,N_4857);
and U5707 (N_5707,N_5328,N_5269);
nor U5708 (N_5708,N_5182,N_5332);
nor U5709 (N_5709,N_5113,N_4868);
nand U5710 (N_5710,N_5111,N_5071);
nor U5711 (N_5711,N_4922,N_5255);
and U5712 (N_5712,N_5173,N_5096);
nand U5713 (N_5713,N_4936,N_5187);
nand U5714 (N_5714,N_4937,N_5267);
or U5715 (N_5715,N_4893,N_4831);
and U5716 (N_5716,N_5021,N_5202);
nand U5717 (N_5717,N_5263,N_5240);
nor U5718 (N_5718,N_4955,N_5274);
nor U5719 (N_5719,N_5236,N_5206);
nand U5720 (N_5720,N_4911,N_5169);
nor U5721 (N_5721,N_4807,N_5369);
nand U5722 (N_5722,N_5348,N_4991);
or U5723 (N_5723,N_4955,N_5156);
and U5724 (N_5724,N_4921,N_4914);
or U5725 (N_5725,N_4943,N_4905);
nand U5726 (N_5726,N_5096,N_4805);
xor U5727 (N_5727,N_5099,N_5340);
and U5728 (N_5728,N_5392,N_5126);
nand U5729 (N_5729,N_5066,N_5197);
and U5730 (N_5730,N_5041,N_5151);
nand U5731 (N_5731,N_5109,N_5036);
nand U5732 (N_5732,N_4971,N_5048);
nor U5733 (N_5733,N_4803,N_5366);
nand U5734 (N_5734,N_4950,N_5292);
or U5735 (N_5735,N_5093,N_5019);
or U5736 (N_5736,N_5110,N_5046);
or U5737 (N_5737,N_5031,N_5021);
nor U5738 (N_5738,N_4892,N_5120);
nand U5739 (N_5739,N_4825,N_5253);
xor U5740 (N_5740,N_5239,N_5267);
nor U5741 (N_5741,N_4815,N_5119);
and U5742 (N_5742,N_5363,N_5353);
or U5743 (N_5743,N_4810,N_5339);
or U5744 (N_5744,N_5137,N_5023);
xor U5745 (N_5745,N_5257,N_4840);
and U5746 (N_5746,N_5175,N_5044);
nor U5747 (N_5747,N_4875,N_5162);
and U5748 (N_5748,N_5354,N_4976);
or U5749 (N_5749,N_5286,N_4962);
or U5750 (N_5750,N_5041,N_5004);
nor U5751 (N_5751,N_5348,N_4982);
and U5752 (N_5752,N_5044,N_5069);
nand U5753 (N_5753,N_4806,N_5182);
nor U5754 (N_5754,N_5019,N_5320);
or U5755 (N_5755,N_5061,N_4808);
or U5756 (N_5756,N_4863,N_4913);
nor U5757 (N_5757,N_4820,N_4901);
or U5758 (N_5758,N_5078,N_5340);
nand U5759 (N_5759,N_5055,N_5354);
or U5760 (N_5760,N_5227,N_5233);
or U5761 (N_5761,N_4887,N_4897);
nand U5762 (N_5762,N_5271,N_4858);
xor U5763 (N_5763,N_4916,N_4938);
or U5764 (N_5764,N_5231,N_5384);
or U5765 (N_5765,N_5030,N_4945);
xnor U5766 (N_5766,N_4837,N_4877);
xnor U5767 (N_5767,N_5079,N_5225);
nor U5768 (N_5768,N_5291,N_5132);
xor U5769 (N_5769,N_5110,N_5271);
nand U5770 (N_5770,N_5365,N_5105);
xnor U5771 (N_5771,N_5064,N_5030);
and U5772 (N_5772,N_5094,N_5318);
and U5773 (N_5773,N_4966,N_4809);
nand U5774 (N_5774,N_4923,N_4889);
nand U5775 (N_5775,N_5383,N_5100);
and U5776 (N_5776,N_4856,N_5256);
or U5777 (N_5777,N_5074,N_5313);
and U5778 (N_5778,N_5368,N_5125);
nand U5779 (N_5779,N_5125,N_5260);
and U5780 (N_5780,N_4941,N_5011);
nand U5781 (N_5781,N_5037,N_5123);
nor U5782 (N_5782,N_4970,N_5098);
nand U5783 (N_5783,N_5390,N_5084);
nor U5784 (N_5784,N_4964,N_5241);
and U5785 (N_5785,N_5135,N_4966);
and U5786 (N_5786,N_5348,N_4862);
nand U5787 (N_5787,N_4824,N_5245);
and U5788 (N_5788,N_5393,N_4831);
or U5789 (N_5789,N_4802,N_4992);
xor U5790 (N_5790,N_5083,N_5130);
or U5791 (N_5791,N_4822,N_4886);
or U5792 (N_5792,N_5244,N_5297);
nor U5793 (N_5793,N_5393,N_4946);
nand U5794 (N_5794,N_5106,N_4978);
nand U5795 (N_5795,N_5187,N_4903);
nor U5796 (N_5796,N_4976,N_5393);
nand U5797 (N_5797,N_4805,N_5377);
nand U5798 (N_5798,N_5295,N_5240);
nand U5799 (N_5799,N_4973,N_4852);
and U5800 (N_5800,N_5189,N_4937);
nand U5801 (N_5801,N_4993,N_4907);
or U5802 (N_5802,N_5284,N_5329);
and U5803 (N_5803,N_4807,N_5316);
and U5804 (N_5804,N_5085,N_4933);
and U5805 (N_5805,N_4956,N_5337);
nor U5806 (N_5806,N_5208,N_5062);
nand U5807 (N_5807,N_5065,N_5176);
nor U5808 (N_5808,N_4809,N_5155);
nor U5809 (N_5809,N_4849,N_4880);
or U5810 (N_5810,N_5221,N_4889);
nand U5811 (N_5811,N_4963,N_4919);
or U5812 (N_5812,N_5085,N_4954);
nand U5813 (N_5813,N_4896,N_5257);
nor U5814 (N_5814,N_5370,N_5086);
or U5815 (N_5815,N_4828,N_5086);
nand U5816 (N_5816,N_4998,N_5194);
nand U5817 (N_5817,N_5300,N_5370);
nor U5818 (N_5818,N_5339,N_5008);
and U5819 (N_5819,N_4918,N_4812);
and U5820 (N_5820,N_5379,N_4843);
nand U5821 (N_5821,N_5388,N_4812);
nand U5822 (N_5822,N_5375,N_4848);
and U5823 (N_5823,N_5037,N_4878);
nand U5824 (N_5824,N_5107,N_5087);
or U5825 (N_5825,N_5063,N_4982);
or U5826 (N_5826,N_5313,N_5012);
nor U5827 (N_5827,N_5241,N_5093);
and U5828 (N_5828,N_5278,N_5314);
nand U5829 (N_5829,N_4876,N_4943);
or U5830 (N_5830,N_4903,N_5068);
and U5831 (N_5831,N_4862,N_5205);
or U5832 (N_5832,N_5186,N_5116);
nand U5833 (N_5833,N_5162,N_5216);
nor U5834 (N_5834,N_5065,N_4938);
nand U5835 (N_5835,N_4973,N_5064);
and U5836 (N_5836,N_5161,N_4897);
nor U5837 (N_5837,N_4861,N_4811);
nor U5838 (N_5838,N_5021,N_5219);
or U5839 (N_5839,N_5084,N_4867);
or U5840 (N_5840,N_5245,N_5059);
and U5841 (N_5841,N_4924,N_5282);
or U5842 (N_5842,N_5102,N_5040);
and U5843 (N_5843,N_5181,N_5003);
nor U5844 (N_5844,N_5206,N_4978);
or U5845 (N_5845,N_4879,N_5355);
nor U5846 (N_5846,N_5111,N_5031);
and U5847 (N_5847,N_4892,N_5238);
nand U5848 (N_5848,N_5310,N_5177);
or U5849 (N_5849,N_5373,N_5223);
or U5850 (N_5850,N_5053,N_5316);
nor U5851 (N_5851,N_5258,N_5155);
nand U5852 (N_5852,N_5090,N_5384);
nand U5853 (N_5853,N_4958,N_5381);
nand U5854 (N_5854,N_5251,N_5238);
nor U5855 (N_5855,N_5376,N_5363);
and U5856 (N_5856,N_5389,N_4959);
nand U5857 (N_5857,N_5134,N_5280);
nor U5858 (N_5858,N_5395,N_5357);
or U5859 (N_5859,N_4836,N_5250);
nor U5860 (N_5860,N_4890,N_5199);
and U5861 (N_5861,N_4953,N_5028);
nor U5862 (N_5862,N_5211,N_5341);
nor U5863 (N_5863,N_4809,N_5141);
and U5864 (N_5864,N_5168,N_5206);
nand U5865 (N_5865,N_4875,N_5131);
nor U5866 (N_5866,N_4863,N_5346);
xor U5867 (N_5867,N_5378,N_4881);
xor U5868 (N_5868,N_4891,N_5150);
nand U5869 (N_5869,N_5089,N_5177);
or U5870 (N_5870,N_5024,N_4897);
and U5871 (N_5871,N_4832,N_5336);
xnor U5872 (N_5872,N_5039,N_5348);
and U5873 (N_5873,N_4977,N_5172);
and U5874 (N_5874,N_5181,N_4984);
nand U5875 (N_5875,N_5195,N_5131);
xnor U5876 (N_5876,N_5224,N_5081);
nand U5877 (N_5877,N_5335,N_5233);
nor U5878 (N_5878,N_5087,N_5297);
and U5879 (N_5879,N_4834,N_5340);
nor U5880 (N_5880,N_5130,N_5248);
nand U5881 (N_5881,N_5240,N_5214);
nand U5882 (N_5882,N_5014,N_5080);
nor U5883 (N_5883,N_5075,N_5210);
and U5884 (N_5884,N_5077,N_5236);
and U5885 (N_5885,N_4849,N_5278);
nand U5886 (N_5886,N_4928,N_5240);
and U5887 (N_5887,N_5259,N_5319);
xor U5888 (N_5888,N_5142,N_5054);
or U5889 (N_5889,N_4976,N_5078);
and U5890 (N_5890,N_5146,N_5373);
and U5891 (N_5891,N_4940,N_5288);
and U5892 (N_5892,N_5304,N_5389);
nand U5893 (N_5893,N_5262,N_5235);
nand U5894 (N_5894,N_4968,N_4884);
and U5895 (N_5895,N_5378,N_5128);
nand U5896 (N_5896,N_5238,N_5165);
and U5897 (N_5897,N_5089,N_5024);
nor U5898 (N_5898,N_4924,N_5073);
nand U5899 (N_5899,N_5160,N_4876);
and U5900 (N_5900,N_5014,N_5205);
nand U5901 (N_5901,N_5309,N_5120);
nand U5902 (N_5902,N_4912,N_4830);
or U5903 (N_5903,N_4885,N_5106);
or U5904 (N_5904,N_5374,N_5165);
or U5905 (N_5905,N_4843,N_4945);
and U5906 (N_5906,N_5273,N_4932);
nand U5907 (N_5907,N_5377,N_4958);
nand U5908 (N_5908,N_5257,N_4885);
or U5909 (N_5909,N_5190,N_5003);
nand U5910 (N_5910,N_5220,N_5263);
and U5911 (N_5911,N_5117,N_5088);
nand U5912 (N_5912,N_4833,N_4886);
and U5913 (N_5913,N_5061,N_4803);
nand U5914 (N_5914,N_5143,N_5286);
nor U5915 (N_5915,N_5175,N_5088);
or U5916 (N_5916,N_5040,N_5139);
or U5917 (N_5917,N_5367,N_5111);
nand U5918 (N_5918,N_4875,N_5089);
xnor U5919 (N_5919,N_4910,N_5337);
nand U5920 (N_5920,N_4974,N_5057);
and U5921 (N_5921,N_5352,N_4966);
nand U5922 (N_5922,N_5092,N_4819);
or U5923 (N_5923,N_4931,N_5039);
nand U5924 (N_5924,N_5259,N_4957);
or U5925 (N_5925,N_4875,N_5308);
or U5926 (N_5926,N_5199,N_5239);
xnor U5927 (N_5927,N_4820,N_5149);
nor U5928 (N_5928,N_5375,N_4994);
nand U5929 (N_5929,N_4901,N_4821);
xnor U5930 (N_5930,N_5272,N_5103);
and U5931 (N_5931,N_5142,N_4861);
nand U5932 (N_5932,N_5152,N_5233);
and U5933 (N_5933,N_5336,N_5154);
or U5934 (N_5934,N_5143,N_4871);
nand U5935 (N_5935,N_5049,N_5295);
or U5936 (N_5936,N_5046,N_5100);
nand U5937 (N_5937,N_5068,N_4843);
nor U5938 (N_5938,N_5373,N_4969);
or U5939 (N_5939,N_4920,N_5311);
nand U5940 (N_5940,N_4806,N_5021);
nor U5941 (N_5941,N_5364,N_5284);
nand U5942 (N_5942,N_5114,N_5253);
nor U5943 (N_5943,N_4813,N_5385);
nand U5944 (N_5944,N_5213,N_5395);
nor U5945 (N_5945,N_5350,N_5112);
nand U5946 (N_5946,N_5082,N_5375);
nand U5947 (N_5947,N_5344,N_4813);
xor U5948 (N_5948,N_5359,N_4983);
and U5949 (N_5949,N_5037,N_5209);
nor U5950 (N_5950,N_5300,N_5279);
or U5951 (N_5951,N_4986,N_5115);
nor U5952 (N_5952,N_5119,N_5041);
and U5953 (N_5953,N_5243,N_4861);
or U5954 (N_5954,N_5198,N_4812);
nand U5955 (N_5955,N_5193,N_4858);
or U5956 (N_5956,N_5015,N_5052);
and U5957 (N_5957,N_5317,N_4998);
and U5958 (N_5958,N_4914,N_5252);
or U5959 (N_5959,N_5178,N_5329);
or U5960 (N_5960,N_4964,N_5393);
or U5961 (N_5961,N_4979,N_4876);
nand U5962 (N_5962,N_5317,N_4896);
and U5963 (N_5963,N_5086,N_5190);
or U5964 (N_5964,N_4883,N_5093);
nand U5965 (N_5965,N_5029,N_5046);
and U5966 (N_5966,N_5052,N_5019);
nor U5967 (N_5967,N_5074,N_5034);
nand U5968 (N_5968,N_5322,N_5057);
or U5969 (N_5969,N_4830,N_4897);
nand U5970 (N_5970,N_4986,N_5051);
and U5971 (N_5971,N_5084,N_5318);
nor U5972 (N_5972,N_5015,N_5150);
nand U5973 (N_5973,N_4888,N_5339);
nor U5974 (N_5974,N_5227,N_5069);
xor U5975 (N_5975,N_5202,N_5340);
nand U5976 (N_5976,N_5334,N_4852);
or U5977 (N_5977,N_5368,N_5023);
xnor U5978 (N_5978,N_5361,N_5368);
or U5979 (N_5979,N_5391,N_5160);
nor U5980 (N_5980,N_5125,N_5085);
nor U5981 (N_5981,N_4954,N_5032);
and U5982 (N_5982,N_4967,N_5156);
nor U5983 (N_5983,N_5253,N_5394);
or U5984 (N_5984,N_5009,N_5156);
or U5985 (N_5985,N_5377,N_5068);
nor U5986 (N_5986,N_5140,N_5316);
nand U5987 (N_5987,N_5060,N_5034);
and U5988 (N_5988,N_4823,N_5128);
nor U5989 (N_5989,N_5298,N_5251);
xnor U5990 (N_5990,N_5294,N_5366);
or U5991 (N_5991,N_4838,N_4963);
xnor U5992 (N_5992,N_4889,N_5280);
or U5993 (N_5993,N_4868,N_5382);
xor U5994 (N_5994,N_5215,N_5114);
nand U5995 (N_5995,N_5225,N_4867);
xnor U5996 (N_5996,N_5255,N_5302);
and U5997 (N_5997,N_4847,N_5290);
and U5998 (N_5998,N_5052,N_4804);
and U5999 (N_5999,N_4903,N_5354);
nor U6000 (N_6000,N_5741,N_5439);
nor U6001 (N_6001,N_5799,N_5459);
and U6002 (N_6002,N_5640,N_5528);
and U6003 (N_6003,N_5539,N_5667);
nand U6004 (N_6004,N_5766,N_5454);
or U6005 (N_6005,N_5639,N_5834);
nand U6006 (N_6006,N_5887,N_5982);
or U6007 (N_6007,N_5425,N_5644);
and U6008 (N_6008,N_5695,N_5960);
or U6009 (N_6009,N_5502,N_5724);
or U6010 (N_6010,N_5926,N_5818);
xnor U6011 (N_6011,N_5694,N_5624);
or U6012 (N_6012,N_5816,N_5487);
nor U6013 (N_6013,N_5819,N_5933);
and U6014 (N_6014,N_5708,N_5714);
or U6015 (N_6015,N_5430,N_5850);
nand U6016 (N_6016,N_5420,N_5770);
nor U6017 (N_6017,N_5451,N_5655);
nand U6018 (N_6018,N_5715,N_5980);
or U6019 (N_6019,N_5495,N_5917);
or U6020 (N_6020,N_5434,N_5597);
or U6021 (N_6021,N_5526,N_5919);
or U6022 (N_6022,N_5757,N_5410);
or U6023 (N_6023,N_5930,N_5900);
nor U6024 (N_6024,N_5879,N_5599);
or U6025 (N_6025,N_5742,N_5636);
nor U6026 (N_6026,N_5939,N_5907);
and U6027 (N_6027,N_5428,N_5914);
and U6028 (N_6028,N_5978,N_5493);
nand U6029 (N_6029,N_5970,N_5929);
and U6030 (N_6030,N_5865,N_5952);
nand U6031 (N_6031,N_5586,N_5617);
or U6032 (N_6032,N_5522,N_5480);
nor U6033 (N_6033,N_5922,N_5553);
and U6034 (N_6034,N_5792,N_5534);
nand U6035 (N_6035,N_5643,N_5657);
or U6036 (N_6036,N_5411,N_5795);
and U6037 (N_6037,N_5844,N_5921);
or U6038 (N_6038,N_5728,N_5533);
or U6039 (N_6039,N_5682,N_5969);
nand U6040 (N_6040,N_5404,N_5532);
or U6041 (N_6041,N_5462,N_5491);
nand U6042 (N_6042,N_5431,N_5693);
nor U6043 (N_6043,N_5854,N_5940);
nor U6044 (N_6044,N_5691,N_5606);
xnor U6045 (N_6045,N_5689,N_5713);
nor U6046 (N_6046,N_5443,N_5506);
nor U6047 (N_6047,N_5497,N_5448);
xnor U6048 (N_6048,N_5492,N_5779);
and U6049 (N_6049,N_5456,N_5958);
nor U6050 (N_6050,N_5482,N_5630);
or U6051 (N_6051,N_5635,N_5992);
nor U6052 (N_6052,N_5609,N_5772);
and U6053 (N_6053,N_5419,N_5886);
or U6054 (N_6054,N_5582,N_5610);
or U6055 (N_6055,N_5863,N_5836);
or U6056 (N_6056,N_5878,N_5883);
nand U6057 (N_6057,N_5452,N_5584);
nand U6058 (N_6058,N_5938,N_5481);
and U6059 (N_6059,N_5463,N_5648);
nor U6060 (N_6060,N_5437,N_5829);
and U6061 (N_6061,N_5801,N_5412);
and U6062 (N_6062,N_5902,N_5875);
and U6063 (N_6063,N_5512,N_5458);
nand U6064 (N_6064,N_5857,N_5824);
or U6065 (N_6065,N_5979,N_5785);
xnor U6066 (N_6066,N_5619,N_5561);
xor U6067 (N_6067,N_5468,N_5686);
nand U6068 (N_6068,N_5861,N_5413);
nand U6069 (N_6069,N_5796,N_5471);
nand U6070 (N_6070,N_5569,N_5706);
and U6071 (N_6071,N_5611,N_5676);
nand U6072 (N_6072,N_5455,N_5935);
nand U6073 (N_6073,N_5725,N_5681);
or U6074 (N_6074,N_5628,N_5418);
nor U6075 (N_6075,N_5759,N_5967);
xor U6076 (N_6076,N_5986,N_5794);
nand U6077 (N_6077,N_5479,N_5751);
nor U6078 (N_6078,N_5531,N_5745);
or U6079 (N_6079,N_5538,N_5906);
nand U6080 (N_6080,N_5548,N_5555);
or U6081 (N_6081,N_5874,N_5777);
and U6082 (N_6082,N_5415,N_5670);
nand U6083 (N_6083,N_5580,N_5445);
nor U6084 (N_6084,N_5600,N_5896);
and U6085 (N_6085,N_5566,N_5918);
nor U6086 (N_6086,N_5767,N_5950);
nand U6087 (N_6087,N_5966,N_5634);
nor U6088 (N_6088,N_5870,N_5525);
nand U6089 (N_6089,N_5898,N_5756);
nor U6090 (N_6090,N_5607,N_5405);
and U6091 (N_6091,N_5421,N_5833);
xnor U6092 (N_6092,N_5780,N_5401);
and U6093 (N_6093,N_5513,N_5965);
or U6094 (N_6094,N_5760,N_5859);
or U6095 (N_6095,N_5438,N_5707);
nand U6096 (N_6096,N_5956,N_5484);
and U6097 (N_6097,N_5647,N_5574);
nor U6098 (N_6098,N_5696,N_5743);
nor U6099 (N_6099,N_5800,N_5503);
xnor U6100 (N_6100,N_5858,N_5633);
or U6101 (N_6101,N_5558,N_5564);
nand U6102 (N_6102,N_5505,N_5987);
or U6103 (N_6103,N_5831,N_5755);
and U6104 (N_6104,N_5614,N_5973);
nor U6105 (N_6105,N_5699,N_5809);
and U6106 (N_6106,N_5923,N_5447);
or U6107 (N_6107,N_5783,N_5465);
and U6108 (N_6108,N_5507,N_5807);
nand U6109 (N_6109,N_5662,N_5910);
nand U6110 (N_6110,N_5478,N_5596);
nand U6111 (N_6111,N_5669,N_5746);
and U6112 (N_6112,N_5901,N_5571);
nor U6113 (N_6113,N_5666,N_5868);
or U6114 (N_6114,N_5748,N_5882);
and U6115 (N_6115,N_5984,N_5905);
xnor U6116 (N_6116,N_5663,N_5638);
nor U6117 (N_6117,N_5664,N_5668);
nor U6118 (N_6118,N_5717,N_5727);
and U6119 (N_6119,N_5521,N_5999);
nand U6120 (N_6120,N_5880,N_5426);
and U6121 (N_6121,N_5559,N_5991);
or U6122 (N_6122,N_5649,N_5613);
and U6123 (N_6123,N_5530,N_5576);
or U6124 (N_6124,N_5869,N_5841);
or U6125 (N_6125,N_5685,N_5890);
or U6126 (N_6126,N_5744,N_5738);
or U6127 (N_6127,N_5400,N_5941);
or U6128 (N_6128,N_5535,N_5828);
nor U6129 (N_6129,N_5771,N_5729);
and U6130 (N_6130,N_5955,N_5943);
or U6131 (N_6131,N_5848,N_5466);
nand U6132 (N_6132,N_5932,N_5954);
or U6133 (N_6133,N_5802,N_5704);
nand U6134 (N_6134,N_5786,N_5435);
nor U6135 (N_6135,N_5523,N_5622);
nor U6136 (N_6136,N_5632,N_5872);
nor U6137 (N_6137,N_5436,N_5823);
nand U6138 (N_6138,N_5461,N_5812);
and U6139 (N_6139,N_5990,N_5838);
and U6140 (N_6140,N_5563,N_5787);
and U6141 (N_6141,N_5881,N_5911);
nor U6142 (N_6142,N_5519,N_5803);
nand U6143 (N_6143,N_5862,N_5402);
nor U6144 (N_6144,N_5683,N_5804);
or U6145 (N_6145,N_5453,N_5722);
and U6146 (N_6146,N_5849,N_5782);
or U6147 (N_6147,N_5605,N_5567);
or U6148 (N_6148,N_5414,N_5602);
and U6149 (N_6149,N_5843,N_5557);
or U6150 (N_6150,N_5540,N_5733);
nor U6151 (N_6151,N_5578,N_5659);
or U6152 (N_6152,N_5688,N_5572);
nor U6153 (N_6153,N_5594,N_5876);
or U6154 (N_6154,N_5855,N_5520);
and U6155 (N_6155,N_5856,N_5731);
and U6156 (N_6156,N_5474,N_5514);
nand U6157 (N_6157,N_5629,N_5705);
and U6158 (N_6158,N_5529,N_5835);
nand U6159 (N_6159,N_5516,N_5702);
nand U6160 (N_6160,N_5994,N_5981);
nand U6161 (N_6161,N_5551,N_5601);
or U6162 (N_6162,N_5737,N_5568);
or U6163 (N_6163,N_5603,N_5920);
and U6164 (N_6164,N_5996,N_5826);
and U6165 (N_6165,N_5498,N_5719);
and U6166 (N_6166,N_5937,N_5690);
nand U6167 (N_6167,N_5953,N_5560);
nor U6168 (N_6168,N_5821,N_5692);
or U6169 (N_6169,N_5813,N_5549);
and U6170 (N_6170,N_5995,N_5416);
nand U6171 (N_6171,N_5997,N_5673);
nor U6172 (N_6172,N_5577,N_5515);
xor U6173 (N_6173,N_5552,N_5974);
nor U6174 (N_6174,N_5944,N_5444);
xor U6175 (N_6175,N_5583,N_5457);
or U6176 (N_6176,N_5543,N_5889);
nand U6177 (N_6177,N_5680,N_5671);
or U6178 (N_6178,N_5562,N_5740);
and U6179 (N_6179,N_5556,N_5499);
nand U6180 (N_6180,N_5627,N_5830);
nor U6181 (N_6181,N_5721,N_5590);
xnor U6182 (N_6182,N_5961,N_5775);
nor U6183 (N_6183,N_5591,N_5726);
xor U6184 (N_6184,N_5537,N_5672);
nand U6185 (N_6185,N_5888,N_5720);
nor U6186 (N_6186,N_5711,N_5931);
xor U6187 (N_6187,N_5485,N_5971);
nor U6188 (N_6188,N_5623,N_5650);
xnor U6189 (N_6189,N_5422,N_5579);
nor U6190 (N_6190,N_5432,N_5697);
nor U6191 (N_6191,N_5749,N_5504);
nor U6192 (N_6192,N_5957,N_5765);
or U6193 (N_6193,N_5710,N_5545);
nor U6194 (N_6194,N_5845,N_5735);
xor U6195 (N_6195,N_5864,N_5524);
xor U6196 (N_6196,N_5962,N_5544);
xor U6197 (N_6197,N_5409,N_5616);
and U6198 (N_6198,N_5550,N_5764);
and U6199 (N_6199,N_5989,N_5976);
xnor U6200 (N_6200,N_5885,N_5518);
or U6201 (N_6201,N_5656,N_5654);
nand U6202 (N_6202,N_5762,N_5815);
and U6203 (N_6203,N_5595,N_5983);
or U6204 (N_6204,N_5449,N_5429);
nor U6205 (N_6205,N_5675,N_5761);
and U6206 (N_6206,N_5768,N_5934);
nand U6207 (N_6207,N_5773,N_5440);
nor U6208 (N_6208,N_5945,N_5651);
nand U6209 (N_6209,N_5985,N_5565);
or U6210 (N_6210,N_5475,N_5959);
nand U6211 (N_6211,N_5892,N_5575);
nand U6212 (N_6212,N_5684,N_5894);
or U6213 (N_6213,N_5631,N_5968);
and U6214 (N_6214,N_5408,N_5608);
nor U6215 (N_6215,N_5903,N_5687);
xnor U6216 (N_6216,N_5433,N_5645);
nand U6217 (N_6217,N_5470,N_5665);
and U6218 (N_6218,N_5946,N_5641);
and U6219 (N_6219,N_5781,N_5486);
and U6220 (N_6220,N_5621,N_5758);
xnor U6221 (N_6221,N_5866,N_5827);
nand U6222 (N_6222,N_5788,N_5403);
and U6223 (N_6223,N_5924,N_5723);
or U6224 (N_6224,N_5912,N_5424);
and U6225 (N_6225,N_5913,N_5776);
nor U6226 (N_6226,N_5677,N_5963);
or U6227 (N_6227,N_5734,N_5851);
or U6228 (N_6228,N_5884,N_5975);
nor U6229 (N_6229,N_5747,N_5825);
xor U6230 (N_6230,N_5700,N_5712);
and U6231 (N_6231,N_5846,N_5951);
and U6232 (N_6232,N_5769,N_5679);
nand U6233 (N_6233,N_5774,N_5853);
or U6234 (N_6234,N_5791,N_5536);
or U6235 (N_6235,N_5573,N_5817);
and U6236 (N_6236,N_5936,N_5646);
nand U6237 (N_6237,N_5446,N_5585);
nor U6238 (N_6238,N_5904,N_5542);
or U6239 (N_6239,N_5750,N_5972);
nor U6240 (N_6240,N_5661,N_5441);
or U6241 (N_6241,N_5652,N_5797);
nand U6242 (N_6242,N_5778,N_5810);
xnor U6243 (N_6243,N_5483,N_5867);
nor U6244 (N_6244,N_5832,N_5500);
and U6245 (N_6245,N_5620,N_5909);
nor U6246 (N_6246,N_5509,N_5942);
xnor U6247 (N_6247,N_5899,N_5626);
nor U6248 (N_6248,N_5489,N_5427);
and U6249 (N_6249,N_5472,N_5837);
nand U6250 (N_6250,N_5998,N_5763);
xnor U6251 (N_6251,N_5798,N_5510);
xnor U6252 (N_6252,N_5842,N_5698);
or U6253 (N_6253,N_5467,N_5893);
and U6254 (N_6254,N_5977,N_5406);
or U6255 (N_6255,N_5716,N_5925);
nor U6256 (N_6256,N_5877,N_5895);
nor U6257 (N_6257,N_5653,N_5752);
or U6258 (N_6258,N_5570,N_5789);
xor U6259 (N_6259,N_5811,N_5820);
or U6260 (N_6260,N_5642,N_5790);
and U6261 (N_6261,N_5547,N_5784);
or U6262 (N_6262,N_5598,N_5477);
xor U6263 (N_6263,N_5476,N_5541);
and U6264 (N_6264,N_5581,N_5674);
or U6265 (N_6265,N_5587,N_5840);
nor U6266 (N_6266,N_5891,N_5948);
or U6267 (N_6267,N_5871,N_5964);
nand U6268 (N_6268,N_5847,N_5860);
and U6269 (N_6269,N_5407,N_5808);
or U6270 (N_6270,N_5908,N_5464);
or U6271 (N_6271,N_5927,N_5916);
and U6272 (N_6272,N_5417,N_5709);
nor U6273 (N_6273,N_5928,N_5814);
nor U6274 (N_6274,N_5469,N_5496);
or U6275 (N_6275,N_5718,N_5615);
nor U6276 (N_6276,N_5915,N_5511);
and U6277 (N_6277,N_5739,N_5546);
or U6278 (N_6278,N_5703,N_5460);
nand U6279 (N_6279,N_5442,N_5618);
or U6280 (N_6280,N_5527,N_5873);
or U6281 (N_6281,N_5949,N_5423);
nand U6282 (N_6282,N_5754,N_5517);
nand U6283 (N_6283,N_5473,N_5637);
and U6284 (N_6284,N_5490,N_5494);
nand U6285 (N_6285,N_5658,N_5839);
nand U6286 (N_6286,N_5501,N_5604);
xor U6287 (N_6287,N_5593,N_5588);
and U6288 (N_6288,N_5736,N_5450);
xor U6289 (N_6289,N_5852,N_5701);
nand U6290 (N_6290,N_5805,N_5732);
or U6291 (N_6291,N_5897,N_5488);
or U6292 (N_6292,N_5592,N_5678);
nor U6293 (N_6293,N_5612,N_5554);
and U6294 (N_6294,N_5660,N_5508);
or U6295 (N_6295,N_5988,N_5625);
xor U6296 (N_6296,N_5753,N_5730);
nand U6297 (N_6297,N_5947,N_5806);
nor U6298 (N_6298,N_5993,N_5589);
and U6299 (N_6299,N_5793,N_5822);
and U6300 (N_6300,N_5424,N_5724);
and U6301 (N_6301,N_5740,N_5879);
nand U6302 (N_6302,N_5603,N_5635);
nor U6303 (N_6303,N_5641,N_5677);
nand U6304 (N_6304,N_5771,N_5734);
and U6305 (N_6305,N_5831,N_5689);
nor U6306 (N_6306,N_5444,N_5581);
nand U6307 (N_6307,N_5484,N_5658);
or U6308 (N_6308,N_5785,N_5980);
nand U6309 (N_6309,N_5765,N_5623);
nand U6310 (N_6310,N_5545,N_5681);
and U6311 (N_6311,N_5880,N_5563);
or U6312 (N_6312,N_5631,N_5420);
or U6313 (N_6313,N_5811,N_5793);
or U6314 (N_6314,N_5475,N_5768);
and U6315 (N_6315,N_5678,N_5996);
nand U6316 (N_6316,N_5543,N_5884);
xor U6317 (N_6317,N_5815,N_5574);
and U6318 (N_6318,N_5876,N_5794);
or U6319 (N_6319,N_5578,N_5896);
nand U6320 (N_6320,N_5770,N_5947);
or U6321 (N_6321,N_5470,N_5709);
nand U6322 (N_6322,N_5554,N_5947);
nor U6323 (N_6323,N_5760,N_5640);
nor U6324 (N_6324,N_5563,N_5641);
xor U6325 (N_6325,N_5441,N_5420);
nand U6326 (N_6326,N_5480,N_5959);
xnor U6327 (N_6327,N_5591,N_5494);
or U6328 (N_6328,N_5564,N_5968);
or U6329 (N_6329,N_5873,N_5569);
and U6330 (N_6330,N_5623,N_5422);
or U6331 (N_6331,N_5901,N_5818);
and U6332 (N_6332,N_5739,N_5755);
and U6333 (N_6333,N_5864,N_5514);
nor U6334 (N_6334,N_5610,N_5652);
xor U6335 (N_6335,N_5516,N_5499);
xnor U6336 (N_6336,N_5919,N_5915);
nand U6337 (N_6337,N_5706,N_5890);
nand U6338 (N_6338,N_5600,N_5665);
and U6339 (N_6339,N_5827,N_5815);
or U6340 (N_6340,N_5589,N_5417);
xor U6341 (N_6341,N_5466,N_5518);
nand U6342 (N_6342,N_5823,N_5594);
xor U6343 (N_6343,N_5843,N_5809);
or U6344 (N_6344,N_5464,N_5694);
or U6345 (N_6345,N_5955,N_5835);
nand U6346 (N_6346,N_5969,N_5561);
nand U6347 (N_6347,N_5981,N_5879);
and U6348 (N_6348,N_5526,N_5941);
or U6349 (N_6349,N_5771,N_5479);
nor U6350 (N_6350,N_5732,N_5657);
nor U6351 (N_6351,N_5585,N_5928);
and U6352 (N_6352,N_5792,N_5907);
or U6353 (N_6353,N_5553,N_5589);
nor U6354 (N_6354,N_5677,N_5753);
nand U6355 (N_6355,N_5514,N_5579);
and U6356 (N_6356,N_5778,N_5831);
or U6357 (N_6357,N_5437,N_5606);
or U6358 (N_6358,N_5427,N_5473);
or U6359 (N_6359,N_5532,N_5772);
or U6360 (N_6360,N_5610,N_5498);
nor U6361 (N_6361,N_5424,N_5703);
or U6362 (N_6362,N_5602,N_5942);
nand U6363 (N_6363,N_5504,N_5617);
nor U6364 (N_6364,N_5638,N_5779);
or U6365 (N_6365,N_5449,N_5481);
xnor U6366 (N_6366,N_5471,N_5821);
nor U6367 (N_6367,N_5927,N_5789);
nor U6368 (N_6368,N_5454,N_5958);
nor U6369 (N_6369,N_5601,N_5620);
nand U6370 (N_6370,N_5765,N_5510);
and U6371 (N_6371,N_5694,N_5475);
xor U6372 (N_6372,N_5677,N_5816);
and U6373 (N_6373,N_5654,N_5800);
nor U6374 (N_6374,N_5541,N_5816);
and U6375 (N_6375,N_5603,N_5935);
or U6376 (N_6376,N_5474,N_5743);
and U6377 (N_6377,N_5943,N_5760);
nor U6378 (N_6378,N_5422,N_5768);
nor U6379 (N_6379,N_5457,N_5948);
or U6380 (N_6380,N_5859,N_5695);
or U6381 (N_6381,N_5710,N_5857);
and U6382 (N_6382,N_5657,N_5670);
nor U6383 (N_6383,N_5542,N_5441);
nand U6384 (N_6384,N_5750,N_5986);
and U6385 (N_6385,N_5775,N_5855);
and U6386 (N_6386,N_5904,N_5660);
and U6387 (N_6387,N_5703,N_5998);
and U6388 (N_6388,N_5432,N_5895);
nand U6389 (N_6389,N_5490,N_5471);
or U6390 (N_6390,N_5442,N_5537);
and U6391 (N_6391,N_5740,N_5631);
nand U6392 (N_6392,N_5852,N_5760);
nor U6393 (N_6393,N_5436,N_5488);
nand U6394 (N_6394,N_5834,N_5439);
and U6395 (N_6395,N_5469,N_5733);
xnor U6396 (N_6396,N_5687,N_5583);
and U6397 (N_6397,N_5469,N_5799);
or U6398 (N_6398,N_5945,N_5545);
xor U6399 (N_6399,N_5587,N_5819);
nand U6400 (N_6400,N_5865,N_5862);
or U6401 (N_6401,N_5687,N_5810);
nor U6402 (N_6402,N_5447,N_5688);
nor U6403 (N_6403,N_5818,N_5987);
and U6404 (N_6404,N_5501,N_5993);
nor U6405 (N_6405,N_5881,N_5698);
nand U6406 (N_6406,N_5762,N_5899);
nor U6407 (N_6407,N_5617,N_5772);
or U6408 (N_6408,N_5818,N_5563);
and U6409 (N_6409,N_5908,N_5466);
and U6410 (N_6410,N_5905,N_5711);
or U6411 (N_6411,N_5568,N_5632);
nand U6412 (N_6412,N_5736,N_5489);
and U6413 (N_6413,N_5899,N_5720);
or U6414 (N_6414,N_5908,N_5884);
and U6415 (N_6415,N_5816,N_5485);
or U6416 (N_6416,N_5459,N_5829);
nor U6417 (N_6417,N_5817,N_5783);
or U6418 (N_6418,N_5504,N_5912);
and U6419 (N_6419,N_5509,N_5534);
and U6420 (N_6420,N_5551,N_5750);
nor U6421 (N_6421,N_5692,N_5452);
or U6422 (N_6422,N_5857,N_5908);
nor U6423 (N_6423,N_5751,N_5968);
and U6424 (N_6424,N_5408,N_5816);
nand U6425 (N_6425,N_5656,N_5925);
xor U6426 (N_6426,N_5960,N_5955);
or U6427 (N_6427,N_5909,N_5835);
xor U6428 (N_6428,N_5490,N_5597);
and U6429 (N_6429,N_5977,N_5871);
or U6430 (N_6430,N_5609,N_5827);
and U6431 (N_6431,N_5893,N_5784);
and U6432 (N_6432,N_5423,N_5881);
or U6433 (N_6433,N_5569,N_5639);
and U6434 (N_6434,N_5539,N_5754);
nand U6435 (N_6435,N_5952,N_5840);
or U6436 (N_6436,N_5584,N_5987);
nor U6437 (N_6437,N_5919,N_5707);
nor U6438 (N_6438,N_5860,N_5653);
or U6439 (N_6439,N_5723,N_5973);
and U6440 (N_6440,N_5686,N_5672);
and U6441 (N_6441,N_5959,N_5776);
nand U6442 (N_6442,N_5861,N_5649);
nand U6443 (N_6443,N_5723,N_5677);
and U6444 (N_6444,N_5738,N_5581);
xor U6445 (N_6445,N_5656,N_5845);
and U6446 (N_6446,N_5789,N_5854);
nor U6447 (N_6447,N_5701,N_5833);
nand U6448 (N_6448,N_5628,N_5585);
or U6449 (N_6449,N_5941,N_5741);
nor U6450 (N_6450,N_5673,N_5710);
nand U6451 (N_6451,N_5636,N_5479);
nor U6452 (N_6452,N_5675,N_5527);
nand U6453 (N_6453,N_5534,N_5500);
and U6454 (N_6454,N_5620,N_5404);
and U6455 (N_6455,N_5666,N_5450);
or U6456 (N_6456,N_5809,N_5979);
and U6457 (N_6457,N_5937,N_5637);
or U6458 (N_6458,N_5978,N_5692);
or U6459 (N_6459,N_5814,N_5727);
and U6460 (N_6460,N_5543,N_5759);
nand U6461 (N_6461,N_5840,N_5697);
xnor U6462 (N_6462,N_5899,N_5832);
nor U6463 (N_6463,N_5491,N_5549);
and U6464 (N_6464,N_5797,N_5491);
xor U6465 (N_6465,N_5627,N_5999);
or U6466 (N_6466,N_5587,N_5589);
nor U6467 (N_6467,N_5764,N_5645);
and U6468 (N_6468,N_5759,N_5748);
and U6469 (N_6469,N_5430,N_5509);
nor U6470 (N_6470,N_5920,N_5545);
and U6471 (N_6471,N_5946,N_5823);
xnor U6472 (N_6472,N_5646,N_5640);
or U6473 (N_6473,N_5777,N_5618);
nand U6474 (N_6474,N_5906,N_5619);
and U6475 (N_6475,N_5804,N_5563);
or U6476 (N_6476,N_5426,N_5959);
nand U6477 (N_6477,N_5747,N_5464);
nor U6478 (N_6478,N_5459,N_5831);
and U6479 (N_6479,N_5830,N_5897);
nor U6480 (N_6480,N_5429,N_5948);
nor U6481 (N_6481,N_5588,N_5750);
and U6482 (N_6482,N_5927,N_5872);
or U6483 (N_6483,N_5697,N_5444);
and U6484 (N_6484,N_5485,N_5490);
nor U6485 (N_6485,N_5419,N_5459);
or U6486 (N_6486,N_5916,N_5871);
nor U6487 (N_6487,N_5587,N_5961);
or U6488 (N_6488,N_5581,N_5484);
nor U6489 (N_6489,N_5921,N_5753);
nor U6490 (N_6490,N_5626,N_5467);
nor U6491 (N_6491,N_5996,N_5745);
nor U6492 (N_6492,N_5632,N_5753);
xnor U6493 (N_6493,N_5624,N_5833);
and U6494 (N_6494,N_5816,N_5516);
nor U6495 (N_6495,N_5960,N_5582);
nand U6496 (N_6496,N_5767,N_5989);
nand U6497 (N_6497,N_5846,N_5629);
nor U6498 (N_6498,N_5873,N_5516);
nand U6499 (N_6499,N_5539,N_5448);
or U6500 (N_6500,N_5572,N_5650);
and U6501 (N_6501,N_5618,N_5778);
nor U6502 (N_6502,N_5614,N_5452);
nand U6503 (N_6503,N_5724,N_5553);
and U6504 (N_6504,N_5953,N_5686);
and U6505 (N_6505,N_5682,N_5815);
nand U6506 (N_6506,N_5655,N_5827);
or U6507 (N_6507,N_5711,N_5679);
and U6508 (N_6508,N_5980,N_5612);
or U6509 (N_6509,N_5794,N_5957);
nand U6510 (N_6510,N_5410,N_5731);
and U6511 (N_6511,N_5871,N_5863);
or U6512 (N_6512,N_5627,N_5930);
nor U6513 (N_6513,N_5496,N_5688);
xnor U6514 (N_6514,N_5431,N_5675);
xor U6515 (N_6515,N_5972,N_5626);
and U6516 (N_6516,N_5781,N_5849);
xor U6517 (N_6517,N_5605,N_5956);
nor U6518 (N_6518,N_5508,N_5980);
nor U6519 (N_6519,N_5436,N_5579);
or U6520 (N_6520,N_5845,N_5641);
and U6521 (N_6521,N_5420,N_5751);
nor U6522 (N_6522,N_5559,N_5656);
nor U6523 (N_6523,N_5669,N_5900);
nand U6524 (N_6524,N_5631,N_5618);
nand U6525 (N_6525,N_5401,N_5931);
and U6526 (N_6526,N_5532,N_5587);
or U6527 (N_6527,N_5911,N_5402);
or U6528 (N_6528,N_5613,N_5863);
or U6529 (N_6529,N_5997,N_5623);
xor U6530 (N_6530,N_5533,N_5497);
or U6531 (N_6531,N_5585,N_5425);
or U6532 (N_6532,N_5507,N_5810);
nand U6533 (N_6533,N_5840,N_5544);
and U6534 (N_6534,N_5841,N_5653);
nor U6535 (N_6535,N_5766,N_5938);
nand U6536 (N_6536,N_5801,N_5567);
and U6537 (N_6537,N_5595,N_5474);
nor U6538 (N_6538,N_5530,N_5735);
or U6539 (N_6539,N_5722,N_5832);
nor U6540 (N_6540,N_5918,N_5883);
or U6541 (N_6541,N_5836,N_5967);
xor U6542 (N_6542,N_5606,N_5674);
nand U6543 (N_6543,N_5580,N_5591);
and U6544 (N_6544,N_5788,N_5644);
nand U6545 (N_6545,N_5888,N_5932);
or U6546 (N_6546,N_5879,N_5935);
and U6547 (N_6547,N_5504,N_5466);
nand U6548 (N_6548,N_5713,N_5887);
and U6549 (N_6549,N_5572,N_5566);
nor U6550 (N_6550,N_5540,N_5652);
or U6551 (N_6551,N_5442,N_5433);
and U6552 (N_6552,N_5882,N_5989);
or U6553 (N_6553,N_5741,N_5695);
or U6554 (N_6554,N_5608,N_5422);
nand U6555 (N_6555,N_5996,N_5434);
and U6556 (N_6556,N_5753,N_5797);
nand U6557 (N_6557,N_5655,N_5600);
or U6558 (N_6558,N_5971,N_5880);
nor U6559 (N_6559,N_5717,N_5564);
and U6560 (N_6560,N_5606,N_5901);
and U6561 (N_6561,N_5709,N_5477);
nand U6562 (N_6562,N_5575,N_5435);
nor U6563 (N_6563,N_5729,N_5597);
nor U6564 (N_6564,N_5457,N_5951);
and U6565 (N_6565,N_5752,N_5903);
and U6566 (N_6566,N_5966,N_5856);
nor U6567 (N_6567,N_5741,N_5707);
xnor U6568 (N_6568,N_5968,N_5406);
or U6569 (N_6569,N_5406,N_5607);
or U6570 (N_6570,N_5682,N_5939);
nand U6571 (N_6571,N_5615,N_5645);
nand U6572 (N_6572,N_5630,N_5831);
and U6573 (N_6573,N_5769,N_5905);
nor U6574 (N_6574,N_5963,N_5901);
xnor U6575 (N_6575,N_5757,N_5439);
nand U6576 (N_6576,N_5800,N_5455);
nor U6577 (N_6577,N_5960,N_5836);
nor U6578 (N_6578,N_5553,N_5544);
nor U6579 (N_6579,N_5434,N_5888);
xnor U6580 (N_6580,N_5550,N_5400);
and U6581 (N_6581,N_5712,N_5711);
or U6582 (N_6582,N_5441,N_5446);
or U6583 (N_6583,N_5653,N_5437);
xor U6584 (N_6584,N_5461,N_5479);
nor U6585 (N_6585,N_5755,N_5445);
and U6586 (N_6586,N_5405,N_5613);
nor U6587 (N_6587,N_5875,N_5440);
nor U6588 (N_6588,N_5527,N_5662);
nand U6589 (N_6589,N_5663,N_5954);
nor U6590 (N_6590,N_5482,N_5529);
and U6591 (N_6591,N_5415,N_5796);
nand U6592 (N_6592,N_5839,N_5481);
and U6593 (N_6593,N_5930,N_5664);
xnor U6594 (N_6594,N_5911,N_5937);
nand U6595 (N_6595,N_5666,N_5408);
xnor U6596 (N_6596,N_5606,N_5621);
nor U6597 (N_6597,N_5491,N_5701);
or U6598 (N_6598,N_5799,N_5893);
nor U6599 (N_6599,N_5896,N_5497);
and U6600 (N_6600,N_6128,N_6533);
nand U6601 (N_6601,N_6268,N_6366);
nand U6602 (N_6602,N_6059,N_6566);
xor U6603 (N_6603,N_6389,N_6392);
and U6604 (N_6604,N_6290,N_6069);
nand U6605 (N_6605,N_6125,N_6191);
xor U6606 (N_6606,N_6467,N_6134);
or U6607 (N_6607,N_6365,N_6204);
or U6608 (N_6608,N_6063,N_6508);
nand U6609 (N_6609,N_6504,N_6295);
nor U6610 (N_6610,N_6198,N_6108);
and U6611 (N_6611,N_6588,N_6439);
and U6612 (N_6612,N_6495,N_6018);
or U6613 (N_6613,N_6115,N_6010);
and U6614 (N_6614,N_6407,N_6346);
nor U6615 (N_6615,N_6254,N_6236);
and U6616 (N_6616,N_6492,N_6273);
and U6617 (N_6617,N_6395,N_6189);
or U6618 (N_6618,N_6517,N_6086);
nand U6619 (N_6619,N_6054,N_6292);
xor U6620 (N_6620,N_6576,N_6451);
or U6621 (N_6621,N_6462,N_6070);
or U6622 (N_6622,N_6399,N_6187);
or U6623 (N_6623,N_6129,N_6412);
nor U6624 (N_6624,N_6406,N_6307);
nor U6625 (N_6625,N_6363,N_6415);
xor U6626 (N_6626,N_6526,N_6170);
nor U6627 (N_6627,N_6417,N_6248);
nand U6628 (N_6628,N_6348,N_6320);
or U6629 (N_6629,N_6057,N_6403);
and U6630 (N_6630,N_6499,N_6515);
nor U6631 (N_6631,N_6209,N_6075);
nor U6632 (N_6632,N_6120,N_6459);
and U6633 (N_6633,N_6240,N_6146);
and U6634 (N_6634,N_6163,N_6225);
nand U6635 (N_6635,N_6545,N_6454);
or U6636 (N_6636,N_6599,N_6507);
or U6637 (N_6637,N_6152,N_6024);
xnor U6638 (N_6638,N_6523,N_6211);
or U6639 (N_6639,N_6172,N_6481);
xor U6640 (N_6640,N_6141,N_6221);
nand U6641 (N_6641,N_6458,N_6592);
and U6642 (N_6642,N_6285,N_6232);
or U6643 (N_6643,N_6247,N_6029);
or U6644 (N_6644,N_6148,N_6357);
and U6645 (N_6645,N_6019,N_6347);
or U6646 (N_6646,N_6231,N_6354);
nand U6647 (N_6647,N_6216,N_6340);
or U6648 (N_6648,N_6337,N_6375);
and U6649 (N_6649,N_6503,N_6561);
nand U6650 (N_6650,N_6360,N_6534);
nor U6651 (N_6651,N_6323,N_6502);
and U6652 (N_6652,N_6262,N_6362);
nor U6653 (N_6653,N_6193,N_6324);
nand U6654 (N_6654,N_6235,N_6530);
and U6655 (N_6655,N_6156,N_6149);
xnor U6656 (N_6656,N_6031,N_6571);
nor U6657 (N_6657,N_6028,N_6103);
or U6658 (N_6658,N_6111,N_6581);
and U6659 (N_6659,N_6005,N_6264);
nand U6660 (N_6660,N_6334,N_6289);
nor U6661 (N_6661,N_6328,N_6388);
nand U6662 (N_6662,N_6577,N_6420);
and U6663 (N_6663,N_6026,N_6107);
or U6664 (N_6664,N_6164,N_6242);
nand U6665 (N_6665,N_6368,N_6060);
and U6666 (N_6666,N_6066,N_6300);
nand U6667 (N_6667,N_6319,N_6233);
nor U6668 (N_6668,N_6280,N_6376);
nand U6669 (N_6669,N_6331,N_6297);
nand U6670 (N_6670,N_6404,N_6578);
and U6671 (N_6671,N_6091,N_6188);
and U6672 (N_6672,N_6222,N_6513);
nor U6673 (N_6673,N_6284,N_6055);
nor U6674 (N_6674,N_6461,N_6097);
xnor U6675 (N_6675,N_6483,N_6243);
or U6676 (N_6676,N_6138,N_6531);
nand U6677 (N_6677,N_6291,N_6118);
xnor U6678 (N_6678,N_6261,N_6355);
nor U6679 (N_6679,N_6474,N_6527);
or U6680 (N_6680,N_6569,N_6586);
nor U6681 (N_6681,N_6093,N_6311);
nand U6682 (N_6682,N_6477,N_6372);
or U6683 (N_6683,N_6329,N_6072);
or U6684 (N_6684,N_6140,N_6007);
nand U6685 (N_6685,N_6001,N_6256);
xor U6686 (N_6686,N_6153,N_6201);
xnor U6687 (N_6687,N_6224,N_6104);
or U6688 (N_6688,N_6064,N_6147);
nand U6689 (N_6689,N_6316,N_6518);
or U6690 (N_6690,N_6246,N_6476);
and U6691 (N_6691,N_6030,N_6312);
or U6692 (N_6692,N_6384,N_6270);
and U6693 (N_6693,N_6597,N_6083);
and U6694 (N_6694,N_6373,N_6550);
or U6695 (N_6695,N_6381,N_6595);
nand U6696 (N_6696,N_6002,N_6500);
and U6697 (N_6697,N_6288,N_6452);
nor U6698 (N_6698,N_6590,N_6326);
or U6699 (N_6699,N_6185,N_6186);
or U6700 (N_6700,N_6370,N_6050);
or U6701 (N_6701,N_6195,N_6468);
and U6702 (N_6702,N_6265,N_6541);
or U6703 (N_6703,N_6298,N_6155);
or U6704 (N_6704,N_6192,N_6315);
or U6705 (N_6705,N_6506,N_6493);
and U6706 (N_6706,N_6151,N_6574);
or U6707 (N_6707,N_6442,N_6339);
or U6708 (N_6708,N_6397,N_6276);
xor U6709 (N_6709,N_6258,N_6434);
xor U6710 (N_6710,N_6208,N_6490);
and U6711 (N_6711,N_6161,N_6519);
nand U6712 (N_6712,N_6321,N_6539);
or U6713 (N_6713,N_6051,N_6441);
xnor U6714 (N_6714,N_6168,N_6520);
nor U6715 (N_6715,N_6165,N_6359);
or U6716 (N_6716,N_6469,N_6127);
and U6717 (N_6717,N_6338,N_6440);
nor U6718 (N_6718,N_6377,N_6088);
and U6719 (N_6719,N_6585,N_6572);
xor U6720 (N_6720,N_6033,N_6343);
nand U6721 (N_6721,N_6532,N_6196);
or U6722 (N_6722,N_6478,N_6325);
xnor U6723 (N_6723,N_6210,N_6090);
or U6724 (N_6724,N_6425,N_6076);
nor U6725 (N_6725,N_6489,N_6011);
or U6726 (N_6726,N_6084,N_6524);
or U6727 (N_6727,N_6383,N_6491);
nand U6728 (N_6728,N_6396,N_6444);
or U6729 (N_6729,N_6047,N_6271);
nand U6730 (N_6730,N_6239,N_6542);
nor U6731 (N_6731,N_6341,N_6302);
xnor U6732 (N_6732,N_6587,N_6040);
or U6733 (N_6733,N_6158,N_6408);
nor U6734 (N_6734,N_6466,N_6299);
and U6735 (N_6735,N_6065,N_6551);
and U6736 (N_6736,N_6294,N_6067);
xor U6737 (N_6737,N_6058,N_6345);
and U6738 (N_6738,N_6277,N_6351);
nor U6739 (N_6739,N_6126,N_6540);
nor U6740 (N_6740,N_6443,N_6037);
and U6741 (N_6741,N_6410,N_6036);
nor U6742 (N_6742,N_6096,N_6145);
nor U6743 (N_6743,N_6528,N_6043);
nor U6744 (N_6744,N_6435,N_6068);
nand U6745 (N_6745,N_6352,N_6332);
and U6746 (N_6746,N_6306,N_6573);
or U6747 (N_6747,N_6203,N_6252);
or U6748 (N_6748,N_6184,N_6350);
xnor U6749 (N_6749,N_6418,N_6480);
and U6750 (N_6750,N_6484,N_6552);
nor U6751 (N_6751,N_6150,N_6385);
and U6752 (N_6752,N_6544,N_6034);
nor U6753 (N_6753,N_6175,N_6053);
nand U6754 (N_6754,N_6035,N_6303);
nand U6755 (N_6755,N_6580,N_6219);
xor U6756 (N_6756,N_6598,N_6546);
or U6757 (N_6757,N_6226,N_6428);
nand U6758 (N_6758,N_6212,N_6485);
nor U6759 (N_6759,N_6358,N_6445);
nor U6760 (N_6760,N_6052,N_6220);
nor U6761 (N_6761,N_6199,N_6259);
nor U6762 (N_6762,N_6085,N_6559);
and U6763 (N_6763,N_6179,N_6041);
nor U6764 (N_6764,N_6049,N_6438);
nor U6765 (N_6765,N_6014,N_6463);
or U6766 (N_6766,N_6078,N_6562);
and U6767 (N_6767,N_6423,N_6369);
or U6768 (N_6768,N_6038,N_6367);
and U6769 (N_6769,N_6594,N_6591);
and U6770 (N_6770,N_6082,N_6465);
or U6771 (N_6771,N_6505,N_6516);
nor U6772 (N_6772,N_6182,N_6080);
and U6773 (N_6773,N_6092,N_6160);
nor U6774 (N_6774,N_6130,N_6249);
or U6775 (N_6775,N_6547,N_6123);
nand U6776 (N_6776,N_6314,N_6565);
nand U6777 (N_6777,N_6121,N_6282);
and U6778 (N_6778,N_6132,N_6206);
nand U6779 (N_6779,N_6529,N_6044);
or U6780 (N_6780,N_6154,N_6456);
or U6781 (N_6781,N_6094,N_6021);
or U6782 (N_6782,N_6426,N_6401);
nor U6783 (N_6783,N_6512,N_6473);
nand U6784 (N_6784,N_6335,N_6062);
nor U6785 (N_6785,N_6475,N_6570);
nor U6786 (N_6786,N_6398,N_6101);
nand U6787 (N_6787,N_6136,N_6116);
nand U6788 (N_6788,N_6230,N_6419);
nor U6789 (N_6789,N_6251,N_6416);
xor U6790 (N_6790,N_6257,N_6488);
or U6791 (N_6791,N_6349,N_6494);
nor U6792 (N_6792,N_6099,N_6455);
and U6793 (N_6793,N_6364,N_6114);
and U6794 (N_6794,N_6133,N_6227);
nand U6795 (N_6795,N_6279,N_6536);
or U6796 (N_6796,N_6174,N_6344);
nor U6797 (N_6797,N_6521,N_6020);
xnor U6798 (N_6798,N_6139,N_6016);
nor U6799 (N_6799,N_6304,N_6336);
or U6800 (N_6800,N_6194,N_6234);
xnor U6801 (N_6801,N_6482,N_6448);
and U6802 (N_6802,N_6087,N_6567);
nor U6803 (N_6803,N_6229,N_6537);
and U6804 (N_6804,N_6217,N_6113);
xnor U6805 (N_6805,N_6190,N_6374);
nor U6806 (N_6806,N_6061,N_6535);
and U6807 (N_6807,N_6549,N_6105);
xnor U6808 (N_6808,N_6414,N_6470);
nand U6809 (N_6809,N_6283,N_6361);
nor U6810 (N_6810,N_6457,N_6584);
and U6811 (N_6811,N_6582,N_6110);
nor U6812 (N_6812,N_6310,N_6322);
nand U6813 (N_6813,N_6244,N_6202);
and U6814 (N_6814,N_6486,N_6032);
or U6815 (N_6815,N_6313,N_6296);
nor U6816 (N_6816,N_6272,N_6342);
nand U6817 (N_6817,N_6556,N_6379);
and U6818 (N_6818,N_6386,N_6487);
and U6819 (N_6819,N_6166,N_6006);
and U6820 (N_6820,N_6137,N_6218);
nor U6821 (N_6821,N_6371,N_6449);
nor U6822 (N_6822,N_6171,N_6238);
nor U6823 (N_6823,N_6197,N_6511);
nand U6824 (N_6824,N_6557,N_6460);
nand U6825 (N_6825,N_6563,N_6109);
or U6826 (N_6826,N_6509,N_6278);
nor U6827 (N_6827,N_6142,N_6112);
or U6828 (N_6828,N_6593,N_6498);
nand U6829 (N_6829,N_6510,N_6079);
or U6830 (N_6830,N_6013,N_6464);
nor U6831 (N_6831,N_6564,N_6387);
nand U6832 (N_6832,N_6437,N_6241);
xnor U6833 (N_6833,N_6213,N_6391);
nand U6834 (N_6834,N_6081,N_6330);
xor U6835 (N_6835,N_6554,N_6178);
nand U6836 (N_6836,N_6012,N_6548);
nor U6837 (N_6837,N_6008,N_6003);
and U6838 (N_6838,N_6453,N_6167);
or U6839 (N_6839,N_6245,N_6575);
and U6840 (N_6840,N_6180,N_6353);
and U6841 (N_6841,N_6327,N_6200);
nand U6842 (N_6842,N_6048,N_6380);
nand U6843 (N_6843,N_6015,N_6402);
and U6844 (N_6844,N_6378,N_6117);
nor U6845 (N_6845,N_6215,N_6422);
xor U6846 (N_6846,N_6432,N_6157);
nor U6847 (N_6847,N_6446,N_6596);
and U6848 (N_6848,N_6553,N_6429);
nand U6849 (N_6849,N_6411,N_6056);
nor U6850 (N_6850,N_6095,N_6207);
or U6851 (N_6851,N_6558,N_6074);
or U6852 (N_6852,N_6046,N_6039);
nand U6853 (N_6853,N_6543,N_6260);
and U6854 (N_6854,N_6555,N_6568);
and U6855 (N_6855,N_6169,N_6159);
or U6856 (N_6856,N_6305,N_6119);
nor U6857 (N_6857,N_6301,N_6253);
or U6858 (N_6858,N_6424,N_6421);
or U6859 (N_6859,N_6089,N_6583);
nor U6860 (N_6860,N_6393,N_6176);
nand U6861 (N_6861,N_6317,N_6025);
or U6862 (N_6862,N_6045,N_6177);
and U6863 (N_6863,N_6356,N_6436);
and U6864 (N_6864,N_6579,N_6022);
or U6865 (N_6865,N_6479,N_6400);
xnor U6866 (N_6866,N_6077,N_6333);
nor U6867 (N_6867,N_6228,N_6560);
nand U6868 (N_6868,N_6223,N_6293);
xnor U6869 (N_6869,N_6004,N_6027);
or U6870 (N_6870,N_6000,N_6522);
xor U6871 (N_6871,N_6394,N_6501);
nand U6872 (N_6872,N_6250,N_6409);
or U6873 (N_6873,N_6106,N_6318);
and U6874 (N_6874,N_6009,N_6135);
nand U6875 (N_6875,N_6205,N_6496);
nor U6876 (N_6876,N_6275,N_6131);
and U6877 (N_6877,N_6181,N_6102);
or U6878 (N_6878,N_6308,N_6173);
or U6879 (N_6879,N_6143,N_6023);
nand U6880 (N_6880,N_6471,N_6427);
or U6881 (N_6881,N_6183,N_6162);
xnor U6882 (N_6882,N_6098,N_6100);
and U6883 (N_6883,N_6497,N_6071);
or U6884 (N_6884,N_6255,N_6214);
nand U6885 (N_6885,N_6405,N_6413);
nand U6886 (N_6886,N_6287,N_6472);
nand U6887 (N_6887,N_6124,N_6122);
or U6888 (N_6888,N_6042,N_6382);
nand U6889 (N_6889,N_6017,N_6538);
nand U6890 (N_6890,N_6269,N_6525);
nor U6891 (N_6891,N_6274,N_6450);
or U6892 (N_6892,N_6430,N_6589);
nor U6893 (N_6893,N_6263,N_6266);
and U6894 (N_6894,N_6514,N_6433);
nand U6895 (N_6895,N_6281,N_6073);
xor U6896 (N_6896,N_6447,N_6144);
nor U6897 (N_6897,N_6237,N_6390);
or U6898 (N_6898,N_6309,N_6267);
or U6899 (N_6899,N_6286,N_6431);
and U6900 (N_6900,N_6518,N_6026);
or U6901 (N_6901,N_6381,N_6013);
nand U6902 (N_6902,N_6223,N_6151);
or U6903 (N_6903,N_6545,N_6276);
nand U6904 (N_6904,N_6508,N_6056);
or U6905 (N_6905,N_6309,N_6521);
or U6906 (N_6906,N_6564,N_6262);
nor U6907 (N_6907,N_6454,N_6408);
nor U6908 (N_6908,N_6175,N_6147);
and U6909 (N_6909,N_6290,N_6038);
and U6910 (N_6910,N_6294,N_6073);
xor U6911 (N_6911,N_6063,N_6121);
and U6912 (N_6912,N_6013,N_6124);
xor U6913 (N_6913,N_6092,N_6118);
nand U6914 (N_6914,N_6148,N_6526);
nand U6915 (N_6915,N_6005,N_6166);
nand U6916 (N_6916,N_6370,N_6203);
and U6917 (N_6917,N_6060,N_6543);
or U6918 (N_6918,N_6480,N_6399);
or U6919 (N_6919,N_6068,N_6043);
nand U6920 (N_6920,N_6273,N_6533);
or U6921 (N_6921,N_6229,N_6059);
or U6922 (N_6922,N_6218,N_6156);
and U6923 (N_6923,N_6304,N_6120);
nand U6924 (N_6924,N_6470,N_6129);
nor U6925 (N_6925,N_6225,N_6323);
nor U6926 (N_6926,N_6385,N_6269);
or U6927 (N_6927,N_6508,N_6437);
and U6928 (N_6928,N_6461,N_6356);
nor U6929 (N_6929,N_6224,N_6002);
and U6930 (N_6930,N_6243,N_6257);
nor U6931 (N_6931,N_6042,N_6328);
xor U6932 (N_6932,N_6463,N_6472);
nor U6933 (N_6933,N_6077,N_6345);
nand U6934 (N_6934,N_6342,N_6042);
and U6935 (N_6935,N_6000,N_6014);
or U6936 (N_6936,N_6546,N_6189);
nand U6937 (N_6937,N_6239,N_6389);
and U6938 (N_6938,N_6200,N_6488);
xor U6939 (N_6939,N_6407,N_6264);
and U6940 (N_6940,N_6546,N_6011);
nor U6941 (N_6941,N_6465,N_6125);
nand U6942 (N_6942,N_6235,N_6553);
nor U6943 (N_6943,N_6007,N_6386);
or U6944 (N_6944,N_6449,N_6353);
nor U6945 (N_6945,N_6012,N_6274);
nand U6946 (N_6946,N_6138,N_6527);
nand U6947 (N_6947,N_6323,N_6116);
nand U6948 (N_6948,N_6085,N_6580);
nor U6949 (N_6949,N_6266,N_6564);
nor U6950 (N_6950,N_6545,N_6093);
nand U6951 (N_6951,N_6094,N_6044);
nand U6952 (N_6952,N_6398,N_6553);
and U6953 (N_6953,N_6555,N_6372);
nand U6954 (N_6954,N_6135,N_6043);
nand U6955 (N_6955,N_6504,N_6487);
xor U6956 (N_6956,N_6046,N_6410);
and U6957 (N_6957,N_6456,N_6308);
or U6958 (N_6958,N_6414,N_6358);
nand U6959 (N_6959,N_6452,N_6450);
nor U6960 (N_6960,N_6396,N_6074);
or U6961 (N_6961,N_6407,N_6156);
and U6962 (N_6962,N_6420,N_6368);
and U6963 (N_6963,N_6297,N_6166);
or U6964 (N_6964,N_6579,N_6391);
nand U6965 (N_6965,N_6009,N_6287);
nor U6966 (N_6966,N_6077,N_6209);
or U6967 (N_6967,N_6385,N_6449);
and U6968 (N_6968,N_6550,N_6264);
xnor U6969 (N_6969,N_6212,N_6318);
nand U6970 (N_6970,N_6364,N_6067);
nand U6971 (N_6971,N_6418,N_6181);
xor U6972 (N_6972,N_6064,N_6463);
xnor U6973 (N_6973,N_6107,N_6361);
and U6974 (N_6974,N_6077,N_6012);
or U6975 (N_6975,N_6438,N_6096);
nand U6976 (N_6976,N_6453,N_6403);
nor U6977 (N_6977,N_6100,N_6561);
or U6978 (N_6978,N_6327,N_6445);
and U6979 (N_6979,N_6219,N_6093);
or U6980 (N_6980,N_6059,N_6109);
nor U6981 (N_6981,N_6087,N_6590);
and U6982 (N_6982,N_6476,N_6148);
or U6983 (N_6983,N_6540,N_6528);
nor U6984 (N_6984,N_6566,N_6345);
xnor U6985 (N_6985,N_6435,N_6046);
or U6986 (N_6986,N_6094,N_6322);
nand U6987 (N_6987,N_6517,N_6188);
nor U6988 (N_6988,N_6506,N_6335);
and U6989 (N_6989,N_6050,N_6470);
and U6990 (N_6990,N_6256,N_6259);
nand U6991 (N_6991,N_6004,N_6063);
or U6992 (N_6992,N_6198,N_6021);
nand U6993 (N_6993,N_6220,N_6502);
or U6994 (N_6994,N_6475,N_6130);
nand U6995 (N_6995,N_6093,N_6533);
and U6996 (N_6996,N_6150,N_6251);
or U6997 (N_6997,N_6458,N_6158);
or U6998 (N_6998,N_6145,N_6223);
nor U6999 (N_6999,N_6445,N_6307);
xnor U7000 (N_7000,N_6280,N_6228);
nand U7001 (N_7001,N_6412,N_6121);
or U7002 (N_7002,N_6159,N_6048);
xor U7003 (N_7003,N_6494,N_6171);
or U7004 (N_7004,N_6299,N_6193);
nor U7005 (N_7005,N_6202,N_6137);
nor U7006 (N_7006,N_6483,N_6359);
nor U7007 (N_7007,N_6360,N_6072);
nor U7008 (N_7008,N_6500,N_6449);
or U7009 (N_7009,N_6010,N_6325);
xnor U7010 (N_7010,N_6503,N_6342);
or U7011 (N_7011,N_6157,N_6295);
xnor U7012 (N_7012,N_6070,N_6039);
or U7013 (N_7013,N_6129,N_6469);
and U7014 (N_7014,N_6032,N_6332);
or U7015 (N_7015,N_6092,N_6029);
nand U7016 (N_7016,N_6211,N_6391);
nand U7017 (N_7017,N_6486,N_6111);
nand U7018 (N_7018,N_6467,N_6421);
nor U7019 (N_7019,N_6277,N_6274);
xor U7020 (N_7020,N_6294,N_6504);
nand U7021 (N_7021,N_6267,N_6505);
and U7022 (N_7022,N_6249,N_6082);
nand U7023 (N_7023,N_6521,N_6235);
or U7024 (N_7024,N_6460,N_6233);
xor U7025 (N_7025,N_6358,N_6305);
or U7026 (N_7026,N_6203,N_6408);
nand U7027 (N_7027,N_6429,N_6016);
nand U7028 (N_7028,N_6233,N_6127);
or U7029 (N_7029,N_6048,N_6214);
nand U7030 (N_7030,N_6496,N_6275);
or U7031 (N_7031,N_6354,N_6039);
or U7032 (N_7032,N_6192,N_6288);
nor U7033 (N_7033,N_6127,N_6117);
nor U7034 (N_7034,N_6017,N_6532);
nand U7035 (N_7035,N_6494,N_6393);
and U7036 (N_7036,N_6404,N_6508);
or U7037 (N_7037,N_6188,N_6460);
or U7038 (N_7038,N_6031,N_6164);
xnor U7039 (N_7039,N_6111,N_6456);
nor U7040 (N_7040,N_6353,N_6054);
nor U7041 (N_7041,N_6104,N_6131);
and U7042 (N_7042,N_6342,N_6205);
nand U7043 (N_7043,N_6368,N_6330);
nor U7044 (N_7044,N_6136,N_6117);
and U7045 (N_7045,N_6100,N_6539);
nor U7046 (N_7046,N_6490,N_6062);
xor U7047 (N_7047,N_6331,N_6144);
nor U7048 (N_7048,N_6585,N_6470);
nor U7049 (N_7049,N_6015,N_6123);
nand U7050 (N_7050,N_6415,N_6465);
nor U7051 (N_7051,N_6491,N_6407);
xor U7052 (N_7052,N_6214,N_6277);
or U7053 (N_7053,N_6133,N_6303);
or U7054 (N_7054,N_6108,N_6003);
nor U7055 (N_7055,N_6158,N_6156);
xnor U7056 (N_7056,N_6382,N_6137);
nand U7057 (N_7057,N_6437,N_6543);
nand U7058 (N_7058,N_6588,N_6044);
nor U7059 (N_7059,N_6026,N_6593);
nand U7060 (N_7060,N_6038,N_6138);
or U7061 (N_7061,N_6488,N_6177);
or U7062 (N_7062,N_6147,N_6089);
nand U7063 (N_7063,N_6321,N_6404);
nor U7064 (N_7064,N_6080,N_6229);
nand U7065 (N_7065,N_6360,N_6244);
or U7066 (N_7066,N_6099,N_6527);
nand U7067 (N_7067,N_6003,N_6276);
nand U7068 (N_7068,N_6506,N_6093);
or U7069 (N_7069,N_6420,N_6231);
xnor U7070 (N_7070,N_6274,N_6474);
and U7071 (N_7071,N_6017,N_6063);
xnor U7072 (N_7072,N_6308,N_6216);
xnor U7073 (N_7073,N_6109,N_6165);
or U7074 (N_7074,N_6398,N_6467);
nand U7075 (N_7075,N_6133,N_6568);
and U7076 (N_7076,N_6448,N_6056);
nand U7077 (N_7077,N_6006,N_6444);
nand U7078 (N_7078,N_6471,N_6201);
nor U7079 (N_7079,N_6431,N_6492);
or U7080 (N_7080,N_6344,N_6351);
and U7081 (N_7081,N_6030,N_6348);
or U7082 (N_7082,N_6569,N_6300);
nor U7083 (N_7083,N_6200,N_6225);
or U7084 (N_7084,N_6167,N_6014);
xnor U7085 (N_7085,N_6216,N_6150);
and U7086 (N_7086,N_6575,N_6322);
nor U7087 (N_7087,N_6195,N_6492);
nor U7088 (N_7088,N_6154,N_6288);
nand U7089 (N_7089,N_6307,N_6064);
nand U7090 (N_7090,N_6094,N_6348);
nor U7091 (N_7091,N_6295,N_6434);
nor U7092 (N_7092,N_6274,N_6360);
and U7093 (N_7093,N_6276,N_6179);
and U7094 (N_7094,N_6336,N_6424);
or U7095 (N_7095,N_6303,N_6587);
or U7096 (N_7096,N_6271,N_6570);
and U7097 (N_7097,N_6067,N_6479);
nor U7098 (N_7098,N_6589,N_6326);
or U7099 (N_7099,N_6207,N_6068);
and U7100 (N_7100,N_6409,N_6246);
nor U7101 (N_7101,N_6562,N_6407);
nor U7102 (N_7102,N_6522,N_6352);
or U7103 (N_7103,N_6208,N_6310);
nor U7104 (N_7104,N_6490,N_6435);
and U7105 (N_7105,N_6449,N_6421);
nand U7106 (N_7106,N_6080,N_6438);
and U7107 (N_7107,N_6430,N_6042);
nor U7108 (N_7108,N_6132,N_6114);
and U7109 (N_7109,N_6497,N_6561);
nand U7110 (N_7110,N_6290,N_6578);
nand U7111 (N_7111,N_6062,N_6089);
and U7112 (N_7112,N_6262,N_6553);
xnor U7113 (N_7113,N_6086,N_6329);
nand U7114 (N_7114,N_6361,N_6174);
and U7115 (N_7115,N_6182,N_6554);
and U7116 (N_7116,N_6599,N_6422);
or U7117 (N_7117,N_6579,N_6397);
and U7118 (N_7118,N_6251,N_6388);
and U7119 (N_7119,N_6596,N_6461);
and U7120 (N_7120,N_6239,N_6512);
xor U7121 (N_7121,N_6107,N_6366);
or U7122 (N_7122,N_6236,N_6564);
nor U7123 (N_7123,N_6550,N_6496);
nand U7124 (N_7124,N_6083,N_6406);
nor U7125 (N_7125,N_6382,N_6497);
or U7126 (N_7126,N_6461,N_6580);
nand U7127 (N_7127,N_6392,N_6539);
xnor U7128 (N_7128,N_6376,N_6295);
or U7129 (N_7129,N_6508,N_6594);
nand U7130 (N_7130,N_6413,N_6246);
and U7131 (N_7131,N_6344,N_6579);
nand U7132 (N_7132,N_6497,N_6366);
nor U7133 (N_7133,N_6398,N_6057);
or U7134 (N_7134,N_6579,N_6445);
xnor U7135 (N_7135,N_6483,N_6242);
xnor U7136 (N_7136,N_6268,N_6576);
nand U7137 (N_7137,N_6205,N_6353);
nor U7138 (N_7138,N_6198,N_6435);
nor U7139 (N_7139,N_6257,N_6157);
and U7140 (N_7140,N_6148,N_6299);
and U7141 (N_7141,N_6030,N_6168);
nor U7142 (N_7142,N_6054,N_6379);
xor U7143 (N_7143,N_6488,N_6065);
and U7144 (N_7144,N_6116,N_6552);
nand U7145 (N_7145,N_6106,N_6548);
or U7146 (N_7146,N_6463,N_6177);
nand U7147 (N_7147,N_6260,N_6449);
nand U7148 (N_7148,N_6330,N_6332);
nand U7149 (N_7149,N_6316,N_6117);
nor U7150 (N_7150,N_6123,N_6262);
and U7151 (N_7151,N_6383,N_6167);
xnor U7152 (N_7152,N_6062,N_6579);
nor U7153 (N_7153,N_6007,N_6206);
and U7154 (N_7154,N_6034,N_6236);
nor U7155 (N_7155,N_6444,N_6406);
and U7156 (N_7156,N_6255,N_6535);
and U7157 (N_7157,N_6591,N_6295);
or U7158 (N_7158,N_6056,N_6556);
nand U7159 (N_7159,N_6068,N_6545);
and U7160 (N_7160,N_6024,N_6390);
nand U7161 (N_7161,N_6230,N_6555);
or U7162 (N_7162,N_6008,N_6129);
nand U7163 (N_7163,N_6248,N_6436);
nor U7164 (N_7164,N_6107,N_6226);
and U7165 (N_7165,N_6522,N_6534);
nand U7166 (N_7166,N_6584,N_6523);
nand U7167 (N_7167,N_6363,N_6269);
nor U7168 (N_7168,N_6028,N_6498);
nor U7169 (N_7169,N_6361,N_6521);
and U7170 (N_7170,N_6147,N_6431);
nor U7171 (N_7171,N_6031,N_6491);
or U7172 (N_7172,N_6450,N_6177);
or U7173 (N_7173,N_6370,N_6289);
and U7174 (N_7174,N_6356,N_6324);
nor U7175 (N_7175,N_6085,N_6159);
nand U7176 (N_7176,N_6474,N_6093);
nand U7177 (N_7177,N_6326,N_6030);
and U7178 (N_7178,N_6058,N_6529);
nand U7179 (N_7179,N_6452,N_6004);
nor U7180 (N_7180,N_6361,N_6352);
nor U7181 (N_7181,N_6323,N_6368);
xor U7182 (N_7182,N_6261,N_6103);
nand U7183 (N_7183,N_6333,N_6344);
nand U7184 (N_7184,N_6582,N_6102);
and U7185 (N_7185,N_6496,N_6230);
or U7186 (N_7186,N_6034,N_6538);
or U7187 (N_7187,N_6576,N_6419);
or U7188 (N_7188,N_6255,N_6415);
nor U7189 (N_7189,N_6076,N_6552);
and U7190 (N_7190,N_6258,N_6032);
or U7191 (N_7191,N_6222,N_6369);
nor U7192 (N_7192,N_6157,N_6456);
nor U7193 (N_7193,N_6392,N_6228);
or U7194 (N_7194,N_6493,N_6461);
and U7195 (N_7195,N_6207,N_6564);
nand U7196 (N_7196,N_6390,N_6548);
xor U7197 (N_7197,N_6188,N_6500);
or U7198 (N_7198,N_6513,N_6153);
nor U7199 (N_7199,N_6040,N_6473);
or U7200 (N_7200,N_6726,N_6837);
and U7201 (N_7201,N_6978,N_7085);
or U7202 (N_7202,N_6681,N_7143);
nor U7203 (N_7203,N_7066,N_6635);
xor U7204 (N_7204,N_7113,N_7021);
nor U7205 (N_7205,N_7073,N_7128);
nand U7206 (N_7206,N_6953,N_7010);
and U7207 (N_7207,N_7058,N_7199);
nor U7208 (N_7208,N_7116,N_6925);
or U7209 (N_7209,N_7072,N_6943);
and U7210 (N_7210,N_6650,N_7093);
or U7211 (N_7211,N_6668,N_7032);
nor U7212 (N_7212,N_6771,N_6696);
nor U7213 (N_7213,N_6753,N_6890);
nor U7214 (N_7214,N_6881,N_6966);
nor U7215 (N_7215,N_6895,N_6908);
nor U7216 (N_7216,N_7151,N_6861);
or U7217 (N_7217,N_6942,N_6945);
or U7218 (N_7218,N_6827,N_6735);
nor U7219 (N_7219,N_6889,N_6995);
or U7220 (N_7220,N_6713,N_7037);
nor U7221 (N_7221,N_6814,N_6644);
nor U7222 (N_7222,N_7098,N_6630);
nor U7223 (N_7223,N_6704,N_7114);
or U7224 (N_7224,N_7124,N_6843);
or U7225 (N_7225,N_7140,N_6677);
or U7226 (N_7226,N_6783,N_7071);
and U7227 (N_7227,N_7180,N_7189);
and U7228 (N_7228,N_6860,N_7193);
and U7229 (N_7229,N_7104,N_6705);
nor U7230 (N_7230,N_7156,N_6817);
nor U7231 (N_7231,N_7059,N_6937);
and U7232 (N_7232,N_7185,N_6980);
xor U7233 (N_7233,N_6679,N_7133);
or U7234 (N_7234,N_7139,N_6897);
and U7235 (N_7235,N_7144,N_7109);
nor U7236 (N_7236,N_6764,N_6812);
and U7237 (N_7237,N_6938,N_7070);
and U7238 (N_7238,N_7042,N_6797);
nand U7239 (N_7239,N_6902,N_7158);
or U7240 (N_7240,N_7017,N_6905);
nor U7241 (N_7241,N_6858,N_6744);
nor U7242 (N_7242,N_7012,N_6687);
and U7243 (N_7243,N_6620,N_6856);
and U7244 (N_7244,N_6605,N_7122);
nand U7245 (N_7245,N_6730,N_7164);
nor U7246 (N_7246,N_6976,N_6907);
nor U7247 (N_7247,N_6693,N_6944);
xor U7248 (N_7248,N_6683,N_6863);
nand U7249 (N_7249,N_6802,N_6854);
nand U7250 (N_7250,N_6891,N_6643);
nor U7251 (N_7251,N_6639,N_6865);
nor U7252 (N_7252,N_6874,N_6940);
nand U7253 (N_7253,N_7147,N_6675);
or U7254 (N_7254,N_7165,N_6707);
or U7255 (N_7255,N_6965,N_7137);
nand U7256 (N_7256,N_6746,N_6714);
nand U7257 (N_7257,N_6997,N_6737);
or U7258 (N_7258,N_6637,N_6975);
nor U7259 (N_7259,N_6694,N_7024);
nand U7260 (N_7260,N_7054,N_7065);
xor U7261 (N_7261,N_7095,N_6653);
and U7262 (N_7262,N_6934,N_7049);
and U7263 (N_7263,N_6826,N_6972);
nor U7264 (N_7264,N_7105,N_6834);
or U7265 (N_7265,N_7050,N_7026);
or U7266 (N_7266,N_6760,N_6723);
and U7267 (N_7267,N_7002,N_6659);
nor U7268 (N_7268,N_6671,N_6959);
nor U7269 (N_7269,N_6821,N_6721);
nand U7270 (N_7270,N_6625,N_6672);
and U7271 (N_7271,N_6724,N_6631);
nand U7272 (N_7272,N_7062,N_7060);
xor U7273 (N_7273,N_6815,N_7061);
xor U7274 (N_7274,N_7029,N_7120);
nor U7275 (N_7275,N_7119,N_7087);
and U7276 (N_7276,N_6948,N_6847);
or U7277 (N_7277,N_6871,N_6801);
xor U7278 (N_7278,N_6919,N_6985);
xnor U7279 (N_7279,N_6602,N_7184);
or U7280 (N_7280,N_7125,N_6646);
or U7281 (N_7281,N_7004,N_6793);
and U7282 (N_7282,N_7076,N_6816);
nor U7283 (N_7283,N_6688,N_6885);
and U7284 (N_7284,N_7097,N_7123);
and U7285 (N_7285,N_7025,N_7134);
xnor U7286 (N_7286,N_6661,N_6851);
nand U7287 (N_7287,N_6647,N_6846);
or U7288 (N_7288,N_6779,N_6917);
or U7289 (N_7289,N_6725,N_6962);
nand U7290 (N_7290,N_6927,N_7051);
nand U7291 (N_7291,N_6869,N_6800);
or U7292 (N_7292,N_7009,N_7039);
nand U7293 (N_7293,N_6669,N_6780);
or U7294 (N_7294,N_6804,N_7179);
xor U7295 (N_7295,N_7118,N_6667);
nor U7296 (N_7296,N_7015,N_6986);
xnor U7297 (N_7297,N_6622,N_6623);
nor U7298 (N_7298,N_6690,N_6989);
and U7299 (N_7299,N_6657,N_6910);
nor U7300 (N_7300,N_6712,N_7044);
and U7301 (N_7301,N_6642,N_6685);
and U7302 (N_7302,N_7033,N_7077);
nand U7303 (N_7303,N_6798,N_7187);
and U7304 (N_7304,N_6952,N_6706);
and U7305 (N_7305,N_6731,N_7078);
and U7306 (N_7306,N_6795,N_6903);
and U7307 (N_7307,N_6619,N_7052);
and U7308 (N_7308,N_6929,N_6673);
nand U7309 (N_7309,N_6709,N_6720);
nand U7310 (N_7310,N_6697,N_6883);
nand U7311 (N_7311,N_6809,N_6762);
nand U7312 (N_7312,N_7074,N_6813);
and U7313 (N_7313,N_7075,N_7023);
nand U7314 (N_7314,N_6752,N_6923);
or U7315 (N_7315,N_6845,N_7106);
and U7316 (N_7316,N_6935,N_7053);
nand U7317 (N_7317,N_7102,N_7013);
and U7318 (N_7318,N_6992,N_6993);
and U7319 (N_7319,N_6634,N_6877);
xor U7320 (N_7320,N_6606,N_7150);
and U7321 (N_7321,N_7145,N_7166);
xnor U7322 (N_7322,N_7048,N_7141);
or U7323 (N_7323,N_6703,N_6930);
or U7324 (N_7324,N_6939,N_6676);
and U7325 (N_7325,N_6699,N_6951);
xor U7326 (N_7326,N_7001,N_6887);
and U7327 (N_7327,N_7090,N_7148);
or U7328 (N_7328,N_6916,N_6828);
nand U7329 (N_7329,N_6880,N_6768);
nand U7330 (N_7330,N_6600,N_6716);
nand U7331 (N_7331,N_7176,N_6777);
xor U7332 (N_7332,N_6769,N_7019);
xnor U7333 (N_7333,N_7082,N_7173);
nand U7334 (N_7334,N_7136,N_6882);
and U7335 (N_7335,N_6741,N_6691);
or U7336 (N_7336,N_6894,N_7038);
or U7337 (N_7337,N_6689,N_6695);
or U7338 (N_7338,N_7080,N_6607);
nor U7339 (N_7339,N_6662,N_6660);
or U7340 (N_7340,N_7055,N_7130);
nand U7341 (N_7341,N_6609,N_6928);
xor U7342 (N_7342,N_6641,N_6901);
nand U7343 (N_7343,N_6784,N_6615);
nor U7344 (N_7344,N_6765,N_6692);
nand U7345 (N_7345,N_7020,N_6864);
nand U7346 (N_7346,N_7110,N_6954);
or U7347 (N_7347,N_6899,N_6651);
nand U7348 (N_7348,N_7043,N_6718);
and U7349 (N_7349,N_7028,N_6983);
or U7350 (N_7350,N_7194,N_6857);
nand U7351 (N_7351,N_6656,N_6808);
xor U7352 (N_7352,N_6742,N_6949);
or U7353 (N_7353,N_6941,N_7132);
or U7354 (N_7354,N_7172,N_7159);
or U7355 (N_7355,N_6610,N_6743);
nor U7356 (N_7356,N_6819,N_7181);
and U7357 (N_7357,N_7153,N_6960);
or U7358 (N_7358,N_6926,N_7067);
and U7359 (N_7359,N_7152,N_7046);
nand U7360 (N_7360,N_6969,N_6727);
xor U7361 (N_7361,N_6790,N_6896);
nor U7362 (N_7362,N_6608,N_6739);
xnor U7363 (N_7363,N_6613,N_6991);
or U7364 (N_7364,N_6789,N_6776);
or U7365 (N_7365,N_7191,N_7197);
xor U7366 (N_7366,N_6849,N_7099);
or U7367 (N_7367,N_6958,N_7107);
nor U7368 (N_7368,N_6898,N_6799);
nand U7369 (N_7369,N_6994,N_7057);
nor U7370 (N_7370,N_6832,N_7040);
or U7371 (N_7371,N_7081,N_6794);
and U7372 (N_7372,N_7036,N_6870);
and U7373 (N_7373,N_6686,N_6875);
nand U7374 (N_7374,N_6604,N_6807);
nand U7375 (N_7375,N_6628,N_7041);
nor U7376 (N_7376,N_7171,N_6868);
or U7377 (N_7377,N_6664,N_6756);
nand U7378 (N_7378,N_6732,N_6838);
nor U7379 (N_7379,N_7192,N_6782);
xnor U7380 (N_7380,N_7167,N_6886);
xnor U7381 (N_7381,N_7175,N_6829);
nor U7382 (N_7382,N_6850,N_7047);
nand U7383 (N_7383,N_6775,N_6663);
or U7384 (N_7384,N_6747,N_7177);
nor U7385 (N_7385,N_6792,N_6633);
or U7386 (N_7386,N_6805,N_6738);
nor U7387 (N_7387,N_6774,N_6648);
and U7388 (N_7388,N_6911,N_6785);
and U7389 (N_7389,N_6974,N_6824);
nand U7390 (N_7390,N_6786,N_6638);
xnor U7391 (N_7391,N_6733,N_6987);
or U7392 (N_7392,N_7084,N_6936);
and U7393 (N_7393,N_7011,N_7092);
nor U7394 (N_7394,N_6766,N_6968);
nand U7395 (N_7395,N_6682,N_7101);
nand U7396 (N_7396,N_6624,N_7121);
and U7397 (N_7397,N_6867,N_6734);
xnor U7398 (N_7398,N_6670,N_6770);
nand U7399 (N_7399,N_6736,N_6893);
nand U7400 (N_7400,N_6754,N_6629);
nor U7401 (N_7401,N_6652,N_6839);
nor U7402 (N_7402,N_7127,N_6618);
nand U7403 (N_7403,N_6666,N_6778);
xor U7404 (N_7404,N_7182,N_6702);
and U7405 (N_7405,N_7045,N_7068);
nand U7406 (N_7406,N_7014,N_6844);
and U7407 (N_7407,N_6900,N_6645);
and U7408 (N_7408,N_6632,N_6866);
and U7409 (N_7409,N_6678,N_6967);
nand U7410 (N_7410,N_6788,N_6708);
or U7411 (N_7411,N_6684,N_6932);
xor U7412 (N_7412,N_6918,N_6921);
nor U7413 (N_7413,N_6914,N_6873);
and U7414 (N_7414,N_7135,N_6823);
or U7415 (N_7415,N_6626,N_7168);
or U7416 (N_7416,N_6970,N_6654);
nand U7417 (N_7417,N_6822,N_7018);
or U7418 (N_7418,N_7196,N_6841);
nand U7419 (N_7419,N_6621,N_7174);
or U7420 (N_7420,N_6761,N_7154);
or U7421 (N_7421,N_7091,N_6950);
nand U7422 (N_7422,N_7146,N_6710);
and U7423 (N_7423,N_6825,N_7142);
and U7424 (N_7424,N_6988,N_6722);
or U7425 (N_7425,N_7183,N_6617);
and U7426 (N_7426,N_7016,N_7169);
and U7427 (N_7427,N_6655,N_7008);
nor U7428 (N_7428,N_7138,N_7086);
nand U7429 (N_7429,N_6998,N_6830);
nor U7430 (N_7430,N_6852,N_6872);
and U7431 (N_7431,N_7035,N_6833);
nand U7432 (N_7432,N_6781,N_6842);
nor U7433 (N_7433,N_6715,N_6755);
nand U7434 (N_7434,N_6749,N_6915);
nand U7435 (N_7435,N_6904,N_7186);
and U7436 (N_7436,N_7160,N_7000);
or U7437 (N_7437,N_7157,N_7103);
nand U7438 (N_7438,N_6946,N_6878);
nand U7439 (N_7439,N_6924,N_7126);
and U7440 (N_7440,N_6674,N_7003);
nand U7441 (N_7441,N_7178,N_6888);
and U7442 (N_7442,N_7027,N_6981);
and U7443 (N_7443,N_6996,N_7115);
nand U7444 (N_7444,N_6748,N_6810);
xor U7445 (N_7445,N_6612,N_6711);
nand U7446 (N_7446,N_6835,N_7155);
nand U7447 (N_7447,N_6611,N_6763);
or U7448 (N_7448,N_6963,N_6811);
xnor U7449 (N_7449,N_6758,N_6719);
nand U7450 (N_7450,N_7149,N_7088);
and U7451 (N_7451,N_6892,N_6853);
or U7452 (N_7452,N_6840,N_7195);
and U7453 (N_7453,N_7131,N_6767);
nor U7454 (N_7454,N_7100,N_6957);
nor U7455 (N_7455,N_7117,N_6717);
and U7456 (N_7456,N_6649,N_6955);
nor U7457 (N_7457,N_7096,N_7112);
nand U7458 (N_7458,N_6999,N_6879);
or U7459 (N_7459,N_7005,N_7089);
and U7460 (N_7460,N_6933,N_7190);
and U7461 (N_7461,N_7034,N_6982);
or U7462 (N_7462,N_6680,N_6836);
nor U7463 (N_7463,N_6990,N_7129);
nand U7464 (N_7464,N_6665,N_6956);
xnor U7465 (N_7465,N_7007,N_6876);
nand U7466 (N_7466,N_7064,N_6701);
and U7467 (N_7467,N_6906,N_6971);
and U7468 (N_7468,N_6796,N_6728);
nor U7469 (N_7469,N_6820,N_7163);
nor U7470 (N_7470,N_7094,N_6787);
nor U7471 (N_7471,N_7031,N_6922);
nand U7472 (N_7472,N_6603,N_6614);
or U7473 (N_7473,N_6658,N_6912);
and U7474 (N_7474,N_6909,N_7162);
nand U7475 (N_7475,N_7063,N_7188);
or U7476 (N_7476,N_6947,N_6848);
xor U7477 (N_7477,N_6698,N_7006);
or U7478 (N_7478,N_6616,N_6803);
nand U7479 (N_7479,N_6979,N_6984);
xor U7480 (N_7480,N_6884,N_6745);
or U7481 (N_7481,N_6751,N_7069);
or U7482 (N_7482,N_6750,N_6791);
nor U7483 (N_7483,N_6740,N_7161);
xor U7484 (N_7484,N_6759,N_6931);
nand U7485 (N_7485,N_6806,N_6627);
or U7486 (N_7486,N_6964,N_6818);
or U7487 (N_7487,N_6640,N_7022);
and U7488 (N_7488,N_7079,N_6729);
nor U7489 (N_7489,N_6920,N_6913);
nor U7490 (N_7490,N_7056,N_6757);
nand U7491 (N_7491,N_6859,N_7108);
nand U7492 (N_7492,N_7111,N_6700);
and U7493 (N_7493,N_6772,N_6855);
nor U7494 (N_7494,N_6973,N_6636);
nand U7495 (N_7495,N_7170,N_6831);
nand U7496 (N_7496,N_7198,N_6977);
nor U7497 (N_7497,N_6601,N_7083);
xor U7498 (N_7498,N_6961,N_6862);
or U7499 (N_7499,N_7030,N_6773);
or U7500 (N_7500,N_6870,N_6816);
or U7501 (N_7501,N_7133,N_6681);
nor U7502 (N_7502,N_6800,N_6833);
nor U7503 (N_7503,N_6781,N_7136);
nor U7504 (N_7504,N_6940,N_7049);
xnor U7505 (N_7505,N_6696,N_6662);
nand U7506 (N_7506,N_6799,N_6675);
and U7507 (N_7507,N_7110,N_6602);
or U7508 (N_7508,N_7099,N_6685);
nor U7509 (N_7509,N_6637,N_6755);
or U7510 (N_7510,N_6723,N_6605);
or U7511 (N_7511,N_6987,N_6939);
and U7512 (N_7512,N_7010,N_7171);
xnor U7513 (N_7513,N_6796,N_7109);
and U7514 (N_7514,N_6989,N_6823);
nand U7515 (N_7515,N_6970,N_6911);
or U7516 (N_7516,N_7051,N_7103);
nand U7517 (N_7517,N_6833,N_6817);
nor U7518 (N_7518,N_7148,N_6991);
nand U7519 (N_7519,N_6775,N_7164);
or U7520 (N_7520,N_7104,N_7091);
and U7521 (N_7521,N_7085,N_6904);
or U7522 (N_7522,N_6648,N_7046);
nand U7523 (N_7523,N_7013,N_7181);
nand U7524 (N_7524,N_6864,N_7081);
nor U7525 (N_7525,N_6728,N_6610);
or U7526 (N_7526,N_7169,N_6969);
and U7527 (N_7527,N_6789,N_6900);
or U7528 (N_7528,N_6966,N_6651);
xnor U7529 (N_7529,N_7120,N_6943);
and U7530 (N_7530,N_7075,N_7000);
nand U7531 (N_7531,N_6826,N_7076);
nor U7532 (N_7532,N_7085,N_6732);
nor U7533 (N_7533,N_6626,N_6723);
nor U7534 (N_7534,N_6835,N_6719);
or U7535 (N_7535,N_6736,N_6715);
or U7536 (N_7536,N_6708,N_6970);
or U7537 (N_7537,N_6859,N_6907);
nand U7538 (N_7538,N_6792,N_6636);
or U7539 (N_7539,N_6809,N_7127);
or U7540 (N_7540,N_7050,N_6619);
and U7541 (N_7541,N_6902,N_7073);
or U7542 (N_7542,N_6814,N_6796);
nand U7543 (N_7543,N_6794,N_6689);
nor U7544 (N_7544,N_7072,N_6629);
and U7545 (N_7545,N_6677,N_6982);
nand U7546 (N_7546,N_6628,N_6651);
and U7547 (N_7547,N_6860,N_7029);
and U7548 (N_7548,N_7090,N_7071);
nand U7549 (N_7549,N_6933,N_6775);
or U7550 (N_7550,N_6797,N_6966);
or U7551 (N_7551,N_7190,N_6865);
nand U7552 (N_7552,N_6735,N_7034);
and U7553 (N_7553,N_6925,N_6638);
nand U7554 (N_7554,N_7151,N_7170);
or U7555 (N_7555,N_6629,N_6778);
or U7556 (N_7556,N_6781,N_7111);
xnor U7557 (N_7557,N_7136,N_6727);
nor U7558 (N_7558,N_6757,N_6712);
nand U7559 (N_7559,N_7116,N_6733);
nand U7560 (N_7560,N_6781,N_6818);
nand U7561 (N_7561,N_6700,N_6749);
and U7562 (N_7562,N_7137,N_6861);
and U7563 (N_7563,N_7169,N_6795);
and U7564 (N_7564,N_6959,N_6874);
nand U7565 (N_7565,N_7027,N_7099);
or U7566 (N_7566,N_6790,N_6651);
or U7567 (N_7567,N_6976,N_7055);
nor U7568 (N_7568,N_7184,N_6917);
or U7569 (N_7569,N_7121,N_6969);
nor U7570 (N_7570,N_6894,N_6620);
or U7571 (N_7571,N_6707,N_6908);
nor U7572 (N_7572,N_6905,N_6837);
nand U7573 (N_7573,N_6776,N_6993);
xor U7574 (N_7574,N_6976,N_6824);
nor U7575 (N_7575,N_7081,N_6648);
and U7576 (N_7576,N_6692,N_6640);
nor U7577 (N_7577,N_6620,N_6731);
nor U7578 (N_7578,N_7058,N_6972);
and U7579 (N_7579,N_6991,N_6917);
nand U7580 (N_7580,N_6726,N_7019);
nor U7581 (N_7581,N_7116,N_6674);
nor U7582 (N_7582,N_7143,N_7105);
nor U7583 (N_7583,N_6673,N_6652);
or U7584 (N_7584,N_7175,N_7184);
or U7585 (N_7585,N_6756,N_6842);
and U7586 (N_7586,N_6922,N_6819);
nor U7587 (N_7587,N_6837,N_6812);
nor U7588 (N_7588,N_6710,N_6783);
nor U7589 (N_7589,N_6700,N_7139);
or U7590 (N_7590,N_7099,N_7091);
xnor U7591 (N_7591,N_6926,N_7125);
and U7592 (N_7592,N_6793,N_6636);
nor U7593 (N_7593,N_7082,N_6914);
nor U7594 (N_7594,N_6903,N_6648);
and U7595 (N_7595,N_6814,N_7157);
or U7596 (N_7596,N_6906,N_6845);
nand U7597 (N_7597,N_6981,N_6647);
and U7598 (N_7598,N_6902,N_7179);
xor U7599 (N_7599,N_7039,N_6859);
nor U7600 (N_7600,N_6638,N_7028);
or U7601 (N_7601,N_6888,N_7048);
or U7602 (N_7602,N_7185,N_6744);
and U7603 (N_7603,N_7072,N_6807);
and U7604 (N_7604,N_7080,N_7097);
nand U7605 (N_7605,N_6956,N_7182);
xor U7606 (N_7606,N_6772,N_7074);
and U7607 (N_7607,N_7115,N_6881);
nand U7608 (N_7608,N_6878,N_7079);
nor U7609 (N_7609,N_7028,N_6803);
nor U7610 (N_7610,N_7147,N_6629);
nand U7611 (N_7611,N_6651,N_6896);
and U7612 (N_7612,N_7055,N_6700);
or U7613 (N_7613,N_7145,N_6845);
xor U7614 (N_7614,N_7188,N_7033);
nor U7615 (N_7615,N_7065,N_6838);
nand U7616 (N_7616,N_7061,N_6770);
and U7617 (N_7617,N_6827,N_6879);
and U7618 (N_7618,N_6999,N_7062);
and U7619 (N_7619,N_6817,N_7176);
or U7620 (N_7620,N_7150,N_6846);
or U7621 (N_7621,N_6748,N_6968);
or U7622 (N_7622,N_6896,N_6805);
nor U7623 (N_7623,N_7199,N_7174);
xnor U7624 (N_7624,N_7005,N_6732);
or U7625 (N_7625,N_6908,N_7002);
and U7626 (N_7626,N_6909,N_6801);
nor U7627 (N_7627,N_6845,N_6700);
nand U7628 (N_7628,N_7032,N_6912);
or U7629 (N_7629,N_6991,N_7157);
nand U7630 (N_7630,N_6709,N_6912);
and U7631 (N_7631,N_7025,N_6645);
nand U7632 (N_7632,N_6802,N_7142);
or U7633 (N_7633,N_6897,N_6867);
nor U7634 (N_7634,N_7018,N_7175);
xor U7635 (N_7635,N_6969,N_7052);
or U7636 (N_7636,N_6705,N_6606);
and U7637 (N_7637,N_6906,N_7080);
nor U7638 (N_7638,N_6864,N_6670);
xnor U7639 (N_7639,N_6610,N_6661);
xnor U7640 (N_7640,N_6730,N_6709);
or U7641 (N_7641,N_6750,N_7087);
nor U7642 (N_7642,N_7139,N_7077);
or U7643 (N_7643,N_7063,N_6867);
or U7644 (N_7644,N_6959,N_7045);
nor U7645 (N_7645,N_6937,N_6715);
or U7646 (N_7646,N_6807,N_7091);
nor U7647 (N_7647,N_7065,N_6720);
nor U7648 (N_7648,N_7090,N_7061);
nand U7649 (N_7649,N_6934,N_7118);
and U7650 (N_7650,N_7042,N_6992);
or U7651 (N_7651,N_6828,N_6797);
nor U7652 (N_7652,N_6719,N_7074);
and U7653 (N_7653,N_7196,N_7064);
and U7654 (N_7654,N_6621,N_6706);
nand U7655 (N_7655,N_6819,N_6608);
nand U7656 (N_7656,N_7103,N_7148);
xor U7657 (N_7657,N_7030,N_7061);
and U7658 (N_7658,N_7052,N_6607);
nand U7659 (N_7659,N_6765,N_6625);
nor U7660 (N_7660,N_7096,N_7097);
nor U7661 (N_7661,N_7141,N_7017);
nor U7662 (N_7662,N_6773,N_7158);
nand U7663 (N_7663,N_6951,N_7195);
nor U7664 (N_7664,N_6733,N_7052);
nor U7665 (N_7665,N_6901,N_7185);
nand U7666 (N_7666,N_6916,N_6610);
and U7667 (N_7667,N_6701,N_6758);
xor U7668 (N_7668,N_6976,N_6973);
or U7669 (N_7669,N_6694,N_6868);
or U7670 (N_7670,N_6907,N_6636);
nor U7671 (N_7671,N_7086,N_6901);
and U7672 (N_7672,N_6893,N_6741);
xnor U7673 (N_7673,N_6964,N_7172);
or U7674 (N_7674,N_6906,N_6730);
nand U7675 (N_7675,N_6650,N_6994);
nor U7676 (N_7676,N_7099,N_7031);
nand U7677 (N_7677,N_6877,N_6935);
nor U7678 (N_7678,N_7061,N_6636);
nand U7679 (N_7679,N_7088,N_7095);
nor U7680 (N_7680,N_6717,N_7130);
or U7681 (N_7681,N_7078,N_6681);
nand U7682 (N_7682,N_6731,N_7023);
and U7683 (N_7683,N_6913,N_6828);
and U7684 (N_7684,N_6668,N_7019);
or U7685 (N_7685,N_6913,N_7024);
or U7686 (N_7686,N_6994,N_7016);
and U7687 (N_7687,N_6951,N_6717);
and U7688 (N_7688,N_6871,N_6830);
or U7689 (N_7689,N_6687,N_7076);
nand U7690 (N_7690,N_6986,N_6664);
and U7691 (N_7691,N_7096,N_7192);
nor U7692 (N_7692,N_7176,N_6808);
and U7693 (N_7693,N_6857,N_6705);
and U7694 (N_7694,N_7120,N_6901);
nand U7695 (N_7695,N_6731,N_7027);
nor U7696 (N_7696,N_6843,N_7015);
xnor U7697 (N_7697,N_7053,N_6955);
nand U7698 (N_7698,N_6744,N_6602);
or U7699 (N_7699,N_7023,N_7197);
or U7700 (N_7700,N_7074,N_6792);
or U7701 (N_7701,N_6951,N_7171);
xnor U7702 (N_7702,N_7046,N_7062);
nor U7703 (N_7703,N_7035,N_6861);
and U7704 (N_7704,N_6850,N_6873);
or U7705 (N_7705,N_7103,N_7173);
or U7706 (N_7706,N_6682,N_6795);
nand U7707 (N_7707,N_6912,N_6990);
or U7708 (N_7708,N_6706,N_7136);
and U7709 (N_7709,N_7199,N_6940);
nor U7710 (N_7710,N_7040,N_6657);
nand U7711 (N_7711,N_6882,N_6886);
and U7712 (N_7712,N_6740,N_6961);
or U7713 (N_7713,N_7124,N_7006);
xor U7714 (N_7714,N_7110,N_6666);
or U7715 (N_7715,N_6614,N_7163);
or U7716 (N_7716,N_7092,N_6909);
and U7717 (N_7717,N_7185,N_7153);
and U7718 (N_7718,N_6671,N_6725);
xnor U7719 (N_7719,N_7180,N_7075);
nand U7720 (N_7720,N_6660,N_7125);
or U7721 (N_7721,N_6729,N_7091);
or U7722 (N_7722,N_7106,N_6732);
and U7723 (N_7723,N_6761,N_7036);
or U7724 (N_7724,N_6947,N_6624);
or U7725 (N_7725,N_6951,N_6782);
or U7726 (N_7726,N_6781,N_7066);
xnor U7727 (N_7727,N_7150,N_6789);
or U7728 (N_7728,N_7180,N_7055);
nor U7729 (N_7729,N_7130,N_6901);
nor U7730 (N_7730,N_6752,N_7060);
nand U7731 (N_7731,N_6663,N_6940);
or U7732 (N_7732,N_7034,N_6694);
nand U7733 (N_7733,N_6872,N_6770);
nand U7734 (N_7734,N_6809,N_7037);
nor U7735 (N_7735,N_6624,N_6965);
or U7736 (N_7736,N_6813,N_6738);
xor U7737 (N_7737,N_6761,N_6662);
nand U7738 (N_7738,N_7068,N_7190);
or U7739 (N_7739,N_7008,N_7142);
and U7740 (N_7740,N_6608,N_7147);
and U7741 (N_7741,N_6903,N_6939);
nand U7742 (N_7742,N_6766,N_6825);
and U7743 (N_7743,N_6608,N_6679);
nor U7744 (N_7744,N_7094,N_6829);
nor U7745 (N_7745,N_6967,N_6912);
and U7746 (N_7746,N_7005,N_6740);
nor U7747 (N_7747,N_7065,N_6999);
nor U7748 (N_7748,N_6760,N_6744);
or U7749 (N_7749,N_6666,N_6765);
or U7750 (N_7750,N_7171,N_6729);
xnor U7751 (N_7751,N_6950,N_7133);
nor U7752 (N_7752,N_7051,N_6934);
xnor U7753 (N_7753,N_7021,N_6932);
xor U7754 (N_7754,N_6876,N_7022);
nor U7755 (N_7755,N_6715,N_7158);
and U7756 (N_7756,N_6688,N_6834);
nand U7757 (N_7757,N_7033,N_6861);
or U7758 (N_7758,N_6971,N_6965);
or U7759 (N_7759,N_7179,N_7100);
nand U7760 (N_7760,N_6908,N_7079);
or U7761 (N_7761,N_7169,N_7046);
nand U7762 (N_7762,N_6665,N_7025);
or U7763 (N_7763,N_6718,N_6757);
or U7764 (N_7764,N_6659,N_6651);
xor U7765 (N_7765,N_6704,N_7074);
xor U7766 (N_7766,N_7067,N_6867);
and U7767 (N_7767,N_6824,N_6796);
nand U7768 (N_7768,N_6958,N_7182);
xnor U7769 (N_7769,N_7043,N_7132);
nand U7770 (N_7770,N_7043,N_6841);
and U7771 (N_7771,N_6686,N_6940);
or U7772 (N_7772,N_6894,N_7049);
nand U7773 (N_7773,N_6782,N_6859);
and U7774 (N_7774,N_7012,N_6990);
or U7775 (N_7775,N_6662,N_7193);
or U7776 (N_7776,N_7085,N_6979);
and U7777 (N_7777,N_6730,N_6943);
and U7778 (N_7778,N_6966,N_7067);
nor U7779 (N_7779,N_6995,N_6735);
and U7780 (N_7780,N_6880,N_6811);
or U7781 (N_7781,N_6665,N_6606);
nand U7782 (N_7782,N_6612,N_6925);
and U7783 (N_7783,N_6927,N_6751);
and U7784 (N_7784,N_6624,N_6665);
and U7785 (N_7785,N_7045,N_7091);
and U7786 (N_7786,N_6807,N_6845);
or U7787 (N_7787,N_6858,N_7067);
or U7788 (N_7788,N_6832,N_6694);
nor U7789 (N_7789,N_6802,N_6963);
or U7790 (N_7790,N_6825,N_6829);
nor U7791 (N_7791,N_6714,N_6665);
and U7792 (N_7792,N_6955,N_7121);
and U7793 (N_7793,N_6833,N_6913);
nand U7794 (N_7794,N_6737,N_6842);
or U7795 (N_7795,N_7194,N_7055);
nor U7796 (N_7796,N_7049,N_6723);
and U7797 (N_7797,N_6957,N_6726);
xnor U7798 (N_7798,N_6770,N_6979);
and U7799 (N_7799,N_6939,N_6764);
xor U7800 (N_7800,N_7335,N_7606);
and U7801 (N_7801,N_7629,N_7741);
nor U7802 (N_7802,N_7429,N_7271);
nand U7803 (N_7803,N_7441,N_7776);
nor U7804 (N_7804,N_7495,N_7544);
or U7805 (N_7805,N_7439,N_7506);
nor U7806 (N_7806,N_7669,N_7386);
or U7807 (N_7807,N_7391,N_7282);
nand U7808 (N_7808,N_7460,N_7650);
or U7809 (N_7809,N_7594,N_7225);
and U7810 (N_7810,N_7234,N_7726);
or U7811 (N_7811,N_7336,N_7605);
nand U7812 (N_7812,N_7372,N_7499);
and U7813 (N_7813,N_7643,N_7436);
xor U7814 (N_7814,N_7292,N_7418);
and U7815 (N_7815,N_7541,N_7223);
nor U7816 (N_7816,N_7485,N_7784);
or U7817 (N_7817,N_7707,N_7573);
xnor U7818 (N_7818,N_7510,N_7297);
or U7819 (N_7819,N_7224,N_7240);
or U7820 (N_7820,N_7533,N_7415);
or U7821 (N_7821,N_7284,N_7320);
and U7822 (N_7822,N_7419,N_7483);
nor U7823 (N_7823,N_7263,N_7652);
nor U7824 (N_7824,N_7554,N_7559);
xnor U7825 (N_7825,N_7360,N_7205);
nand U7826 (N_7826,N_7422,N_7376);
xor U7827 (N_7827,N_7791,N_7508);
or U7828 (N_7828,N_7327,N_7574);
nand U7829 (N_7829,N_7789,N_7531);
xor U7830 (N_7830,N_7575,N_7231);
or U7831 (N_7831,N_7543,N_7752);
and U7832 (N_7832,N_7395,N_7494);
or U7833 (N_7833,N_7361,N_7614);
nand U7834 (N_7834,N_7480,N_7555);
or U7835 (N_7835,N_7708,N_7215);
or U7836 (N_7836,N_7449,N_7524);
nand U7837 (N_7837,N_7468,N_7276);
nand U7838 (N_7838,N_7238,N_7763);
nor U7839 (N_7839,N_7298,N_7280);
or U7840 (N_7840,N_7551,N_7651);
nor U7841 (N_7841,N_7775,N_7484);
xor U7842 (N_7842,N_7749,N_7507);
nor U7843 (N_7843,N_7730,N_7232);
nor U7844 (N_7844,N_7607,N_7431);
and U7845 (N_7845,N_7404,N_7777);
nor U7846 (N_7846,N_7388,N_7637);
nor U7847 (N_7847,N_7330,N_7200);
nand U7848 (N_7848,N_7472,N_7665);
and U7849 (N_7849,N_7713,N_7583);
or U7850 (N_7850,N_7244,N_7355);
nor U7851 (N_7851,N_7247,N_7538);
or U7852 (N_7852,N_7307,N_7743);
or U7853 (N_7853,N_7517,N_7679);
nand U7854 (N_7854,N_7430,N_7671);
xor U7855 (N_7855,N_7349,N_7635);
nand U7856 (N_7856,N_7370,N_7414);
nor U7857 (N_7857,N_7359,N_7382);
and U7858 (N_7858,N_7557,N_7778);
or U7859 (N_7859,N_7217,N_7329);
nand U7860 (N_7860,N_7413,N_7765);
nand U7861 (N_7861,N_7619,N_7364);
xnor U7862 (N_7862,N_7428,N_7590);
and U7863 (N_7863,N_7695,N_7731);
xor U7864 (N_7864,N_7464,N_7350);
nor U7865 (N_7865,N_7287,N_7689);
and U7866 (N_7866,N_7666,N_7511);
nand U7867 (N_7867,N_7660,N_7545);
or U7868 (N_7868,N_7337,N_7339);
xor U7869 (N_7869,N_7714,N_7211);
and U7870 (N_7870,N_7332,N_7600);
and U7871 (N_7871,N_7352,N_7257);
nor U7872 (N_7872,N_7486,N_7702);
nor U7873 (N_7873,N_7737,N_7270);
or U7874 (N_7874,N_7539,N_7560);
nor U7875 (N_7875,N_7394,N_7401);
nor U7876 (N_7876,N_7226,N_7479);
and U7877 (N_7877,N_7291,N_7780);
xnor U7878 (N_7878,N_7410,N_7520);
nor U7879 (N_7879,N_7347,N_7723);
or U7880 (N_7880,N_7795,N_7487);
and U7881 (N_7881,N_7721,N_7724);
nor U7882 (N_7882,N_7586,N_7754);
nor U7883 (N_7883,N_7739,N_7374);
or U7884 (N_7884,N_7323,N_7732);
xnor U7885 (N_7885,N_7405,N_7773);
xnor U7886 (N_7886,N_7761,N_7283);
or U7887 (N_7887,N_7406,N_7345);
nand U7888 (N_7888,N_7239,N_7728);
or U7889 (N_7889,N_7546,N_7313);
nor U7890 (N_7890,N_7736,N_7766);
nor U7891 (N_7891,N_7658,N_7326);
nand U7892 (N_7892,N_7793,N_7351);
nand U7893 (N_7893,N_7467,N_7755);
nor U7894 (N_7894,N_7504,N_7624);
nand U7895 (N_7895,N_7657,N_7518);
nor U7896 (N_7896,N_7672,N_7768);
nand U7897 (N_7897,N_7727,N_7204);
nand U7898 (N_7898,N_7709,N_7375);
nand U7899 (N_7899,N_7218,N_7542);
xnor U7900 (N_7900,N_7319,N_7342);
xnor U7901 (N_7901,N_7354,N_7434);
or U7902 (N_7902,N_7309,N_7751);
or U7903 (N_7903,N_7267,N_7403);
or U7904 (N_7904,N_7272,N_7634);
or U7905 (N_7905,N_7278,N_7492);
nor U7906 (N_7906,N_7237,N_7748);
and U7907 (N_7907,N_7788,N_7670);
or U7908 (N_7908,N_7365,N_7409);
nor U7909 (N_7909,N_7633,N_7221);
xor U7910 (N_7910,N_7259,N_7343);
nor U7911 (N_7911,N_7235,N_7601);
and U7912 (N_7912,N_7740,N_7562);
nor U7913 (N_7913,N_7245,N_7710);
nor U7914 (N_7914,N_7774,N_7502);
nand U7915 (N_7915,N_7530,N_7392);
nand U7916 (N_7916,N_7623,N_7536);
xor U7917 (N_7917,N_7233,N_7227);
or U7918 (N_7918,N_7399,N_7592);
xor U7919 (N_7919,N_7498,N_7302);
and U7920 (N_7920,N_7322,N_7346);
nand U7921 (N_7921,N_7523,N_7792);
xnor U7922 (N_7922,N_7423,N_7753);
nand U7923 (N_7923,N_7663,N_7580);
nor U7924 (N_7924,N_7598,N_7703);
nand U7925 (N_7925,N_7675,N_7610);
and U7926 (N_7926,N_7344,N_7328);
nand U7927 (N_7927,N_7496,N_7734);
or U7928 (N_7928,N_7261,N_7550);
nor U7929 (N_7929,N_7626,N_7260);
nand U7930 (N_7930,N_7471,N_7312);
nand U7931 (N_7931,N_7692,N_7785);
or U7932 (N_7932,N_7698,N_7251);
or U7933 (N_7933,N_7742,N_7432);
nor U7934 (N_7934,N_7407,N_7688);
xor U7935 (N_7935,N_7682,N_7293);
xor U7936 (N_7936,N_7604,N_7595);
nor U7937 (N_7937,N_7579,N_7402);
and U7938 (N_7938,N_7602,N_7653);
or U7939 (N_7939,N_7733,N_7711);
and U7940 (N_7940,N_7639,N_7474);
nor U7941 (N_7941,N_7202,N_7760);
or U7942 (N_7942,N_7219,N_7490);
nand U7943 (N_7943,N_7249,N_7582);
or U7944 (N_7944,N_7525,N_7443);
nor U7945 (N_7945,N_7389,N_7717);
nand U7946 (N_7946,N_7540,N_7236);
or U7947 (N_7947,N_7589,N_7676);
or U7948 (N_7948,N_7640,N_7482);
xor U7949 (N_7949,N_7489,N_7662);
nand U7950 (N_7950,N_7248,N_7796);
or U7951 (N_7951,N_7357,N_7288);
or U7952 (N_7952,N_7424,N_7781);
and U7953 (N_7953,N_7253,N_7674);
or U7954 (N_7954,N_7649,N_7201);
and U7955 (N_7955,N_7593,N_7274);
nor U7956 (N_7956,N_7367,N_7447);
nor U7957 (N_7957,N_7497,N_7268);
or U7958 (N_7958,N_7442,N_7416);
nand U7959 (N_7959,N_7371,N_7700);
or U7960 (N_7960,N_7385,N_7456);
xnor U7961 (N_7961,N_7252,N_7577);
xnor U7962 (N_7962,N_7572,N_7515);
nor U7963 (N_7963,N_7420,N_7438);
or U7964 (N_7964,N_7779,N_7631);
and U7965 (N_7965,N_7585,N_7664);
and U7966 (N_7966,N_7750,N_7556);
xor U7967 (N_7967,N_7632,N_7587);
or U7968 (N_7968,N_7308,N_7783);
or U7969 (N_7969,N_7481,N_7466);
and U7970 (N_7970,N_7738,N_7390);
or U7971 (N_7971,N_7417,N_7786);
or U7972 (N_7972,N_7615,N_7501);
nand U7973 (N_7973,N_7668,N_7368);
or U7974 (N_7974,N_7279,N_7565);
or U7975 (N_7975,N_7706,N_7790);
nand U7976 (N_7976,N_7493,N_7620);
and U7977 (N_7977,N_7314,N_7684);
xnor U7978 (N_7978,N_7787,N_7286);
and U7979 (N_7979,N_7210,N_7527);
nand U7980 (N_7980,N_7300,N_7408);
nor U7981 (N_7981,N_7797,N_7655);
nor U7982 (N_7982,N_7681,N_7448);
nor U7983 (N_7983,N_7397,N_7529);
xnor U7984 (N_7984,N_7642,N_7552);
and U7985 (N_7985,N_7597,N_7455);
xor U7986 (N_7986,N_7528,N_7722);
and U7987 (N_7987,N_7366,N_7318);
nor U7988 (N_7988,N_7558,N_7799);
nand U7989 (N_7989,N_7454,N_7720);
or U7990 (N_7990,N_7758,N_7646);
nand U7991 (N_7991,N_7519,N_7680);
and U7992 (N_7992,N_7222,N_7289);
or U7993 (N_7993,N_7630,N_7333);
or U7994 (N_7994,N_7612,N_7609);
and U7995 (N_7995,N_7696,N_7534);
nor U7996 (N_7996,N_7678,N_7697);
nor U7997 (N_7997,N_7563,N_7220);
nor U7998 (N_7998,N_7656,N_7603);
and U7999 (N_7999,N_7522,N_7654);
nor U8000 (N_8000,N_7459,N_7362);
nand U8001 (N_8001,N_7383,N_7453);
nand U8002 (N_8002,N_7532,N_7636);
nand U8003 (N_8003,N_7683,N_7281);
xor U8004 (N_8004,N_7770,N_7452);
nand U8005 (N_8005,N_7621,N_7568);
and U8006 (N_8006,N_7744,N_7513);
and U8007 (N_8007,N_7627,N_7311);
and U8008 (N_8008,N_7509,N_7581);
xor U8009 (N_8009,N_7576,N_7250);
nor U8010 (N_8010,N_7317,N_7491);
nor U8011 (N_8011,N_7353,N_7207);
and U8012 (N_8012,N_7356,N_7378);
nor U8013 (N_8013,N_7475,N_7444);
nor U8014 (N_8014,N_7735,N_7747);
or U8015 (N_8015,N_7659,N_7667);
nand U8016 (N_8016,N_7358,N_7591);
nand U8017 (N_8017,N_7258,N_7704);
nor U8018 (N_8018,N_7798,N_7617);
xnor U8019 (N_8019,N_7771,N_7553);
or U8020 (N_8020,N_7561,N_7254);
or U8021 (N_8021,N_7457,N_7756);
nor U8022 (N_8022,N_7772,N_7571);
or U8023 (N_8023,N_7310,N_7746);
nor U8024 (N_8024,N_7564,N_7321);
xor U8025 (N_8025,N_7398,N_7759);
nor U8026 (N_8026,N_7537,N_7304);
and U8027 (N_8027,N_7569,N_7693);
nand U8028 (N_8028,N_7725,N_7305);
and U8029 (N_8029,N_7584,N_7616);
nand U8030 (N_8030,N_7648,N_7673);
or U8031 (N_8031,N_7295,N_7608);
and U8032 (N_8032,N_7599,N_7285);
nor U8033 (N_8033,N_7451,N_7762);
nor U8034 (N_8034,N_7348,N_7465);
nor U8035 (N_8035,N_7435,N_7387);
nor U8036 (N_8036,N_7625,N_7476);
nor U8037 (N_8037,N_7596,N_7246);
and U8038 (N_8038,N_7265,N_7228);
or U8039 (N_8039,N_7677,N_7477);
or U8040 (N_8040,N_7567,N_7369);
and U8041 (N_8041,N_7208,N_7243);
nand U8042 (N_8042,N_7488,N_7324);
or U8043 (N_8043,N_7463,N_7421);
or U8044 (N_8044,N_7264,N_7549);
nand U8045 (N_8045,N_7478,N_7212);
or U8046 (N_8046,N_7450,N_7437);
xor U8047 (N_8047,N_7690,N_7461);
and U8048 (N_8048,N_7203,N_7262);
nand U8049 (N_8049,N_7611,N_7277);
nor U8050 (N_8050,N_7373,N_7699);
and U8051 (N_8051,N_7715,N_7769);
or U8052 (N_8052,N_7296,N_7411);
or U8053 (N_8053,N_7425,N_7325);
or U8054 (N_8054,N_7315,N_7729);
and U8055 (N_8055,N_7647,N_7712);
nor U8056 (N_8056,N_7214,N_7691);
and U8057 (N_8057,N_7334,N_7381);
nand U8058 (N_8058,N_7213,N_7578);
nand U8059 (N_8059,N_7686,N_7229);
nor U8060 (N_8060,N_7638,N_7618);
or U8061 (N_8061,N_7473,N_7380);
or U8062 (N_8062,N_7782,N_7216);
nand U8063 (N_8063,N_7269,N_7745);
nand U8064 (N_8064,N_7547,N_7719);
xnor U8065 (N_8065,N_7396,N_7256);
xnor U8066 (N_8066,N_7512,N_7427);
or U8067 (N_8067,N_7521,N_7685);
and U8068 (N_8068,N_7303,N_7242);
nor U8069 (N_8069,N_7273,N_7767);
nor U8070 (N_8070,N_7412,N_7230);
nand U8071 (N_8071,N_7458,N_7514);
or U8072 (N_8072,N_7462,N_7400);
and U8073 (N_8073,N_7694,N_7363);
or U8074 (N_8074,N_7379,N_7566);
and U8075 (N_8075,N_7426,N_7469);
or U8076 (N_8076,N_7628,N_7516);
or U8077 (N_8077,N_7433,N_7687);
or U8078 (N_8078,N_7266,N_7301);
or U8079 (N_8079,N_7341,N_7718);
nor U8080 (N_8080,N_7331,N_7526);
nand U8081 (N_8081,N_7306,N_7570);
nor U8082 (N_8082,N_7209,N_7794);
nor U8083 (N_8083,N_7340,N_7548);
nand U8084 (N_8084,N_7535,N_7290);
and U8085 (N_8085,N_7384,N_7338);
nand U8086 (N_8086,N_7299,N_7622);
nand U8087 (N_8087,N_7641,N_7440);
nor U8088 (N_8088,N_7377,N_7505);
nor U8089 (N_8089,N_7470,N_7316);
nand U8090 (N_8090,N_7701,N_7206);
nand U8091 (N_8091,N_7613,N_7503);
or U8092 (N_8092,N_7446,N_7445);
nor U8093 (N_8093,N_7393,N_7645);
and U8094 (N_8094,N_7705,N_7500);
or U8095 (N_8095,N_7644,N_7757);
nor U8096 (N_8096,N_7716,N_7661);
nor U8097 (N_8097,N_7294,N_7764);
xnor U8098 (N_8098,N_7255,N_7275);
nand U8099 (N_8099,N_7241,N_7588);
xor U8100 (N_8100,N_7476,N_7465);
or U8101 (N_8101,N_7492,N_7336);
or U8102 (N_8102,N_7391,N_7524);
or U8103 (N_8103,N_7415,N_7602);
or U8104 (N_8104,N_7546,N_7727);
xor U8105 (N_8105,N_7482,N_7736);
nand U8106 (N_8106,N_7434,N_7660);
or U8107 (N_8107,N_7657,N_7387);
nor U8108 (N_8108,N_7772,N_7524);
nand U8109 (N_8109,N_7235,N_7323);
and U8110 (N_8110,N_7469,N_7665);
nand U8111 (N_8111,N_7695,N_7679);
or U8112 (N_8112,N_7746,N_7762);
and U8113 (N_8113,N_7227,N_7342);
or U8114 (N_8114,N_7409,N_7535);
or U8115 (N_8115,N_7756,N_7539);
nand U8116 (N_8116,N_7293,N_7559);
nand U8117 (N_8117,N_7631,N_7511);
nor U8118 (N_8118,N_7779,N_7308);
nor U8119 (N_8119,N_7613,N_7504);
or U8120 (N_8120,N_7309,N_7738);
xor U8121 (N_8121,N_7727,N_7778);
and U8122 (N_8122,N_7268,N_7718);
xor U8123 (N_8123,N_7768,N_7773);
nand U8124 (N_8124,N_7313,N_7642);
xnor U8125 (N_8125,N_7631,N_7758);
and U8126 (N_8126,N_7663,N_7529);
or U8127 (N_8127,N_7299,N_7742);
nor U8128 (N_8128,N_7578,N_7648);
or U8129 (N_8129,N_7375,N_7233);
and U8130 (N_8130,N_7406,N_7576);
nand U8131 (N_8131,N_7702,N_7361);
or U8132 (N_8132,N_7556,N_7664);
and U8133 (N_8133,N_7407,N_7540);
nor U8134 (N_8134,N_7256,N_7260);
xor U8135 (N_8135,N_7422,N_7323);
nand U8136 (N_8136,N_7546,N_7720);
nand U8137 (N_8137,N_7548,N_7375);
nor U8138 (N_8138,N_7254,N_7304);
nor U8139 (N_8139,N_7539,N_7487);
nor U8140 (N_8140,N_7386,N_7562);
nor U8141 (N_8141,N_7705,N_7704);
or U8142 (N_8142,N_7336,N_7548);
and U8143 (N_8143,N_7582,N_7265);
nor U8144 (N_8144,N_7521,N_7377);
xor U8145 (N_8145,N_7212,N_7685);
nor U8146 (N_8146,N_7267,N_7534);
or U8147 (N_8147,N_7340,N_7602);
and U8148 (N_8148,N_7679,N_7549);
nand U8149 (N_8149,N_7338,N_7489);
or U8150 (N_8150,N_7323,N_7478);
or U8151 (N_8151,N_7242,N_7639);
nor U8152 (N_8152,N_7688,N_7303);
and U8153 (N_8153,N_7590,N_7214);
nor U8154 (N_8154,N_7454,N_7499);
nor U8155 (N_8155,N_7555,N_7630);
and U8156 (N_8156,N_7265,N_7535);
or U8157 (N_8157,N_7692,N_7299);
xnor U8158 (N_8158,N_7704,N_7599);
nand U8159 (N_8159,N_7535,N_7557);
and U8160 (N_8160,N_7690,N_7200);
xor U8161 (N_8161,N_7285,N_7247);
nand U8162 (N_8162,N_7252,N_7712);
or U8163 (N_8163,N_7271,N_7550);
xnor U8164 (N_8164,N_7202,N_7363);
and U8165 (N_8165,N_7767,N_7266);
nor U8166 (N_8166,N_7593,N_7457);
nand U8167 (N_8167,N_7680,N_7753);
nor U8168 (N_8168,N_7679,N_7625);
and U8169 (N_8169,N_7320,N_7429);
nand U8170 (N_8170,N_7485,N_7721);
and U8171 (N_8171,N_7613,N_7759);
and U8172 (N_8172,N_7720,N_7618);
nand U8173 (N_8173,N_7323,N_7227);
or U8174 (N_8174,N_7223,N_7518);
or U8175 (N_8175,N_7466,N_7217);
nor U8176 (N_8176,N_7260,N_7380);
and U8177 (N_8177,N_7717,N_7206);
or U8178 (N_8178,N_7494,N_7417);
or U8179 (N_8179,N_7633,N_7210);
nor U8180 (N_8180,N_7358,N_7486);
nor U8181 (N_8181,N_7407,N_7435);
nand U8182 (N_8182,N_7613,N_7475);
nor U8183 (N_8183,N_7742,N_7526);
or U8184 (N_8184,N_7426,N_7327);
nand U8185 (N_8185,N_7516,N_7650);
and U8186 (N_8186,N_7748,N_7230);
or U8187 (N_8187,N_7625,N_7542);
and U8188 (N_8188,N_7406,N_7768);
or U8189 (N_8189,N_7477,N_7298);
and U8190 (N_8190,N_7380,N_7689);
nor U8191 (N_8191,N_7383,N_7717);
nor U8192 (N_8192,N_7442,N_7428);
xor U8193 (N_8193,N_7373,N_7653);
nand U8194 (N_8194,N_7783,N_7462);
nand U8195 (N_8195,N_7568,N_7361);
nor U8196 (N_8196,N_7513,N_7662);
nand U8197 (N_8197,N_7498,N_7375);
nor U8198 (N_8198,N_7753,N_7747);
nor U8199 (N_8199,N_7434,N_7284);
nor U8200 (N_8200,N_7224,N_7690);
xor U8201 (N_8201,N_7222,N_7320);
and U8202 (N_8202,N_7440,N_7653);
nand U8203 (N_8203,N_7257,N_7782);
xor U8204 (N_8204,N_7596,N_7440);
and U8205 (N_8205,N_7443,N_7418);
nand U8206 (N_8206,N_7567,N_7552);
nor U8207 (N_8207,N_7733,N_7500);
nor U8208 (N_8208,N_7557,N_7797);
or U8209 (N_8209,N_7774,N_7572);
nor U8210 (N_8210,N_7667,N_7409);
or U8211 (N_8211,N_7619,N_7738);
or U8212 (N_8212,N_7587,N_7798);
and U8213 (N_8213,N_7727,N_7642);
and U8214 (N_8214,N_7223,N_7276);
nor U8215 (N_8215,N_7772,N_7507);
and U8216 (N_8216,N_7415,N_7474);
nor U8217 (N_8217,N_7730,N_7540);
nor U8218 (N_8218,N_7634,N_7743);
nand U8219 (N_8219,N_7463,N_7287);
or U8220 (N_8220,N_7282,N_7594);
nand U8221 (N_8221,N_7621,N_7352);
xor U8222 (N_8222,N_7724,N_7593);
nand U8223 (N_8223,N_7625,N_7769);
nand U8224 (N_8224,N_7711,N_7700);
or U8225 (N_8225,N_7574,N_7509);
nor U8226 (N_8226,N_7520,N_7773);
nand U8227 (N_8227,N_7482,N_7501);
nor U8228 (N_8228,N_7725,N_7687);
xnor U8229 (N_8229,N_7406,N_7690);
and U8230 (N_8230,N_7593,N_7630);
or U8231 (N_8231,N_7395,N_7632);
and U8232 (N_8232,N_7793,N_7771);
xnor U8233 (N_8233,N_7799,N_7322);
or U8234 (N_8234,N_7212,N_7776);
nand U8235 (N_8235,N_7416,N_7346);
xnor U8236 (N_8236,N_7563,N_7494);
or U8237 (N_8237,N_7552,N_7471);
nor U8238 (N_8238,N_7748,N_7771);
xnor U8239 (N_8239,N_7784,N_7720);
and U8240 (N_8240,N_7794,N_7708);
nand U8241 (N_8241,N_7314,N_7313);
nand U8242 (N_8242,N_7734,N_7205);
and U8243 (N_8243,N_7575,N_7444);
nor U8244 (N_8244,N_7468,N_7666);
or U8245 (N_8245,N_7724,N_7349);
or U8246 (N_8246,N_7753,N_7603);
xnor U8247 (N_8247,N_7439,N_7422);
xnor U8248 (N_8248,N_7538,N_7342);
or U8249 (N_8249,N_7372,N_7752);
nand U8250 (N_8250,N_7308,N_7457);
nand U8251 (N_8251,N_7430,N_7395);
or U8252 (N_8252,N_7298,N_7700);
and U8253 (N_8253,N_7536,N_7290);
and U8254 (N_8254,N_7214,N_7797);
nand U8255 (N_8255,N_7438,N_7245);
xnor U8256 (N_8256,N_7734,N_7248);
nor U8257 (N_8257,N_7244,N_7711);
xnor U8258 (N_8258,N_7363,N_7426);
or U8259 (N_8259,N_7546,N_7469);
xor U8260 (N_8260,N_7432,N_7461);
or U8261 (N_8261,N_7385,N_7659);
nor U8262 (N_8262,N_7493,N_7353);
or U8263 (N_8263,N_7577,N_7203);
and U8264 (N_8264,N_7415,N_7341);
xor U8265 (N_8265,N_7219,N_7320);
and U8266 (N_8266,N_7282,N_7712);
nor U8267 (N_8267,N_7689,N_7468);
and U8268 (N_8268,N_7758,N_7524);
nor U8269 (N_8269,N_7613,N_7737);
nand U8270 (N_8270,N_7700,N_7499);
or U8271 (N_8271,N_7655,N_7653);
and U8272 (N_8272,N_7294,N_7669);
or U8273 (N_8273,N_7247,N_7687);
nor U8274 (N_8274,N_7764,N_7738);
nand U8275 (N_8275,N_7355,N_7762);
nor U8276 (N_8276,N_7214,N_7735);
nand U8277 (N_8277,N_7640,N_7528);
xnor U8278 (N_8278,N_7503,N_7745);
nand U8279 (N_8279,N_7419,N_7314);
nand U8280 (N_8280,N_7668,N_7481);
nand U8281 (N_8281,N_7355,N_7612);
and U8282 (N_8282,N_7776,N_7296);
nor U8283 (N_8283,N_7482,N_7597);
or U8284 (N_8284,N_7625,N_7649);
or U8285 (N_8285,N_7388,N_7473);
xnor U8286 (N_8286,N_7686,N_7448);
and U8287 (N_8287,N_7524,N_7612);
and U8288 (N_8288,N_7336,N_7275);
nor U8289 (N_8289,N_7573,N_7506);
and U8290 (N_8290,N_7717,N_7265);
and U8291 (N_8291,N_7781,N_7220);
nand U8292 (N_8292,N_7489,N_7484);
or U8293 (N_8293,N_7424,N_7788);
or U8294 (N_8294,N_7260,N_7669);
or U8295 (N_8295,N_7798,N_7566);
nand U8296 (N_8296,N_7475,N_7455);
nor U8297 (N_8297,N_7456,N_7207);
or U8298 (N_8298,N_7376,N_7497);
and U8299 (N_8299,N_7293,N_7434);
xor U8300 (N_8300,N_7548,N_7480);
nor U8301 (N_8301,N_7528,N_7774);
nor U8302 (N_8302,N_7730,N_7400);
and U8303 (N_8303,N_7457,N_7512);
and U8304 (N_8304,N_7774,N_7339);
nor U8305 (N_8305,N_7536,N_7323);
nor U8306 (N_8306,N_7766,N_7512);
nor U8307 (N_8307,N_7282,N_7411);
or U8308 (N_8308,N_7267,N_7396);
xor U8309 (N_8309,N_7694,N_7557);
xor U8310 (N_8310,N_7321,N_7544);
or U8311 (N_8311,N_7403,N_7234);
and U8312 (N_8312,N_7529,N_7380);
and U8313 (N_8313,N_7730,N_7721);
and U8314 (N_8314,N_7761,N_7612);
and U8315 (N_8315,N_7740,N_7748);
and U8316 (N_8316,N_7373,N_7365);
and U8317 (N_8317,N_7596,N_7640);
or U8318 (N_8318,N_7501,N_7591);
nand U8319 (N_8319,N_7602,N_7591);
or U8320 (N_8320,N_7550,N_7336);
xnor U8321 (N_8321,N_7420,N_7315);
and U8322 (N_8322,N_7793,N_7569);
nand U8323 (N_8323,N_7516,N_7459);
or U8324 (N_8324,N_7453,N_7708);
nor U8325 (N_8325,N_7668,N_7527);
nand U8326 (N_8326,N_7699,N_7578);
xnor U8327 (N_8327,N_7778,N_7586);
or U8328 (N_8328,N_7481,N_7669);
nor U8329 (N_8329,N_7334,N_7737);
and U8330 (N_8330,N_7426,N_7444);
nand U8331 (N_8331,N_7535,N_7448);
and U8332 (N_8332,N_7273,N_7338);
or U8333 (N_8333,N_7264,N_7656);
nand U8334 (N_8334,N_7218,N_7481);
xnor U8335 (N_8335,N_7405,N_7588);
nor U8336 (N_8336,N_7725,N_7370);
nor U8337 (N_8337,N_7417,N_7259);
or U8338 (N_8338,N_7790,N_7664);
nand U8339 (N_8339,N_7535,N_7217);
and U8340 (N_8340,N_7697,N_7329);
and U8341 (N_8341,N_7528,N_7695);
xnor U8342 (N_8342,N_7634,N_7417);
nor U8343 (N_8343,N_7472,N_7564);
or U8344 (N_8344,N_7531,N_7533);
and U8345 (N_8345,N_7603,N_7405);
or U8346 (N_8346,N_7755,N_7547);
nand U8347 (N_8347,N_7247,N_7561);
nor U8348 (N_8348,N_7239,N_7201);
or U8349 (N_8349,N_7479,N_7605);
and U8350 (N_8350,N_7535,N_7735);
xnor U8351 (N_8351,N_7458,N_7673);
and U8352 (N_8352,N_7488,N_7540);
xnor U8353 (N_8353,N_7638,N_7522);
or U8354 (N_8354,N_7455,N_7526);
nand U8355 (N_8355,N_7449,N_7629);
nor U8356 (N_8356,N_7706,N_7626);
nor U8357 (N_8357,N_7793,N_7787);
and U8358 (N_8358,N_7560,N_7778);
and U8359 (N_8359,N_7571,N_7598);
nor U8360 (N_8360,N_7258,N_7727);
xnor U8361 (N_8361,N_7245,N_7546);
nand U8362 (N_8362,N_7404,N_7742);
nand U8363 (N_8363,N_7214,N_7722);
or U8364 (N_8364,N_7202,N_7232);
or U8365 (N_8365,N_7415,N_7567);
nor U8366 (N_8366,N_7771,N_7594);
or U8367 (N_8367,N_7761,N_7474);
and U8368 (N_8368,N_7545,N_7623);
nand U8369 (N_8369,N_7796,N_7462);
or U8370 (N_8370,N_7427,N_7607);
nor U8371 (N_8371,N_7560,N_7640);
and U8372 (N_8372,N_7512,N_7792);
nor U8373 (N_8373,N_7612,N_7591);
nor U8374 (N_8374,N_7210,N_7429);
or U8375 (N_8375,N_7374,N_7537);
or U8376 (N_8376,N_7799,N_7713);
or U8377 (N_8377,N_7760,N_7767);
or U8378 (N_8378,N_7567,N_7690);
and U8379 (N_8379,N_7686,N_7243);
nand U8380 (N_8380,N_7673,N_7504);
or U8381 (N_8381,N_7454,N_7236);
nor U8382 (N_8382,N_7643,N_7568);
nand U8383 (N_8383,N_7667,N_7765);
and U8384 (N_8384,N_7291,N_7467);
or U8385 (N_8385,N_7643,N_7411);
nand U8386 (N_8386,N_7746,N_7694);
or U8387 (N_8387,N_7324,N_7329);
nand U8388 (N_8388,N_7416,N_7408);
nor U8389 (N_8389,N_7307,N_7582);
nor U8390 (N_8390,N_7729,N_7427);
or U8391 (N_8391,N_7705,N_7388);
nand U8392 (N_8392,N_7480,N_7448);
nand U8393 (N_8393,N_7226,N_7273);
and U8394 (N_8394,N_7677,N_7763);
or U8395 (N_8395,N_7774,N_7487);
nor U8396 (N_8396,N_7788,N_7285);
and U8397 (N_8397,N_7571,N_7343);
nand U8398 (N_8398,N_7305,N_7536);
nor U8399 (N_8399,N_7592,N_7496);
xor U8400 (N_8400,N_7905,N_8111);
xnor U8401 (N_8401,N_8327,N_7850);
or U8402 (N_8402,N_7948,N_8348);
or U8403 (N_8403,N_8063,N_7825);
nor U8404 (N_8404,N_7904,N_8231);
or U8405 (N_8405,N_8219,N_8261);
xor U8406 (N_8406,N_7930,N_8113);
nor U8407 (N_8407,N_8095,N_8302);
nand U8408 (N_8408,N_8055,N_7924);
nor U8409 (N_8409,N_8036,N_8286);
nand U8410 (N_8410,N_8053,N_7859);
nand U8411 (N_8411,N_7967,N_8315);
nor U8412 (N_8412,N_8265,N_8382);
nand U8413 (N_8413,N_7835,N_7839);
or U8414 (N_8414,N_8125,N_8180);
and U8415 (N_8415,N_8133,N_8372);
and U8416 (N_8416,N_8078,N_8234);
and U8417 (N_8417,N_8086,N_8105);
nand U8418 (N_8418,N_8209,N_7970);
nor U8419 (N_8419,N_8397,N_8291);
nor U8420 (N_8420,N_8274,N_8168);
xor U8421 (N_8421,N_8172,N_7806);
nand U8422 (N_8422,N_7808,N_8325);
xor U8423 (N_8423,N_8293,N_7996);
and U8424 (N_8424,N_8260,N_7931);
or U8425 (N_8425,N_8049,N_7897);
nor U8426 (N_8426,N_8370,N_7849);
and U8427 (N_8427,N_8004,N_8340);
and U8428 (N_8428,N_7801,N_8159);
or U8429 (N_8429,N_8061,N_7807);
and U8430 (N_8430,N_8236,N_7978);
nand U8431 (N_8431,N_8363,N_7809);
nand U8432 (N_8432,N_8115,N_8385);
nand U8433 (N_8433,N_8203,N_8120);
nand U8434 (N_8434,N_7911,N_7915);
nand U8435 (N_8435,N_8319,N_8222);
and U8436 (N_8436,N_8106,N_8303);
or U8437 (N_8437,N_8289,N_7824);
nand U8438 (N_8438,N_8237,N_7896);
xor U8439 (N_8439,N_8022,N_8057);
nor U8440 (N_8440,N_7995,N_8183);
or U8441 (N_8441,N_7891,N_8322);
and U8442 (N_8442,N_8150,N_8028);
nor U8443 (N_8443,N_8141,N_8254);
or U8444 (N_8444,N_8093,N_8054);
nor U8445 (N_8445,N_8112,N_8332);
nor U8446 (N_8446,N_8246,N_7987);
nor U8447 (N_8447,N_7823,N_8085);
nor U8448 (N_8448,N_8084,N_7984);
nor U8449 (N_8449,N_8077,N_8296);
or U8450 (N_8450,N_8352,N_8301);
nand U8451 (N_8451,N_7886,N_8233);
nand U8452 (N_8452,N_8228,N_8051);
nand U8453 (N_8453,N_7954,N_8288);
nand U8454 (N_8454,N_8094,N_7818);
and U8455 (N_8455,N_8017,N_8074);
xor U8456 (N_8456,N_7854,N_8257);
or U8457 (N_8457,N_8043,N_7945);
nand U8458 (N_8458,N_8294,N_8364);
and U8459 (N_8459,N_7840,N_8258);
or U8460 (N_8460,N_8032,N_8013);
or U8461 (N_8461,N_7941,N_8187);
nor U8462 (N_8462,N_7899,N_7864);
or U8463 (N_8463,N_8048,N_8379);
nand U8464 (N_8464,N_8316,N_8116);
nand U8465 (N_8465,N_8376,N_8267);
nor U8466 (N_8466,N_7884,N_7990);
nor U8467 (N_8467,N_8156,N_7933);
nand U8468 (N_8468,N_8123,N_8068);
nand U8469 (N_8469,N_7985,N_8157);
nand U8470 (N_8470,N_8244,N_8114);
or U8471 (N_8471,N_7857,N_8005);
xnor U8472 (N_8472,N_8213,N_8015);
nor U8473 (N_8473,N_8240,N_8071);
or U8474 (N_8474,N_7953,N_7947);
xor U8475 (N_8475,N_8119,N_7980);
xor U8476 (N_8476,N_8298,N_8135);
and U8477 (N_8477,N_7865,N_8158);
and U8478 (N_8478,N_8179,N_8142);
or U8479 (N_8479,N_8174,N_7964);
or U8480 (N_8480,N_8239,N_8276);
or U8481 (N_8481,N_7977,N_8198);
and U8482 (N_8482,N_8249,N_8349);
and U8483 (N_8483,N_8065,N_8259);
or U8484 (N_8484,N_8290,N_7812);
xor U8485 (N_8485,N_8247,N_8129);
nand U8486 (N_8486,N_7907,N_7895);
nand U8487 (N_8487,N_7830,N_7855);
or U8488 (N_8488,N_8050,N_8381);
xor U8489 (N_8489,N_8147,N_7922);
or U8490 (N_8490,N_8137,N_8058);
nor U8491 (N_8491,N_8285,N_7898);
nand U8492 (N_8492,N_8241,N_7908);
nor U8493 (N_8493,N_7810,N_8171);
nor U8494 (N_8494,N_8270,N_8323);
and U8495 (N_8495,N_8354,N_7943);
nand U8496 (N_8496,N_7975,N_8358);
nand U8497 (N_8497,N_8104,N_7916);
or U8498 (N_8498,N_8040,N_7815);
or U8499 (N_8499,N_8153,N_8221);
nor U8500 (N_8500,N_7923,N_7968);
xor U8501 (N_8501,N_8202,N_8380);
nand U8502 (N_8502,N_8225,N_7860);
nand U8503 (N_8503,N_8357,N_8378);
and U8504 (N_8504,N_8169,N_8072);
nand U8505 (N_8505,N_8038,N_8282);
nand U8506 (N_8506,N_8165,N_7842);
and U8507 (N_8507,N_7955,N_8321);
and U8508 (N_8508,N_8060,N_8229);
nor U8509 (N_8509,N_8096,N_8181);
or U8510 (N_8510,N_8251,N_8278);
nand U8511 (N_8511,N_8189,N_8103);
or U8512 (N_8512,N_8008,N_8374);
and U8513 (N_8513,N_8132,N_7971);
or U8514 (N_8514,N_8182,N_8214);
nor U8515 (N_8515,N_7803,N_8118);
nor U8516 (N_8516,N_7893,N_8018);
or U8517 (N_8517,N_8194,N_8011);
xnor U8518 (N_8518,N_8184,N_7934);
and U8519 (N_8519,N_8064,N_8099);
and U8520 (N_8520,N_7874,N_8305);
and U8521 (N_8521,N_7866,N_7817);
and U8522 (N_8522,N_7832,N_7877);
nor U8523 (N_8523,N_7834,N_8317);
and U8524 (N_8524,N_8146,N_8021);
nor U8525 (N_8525,N_8160,N_7826);
xor U8526 (N_8526,N_7939,N_8083);
and U8527 (N_8527,N_8009,N_8201);
and U8528 (N_8528,N_8207,N_8088);
nand U8529 (N_8529,N_8102,N_8029);
or U8530 (N_8530,N_8066,N_8396);
nand U8531 (N_8531,N_8208,N_8320);
nor U8532 (N_8532,N_8314,N_8101);
or U8533 (N_8533,N_8351,N_8010);
nor U8534 (N_8534,N_7845,N_7997);
nand U8535 (N_8535,N_7982,N_8226);
or U8536 (N_8536,N_8091,N_7833);
nand U8537 (N_8537,N_8131,N_8304);
nand U8538 (N_8538,N_8386,N_8346);
or U8539 (N_8539,N_7813,N_8173);
and U8540 (N_8540,N_7989,N_8359);
and U8541 (N_8541,N_8269,N_8047);
nor U8542 (N_8542,N_7814,N_8324);
nand U8543 (N_8543,N_8161,N_8394);
nor U8544 (N_8544,N_8262,N_8362);
nand U8545 (N_8545,N_8341,N_7862);
xor U8546 (N_8546,N_8309,N_8034);
or U8547 (N_8547,N_7882,N_8069);
or U8548 (N_8548,N_8350,N_8046);
nor U8549 (N_8549,N_8271,N_7991);
nand U8550 (N_8550,N_7951,N_8177);
xnor U8551 (N_8551,N_8395,N_7831);
and U8552 (N_8552,N_7998,N_7875);
nor U8553 (N_8553,N_7868,N_7960);
and U8554 (N_8554,N_8281,N_8242);
nor U8555 (N_8555,N_8031,N_8140);
and U8556 (N_8556,N_7838,N_8090);
or U8557 (N_8557,N_7836,N_8264);
xor U8558 (N_8558,N_7906,N_7867);
nand U8559 (N_8559,N_8188,N_7844);
nand U8560 (N_8560,N_8217,N_7841);
and U8561 (N_8561,N_8126,N_8252);
nor U8562 (N_8562,N_7950,N_8143);
and U8563 (N_8563,N_8330,N_7822);
xor U8564 (N_8564,N_7913,N_8275);
nand U8565 (N_8565,N_8138,N_8014);
nor U8566 (N_8566,N_8367,N_7894);
and U8567 (N_8567,N_7871,N_7914);
or U8568 (N_8568,N_8366,N_8030);
or U8569 (N_8569,N_8124,N_7992);
or U8570 (N_8570,N_7816,N_7974);
nand U8571 (N_8571,N_7940,N_7918);
nor U8572 (N_8572,N_8393,N_8292);
xor U8573 (N_8573,N_8148,N_8307);
and U8574 (N_8574,N_8223,N_7821);
nand U8575 (N_8575,N_8310,N_8154);
nand U8576 (N_8576,N_8087,N_8279);
or U8577 (N_8577,N_7883,N_8335);
and U8578 (N_8578,N_8287,N_7828);
nor U8579 (N_8579,N_8283,N_7928);
nand U8580 (N_8580,N_8311,N_8195);
nor U8581 (N_8581,N_7958,N_7881);
or U8582 (N_8582,N_7851,N_8344);
xnor U8583 (N_8583,N_8206,N_8299);
nor U8584 (N_8584,N_8383,N_8248);
nand U8585 (N_8585,N_8136,N_7843);
nand U8586 (N_8586,N_8334,N_8079);
and U8587 (N_8587,N_7885,N_8243);
nand U8588 (N_8588,N_8059,N_7872);
xor U8589 (N_8589,N_8300,N_7986);
or U8590 (N_8590,N_8062,N_8016);
nor U8591 (N_8591,N_8127,N_8353);
nand U8592 (N_8592,N_7909,N_8277);
xor U8593 (N_8593,N_7935,N_8070);
and U8594 (N_8594,N_8073,N_7936);
nand U8595 (N_8595,N_7863,N_8200);
nor U8596 (N_8596,N_8002,N_8144);
nor U8597 (N_8597,N_8041,N_8220);
nor U8598 (N_8598,N_8199,N_7888);
nor U8599 (N_8599,N_8108,N_7942);
nor U8600 (N_8600,N_8313,N_8109);
or U8601 (N_8601,N_7969,N_7999);
and U8602 (N_8602,N_7861,N_8371);
and U8603 (N_8603,N_8186,N_8192);
xor U8604 (N_8604,N_8333,N_7932);
or U8605 (N_8605,N_8044,N_7912);
or U8606 (N_8606,N_8205,N_8398);
and U8607 (N_8607,N_8045,N_8026);
or U8608 (N_8608,N_7961,N_7889);
or U8609 (N_8609,N_8023,N_8052);
and U8610 (N_8610,N_8175,N_7972);
nor U8611 (N_8611,N_8039,N_7880);
and U8612 (N_8612,N_7827,N_7837);
nor U8613 (N_8613,N_8149,N_8210);
nor U8614 (N_8614,N_8365,N_8295);
nor U8615 (N_8615,N_8284,N_8128);
nand U8616 (N_8616,N_7820,N_7856);
or U8617 (N_8617,N_8092,N_8100);
and U8618 (N_8618,N_8056,N_8339);
and U8619 (N_8619,N_8080,N_8190);
nor U8620 (N_8620,N_7901,N_8193);
nor U8621 (N_8621,N_8391,N_7802);
nand U8622 (N_8622,N_8328,N_7983);
nor U8623 (N_8623,N_8272,N_8117);
nor U8624 (N_8624,N_8042,N_7927);
and U8625 (N_8625,N_7917,N_7946);
and U8626 (N_8626,N_7957,N_7921);
and U8627 (N_8627,N_7965,N_8336);
nor U8628 (N_8628,N_8006,N_7876);
nand U8629 (N_8629,N_8204,N_7829);
nor U8630 (N_8630,N_7902,N_8035);
and U8631 (N_8631,N_7900,N_8268);
or U8632 (N_8632,N_7920,N_8343);
or U8633 (N_8633,N_8347,N_7952);
or U8634 (N_8634,N_8020,N_7994);
or U8635 (N_8635,N_7852,N_8392);
or U8636 (N_8636,N_8176,N_8218);
and U8637 (N_8637,N_8369,N_7944);
and U8638 (N_8638,N_8139,N_8166);
nor U8639 (N_8639,N_8075,N_7976);
and U8640 (N_8640,N_7903,N_8216);
or U8641 (N_8641,N_8297,N_8122);
nand U8642 (N_8642,N_8107,N_7993);
or U8643 (N_8643,N_8110,N_8097);
and U8644 (N_8644,N_7847,N_8329);
and U8645 (N_8645,N_8338,N_8037);
nand U8646 (N_8646,N_8390,N_7800);
xor U8647 (N_8647,N_8191,N_8196);
nand U8648 (N_8648,N_7963,N_8121);
or U8649 (N_8649,N_8253,N_8185);
nand U8650 (N_8650,N_7937,N_7925);
nand U8651 (N_8651,N_7846,N_8388);
xnor U8652 (N_8652,N_8355,N_8326);
or U8653 (N_8653,N_7966,N_7892);
and U8654 (N_8654,N_8361,N_7811);
and U8655 (N_8655,N_8373,N_8306);
xnor U8656 (N_8656,N_8164,N_8081);
nand U8657 (N_8657,N_8375,N_8033);
or U8658 (N_8658,N_7890,N_8163);
and U8659 (N_8659,N_8197,N_7879);
nand U8660 (N_8660,N_7805,N_8001);
and U8661 (N_8661,N_7873,N_7848);
or U8662 (N_8662,N_7959,N_8263);
or U8663 (N_8663,N_7819,N_8337);
or U8664 (N_8664,N_7973,N_8266);
or U8665 (N_8665,N_8356,N_7887);
or U8666 (N_8666,N_8152,N_8318);
nor U8667 (N_8667,N_8003,N_8256);
nand U8668 (N_8668,N_8167,N_7919);
and U8669 (N_8669,N_7979,N_8232);
or U8670 (N_8670,N_8255,N_8089);
nand U8671 (N_8671,N_7938,N_8145);
nor U8672 (N_8672,N_7878,N_7929);
nand U8673 (N_8673,N_8134,N_8211);
nor U8674 (N_8674,N_8389,N_7870);
nand U8675 (N_8675,N_8250,N_8025);
nand U8676 (N_8676,N_7858,N_7853);
or U8677 (N_8677,N_8235,N_8384);
or U8678 (N_8678,N_8162,N_8155);
nand U8679 (N_8679,N_7988,N_8215);
nand U8680 (N_8680,N_8345,N_8212);
nand U8681 (N_8681,N_8387,N_8227);
and U8682 (N_8682,N_7804,N_8224);
nor U8683 (N_8683,N_8098,N_8007);
and U8684 (N_8684,N_8312,N_8230);
nand U8685 (N_8685,N_7962,N_7949);
or U8686 (N_8686,N_8280,N_8273);
nor U8687 (N_8687,N_8019,N_8027);
xnor U8688 (N_8688,N_7956,N_8377);
nor U8689 (N_8689,N_8082,N_8178);
nand U8690 (N_8690,N_8151,N_8012);
xnor U8691 (N_8691,N_8238,N_8024);
and U8692 (N_8692,N_8130,N_8331);
nand U8693 (N_8693,N_8360,N_8368);
and U8694 (N_8694,N_8399,N_7910);
nor U8695 (N_8695,N_8000,N_7981);
nand U8696 (N_8696,N_8342,N_8076);
nor U8697 (N_8697,N_8308,N_8067);
xnor U8698 (N_8698,N_8245,N_7926);
nor U8699 (N_8699,N_7869,N_8170);
or U8700 (N_8700,N_8151,N_8098);
nand U8701 (N_8701,N_8380,N_8087);
nor U8702 (N_8702,N_8318,N_7996);
nand U8703 (N_8703,N_7818,N_8178);
nand U8704 (N_8704,N_8226,N_8166);
xnor U8705 (N_8705,N_8014,N_7957);
xnor U8706 (N_8706,N_8253,N_7971);
nand U8707 (N_8707,N_7816,N_8243);
or U8708 (N_8708,N_8161,N_8127);
and U8709 (N_8709,N_8314,N_8358);
or U8710 (N_8710,N_7890,N_7956);
or U8711 (N_8711,N_7848,N_7978);
nand U8712 (N_8712,N_7951,N_8171);
nor U8713 (N_8713,N_8022,N_8180);
nand U8714 (N_8714,N_8255,N_8167);
or U8715 (N_8715,N_8287,N_7924);
or U8716 (N_8716,N_7835,N_8357);
nand U8717 (N_8717,N_8328,N_8292);
or U8718 (N_8718,N_7913,N_8003);
nor U8719 (N_8719,N_8088,N_8290);
nand U8720 (N_8720,N_7811,N_7813);
nand U8721 (N_8721,N_8370,N_8313);
or U8722 (N_8722,N_7871,N_7925);
and U8723 (N_8723,N_8113,N_8108);
nor U8724 (N_8724,N_7811,N_7907);
xor U8725 (N_8725,N_8394,N_8173);
or U8726 (N_8726,N_8164,N_8133);
nand U8727 (N_8727,N_7877,N_7936);
and U8728 (N_8728,N_8025,N_8178);
or U8729 (N_8729,N_7897,N_8125);
and U8730 (N_8730,N_7991,N_8128);
nand U8731 (N_8731,N_7899,N_8360);
nor U8732 (N_8732,N_8337,N_7815);
nand U8733 (N_8733,N_8281,N_7874);
nor U8734 (N_8734,N_8231,N_8216);
xor U8735 (N_8735,N_8253,N_7942);
nor U8736 (N_8736,N_8320,N_8046);
and U8737 (N_8737,N_8043,N_8187);
or U8738 (N_8738,N_7925,N_7928);
or U8739 (N_8739,N_7861,N_8294);
and U8740 (N_8740,N_8087,N_7874);
xnor U8741 (N_8741,N_8000,N_8152);
nor U8742 (N_8742,N_8354,N_8189);
and U8743 (N_8743,N_8055,N_8032);
and U8744 (N_8744,N_7904,N_7877);
nor U8745 (N_8745,N_8167,N_8226);
nor U8746 (N_8746,N_8388,N_8156);
nand U8747 (N_8747,N_8070,N_7952);
or U8748 (N_8748,N_8177,N_7926);
xnor U8749 (N_8749,N_8345,N_8128);
xnor U8750 (N_8750,N_7821,N_8002);
nand U8751 (N_8751,N_7847,N_7872);
and U8752 (N_8752,N_8061,N_8265);
nor U8753 (N_8753,N_8048,N_7894);
nor U8754 (N_8754,N_7950,N_8250);
or U8755 (N_8755,N_8166,N_7811);
nor U8756 (N_8756,N_7939,N_8022);
and U8757 (N_8757,N_8191,N_7856);
nand U8758 (N_8758,N_8056,N_8383);
xnor U8759 (N_8759,N_8155,N_8386);
and U8760 (N_8760,N_7842,N_7963);
nor U8761 (N_8761,N_8303,N_8239);
nand U8762 (N_8762,N_7900,N_7942);
nand U8763 (N_8763,N_7867,N_8324);
nor U8764 (N_8764,N_7838,N_8214);
nor U8765 (N_8765,N_8370,N_8390);
nor U8766 (N_8766,N_8001,N_8183);
and U8767 (N_8767,N_8071,N_7954);
nor U8768 (N_8768,N_8219,N_8018);
and U8769 (N_8769,N_8224,N_8099);
and U8770 (N_8770,N_7865,N_8149);
nor U8771 (N_8771,N_8031,N_8387);
and U8772 (N_8772,N_8029,N_7832);
nor U8773 (N_8773,N_7825,N_7993);
and U8774 (N_8774,N_7973,N_8313);
nand U8775 (N_8775,N_8343,N_8303);
or U8776 (N_8776,N_7870,N_7990);
nor U8777 (N_8777,N_8357,N_8230);
nor U8778 (N_8778,N_8091,N_7861);
nand U8779 (N_8779,N_7847,N_8118);
nor U8780 (N_8780,N_8010,N_8259);
nor U8781 (N_8781,N_8222,N_8364);
nand U8782 (N_8782,N_8205,N_8263);
and U8783 (N_8783,N_8317,N_8037);
nor U8784 (N_8784,N_8104,N_7805);
or U8785 (N_8785,N_7939,N_7928);
nor U8786 (N_8786,N_8303,N_8093);
xnor U8787 (N_8787,N_8334,N_8080);
nor U8788 (N_8788,N_8069,N_8010);
and U8789 (N_8789,N_7985,N_7995);
and U8790 (N_8790,N_8219,N_8004);
xor U8791 (N_8791,N_8284,N_8315);
or U8792 (N_8792,N_8129,N_8024);
nand U8793 (N_8793,N_8361,N_8398);
and U8794 (N_8794,N_8066,N_8125);
and U8795 (N_8795,N_8223,N_7896);
nor U8796 (N_8796,N_8002,N_8141);
and U8797 (N_8797,N_8063,N_8058);
nand U8798 (N_8798,N_8119,N_7890);
xnor U8799 (N_8799,N_8389,N_7842);
nor U8800 (N_8800,N_8082,N_8020);
nand U8801 (N_8801,N_8248,N_8220);
or U8802 (N_8802,N_8197,N_8083);
nand U8803 (N_8803,N_7931,N_7991);
nand U8804 (N_8804,N_8302,N_8334);
xor U8805 (N_8805,N_8292,N_8376);
and U8806 (N_8806,N_8236,N_7973);
xnor U8807 (N_8807,N_8007,N_8072);
nand U8808 (N_8808,N_8272,N_7804);
and U8809 (N_8809,N_7943,N_7929);
or U8810 (N_8810,N_8103,N_8237);
and U8811 (N_8811,N_7955,N_8173);
xnor U8812 (N_8812,N_8003,N_8389);
nor U8813 (N_8813,N_8348,N_8129);
or U8814 (N_8814,N_8317,N_8201);
or U8815 (N_8815,N_8390,N_8325);
and U8816 (N_8816,N_8031,N_8321);
or U8817 (N_8817,N_8338,N_8052);
or U8818 (N_8818,N_7905,N_7829);
nand U8819 (N_8819,N_8141,N_7807);
and U8820 (N_8820,N_7935,N_8218);
nor U8821 (N_8821,N_8016,N_8185);
and U8822 (N_8822,N_8020,N_8070);
or U8823 (N_8823,N_7942,N_8129);
and U8824 (N_8824,N_8373,N_8105);
or U8825 (N_8825,N_8081,N_7971);
or U8826 (N_8826,N_7894,N_7857);
and U8827 (N_8827,N_8276,N_7949);
and U8828 (N_8828,N_8127,N_7939);
or U8829 (N_8829,N_8000,N_7845);
and U8830 (N_8830,N_8290,N_7923);
nor U8831 (N_8831,N_7898,N_8329);
nor U8832 (N_8832,N_7959,N_7883);
or U8833 (N_8833,N_7944,N_7958);
xnor U8834 (N_8834,N_8230,N_7915);
nor U8835 (N_8835,N_8345,N_8049);
and U8836 (N_8836,N_7959,N_8260);
nor U8837 (N_8837,N_8070,N_7826);
xnor U8838 (N_8838,N_8204,N_8376);
and U8839 (N_8839,N_7915,N_8152);
nand U8840 (N_8840,N_8367,N_8261);
nor U8841 (N_8841,N_7844,N_7991);
and U8842 (N_8842,N_8385,N_7823);
or U8843 (N_8843,N_8080,N_8343);
nor U8844 (N_8844,N_8088,N_7930);
or U8845 (N_8845,N_7913,N_8253);
nand U8846 (N_8846,N_8168,N_8365);
and U8847 (N_8847,N_7887,N_8312);
and U8848 (N_8848,N_7995,N_7970);
or U8849 (N_8849,N_8223,N_8126);
and U8850 (N_8850,N_8052,N_7878);
nor U8851 (N_8851,N_8374,N_8234);
and U8852 (N_8852,N_8254,N_8043);
and U8853 (N_8853,N_7923,N_8129);
or U8854 (N_8854,N_8333,N_8215);
or U8855 (N_8855,N_7830,N_8214);
or U8856 (N_8856,N_8354,N_8265);
nand U8857 (N_8857,N_7916,N_7893);
xor U8858 (N_8858,N_7814,N_8147);
nand U8859 (N_8859,N_8047,N_7837);
nor U8860 (N_8860,N_7833,N_8145);
nor U8861 (N_8861,N_7992,N_8159);
or U8862 (N_8862,N_8072,N_8180);
nand U8863 (N_8863,N_8065,N_8132);
and U8864 (N_8864,N_7966,N_8223);
nor U8865 (N_8865,N_7918,N_7894);
nor U8866 (N_8866,N_7939,N_8095);
or U8867 (N_8867,N_7841,N_7813);
xnor U8868 (N_8868,N_8250,N_8371);
xnor U8869 (N_8869,N_7891,N_7861);
and U8870 (N_8870,N_7972,N_8223);
nand U8871 (N_8871,N_8021,N_8088);
or U8872 (N_8872,N_8329,N_8159);
xor U8873 (N_8873,N_8248,N_8292);
and U8874 (N_8874,N_7975,N_8149);
nor U8875 (N_8875,N_7915,N_8372);
and U8876 (N_8876,N_8326,N_7853);
nand U8877 (N_8877,N_8231,N_8037);
nand U8878 (N_8878,N_8271,N_8020);
nand U8879 (N_8879,N_7930,N_7880);
or U8880 (N_8880,N_8100,N_8354);
or U8881 (N_8881,N_8354,N_7890);
nor U8882 (N_8882,N_8356,N_8302);
nor U8883 (N_8883,N_8256,N_8212);
nor U8884 (N_8884,N_8251,N_8334);
nor U8885 (N_8885,N_8188,N_7878);
nand U8886 (N_8886,N_8233,N_8269);
or U8887 (N_8887,N_8356,N_8137);
or U8888 (N_8888,N_8148,N_7809);
or U8889 (N_8889,N_8208,N_7925);
nor U8890 (N_8890,N_7816,N_8088);
and U8891 (N_8891,N_7984,N_8138);
and U8892 (N_8892,N_8343,N_8134);
or U8893 (N_8893,N_7961,N_8285);
nor U8894 (N_8894,N_7814,N_8373);
nand U8895 (N_8895,N_7827,N_8055);
and U8896 (N_8896,N_8372,N_7992);
or U8897 (N_8897,N_7936,N_8345);
and U8898 (N_8898,N_8275,N_8166);
and U8899 (N_8899,N_8027,N_7810);
or U8900 (N_8900,N_7989,N_7919);
or U8901 (N_8901,N_8237,N_7876);
nor U8902 (N_8902,N_8125,N_8110);
nor U8903 (N_8903,N_7801,N_7965);
nand U8904 (N_8904,N_8170,N_7929);
xnor U8905 (N_8905,N_8207,N_8115);
and U8906 (N_8906,N_7990,N_8074);
and U8907 (N_8907,N_7801,N_7941);
nor U8908 (N_8908,N_7938,N_7913);
xnor U8909 (N_8909,N_8331,N_8080);
or U8910 (N_8910,N_8066,N_8210);
or U8911 (N_8911,N_8274,N_8306);
nor U8912 (N_8912,N_7970,N_7846);
or U8913 (N_8913,N_7859,N_8331);
nor U8914 (N_8914,N_8029,N_8197);
nand U8915 (N_8915,N_8357,N_8151);
and U8916 (N_8916,N_7950,N_8297);
nand U8917 (N_8917,N_8029,N_7988);
and U8918 (N_8918,N_8196,N_7877);
nor U8919 (N_8919,N_8065,N_7946);
and U8920 (N_8920,N_7813,N_8225);
nor U8921 (N_8921,N_8372,N_8255);
nor U8922 (N_8922,N_8146,N_8255);
nor U8923 (N_8923,N_8158,N_7915);
nor U8924 (N_8924,N_8091,N_7820);
and U8925 (N_8925,N_8062,N_8071);
and U8926 (N_8926,N_8019,N_7849);
nand U8927 (N_8927,N_8239,N_7802);
nand U8928 (N_8928,N_8049,N_8284);
and U8929 (N_8929,N_8361,N_7977);
nand U8930 (N_8930,N_8220,N_7820);
or U8931 (N_8931,N_8050,N_7967);
or U8932 (N_8932,N_8108,N_7946);
nor U8933 (N_8933,N_8154,N_8376);
nor U8934 (N_8934,N_8163,N_8074);
and U8935 (N_8935,N_7960,N_7839);
or U8936 (N_8936,N_8312,N_8265);
or U8937 (N_8937,N_8210,N_8208);
nand U8938 (N_8938,N_8266,N_7821);
or U8939 (N_8939,N_7962,N_7816);
or U8940 (N_8940,N_8236,N_8039);
nor U8941 (N_8941,N_7909,N_8082);
nand U8942 (N_8942,N_8156,N_8176);
nand U8943 (N_8943,N_8104,N_7819);
xor U8944 (N_8944,N_7919,N_7963);
xnor U8945 (N_8945,N_8259,N_8265);
nand U8946 (N_8946,N_8304,N_7937);
nand U8947 (N_8947,N_8204,N_8245);
nor U8948 (N_8948,N_8054,N_7877);
nand U8949 (N_8949,N_7802,N_8131);
and U8950 (N_8950,N_7924,N_8264);
nor U8951 (N_8951,N_8335,N_7994);
nand U8952 (N_8952,N_7944,N_7809);
or U8953 (N_8953,N_7836,N_8104);
nand U8954 (N_8954,N_8340,N_8031);
xnor U8955 (N_8955,N_8279,N_8375);
nor U8956 (N_8956,N_7845,N_8007);
xor U8957 (N_8957,N_8169,N_8178);
nand U8958 (N_8958,N_8302,N_7835);
and U8959 (N_8959,N_7853,N_8314);
or U8960 (N_8960,N_7870,N_8300);
and U8961 (N_8961,N_8168,N_8084);
nor U8962 (N_8962,N_8034,N_8145);
and U8963 (N_8963,N_7927,N_8065);
or U8964 (N_8964,N_7900,N_8389);
xor U8965 (N_8965,N_8239,N_8200);
nand U8966 (N_8966,N_7918,N_7908);
nand U8967 (N_8967,N_8310,N_8334);
nand U8968 (N_8968,N_8312,N_8171);
xnor U8969 (N_8969,N_8210,N_7908);
and U8970 (N_8970,N_8175,N_8134);
or U8971 (N_8971,N_7865,N_7849);
and U8972 (N_8972,N_7994,N_8260);
and U8973 (N_8973,N_7883,N_7848);
and U8974 (N_8974,N_8389,N_7978);
xnor U8975 (N_8975,N_7836,N_7893);
nand U8976 (N_8976,N_7903,N_8062);
nor U8977 (N_8977,N_7952,N_7852);
or U8978 (N_8978,N_8238,N_8199);
nor U8979 (N_8979,N_8321,N_8101);
nor U8980 (N_8980,N_8008,N_8386);
nor U8981 (N_8981,N_7817,N_8301);
and U8982 (N_8982,N_8269,N_8219);
nand U8983 (N_8983,N_8244,N_8331);
and U8984 (N_8984,N_7910,N_8084);
or U8985 (N_8985,N_7894,N_8036);
and U8986 (N_8986,N_8112,N_8175);
nor U8987 (N_8987,N_8246,N_7862);
nand U8988 (N_8988,N_7870,N_7865);
and U8989 (N_8989,N_7980,N_7849);
and U8990 (N_8990,N_8272,N_8177);
nand U8991 (N_8991,N_8307,N_7826);
nor U8992 (N_8992,N_7919,N_8026);
nand U8993 (N_8993,N_8045,N_8172);
and U8994 (N_8994,N_8308,N_8182);
xor U8995 (N_8995,N_8154,N_8245);
or U8996 (N_8996,N_8321,N_8234);
xor U8997 (N_8997,N_8127,N_8217);
or U8998 (N_8998,N_8358,N_8111);
nand U8999 (N_8999,N_8261,N_8191);
nand U9000 (N_9000,N_8697,N_8546);
and U9001 (N_9001,N_8753,N_8643);
xnor U9002 (N_9002,N_8930,N_8843);
and U9003 (N_9003,N_8519,N_8590);
nand U9004 (N_9004,N_8940,N_8598);
or U9005 (N_9005,N_8887,N_8947);
and U9006 (N_9006,N_8589,N_8527);
nor U9007 (N_9007,N_8858,N_8632);
xnor U9008 (N_9008,N_8815,N_8418);
nand U9009 (N_9009,N_8464,N_8477);
or U9010 (N_9010,N_8535,N_8606);
and U9011 (N_9011,N_8439,N_8763);
nor U9012 (N_9012,N_8859,N_8939);
or U9013 (N_9013,N_8718,N_8489);
nand U9014 (N_9014,N_8921,N_8537);
nor U9015 (N_9015,N_8757,N_8716);
nand U9016 (N_9016,N_8918,N_8719);
xnor U9017 (N_9017,N_8827,N_8454);
and U9018 (N_9018,N_8510,N_8877);
and U9019 (N_9019,N_8754,N_8710);
and U9020 (N_9020,N_8514,N_8731);
or U9021 (N_9021,N_8969,N_8695);
nor U9022 (N_9022,N_8430,N_8875);
nand U9023 (N_9023,N_8442,N_8528);
nor U9024 (N_9024,N_8771,N_8401);
or U9025 (N_9025,N_8825,N_8983);
and U9026 (N_9026,N_8652,N_8686);
nand U9027 (N_9027,N_8416,N_8425);
or U9028 (N_9028,N_8903,N_8673);
or U9029 (N_9029,N_8573,N_8547);
nor U9030 (N_9030,N_8961,N_8642);
or U9031 (N_9031,N_8511,N_8582);
and U9032 (N_9032,N_8654,N_8832);
or U9033 (N_9033,N_8491,N_8865);
nor U9034 (N_9034,N_8678,N_8945);
nor U9035 (N_9035,N_8839,N_8826);
and U9036 (N_9036,N_8923,N_8612);
nor U9037 (N_9037,N_8460,N_8506);
nand U9038 (N_9038,N_8737,N_8626);
and U9039 (N_9039,N_8487,N_8524);
and U9040 (N_9040,N_8583,N_8805);
or U9041 (N_9041,N_8772,N_8905);
and U9042 (N_9042,N_8861,N_8882);
and U9043 (N_9043,N_8835,N_8620);
or U9044 (N_9044,N_8931,N_8950);
and U9045 (N_9045,N_8540,N_8848);
or U9046 (N_9046,N_8680,N_8692);
nor U9047 (N_9047,N_8521,N_8989);
nand U9048 (N_9048,N_8787,N_8899);
and U9049 (N_9049,N_8976,N_8978);
nor U9050 (N_9050,N_8896,N_8560);
nor U9051 (N_9051,N_8550,N_8586);
or U9052 (N_9052,N_8480,N_8709);
and U9053 (N_9053,N_8470,N_8972);
nand U9054 (N_9054,N_8912,N_8595);
and U9055 (N_9055,N_8810,N_8580);
or U9056 (N_9056,N_8769,N_8513);
and U9057 (N_9057,N_8981,N_8419);
xnor U9058 (N_9058,N_8414,N_8893);
nand U9059 (N_9059,N_8706,N_8596);
and U9060 (N_9060,N_8760,N_8641);
nor U9061 (N_9061,N_8833,N_8762);
or U9062 (N_9062,N_8744,N_8597);
nand U9063 (N_9063,N_8986,N_8503);
and U9064 (N_9064,N_8587,N_8474);
or U9065 (N_9065,N_8855,N_8942);
or U9066 (N_9066,N_8866,N_8475);
or U9067 (N_9067,N_8886,N_8800);
or U9068 (N_9068,N_8473,N_8929);
nor U9069 (N_9069,N_8911,N_8995);
or U9070 (N_9070,N_8427,N_8496);
nor U9071 (N_9071,N_8651,N_8993);
or U9072 (N_9072,N_8765,N_8990);
or U9073 (N_9073,N_8617,N_8533);
or U9074 (N_9074,N_8438,N_8638);
or U9075 (N_9075,N_8406,N_8846);
or U9076 (N_9076,N_8694,N_8852);
xor U9077 (N_9077,N_8426,N_8463);
or U9078 (N_9078,N_8639,N_8417);
or U9079 (N_9079,N_8630,N_8723);
nand U9080 (N_9080,N_8831,N_8851);
nor U9081 (N_9081,N_8732,N_8532);
nor U9082 (N_9082,N_8946,N_8613);
nor U9083 (N_9083,N_8455,N_8655);
or U9084 (N_9084,N_8538,N_8530);
or U9085 (N_9085,N_8637,N_8705);
or U9086 (N_9086,N_8883,N_8663);
and U9087 (N_9087,N_8818,N_8925);
nand U9088 (N_9088,N_8792,N_8486);
or U9089 (N_9089,N_8975,N_8994);
and U9090 (N_9090,N_8581,N_8555);
nand U9091 (N_9091,N_8724,N_8715);
or U9092 (N_9092,N_8508,N_8447);
xor U9093 (N_9093,N_8752,N_8435);
or U9094 (N_9094,N_8433,N_8421);
nand U9095 (N_9095,N_8897,N_8434);
nor U9096 (N_9096,N_8681,N_8482);
or U9097 (N_9097,N_8864,N_8730);
and U9098 (N_9098,N_8400,N_8954);
nor U9099 (N_9099,N_8955,N_8944);
nor U9100 (N_9100,N_8774,N_8777);
or U9101 (N_9101,N_8666,N_8713);
nor U9102 (N_9102,N_8539,N_8922);
xor U9103 (N_9103,N_8608,N_8572);
or U9104 (N_9104,N_8614,N_8646);
and U9105 (N_9105,N_8756,N_8634);
nand U9106 (N_9106,N_8982,N_8959);
nand U9107 (N_9107,N_8523,N_8687);
xnor U9108 (N_9108,N_8428,N_8938);
and U9109 (N_9109,N_8668,N_8962);
nor U9110 (N_9110,N_8570,N_8968);
nor U9111 (N_9111,N_8602,N_8577);
nor U9112 (N_9112,N_8704,N_8431);
nor U9113 (N_9113,N_8682,N_8664);
nor U9114 (N_9114,N_8812,N_8786);
or U9115 (N_9115,N_8776,N_8952);
nand U9116 (N_9116,N_8564,N_8770);
and U9117 (N_9117,N_8522,N_8661);
nor U9118 (N_9118,N_8780,N_8472);
and U9119 (N_9119,N_8747,N_8804);
nor U9120 (N_9120,N_8735,N_8880);
and U9121 (N_9121,N_8948,N_8917);
nor U9122 (N_9122,N_8838,N_8551);
nor U9123 (N_9123,N_8902,N_8504);
and U9124 (N_9124,N_8567,N_8534);
and U9125 (N_9125,N_8565,N_8868);
nor U9126 (N_9126,N_8621,N_8913);
nor U9127 (N_9127,N_8543,N_8649);
or U9128 (N_9128,N_8980,N_8520);
and U9129 (N_9129,N_8615,N_8958);
xnor U9130 (N_9130,N_8984,N_8928);
xor U9131 (N_9131,N_8801,N_8793);
or U9132 (N_9132,N_8700,N_8915);
nor U9133 (N_9133,N_8701,N_8802);
nor U9134 (N_9134,N_8645,N_8484);
and U9135 (N_9135,N_8488,N_8884);
nor U9136 (N_9136,N_8548,N_8808);
or U9137 (N_9137,N_8610,N_8854);
or U9138 (N_9138,N_8919,N_8726);
xnor U9139 (N_9139,N_8479,N_8750);
or U9140 (N_9140,N_8494,N_8782);
or U9141 (N_9141,N_8767,N_8594);
nor U9142 (N_9142,N_8736,N_8690);
or U9143 (N_9143,N_8790,N_8725);
nand U9144 (N_9144,N_8499,N_8721);
or U9145 (N_9145,N_8844,N_8562);
nand U9146 (N_9146,N_8451,N_8809);
and U9147 (N_9147,N_8557,N_8653);
and U9148 (N_9148,N_8525,N_8849);
and U9149 (N_9149,N_8405,N_8888);
nand U9150 (N_9150,N_8881,N_8457);
nor U9151 (N_9151,N_8691,N_8600);
nor U9152 (N_9152,N_8604,N_8609);
nor U9153 (N_9153,N_8449,N_8498);
xnor U9154 (N_9154,N_8941,N_8437);
nand U9155 (N_9155,N_8907,N_8552);
nand U9156 (N_9156,N_8906,N_8773);
nand U9157 (N_9157,N_8640,N_8734);
nor U9158 (N_9158,N_8998,N_8627);
xor U9159 (N_9159,N_8461,N_8956);
and U9160 (N_9160,N_8837,N_8970);
and U9161 (N_9161,N_8670,N_8512);
or U9162 (N_9162,N_8977,N_8828);
or U9163 (N_9163,N_8830,N_8728);
nor U9164 (N_9164,N_8748,N_8836);
nand U9165 (N_9165,N_8824,N_8797);
xnor U9166 (N_9166,N_8440,N_8926);
and U9167 (N_9167,N_8829,N_8967);
and U9168 (N_9168,N_8795,N_8683);
or U9169 (N_9169,N_8711,N_8415);
nor U9170 (N_9170,N_8660,N_8739);
nor U9171 (N_9171,N_8650,N_8784);
nor U9172 (N_9172,N_8820,N_8554);
and U9173 (N_9173,N_8714,N_8500);
nor U9174 (N_9174,N_8814,N_8413);
nor U9175 (N_9175,N_8624,N_8591);
nand U9176 (N_9176,N_8569,N_8526);
nand U9177 (N_9177,N_8529,N_8404);
or U9178 (N_9178,N_8746,N_8799);
xnor U9179 (N_9179,N_8493,N_8789);
and U9180 (N_9180,N_8932,N_8698);
and U9181 (N_9181,N_8676,N_8974);
and U9182 (N_9182,N_8885,N_8625);
and U9183 (N_9183,N_8823,N_8631);
or U9184 (N_9184,N_8965,N_8432);
xnor U9185 (N_9185,N_8616,N_8966);
and U9186 (N_9186,N_8476,N_8857);
nand U9187 (N_9187,N_8758,N_8408);
or U9188 (N_9188,N_8991,N_8515);
nor U9189 (N_9189,N_8850,N_8891);
nand U9190 (N_9190,N_8764,N_8545);
nand U9191 (N_9191,N_8657,N_8775);
nor U9192 (N_9192,N_8894,N_8662);
nor U9193 (N_9193,N_8712,N_8807);
and U9194 (N_9194,N_8509,N_8901);
and U9195 (N_9195,N_8916,N_8622);
nor U9196 (N_9196,N_8563,N_8443);
nor U9197 (N_9197,N_8648,N_8465);
and U9198 (N_9198,N_8908,N_8481);
and U9199 (N_9199,N_8536,N_8490);
and U9200 (N_9200,N_8949,N_8819);
xor U9201 (N_9201,N_8665,N_8909);
nand U9202 (N_9202,N_8768,N_8935);
nor U9203 (N_9203,N_8456,N_8483);
or U9204 (N_9204,N_8953,N_8679);
nand U9205 (N_9205,N_8834,N_8497);
nor U9206 (N_9206,N_8559,N_8997);
nor U9207 (N_9207,N_8707,N_8856);
nand U9208 (N_9208,N_8862,N_8755);
nor U9209 (N_9209,N_8517,N_8671);
nand U9210 (N_9210,N_8816,N_8717);
nand U9211 (N_9211,N_8633,N_8727);
nand U9212 (N_9212,N_8677,N_8878);
and U9213 (N_9213,N_8605,N_8684);
and U9214 (N_9214,N_8822,N_8412);
nand U9215 (N_9215,N_8599,N_8749);
or U9216 (N_9216,N_8813,N_8936);
nor U9217 (N_9217,N_8492,N_8448);
and U9218 (N_9218,N_8429,N_8674);
xnor U9219 (N_9219,N_8853,N_8996);
and U9220 (N_9220,N_8458,N_8672);
nand U9221 (N_9221,N_8879,N_8870);
and U9222 (N_9222,N_8636,N_8895);
xor U9223 (N_9223,N_8542,N_8601);
nor U9224 (N_9224,N_8867,N_8863);
nand U9225 (N_9225,N_8992,N_8933);
nor U9226 (N_9226,N_8574,N_8740);
xnor U9227 (N_9227,N_8794,N_8585);
or U9228 (N_9228,N_8960,N_8607);
or U9229 (N_9229,N_8871,N_8424);
nand U9230 (N_9230,N_8495,N_8741);
or U9231 (N_9231,N_8628,N_8688);
and U9232 (N_9232,N_8811,N_8779);
nand U9233 (N_9233,N_8708,N_8578);
or U9234 (N_9234,N_8409,N_8873);
and U9235 (N_9235,N_8453,N_8531);
nor U9236 (N_9236,N_8423,N_8898);
nand U9237 (N_9237,N_8445,N_8450);
or U9238 (N_9238,N_8619,N_8876);
nor U9239 (N_9239,N_8841,N_8842);
or U9240 (N_9240,N_8566,N_8549);
xnor U9241 (N_9241,N_8611,N_8910);
nand U9242 (N_9242,N_8576,N_8788);
or U9243 (N_9243,N_8647,N_8702);
nor U9244 (N_9244,N_8759,N_8593);
or U9245 (N_9245,N_8603,N_8592);
nor U9246 (N_9246,N_8507,N_8927);
nand U9247 (N_9247,N_8934,N_8937);
or U9248 (N_9248,N_8973,N_8685);
nor U9249 (N_9249,N_8943,N_8892);
or U9250 (N_9250,N_8987,N_8544);
nor U9251 (N_9251,N_8778,N_8469);
and U9252 (N_9252,N_8817,N_8644);
and U9253 (N_9253,N_8971,N_8840);
and U9254 (N_9254,N_8785,N_8407);
nor U9255 (N_9255,N_8845,N_8667);
nand U9256 (N_9256,N_8452,N_8964);
and U9257 (N_9257,N_8618,N_8729);
and U9258 (N_9258,N_8422,N_8890);
and U9259 (N_9259,N_8791,N_8410);
xnor U9260 (N_9260,N_8669,N_8518);
xor U9261 (N_9261,N_8485,N_8459);
and U9262 (N_9262,N_8571,N_8920);
nand U9263 (N_9263,N_8558,N_8588);
nand U9264 (N_9264,N_8999,N_8847);
nand U9265 (N_9265,N_8516,N_8462);
nand U9266 (N_9266,N_8502,N_8411);
or U9267 (N_9267,N_8796,N_8444);
and U9268 (N_9268,N_8556,N_8436);
and U9269 (N_9269,N_8745,N_8806);
nand U9270 (N_9270,N_8468,N_8783);
xnor U9271 (N_9271,N_8402,N_8446);
nor U9272 (N_9272,N_8781,N_8798);
nand U9273 (N_9273,N_8696,N_8579);
and U9274 (N_9274,N_8979,N_8957);
nor U9275 (N_9275,N_8659,N_8693);
or U9276 (N_9276,N_8951,N_8699);
nand U9277 (N_9277,N_8743,N_8985);
xnor U9278 (N_9278,N_8869,N_8505);
nor U9279 (N_9279,N_8568,N_8501);
and U9280 (N_9280,N_8722,N_8467);
nor U9281 (N_9281,N_8874,N_8924);
nand U9282 (N_9282,N_8860,N_8629);
nor U9283 (N_9283,N_8403,N_8742);
or U9284 (N_9284,N_8541,N_8720);
and U9285 (N_9285,N_8420,N_8904);
nand U9286 (N_9286,N_8623,N_8689);
or U9287 (N_9287,N_8441,N_8821);
nand U9288 (N_9288,N_8963,N_8988);
and U9289 (N_9289,N_8635,N_8584);
nor U9290 (N_9290,N_8761,N_8561);
and U9291 (N_9291,N_8889,N_8803);
and U9292 (N_9292,N_8751,N_8766);
xnor U9293 (N_9293,N_8675,N_8738);
nor U9294 (N_9294,N_8914,N_8733);
nor U9295 (N_9295,N_8656,N_8703);
or U9296 (N_9296,N_8478,N_8553);
nand U9297 (N_9297,N_8466,N_8575);
nor U9298 (N_9298,N_8900,N_8872);
and U9299 (N_9299,N_8471,N_8658);
nor U9300 (N_9300,N_8629,N_8822);
and U9301 (N_9301,N_8711,N_8954);
nand U9302 (N_9302,N_8506,N_8864);
or U9303 (N_9303,N_8600,N_8668);
nor U9304 (N_9304,N_8899,N_8548);
xnor U9305 (N_9305,N_8528,N_8456);
and U9306 (N_9306,N_8718,N_8479);
and U9307 (N_9307,N_8598,N_8681);
nand U9308 (N_9308,N_8989,N_8919);
and U9309 (N_9309,N_8409,N_8832);
and U9310 (N_9310,N_8950,N_8596);
nand U9311 (N_9311,N_8803,N_8962);
and U9312 (N_9312,N_8525,N_8965);
nor U9313 (N_9313,N_8809,N_8581);
nor U9314 (N_9314,N_8502,N_8849);
and U9315 (N_9315,N_8964,N_8693);
nor U9316 (N_9316,N_8578,N_8445);
nor U9317 (N_9317,N_8889,N_8504);
and U9318 (N_9318,N_8909,N_8425);
xnor U9319 (N_9319,N_8837,N_8569);
nor U9320 (N_9320,N_8848,N_8593);
nand U9321 (N_9321,N_8966,N_8543);
nand U9322 (N_9322,N_8909,N_8875);
nand U9323 (N_9323,N_8511,N_8541);
nand U9324 (N_9324,N_8602,N_8540);
nor U9325 (N_9325,N_8511,N_8401);
or U9326 (N_9326,N_8951,N_8453);
nor U9327 (N_9327,N_8450,N_8945);
nor U9328 (N_9328,N_8412,N_8913);
and U9329 (N_9329,N_8490,N_8603);
or U9330 (N_9330,N_8579,N_8623);
nor U9331 (N_9331,N_8588,N_8765);
nand U9332 (N_9332,N_8635,N_8486);
and U9333 (N_9333,N_8478,N_8782);
nor U9334 (N_9334,N_8559,N_8409);
nor U9335 (N_9335,N_8480,N_8989);
and U9336 (N_9336,N_8882,N_8627);
and U9337 (N_9337,N_8407,N_8792);
or U9338 (N_9338,N_8863,N_8417);
nor U9339 (N_9339,N_8811,N_8568);
nand U9340 (N_9340,N_8917,N_8647);
xnor U9341 (N_9341,N_8567,N_8846);
or U9342 (N_9342,N_8604,N_8799);
nand U9343 (N_9343,N_8837,N_8921);
nand U9344 (N_9344,N_8646,N_8846);
nand U9345 (N_9345,N_8654,N_8976);
nor U9346 (N_9346,N_8874,N_8645);
and U9347 (N_9347,N_8475,N_8998);
nor U9348 (N_9348,N_8526,N_8920);
xnor U9349 (N_9349,N_8659,N_8910);
nor U9350 (N_9350,N_8594,N_8559);
nand U9351 (N_9351,N_8883,N_8514);
and U9352 (N_9352,N_8402,N_8729);
or U9353 (N_9353,N_8629,N_8866);
nor U9354 (N_9354,N_8552,N_8850);
or U9355 (N_9355,N_8615,N_8734);
nand U9356 (N_9356,N_8916,N_8667);
or U9357 (N_9357,N_8452,N_8588);
or U9358 (N_9358,N_8823,N_8662);
xnor U9359 (N_9359,N_8437,N_8922);
and U9360 (N_9360,N_8720,N_8973);
or U9361 (N_9361,N_8933,N_8623);
or U9362 (N_9362,N_8736,N_8870);
and U9363 (N_9363,N_8918,N_8583);
and U9364 (N_9364,N_8777,N_8971);
and U9365 (N_9365,N_8908,N_8806);
and U9366 (N_9366,N_8436,N_8552);
and U9367 (N_9367,N_8805,N_8886);
nand U9368 (N_9368,N_8934,N_8408);
nand U9369 (N_9369,N_8902,N_8814);
nand U9370 (N_9370,N_8456,N_8672);
nor U9371 (N_9371,N_8586,N_8861);
nor U9372 (N_9372,N_8508,N_8763);
nor U9373 (N_9373,N_8995,N_8822);
nor U9374 (N_9374,N_8940,N_8941);
nor U9375 (N_9375,N_8559,N_8716);
or U9376 (N_9376,N_8544,N_8492);
nand U9377 (N_9377,N_8458,N_8950);
nor U9378 (N_9378,N_8847,N_8785);
nand U9379 (N_9379,N_8424,N_8720);
and U9380 (N_9380,N_8994,N_8585);
and U9381 (N_9381,N_8886,N_8591);
or U9382 (N_9382,N_8479,N_8414);
xnor U9383 (N_9383,N_8988,N_8428);
and U9384 (N_9384,N_8989,N_8485);
and U9385 (N_9385,N_8743,N_8516);
nor U9386 (N_9386,N_8888,N_8506);
or U9387 (N_9387,N_8763,N_8810);
nor U9388 (N_9388,N_8765,N_8511);
and U9389 (N_9389,N_8990,N_8823);
xor U9390 (N_9390,N_8729,N_8639);
xnor U9391 (N_9391,N_8901,N_8729);
and U9392 (N_9392,N_8876,N_8539);
nor U9393 (N_9393,N_8540,N_8912);
and U9394 (N_9394,N_8568,N_8976);
and U9395 (N_9395,N_8761,N_8679);
nor U9396 (N_9396,N_8521,N_8778);
nor U9397 (N_9397,N_8861,N_8435);
or U9398 (N_9398,N_8929,N_8549);
or U9399 (N_9399,N_8680,N_8868);
and U9400 (N_9400,N_8896,N_8412);
and U9401 (N_9401,N_8610,N_8566);
xnor U9402 (N_9402,N_8432,N_8561);
or U9403 (N_9403,N_8762,N_8479);
and U9404 (N_9404,N_8775,N_8922);
and U9405 (N_9405,N_8636,N_8473);
xnor U9406 (N_9406,N_8602,N_8862);
xnor U9407 (N_9407,N_8613,N_8543);
and U9408 (N_9408,N_8492,N_8659);
and U9409 (N_9409,N_8553,N_8459);
and U9410 (N_9410,N_8538,N_8616);
nor U9411 (N_9411,N_8792,N_8898);
nor U9412 (N_9412,N_8441,N_8928);
xnor U9413 (N_9413,N_8733,N_8412);
or U9414 (N_9414,N_8455,N_8636);
nand U9415 (N_9415,N_8730,N_8834);
nor U9416 (N_9416,N_8742,N_8560);
nand U9417 (N_9417,N_8855,N_8810);
xor U9418 (N_9418,N_8470,N_8683);
nand U9419 (N_9419,N_8999,N_8595);
nand U9420 (N_9420,N_8638,N_8775);
xnor U9421 (N_9421,N_8665,N_8513);
nand U9422 (N_9422,N_8413,N_8960);
or U9423 (N_9423,N_8582,N_8402);
or U9424 (N_9424,N_8817,N_8871);
nor U9425 (N_9425,N_8781,N_8776);
or U9426 (N_9426,N_8928,N_8708);
or U9427 (N_9427,N_8761,N_8946);
or U9428 (N_9428,N_8698,N_8835);
xor U9429 (N_9429,N_8944,N_8785);
or U9430 (N_9430,N_8847,N_8586);
and U9431 (N_9431,N_8837,N_8457);
and U9432 (N_9432,N_8483,N_8742);
or U9433 (N_9433,N_8737,N_8576);
or U9434 (N_9434,N_8683,N_8516);
xor U9435 (N_9435,N_8645,N_8754);
and U9436 (N_9436,N_8440,N_8728);
or U9437 (N_9437,N_8516,N_8693);
nor U9438 (N_9438,N_8718,N_8508);
and U9439 (N_9439,N_8581,N_8982);
or U9440 (N_9440,N_8526,N_8944);
and U9441 (N_9441,N_8754,N_8558);
or U9442 (N_9442,N_8977,N_8712);
nor U9443 (N_9443,N_8609,N_8981);
or U9444 (N_9444,N_8796,N_8759);
nor U9445 (N_9445,N_8811,N_8754);
and U9446 (N_9446,N_8826,N_8907);
and U9447 (N_9447,N_8832,N_8550);
and U9448 (N_9448,N_8692,N_8830);
or U9449 (N_9449,N_8552,N_8764);
or U9450 (N_9450,N_8938,N_8846);
nand U9451 (N_9451,N_8688,N_8508);
nand U9452 (N_9452,N_8412,N_8973);
nand U9453 (N_9453,N_8641,N_8970);
or U9454 (N_9454,N_8888,N_8849);
or U9455 (N_9455,N_8824,N_8821);
xor U9456 (N_9456,N_8547,N_8793);
nand U9457 (N_9457,N_8575,N_8957);
xor U9458 (N_9458,N_8976,N_8555);
nand U9459 (N_9459,N_8525,N_8858);
or U9460 (N_9460,N_8992,N_8846);
and U9461 (N_9461,N_8748,N_8405);
or U9462 (N_9462,N_8444,N_8431);
nor U9463 (N_9463,N_8552,N_8628);
or U9464 (N_9464,N_8551,N_8530);
xnor U9465 (N_9465,N_8431,N_8536);
nor U9466 (N_9466,N_8952,N_8412);
and U9467 (N_9467,N_8732,N_8783);
nand U9468 (N_9468,N_8746,N_8865);
nor U9469 (N_9469,N_8721,N_8915);
or U9470 (N_9470,N_8941,N_8505);
nand U9471 (N_9471,N_8516,N_8763);
or U9472 (N_9472,N_8827,N_8848);
nor U9473 (N_9473,N_8592,N_8593);
nand U9474 (N_9474,N_8599,N_8670);
nor U9475 (N_9475,N_8896,N_8953);
or U9476 (N_9476,N_8988,N_8873);
xor U9477 (N_9477,N_8660,N_8776);
and U9478 (N_9478,N_8794,N_8420);
and U9479 (N_9479,N_8648,N_8665);
or U9480 (N_9480,N_8568,N_8818);
nor U9481 (N_9481,N_8559,N_8616);
nor U9482 (N_9482,N_8608,N_8410);
nor U9483 (N_9483,N_8575,N_8441);
or U9484 (N_9484,N_8424,N_8762);
or U9485 (N_9485,N_8489,N_8734);
and U9486 (N_9486,N_8796,N_8902);
nor U9487 (N_9487,N_8730,N_8930);
or U9488 (N_9488,N_8611,N_8469);
xor U9489 (N_9489,N_8494,N_8515);
and U9490 (N_9490,N_8681,N_8845);
and U9491 (N_9491,N_8917,N_8924);
and U9492 (N_9492,N_8814,N_8883);
nor U9493 (N_9493,N_8781,N_8983);
nand U9494 (N_9494,N_8668,N_8785);
nor U9495 (N_9495,N_8455,N_8973);
nand U9496 (N_9496,N_8764,N_8535);
nand U9497 (N_9497,N_8816,N_8954);
nand U9498 (N_9498,N_8433,N_8893);
nand U9499 (N_9499,N_8988,N_8439);
or U9500 (N_9500,N_8790,N_8540);
nand U9501 (N_9501,N_8419,N_8476);
or U9502 (N_9502,N_8596,N_8754);
and U9503 (N_9503,N_8664,N_8769);
and U9504 (N_9504,N_8536,N_8844);
or U9505 (N_9505,N_8613,N_8671);
and U9506 (N_9506,N_8754,N_8430);
or U9507 (N_9507,N_8583,N_8772);
and U9508 (N_9508,N_8699,N_8882);
nand U9509 (N_9509,N_8907,N_8919);
nor U9510 (N_9510,N_8679,N_8884);
nand U9511 (N_9511,N_8492,N_8440);
nor U9512 (N_9512,N_8477,N_8778);
or U9513 (N_9513,N_8823,N_8440);
or U9514 (N_9514,N_8714,N_8520);
nor U9515 (N_9515,N_8516,N_8785);
nor U9516 (N_9516,N_8891,N_8806);
nand U9517 (N_9517,N_8743,N_8541);
xor U9518 (N_9518,N_8587,N_8432);
or U9519 (N_9519,N_8628,N_8461);
and U9520 (N_9520,N_8677,N_8819);
and U9521 (N_9521,N_8955,N_8929);
or U9522 (N_9522,N_8961,N_8673);
and U9523 (N_9523,N_8442,N_8978);
xnor U9524 (N_9524,N_8995,N_8906);
or U9525 (N_9525,N_8694,N_8569);
xnor U9526 (N_9526,N_8731,N_8618);
nor U9527 (N_9527,N_8765,N_8811);
nor U9528 (N_9528,N_8403,N_8561);
or U9529 (N_9529,N_8429,N_8473);
or U9530 (N_9530,N_8882,N_8704);
xor U9531 (N_9531,N_8518,N_8618);
or U9532 (N_9532,N_8447,N_8706);
and U9533 (N_9533,N_8926,N_8981);
and U9534 (N_9534,N_8615,N_8682);
or U9535 (N_9535,N_8637,N_8526);
nor U9536 (N_9536,N_8491,N_8686);
and U9537 (N_9537,N_8752,N_8658);
and U9538 (N_9538,N_8745,N_8918);
or U9539 (N_9539,N_8429,N_8990);
xor U9540 (N_9540,N_8852,N_8879);
nor U9541 (N_9541,N_8451,N_8755);
or U9542 (N_9542,N_8743,N_8657);
and U9543 (N_9543,N_8587,N_8684);
nand U9544 (N_9544,N_8616,N_8732);
nand U9545 (N_9545,N_8602,N_8459);
and U9546 (N_9546,N_8681,N_8705);
and U9547 (N_9547,N_8900,N_8743);
and U9548 (N_9548,N_8899,N_8421);
or U9549 (N_9549,N_8492,N_8496);
nand U9550 (N_9550,N_8885,N_8432);
or U9551 (N_9551,N_8702,N_8492);
or U9552 (N_9552,N_8748,N_8766);
and U9553 (N_9553,N_8598,N_8454);
nand U9554 (N_9554,N_8987,N_8656);
or U9555 (N_9555,N_8440,N_8739);
nand U9556 (N_9556,N_8464,N_8753);
nand U9557 (N_9557,N_8867,N_8571);
or U9558 (N_9558,N_8500,N_8523);
nand U9559 (N_9559,N_8459,N_8518);
nand U9560 (N_9560,N_8773,N_8952);
xnor U9561 (N_9561,N_8649,N_8681);
xor U9562 (N_9562,N_8526,N_8524);
xnor U9563 (N_9563,N_8846,N_8597);
nand U9564 (N_9564,N_8778,N_8897);
xnor U9565 (N_9565,N_8523,N_8670);
nor U9566 (N_9566,N_8464,N_8597);
nor U9567 (N_9567,N_8887,N_8860);
nand U9568 (N_9568,N_8605,N_8878);
nand U9569 (N_9569,N_8717,N_8754);
nor U9570 (N_9570,N_8681,N_8535);
or U9571 (N_9571,N_8681,N_8732);
or U9572 (N_9572,N_8994,N_8539);
nand U9573 (N_9573,N_8952,N_8562);
or U9574 (N_9574,N_8656,N_8940);
or U9575 (N_9575,N_8920,N_8777);
nor U9576 (N_9576,N_8726,N_8924);
xnor U9577 (N_9577,N_8581,N_8835);
nand U9578 (N_9578,N_8494,N_8978);
and U9579 (N_9579,N_8830,N_8734);
or U9580 (N_9580,N_8648,N_8964);
nor U9581 (N_9581,N_8889,N_8706);
xor U9582 (N_9582,N_8799,N_8942);
nor U9583 (N_9583,N_8547,N_8892);
and U9584 (N_9584,N_8699,N_8420);
xor U9585 (N_9585,N_8765,N_8973);
and U9586 (N_9586,N_8463,N_8500);
nor U9587 (N_9587,N_8996,N_8663);
or U9588 (N_9588,N_8491,N_8528);
and U9589 (N_9589,N_8611,N_8766);
nand U9590 (N_9590,N_8429,N_8724);
nand U9591 (N_9591,N_8884,N_8971);
and U9592 (N_9592,N_8879,N_8698);
and U9593 (N_9593,N_8528,N_8650);
nor U9594 (N_9594,N_8590,N_8622);
nor U9595 (N_9595,N_8925,N_8776);
nand U9596 (N_9596,N_8710,N_8556);
or U9597 (N_9597,N_8527,N_8721);
and U9598 (N_9598,N_8932,N_8852);
xnor U9599 (N_9599,N_8825,N_8732);
and U9600 (N_9600,N_9036,N_9104);
nor U9601 (N_9601,N_9155,N_9367);
xnor U9602 (N_9602,N_9166,N_9421);
and U9603 (N_9603,N_9030,N_9248);
and U9604 (N_9604,N_9083,N_9056);
nand U9605 (N_9605,N_9289,N_9029);
nor U9606 (N_9606,N_9346,N_9426);
nand U9607 (N_9607,N_9245,N_9496);
or U9608 (N_9608,N_9588,N_9106);
or U9609 (N_9609,N_9471,N_9159);
nor U9610 (N_9610,N_9061,N_9050);
or U9611 (N_9611,N_9534,N_9559);
xnor U9612 (N_9612,N_9208,N_9413);
and U9613 (N_9613,N_9277,N_9086);
nor U9614 (N_9614,N_9291,N_9423);
nor U9615 (N_9615,N_9101,N_9156);
nor U9616 (N_9616,N_9154,N_9254);
xnor U9617 (N_9617,N_9008,N_9121);
nor U9618 (N_9618,N_9337,N_9284);
nor U9619 (N_9619,N_9480,N_9206);
nand U9620 (N_9620,N_9386,N_9409);
or U9621 (N_9621,N_9529,N_9225);
nor U9622 (N_9622,N_9515,N_9473);
nand U9623 (N_9623,N_9552,N_9280);
or U9624 (N_9624,N_9356,N_9385);
or U9625 (N_9625,N_9241,N_9115);
nand U9626 (N_9626,N_9293,N_9103);
nor U9627 (N_9627,N_9308,N_9594);
or U9628 (N_9628,N_9422,N_9541);
xnor U9629 (N_9629,N_9412,N_9143);
nand U9630 (N_9630,N_9249,N_9545);
xor U9631 (N_9631,N_9393,N_9077);
or U9632 (N_9632,N_9438,N_9466);
or U9633 (N_9633,N_9485,N_9417);
nand U9634 (N_9634,N_9449,N_9040);
or U9635 (N_9635,N_9137,N_9052);
nand U9636 (N_9636,N_9316,N_9470);
nor U9637 (N_9637,N_9467,N_9437);
nand U9638 (N_9638,N_9502,N_9020);
or U9639 (N_9639,N_9445,N_9063);
xor U9640 (N_9640,N_9345,N_9178);
nand U9641 (N_9641,N_9114,N_9370);
and U9642 (N_9642,N_9318,N_9003);
and U9643 (N_9643,N_9105,N_9142);
nor U9644 (N_9644,N_9011,N_9398);
or U9645 (N_9645,N_9285,N_9487);
and U9646 (N_9646,N_9082,N_9573);
or U9647 (N_9647,N_9574,N_9332);
and U9648 (N_9648,N_9296,N_9294);
nand U9649 (N_9649,N_9149,N_9129);
nor U9650 (N_9650,N_9022,N_9381);
nor U9651 (N_9651,N_9257,N_9322);
or U9652 (N_9652,N_9012,N_9581);
nand U9653 (N_9653,N_9298,N_9251);
xor U9654 (N_9654,N_9392,N_9582);
nand U9655 (N_9655,N_9435,N_9067);
nor U9656 (N_9656,N_9055,N_9317);
nor U9657 (N_9657,N_9116,N_9465);
or U9658 (N_9658,N_9150,N_9428);
xnor U9659 (N_9659,N_9474,N_9505);
nand U9660 (N_9660,N_9202,N_9094);
and U9661 (N_9661,N_9450,N_9233);
or U9662 (N_9662,N_9580,N_9136);
xor U9663 (N_9663,N_9200,N_9507);
or U9664 (N_9664,N_9306,N_9263);
and U9665 (N_9665,N_9522,N_9407);
nor U9666 (N_9666,N_9272,N_9042);
nand U9667 (N_9667,N_9152,N_9181);
and U9668 (N_9668,N_9504,N_9535);
xor U9669 (N_9669,N_9509,N_9433);
or U9670 (N_9670,N_9087,N_9369);
nor U9671 (N_9671,N_9388,N_9425);
nand U9672 (N_9672,N_9468,N_9560);
nor U9673 (N_9673,N_9039,N_9447);
nand U9674 (N_9674,N_9000,N_9547);
and U9675 (N_9675,N_9274,N_9376);
or U9676 (N_9676,N_9500,N_9219);
nand U9677 (N_9677,N_9402,N_9429);
nor U9678 (N_9678,N_9344,N_9002);
and U9679 (N_9679,N_9355,N_9451);
nor U9680 (N_9680,N_9244,N_9589);
and U9681 (N_9681,N_9228,N_9472);
and U9682 (N_9682,N_9045,N_9278);
nand U9683 (N_9683,N_9389,N_9273);
nand U9684 (N_9684,N_9328,N_9361);
or U9685 (N_9685,N_9239,N_9518);
or U9686 (N_9686,N_9536,N_9238);
nand U9687 (N_9687,N_9310,N_9096);
or U9688 (N_9688,N_9569,N_9215);
or U9689 (N_9689,N_9434,N_9302);
and U9690 (N_9690,N_9524,N_9259);
nand U9691 (N_9691,N_9183,N_9243);
nor U9692 (N_9692,N_9368,N_9198);
nor U9693 (N_9693,N_9453,N_9312);
nand U9694 (N_9694,N_9210,N_9269);
nand U9695 (N_9695,N_9304,N_9439);
and U9696 (N_9696,N_9349,N_9194);
or U9697 (N_9697,N_9598,N_9410);
nor U9698 (N_9698,N_9532,N_9148);
or U9699 (N_9699,N_9135,N_9138);
nand U9700 (N_9700,N_9575,N_9576);
or U9701 (N_9701,N_9120,N_9572);
nand U9702 (N_9702,N_9197,N_9174);
or U9703 (N_9703,N_9224,N_9384);
and U9704 (N_9704,N_9054,N_9549);
nand U9705 (N_9705,N_9169,N_9283);
nand U9706 (N_9706,N_9373,N_9246);
nand U9707 (N_9707,N_9334,N_9131);
nand U9708 (N_9708,N_9360,N_9134);
nor U9709 (N_9709,N_9424,N_9184);
nand U9710 (N_9710,N_9185,N_9146);
and U9711 (N_9711,N_9544,N_9226);
nor U9712 (N_9712,N_9590,N_9320);
or U9713 (N_9713,N_9001,N_9191);
or U9714 (N_9714,N_9462,N_9481);
or U9715 (N_9715,N_9394,N_9578);
nor U9716 (N_9716,N_9330,N_9141);
nand U9717 (N_9717,N_9080,N_9062);
and U9718 (N_9718,N_9007,N_9498);
or U9719 (N_9719,N_9119,N_9160);
or U9720 (N_9720,N_9300,N_9523);
or U9721 (N_9721,N_9546,N_9187);
or U9722 (N_9722,N_9309,N_9315);
or U9723 (N_9723,N_9483,N_9041);
nor U9724 (N_9724,N_9161,N_9072);
and U9725 (N_9725,N_9190,N_9555);
or U9726 (N_9726,N_9400,N_9526);
nor U9727 (N_9727,N_9478,N_9108);
nand U9728 (N_9728,N_9223,N_9034);
and U9729 (N_9729,N_9265,N_9493);
nand U9730 (N_9730,N_9299,N_9199);
nor U9731 (N_9731,N_9324,N_9495);
nand U9732 (N_9732,N_9548,N_9490);
nand U9733 (N_9733,N_9222,N_9021);
or U9734 (N_9734,N_9554,N_9557);
nand U9735 (N_9735,N_9416,N_9046);
and U9736 (N_9736,N_9357,N_9538);
nand U9737 (N_9737,N_9093,N_9097);
or U9738 (N_9738,N_9209,N_9033);
nand U9739 (N_9739,N_9562,N_9207);
nor U9740 (N_9740,N_9095,N_9023);
nor U9741 (N_9741,N_9365,N_9252);
nor U9742 (N_9742,N_9511,N_9015);
or U9743 (N_9743,N_9024,N_9377);
nand U9744 (N_9744,N_9517,N_9031);
nor U9745 (N_9745,N_9347,N_9125);
nor U9746 (N_9746,N_9459,N_9537);
and U9747 (N_9747,N_9372,N_9139);
and U9748 (N_9748,N_9004,N_9596);
and U9749 (N_9749,N_9270,N_9411);
and U9750 (N_9750,N_9297,N_9469);
nand U9751 (N_9751,N_9338,N_9446);
or U9752 (N_9752,N_9235,N_9510);
or U9753 (N_9753,N_9068,N_9343);
and U9754 (N_9754,N_9436,N_9242);
and U9755 (N_9755,N_9455,N_9162);
nand U9756 (N_9756,N_9196,N_9216);
and U9757 (N_9757,N_9076,N_9336);
and U9758 (N_9758,N_9229,N_9484);
nand U9759 (N_9759,N_9218,N_9567);
nand U9760 (N_9760,N_9193,N_9234);
xor U9761 (N_9761,N_9432,N_9153);
and U9762 (N_9762,N_9414,N_9028);
nand U9763 (N_9763,N_9440,N_9499);
nor U9764 (N_9764,N_9281,N_9543);
xnor U9765 (N_9765,N_9205,N_9032);
nor U9766 (N_9766,N_9073,N_9171);
nand U9767 (N_9767,N_9497,N_9339);
and U9768 (N_9768,N_9565,N_9528);
nor U9769 (N_9769,N_9126,N_9371);
and U9770 (N_9770,N_9237,N_9527);
nor U9771 (N_9771,N_9069,N_9454);
nor U9772 (N_9772,N_9057,N_9078);
nand U9773 (N_9773,N_9482,N_9333);
and U9774 (N_9774,N_9305,N_9013);
xnor U9775 (N_9775,N_9570,N_9531);
and U9776 (N_9776,N_9597,N_9089);
xnor U9777 (N_9777,N_9383,N_9211);
nand U9778 (N_9778,N_9390,N_9144);
nand U9779 (N_9779,N_9519,N_9088);
or U9780 (N_9780,N_9494,N_9109);
nor U9781 (N_9781,N_9592,N_9362);
or U9782 (N_9782,N_9227,N_9418);
or U9783 (N_9783,N_9147,N_9085);
nand U9784 (N_9784,N_9331,N_9431);
and U9785 (N_9785,N_9195,N_9044);
or U9786 (N_9786,N_9186,N_9271);
nor U9787 (N_9787,N_9026,N_9006);
and U9788 (N_9788,N_9508,N_9404);
xor U9789 (N_9789,N_9327,N_9550);
nand U9790 (N_9790,N_9420,N_9158);
xnor U9791 (N_9791,N_9525,N_9475);
nand U9792 (N_9792,N_9521,N_9163);
and U9793 (N_9793,N_9348,N_9479);
or U9794 (N_9794,N_9240,N_9568);
nand U9795 (N_9795,N_9571,N_9307);
nand U9796 (N_9796,N_9010,N_9364);
and U9797 (N_9797,N_9342,N_9444);
xnor U9798 (N_9798,N_9399,N_9016);
nand U9799 (N_9799,N_9520,N_9311);
and U9800 (N_9800,N_9512,N_9395);
and U9801 (N_9801,N_9130,N_9366);
nand U9802 (N_9802,N_9443,N_9090);
xnor U9803 (N_9803,N_9075,N_9151);
nand U9804 (N_9804,N_9018,N_9584);
nand U9805 (N_9805,N_9401,N_9441);
and U9806 (N_9806,N_9236,N_9047);
and U9807 (N_9807,N_9081,N_9477);
or U9808 (N_9808,N_9204,N_9403);
xnor U9809 (N_9809,N_9396,N_9168);
nand U9810 (N_9810,N_9124,N_9221);
and U9811 (N_9811,N_9164,N_9326);
or U9812 (N_9812,N_9043,N_9288);
or U9813 (N_9813,N_9516,N_9286);
nor U9814 (N_9814,N_9058,N_9048);
xnor U9815 (N_9815,N_9127,N_9292);
nor U9816 (N_9816,N_9301,N_9556);
nand U9817 (N_9817,N_9489,N_9071);
xnor U9818 (N_9818,N_9091,N_9260);
nand U9819 (N_9819,N_9102,N_9099);
nor U9820 (N_9820,N_9340,N_9583);
nor U9821 (N_9821,N_9488,N_9303);
nor U9822 (N_9822,N_9353,N_9354);
and U9823 (N_9823,N_9123,N_9586);
nor U9824 (N_9824,N_9513,N_9458);
nand U9825 (N_9825,N_9397,N_9341);
or U9826 (N_9826,N_9182,N_9059);
and U9827 (N_9827,N_9378,N_9530);
nand U9828 (N_9828,N_9213,N_9179);
nor U9829 (N_9829,N_9037,N_9201);
and U9830 (N_9830,N_9491,N_9255);
or U9831 (N_9831,N_9092,N_9192);
and U9832 (N_9832,N_9111,N_9025);
or U9833 (N_9833,N_9230,N_9250);
nand U9834 (N_9834,N_9501,N_9587);
xnor U9835 (N_9835,N_9167,N_9217);
nand U9836 (N_9836,N_9448,N_9533);
or U9837 (N_9837,N_9290,N_9351);
xor U9838 (N_9838,N_9358,N_9170);
nand U9839 (N_9839,N_9593,N_9232);
xnor U9840 (N_9840,N_9514,N_9188);
and U9841 (N_9841,N_9140,N_9551);
nor U9842 (N_9842,N_9379,N_9405);
and U9843 (N_9843,N_9313,N_9314);
and U9844 (N_9844,N_9107,N_9066);
nand U9845 (N_9845,N_9319,N_9540);
nor U9846 (N_9846,N_9261,N_9049);
or U9847 (N_9847,N_9408,N_9282);
or U9848 (N_9848,N_9503,N_9014);
nand U9849 (N_9849,N_9476,N_9157);
or U9850 (N_9850,N_9100,N_9180);
and U9851 (N_9851,N_9599,N_9133);
and U9852 (N_9852,N_9038,N_9323);
nand U9853 (N_9853,N_9427,N_9350);
nor U9854 (N_9854,N_9005,N_9352);
nor U9855 (N_9855,N_9359,N_9214);
or U9856 (N_9856,N_9079,N_9256);
and U9857 (N_9857,N_9463,N_9553);
nand U9858 (N_9858,N_9173,N_9253);
xor U9859 (N_9859,N_9287,N_9335);
nand U9860 (N_9860,N_9295,N_9267);
or U9861 (N_9861,N_9070,N_9492);
nand U9862 (N_9862,N_9430,N_9564);
nand U9863 (N_9863,N_9585,N_9566);
and U9864 (N_9864,N_9027,N_9189);
nand U9865 (N_9865,N_9380,N_9452);
and U9866 (N_9866,N_9231,N_9415);
and U9867 (N_9867,N_9591,N_9275);
and U9868 (N_9868,N_9065,N_9375);
and U9869 (N_9869,N_9391,N_9461);
nand U9870 (N_9870,N_9177,N_9579);
or U9871 (N_9871,N_9264,N_9387);
nor U9872 (N_9872,N_9321,N_9084);
nor U9873 (N_9873,N_9203,N_9118);
or U9874 (N_9874,N_9577,N_9460);
nor U9875 (N_9875,N_9258,N_9128);
nand U9876 (N_9876,N_9064,N_9464);
or U9877 (N_9877,N_9558,N_9406);
nor U9878 (N_9878,N_9276,N_9266);
nor U9879 (N_9879,N_9051,N_9074);
and U9880 (N_9880,N_9035,N_9561);
and U9881 (N_9881,N_9112,N_9363);
or U9882 (N_9882,N_9176,N_9060);
and U9883 (N_9883,N_9019,N_9145);
and U9884 (N_9884,N_9113,N_9419);
and U9885 (N_9885,N_9122,N_9247);
nor U9886 (N_9886,N_9457,N_9110);
and U9887 (N_9887,N_9098,N_9325);
nor U9888 (N_9888,N_9506,N_9220);
xor U9889 (N_9889,N_9165,N_9053);
nor U9890 (N_9890,N_9539,N_9486);
or U9891 (N_9891,N_9382,N_9456);
and U9892 (N_9892,N_9595,N_9212);
or U9893 (N_9893,N_9175,N_9262);
xor U9894 (N_9894,N_9374,N_9442);
nor U9895 (N_9895,N_9329,N_9132);
xnor U9896 (N_9896,N_9563,N_9172);
or U9897 (N_9897,N_9268,N_9009);
and U9898 (N_9898,N_9279,N_9017);
nand U9899 (N_9899,N_9117,N_9542);
and U9900 (N_9900,N_9285,N_9371);
nor U9901 (N_9901,N_9373,N_9476);
nor U9902 (N_9902,N_9423,N_9332);
or U9903 (N_9903,N_9256,N_9588);
nand U9904 (N_9904,N_9033,N_9350);
nor U9905 (N_9905,N_9484,N_9593);
nor U9906 (N_9906,N_9500,N_9261);
nand U9907 (N_9907,N_9560,N_9575);
nor U9908 (N_9908,N_9586,N_9232);
nand U9909 (N_9909,N_9280,N_9307);
and U9910 (N_9910,N_9334,N_9054);
nor U9911 (N_9911,N_9205,N_9237);
nand U9912 (N_9912,N_9164,N_9490);
and U9913 (N_9913,N_9030,N_9223);
and U9914 (N_9914,N_9042,N_9582);
nand U9915 (N_9915,N_9245,N_9294);
xnor U9916 (N_9916,N_9512,N_9022);
and U9917 (N_9917,N_9019,N_9275);
xor U9918 (N_9918,N_9352,N_9351);
or U9919 (N_9919,N_9433,N_9469);
nor U9920 (N_9920,N_9441,N_9472);
nor U9921 (N_9921,N_9125,N_9599);
or U9922 (N_9922,N_9013,N_9459);
nor U9923 (N_9923,N_9223,N_9094);
nand U9924 (N_9924,N_9108,N_9555);
or U9925 (N_9925,N_9069,N_9172);
nand U9926 (N_9926,N_9200,N_9013);
xor U9927 (N_9927,N_9072,N_9093);
and U9928 (N_9928,N_9503,N_9274);
nand U9929 (N_9929,N_9509,N_9315);
nor U9930 (N_9930,N_9474,N_9472);
and U9931 (N_9931,N_9306,N_9587);
or U9932 (N_9932,N_9539,N_9091);
nand U9933 (N_9933,N_9102,N_9576);
and U9934 (N_9934,N_9149,N_9055);
nand U9935 (N_9935,N_9474,N_9092);
nor U9936 (N_9936,N_9075,N_9431);
and U9937 (N_9937,N_9247,N_9460);
and U9938 (N_9938,N_9326,N_9156);
nor U9939 (N_9939,N_9023,N_9417);
xor U9940 (N_9940,N_9467,N_9582);
nor U9941 (N_9941,N_9106,N_9189);
nor U9942 (N_9942,N_9522,N_9202);
xnor U9943 (N_9943,N_9566,N_9273);
and U9944 (N_9944,N_9077,N_9221);
nand U9945 (N_9945,N_9564,N_9004);
or U9946 (N_9946,N_9274,N_9318);
or U9947 (N_9947,N_9291,N_9006);
nand U9948 (N_9948,N_9422,N_9539);
nor U9949 (N_9949,N_9138,N_9112);
nor U9950 (N_9950,N_9561,N_9253);
or U9951 (N_9951,N_9483,N_9104);
and U9952 (N_9952,N_9161,N_9399);
nor U9953 (N_9953,N_9329,N_9308);
nand U9954 (N_9954,N_9195,N_9346);
and U9955 (N_9955,N_9120,N_9096);
and U9956 (N_9956,N_9115,N_9207);
and U9957 (N_9957,N_9319,N_9559);
or U9958 (N_9958,N_9468,N_9133);
nand U9959 (N_9959,N_9325,N_9145);
or U9960 (N_9960,N_9217,N_9085);
and U9961 (N_9961,N_9406,N_9364);
or U9962 (N_9962,N_9211,N_9384);
nor U9963 (N_9963,N_9075,N_9095);
nand U9964 (N_9964,N_9162,N_9283);
or U9965 (N_9965,N_9518,N_9044);
nor U9966 (N_9966,N_9443,N_9507);
and U9967 (N_9967,N_9131,N_9010);
nor U9968 (N_9968,N_9247,N_9346);
nor U9969 (N_9969,N_9374,N_9553);
nor U9970 (N_9970,N_9002,N_9206);
or U9971 (N_9971,N_9029,N_9077);
or U9972 (N_9972,N_9168,N_9103);
nor U9973 (N_9973,N_9497,N_9019);
nor U9974 (N_9974,N_9153,N_9047);
nand U9975 (N_9975,N_9044,N_9390);
or U9976 (N_9976,N_9117,N_9448);
and U9977 (N_9977,N_9149,N_9228);
and U9978 (N_9978,N_9278,N_9426);
nor U9979 (N_9979,N_9487,N_9074);
and U9980 (N_9980,N_9477,N_9518);
nor U9981 (N_9981,N_9315,N_9414);
nand U9982 (N_9982,N_9547,N_9108);
nor U9983 (N_9983,N_9475,N_9551);
xor U9984 (N_9984,N_9144,N_9089);
or U9985 (N_9985,N_9341,N_9411);
and U9986 (N_9986,N_9299,N_9526);
and U9987 (N_9987,N_9395,N_9138);
and U9988 (N_9988,N_9549,N_9415);
nor U9989 (N_9989,N_9069,N_9132);
and U9990 (N_9990,N_9284,N_9383);
xnor U9991 (N_9991,N_9450,N_9090);
or U9992 (N_9992,N_9369,N_9015);
nor U9993 (N_9993,N_9249,N_9468);
xor U9994 (N_9994,N_9349,N_9249);
nor U9995 (N_9995,N_9246,N_9191);
or U9996 (N_9996,N_9528,N_9431);
nor U9997 (N_9997,N_9522,N_9588);
xnor U9998 (N_9998,N_9592,N_9204);
nor U9999 (N_9999,N_9379,N_9396);
and U10000 (N_10000,N_9097,N_9364);
or U10001 (N_10001,N_9166,N_9590);
and U10002 (N_10002,N_9387,N_9497);
nor U10003 (N_10003,N_9182,N_9260);
and U10004 (N_10004,N_9112,N_9480);
nand U10005 (N_10005,N_9271,N_9108);
nand U10006 (N_10006,N_9284,N_9121);
and U10007 (N_10007,N_9508,N_9156);
nor U10008 (N_10008,N_9595,N_9040);
nand U10009 (N_10009,N_9040,N_9356);
and U10010 (N_10010,N_9405,N_9018);
nand U10011 (N_10011,N_9313,N_9320);
and U10012 (N_10012,N_9173,N_9394);
nand U10013 (N_10013,N_9577,N_9129);
xor U10014 (N_10014,N_9433,N_9108);
or U10015 (N_10015,N_9153,N_9068);
nor U10016 (N_10016,N_9302,N_9367);
nor U10017 (N_10017,N_9051,N_9296);
and U10018 (N_10018,N_9425,N_9595);
or U10019 (N_10019,N_9152,N_9436);
nand U10020 (N_10020,N_9546,N_9191);
nor U10021 (N_10021,N_9575,N_9144);
and U10022 (N_10022,N_9508,N_9172);
nor U10023 (N_10023,N_9034,N_9193);
or U10024 (N_10024,N_9091,N_9434);
and U10025 (N_10025,N_9494,N_9387);
and U10026 (N_10026,N_9517,N_9191);
nand U10027 (N_10027,N_9163,N_9421);
nand U10028 (N_10028,N_9514,N_9065);
or U10029 (N_10029,N_9015,N_9471);
and U10030 (N_10030,N_9075,N_9278);
nor U10031 (N_10031,N_9439,N_9147);
or U10032 (N_10032,N_9308,N_9356);
nor U10033 (N_10033,N_9108,N_9386);
nor U10034 (N_10034,N_9552,N_9293);
nor U10035 (N_10035,N_9199,N_9109);
and U10036 (N_10036,N_9047,N_9195);
nand U10037 (N_10037,N_9049,N_9334);
nand U10038 (N_10038,N_9463,N_9211);
nand U10039 (N_10039,N_9007,N_9578);
xor U10040 (N_10040,N_9244,N_9158);
nand U10041 (N_10041,N_9470,N_9544);
xnor U10042 (N_10042,N_9067,N_9426);
and U10043 (N_10043,N_9532,N_9027);
nand U10044 (N_10044,N_9414,N_9244);
nor U10045 (N_10045,N_9351,N_9585);
nor U10046 (N_10046,N_9495,N_9453);
or U10047 (N_10047,N_9425,N_9014);
xnor U10048 (N_10048,N_9557,N_9340);
xor U10049 (N_10049,N_9083,N_9143);
and U10050 (N_10050,N_9378,N_9059);
or U10051 (N_10051,N_9336,N_9073);
nor U10052 (N_10052,N_9124,N_9471);
and U10053 (N_10053,N_9008,N_9498);
or U10054 (N_10054,N_9220,N_9333);
and U10055 (N_10055,N_9039,N_9491);
and U10056 (N_10056,N_9054,N_9372);
and U10057 (N_10057,N_9551,N_9395);
and U10058 (N_10058,N_9148,N_9493);
and U10059 (N_10059,N_9398,N_9136);
and U10060 (N_10060,N_9328,N_9548);
or U10061 (N_10061,N_9022,N_9583);
and U10062 (N_10062,N_9513,N_9500);
and U10063 (N_10063,N_9005,N_9042);
or U10064 (N_10064,N_9169,N_9083);
and U10065 (N_10065,N_9548,N_9252);
or U10066 (N_10066,N_9454,N_9551);
nor U10067 (N_10067,N_9551,N_9455);
or U10068 (N_10068,N_9059,N_9430);
nand U10069 (N_10069,N_9499,N_9088);
nor U10070 (N_10070,N_9346,N_9505);
nand U10071 (N_10071,N_9216,N_9132);
xor U10072 (N_10072,N_9116,N_9102);
nor U10073 (N_10073,N_9156,N_9065);
and U10074 (N_10074,N_9521,N_9526);
nand U10075 (N_10075,N_9198,N_9590);
and U10076 (N_10076,N_9264,N_9331);
and U10077 (N_10077,N_9504,N_9006);
nand U10078 (N_10078,N_9434,N_9064);
and U10079 (N_10079,N_9226,N_9334);
and U10080 (N_10080,N_9021,N_9385);
nand U10081 (N_10081,N_9401,N_9300);
or U10082 (N_10082,N_9407,N_9401);
or U10083 (N_10083,N_9492,N_9547);
nand U10084 (N_10084,N_9079,N_9095);
nand U10085 (N_10085,N_9182,N_9045);
or U10086 (N_10086,N_9531,N_9423);
nand U10087 (N_10087,N_9354,N_9529);
or U10088 (N_10088,N_9058,N_9529);
xnor U10089 (N_10089,N_9489,N_9537);
or U10090 (N_10090,N_9154,N_9401);
nand U10091 (N_10091,N_9533,N_9334);
nand U10092 (N_10092,N_9088,N_9467);
nand U10093 (N_10093,N_9010,N_9374);
xor U10094 (N_10094,N_9392,N_9380);
and U10095 (N_10095,N_9319,N_9576);
and U10096 (N_10096,N_9226,N_9280);
or U10097 (N_10097,N_9424,N_9207);
and U10098 (N_10098,N_9101,N_9164);
and U10099 (N_10099,N_9597,N_9407);
nor U10100 (N_10100,N_9470,N_9407);
or U10101 (N_10101,N_9253,N_9303);
nand U10102 (N_10102,N_9096,N_9239);
nand U10103 (N_10103,N_9468,N_9140);
nand U10104 (N_10104,N_9348,N_9201);
nor U10105 (N_10105,N_9386,N_9408);
and U10106 (N_10106,N_9524,N_9166);
or U10107 (N_10107,N_9585,N_9436);
nand U10108 (N_10108,N_9287,N_9575);
or U10109 (N_10109,N_9285,N_9016);
or U10110 (N_10110,N_9223,N_9460);
or U10111 (N_10111,N_9282,N_9023);
nand U10112 (N_10112,N_9588,N_9136);
and U10113 (N_10113,N_9564,N_9455);
nand U10114 (N_10114,N_9186,N_9534);
nor U10115 (N_10115,N_9587,N_9383);
or U10116 (N_10116,N_9358,N_9283);
nand U10117 (N_10117,N_9133,N_9260);
nor U10118 (N_10118,N_9002,N_9545);
or U10119 (N_10119,N_9532,N_9335);
or U10120 (N_10120,N_9424,N_9575);
nor U10121 (N_10121,N_9177,N_9525);
and U10122 (N_10122,N_9521,N_9338);
or U10123 (N_10123,N_9005,N_9534);
and U10124 (N_10124,N_9459,N_9042);
nor U10125 (N_10125,N_9227,N_9426);
nor U10126 (N_10126,N_9597,N_9055);
or U10127 (N_10127,N_9129,N_9462);
or U10128 (N_10128,N_9373,N_9263);
and U10129 (N_10129,N_9425,N_9515);
nand U10130 (N_10130,N_9394,N_9343);
xnor U10131 (N_10131,N_9588,N_9396);
xnor U10132 (N_10132,N_9090,N_9059);
and U10133 (N_10133,N_9443,N_9537);
nor U10134 (N_10134,N_9455,N_9308);
and U10135 (N_10135,N_9047,N_9188);
nor U10136 (N_10136,N_9404,N_9038);
or U10137 (N_10137,N_9091,N_9115);
nand U10138 (N_10138,N_9203,N_9241);
or U10139 (N_10139,N_9391,N_9214);
nor U10140 (N_10140,N_9379,N_9016);
nand U10141 (N_10141,N_9364,N_9021);
nand U10142 (N_10142,N_9035,N_9229);
nor U10143 (N_10143,N_9249,N_9548);
nor U10144 (N_10144,N_9417,N_9591);
or U10145 (N_10145,N_9394,N_9448);
and U10146 (N_10146,N_9328,N_9109);
or U10147 (N_10147,N_9352,N_9316);
nand U10148 (N_10148,N_9383,N_9503);
nor U10149 (N_10149,N_9067,N_9517);
xor U10150 (N_10150,N_9545,N_9412);
and U10151 (N_10151,N_9497,N_9266);
nand U10152 (N_10152,N_9225,N_9209);
xor U10153 (N_10153,N_9579,N_9254);
or U10154 (N_10154,N_9543,N_9045);
or U10155 (N_10155,N_9092,N_9523);
or U10156 (N_10156,N_9427,N_9187);
nor U10157 (N_10157,N_9319,N_9080);
nor U10158 (N_10158,N_9197,N_9531);
nand U10159 (N_10159,N_9113,N_9123);
or U10160 (N_10160,N_9377,N_9040);
xor U10161 (N_10161,N_9476,N_9187);
nor U10162 (N_10162,N_9328,N_9459);
xor U10163 (N_10163,N_9193,N_9059);
nand U10164 (N_10164,N_9156,N_9294);
and U10165 (N_10165,N_9594,N_9573);
nand U10166 (N_10166,N_9293,N_9043);
and U10167 (N_10167,N_9544,N_9510);
nand U10168 (N_10168,N_9537,N_9518);
nand U10169 (N_10169,N_9298,N_9235);
nand U10170 (N_10170,N_9345,N_9424);
nand U10171 (N_10171,N_9284,N_9421);
nor U10172 (N_10172,N_9108,N_9365);
or U10173 (N_10173,N_9028,N_9432);
nor U10174 (N_10174,N_9426,N_9292);
nor U10175 (N_10175,N_9509,N_9258);
nand U10176 (N_10176,N_9526,N_9162);
nor U10177 (N_10177,N_9208,N_9175);
xnor U10178 (N_10178,N_9500,N_9199);
and U10179 (N_10179,N_9207,N_9168);
nand U10180 (N_10180,N_9257,N_9127);
nor U10181 (N_10181,N_9482,N_9353);
and U10182 (N_10182,N_9312,N_9153);
or U10183 (N_10183,N_9537,N_9244);
or U10184 (N_10184,N_9034,N_9122);
or U10185 (N_10185,N_9118,N_9085);
nor U10186 (N_10186,N_9119,N_9349);
xnor U10187 (N_10187,N_9024,N_9376);
nand U10188 (N_10188,N_9355,N_9359);
xor U10189 (N_10189,N_9407,N_9520);
and U10190 (N_10190,N_9475,N_9268);
nand U10191 (N_10191,N_9015,N_9163);
and U10192 (N_10192,N_9271,N_9163);
nor U10193 (N_10193,N_9301,N_9107);
xor U10194 (N_10194,N_9041,N_9049);
nand U10195 (N_10195,N_9125,N_9288);
and U10196 (N_10196,N_9171,N_9475);
or U10197 (N_10197,N_9159,N_9014);
or U10198 (N_10198,N_9529,N_9541);
nand U10199 (N_10199,N_9189,N_9243);
nor U10200 (N_10200,N_10080,N_9768);
or U10201 (N_10201,N_10031,N_9693);
nand U10202 (N_10202,N_10090,N_9675);
nand U10203 (N_10203,N_10182,N_10169);
xor U10204 (N_10204,N_10128,N_10092);
nor U10205 (N_10205,N_10006,N_10066);
xnor U10206 (N_10206,N_10039,N_9850);
nor U10207 (N_10207,N_10180,N_9866);
and U10208 (N_10208,N_9940,N_9791);
or U10209 (N_10209,N_9824,N_9711);
and U10210 (N_10210,N_9612,N_9947);
or U10211 (N_10211,N_10196,N_9935);
nor U10212 (N_10212,N_10011,N_10168);
or U10213 (N_10213,N_9702,N_10094);
or U10214 (N_10214,N_9857,N_10042);
xor U10215 (N_10215,N_10164,N_9709);
or U10216 (N_10216,N_9622,N_10149);
and U10217 (N_10217,N_9881,N_9821);
nor U10218 (N_10218,N_10097,N_9671);
nand U10219 (N_10219,N_9945,N_9964);
nor U10220 (N_10220,N_10134,N_9925);
xor U10221 (N_10221,N_9831,N_9839);
xor U10222 (N_10222,N_9764,N_10067);
and U10223 (N_10223,N_9782,N_9994);
and U10224 (N_10224,N_10010,N_9962);
and U10225 (N_10225,N_10107,N_9752);
or U10226 (N_10226,N_9636,N_10142);
nand U10227 (N_10227,N_9692,N_9921);
nor U10228 (N_10228,N_9713,N_10029);
and U10229 (N_10229,N_9859,N_9984);
and U10230 (N_10230,N_10102,N_9733);
xor U10231 (N_10231,N_9797,N_10181);
nor U10232 (N_10232,N_9919,N_9851);
nor U10233 (N_10233,N_9684,N_9965);
nand U10234 (N_10234,N_10130,N_10028);
nor U10235 (N_10235,N_9981,N_9832);
nor U10236 (N_10236,N_9785,N_9882);
nand U10237 (N_10237,N_9651,N_9760);
xor U10238 (N_10238,N_9813,N_10157);
and U10239 (N_10239,N_10001,N_9941);
xnor U10240 (N_10240,N_10139,N_10162);
or U10241 (N_10241,N_9890,N_10171);
nor U10242 (N_10242,N_9732,N_9986);
or U10243 (N_10243,N_9877,N_10145);
or U10244 (N_10244,N_9619,N_9845);
xnor U10245 (N_10245,N_9765,N_9812);
or U10246 (N_10246,N_9611,N_10060);
nand U10247 (N_10247,N_9840,N_9978);
or U10248 (N_10248,N_9663,N_9817);
nor U10249 (N_10249,N_9911,N_9932);
and U10250 (N_10250,N_9971,N_10193);
nand U10251 (N_10251,N_9621,N_9718);
or U10252 (N_10252,N_9977,N_10043);
or U10253 (N_10253,N_9893,N_9920);
and U10254 (N_10254,N_9620,N_10105);
nand U10255 (N_10255,N_9873,N_10106);
nand U10256 (N_10256,N_9694,N_9686);
nor U10257 (N_10257,N_10146,N_9799);
nand U10258 (N_10258,N_9802,N_10199);
nand U10259 (N_10259,N_9604,N_9959);
or U10260 (N_10260,N_10034,N_9916);
nor U10261 (N_10261,N_9735,N_10174);
nand U10262 (N_10262,N_10095,N_10191);
xor U10263 (N_10263,N_10023,N_10100);
and U10264 (N_10264,N_9901,N_9938);
and U10265 (N_10265,N_9736,N_9892);
xor U10266 (N_10266,N_9753,N_9697);
or U10267 (N_10267,N_9703,N_9979);
xnor U10268 (N_10268,N_9862,N_10198);
or U10269 (N_10269,N_9689,N_9673);
nand U10270 (N_10270,N_10190,N_9654);
nor U10271 (N_10271,N_9951,N_9679);
nor U10272 (N_10272,N_10115,N_10004);
and U10273 (N_10273,N_9770,N_9647);
and U10274 (N_10274,N_9649,N_10108);
or U10275 (N_10275,N_9833,N_9741);
and U10276 (N_10276,N_10120,N_9909);
and U10277 (N_10277,N_9665,N_10084);
and U10278 (N_10278,N_9742,N_9615);
nand U10279 (N_10279,N_9894,N_10113);
nand U10280 (N_10280,N_9754,N_9729);
or U10281 (N_10281,N_10119,N_10082);
nand U10282 (N_10282,N_9837,N_9633);
and U10283 (N_10283,N_9625,N_9639);
nor U10284 (N_10284,N_10192,N_9670);
nor U10285 (N_10285,N_10148,N_10132);
nand U10286 (N_10286,N_10059,N_9931);
or U10287 (N_10287,N_9823,N_9895);
or U10288 (N_10288,N_10177,N_9744);
or U10289 (N_10289,N_9800,N_9776);
or U10290 (N_10290,N_10026,N_10194);
nand U10291 (N_10291,N_9769,N_10050);
nor U10292 (N_10292,N_9674,N_9705);
xnor U10293 (N_10293,N_10047,N_9721);
xor U10294 (N_10294,N_10065,N_9726);
nor U10295 (N_10295,N_10159,N_9700);
xor U10296 (N_10296,N_10014,N_10013);
or U10297 (N_10297,N_10183,N_9676);
and U10298 (N_10298,N_10165,N_9956);
nand U10299 (N_10299,N_9645,N_10179);
or U10300 (N_10300,N_9614,N_10027);
nand U10301 (N_10301,N_9870,N_9999);
or U10302 (N_10302,N_10144,N_9723);
and U10303 (N_10303,N_9610,N_10071);
and U10304 (N_10304,N_9695,N_9655);
or U10305 (N_10305,N_9637,N_9880);
nor U10306 (N_10306,N_9899,N_9788);
or U10307 (N_10307,N_9868,N_9953);
nor U10308 (N_10308,N_9680,N_9662);
and U10309 (N_10309,N_9943,N_10051);
xnor U10310 (N_10310,N_9808,N_9898);
or U10311 (N_10311,N_9929,N_10086);
nor U10312 (N_10312,N_9838,N_9657);
and U10313 (N_10313,N_9900,N_10055);
nand U10314 (N_10314,N_9896,N_9747);
nand U10315 (N_10315,N_9653,N_10061);
nand U10316 (N_10316,N_9728,N_10103);
and U10317 (N_10317,N_9714,N_9988);
or U10318 (N_10318,N_10155,N_9950);
and U10319 (N_10319,N_10138,N_9716);
xor U10320 (N_10320,N_10070,N_9652);
and U10321 (N_10321,N_9822,N_9827);
or U10322 (N_10322,N_9624,N_9631);
and U10323 (N_10323,N_10158,N_9740);
xnor U10324 (N_10324,N_9967,N_9779);
or U10325 (N_10325,N_9889,N_9973);
and U10326 (N_10326,N_9816,N_9918);
and U10327 (N_10327,N_9660,N_9915);
and U10328 (N_10328,N_9600,N_9616);
nor U10329 (N_10329,N_9961,N_9640);
or U10330 (N_10330,N_10077,N_10019);
nor U10331 (N_10331,N_9972,N_10046);
nor U10332 (N_10332,N_9887,N_10007);
nand U10333 (N_10333,N_9980,N_9609);
or U10334 (N_10334,N_10154,N_10140);
nor U10335 (N_10335,N_10135,N_9623);
or U10336 (N_10336,N_9668,N_9603);
and U10337 (N_10337,N_9731,N_9939);
nor U10338 (N_10338,N_9884,N_9745);
and U10339 (N_10339,N_10081,N_10064);
xor U10340 (N_10340,N_9917,N_9794);
or U10341 (N_10341,N_10121,N_10189);
nor U10342 (N_10342,N_9869,N_10116);
or U10343 (N_10343,N_9613,N_9946);
nor U10344 (N_10344,N_10101,N_9682);
or U10345 (N_10345,N_9722,N_9825);
nor U10346 (N_10346,N_10003,N_9989);
and U10347 (N_10347,N_9725,N_9948);
and U10348 (N_10348,N_9853,N_9960);
or U10349 (N_10349,N_10187,N_9908);
and U10350 (N_10350,N_9867,N_10000);
and U10351 (N_10351,N_10052,N_9914);
xnor U10352 (N_10352,N_9963,N_9834);
and U10353 (N_10353,N_9991,N_9927);
and U10354 (N_10354,N_10131,N_9706);
and U10355 (N_10355,N_9924,N_9875);
and U10356 (N_10356,N_9987,N_9701);
nand U10357 (N_10357,N_10170,N_10127);
xor U10358 (N_10358,N_10020,N_9997);
nand U10359 (N_10359,N_10163,N_9803);
nand U10360 (N_10360,N_10160,N_9712);
nand U10361 (N_10361,N_10037,N_9661);
or U10362 (N_10362,N_10109,N_9758);
nor U10363 (N_10363,N_10150,N_9638);
xor U10364 (N_10364,N_9974,N_9798);
and U10365 (N_10365,N_9677,N_10173);
nand U10366 (N_10366,N_10074,N_10078);
nand U10367 (N_10367,N_10035,N_9905);
or U10368 (N_10368,N_9605,N_10175);
nor U10369 (N_10369,N_9687,N_9781);
xor U10370 (N_10370,N_9936,N_9757);
and U10371 (N_10371,N_9790,N_9910);
and U10372 (N_10372,N_9944,N_9763);
xnor U10373 (N_10373,N_9952,N_9678);
and U10374 (N_10374,N_10056,N_10021);
xor U10375 (N_10375,N_10033,N_9830);
nor U10376 (N_10376,N_10125,N_9902);
and U10377 (N_10377,N_9975,N_9658);
xnor U10378 (N_10378,N_10025,N_9930);
or U10379 (N_10379,N_10091,N_10118);
nand U10380 (N_10380,N_9617,N_9864);
xnor U10381 (N_10381,N_10012,N_9897);
or U10382 (N_10382,N_9937,N_9985);
nor U10383 (N_10383,N_9828,N_9659);
nor U10384 (N_10384,N_9844,N_10188);
and U10385 (N_10385,N_10040,N_9771);
nor U10386 (N_10386,N_9811,N_9842);
and U10387 (N_10387,N_9883,N_9871);
nand U10388 (N_10388,N_9970,N_9778);
xor U10389 (N_10389,N_9809,N_10104);
nor U10390 (N_10390,N_9826,N_10110);
nor U10391 (N_10391,N_9847,N_9724);
nor U10392 (N_10392,N_10072,N_10076);
nor U10393 (N_10393,N_10141,N_10186);
nor U10394 (N_10394,N_10147,N_9786);
or U10395 (N_10395,N_9957,N_9983);
or U10396 (N_10396,N_10063,N_10195);
nand U10397 (N_10397,N_9632,N_10032);
or U10398 (N_10398,N_10111,N_9669);
nand U10399 (N_10399,N_10112,N_9629);
nand U10400 (N_10400,N_10041,N_9904);
nor U10401 (N_10401,N_9843,N_9969);
and U10402 (N_10402,N_9933,N_9708);
or U10403 (N_10403,N_9698,N_10079);
nand U10404 (N_10404,N_10178,N_9998);
and U10405 (N_10405,N_10185,N_9751);
nor U10406 (N_10406,N_9648,N_10015);
nor U10407 (N_10407,N_10114,N_9688);
and U10408 (N_10408,N_10049,N_9903);
nor U10409 (N_10409,N_9681,N_9642);
xor U10410 (N_10410,N_10083,N_9804);
nand U10411 (N_10411,N_9913,N_10089);
or U10412 (N_10412,N_9734,N_9759);
nand U10413 (N_10413,N_9926,N_9955);
nand U10414 (N_10414,N_10133,N_9958);
or U10415 (N_10415,N_9923,N_10129);
or U10416 (N_10416,N_9618,N_10093);
or U10417 (N_10417,N_9691,N_9646);
or U10418 (N_10418,N_10058,N_9772);
xor U10419 (N_10419,N_9699,N_9942);
nor U10420 (N_10420,N_10017,N_10124);
nand U10421 (N_10421,N_10151,N_9750);
or U10422 (N_10422,N_9710,N_9690);
and U10423 (N_10423,N_9746,N_9849);
nor U10424 (N_10424,N_9879,N_9641);
xnor U10425 (N_10425,N_9878,N_10024);
and U10426 (N_10426,N_10016,N_9861);
nor U10427 (N_10427,N_9773,N_10172);
or U10428 (N_10428,N_10096,N_10156);
or U10429 (N_10429,N_9966,N_9891);
or U10430 (N_10430,N_9995,N_9912);
nor U10431 (N_10431,N_9719,N_9818);
nor U10432 (N_10432,N_9730,N_9715);
nor U10433 (N_10433,N_9643,N_9886);
and U10434 (N_10434,N_9819,N_9787);
nor U10435 (N_10435,N_9801,N_9792);
and U10436 (N_10436,N_9874,N_9820);
nand U10437 (N_10437,N_9656,N_9876);
or U10438 (N_10438,N_9888,N_9858);
or U10439 (N_10439,N_9872,N_10008);
or U10440 (N_10440,N_9806,N_9644);
and U10441 (N_10441,N_10038,N_9755);
or U10442 (N_10442,N_10068,N_9739);
and U10443 (N_10443,N_9934,N_9990);
and U10444 (N_10444,N_9907,N_9696);
nand U10445 (N_10445,N_10153,N_10184);
and U10446 (N_10446,N_9780,N_9627);
or U10447 (N_10447,N_9727,N_9650);
or U10448 (N_10448,N_10062,N_10044);
or U10449 (N_10449,N_9683,N_9664);
nand U10450 (N_10450,N_9704,N_10002);
or U10451 (N_10451,N_9814,N_10167);
or U10452 (N_10452,N_10030,N_9863);
xnor U10453 (N_10453,N_9717,N_10054);
nor U10454 (N_10454,N_10088,N_10087);
nor U10455 (N_10455,N_10018,N_9628);
or U10456 (N_10456,N_9992,N_9855);
and U10457 (N_10457,N_9738,N_9602);
nor U10458 (N_10458,N_9666,N_9885);
and U10459 (N_10459,N_9793,N_9626);
nor U10460 (N_10460,N_10137,N_9836);
or U10461 (N_10461,N_9749,N_9634);
or U10462 (N_10462,N_9685,N_9852);
nor U10463 (N_10463,N_9607,N_10073);
and U10464 (N_10464,N_9635,N_10117);
nand U10465 (N_10465,N_9982,N_9996);
nor U10466 (N_10466,N_9796,N_9954);
nand U10467 (N_10467,N_9810,N_9928);
and U10468 (N_10468,N_10053,N_9761);
nor U10469 (N_10469,N_9795,N_9672);
and U10470 (N_10470,N_9829,N_9968);
and U10471 (N_10471,N_10122,N_9846);
or U10472 (N_10472,N_9630,N_10009);
or U10473 (N_10473,N_9766,N_9922);
xnor U10474 (N_10474,N_10022,N_9601);
or U10475 (N_10475,N_10166,N_10048);
and U10476 (N_10476,N_10152,N_9854);
nor U10477 (N_10477,N_10143,N_9848);
nor U10478 (N_10478,N_9667,N_10045);
or U10479 (N_10479,N_9606,N_9865);
nor U10480 (N_10480,N_9835,N_9748);
nor U10481 (N_10481,N_10036,N_10057);
and U10482 (N_10482,N_9976,N_9743);
xnor U10483 (N_10483,N_9784,N_10075);
xnor U10484 (N_10484,N_9807,N_9756);
nor U10485 (N_10485,N_9860,N_10099);
nand U10486 (N_10486,N_9949,N_10069);
nor U10487 (N_10487,N_10085,N_9762);
nand U10488 (N_10488,N_10197,N_9720);
xor U10489 (N_10489,N_9805,N_10098);
and U10490 (N_10490,N_10123,N_9775);
nor U10491 (N_10491,N_10161,N_10126);
nor U10492 (N_10492,N_9789,N_10136);
nand U10493 (N_10493,N_9774,N_9777);
nor U10494 (N_10494,N_9767,N_9993);
nand U10495 (N_10495,N_9707,N_9841);
xnor U10496 (N_10496,N_9815,N_9783);
xnor U10497 (N_10497,N_9856,N_9737);
nand U10498 (N_10498,N_10005,N_9608);
nor U10499 (N_10499,N_10176,N_9906);
or U10500 (N_10500,N_9904,N_9812);
or U10501 (N_10501,N_9683,N_10048);
nor U10502 (N_10502,N_10152,N_9758);
and U10503 (N_10503,N_9800,N_10125);
and U10504 (N_10504,N_9982,N_9925);
or U10505 (N_10505,N_9929,N_10090);
or U10506 (N_10506,N_9787,N_9734);
or U10507 (N_10507,N_9603,N_10016);
xor U10508 (N_10508,N_9918,N_10002);
and U10509 (N_10509,N_9794,N_9947);
nor U10510 (N_10510,N_9931,N_10099);
xnor U10511 (N_10511,N_9734,N_9907);
xor U10512 (N_10512,N_10011,N_10027);
and U10513 (N_10513,N_9757,N_9697);
xnor U10514 (N_10514,N_10048,N_9751);
nor U10515 (N_10515,N_10033,N_10018);
or U10516 (N_10516,N_9736,N_10023);
nand U10517 (N_10517,N_9916,N_9843);
xnor U10518 (N_10518,N_9728,N_9966);
and U10519 (N_10519,N_9847,N_9772);
xnor U10520 (N_10520,N_9703,N_9710);
nand U10521 (N_10521,N_9712,N_9815);
and U10522 (N_10522,N_9775,N_10008);
nor U10523 (N_10523,N_9846,N_9792);
nand U10524 (N_10524,N_10028,N_10035);
or U10525 (N_10525,N_10184,N_10179);
and U10526 (N_10526,N_10114,N_10130);
nor U10527 (N_10527,N_9905,N_10084);
nor U10528 (N_10528,N_10054,N_10138);
or U10529 (N_10529,N_9960,N_9607);
nor U10530 (N_10530,N_9776,N_9986);
nor U10531 (N_10531,N_9752,N_9934);
or U10532 (N_10532,N_9976,N_10194);
or U10533 (N_10533,N_9882,N_10115);
nand U10534 (N_10534,N_9916,N_9853);
xnor U10535 (N_10535,N_9910,N_9948);
xor U10536 (N_10536,N_10193,N_10174);
nor U10537 (N_10537,N_10163,N_9823);
nand U10538 (N_10538,N_9632,N_10163);
nor U10539 (N_10539,N_9623,N_10183);
nor U10540 (N_10540,N_9941,N_10153);
nor U10541 (N_10541,N_10100,N_10014);
nand U10542 (N_10542,N_9929,N_9608);
xnor U10543 (N_10543,N_9715,N_10141);
or U10544 (N_10544,N_9885,N_9989);
xnor U10545 (N_10545,N_10131,N_9784);
or U10546 (N_10546,N_10137,N_9879);
nor U10547 (N_10547,N_9752,N_9630);
nor U10548 (N_10548,N_10023,N_10049);
nand U10549 (N_10549,N_10002,N_9818);
xnor U10550 (N_10550,N_10109,N_10131);
and U10551 (N_10551,N_9827,N_10001);
and U10552 (N_10552,N_9920,N_9962);
nor U10553 (N_10553,N_9999,N_10013);
or U10554 (N_10554,N_9904,N_9640);
nand U10555 (N_10555,N_10144,N_10193);
and U10556 (N_10556,N_10158,N_9617);
and U10557 (N_10557,N_9731,N_10161);
nand U10558 (N_10558,N_9874,N_10059);
nand U10559 (N_10559,N_9768,N_9793);
nor U10560 (N_10560,N_9694,N_9628);
nor U10561 (N_10561,N_10158,N_10150);
and U10562 (N_10562,N_9679,N_10062);
nor U10563 (N_10563,N_10002,N_10034);
nor U10564 (N_10564,N_10142,N_9640);
and U10565 (N_10565,N_9877,N_9655);
nand U10566 (N_10566,N_10043,N_9805);
xor U10567 (N_10567,N_10028,N_9662);
and U10568 (N_10568,N_9642,N_9609);
or U10569 (N_10569,N_10122,N_9912);
or U10570 (N_10570,N_9620,N_9736);
or U10571 (N_10571,N_9997,N_10130);
or U10572 (N_10572,N_10020,N_9608);
nor U10573 (N_10573,N_10181,N_9879);
or U10574 (N_10574,N_9661,N_10063);
and U10575 (N_10575,N_9762,N_10019);
and U10576 (N_10576,N_9704,N_9992);
nand U10577 (N_10577,N_9758,N_9605);
and U10578 (N_10578,N_9897,N_9860);
or U10579 (N_10579,N_9827,N_10199);
or U10580 (N_10580,N_9689,N_9659);
and U10581 (N_10581,N_10120,N_9841);
nor U10582 (N_10582,N_10019,N_9836);
nand U10583 (N_10583,N_9683,N_9710);
or U10584 (N_10584,N_10023,N_9643);
nand U10585 (N_10585,N_9788,N_10081);
xnor U10586 (N_10586,N_10032,N_9776);
or U10587 (N_10587,N_9754,N_9931);
or U10588 (N_10588,N_9933,N_9795);
or U10589 (N_10589,N_9657,N_9976);
nor U10590 (N_10590,N_10042,N_10152);
and U10591 (N_10591,N_10189,N_10158);
and U10592 (N_10592,N_10132,N_9652);
or U10593 (N_10593,N_9739,N_9664);
and U10594 (N_10594,N_10058,N_10147);
or U10595 (N_10595,N_9847,N_10037);
xor U10596 (N_10596,N_9613,N_9681);
xor U10597 (N_10597,N_10026,N_9772);
or U10598 (N_10598,N_9616,N_10100);
or U10599 (N_10599,N_9758,N_9743);
nand U10600 (N_10600,N_9693,N_10137);
nor U10601 (N_10601,N_9719,N_9956);
nor U10602 (N_10602,N_9668,N_9723);
and U10603 (N_10603,N_10089,N_10040);
xor U10604 (N_10604,N_9963,N_9936);
and U10605 (N_10605,N_10017,N_9810);
nor U10606 (N_10606,N_10111,N_9962);
nand U10607 (N_10607,N_9808,N_10033);
nand U10608 (N_10608,N_10082,N_9923);
nor U10609 (N_10609,N_9611,N_9755);
and U10610 (N_10610,N_10031,N_9700);
nand U10611 (N_10611,N_10023,N_9613);
xnor U10612 (N_10612,N_9829,N_10034);
and U10613 (N_10613,N_10017,N_9737);
nor U10614 (N_10614,N_9662,N_9895);
nand U10615 (N_10615,N_9891,N_9929);
xor U10616 (N_10616,N_9884,N_9998);
nand U10617 (N_10617,N_9955,N_9672);
nor U10618 (N_10618,N_10091,N_10134);
or U10619 (N_10619,N_9797,N_10086);
or U10620 (N_10620,N_9943,N_9979);
nor U10621 (N_10621,N_9882,N_9755);
and U10622 (N_10622,N_9834,N_9629);
nor U10623 (N_10623,N_9638,N_10179);
nor U10624 (N_10624,N_10114,N_9799);
xnor U10625 (N_10625,N_9717,N_9842);
xor U10626 (N_10626,N_9814,N_10186);
or U10627 (N_10627,N_10150,N_10089);
xnor U10628 (N_10628,N_9625,N_9815);
or U10629 (N_10629,N_10173,N_9792);
or U10630 (N_10630,N_9825,N_10074);
or U10631 (N_10631,N_10153,N_10190);
and U10632 (N_10632,N_9967,N_10118);
nand U10633 (N_10633,N_10116,N_9960);
and U10634 (N_10634,N_9933,N_10010);
or U10635 (N_10635,N_9633,N_10178);
or U10636 (N_10636,N_9776,N_9900);
xnor U10637 (N_10637,N_9611,N_9920);
xnor U10638 (N_10638,N_9734,N_9834);
nand U10639 (N_10639,N_9815,N_9689);
and U10640 (N_10640,N_9952,N_9630);
nor U10641 (N_10641,N_9901,N_10073);
nand U10642 (N_10642,N_9938,N_10116);
xnor U10643 (N_10643,N_9815,N_9914);
and U10644 (N_10644,N_9823,N_9903);
and U10645 (N_10645,N_9870,N_9702);
xor U10646 (N_10646,N_9813,N_9645);
nand U10647 (N_10647,N_9686,N_10132);
nor U10648 (N_10648,N_9632,N_9755);
and U10649 (N_10649,N_10037,N_9720);
nand U10650 (N_10650,N_10094,N_10183);
xor U10651 (N_10651,N_9951,N_9815);
or U10652 (N_10652,N_10075,N_10162);
and U10653 (N_10653,N_9809,N_9703);
or U10654 (N_10654,N_9634,N_10074);
nand U10655 (N_10655,N_9831,N_9838);
or U10656 (N_10656,N_10021,N_10101);
and U10657 (N_10657,N_10193,N_9749);
xnor U10658 (N_10658,N_10112,N_10151);
nor U10659 (N_10659,N_10031,N_10114);
nor U10660 (N_10660,N_9665,N_9697);
and U10661 (N_10661,N_10026,N_9617);
nand U10662 (N_10662,N_10179,N_10007);
and U10663 (N_10663,N_10188,N_9600);
or U10664 (N_10664,N_10047,N_10173);
nand U10665 (N_10665,N_10004,N_9980);
or U10666 (N_10666,N_9960,N_10028);
or U10667 (N_10667,N_9711,N_10077);
nor U10668 (N_10668,N_10148,N_9862);
and U10669 (N_10669,N_9792,N_9912);
nor U10670 (N_10670,N_9679,N_9864);
nand U10671 (N_10671,N_9828,N_9817);
nor U10672 (N_10672,N_10145,N_10090);
and U10673 (N_10673,N_9646,N_10009);
nand U10674 (N_10674,N_10136,N_9885);
and U10675 (N_10675,N_9655,N_9788);
nand U10676 (N_10676,N_10167,N_10080);
nand U10677 (N_10677,N_10139,N_10199);
nor U10678 (N_10678,N_10127,N_10123);
nand U10679 (N_10679,N_10195,N_10163);
nor U10680 (N_10680,N_9652,N_9635);
or U10681 (N_10681,N_9935,N_9646);
and U10682 (N_10682,N_9885,N_9700);
nand U10683 (N_10683,N_9913,N_9874);
nand U10684 (N_10684,N_9711,N_9776);
xnor U10685 (N_10685,N_9953,N_9883);
xnor U10686 (N_10686,N_10063,N_9668);
xor U10687 (N_10687,N_9864,N_9994);
nand U10688 (N_10688,N_9958,N_9686);
or U10689 (N_10689,N_10146,N_10110);
nor U10690 (N_10690,N_10134,N_10078);
xor U10691 (N_10691,N_10049,N_10139);
or U10692 (N_10692,N_10059,N_10093);
xor U10693 (N_10693,N_10140,N_9921);
and U10694 (N_10694,N_9674,N_9824);
nor U10695 (N_10695,N_9889,N_9875);
nor U10696 (N_10696,N_9702,N_10072);
or U10697 (N_10697,N_9688,N_10062);
nor U10698 (N_10698,N_9627,N_10151);
nand U10699 (N_10699,N_10166,N_9652);
and U10700 (N_10700,N_10171,N_9776);
nand U10701 (N_10701,N_10068,N_9667);
xnor U10702 (N_10702,N_9848,N_9694);
or U10703 (N_10703,N_9629,N_9674);
nand U10704 (N_10704,N_9622,N_9699);
or U10705 (N_10705,N_9888,N_9613);
nand U10706 (N_10706,N_10046,N_10131);
and U10707 (N_10707,N_10117,N_10178);
or U10708 (N_10708,N_9831,N_10093);
or U10709 (N_10709,N_9812,N_10131);
or U10710 (N_10710,N_9669,N_9723);
and U10711 (N_10711,N_10139,N_9900);
nor U10712 (N_10712,N_9604,N_9769);
and U10713 (N_10713,N_10192,N_9925);
or U10714 (N_10714,N_9787,N_9612);
nand U10715 (N_10715,N_10073,N_9983);
nand U10716 (N_10716,N_9947,N_9941);
nor U10717 (N_10717,N_9714,N_9841);
and U10718 (N_10718,N_9727,N_9695);
nand U10719 (N_10719,N_9749,N_9759);
nand U10720 (N_10720,N_9707,N_9862);
nor U10721 (N_10721,N_9967,N_10166);
nand U10722 (N_10722,N_10017,N_9869);
or U10723 (N_10723,N_9895,N_9830);
nor U10724 (N_10724,N_10112,N_9886);
or U10725 (N_10725,N_9643,N_10190);
or U10726 (N_10726,N_9752,N_10081);
or U10727 (N_10727,N_10092,N_9902);
and U10728 (N_10728,N_9635,N_9929);
xor U10729 (N_10729,N_9707,N_10118);
and U10730 (N_10730,N_9692,N_10168);
and U10731 (N_10731,N_10062,N_9780);
nand U10732 (N_10732,N_10026,N_10187);
nor U10733 (N_10733,N_9941,N_10144);
or U10734 (N_10734,N_9764,N_9845);
or U10735 (N_10735,N_9720,N_9874);
or U10736 (N_10736,N_9839,N_10153);
nand U10737 (N_10737,N_10143,N_10054);
or U10738 (N_10738,N_9809,N_10002);
xnor U10739 (N_10739,N_10124,N_9902);
xnor U10740 (N_10740,N_9631,N_9848);
nand U10741 (N_10741,N_10141,N_9705);
or U10742 (N_10742,N_9885,N_9652);
nor U10743 (N_10743,N_9854,N_9879);
nor U10744 (N_10744,N_10062,N_10085);
and U10745 (N_10745,N_10121,N_10146);
nand U10746 (N_10746,N_9682,N_10084);
nand U10747 (N_10747,N_9880,N_9974);
or U10748 (N_10748,N_9610,N_9981);
xor U10749 (N_10749,N_9891,N_9802);
or U10750 (N_10750,N_9893,N_10166);
nor U10751 (N_10751,N_10101,N_10143);
or U10752 (N_10752,N_9918,N_10062);
nand U10753 (N_10753,N_9608,N_9773);
nand U10754 (N_10754,N_9681,N_9965);
xnor U10755 (N_10755,N_9624,N_9704);
or U10756 (N_10756,N_9622,N_10183);
nor U10757 (N_10757,N_9889,N_10127);
or U10758 (N_10758,N_9616,N_9801);
and U10759 (N_10759,N_10186,N_9773);
nand U10760 (N_10760,N_9926,N_9603);
or U10761 (N_10761,N_10099,N_9997);
and U10762 (N_10762,N_9735,N_9993);
nand U10763 (N_10763,N_10086,N_9796);
nor U10764 (N_10764,N_9744,N_9673);
nor U10765 (N_10765,N_9693,N_9942);
nand U10766 (N_10766,N_9945,N_9831);
and U10767 (N_10767,N_9634,N_9751);
or U10768 (N_10768,N_9856,N_9943);
or U10769 (N_10769,N_9809,N_10073);
and U10770 (N_10770,N_10029,N_9817);
xor U10771 (N_10771,N_10041,N_9800);
xnor U10772 (N_10772,N_10038,N_9697);
nand U10773 (N_10773,N_10138,N_9720);
nand U10774 (N_10774,N_9911,N_10142);
or U10775 (N_10775,N_10063,N_9689);
nor U10776 (N_10776,N_10085,N_9817);
and U10777 (N_10777,N_9755,N_10030);
or U10778 (N_10778,N_9855,N_10134);
or U10779 (N_10779,N_10079,N_9955);
xnor U10780 (N_10780,N_10135,N_9752);
nor U10781 (N_10781,N_9665,N_9843);
xor U10782 (N_10782,N_9656,N_10197);
nor U10783 (N_10783,N_9667,N_9941);
and U10784 (N_10784,N_9920,N_10075);
and U10785 (N_10785,N_9777,N_9789);
nor U10786 (N_10786,N_9719,N_9943);
nand U10787 (N_10787,N_10068,N_9967);
and U10788 (N_10788,N_9844,N_10105);
nor U10789 (N_10789,N_9856,N_9734);
and U10790 (N_10790,N_9720,N_9846);
or U10791 (N_10791,N_9685,N_9809);
and U10792 (N_10792,N_9747,N_9891);
or U10793 (N_10793,N_9659,N_10154);
or U10794 (N_10794,N_9795,N_9914);
or U10795 (N_10795,N_9900,N_10032);
xor U10796 (N_10796,N_10017,N_9735);
nor U10797 (N_10797,N_9803,N_9721);
xor U10798 (N_10798,N_9679,N_9971);
and U10799 (N_10799,N_10040,N_9866);
or U10800 (N_10800,N_10753,N_10763);
xnor U10801 (N_10801,N_10252,N_10262);
and U10802 (N_10802,N_10237,N_10224);
nor U10803 (N_10803,N_10661,N_10527);
xnor U10804 (N_10804,N_10694,N_10256);
xor U10805 (N_10805,N_10208,N_10706);
and U10806 (N_10806,N_10647,N_10730);
nor U10807 (N_10807,N_10359,N_10350);
or U10808 (N_10808,N_10562,N_10475);
or U10809 (N_10809,N_10419,N_10717);
nand U10810 (N_10810,N_10467,N_10388);
and U10811 (N_10811,N_10689,N_10269);
nor U10812 (N_10812,N_10457,N_10234);
or U10813 (N_10813,N_10557,N_10501);
nand U10814 (N_10814,N_10740,N_10746);
nand U10815 (N_10815,N_10522,N_10623);
or U10816 (N_10816,N_10507,N_10679);
nand U10817 (N_10817,N_10701,N_10541);
or U10818 (N_10818,N_10500,N_10751);
xnor U10819 (N_10819,N_10696,N_10456);
nand U10820 (N_10820,N_10630,N_10596);
nor U10821 (N_10821,N_10211,N_10606);
nor U10822 (N_10822,N_10330,N_10563);
nand U10823 (N_10823,N_10555,N_10727);
xnor U10824 (N_10824,N_10624,N_10705);
or U10825 (N_10825,N_10474,N_10543);
nand U10826 (N_10826,N_10473,N_10495);
xnor U10827 (N_10827,N_10690,N_10489);
and U10828 (N_10828,N_10616,N_10514);
xnor U10829 (N_10829,N_10564,N_10317);
and U10830 (N_10830,N_10712,N_10586);
or U10831 (N_10831,N_10212,N_10568);
or U10832 (N_10832,N_10481,N_10447);
nor U10833 (N_10833,N_10608,N_10750);
nand U10834 (N_10834,N_10280,N_10595);
or U10835 (N_10835,N_10486,N_10675);
or U10836 (N_10836,N_10699,N_10780);
xnor U10837 (N_10837,N_10505,N_10542);
nor U10838 (N_10838,N_10321,N_10633);
xor U10839 (N_10839,N_10381,N_10778);
nand U10840 (N_10840,N_10272,N_10358);
nand U10841 (N_10841,N_10508,N_10723);
and U10842 (N_10842,N_10663,N_10498);
nand U10843 (N_10843,N_10270,N_10493);
and U10844 (N_10844,N_10782,N_10697);
xor U10845 (N_10845,N_10672,N_10503);
or U10846 (N_10846,N_10646,N_10353);
and U10847 (N_10847,N_10504,N_10776);
and U10848 (N_10848,N_10335,N_10682);
nor U10849 (N_10849,N_10588,N_10627);
or U10850 (N_10850,N_10768,N_10573);
xor U10851 (N_10851,N_10619,N_10389);
nand U10852 (N_10852,N_10228,N_10214);
or U10853 (N_10853,N_10472,N_10253);
nor U10854 (N_10854,N_10202,N_10668);
nor U10855 (N_10855,N_10366,N_10714);
or U10856 (N_10856,N_10632,N_10655);
nor U10857 (N_10857,N_10677,N_10391);
nand U10858 (N_10858,N_10692,N_10683);
nor U10859 (N_10859,N_10653,N_10297);
nor U10860 (N_10860,N_10725,N_10521);
and U10861 (N_10861,N_10615,N_10238);
nand U10862 (N_10862,N_10468,N_10511);
or U10863 (N_10863,N_10652,N_10748);
or U10864 (N_10864,N_10572,N_10332);
or U10865 (N_10865,N_10245,N_10276);
or U10866 (N_10866,N_10334,N_10518);
nor U10867 (N_10867,N_10392,N_10715);
nor U10868 (N_10868,N_10759,N_10409);
nand U10869 (N_10869,N_10635,N_10546);
or U10870 (N_10870,N_10517,N_10614);
xnor U10871 (N_10871,N_10303,N_10470);
or U10872 (N_10872,N_10769,N_10549);
nor U10873 (N_10873,N_10729,N_10399);
nor U10874 (N_10874,N_10600,N_10241);
nor U10875 (N_10875,N_10316,N_10434);
and U10876 (N_10876,N_10482,N_10320);
and U10877 (N_10877,N_10658,N_10345);
xnor U10878 (N_10878,N_10499,N_10580);
and U10879 (N_10879,N_10250,N_10449);
or U10880 (N_10880,N_10758,N_10306);
or U10881 (N_10881,N_10414,N_10743);
nand U10882 (N_10882,N_10342,N_10469);
xor U10883 (N_10883,N_10213,N_10446);
nor U10884 (N_10884,N_10719,N_10516);
or U10885 (N_10885,N_10754,N_10631);
nand U10886 (N_10886,N_10257,N_10230);
and U10887 (N_10887,N_10556,N_10322);
nor U10888 (N_10888,N_10403,N_10298);
or U10889 (N_10889,N_10536,N_10310);
nand U10890 (N_10890,N_10458,N_10231);
or U10891 (N_10891,N_10251,N_10464);
nand U10892 (N_10892,N_10533,N_10369);
or U10893 (N_10893,N_10311,N_10361);
or U10894 (N_10894,N_10355,N_10590);
and U10895 (N_10895,N_10227,N_10520);
nand U10896 (N_10896,N_10534,N_10747);
nor U10897 (N_10897,N_10233,N_10745);
or U10898 (N_10898,N_10724,N_10432);
and U10899 (N_10899,N_10477,N_10589);
nor U10900 (N_10900,N_10360,N_10574);
nand U10901 (N_10901,N_10279,N_10277);
or U10902 (N_10902,N_10378,N_10443);
or U10903 (N_10903,N_10436,N_10703);
or U10904 (N_10904,N_10288,N_10762);
xor U10905 (N_10905,N_10643,N_10576);
nand U10906 (N_10906,N_10741,N_10215);
nor U10907 (N_10907,N_10738,N_10259);
nor U10908 (N_10908,N_10242,N_10220);
nor U10909 (N_10909,N_10203,N_10711);
nand U10910 (N_10910,N_10347,N_10771);
or U10911 (N_10911,N_10471,N_10532);
nand U10912 (N_10912,N_10509,N_10271);
nor U10913 (N_10913,N_10581,N_10790);
xor U10914 (N_10914,N_10236,N_10396);
and U10915 (N_10915,N_10433,N_10798);
and U10916 (N_10916,N_10226,N_10638);
nor U10917 (N_10917,N_10451,N_10216);
or U10918 (N_10918,N_10368,N_10340);
xor U10919 (N_10919,N_10229,N_10654);
or U10920 (N_10920,N_10352,N_10752);
nor U10921 (N_10921,N_10268,N_10283);
or U10922 (N_10922,N_10626,N_10726);
and U10923 (N_10923,N_10793,N_10442);
nor U10924 (N_10924,N_10485,N_10222);
nand U10925 (N_10925,N_10554,N_10328);
nand U10926 (N_10926,N_10372,N_10487);
or U10927 (N_10927,N_10354,N_10367);
nand U10928 (N_10928,N_10435,N_10687);
and U10929 (N_10929,N_10707,N_10666);
and U10930 (N_10930,N_10788,N_10585);
or U10931 (N_10931,N_10651,N_10783);
nand U10932 (N_10932,N_10480,N_10244);
or U10933 (N_10933,N_10329,N_10286);
nand U10934 (N_10934,N_10429,N_10767);
nor U10935 (N_10935,N_10376,N_10620);
nand U10936 (N_10936,N_10698,N_10667);
xor U10937 (N_10937,N_10761,N_10789);
xor U10938 (N_10938,N_10544,N_10278);
xnor U10939 (N_10939,N_10406,N_10284);
nand U10940 (N_10940,N_10383,N_10225);
and U10941 (N_10941,N_10559,N_10611);
or U10942 (N_10942,N_10219,N_10774);
nor U10943 (N_10943,N_10281,N_10301);
xor U10944 (N_10944,N_10425,N_10295);
nand U10945 (N_10945,N_10304,N_10773);
or U10946 (N_10946,N_10408,N_10326);
or U10947 (N_10947,N_10263,N_10410);
and U10948 (N_10948,N_10343,N_10318);
or U10949 (N_10949,N_10599,N_10494);
nor U10950 (N_10950,N_10609,N_10642);
nor U10951 (N_10951,N_10421,N_10604);
nor U10952 (N_10952,N_10413,N_10398);
and U10953 (N_10953,N_10681,N_10657);
and U10954 (N_10954,N_10323,N_10339);
xor U10955 (N_10955,N_10426,N_10374);
or U10956 (N_10956,N_10382,N_10377);
or U10957 (N_10957,N_10757,N_10201);
nor U10958 (N_10958,N_10553,N_10356);
nor U10959 (N_10959,N_10441,N_10660);
and U10960 (N_10960,N_10756,N_10478);
or U10961 (N_10961,N_10584,N_10267);
nand U10962 (N_10962,N_10733,N_10274);
or U10963 (N_10963,N_10404,N_10292);
xnor U10964 (N_10964,N_10445,N_10363);
nor U10965 (N_10965,N_10770,N_10387);
xnor U10966 (N_10966,N_10612,N_10415);
nand U10967 (N_10967,N_10315,N_10693);
xor U10968 (N_10968,N_10560,N_10338);
nand U10969 (N_10969,N_10607,N_10598);
or U10970 (N_10970,N_10314,N_10716);
or U10971 (N_10971,N_10566,N_10465);
or U10972 (N_10972,N_10676,N_10275);
and U10973 (N_10973,N_10680,N_10497);
and U10974 (N_10974,N_10254,N_10325);
or U10975 (N_10975,N_10764,N_10476);
and U10976 (N_10976,N_10571,N_10351);
nor U10977 (N_10977,N_10791,N_10591);
nor U10978 (N_10978,N_10248,N_10308);
xor U10979 (N_10979,N_10496,N_10309);
and U10980 (N_10980,N_10427,N_10385);
nor U10981 (N_10981,N_10512,N_10362);
or U10982 (N_10982,N_10760,N_10649);
or U10983 (N_10983,N_10695,N_10390);
xor U10984 (N_10984,N_10529,N_10735);
or U10985 (N_10985,N_10484,N_10491);
xnor U10986 (N_10986,N_10772,N_10299);
and U10987 (N_10987,N_10691,N_10221);
nor U10988 (N_10988,N_10466,N_10266);
nor U10989 (N_10989,N_10525,N_10794);
and U10990 (N_10990,N_10287,N_10765);
and U10991 (N_10991,N_10420,N_10327);
nand U10992 (N_10992,N_10538,N_10460);
or U10993 (N_10993,N_10290,N_10684);
and U10994 (N_10994,N_10438,N_10784);
nor U10995 (N_10995,N_10702,N_10582);
nor U10996 (N_10996,N_10722,N_10688);
nand U10997 (N_10997,N_10336,N_10218);
xnor U10998 (N_10998,N_10437,N_10289);
nor U10999 (N_10999,N_10502,N_10708);
and U11000 (N_11000,N_10239,N_10463);
nand U11001 (N_11001,N_10384,N_10704);
nor U11002 (N_11002,N_10461,N_10728);
nand U11003 (N_11003,N_10319,N_10312);
or U11004 (N_11004,N_10775,N_10428);
or U11005 (N_11005,N_10488,N_10397);
nand U11006 (N_11006,N_10592,N_10510);
nor U11007 (N_11007,N_10575,N_10513);
or U11008 (N_11008,N_10785,N_10720);
nor U11009 (N_11009,N_10417,N_10731);
or U11010 (N_11010,N_10613,N_10567);
and U11011 (N_11011,N_10291,N_10550);
and U11012 (N_11012,N_10313,N_10344);
nand U11013 (N_11013,N_10302,N_10641);
and U11014 (N_11014,N_10204,N_10261);
nand U11015 (N_11015,N_10373,N_10786);
and U11016 (N_11016,N_10346,N_10686);
nor U11017 (N_11017,N_10331,N_10605);
or U11018 (N_11018,N_10732,N_10395);
nand U11019 (N_11019,N_10210,N_10526);
nor U11020 (N_11020,N_10552,N_10602);
and U11021 (N_11021,N_10640,N_10570);
nand U11022 (N_11022,N_10370,N_10670);
nor U11023 (N_11023,N_10448,N_10659);
nor U11024 (N_11024,N_10375,N_10673);
nor U11025 (N_11025,N_10401,N_10781);
nor U11026 (N_11026,N_10528,N_10737);
or U11027 (N_11027,N_10324,N_10547);
and U11028 (N_11028,N_10603,N_10418);
and U11029 (N_11029,N_10628,N_10593);
nor U11030 (N_11030,N_10796,N_10246);
nor U11031 (N_11031,N_10411,N_10223);
or U11032 (N_11032,N_10755,N_10561);
xnor U11033 (N_11033,N_10709,N_10405);
nor U11034 (N_11034,N_10424,N_10459);
and U11035 (N_11035,N_10664,N_10380);
or U11036 (N_11036,N_10548,N_10545);
nand U11037 (N_11037,N_10365,N_10371);
or U11038 (N_11038,N_10622,N_10787);
xor U11039 (N_11039,N_10749,N_10742);
and U11040 (N_11040,N_10407,N_10402);
nand U11041 (N_11041,N_10296,N_10453);
and U11042 (N_11042,N_10379,N_10454);
or U11043 (N_11043,N_10255,N_10247);
and U11044 (N_11044,N_10639,N_10293);
xnor U11045 (N_11045,N_10618,N_10535);
nand U11046 (N_11046,N_10569,N_10349);
or U11047 (N_11047,N_10671,N_10430);
xor U11048 (N_11048,N_10656,N_10779);
nor U11049 (N_11049,N_10736,N_10386);
nand U11050 (N_11050,N_10439,N_10718);
nand U11051 (N_11051,N_10634,N_10440);
or U11052 (N_11052,N_10523,N_10739);
nor U11053 (N_11053,N_10209,N_10610);
nor U11054 (N_11054,N_10583,N_10594);
xnor U11055 (N_11055,N_10205,N_10455);
nor U11056 (N_11056,N_10294,N_10799);
xnor U11057 (N_11057,N_10565,N_10357);
nor U11058 (N_11058,N_10530,N_10282);
nand U11059 (N_11059,N_10539,N_10483);
and U11060 (N_11060,N_10744,N_10524);
nor U11061 (N_11061,N_10700,N_10577);
nor U11062 (N_11062,N_10601,N_10797);
and U11063 (N_11063,N_10551,N_10579);
nor U11064 (N_11064,N_10235,N_10685);
nor U11065 (N_11065,N_10423,N_10207);
nand U11066 (N_11066,N_10249,N_10333);
xor U11067 (N_11067,N_10260,N_10777);
and U11068 (N_11068,N_10531,N_10674);
and U11069 (N_11069,N_10669,N_10490);
or U11070 (N_11070,N_10264,N_10597);
and U11071 (N_11071,N_10393,N_10506);
nand U11072 (N_11072,N_10412,N_10515);
and U11073 (N_11073,N_10452,N_10625);
and U11074 (N_11074,N_10431,N_10519);
and U11075 (N_11075,N_10678,N_10273);
and U11076 (N_11076,N_10400,N_10587);
and U11077 (N_11077,N_10462,N_10710);
or U11078 (N_11078,N_10617,N_10232);
or U11079 (N_11079,N_10578,N_10662);
xnor U11080 (N_11080,N_10665,N_10422);
or U11081 (N_11081,N_10416,N_10265);
and U11082 (N_11082,N_10206,N_10637);
or U11083 (N_11083,N_10450,N_10305);
and U11084 (N_11084,N_10479,N_10537);
nor U11085 (N_11085,N_10348,N_10734);
and U11086 (N_11086,N_10645,N_10492);
xor U11087 (N_11087,N_10285,N_10650);
or U11088 (N_11088,N_10648,N_10644);
xor U11089 (N_11089,N_10217,N_10200);
nand U11090 (N_11090,N_10243,N_10341);
nand U11091 (N_11091,N_10240,N_10558);
nor U11092 (N_11092,N_10795,N_10721);
nand U11093 (N_11093,N_10337,N_10792);
nor U11094 (N_11094,N_10629,N_10300);
nand U11095 (N_11095,N_10636,N_10258);
xor U11096 (N_11096,N_10307,N_10444);
nand U11097 (N_11097,N_10364,N_10540);
nand U11098 (N_11098,N_10621,N_10394);
nor U11099 (N_11099,N_10766,N_10713);
xor U11100 (N_11100,N_10205,N_10574);
nand U11101 (N_11101,N_10368,N_10287);
and U11102 (N_11102,N_10345,N_10537);
nand U11103 (N_11103,N_10234,N_10289);
and U11104 (N_11104,N_10279,N_10329);
and U11105 (N_11105,N_10203,N_10701);
or U11106 (N_11106,N_10362,N_10697);
or U11107 (N_11107,N_10434,N_10219);
nand U11108 (N_11108,N_10645,N_10679);
nor U11109 (N_11109,N_10275,N_10509);
and U11110 (N_11110,N_10627,N_10273);
nand U11111 (N_11111,N_10545,N_10754);
and U11112 (N_11112,N_10494,N_10754);
nand U11113 (N_11113,N_10605,N_10617);
nor U11114 (N_11114,N_10791,N_10481);
or U11115 (N_11115,N_10780,N_10737);
nor U11116 (N_11116,N_10470,N_10365);
nor U11117 (N_11117,N_10730,N_10234);
nand U11118 (N_11118,N_10496,N_10392);
and U11119 (N_11119,N_10406,N_10789);
and U11120 (N_11120,N_10441,N_10253);
or U11121 (N_11121,N_10475,N_10269);
nand U11122 (N_11122,N_10383,N_10215);
xnor U11123 (N_11123,N_10204,N_10789);
or U11124 (N_11124,N_10370,N_10686);
and U11125 (N_11125,N_10406,N_10555);
xnor U11126 (N_11126,N_10226,N_10746);
and U11127 (N_11127,N_10700,N_10468);
nor U11128 (N_11128,N_10789,N_10750);
or U11129 (N_11129,N_10588,N_10544);
or U11130 (N_11130,N_10725,N_10514);
or U11131 (N_11131,N_10728,N_10297);
and U11132 (N_11132,N_10549,N_10683);
or U11133 (N_11133,N_10791,N_10673);
xor U11134 (N_11134,N_10785,N_10472);
nand U11135 (N_11135,N_10558,N_10633);
or U11136 (N_11136,N_10762,N_10269);
nor U11137 (N_11137,N_10631,N_10272);
or U11138 (N_11138,N_10715,N_10659);
nor U11139 (N_11139,N_10263,N_10271);
and U11140 (N_11140,N_10364,N_10725);
or U11141 (N_11141,N_10317,N_10300);
or U11142 (N_11142,N_10354,N_10593);
nand U11143 (N_11143,N_10622,N_10262);
and U11144 (N_11144,N_10444,N_10530);
or U11145 (N_11145,N_10223,N_10420);
or U11146 (N_11146,N_10554,N_10765);
nor U11147 (N_11147,N_10502,N_10649);
xnor U11148 (N_11148,N_10768,N_10277);
nand U11149 (N_11149,N_10531,N_10219);
or U11150 (N_11150,N_10348,N_10532);
nor U11151 (N_11151,N_10624,N_10617);
and U11152 (N_11152,N_10492,N_10607);
or U11153 (N_11153,N_10490,N_10572);
or U11154 (N_11154,N_10761,N_10304);
nor U11155 (N_11155,N_10617,N_10432);
nor U11156 (N_11156,N_10677,N_10483);
nand U11157 (N_11157,N_10547,N_10231);
nor U11158 (N_11158,N_10330,N_10390);
nor U11159 (N_11159,N_10434,N_10685);
nor U11160 (N_11160,N_10760,N_10276);
nand U11161 (N_11161,N_10501,N_10750);
nand U11162 (N_11162,N_10565,N_10799);
xnor U11163 (N_11163,N_10616,N_10351);
xor U11164 (N_11164,N_10263,N_10627);
nand U11165 (N_11165,N_10678,N_10366);
or U11166 (N_11166,N_10214,N_10274);
and U11167 (N_11167,N_10772,N_10458);
nand U11168 (N_11168,N_10662,N_10533);
nor U11169 (N_11169,N_10257,N_10349);
or U11170 (N_11170,N_10477,N_10231);
and U11171 (N_11171,N_10203,N_10325);
nor U11172 (N_11172,N_10506,N_10639);
nand U11173 (N_11173,N_10417,N_10248);
xor U11174 (N_11174,N_10333,N_10782);
nand U11175 (N_11175,N_10641,N_10578);
and U11176 (N_11176,N_10765,N_10783);
or U11177 (N_11177,N_10684,N_10280);
nor U11178 (N_11178,N_10797,N_10431);
and U11179 (N_11179,N_10647,N_10377);
nand U11180 (N_11180,N_10693,N_10427);
nor U11181 (N_11181,N_10792,N_10590);
nor U11182 (N_11182,N_10348,N_10788);
and U11183 (N_11183,N_10547,N_10388);
nand U11184 (N_11184,N_10637,N_10676);
nor U11185 (N_11185,N_10459,N_10421);
xor U11186 (N_11186,N_10524,N_10645);
nand U11187 (N_11187,N_10276,N_10237);
nor U11188 (N_11188,N_10410,N_10294);
nor U11189 (N_11189,N_10239,N_10387);
nand U11190 (N_11190,N_10387,N_10589);
nand U11191 (N_11191,N_10433,N_10417);
nor U11192 (N_11192,N_10788,N_10451);
and U11193 (N_11193,N_10740,N_10576);
and U11194 (N_11194,N_10497,N_10634);
nor U11195 (N_11195,N_10250,N_10444);
xor U11196 (N_11196,N_10608,N_10485);
nor U11197 (N_11197,N_10342,N_10378);
xnor U11198 (N_11198,N_10468,N_10781);
xor U11199 (N_11199,N_10472,N_10481);
nor U11200 (N_11200,N_10393,N_10436);
xnor U11201 (N_11201,N_10543,N_10418);
nor U11202 (N_11202,N_10478,N_10465);
nor U11203 (N_11203,N_10255,N_10398);
or U11204 (N_11204,N_10783,N_10500);
or U11205 (N_11205,N_10330,N_10526);
or U11206 (N_11206,N_10790,N_10767);
nor U11207 (N_11207,N_10610,N_10289);
xor U11208 (N_11208,N_10604,N_10632);
or U11209 (N_11209,N_10634,N_10318);
or U11210 (N_11210,N_10403,N_10719);
nand U11211 (N_11211,N_10336,N_10456);
or U11212 (N_11212,N_10345,N_10686);
nand U11213 (N_11213,N_10427,N_10200);
or U11214 (N_11214,N_10509,N_10763);
or U11215 (N_11215,N_10495,N_10788);
nand U11216 (N_11216,N_10444,N_10686);
nor U11217 (N_11217,N_10688,N_10473);
and U11218 (N_11218,N_10393,N_10649);
nor U11219 (N_11219,N_10242,N_10746);
nor U11220 (N_11220,N_10516,N_10305);
and U11221 (N_11221,N_10792,N_10474);
nand U11222 (N_11222,N_10233,N_10644);
or U11223 (N_11223,N_10354,N_10427);
nand U11224 (N_11224,N_10695,N_10344);
and U11225 (N_11225,N_10336,N_10458);
xnor U11226 (N_11226,N_10322,N_10216);
or U11227 (N_11227,N_10542,N_10797);
or U11228 (N_11228,N_10713,N_10283);
nor U11229 (N_11229,N_10713,N_10445);
nor U11230 (N_11230,N_10476,N_10403);
and U11231 (N_11231,N_10453,N_10540);
nor U11232 (N_11232,N_10730,N_10210);
or U11233 (N_11233,N_10514,N_10724);
or U11234 (N_11234,N_10561,N_10284);
nand U11235 (N_11235,N_10249,N_10361);
xor U11236 (N_11236,N_10473,N_10482);
and U11237 (N_11237,N_10342,N_10798);
or U11238 (N_11238,N_10594,N_10213);
and U11239 (N_11239,N_10305,N_10415);
nand U11240 (N_11240,N_10519,N_10595);
xor U11241 (N_11241,N_10475,N_10598);
nor U11242 (N_11242,N_10491,N_10204);
and U11243 (N_11243,N_10279,N_10591);
and U11244 (N_11244,N_10757,N_10405);
or U11245 (N_11245,N_10723,N_10227);
nor U11246 (N_11246,N_10714,N_10690);
xnor U11247 (N_11247,N_10591,N_10309);
nand U11248 (N_11248,N_10340,N_10201);
and U11249 (N_11249,N_10526,N_10504);
nor U11250 (N_11250,N_10296,N_10313);
or U11251 (N_11251,N_10223,N_10640);
xor U11252 (N_11252,N_10646,N_10432);
or U11253 (N_11253,N_10209,N_10515);
or U11254 (N_11254,N_10444,N_10224);
nor U11255 (N_11255,N_10715,N_10768);
and U11256 (N_11256,N_10778,N_10625);
nor U11257 (N_11257,N_10673,N_10691);
nand U11258 (N_11258,N_10686,N_10680);
nor U11259 (N_11259,N_10418,N_10208);
nor U11260 (N_11260,N_10498,N_10412);
and U11261 (N_11261,N_10431,N_10384);
nand U11262 (N_11262,N_10223,N_10575);
and U11263 (N_11263,N_10785,N_10690);
or U11264 (N_11264,N_10762,N_10478);
nor U11265 (N_11265,N_10281,N_10586);
or U11266 (N_11266,N_10789,N_10729);
or U11267 (N_11267,N_10779,N_10435);
nor U11268 (N_11268,N_10440,N_10754);
nor U11269 (N_11269,N_10363,N_10698);
nor U11270 (N_11270,N_10449,N_10366);
nand U11271 (N_11271,N_10534,N_10568);
nand U11272 (N_11272,N_10714,N_10406);
or U11273 (N_11273,N_10575,N_10619);
and U11274 (N_11274,N_10313,N_10676);
nand U11275 (N_11275,N_10721,N_10780);
nor U11276 (N_11276,N_10748,N_10440);
and U11277 (N_11277,N_10473,N_10255);
or U11278 (N_11278,N_10419,N_10407);
nand U11279 (N_11279,N_10767,N_10776);
and U11280 (N_11280,N_10294,N_10272);
and U11281 (N_11281,N_10311,N_10285);
nor U11282 (N_11282,N_10207,N_10770);
and U11283 (N_11283,N_10663,N_10555);
nand U11284 (N_11284,N_10405,N_10699);
or U11285 (N_11285,N_10302,N_10408);
nor U11286 (N_11286,N_10227,N_10572);
or U11287 (N_11287,N_10224,N_10434);
and U11288 (N_11288,N_10496,N_10284);
nor U11289 (N_11289,N_10540,N_10243);
nand U11290 (N_11290,N_10411,N_10215);
and U11291 (N_11291,N_10412,N_10615);
and U11292 (N_11292,N_10224,N_10518);
or U11293 (N_11293,N_10205,N_10682);
nand U11294 (N_11294,N_10631,N_10461);
nand U11295 (N_11295,N_10780,N_10637);
and U11296 (N_11296,N_10209,N_10660);
and U11297 (N_11297,N_10539,N_10207);
and U11298 (N_11298,N_10410,N_10513);
nor U11299 (N_11299,N_10519,N_10447);
and U11300 (N_11300,N_10334,N_10499);
nor U11301 (N_11301,N_10615,N_10658);
nor U11302 (N_11302,N_10360,N_10281);
xor U11303 (N_11303,N_10463,N_10469);
or U11304 (N_11304,N_10473,N_10743);
and U11305 (N_11305,N_10217,N_10389);
or U11306 (N_11306,N_10516,N_10598);
nand U11307 (N_11307,N_10399,N_10491);
or U11308 (N_11308,N_10431,N_10265);
or U11309 (N_11309,N_10249,N_10586);
nor U11310 (N_11310,N_10747,N_10319);
and U11311 (N_11311,N_10689,N_10552);
or U11312 (N_11312,N_10592,N_10670);
or U11313 (N_11313,N_10320,N_10651);
or U11314 (N_11314,N_10770,N_10260);
nand U11315 (N_11315,N_10663,N_10239);
or U11316 (N_11316,N_10284,N_10316);
or U11317 (N_11317,N_10336,N_10511);
or U11318 (N_11318,N_10725,N_10263);
and U11319 (N_11319,N_10730,N_10512);
or U11320 (N_11320,N_10746,N_10418);
and U11321 (N_11321,N_10557,N_10527);
xor U11322 (N_11322,N_10441,N_10464);
and U11323 (N_11323,N_10697,N_10300);
nor U11324 (N_11324,N_10549,N_10744);
xor U11325 (N_11325,N_10729,N_10582);
xor U11326 (N_11326,N_10755,N_10502);
or U11327 (N_11327,N_10780,N_10716);
and U11328 (N_11328,N_10309,N_10240);
or U11329 (N_11329,N_10448,N_10620);
or U11330 (N_11330,N_10356,N_10635);
nand U11331 (N_11331,N_10410,N_10507);
nand U11332 (N_11332,N_10655,N_10732);
nand U11333 (N_11333,N_10569,N_10269);
or U11334 (N_11334,N_10348,N_10360);
nor U11335 (N_11335,N_10473,N_10219);
nor U11336 (N_11336,N_10506,N_10783);
or U11337 (N_11337,N_10768,N_10220);
nor U11338 (N_11338,N_10272,N_10442);
or U11339 (N_11339,N_10445,N_10781);
or U11340 (N_11340,N_10343,N_10620);
or U11341 (N_11341,N_10783,N_10413);
or U11342 (N_11342,N_10605,N_10562);
xnor U11343 (N_11343,N_10752,N_10585);
and U11344 (N_11344,N_10234,N_10236);
xor U11345 (N_11345,N_10420,N_10402);
and U11346 (N_11346,N_10360,N_10297);
or U11347 (N_11347,N_10327,N_10759);
and U11348 (N_11348,N_10216,N_10775);
xor U11349 (N_11349,N_10361,N_10707);
nand U11350 (N_11350,N_10378,N_10627);
nor U11351 (N_11351,N_10775,N_10632);
xnor U11352 (N_11352,N_10475,N_10408);
and U11353 (N_11353,N_10432,N_10241);
nor U11354 (N_11354,N_10571,N_10498);
nand U11355 (N_11355,N_10747,N_10244);
nor U11356 (N_11356,N_10478,N_10272);
nor U11357 (N_11357,N_10225,N_10541);
or U11358 (N_11358,N_10797,N_10792);
nand U11359 (N_11359,N_10461,N_10673);
nor U11360 (N_11360,N_10202,N_10723);
or U11361 (N_11361,N_10437,N_10631);
or U11362 (N_11362,N_10440,N_10503);
and U11363 (N_11363,N_10484,N_10216);
or U11364 (N_11364,N_10755,N_10283);
and U11365 (N_11365,N_10454,N_10458);
nor U11366 (N_11366,N_10765,N_10620);
xnor U11367 (N_11367,N_10767,N_10320);
nand U11368 (N_11368,N_10559,N_10780);
or U11369 (N_11369,N_10264,N_10505);
and U11370 (N_11370,N_10635,N_10699);
or U11371 (N_11371,N_10234,N_10696);
and U11372 (N_11372,N_10554,N_10643);
nand U11373 (N_11373,N_10200,N_10288);
and U11374 (N_11374,N_10488,N_10478);
and U11375 (N_11375,N_10293,N_10397);
and U11376 (N_11376,N_10216,N_10793);
and U11377 (N_11377,N_10733,N_10366);
and U11378 (N_11378,N_10362,N_10413);
nor U11379 (N_11379,N_10318,N_10311);
nor U11380 (N_11380,N_10749,N_10510);
nand U11381 (N_11381,N_10575,N_10792);
or U11382 (N_11382,N_10261,N_10705);
nor U11383 (N_11383,N_10610,N_10200);
or U11384 (N_11384,N_10293,N_10573);
or U11385 (N_11385,N_10402,N_10570);
xor U11386 (N_11386,N_10466,N_10448);
xnor U11387 (N_11387,N_10363,N_10577);
nand U11388 (N_11388,N_10548,N_10491);
nor U11389 (N_11389,N_10518,N_10503);
nor U11390 (N_11390,N_10229,N_10500);
nand U11391 (N_11391,N_10232,N_10217);
or U11392 (N_11392,N_10597,N_10755);
or U11393 (N_11393,N_10396,N_10522);
nand U11394 (N_11394,N_10265,N_10601);
nor U11395 (N_11395,N_10666,N_10646);
nor U11396 (N_11396,N_10442,N_10233);
or U11397 (N_11397,N_10733,N_10616);
and U11398 (N_11398,N_10457,N_10799);
xnor U11399 (N_11399,N_10393,N_10263);
and U11400 (N_11400,N_10901,N_10961);
or U11401 (N_11401,N_11258,N_10960);
xor U11402 (N_11402,N_10892,N_11194);
or U11403 (N_11403,N_10885,N_11332);
nand U11404 (N_11404,N_10948,N_10821);
and U11405 (N_11405,N_11054,N_11372);
nor U11406 (N_11406,N_10902,N_11065);
nand U11407 (N_11407,N_11027,N_11102);
or U11408 (N_11408,N_10816,N_10887);
nor U11409 (N_11409,N_11312,N_11385);
and U11410 (N_11410,N_11213,N_10843);
and U11411 (N_11411,N_10943,N_11394);
nor U11412 (N_11412,N_11058,N_10989);
nor U11413 (N_11413,N_10879,N_10907);
xnor U11414 (N_11414,N_10933,N_10818);
nand U11415 (N_11415,N_11056,N_11141);
or U11416 (N_11416,N_11029,N_10815);
nand U11417 (N_11417,N_11344,N_11180);
and U11418 (N_11418,N_11123,N_10840);
nand U11419 (N_11419,N_10918,N_11093);
and U11420 (N_11420,N_11224,N_11092);
nand U11421 (N_11421,N_11111,N_11179);
and U11422 (N_11422,N_10900,N_11061);
nor U11423 (N_11423,N_11361,N_11208);
or U11424 (N_11424,N_11324,N_11059);
nand U11425 (N_11425,N_11013,N_11295);
or U11426 (N_11426,N_11158,N_10847);
nor U11427 (N_11427,N_10866,N_11221);
or U11428 (N_11428,N_11302,N_11209);
or U11429 (N_11429,N_10986,N_11098);
and U11430 (N_11430,N_11137,N_11348);
nand U11431 (N_11431,N_10920,N_11002);
or U11432 (N_11432,N_10898,N_11185);
and U11433 (N_11433,N_10993,N_11379);
nand U11434 (N_11434,N_11251,N_10959);
nor U11435 (N_11435,N_11125,N_11286);
nand U11436 (N_11436,N_11087,N_11193);
nor U11437 (N_11437,N_10809,N_10876);
and U11438 (N_11438,N_11364,N_10908);
nand U11439 (N_11439,N_10995,N_11319);
or U11440 (N_11440,N_11161,N_10917);
nor U11441 (N_11441,N_11060,N_10880);
and U11442 (N_11442,N_11287,N_11064);
and U11443 (N_11443,N_10865,N_11167);
or U11444 (N_11444,N_11025,N_10988);
nand U11445 (N_11445,N_11078,N_11274);
nand U11446 (N_11446,N_11046,N_10916);
nand U11447 (N_11447,N_10859,N_11207);
or U11448 (N_11448,N_10946,N_10983);
nand U11449 (N_11449,N_10934,N_11103);
nand U11450 (N_11450,N_11227,N_11032);
nand U11451 (N_11451,N_10942,N_10911);
or U11452 (N_11452,N_11067,N_11055);
or U11453 (N_11453,N_11266,N_10957);
and U11454 (N_11454,N_10998,N_11333);
and U11455 (N_11455,N_11139,N_11031);
or U11456 (N_11456,N_11144,N_11198);
or U11457 (N_11457,N_11349,N_10929);
nor U11458 (N_11458,N_11285,N_10894);
nor U11459 (N_11459,N_10994,N_11343);
xnor U11460 (N_11460,N_10928,N_11006);
or U11461 (N_11461,N_10975,N_10968);
or U11462 (N_11462,N_11101,N_11359);
nor U11463 (N_11463,N_11143,N_11278);
or U11464 (N_11464,N_10877,N_11126);
nor U11465 (N_11465,N_11217,N_11253);
or U11466 (N_11466,N_11118,N_11378);
and U11467 (N_11467,N_11398,N_11244);
and U11468 (N_11468,N_11355,N_11300);
nand U11469 (N_11469,N_10996,N_11083);
or U11470 (N_11470,N_11140,N_11282);
or U11471 (N_11471,N_11195,N_11129);
nand U11472 (N_11472,N_10811,N_11063);
nand U11473 (N_11473,N_10914,N_11089);
nor U11474 (N_11474,N_11202,N_10997);
nand U11475 (N_11475,N_11232,N_11201);
nor U11476 (N_11476,N_11340,N_11238);
nor U11477 (N_11477,N_10991,N_11135);
xor U11478 (N_11478,N_11149,N_11357);
and U11479 (N_11479,N_11218,N_11296);
nand U11480 (N_11480,N_11279,N_10965);
and U11481 (N_11481,N_11346,N_11381);
nor U11482 (N_11482,N_10947,N_10819);
nor U11483 (N_11483,N_11088,N_10856);
or U11484 (N_11484,N_11231,N_11393);
or U11485 (N_11485,N_11206,N_11016);
xnor U11486 (N_11486,N_11106,N_11337);
or U11487 (N_11487,N_10939,N_11336);
nand U11488 (N_11488,N_11003,N_11113);
nor U11489 (N_11489,N_11192,N_10823);
or U11490 (N_11490,N_11223,N_11384);
xnor U11491 (N_11491,N_11362,N_11081);
nand U11492 (N_11492,N_10814,N_10800);
nand U11493 (N_11493,N_10871,N_10904);
and U11494 (N_11494,N_11110,N_10861);
nor U11495 (N_11495,N_11270,N_10966);
xnor U11496 (N_11496,N_10919,N_11052);
and U11497 (N_11497,N_11159,N_11397);
nand U11498 (N_11498,N_10897,N_10912);
or U11499 (N_11499,N_10921,N_11255);
xnor U11500 (N_11500,N_10972,N_11241);
and U11501 (N_11501,N_11094,N_11001);
or U11502 (N_11502,N_11304,N_11035);
or U11503 (N_11503,N_11387,N_11354);
nor U11504 (N_11504,N_11045,N_11164);
or U11505 (N_11505,N_11289,N_11327);
nand U11506 (N_11506,N_10829,N_11261);
nor U11507 (N_11507,N_11199,N_10801);
or U11508 (N_11508,N_11099,N_11022);
xor U11509 (N_11509,N_10850,N_11328);
nand U11510 (N_11510,N_11248,N_11292);
and U11511 (N_11511,N_11095,N_10831);
and U11512 (N_11512,N_11112,N_11020);
or U11513 (N_11513,N_11386,N_10833);
nor U11514 (N_11514,N_10834,N_10930);
nand U11515 (N_11515,N_11351,N_11062);
and U11516 (N_11516,N_10982,N_11107);
nand U11517 (N_11517,N_11247,N_11146);
or U11518 (N_11518,N_11222,N_10905);
xor U11519 (N_11519,N_11173,N_11272);
or U11520 (N_11520,N_11196,N_10958);
and U11521 (N_11521,N_11047,N_11155);
and U11522 (N_11522,N_10870,N_10967);
or U11523 (N_11523,N_10863,N_11160);
xnor U11524 (N_11524,N_11352,N_11363);
or U11525 (N_11525,N_10810,N_11100);
nor U11526 (N_11526,N_11148,N_11169);
and U11527 (N_11527,N_11115,N_11066);
and U11528 (N_11528,N_10804,N_11392);
or U11529 (N_11529,N_11197,N_10842);
or U11530 (N_11530,N_11007,N_10970);
nand U11531 (N_11531,N_11283,N_11042);
or U11532 (N_11532,N_11040,N_10915);
and U11533 (N_11533,N_11358,N_11152);
and U11534 (N_11534,N_11373,N_11234);
or U11535 (N_11535,N_11273,N_11172);
nand U11536 (N_11536,N_11011,N_10932);
or U11537 (N_11537,N_10881,N_11243);
and U11538 (N_11538,N_11230,N_10895);
nor U11539 (N_11539,N_10969,N_11153);
nand U11540 (N_11540,N_11163,N_11331);
and U11541 (N_11541,N_11281,N_11130);
or U11542 (N_11542,N_10903,N_10926);
or U11543 (N_11543,N_10875,N_10938);
nand U11544 (N_11544,N_10923,N_11077);
or U11545 (N_11545,N_11084,N_11018);
or U11546 (N_11546,N_11096,N_11311);
nor U11547 (N_11547,N_11334,N_11395);
xor U11548 (N_11548,N_11043,N_10990);
nand U11549 (N_11549,N_11391,N_10869);
nor U11550 (N_11550,N_10872,N_11325);
nor U11551 (N_11551,N_10839,N_11254);
nor U11552 (N_11552,N_10978,N_10906);
or U11553 (N_11553,N_11069,N_11382);
and U11554 (N_11554,N_11298,N_11293);
or U11555 (N_11555,N_10852,N_11105);
nand U11556 (N_11556,N_11182,N_11313);
nand U11557 (N_11557,N_10953,N_11330);
xor U11558 (N_11558,N_11318,N_11271);
xor U11559 (N_11559,N_10858,N_10981);
nor U11560 (N_11560,N_11120,N_11051);
and U11561 (N_11561,N_11277,N_11367);
or U11562 (N_11562,N_11246,N_10941);
and U11563 (N_11563,N_11245,N_11229);
and U11564 (N_11564,N_10851,N_10955);
or U11565 (N_11565,N_10836,N_10862);
xor U11566 (N_11566,N_11291,N_10913);
and U11567 (N_11567,N_11301,N_10977);
or U11568 (N_11568,N_10974,N_11133);
and U11569 (N_11569,N_10882,N_11260);
nand U11570 (N_11570,N_10828,N_10937);
xnor U11571 (N_11571,N_11005,N_10951);
and U11572 (N_11572,N_11116,N_11323);
or U11573 (N_11573,N_10807,N_11171);
or U11574 (N_11574,N_11347,N_10848);
xnor U11575 (N_11575,N_11200,N_11122);
and U11576 (N_11576,N_10824,N_11085);
and U11577 (N_11577,N_10980,N_11010);
and U11578 (N_11578,N_11263,N_11117);
nand U11579 (N_11579,N_11262,N_11039);
nand U11580 (N_11580,N_10867,N_11306);
or U11581 (N_11581,N_11075,N_10878);
nand U11582 (N_11582,N_11033,N_10832);
and U11583 (N_11583,N_11380,N_11189);
and U11584 (N_11584,N_11370,N_11136);
xnor U11585 (N_11585,N_11186,N_11239);
or U11586 (N_11586,N_10826,N_10802);
nand U11587 (N_11587,N_11121,N_11134);
or U11588 (N_11588,N_10812,N_11034);
and U11589 (N_11589,N_11335,N_10909);
nor U11590 (N_11590,N_11314,N_11290);
nand U11591 (N_11591,N_11168,N_10973);
nand U11592 (N_11592,N_10846,N_10945);
and U11593 (N_11593,N_11226,N_11124);
nand U11594 (N_11594,N_11050,N_10956);
or U11595 (N_11595,N_11299,N_11276);
and U11596 (N_11596,N_10922,N_11396);
nand U11597 (N_11597,N_11080,N_11017);
or U11598 (N_11598,N_10853,N_11307);
or U11599 (N_11599,N_10992,N_11119);
and U11600 (N_11600,N_11014,N_11321);
and U11601 (N_11601,N_10962,N_10874);
nand U11602 (N_11602,N_11256,N_10813);
or U11603 (N_11603,N_11297,N_11383);
and U11604 (N_11604,N_11210,N_11151);
and U11605 (N_11605,N_11203,N_10963);
or U11606 (N_11606,N_11154,N_11165);
nand U11607 (N_11607,N_10844,N_11215);
nor U11608 (N_11608,N_11021,N_11356);
and U11609 (N_11609,N_11181,N_11086);
or U11610 (N_11610,N_11127,N_10825);
and U11611 (N_11611,N_10806,N_11038);
xnor U11612 (N_11612,N_11079,N_11216);
xor U11613 (N_11613,N_11175,N_11024);
nor U11614 (N_11614,N_11350,N_11390);
nand U11615 (N_11615,N_10890,N_11371);
nor U11616 (N_11616,N_11166,N_10891);
xnor U11617 (N_11617,N_11082,N_11004);
or U11618 (N_11618,N_11183,N_10883);
nand U11619 (N_11619,N_11249,N_10985);
or U11620 (N_11620,N_11109,N_11128);
or U11621 (N_11621,N_10827,N_11000);
or U11622 (N_11622,N_11131,N_10820);
and U11623 (N_11623,N_11369,N_11342);
nand U11624 (N_11624,N_10835,N_11205);
nand U11625 (N_11625,N_11288,N_11338);
or U11626 (N_11626,N_11156,N_10808);
and U11627 (N_11627,N_10860,N_11072);
xor U11628 (N_11628,N_10924,N_11280);
nor U11629 (N_11629,N_11041,N_10857);
nand U11630 (N_11630,N_11303,N_10837);
or U11631 (N_11631,N_11365,N_11320);
and U11632 (N_11632,N_11315,N_10884);
nor U11633 (N_11633,N_11023,N_11310);
or U11634 (N_11634,N_11259,N_11132);
or U11635 (N_11635,N_10936,N_11368);
or U11636 (N_11636,N_11068,N_11076);
and U11637 (N_11637,N_11237,N_10949);
xnor U11638 (N_11638,N_11019,N_10954);
nor U11639 (N_11639,N_11294,N_10976);
or U11640 (N_11640,N_11157,N_11162);
and U11641 (N_11641,N_11048,N_11322);
nor U11642 (N_11642,N_10886,N_10952);
xnor U11643 (N_11643,N_10803,N_10889);
and U11644 (N_11644,N_11036,N_11376);
and U11645 (N_11645,N_11037,N_11399);
and U11646 (N_11646,N_11176,N_11366);
and U11647 (N_11647,N_10971,N_11170);
and U11648 (N_11648,N_11074,N_11284);
or U11649 (N_11649,N_11329,N_10979);
or U11650 (N_11650,N_11316,N_10931);
and U11651 (N_11651,N_11178,N_10950);
and U11652 (N_11652,N_10896,N_11317);
and U11653 (N_11653,N_11044,N_11026);
nor U11654 (N_11654,N_11353,N_11269);
nand U11655 (N_11655,N_11214,N_11360);
or U11656 (N_11656,N_11236,N_11308);
nor U11657 (N_11657,N_11177,N_11070);
nor U11658 (N_11658,N_11187,N_11264);
or U11659 (N_11659,N_11104,N_11389);
or U11660 (N_11660,N_10984,N_11028);
nor U11661 (N_11661,N_10868,N_11108);
nor U11662 (N_11662,N_10864,N_11174);
nor U11663 (N_11663,N_11268,N_10817);
nand U11664 (N_11664,N_11114,N_11053);
nor U11665 (N_11665,N_11147,N_11235);
nor U11666 (N_11666,N_11375,N_11219);
nand U11667 (N_11667,N_10935,N_11009);
and U11668 (N_11668,N_11242,N_10925);
and U11669 (N_11669,N_11265,N_11228);
nand U11670 (N_11670,N_10927,N_10999);
and U11671 (N_11671,N_11220,N_11339);
xnor U11672 (N_11672,N_11145,N_11377);
nor U11673 (N_11673,N_11091,N_10944);
nor U11674 (N_11674,N_10841,N_11309);
or U11675 (N_11675,N_11233,N_11252);
and U11676 (N_11676,N_11190,N_10822);
nor U11677 (N_11677,N_11225,N_10964);
xnor U11678 (N_11678,N_11138,N_10855);
or U11679 (N_11679,N_11204,N_10940);
nor U11680 (N_11680,N_11008,N_11097);
nor U11681 (N_11681,N_11012,N_11275);
xor U11682 (N_11682,N_10893,N_11326);
nor U11683 (N_11683,N_10854,N_11142);
and U11684 (N_11684,N_11388,N_11184);
or U11685 (N_11685,N_10888,N_11188);
xor U11686 (N_11686,N_11073,N_11305);
nand U11687 (N_11687,N_10987,N_11191);
and U11688 (N_11688,N_10830,N_11240);
xor U11689 (N_11689,N_10838,N_10873);
nor U11690 (N_11690,N_11345,N_11250);
nor U11691 (N_11691,N_10910,N_11090);
nand U11692 (N_11692,N_11071,N_10845);
nand U11693 (N_11693,N_11341,N_11257);
nor U11694 (N_11694,N_11374,N_11057);
or U11695 (N_11695,N_10899,N_10849);
nand U11696 (N_11696,N_10805,N_11211);
and U11697 (N_11697,N_11015,N_11212);
nor U11698 (N_11698,N_11267,N_11150);
or U11699 (N_11699,N_11030,N_11049);
and U11700 (N_11700,N_11236,N_11295);
and U11701 (N_11701,N_10815,N_10989);
xnor U11702 (N_11702,N_10998,N_10820);
or U11703 (N_11703,N_11127,N_11011);
and U11704 (N_11704,N_10987,N_11259);
nand U11705 (N_11705,N_11049,N_10979);
and U11706 (N_11706,N_10984,N_11171);
nand U11707 (N_11707,N_10953,N_10950);
nand U11708 (N_11708,N_11276,N_11254);
and U11709 (N_11709,N_11365,N_10805);
and U11710 (N_11710,N_10804,N_11327);
or U11711 (N_11711,N_11259,N_11163);
nand U11712 (N_11712,N_10816,N_11307);
xnor U11713 (N_11713,N_10963,N_11103);
nor U11714 (N_11714,N_11371,N_11151);
nor U11715 (N_11715,N_10843,N_11082);
and U11716 (N_11716,N_10951,N_11060);
and U11717 (N_11717,N_11287,N_11132);
nor U11718 (N_11718,N_10995,N_11021);
or U11719 (N_11719,N_11207,N_10880);
nor U11720 (N_11720,N_11342,N_11258);
or U11721 (N_11721,N_11391,N_10991);
and U11722 (N_11722,N_10870,N_10831);
nand U11723 (N_11723,N_10879,N_11108);
and U11724 (N_11724,N_11094,N_10935);
nand U11725 (N_11725,N_11322,N_11240);
or U11726 (N_11726,N_10966,N_11179);
nor U11727 (N_11727,N_11328,N_11362);
nor U11728 (N_11728,N_10893,N_11262);
nand U11729 (N_11729,N_10825,N_10856);
or U11730 (N_11730,N_11000,N_11323);
or U11731 (N_11731,N_11229,N_11121);
nand U11732 (N_11732,N_11137,N_10881);
nor U11733 (N_11733,N_11018,N_10915);
xor U11734 (N_11734,N_10918,N_11157);
nand U11735 (N_11735,N_10886,N_11080);
xor U11736 (N_11736,N_10865,N_10858);
and U11737 (N_11737,N_10824,N_11292);
and U11738 (N_11738,N_11099,N_11399);
and U11739 (N_11739,N_11292,N_11239);
nand U11740 (N_11740,N_11235,N_11004);
or U11741 (N_11741,N_10920,N_11231);
and U11742 (N_11742,N_11182,N_11358);
or U11743 (N_11743,N_10979,N_11142);
and U11744 (N_11744,N_11355,N_10930);
nand U11745 (N_11745,N_11132,N_11177);
or U11746 (N_11746,N_10827,N_11024);
nand U11747 (N_11747,N_10936,N_11026);
or U11748 (N_11748,N_10821,N_11000);
xnor U11749 (N_11749,N_11168,N_11307);
nand U11750 (N_11750,N_11208,N_11073);
nor U11751 (N_11751,N_10932,N_11348);
nor U11752 (N_11752,N_11328,N_11193);
and U11753 (N_11753,N_11285,N_11170);
nor U11754 (N_11754,N_10990,N_10862);
nor U11755 (N_11755,N_11321,N_11278);
and U11756 (N_11756,N_11286,N_10867);
nand U11757 (N_11757,N_11107,N_11012);
nand U11758 (N_11758,N_10938,N_10908);
or U11759 (N_11759,N_10995,N_11371);
nand U11760 (N_11760,N_10985,N_11081);
and U11761 (N_11761,N_10846,N_11338);
nor U11762 (N_11762,N_11316,N_11083);
xor U11763 (N_11763,N_10859,N_11288);
or U11764 (N_11764,N_11322,N_11226);
and U11765 (N_11765,N_10980,N_11006);
nand U11766 (N_11766,N_10923,N_10947);
nor U11767 (N_11767,N_11191,N_11312);
nor U11768 (N_11768,N_11214,N_10839);
nor U11769 (N_11769,N_10953,N_10921);
and U11770 (N_11770,N_11052,N_11178);
or U11771 (N_11771,N_11349,N_11364);
and U11772 (N_11772,N_10884,N_10931);
nand U11773 (N_11773,N_10852,N_11242);
nand U11774 (N_11774,N_11103,N_11364);
and U11775 (N_11775,N_11134,N_11395);
nand U11776 (N_11776,N_11116,N_11397);
nor U11777 (N_11777,N_10817,N_11041);
nor U11778 (N_11778,N_10890,N_11041);
nor U11779 (N_11779,N_11091,N_11074);
nand U11780 (N_11780,N_11001,N_11076);
and U11781 (N_11781,N_10809,N_10969);
and U11782 (N_11782,N_11178,N_10919);
and U11783 (N_11783,N_10975,N_10905);
or U11784 (N_11784,N_10820,N_10809);
and U11785 (N_11785,N_10912,N_11399);
or U11786 (N_11786,N_10975,N_11152);
nand U11787 (N_11787,N_11356,N_11141);
and U11788 (N_11788,N_11373,N_10832);
nor U11789 (N_11789,N_11314,N_10960);
nand U11790 (N_11790,N_11015,N_11275);
nor U11791 (N_11791,N_10903,N_11012);
xor U11792 (N_11792,N_11122,N_10820);
and U11793 (N_11793,N_10826,N_11064);
nand U11794 (N_11794,N_11290,N_11352);
nor U11795 (N_11795,N_11002,N_11238);
nor U11796 (N_11796,N_10876,N_10899);
nand U11797 (N_11797,N_11255,N_10988);
xnor U11798 (N_11798,N_11318,N_11091);
and U11799 (N_11799,N_11106,N_11237);
and U11800 (N_11800,N_11204,N_11270);
nand U11801 (N_11801,N_10941,N_10903);
or U11802 (N_11802,N_11077,N_11244);
and U11803 (N_11803,N_10876,N_11387);
and U11804 (N_11804,N_10835,N_11377);
or U11805 (N_11805,N_11295,N_11273);
nand U11806 (N_11806,N_11327,N_11033);
nor U11807 (N_11807,N_11369,N_10962);
or U11808 (N_11808,N_10807,N_10864);
nor U11809 (N_11809,N_11192,N_10843);
nor U11810 (N_11810,N_11020,N_11359);
or U11811 (N_11811,N_11038,N_11231);
and U11812 (N_11812,N_11134,N_10803);
nand U11813 (N_11813,N_11208,N_10987);
or U11814 (N_11814,N_11091,N_11286);
or U11815 (N_11815,N_10942,N_11127);
nor U11816 (N_11816,N_11371,N_11225);
and U11817 (N_11817,N_11260,N_10945);
nor U11818 (N_11818,N_11263,N_10998);
nor U11819 (N_11819,N_11294,N_11158);
and U11820 (N_11820,N_11005,N_11058);
and U11821 (N_11821,N_10919,N_11398);
nand U11822 (N_11822,N_11073,N_10939);
nor U11823 (N_11823,N_11155,N_11027);
nand U11824 (N_11824,N_11000,N_11383);
or U11825 (N_11825,N_10906,N_11342);
nor U11826 (N_11826,N_10843,N_11311);
nor U11827 (N_11827,N_10984,N_11238);
nand U11828 (N_11828,N_11301,N_11346);
nor U11829 (N_11829,N_10928,N_11299);
nor U11830 (N_11830,N_11111,N_11303);
nand U11831 (N_11831,N_11003,N_11356);
or U11832 (N_11832,N_10956,N_11395);
and U11833 (N_11833,N_11231,N_11353);
and U11834 (N_11834,N_11306,N_11155);
xor U11835 (N_11835,N_10833,N_11050);
nor U11836 (N_11836,N_10800,N_11023);
or U11837 (N_11837,N_11130,N_11233);
nand U11838 (N_11838,N_10966,N_11382);
nor U11839 (N_11839,N_10976,N_11361);
and U11840 (N_11840,N_10874,N_11197);
nand U11841 (N_11841,N_10971,N_11343);
nand U11842 (N_11842,N_11223,N_11244);
xor U11843 (N_11843,N_10875,N_11273);
nor U11844 (N_11844,N_10956,N_11318);
and U11845 (N_11845,N_11176,N_10893);
nand U11846 (N_11846,N_10889,N_11288);
nand U11847 (N_11847,N_11279,N_11334);
nor U11848 (N_11848,N_11319,N_11006);
nand U11849 (N_11849,N_11293,N_10963);
xor U11850 (N_11850,N_10925,N_11361);
and U11851 (N_11851,N_10969,N_11012);
nand U11852 (N_11852,N_11139,N_11018);
xnor U11853 (N_11853,N_11236,N_10931);
nor U11854 (N_11854,N_11385,N_10926);
nand U11855 (N_11855,N_10970,N_11109);
nand U11856 (N_11856,N_11258,N_10909);
or U11857 (N_11857,N_11273,N_11036);
nand U11858 (N_11858,N_11073,N_10976);
nor U11859 (N_11859,N_11026,N_11134);
nand U11860 (N_11860,N_10885,N_11069);
nand U11861 (N_11861,N_11003,N_11120);
or U11862 (N_11862,N_11112,N_11386);
and U11863 (N_11863,N_10901,N_11298);
nor U11864 (N_11864,N_11090,N_10914);
xnor U11865 (N_11865,N_11335,N_10873);
nor U11866 (N_11866,N_11078,N_11369);
nand U11867 (N_11867,N_11163,N_10918);
or U11868 (N_11868,N_10881,N_10911);
xnor U11869 (N_11869,N_11025,N_10898);
and U11870 (N_11870,N_11114,N_10907);
or U11871 (N_11871,N_10851,N_10840);
nor U11872 (N_11872,N_11164,N_10829);
nand U11873 (N_11873,N_11203,N_11211);
nor U11874 (N_11874,N_11113,N_10999);
and U11875 (N_11875,N_10905,N_11121);
or U11876 (N_11876,N_11180,N_11253);
nor U11877 (N_11877,N_10888,N_10827);
nand U11878 (N_11878,N_10954,N_11349);
nor U11879 (N_11879,N_11214,N_11040);
nor U11880 (N_11880,N_11394,N_10865);
xor U11881 (N_11881,N_10998,N_11038);
or U11882 (N_11882,N_11289,N_11326);
xnor U11883 (N_11883,N_11222,N_11041);
xor U11884 (N_11884,N_11284,N_11228);
or U11885 (N_11885,N_11229,N_10950);
or U11886 (N_11886,N_11122,N_11309);
nor U11887 (N_11887,N_10929,N_10803);
or U11888 (N_11888,N_11020,N_10962);
and U11889 (N_11889,N_11316,N_10904);
and U11890 (N_11890,N_11042,N_10804);
nor U11891 (N_11891,N_11223,N_11089);
xnor U11892 (N_11892,N_10808,N_10886);
and U11893 (N_11893,N_11161,N_10834);
nor U11894 (N_11894,N_11043,N_10816);
or U11895 (N_11895,N_10958,N_11181);
and U11896 (N_11896,N_11323,N_10911);
xor U11897 (N_11897,N_11394,N_11170);
or U11898 (N_11898,N_10936,N_11297);
or U11899 (N_11899,N_10939,N_11079);
nor U11900 (N_11900,N_10997,N_11304);
or U11901 (N_11901,N_10952,N_11106);
nand U11902 (N_11902,N_11383,N_10886);
or U11903 (N_11903,N_10848,N_10965);
nand U11904 (N_11904,N_11026,N_11365);
nor U11905 (N_11905,N_11103,N_11396);
or U11906 (N_11906,N_11174,N_11188);
nor U11907 (N_11907,N_11305,N_11035);
nand U11908 (N_11908,N_10893,N_10811);
nand U11909 (N_11909,N_11276,N_11279);
nand U11910 (N_11910,N_11314,N_11096);
nand U11911 (N_11911,N_11224,N_11061);
and U11912 (N_11912,N_11104,N_10876);
xnor U11913 (N_11913,N_11123,N_11256);
or U11914 (N_11914,N_11369,N_11304);
and U11915 (N_11915,N_11037,N_11386);
or U11916 (N_11916,N_11213,N_10859);
nor U11917 (N_11917,N_10939,N_10956);
or U11918 (N_11918,N_11193,N_11201);
xnor U11919 (N_11919,N_10979,N_11261);
or U11920 (N_11920,N_11095,N_11268);
and U11921 (N_11921,N_11244,N_11213);
and U11922 (N_11922,N_10815,N_11332);
nand U11923 (N_11923,N_11350,N_11364);
and U11924 (N_11924,N_11020,N_11398);
nand U11925 (N_11925,N_11083,N_10988);
nor U11926 (N_11926,N_11090,N_11036);
nor U11927 (N_11927,N_10879,N_11054);
nor U11928 (N_11928,N_11270,N_10874);
and U11929 (N_11929,N_10861,N_10874);
nand U11930 (N_11930,N_11200,N_10885);
nor U11931 (N_11931,N_10928,N_11107);
and U11932 (N_11932,N_10994,N_10858);
nand U11933 (N_11933,N_11175,N_11205);
nand U11934 (N_11934,N_11300,N_11157);
nand U11935 (N_11935,N_11274,N_11131);
nand U11936 (N_11936,N_10947,N_11149);
nor U11937 (N_11937,N_11155,N_11000);
xnor U11938 (N_11938,N_11135,N_11103);
or U11939 (N_11939,N_10957,N_11301);
and U11940 (N_11940,N_10869,N_11120);
or U11941 (N_11941,N_11287,N_11046);
and U11942 (N_11942,N_11359,N_11292);
and U11943 (N_11943,N_10813,N_11132);
or U11944 (N_11944,N_11263,N_11286);
or U11945 (N_11945,N_11325,N_11021);
nand U11946 (N_11946,N_10827,N_11107);
nand U11947 (N_11947,N_11211,N_10830);
nand U11948 (N_11948,N_11239,N_10909);
and U11949 (N_11949,N_11011,N_11082);
or U11950 (N_11950,N_11176,N_11149);
and U11951 (N_11951,N_11034,N_10835);
or U11952 (N_11952,N_11233,N_10932);
and U11953 (N_11953,N_11136,N_11160);
or U11954 (N_11954,N_10901,N_10930);
nor U11955 (N_11955,N_11310,N_10889);
and U11956 (N_11956,N_11089,N_11310);
nor U11957 (N_11957,N_11350,N_11175);
nand U11958 (N_11958,N_11269,N_10843);
and U11959 (N_11959,N_11372,N_11186);
and U11960 (N_11960,N_11103,N_11138);
or U11961 (N_11961,N_10915,N_11111);
or U11962 (N_11962,N_10991,N_11392);
and U11963 (N_11963,N_11064,N_11000);
nor U11964 (N_11964,N_11121,N_11267);
or U11965 (N_11965,N_10842,N_11361);
and U11966 (N_11966,N_10934,N_10959);
nor U11967 (N_11967,N_11093,N_11090);
and U11968 (N_11968,N_11108,N_11229);
and U11969 (N_11969,N_10947,N_10830);
and U11970 (N_11970,N_11004,N_11272);
nor U11971 (N_11971,N_10872,N_10825);
nor U11972 (N_11972,N_11213,N_11154);
nor U11973 (N_11973,N_11194,N_10857);
and U11974 (N_11974,N_10948,N_11039);
xnor U11975 (N_11975,N_11211,N_11019);
or U11976 (N_11976,N_11016,N_11028);
and U11977 (N_11977,N_11132,N_11089);
and U11978 (N_11978,N_11204,N_11198);
or U11979 (N_11979,N_11059,N_10968);
and U11980 (N_11980,N_11192,N_11285);
nand U11981 (N_11981,N_11134,N_10944);
and U11982 (N_11982,N_11044,N_11167);
nor U11983 (N_11983,N_11292,N_11356);
xnor U11984 (N_11984,N_11370,N_11120);
nand U11985 (N_11985,N_11237,N_10840);
nand U11986 (N_11986,N_11169,N_10930);
and U11987 (N_11987,N_11088,N_11008);
or U11988 (N_11988,N_11347,N_11241);
nand U11989 (N_11989,N_11157,N_11166);
or U11990 (N_11990,N_11134,N_10919);
or U11991 (N_11991,N_11241,N_11103);
or U11992 (N_11992,N_11161,N_11052);
or U11993 (N_11993,N_11365,N_10853);
or U11994 (N_11994,N_11339,N_11271);
xnor U11995 (N_11995,N_11086,N_11126);
nand U11996 (N_11996,N_10833,N_10921);
and U11997 (N_11997,N_11091,N_11322);
and U11998 (N_11998,N_10929,N_10908);
nand U11999 (N_11999,N_10880,N_11326);
nor U12000 (N_12000,N_11680,N_11962);
and U12001 (N_12001,N_11946,N_11665);
nand U12002 (N_12002,N_11560,N_11501);
or U12003 (N_12003,N_11416,N_11589);
and U12004 (N_12004,N_11704,N_11664);
nor U12005 (N_12005,N_11497,N_11420);
nor U12006 (N_12006,N_11462,N_11676);
nor U12007 (N_12007,N_11949,N_11641);
xor U12008 (N_12008,N_11604,N_11563);
and U12009 (N_12009,N_11469,N_11580);
xnor U12010 (N_12010,N_11649,N_11774);
nor U12011 (N_12011,N_11653,N_11490);
and U12012 (N_12012,N_11900,N_11833);
nor U12013 (N_12013,N_11619,N_11481);
nor U12014 (N_12014,N_11724,N_11617);
or U12015 (N_12015,N_11922,N_11824);
nor U12016 (N_12016,N_11738,N_11981);
and U12017 (N_12017,N_11628,N_11867);
xor U12018 (N_12018,N_11770,N_11899);
nand U12019 (N_12019,N_11422,N_11412);
nor U12020 (N_12020,N_11575,N_11541);
nor U12021 (N_12021,N_11647,N_11418);
nand U12022 (N_12022,N_11532,N_11616);
and U12023 (N_12023,N_11817,N_11950);
nand U12024 (N_12024,N_11531,N_11546);
xor U12025 (N_12025,N_11703,N_11702);
nor U12026 (N_12026,N_11593,N_11442);
xor U12027 (N_12027,N_11947,N_11999);
and U12028 (N_12028,N_11431,N_11594);
nand U12029 (N_12029,N_11956,N_11727);
or U12030 (N_12030,N_11712,N_11449);
nor U12031 (N_12031,N_11830,N_11719);
and U12032 (N_12032,N_11916,N_11600);
or U12033 (N_12033,N_11540,N_11809);
and U12034 (N_12034,N_11735,N_11974);
and U12035 (N_12035,N_11843,N_11569);
and U12036 (N_12036,N_11706,N_11944);
nand U12037 (N_12037,N_11829,N_11610);
or U12038 (N_12038,N_11714,N_11476);
nand U12039 (N_12039,N_11739,N_11957);
or U12040 (N_12040,N_11749,N_11646);
nor U12041 (N_12041,N_11761,N_11777);
nor U12042 (N_12042,N_11440,N_11545);
or U12043 (N_12043,N_11517,N_11447);
nand U12044 (N_12044,N_11758,N_11623);
or U12045 (N_12045,N_11984,N_11556);
and U12046 (N_12046,N_11640,N_11669);
nand U12047 (N_12047,N_11652,N_11692);
or U12048 (N_12048,N_11553,N_11891);
nand U12049 (N_12049,N_11784,N_11686);
nor U12050 (N_12050,N_11723,N_11812);
or U12051 (N_12051,N_11868,N_11675);
or U12052 (N_12052,N_11695,N_11880);
nor U12053 (N_12053,N_11499,N_11919);
nand U12054 (N_12054,N_11456,N_11662);
and U12055 (N_12055,N_11544,N_11608);
or U12056 (N_12056,N_11612,N_11760);
xnor U12057 (N_12057,N_11658,N_11525);
nand U12058 (N_12058,N_11504,N_11907);
xnor U12059 (N_12059,N_11890,N_11659);
nand U12060 (N_12060,N_11808,N_11883);
nand U12061 (N_12061,N_11898,N_11786);
nand U12062 (N_12062,N_11578,N_11762);
nand U12063 (N_12063,N_11684,N_11559);
xnor U12064 (N_12064,N_11666,N_11987);
nand U12065 (N_12065,N_11415,N_11773);
nand U12066 (N_12066,N_11794,N_11534);
nand U12067 (N_12067,N_11421,N_11783);
and U12068 (N_12068,N_11795,N_11607);
nor U12069 (N_12069,N_11953,N_11926);
nand U12070 (N_12070,N_11690,N_11861);
and U12071 (N_12071,N_11570,N_11820);
or U12072 (N_12072,N_11862,N_11561);
nor U12073 (N_12073,N_11764,N_11535);
nor U12074 (N_12074,N_11838,N_11400);
and U12075 (N_12075,N_11627,N_11805);
nand U12076 (N_12076,N_11423,N_11876);
nand U12077 (N_12077,N_11878,N_11800);
nor U12078 (N_12078,N_11753,N_11509);
xor U12079 (N_12079,N_11537,N_11973);
and U12080 (N_12080,N_11603,N_11539);
nand U12081 (N_12081,N_11840,N_11920);
and U12082 (N_12082,N_11458,N_11495);
or U12083 (N_12083,N_11419,N_11661);
and U12084 (N_12084,N_11657,N_11466);
and U12085 (N_12085,N_11624,N_11547);
nand U12086 (N_12086,N_11485,N_11810);
and U12087 (N_12087,N_11970,N_11637);
nor U12088 (N_12088,N_11611,N_11551);
and U12089 (N_12089,N_11598,N_11945);
nand U12090 (N_12090,N_11498,N_11799);
nand U12091 (N_12091,N_11752,N_11976);
nor U12092 (N_12092,N_11983,N_11825);
nor U12093 (N_12093,N_11663,N_11564);
nand U12094 (N_12094,N_11672,N_11912);
and U12095 (N_12095,N_11814,N_11679);
and U12096 (N_12096,N_11816,N_11965);
and U12097 (N_12097,N_11555,N_11884);
or U12098 (N_12098,N_11631,N_11474);
nor U12099 (N_12099,N_11635,N_11767);
and U12100 (N_12100,N_11668,N_11917);
nand U12101 (N_12101,N_11896,N_11892);
and U12102 (N_12102,N_11938,N_11996);
and U12103 (N_12103,N_11413,N_11590);
xor U12104 (N_12104,N_11461,N_11971);
xnor U12105 (N_12105,N_11697,N_11444);
nand U12106 (N_12106,N_11903,N_11656);
xor U12107 (N_12107,N_11885,N_11813);
and U12108 (N_12108,N_11491,N_11518);
or U12109 (N_12109,N_11549,N_11626);
nand U12110 (N_12110,N_11568,N_11595);
or U12111 (N_12111,N_11685,N_11873);
and U12112 (N_12112,N_11828,N_11855);
nand U12113 (N_12113,N_11853,N_11417);
and U12114 (N_12114,N_11448,N_11857);
and U12115 (N_12115,N_11879,N_11565);
nand U12116 (N_12116,N_11599,N_11745);
xnor U12117 (N_12117,N_11503,N_11645);
and U12118 (N_12118,N_11660,N_11487);
or U12119 (N_12119,N_11486,N_11914);
nand U12120 (N_12120,N_11506,N_11542);
nor U12121 (N_12121,N_11835,N_11975);
and U12122 (N_12122,N_11798,N_11730);
nor U12123 (N_12123,N_11582,N_11615);
xnor U12124 (N_12124,N_11988,N_11522);
nor U12125 (N_12125,N_11927,N_11923);
or U12126 (N_12126,N_11797,N_11682);
xor U12127 (N_12127,N_11577,N_11841);
nand U12128 (N_12128,N_11769,N_11948);
xor U12129 (N_12129,N_11865,N_11404);
nor U12130 (N_12130,N_11587,N_11740);
xor U12131 (N_12131,N_11915,N_11677);
nand U12132 (N_12132,N_11633,N_11543);
and U12133 (N_12133,N_11614,N_11583);
and U12134 (N_12134,N_11781,N_11602);
and U12135 (N_12135,N_11477,N_11750);
or U12136 (N_12136,N_11964,N_11882);
nand U12137 (N_12137,N_11854,N_11952);
and U12138 (N_12138,N_11478,N_11674);
nand U12139 (N_12139,N_11699,N_11910);
and U12140 (N_12140,N_11832,N_11457);
nand U12141 (N_12141,N_11573,N_11893);
nor U12142 (N_12142,N_11844,N_11407);
and U12143 (N_12143,N_11791,N_11822);
and U12144 (N_12144,N_11597,N_11521);
nor U12145 (N_12145,N_11966,N_11566);
and U12146 (N_12146,N_11642,N_11827);
xnor U12147 (N_12147,N_11698,N_11480);
nand U12148 (N_12148,N_11776,N_11718);
nor U12149 (N_12149,N_11622,N_11918);
nor U12150 (N_12150,N_11567,N_11789);
nor U12151 (N_12151,N_11992,N_11778);
nor U12152 (N_12152,N_11801,N_11572);
and U12153 (N_12153,N_11629,N_11989);
or U12154 (N_12154,N_11870,N_11494);
nor U12155 (N_12155,N_11508,N_11639);
or U12156 (N_12156,N_11405,N_11694);
and U12157 (N_12157,N_11823,N_11925);
nor U12158 (N_12158,N_11632,N_11995);
or U12159 (N_12159,N_11414,N_11515);
or U12160 (N_12160,N_11860,N_11606);
nor U12161 (N_12161,N_11455,N_11863);
or U12162 (N_12162,N_11401,N_11529);
xor U12163 (N_12163,N_11500,N_11467);
and U12164 (N_12164,N_11759,N_11874);
and U12165 (N_12165,N_11856,N_11681);
nand U12166 (N_12166,N_11450,N_11887);
nand U12167 (N_12167,N_11426,N_11731);
nor U12168 (N_12168,N_11492,N_11691);
or U12169 (N_12169,N_11831,N_11479);
or U12170 (N_12170,N_11687,N_11725);
or U12171 (N_12171,N_11678,N_11715);
or U12172 (N_12172,N_11630,N_11852);
nor U12173 (N_12173,N_11746,N_11889);
or U12174 (N_12174,N_11470,N_11696);
nor U12175 (N_12175,N_11772,N_11650);
and U12176 (N_12176,N_11402,N_11963);
nand U12177 (N_12177,N_11493,N_11780);
nor U12178 (N_12178,N_11768,N_11836);
xnor U12179 (N_12179,N_11756,N_11941);
nand U12180 (N_12180,N_11667,N_11787);
nand U12181 (N_12181,N_11558,N_11807);
or U12182 (N_12182,N_11848,N_11516);
nand U12183 (N_12183,N_11460,N_11707);
nand U12184 (N_12184,N_11908,N_11864);
or U12185 (N_12185,N_11804,N_11519);
nor U12186 (N_12186,N_11958,N_11708);
nor U12187 (N_12187,N_11489,N_11453);
nand U12188 (N_12188,N_11837,N_11913);
or U12189 (N_12189,N_11788,N_11755);
nand U12190 (N_12190,N_11819,N_11654);
xnor U12191 (N_12191,N_11871,N_11536);
nand U12192 (N_12192,N_11550,N_11557);
or U12193 (N_12193,N_11562,N_11451);
and U12194 (N_12194,N_11729,N_11728);
and U12195 (N_12195,N_11574,N_11530);
nor U12196 (N_12196,N_11961,N_11634);
and U12197 (N_12197,N_11937,N_11432);
xor U12198 (N_12198,N_11901,N_11811);
or U12199 (N_12199,N_11886,N_11584);
and U12200 (N_12200,N_11998,N_11511);
nand U12201 (N_12201,N_11700,N_11775);
or U12202 (N_12202,N_11960,N_11748);
nand U12203 (N_12203,N_11904,N_11932);
xnor U12204 (N_12204,N_11842,N_11510);
nand U12205 (N_12205,N_11717,N_11977);
nand U12206 (N_12206,N_11496,N_11552);
or U12207 (N_12207,N_11505,N_11834);
and U12208 (N_12208,N_11881,N_11726);
or U12209 (N_12209,N_11513,N_11428);
nor U12210 (N_12210,N_11482,N_11403);
and U12211 (N_12211,N_11721,N_11994);
nand U12212 (N_12212,N_11921,N_11894);
or U12213 (N_12213,N_11931,N_11528);
nor U12214 (N_12214,N_11747,N_11651);
nor U12215 (N_12215,N_11483,N_11710);
or U12216 (N_12216,N_11571,N_11826);
nor U12217 (N_12217,N_11512,N_11736);
nand U12218 (N_12218,N_11982,N_11644);
nor U12219 (N_12219,N_11928,N_11782);
and U12220 (N_12220,N_11934,N_11845);
nor U12221 (N_12221,N_11688,N_11588);
or U12222 (N_12222,N_11576,N_11978);
xnor U12223 (N_12223,N_11514,N_11954);
nand U12224 (N_12224,N_11411,N_11765);
xor U12225 (N_12225,N_11524,N_11548);
and U12226 (N_12226,N_11427,N_11406);
xnor U12227 (N_12227,N_11713,N_11648);
nor U12228 (N_12228,N_11452,N_11625);
nand U12229 (N_12229,N_11897,N_11754);
nor U12230 (N_12230,N_11930,N_11579);
nor U12231 (N_12231,N_11409,N_11858);
nor U12232 (N_12232,N_11935,N_11859);
xnor U12233 (N_12233,N_11790,N_11502);
nand U12234 (N_12234,N_11991,N_11888);
xor U12235 (N_12235,N_11596,N_11803);
nor U12236 (N_12236,N_11554,N_11929);
nand U12237 (N_12237,N_11875,N_11671);
nor U12238 (N_12238,N_11818,N_11851);
nand U12239 (N_12239,N_11895,N_11673);
or U12240 (N_12240,N_11463,N_11429);
nand U12241 (N_12241,N_11969,N_11716);
xnor U12242 (N_12242,N_11720,N_11849);
or U12243 (N_12243,N_11951,N_11711);
nor U12244 (N_12244,N_11586,N_11742);
and U12245 (N_12245,N_11472,N_11655);
or U12246 (N_12246,N_11410,N_11939);
and U12247 (N_12247,N_11737,N_11943);
nand U12248 (N_12248,N_11846,N_11520);
or U12249 (N_12249,N_11990,N_11538);
or U12250 (N_12250,N_11445,N_11940);
xnor U12251 (N_12251,N_11959,N_11705);
nor U12252 (N_12252,N_11744,N_11437);
nand U12253 (N_12253,N_11446,N_11683);
or U12254 (N_12254,N_11454,N_11609);
and U12255 (N_12255,N_11592,N_11585);
nor U12256 (N_12256,N_11526,N_11613);
nor U12257 (N_12257,N_11701,N_11909);
or U12258 (N_12258,N_11936,N_11847);
nor U12259 (N_12259,N_11839,N_11821);
nor U12260 (N_12260,N_11425,N_11733);
or U12261 (N_12261,N_11986,N_11638);
or U12262 (N_12262,N_11605,N_11689);
nor U12263 (N_12263,N_11751,N_11979);
and U12264 (N_12264,N_11424,N_11763);
nor U12265 (N_12265,N_11473,N_11471);
nand U12266 (N_12266,N_11796,N_11993);
nand U12267 (N_12267,N_11443,N_11527);
and U12268 (N_12268,N_11933,N_11877);
nand U12269 (N_12269,N_11967,N_11793);
xnor U12270 (N_12270,N_11997,N_11743);
and U12271 (N_12271,N_11872,N_11866);
nor U12272 (N_12272,N_11766,N_11621);
nand U12273 (N_12273,N_11815,N_11581);
and U12274 (N_12274,N_11732,N_11488);
nor U12275 (N_12275,N_11924,N_11771);
nand U12276 (N_12276,N_11670,N_11618);
nand U12277 (N_12277,N_11806,N_11968);
nand U12278 (N_12278,N_11792,N_11433);
nor U12279 (N_12279,N_11533,N_11408);
and U12280 (N_12280,N_11464,N_11785);
and U12281 (N_12281,N_11475,N_11906);
nor U12282 (N_12282,N_11434,N_11734);
xor U12283 (N_12283,N_11523,N_11902);
and U12284 (N_12284,N_11980,N_11438);
xnor U12285 (N_12285,N_11972,N_11591);
and U12286 (N_12286,N_11869,N_11905);
or U12287 (N_12287,N_11436,N_11911);
or U12288 (N_12288,N_11430,N_11779);
or U12289 (N_12289,N_11484,N_11620);
or U12290 (N_12290,N_11942,N_11636);
nand U12291 (N_12291,N_11507,N_11643);
nand U12292 (N_12292,N_11802,N_11985);
nor U12293 (N_12293,N_11850,N_11441);
nor U12294 (N_12294,N_11439,N_11601);
nor U12295 (N_12295,N_11465,N_11741);
nor U12296 (N_12296,N_11468,N_11435);
and U12297 (N_12297,N_11722,N_11709);
nand U12298 (N_12298,N_11693,N_11459);
or U12299 (N_12299,N_11955,N_11757);
and U12300 (N_12300,N_11907,N_11649);
nor U12301 (N_12301,N_11527,N_11722);
nor U12302 (N_12302,N_11487,N_11627);
nor U12303 (N_12303,N_11956,N_11986);
or U12304 (N_12304,N_11647,N_11632);
or U12305 (N_12305,N_11959,N_11586);
or U12306 (N_12306,N_11749,N_11436);
or U12307 (N_12307,N_11550,N_11821);
nor U12308 (N_12308,N_11417,N_11983);
nor U12309 (N_12309,N_11917,N_11972);
nor U12310 (N_12310,N_11651,N_11483);
nand U12311 (N_12311,N_11816,N_11930);
xnor U12312 (N_12312,N_11933,N_11649);
nor U12313 (N_12313,N_11873,N_11983);
or U12314 (N_12314,N_11631,N_11945);
nor U12315 (N_12315,N_11902,N_11597);
nor U12316 (N_12316,N_11575,N_11989);
and U12317 (N_12317,N_11672,N_11614);
and U12318 (N_12318,N_11803,N_11807);
and U12319 (N_12319,N_11813,N_11404);
nand U12320 (N_12320,N_11528,N_11930);
or U12321 (N_12321,N_11405,N_11669);
and U12322 (N_12322,N_11616,N_11988);
and U12323 (N_12323,N_11954,N_11703);
nor U12324 (N_12324,N_11485,N_11926);
and U12325 (N_12325,N_11775,N_11952);
nor U12326 (N_12326,N_11932,N_11717);
and U12327 (N_12327,N_11673,N_11884);
xnor U12328 (N_12328,N_11710,N_11784);
and U12329 (N_12329,N_11548,N_11732);
xor U12330 (N_12330,N_11964,N_11435);
nand U12331 (N_12331,N_11418,N_11525);
nor U12332 (N_12332,N_11401,N_11717);
and U12333 (N_12333,N_11647,N_11556);
or U12334 (N_12334,N_11446,N_11591);
xor U12335 (N_12335,N_11451,N_11888);
nor U12336 (N_12336,N_11646,N_11654);
xor U12337 (N_12337,N_11499,N_11588);
nand U12338 (N_12338,N_11642,N_11985);
xnor U12339 (N_12339,N_11716,N_11448);
and U12340 (N_12340,N_11893,N_11524);
xnor U12341 (N_12341,N_11687,N_11680);
nor U12342 (N_12342,N_11619,N_11741);
nand U12343 (N_12343,N_11984,N_11964);
nand U12344 (N_12344,N_11840,N_11730);
and U12345 (N_12345,N_11545,N_11604);
nor U12346 (N_12346,N_11787,N_11864);
xnor U12347 (N_12347,N_11912,N_11534);
and U12348 (N_12348,N_11786,N_11744);
nand U12349 (N_12349,N_11592,N_11449);
and U12350 (N_12350,N_11446,N_11827);
nand U12351 (N_12351,N_11505,N_11683);
or U12352 (N_12352,N_11413,N_11614);
nor U12353 (N_12353,N_11900,N_11782);
and U12354 (N_12354,N_11855,N_11512);
nor U12355 (N_12355,N_11443,N_11415);
nor U12356 (N_12356,N_11960,N_11528);
or U12357 (N_12357,N_11949,N_11562);
and U12358 (N_12358,N_11905,N_11703);
nor U12359 (N_12359,N_11613,N_11451);
xor U12360 (N_12360,N_11412,N_11631);
nand U12361 (N_12361,N_11651,N_11488);
or U12362 (N_12362,N_11777,N_11624);
nor U12363 (N_12363,N_11880,N_11453);
nor U12364 (N_12364,N_11781,N_11437);
nor U12365 (N_12365,N_11783,N_11664);
xor U12366 (N_12366,N_11839,N_11910);
xor U12367 (N_12367,N_11572,N_11551);
and U12368 (N_12368,N_11515,N_11687);
xnor U12369 (N_12369,N_11611,N_11903);
or U12370 (N_12370,N_11475,N_11749);
nor U12371 (N_12371,N_11742,N_11713);
nor U12372 (N_12372,N_11897,N_11566);
xor U12373 (N_12373,N_11675,N_11612);
nand U12374 (N_12374,N_11971,N_11451);
nor U12375 (N_12375,N_11490,N_11745);
nor U12376 (N_12376,N_11688,N_11805);
nor U12377 (N_12377,N_11509,N_11825);
nand U12378 (N_12378,N_11764,N_11708);
nor U12379 (N_12379,N_11952,N_11763);
nand U12380 (N_12380,N_11892,N_11929);
xor U12381 (N_12381,N_11426,N_11982);
or U12382 (N_12382,N_11547,N_11445);
nor U12383 (N_12383,N_11403,N_11924);
nor U12384 (N_12384,N_11983,N_11998);
and U12385 (N_12385,N_11534,N_11862);
nand U12386 (N_12386,N_11781,N_11612);
and U12387 (N_12387,N_11599,N_11910);
and U12388 (N_12388,N_11724,N_11919);
and U12389 (N_12389,N_11775,N_11918);
or U12390 (N_12390,N_11739,N_11801);
nor U12391 (N_12391,N_11662,N_11472);
and U12392 (N_12392,N_11525,N_11690);
or U12393 (N_12393,N_11818,N_11998);
nand U12394 (N_12394,N_11781,N_11549);
nor U12395 (N_12395,N_11873,N_11862);
and U12396 (N_12396,N_11630,N_11706);
or U12397 (N_12397,N_11969,N_11533);
nand U12398 (N_12398,N_11719,N_11550);
or U12399 (N_12399,N_11409,N_11745);
and U12400 (N_12400,N_11960,N_11716);
nand U12401 (N_12401,N_11454,N_11853);
nand U12402 (N_12402,N_11866,N_11561);
nand U12403 (N_12403,N_11540,N_11676);
and U12404 (N_12404,N_11441,N_11960);
and U12405 (N_12405,N_11908,N_11698);
and U12406 (N_12406,N_11400,N_11839);
nand U12407 (N_12407,N_11701,N_11523);
and U12408 (N_12408,N_11976,N_11957);
or U12409 (N_12409,N_11938,N_11649);
or U12410 (N_12410,N_11474,N_11514);
or U12411 (N_12411,N_11869,N_11743);
nor U12412 (N_12412,N_11731,N_11803);
or U12413 (N_12413,N_11678,N_11653);
nand U12414 (N_12414,N_11975,N_11545);
nand U12415 (N_12415,N_11602,N_11712);
and U12416 (N_12416,N_11597,N_11911);
xnor U12417 (N_12417,N_11594,N_11465);
nand U12418 (N_12418,N_11884,N_11640);
or U12419 (N_12419,N_11863,N_11972);
nor U12420 (N_12420,N_11810,N_11611);
nor U12421 (N_12421,N_11662,N_11872);
and U12422 (N_12422,N_11406,N_11834);
nand U12423 (N_12423,N_11717,N_11816);
nor U12424 (N_12424,N_11618,N_11602);
xnor U12425 (N_12425,N_11589,N_11478);
xor U12426 (N_12426,N_11704,N_11870);
nand U12427 (N_12427,N_11857,N_11693);
xor U12428 (N_12428,N_11660,N_11954);
nor U12429 (N_12429,N_11426,N_11767);
nand U12430 (N_12430,N_11959,N_11631);
nor U12431 (N_12431,N_11811,N_11543);
nand U12432 (N_12432,N_11641,N_11640);
nand U12433 (N_12433,N_11909,N_11768);
nor U12434 (N_12434,N_11830,N_11951);
nor U12435 (N_12435,N_11724,N_11846);
or U12436 (N_12436,N_11616,N_11438);
nor U12437 (N_12437,N_11567,N_11916);
or U12438 (N_12438,N_11510,N_11430);
or U12439 (N_12439,N_11754,N_11634);
xnor U12440 (N_12440,N_11801,N_11890);
and U12441 (N_12441,N_11877,N_11789);
xor U12442 (N_12442,N_11691,N_11858);
and U12443 (N_12443,N_11779,N_11618);
or U12444 (N_12444,N_11965,N_11876);
and U12445 (N_12445,N_11467,N_11649);
nor U12446 (N_12446,N_11852,N_11550);
and U12447 (N_12447,N_11892,N_11566);
and U12448 (N_12448,N_11434,N_11664);
and U12449 (N_12449,N_11950,N_11947);
nand U12450 (N_12450,N_11933,N_11589);
or U12451 (N_12451,N_11812,N_11407);
or U12452 (N_12452,N_11823,N_11557);
nor U12453 (N_12453,N_11810,N_11992);
and U12454 (N_12454,N_11716,N_11490);
nand U12455 (N_12455,N_11797,N_11619);
and U12456 (N_12456,N_11700,N_11778);
or U12457 (N_12457,N_11922,N_11456);
and U12458 (N_12458,N_11776,N_11970);
nand U12459 (N_12459,N_11573,N_11422);
and U12460 (N_12460,N_11836,N_11547);
and U12461 (N_12461,N_11991,N_11707);
nor U12462 (N_12462,N_11472,N_11417);
nor U12463 (N_12463,N_11466,N_11969);
nor U12464 (N_12464,N_11653,N_11729);
xor U12465 (N_12465,N_11434,N_11880);
xnor U12466 (N_12466,N_11805,N_11741);
nand U12467 (N_12467,N_11565,N_11585);
nand U12468 (N_12468,N_11649,N_11986);
and U12469 (N_12469,N_11962,N_11775);
xnor U12470 (N_12470,N_11714,N_11751);
nand U12471 (N_12471,N_11608,N_11407);
nand U12472 (N_12472,N_11777,N_11430);
nand U12473 (N_12473,N_11433,N_11938);
nand U12474 (N_12474,N_11465,N_11539);
or U12475 (N_12475,N_11882,N_11459);
or U12476 (N_12476,N_11887,N_11856);
or U12477 (N_12477,N_11920,N_11553);
nor U12478 (N_12478,N_11844,N_11470);
or U12479 (N_12479,N_11401,N_11742);
nand U12480 (N_12480,N_11732,N_11701);
nand U12481 (N_12481,N_11488,N_11795);
and U12482 (N_12482,N_11910,N_11529);
or U12483 (N_12483,N_11458,N_11967);
or U12484 (N_12484,N_11422,N_11815);
nor U12485 (N_12485,N_11481,N_11965);
or U12486 (N_12486,N_11952,N_11804);
nor U12487 (N_12487,N_11812,N_11481);
or U12488 (N_12488,N_11446,N_11436);
nor U12489 (N_12489,N_11631,N_11606);
and U12490 (N_12490,N_11919,N_11412);
nor U12491 (N_12491,N_11529,N_11778);
or U12492 (N_12492,N_11440,N_11792);
or U12493 (N_12493,N_11446,N_11716);
or U12494 (N_12494,N_11884,N_11585);
and U12495 (N_12495,N_11693,N_11810);
nor U12496 (N_12496,N_11836,N_11500);
or U12497 (N_12497,N_11766,N_11850);
nand U12498 (N_12498,N_11508,N_11920);
xnor U12499 (N_12499,N_11820,N_11845);
and U12500 (N_12500,N_11685,N_11499);
or U12501 (N_12501,N_11493,N_11893);
xor U12502 (N_12502,N_11964,N_11840);
nand U12503 (N_12503,N_11996,N_11414);
or U12504 (N_12504,N_11967,N_11674);
xor U12505 (N_12505,N_11556,N_11629);
or U12506 (N_12506,N_11426,N_11759);
xor U12507 (N_12507,N_11627,N_11549);
nor U12508 (N_12508,N_11963,N_11892);
nor U12509 (N_12509,N_11695,N_11495);
or U12510 (N_12510,N_11754,N_11963);
nand U12511 (N_12511,N_11802,N_11732);
nand U12512 (N_12512,N_11936,N_11985);
nor U12513 (N_12513,N_11998,N_11664);
nor U12514 (N_12514,N_11633,N_11926);
and U12515 (N_12515,N_11482,N_11871);
or U12516 (N_12516,N_11907,N_11710);
nor U12517 (N_12517,N_11840,N_11470);
and U12518 (N_12518,N_11675,N_11650);
or U12519 (N_12519,N_11814,N_11493);
and U12520 (N_12520,N_11430,N_11674);
nand U12521 (N_12521,N_11665,N_11505);
and U12522 (N_12522,N_11684,N_11877);
nor U12523 (N_12523,N_11920,N_11650);
and U12524 (N_12524,N_11671,N_11617);
or U12525 (N_12525,N_11942,N_11970);
nand U12526 (N_12526,N_11943,N_11463);
nor U12527 (N_12527,N_11433,N_11987);
or U12528 (N_12528,N_11400,N_11901);
nor U12529 (N_12529,N_11427,N_11876);
and U12530 (N_12530,N_11509,N_11676);
and U12531 (N_12531,N_11806,N_11579);
and U12532 (N_12532,N_11812,N_11885);
or U12533 (N_12533,N_11697,N_11656);
and U12534 (N_12534,N_11884,N_11709);
and U12535 (N_12535,N_11655,N_11661);
xnor U12536 (N_12536,N_11510,N_11454);
xor U12537 (N_12537,N_11479,N_11629);
and U12538 (N_12538,N_11470,N_11866);
or U12539 (N_12539,N_11697,N_11647);
nor U12540 (N_12540,N_11557,N_11749);
nand U12541 (N_12541,N_11569,N_11472);
or U12542 (N_12542,N_11668,N_11810);
and U12543 (N_12543,N_11953,N_11525);
or U12544 (N_12544,N_11529,N_11632);
or U12545 (N_12545,N_11574,N_11565);
nor U12546 (N_12546,N_11746,N_11935);
nand U12547 (N_12547,N_11713,N_11479);
nand U12548 (N_12548,N_11661,N_11928);
and U12549 (N_12549,N_11472,N_11999);
or U12550 (N_12550,N_11458,N_11922);
nand U12551 (N_12551,N_11931,N_11488);
nand U12552 (N_12552,N_11546,N_11777);
or U12553 (N_12553,N_11484,N_11936);
nand U12554 (N_12554,N_11888,N_11923);
nand U12555 (N_12555,N_11836,N_11928);
nor U12556 (N_12556,N_11893,N_11836);
nand U12557 (N_12557,N_11983,N_11664);
or U12558 (N_12558,N_11822,N_11604);
or U12559 (N_12559,N_11678,N_11803);
nand U12560 (N_12560,N_11595,N_11405);
or U12561 (N_12561,N_11530,N_11716);
nor U12562 (N_12562,N_11440,N_11919);
xnor U12563 (N_12563,N_11482,N_11825);
nor U12564 (N_12564,N_11851,N_11843);
nand U12565 (N_12565,N_11455,N_11755);
or U12566 (N_12566,N_11800,N_11541);
or U12567 (N_12567,N_11413,N_11573);
and U12568 (N_12568,N_11548,N_11651);
or U12569 (N_12569,N_11684,N_11704);
xor U12570 (N_12570,N_11746,N_11836);
or U12571 (N_12571,N_11947,N_11635);
or U12572 (N_12572,N_11620,N_11488);
nand U12573 (N_12573,N_11951,N_11980);
nor U12574 (N_12574,N_11726,N_11980);
and U12575 (N_12575,N_11927,N_11777);
or U12576 (N_12576,N_11694,N_11434);
nor U12577 (N_12577,N_11458,N_11454);
or U12578 (N_12578,N_11585,N_11687);
nand U12579 (N_12579,N_11566,N_11499);
nand U12580 (N_12580,N_11445,N_11500);
or U12581 (N_12581,N_11900,N_11541);
or U12582 (N_12582,N_11925,N_11948);
or U12583 (N_12583,N_11448,N_11837);
xor U12584 (N_12584,N_11645,N_11669);
nor U12585 (N_12585,N_11705,N_11823);
nor U12586 (N_12586,N_11783,N_11753);
nor U12587 (N_12587,N_11803,N_11703);
nor U12588 (N_12588,N_11525,N_11909);
xor U12589 (N_12589,N_11493,N_11580);
and U12590 (N_12590,N_11701,N_11609);
nand U12591 (N_12591,N_11887,N_11945);
xnor U12592 (N_12592,N_11600,N_11958);
xnor U12593 (N_12593,N_11885,N_11692);
nor U12594 (N_12594,N_11981,N_11937);
nand U12595 (N_12595,N_11540,N_11862);
or U12596 (N_12596,N_11989,N_11577);
and U12597 (N_12597,N_11410,N_11959);
or U12598 (N_12598,N_11672,N_11676);
nand U12599 (N_12599,N_11600,N_11845);
nand U12600 (N_12600,N_12425,N_12236);
and U12601 (N_12601,N_12054,N_12583);
nor U12602 (N_12602,N_12412,N_12446);
or U12603 (N_12603,N_12521,N_12165);
nor U12604 (N_12604,N_12438,N_12286);
xnor U12605 (N_12605,N_12411,N_12120);
nor U12606 (N_12606,N_12492,N_12262);
nor U12607 (N_12607,N_12226,N_12440);
or U12608 (N_12608,N_12554,N_12366);
nor U12609 (N_12609,N_12448,N_12156);
or U12610 (N_12610,N_12490,N_12562);
nand U12611 (N_12611,N_12198,N_12399);
nand U12612 (N_12612,N_12215,N_12373);
xnor U12613 (N_12613,N_12190,N_12151);
or U12614 (N_12614,N_12204,N_12536);
nor U12615 (N_12615,N_12248,N_12240);
or U12616 (N_12616,N_12047,N_12517);
nand U12617 (N_12617,N_12402,N_12300);
nand U12618 (N_12618,N_12181,N_12103);
and U12619 (N_12619,N_12244,N_12046);
nand U12620 (N_12620,N_12529,N_12026);
nand U12621 (N_12621,N_12436,N_12235);
nand U12622 (N_12622,N_12586,N_12432);
or U12623 (N_12623,N_12407,N_12036);
nor U12624 (N_12624,N_12596,N_12258);
or U12625 (N_12625,N_12506,N_12219);
nor U12626 (N_12626,N_12343,N_12463);
or U12627 (N_12627,N_12063,N_12158);
nand U12628 (N_12628,N_12309,N_12024);
and U12629 (N_12629,N_12322,N_12572);
nand U12630 (N_12630,N_12450,N_12106);
nor U12631 (N_12631,N_12289,N_12569);
and U12632 (N_12632,N_12419,N_12480);
and U12633 (N_12633,N_12067,N_12060);
nand U12634 (N_12634,N_12290,N_12221);
and U12635 (N_12635,N_12305,N_12088);
nor U12636 (N_12636,N_12050,N_12332);
nand U12637 (N_12637,N_12380,N_12141);
and U12638 (N_12638,N_12002,N_12137);
and U12639 (N_12639,N_12145,N_12186);
nor U12640 (N_12640,N_12382,N_12144);
nor U12641 (N_12641,N_12350,N_12577);
nand U12642 (N_12642,N_12581,N_12007);
or U12643 (N_12643,N_12033,N_12409);
nor U12644 (N_12644,N_12514,N_12293);
or U12645 (N_12645,N_12140,N_12534);
and U12646 (N_12646,N_12483,N_12231);
nand U12647 (N_12647,N_12157,N_12593);
nand U12648 (N_12648,N_12225,N_12573);
and U12649 (N_12649,N_12056,N_12051);
and U12650 (N_12650,N_12169,N_12539);
or U12651 (N_12651,N_12361,N_12449);
nand U12652 (N_12652,N_12164,N_12201);
nor U12653 (N_12653,N_12335,N_12223);
and U12654 (N_12654,N_12153,N_12388);
nor U12655 (N_12655,N_12178,N_12229);
nor U12656 (N_12656,N_12136,N_12001);
and U12657 (N_12657,N_12368,N_12179);
nor U12658 (N_12658,N_12207,N_12092);
nor U12659 (N_12659,N_12008,N_12540);
nand U12660 (N_12660,N_12365,N_12414);
or U12661 (N_12661,N_12516,N_12531);
and U12662 (N_12662,N_12148,N_12102);
nor U12663 (N_12663,N_12424,N_12538);
or U12664 (N_12664,N_12316,N_12591);
nor U12665 (N_12665,N_12321,N_12196);
or U12666 (N_12666,N_12356,N_12167);
and U12667 (N_12667,N_12405,N_12049);
and U12668 (N_12668,N_12563,N_12549);
or U12669 (N_12669,N_12061,N_12502);
nor U12670 (N_12670,N_12441,N_12401);
or U12671 (N_12671,N_12325,N_12482);
xnor U12672 (N_12672,N_12452,N_12358);
or U12673 (N_12673,N_12394,N_12101);
or U12674 (N_12674,N_12344,N_12110);
nor U12675 (N_12675,N_12210,N_12097);
nor U12676 (N_12676,N_12149,N_12280);
xor U12677 (N_12677,N_12333,N_12326);
nor U12678 (N_12678,N_12218,N_12121);
xor U12679 (N_12679,N_12413,N_12447);
nor U12680 (N_12680,N_12561,N_12513);
nand U12681 (N_12681,N_12509,N_12014);
and U12682 (N_12682,N_12415,N_12057);
nand U12683 (N_12683,N_12484,N_12062);
nand U12684 (N_12684,N_12515,N_12111);
or U12685 (N_12685,N_12579,N_12260);
or U12686 (N_12686,N_12160,N_12000);
nor U12687 (N_12687,N_12195,N_12220);
nor U12688 (N_12688,N_12085,N_12594);
or U12689 (N_12689,N_12304,N_12255);
nand U12690 (N_12690,N_12267,N_12533);
xor U12691 (N_12691,N_12458,N_12232);
nand U12692 (N_12692,N_12565,N_12445);
nand U12693 (N_12693,N_12173,N_12161);
or U12694 (N_12694,N_12078,N_12574);
or U12695 (N_12695,N_12227,N_12071);
nor U12696 (N_12696,N_12084,N_12471);
xnor U12697 (N_12697,N_12087,N_12090);
and U12698 (N_12698,N_12059,N_12108);
and U12699 (N_12699,N_12212,N_12354);
or U12700 (N_12700,N_12474,N_12155);
and U12701 (N_12701,N_12077,N_12567);
nor U12702 (N_12702,N_12488,N_12177);
nor U12703 (N_12703,N_12132,N_12389);
nor U12704 (N_12704,N_12105,N_12222);
and U12705 (N_12705,N_12434,N_12575);
and U12706 (N_12706,N_12194,N_12557);
nor U12707 (N_12707,N_12597,N_12296);
and U12708 (N_12708,N_12346,N_12537);
or U12709 (N_12709,N_12599,N_12543);
nor U12710 (N_12710,N_12298,N_12393);
xnor U12711 (N_12711,N_12184,N_12152);
or U12712 (N_12712,N_12442,N_12422);
and U12713 (N_12713,N_12009,N_12327);
and U12714 (N_12714,N_12323,N_12498);
and U12715 (N_12715,N_12291,N_12455);
and U12716 (N_12716,N_12328,N_12216);
and U12717 (N_12717,N_12369,N_12270);
or U12718 (N_12718,N_12125,N_12163);
xor U12719 (N_12719,N_12276,N_12138);
or U12720 (N_12720,N_12279,N_12370);
nor U12721 (N_12721,N_12131,N_12428);
nor U12722 (N_12722,N_12550,N_12541);
or U12723 (N_12723,N_12443,N_12199);
and U12724 (N_12724,N_12233,N_12427);
xnor U12725 (N_12725,N_12384,N_12068);
or U12726 (N_12726,N_12004,N_12473);
nand U12727 (N_12727,N_12396,N_12497);
or U12728 (N_12728,N_12080,N_12189);
nor U12729 (N_12729,N_12351,N_12032);
and U12730 (N_12730,N_12025,N_12193);
or U12731 (N_12731,N_12383,N_12525);
and U12732 (N_12732,N_12417,N_12021);
or U12733 (N_12733,N_12238,N_12459);
nand U12734 (N_12734,N_12364,N_12100);
nor U12735 (N_12735,N_12107,N_12268);
nor U12736 (N_12736,N_12188,N_12075);
or U12737 (N_12737,N_12377,N_12392);
xor U12738 (N_12738,N_12421,N_12360);
and U12739 (N_12739,N_12171,N_12493);
nor U12740 (N_12740,N_12578,N_12329);
or U12741 (N_12741,N_12367,N_12083);
xor U12742 (N_12742,N_12315,N_12082);
xor U12743 (N_12743,N_12387,N_12526);
nor U12744 (N_12744,N_12037,N_12451);
xnor U12745 (N_12745,N_12324,N_12313);
or U12746 (N_12746,N_12045,N_12330);
nand U12747 (N_12747,N_12123,N_12041);
or U12748 (N_12748,N_12457,N_12266);
and U12749 (N_12749,N_12499,N_12423);
nor U12750 (N_12750,N_12175,N_12391);
or U12751 (N_12751,N_12522,N_12070);
nand U12752 (N_12752,N_12200,N_12053);
xor U12753 (N_12753,N_12288,N_12371);
or U12754 (N_12754,N_12109,N_12073);
or U12755 (N_12755,N_12485,N_12205);
xor U12756 (N_12756,N_12406,N_12560);
and U12757 (N_12757,N_12456,N_12104);
and U12758 (N_12758,N_12076,N_12507);
nor U12759 (N_12759,N_12020,N_12306);
nor U12760 (N_12760,N_12042,N_12016);
and U12761 (N_12761,N_12019,N_12466);
nand U12762 (N_12762,N_12297,N_12386);
and U12763 (N_12763,N_12079,N_12299);
nand U12764 (N_12764,N_12034,N_12012);
nor U12765 (N_12765,N_12172,N_12095);
nand U12766 (N_12766,N_12501,N_12310);
nor U12767 (N_12767,N_12566,N_12495);
xnor U12768 (N_12768,N_12113,N_12410);
and U12769 (N_12769,N_12242,N_12117);
nand U12770 (N_12770,N_12379,N_12571);
and U12771 (N_12771,N_12269,N_12209);
xor U12772 (N_12772,N_12159,N_12211);
and U12773 (N_12773,N_12408,N_12126);
and U12774 (N_12774,N_12372,N_12069);
and U12775 (N_12775,N_12580,N_12564);
and U12776 (N_12776,N_12547,N_12249);
and U12777 (N_12777,N_12129,N_12086);
or U12778 (N_12778,N_12433,N_12504);
nand U12779 (N_12779,N_12230,N_12055);
nand U12780 (N_12780,N_12314,N_12048);
nand U12781 (N_12781,N_12252,N_12319);
and U12782 (N_12782,N_12342,N_12187);
and U12783 (N_12783,N_12256,N_12264);
nand U12784 (N_12784,N_12524,N_12214);
nand U12785 (N_12785,N_12302,N_12295);
nand U12786 (N_12786,N_12038,N_12303);
nand U12787 (N_12787,N_12588,N_12089);
or U12788 (N_12788,N_12528,N_12185);
and U12789 (N_12789,N_12331,N_12431);
nor U12790 (N_12790,N_12027,N_12228);
nor U12791 (N_12791,N_12239,N_12183);
and U12792 (N_12792,N_12486,N_12548);
and U12793 (N_12793,N_12510,N_12553);
and U12794 (N_12794,N_12162,N_12544);
xor U12795 (N_12795,N_12285,N_12584);
and U12796 (N_12796,N_12017,N_12301);
and U12797 (N_12797,N_12355,N_12166);
and U12798 (N_12798,N_12362,N_12336);
nand U12799 (N_12799,N_12135,N_12124);
or U12800 (N_12800,N_12170,N_12005);
xor U12801 (N_12801,N_12420,N_12479);
nand U12802 (N_12802,N_12527,N_12180);
nor U12803 (N_12803,N_12023,N_12147);
nand U12804 (N_12804,N_12339,N_12146);
nor U12805 (N_12805,N_12418,N_12559);
nor U12806 (N_12806,N_12467,N_12481);
nand U12807 (N_12807,N_12202,N_12203);
nand U12808 (N_12808,N_12378,N_12439);
and U12809 (N_12809,N_12287,N_12546);
nor U12810 (N_12810,N_12568,N_12099);
xnor U12811 (N_12811,N_12592,N_12337);
or U12812 (N_12812,N_12259,N_12503);
and U12813 (N_12813,N_12318,N_12119);
xnor U12814 (N_12814,N_12191,N_12558);
xnor U12815 (N_12815,N_12247,N_12028);
xor U12816 (N_12816,N_12472,N_12555);
nand U12817 (N_12817,N_12031,N_12395);
or U12818 (N_12818,N_12091,N_12345);
and U12819 (N_12819,N_12454,N_12030);
nand U12820 (N_12820,N_12453,N_12081);
nor U12821 (N_12821,N_12074,N_12013);
nor U12822 (N_12822,N_12487,N_12334);
and U12823 (N_12823,N_12064,N_12430);
and U12824 (N_12824,N_12341,N_12251);
or U12825 (N_12825,N_12237,N_12400);
or U12826 (N_12826,N_12530,N_12206);
nand U12827 (N_12827,N_12556,N_12519);
or U12828 (N_12828,N_12347,N_12461);
nor U12829 (N_12829,N_12066,N_12523);
nor U12830 (N_12830,N_12246,N_12176);
nor U12831 (N_12831,N_12311,N_12429);
or U12832 (N_12832,N_12348,N_12403);
or U12833 (N_12833,N_12532,N_12464);
and U12834 (N_12834,N_12508,N_12489);
xor U12835 (N_12835,N_12022,N_12282);
or U12836 (N_12836,N_12312,N_12243);
and U12837 (N_12837,N_12283,N_12093);
and U12838 (N_12838,N_12477,N_12116);
or U12839 (N_12839,N_12254,N_12011);
and U12840 (N_12840,N_12272,N_12468);
nor U12841 (N_12841,N_12128,N_12006);
xor U12842 (N_12842,N_12208,N_12462);
or U12843 (N_12843,N_12234,N_12496);
or U12844 (N_12844,N_12065,N_12435);
nand U12845 (N_12845,N_12320,N_12273);
nor U12846 (N_12846,N_12476,N_12582);
xnor U12847 (N_12847,N_12275,N_12174);
nand U12848 (N_12848,N_12044,N_12197);
nand U12849 (N_12849,N_12150,N_12512);
or U12850 (N_12850,N_12010,N_12122);
or U12851 (N_12851,N_12585,N_12168);
nand U12852 (N_12852,N_12182,N_12317);
and U12853 (N_12853,N_12374,N_12098);
or U12854 (N_12854,N_12587,N_12261);
and U12855 (N_12855,N_12281,N_12294);
nor U12856 (N_12856,N_12217,N_12250);
nor U12857 (N_12857,N_12437,N_12520);
nor U12858 (N_12858,N_12404,N_12511);
or U12859 (N_12859,N_12470,N_12469);
and U12860 (N_12860,N_12551,N_12570);
nand U12861 (N_12861,N_12385,N_12277);
and U12862 (N_12862,N_12213,N_12465);
nand U12863 (N_12863,N_12426,N_12274);
nand U12864 (N_12864,N_12359,N_12154);
or U12865 (N_12865,N_12576,N_12505);
or U12866 (N_12866,N_12003,N_12253);
nand U12867 (N_12867,N_12094,N_12542);
xnor U12868 (N_12868,N_12224,N_12494);
nand U12869 (N_12869,N_12134,N_12444);
nand U12870 (N_12870,N_12015,N_12363);
or U12871 (N_12871,N_12278,N_12352);
and U12872 (N_12872,N_12308,N_12114);
nor U12873 (N_12873,N_12416,N_12595);
and U12874 (N_12874,N_12589,N_12029);
nor U12875 (N_12875,N_12072,N_12143);
or U12876 (N_12876,N_12353,N_12115);
xor U12877 (N_12877,N_12518,N_12307);
nor U12878 (N_12878,N_12381,N_12500);
xnor U12879 (N_12879,N_12130,N_12292);
nand U12880 (N_12880,N_12535,N_12118);
and U12881 (N_12881,N_12375,N_12142);
nand U12882 (N_12882,N_12133,N_12043);
nand U12883 (N_12883,N_12590,N_12397);
nor U12884 (N_12884,N_12357,N_12390);
nor U12885 (N_12885,N_12398,N_12139);
and U12886 (N_12886,N_12475,N_12096);
nor U12887 (N_12887,N_12263,N_12035);
nor U12888 (N_12888,N_12018,N_12245);
nand U12889 (N_12889,N_12340,N_12039);
or U12890 (N_12890,N_12271,N_12478);
nand U12891 (N_12891,N_12545,N_12040);
nand U12892 (N_12892,N_12460,N_12265);
and U12893 (N_12893,N_12112,N_12376);
and U12894 (N_12894,N_12058,N_12052);
nand U12895 (N_12895,N_12241,N_12552);
nand U12896 (N_12896,N_12284,N_12127);
and U12897 (N_12897,N_12192,N_12598);
and U12898 (N_12898,N_12257,N_12338);
or U12899 (N_12899,N_12349,N_12491);
or U12900 (N_12900,N_12230,N_12566);
nor U12901 (N_12901,N_12550,N_12265);
and U12902 (N_12902,N_12067,N_12489);
nor U12903 (N_12903,N_12009,N_12221);
or U12904 (N_12904,N_12475,N_12324);
or U12905 (N_12905,N_12538,N_12201);
nand U12906 (N_12906,N_12540,N_12172);
and U12907 (N_12907,N_12365,N_12159);
or U12908 (N_12908,N_12085,N_12308);
and U12909 (N_12909,N_12008,N_12014);
nand U12910 (N_12910,N_12454,N_12405);
and U12911 (N_12911,N_12473,N_12016);
and U12912 (N_12912,N_12210,N_12266);
or U12913 (N_12913,N_12390,N_12255);
xor U12914 (N_12914,N_12073,N_12186);
or U12915 (N_12915,N_12596,N_12052);
xor U12916 (N_12916,N_12291,N_12063);
or U12917 (N_12917,N_12350,N_12219);
or U12918 (N_12918,N_12224,N_12326);
nand U12919 (N_12919,N_12393,N_12472);
and U12920 (N_12920,N_12013,N_12322);
xor U12921 (N_12921,N_12349,N_12132);
and U12922 (N_12922,N_12123,N_12205);
nor U12923 (N_12923,N_12214,N_12116);
nand U12924 (N_12924,N_12572,N_12201);
nand U12925 (N_12925,N_12480,N_12128);
nor U12926 (N_12926,N_12113,N_12264);
or U12927 (N_12927,N_12153,N_12570);
xnor U12928 (N_12928,N_12565,N_12236);
or U12929 (N_12929,N_12103,N_12427);
nor U12930 (N_12930,N_12319,N_12283);
and U12931 (N_12931,N_12427,N_12449);
or U12932 (N_12932,N_12520,N_12031);
and U12933 (N_12933,N_12336,N_12320);
and U12934 (N_12934,N_12075,N_12392);
or U12935 (N_12935,N_12167,N_12126);
nand U12936 (N_12936,N_12346,N_12220);
and U12937 (N_12937,N_12006,N_12097);
nor U12938 (N_12938,N_12327,N_12035);
nand U12939 (N_12939,N_12557,N_12403);
nor U12940 (N_12940,N_12025,N_12066);
nand U12941 (N_12941,N_12457,N_12372);
or U12942 (N_12942,N_12176,N_12116);
and U12943 (N_12943,N_12590,N_12341);
or U12944 (N_12944,N_12508,N_12022);
xnor U12945 (N_12945,N_12121,N_12518);
and U12946 (N_12946,N_12382,N_12073);
nand U12947 (N_12947,N_12242,N_12429);
and U12948 (N_12948,N_12583,N_12278);
nand U12949 (N_12949,N_12148,N_12025);
or U12950 (N_12950,N_12471,N_12580);
and U12951 (N_12951,N_12526,N_12245);
nand U12952 (N_12952,N_12509,N_12137);
nor U12953 (N_12953,N_12432,N_12463);
nand U12954 (N_12954,N_12052,N_12555);
xor U12955 (N_12955,N_12127,N_12068);
or U12956 (N_12956,N_12275,N_12398);
and U12957 (N_12957,N_12278,N_12574);
or U12958 (N_12958,N_12003,N_12339);
or U12959 (N_12959,N_12477,N_12520);
nand U12960 (N_12960,N_12295,N_12169);
nand U12961 (N_12961,N_12564,N_12248);
xor U12962 (N_12962,N_12293,N_12510);
nand U12963 (N_12963,N_12074,N_12420);
nor U12964 (N_12964,N_12255,N_12122);
and U12965 (N_12965,N_12028,N_12218);
and U12966 (N_12966,N_12106,N_12475);
nand U12967 (N_12967,N_12546,N_12201);
nor U12968 (N_12968,N_12165,N_12390);
or U12969 (N_12969,N_12492,N_12112);
or U12970 (N_12970,N_12131,N_12298);
xnor U12971 (N_12971,N_12582,N_12099);
nand U12972 (N_12972,N_12049,N_12249);
nand U12973 (N_12973,N_12298,N_12508);
nor U12974 (N_12974,N_12105,N_12534);
xnor U12975 (N_12975,N_12136,N_12538);
or U12976 (N_12976,N_12506,N_12172);
and U12977 (N_12977,N_12179,N_12054);
nand U12978 (N_12978,N_12458,N_12253);
nor U12979 (N_12979,N_12031,N_12491);
nor U12980 (N_12980,N_12078,N_12018);
and U12981 (N_12981,N_12137,N_12451);
or U12982 (N_12982,N_12282,N_12089);
nand U12983 (N_12983,N_12512,N_12070);
xnor U12984 (N_12984,N_12594,N_12477);
nor U12985 (N_12985,N_12597,N_12045);
or U12986 (N_12986,N_12126,N_12404);
nand U12987 (N_12987,N_12177,N_12386);
or U12988 (N_12988,N_12133,N_12499);
nor U12989 (N_12989,N_12376,N_12480);
and U12990 (N_12990,N_12578,N_12001);
or U12991 (N_12991,N_12128,N_12382);
or U12992 (N_12992,N_12064,N_12321);
or U12993 (N_12993,N_12374,N_12397);
or U12994 (N_12994,N_12218,N_12556);
or U12995 (N_12995,N_12002,N_12128);
xor U12996 (N_12996,N_12596,N_12049);
xor U12997 (N_12997,N_12575,N_12428);
and U12998 (N_12998,N_12395,N_12200);
or U12999 (N_12999,N_12242,N_12182);
nor U13000 (N_13000,N_12265,N_12105);
xnor U13001 (N_13001,N_12165,N_12191);
and U13002 (N_13002,N_12395,N_12593);
and U13003 (N_13003,N_12502,N_12575);
or U13004 (N_13004,N_12203,N_12267);
nor U13005 (N_13005,N_12082,N_12320);
and U13006 (N_13006,N_12489,N_12569);
or U13007 (N_13007,N_12417,N_12249);
and U13008 (N_13008,N_12060,N_12324);
xor U13009 (N_13009,N_12013,N_12057);
nor U13010 (N_13010,N_12188,N_12492);
or U13011 (N_13011,N_12039,N_12095);
or U13012 (N_13012,N_12292,N_12373);
xor U13013 (N_13013,N_12388,N_12346);
or U13014 (N_13014,N_12011,N_12283);
nor U13015 (N_13015,N_12080,N_12265);
nand U13016 (N_13016,N_12460,N_12443);
nand U13017 (N_13017,N_12010,N_12036);
nand U13018 (N_13018,N_12135,N_12194);
nor U13019 (N_13019,N_12491,N_12586);
nor U13020 (N_13020,N_12489,N_12139);
nand U13021 (N_13021,N_12353,N_12130);
or U13022 (N_13022,N_12185,N_12009);
nand U13023 (N_13023,N_12028,N_12584);
xor U13024 (N_13024,N_12518,N_12493);
nor U13025 (N_13025,N_12188,N_12071);
or U13026 (N_13026,N_12110,N_12125);
or U13027 (N_13027,N_12275,N_12192);
nand U13028 (N_13028,N_12551,N_12515);
and U13029 (N_13029,N_12012,N_12418);
xnor U13030 (N_13030,N_12320,N_12487);
and U13031 (N_13031,N_12183,N_12140);
nor U13032 (N_13032,N_12067,N_12477);
xor U13033 (N_13033,N_12488,N_12533);
or U13034 (N_13034,N_12302,N_12484);
xor U13035 (N_13035,N_12223,N_12302);
and U13036 (N_13036,N_12072,N_12450);
and U13037 (N_13037,N_12331,N_12391);
or U13038 (N_13038,N_12186,N_12546);
nor U13039 (N_13039,N_12407,N_12377);
and U13040 (N_13040,N_12240,N_12133);
or U13041 (N_13041,N_12532,N_12358);
and U13042 (N_13042,N_12361,N_12589);
nor U13043 (N_13043,N_12393,N_12241);
nand U13044 (N_13044,N_12161,N_12522);
xnor U13045 (N_13045,N_12297,N_12259);
and U13046 (N_13046,N_12580,N_12425);
nor U13047 (N_13047,N_12052,N_12390);
and U13048 (N_13048,N_12144,N_12054);
xnor U13049 (N_13049,N_12204,N_12358);
and U13050 (N_13050,N_12391,N_12019);
or U13051 (N_13051,N_12004,N_12388);
xnor U13052 (N_13052,N_12157,N_12068);
nor U13053 (N_13053,N_12348,N_12011);
or U13054 (N_13054,N_12299,N_12067);
or U13055 (N_13055,N_12414,N_12275);
or U13056 (N_13056,N_12316,N_12575);
nand U13057 (N_13057,N_12081,N_12189);
nand U13058 (N_13058,N_12117,N_12582);
or U13059 (N_13059,N_12415,N_12034);
nand U13060 (N_13060,N_12316,N_12550);
xnor U13061 (N_13061,N_12595,N_12227);
and U13062 (N_13062,N_12139,N_12471);
nor U13063 (N_13063,N_12230,N_12105);
nand U13064 (N_13064,N_12040,N_12453);
nand U13065 (N_13065,N_12278,N_12415);
and U13066 (N_13066,N_12564,N_12361);
nand U13067 (N_13067,N_12556,N_12541);
nand U13068 (N_13068,N_12281,N_12082);
and U13069 (N_13069,N_12595,N_12590);
and U13070 (N_13070,N_12464,N_12597);
and U13071 (N_13071,N_12230,N_12093);
and U13072 (N_13072,N_12131,N_12083);
and U13073 (N_13073,N_12377,N_12587);
or U13074 (N_13074,N_12095,N_12012);
nand U13075 (N_13075,N_12157,N_12043);
and U13076 (N_13076,N_12368,N_12180);
and U13077 (N_13077,N_12439,N_12222);
nor U13078 (N_13078,N_12479,N_12545);
or U13079 (N_13079,N_12166,N_12084);
nor U13080 (N_13080,N_12462,N_12130);
or U13081 (N_13081,N_12031,N_12411);
nor U13082 (N_13082,N_12270,N_12060);
nor U13083 (N_13083,N_12357,N_12277);
nand U13084 (N_13084,N_12528,N_12246);
or U13085 (N_13085,N_12355,N_12005);
nor U13086 (N_13086,N_12056,N_12478);
or U13087 (N_13087,N_12203,N_12260);
or U13088 (N_13088,N_12282,N_12244);
or U13089 (N_13089,N_12530,N_12443);
nand U13090 (N_13090,N_12384,N_12546);
and U13091 (N_13091,N_12591,N_12534);
nand U13092 (N_13092,N_12035,N_12227);
or U13093 (N_13093,N_12205,N_12014);
and U13094 (N_13094,N_12438,N_12387);
or U13095 (N_13095,N_12178,N_12180);
nor U13096 (N_13096,N_12140,N_12473);
nor U13097 (N_13097,N_12406,N_12547);
nand U13098 (N_13098,N_12090,N_12199);
and U13099 (N_13099,N_12010,N_12496);
or U13100 (N_13100,N_12230,N_12540);
nand U13101 (N_13101,N_12576,N_12147);
nor U13102 (N_13102,N_12054,N_12189);
and U13103 (N_13103,N_12316,N_12538);
and U13104 (N_13104,N_12146,N_12563);
nor U13105 (N_13105,N_12448,N_12530);
or U13106 (N_13106,N_12502,N_12099);
or U13107 (N_13107,N_12144,N_12106);
nor U13108 (N_13108,N_12433,N_12144);
and U13109 (N_13109,N_12230,N_12469);
xor U13110 (N_13110,N_12571,N_12245);
and U13111 (N_13111,N_12287,N_12101);
or U13112 (N_13112,N_12103,N_12508);
nand U13113 (N_13113,N_12133,N_12286);
nand U13114 (N_13114,N_12316,N_12255);
nand U13115 (N_13115,N_12220,N_12591);
xnor U13116 (N_13116,N_12589,N_12333);
or U13117 (N_13117,N_12387,N_12419);
and U13118 (N_13118,N_12045,N_12561);
and U13119 (N_13119,N_12383,N_12152);
and U13120 (N_13120,N_12364,N_12414);
or U13121 (N_13121,N_12243,N_12106);
and U13122 (N_13122,N_12134,N_12217);
xor U13123 (N_13123,N_12453,N_12210);
and U13124 (N_13124,N_12372,N_12329);
nand U13125 (N_13125,N_12457,N_12463);
nand U13126 (N_13126,N_12226,N_12373);
and U13127 (N_13127,N_12328,N_12378);
or U13128 (N_13128,N_12556,N_12436);
nor U13129 (N_13129,N_12275,N_12130);
and U13130 (N_13130,N_12294,N_12058);
nor U13131 (N_13131,N_12076,N_12021);
or U13132 (N_13132,N_12482,N_12078);
nor U13133 (N_13133,N_12142,N_12373);
nand U13134 (N_13134,N_12269,N_12433);
nor U13135 (N_13135,N_12500,N_12471);
nand U13136 (N_13136,N_12315,N_12480);
and U13137 (N_13137,N_12232,N_12179);
or U13138 (N_13138,N_12112,N_12027);
nor U13139 (N_13139,N_12150,N_12035);
nand U13140 (N_13140,N_12474,N_12396);
nor U13141 (N_13141,N_12351,N_12080);
nand U13142 (N_13142,N_12060,N_12316);
nor U13143 (N_13143,N_12033,N_12070);
xor U13144 (N_13144,N_12461,N_12469);
or U13145 (N_13145,N_12474,N_12271);
or U13146 (N_13146,N_12091,N_12164);
nand U13147 (N_13147,N_12262,N_12218);
xnor U13148 (N_13148,N_12189,N_12339);
or U13149 (N_13149,N_12080,N_12131);
and U13150 (N_13150,N_12433,N_12082);
or U13151 (N_13151,N_12327,N_12164);
or U13152 (N_13152,N_12225,N_12285);
nand U13153 (N_13153,N_12069,N_12361);
or U13154 (N_13154,N_12222,N_12216);
nor U13155 (N_13155,N_12278,N_12076);
xor U13156 (N_13156,N_12068,N_12023);
nand U13157 (N_13157,N_12335,N_12473);
or U13158 (N_13158,N_12549,N_12462);
and U13159 (N_13159,N_12048,N_12448);
nor U13160 (N_13160,N_12261,N_12008);
xnor U13161 (N_13161,N_12260,N_12003);
nand U13162 (N_13162,N_12257,N_12218);
or U13163 (N_13163,N_12315,N_12347);
nor U13164 (N_13164,N_12332,N_12219);
xor U13165 (N_13165,N_12594,N_12206);
xnor U13166 (N_13166,N_12258,N_12337);
xor U13167 (N_13167,N_12347,N_12393);
nor U13168 (N_13168,N_12419,N_12432);
or U13169 (N_13169,N_12504,N_12493);
and U13170 (N_13170,N_12254,N_12539);
nand U13171 (N_13171,N_12385,N_12448);
nor U13172 (N_13172,N_12378,N_12182);
or U13173 (N_13173,N_12002,N_12281);
nand U13174 (N_13174,N_12457,N_12306);
nand U13175 (N_13175,N_12335,N_12013);
and U13176 (N_13176,N_12537,N_12076);
nand U13177 (N_13177,N_12208,N_12133);
xor U13178 (N_13178,N_12536,N_12318);
or U13179 (N_13179,N_12176,N_12026);
xor U13180 (N_13180,N_12408,N_12519);
xnor U13181 (N_13181,N_12510,N_12176);
and U13182 (N_13182,N_12026,N_12192);
and U13183 (N_13183,N_12015,N_12019);
nor U13184 (N_13184,N_12528,N_12191);
and U13185 (N_13185,N_12431,N_12374);
nor U13186 (N_13186,N_12121,N_12193);
xor U13187 (N_13187,N_12366,N_12252);
nor U13188 (N_13188,N_12207,N_12521);
or U13189 (N_13189,N_12350,N_12340);
nor U13190 (N_13190,N_12552,N_12157);
and U13191 (N_13191,N_12149,N_12228);
nand U13192 (N_13192,N_12485,N_12230);
or U13193 (N_13193,N_12287,N_12014);
nand U13194 (N_13194,N_12080,N_12241);
xnor U13195 (N_13195,N_12241,N_12221);
and U13196 (N_13196,N_12497,N_12255);
or U13197 (N_13197,N_12210,N_12376);
and U13198 (N_13198,N_12085,N_12020);
nor U13199 (N_13199,N_12479,N_12492);
nand U13200 (N_13200,N_12857,N_13155);
nor U13201 (N_13201,N_12909,N_12939);
or U13202 (N_13202,N_13165,N_13088);
and U13203 (N_13203,N_13098,N_12675);
or U13204 (N_13204,N_13034,N_12902);
and U13205 (N_13205,N_12933,N_12922);
or U13206 (N_13206,N_12987,N_12839);
nand U13207 (N_13207,N_12957,N_12782);
nor U13208 (N_13208,N_12806,N_13141);
nor U13209 (N_13209,N_12934,N_12709);
nor U13210 (N_13210,N_12965,N_12668);
nor U13211 (N_13211,N_12702,N_12863);
and U13212 (N_13212,N_13095,N_12884);
or U13213 (N_13213,N_12606,N_13049);
nand U13214 (N_13214,N_12836,N_12880);
xnor U13215 (N_13215,N_12680,N_12859);
or U13216 (N_13216,N_13057,N_13009);
nor U13217 (N_13217,N_12755,N_12916);
and U13218 (N_13218,N_12866,N_12911);
and U13219 (N_13219,N_13132,N_12918);
or U13220 (N_13220,N_12984,N_13094);
nor U13221 (N_13221,N_13025,N_12868);
or U13222 (N_13222,N_13153,N_13100);
nor U13223 (N_13223,N_12627,N_12721);
or U13224 (N_13224,N_13037,N_12813);
or U13225 (N_13225,N_12960,N_13156);
nand U13226 (N_13226,N_12601,N_12656);
nand U13227 (N_13227,N_12614,N_13067);
nor U13228 (N_13228,N_12788,N_12847);
xor U13229 (N_13229,N_12958,N_12753);
nand U13230 (N_13230,N_12695,N_12797);
nand U13231 (N_13231,N_12832,N_12658);
and U13232 (N_13232,N_13041,N_12890);
nor U13233 (N_13233,N_12993,N_13096);
xor U13234 (N_13234,N_13086,N_12981);
nand U13235 (N_13235,N_12701,N_12693);
or U13236 (N_13236,N_13070,N_12745);
nor U13237 (N_13237,N_12897,N_12842);
nand U13238 (N_13238,N_13176,N_13074);
or U13239 (N_13239,N_12698,N_13033);
and U13240 (N_13240,N_13027,N_13131);
or U13241 (N_13241,N_13022,N_12643);
nor U13242 (N_13242,N_12878,N_12792);
or U13243 (N_13243,N_13197,N_13196);
and U13244 (N_13244,N_12864,N_13122);
nand U13245 (N_13245,N_13105,N_12600);
nand U13246 (N_13246,N_13136,N_13108);
nor U13247 (N_13247,N_13147,N_13007);
and U13248 (N_13248,N_13056,N_12616);
and U13249 (N_13249,N_12858,N_12715);
or U13250 (N_13250,N_13188,N_12853);
nand U13251 (N_13251,N_13183,N_12964);
or U13252 (N_13252,N_13148,N_13015);
or U13253 (N_13253,N_12850,N_12990);
nand U13254 (N_13254,N_13043,N_12659);
and U13255 (N_13255,N_12881,N_13128);
nand U13256 (N_13256,N_12920,N_12846);
nor U13257 (N_13257,N_12952,N_13054);
nor U13258 (N_13258,N_12812,N_12899);
and U13259 (N_13259,N_13115,N_13039);
or U13260 (N_13260,N_12891,N_13012);
nor U13261 (N_13261,N_12720,N_12672);
nor U13262 (N_13262,N_13016,N_13199);
or U13263 (N_13263,N_12856,N_12996);
and U13264 (N_13264,N_13004,N_12908);
nor U13265 (N_13265,N_13006,N_12862);
xor U13266 (N_13266,N_12674,N_12626);
nor U13267 (N_13267,N_12946,N_12975);
xor U13268 (N_13268,N_13024,N_12982);
nand U13269 (N_13269,N_13064,N_12795);
nand U13270 (N_13270,N_12738,N_13083);
nand U13271 (N_13271,N_13110,N_12855);
nor U13272 (N_13272,N_12811,N_12630);
and U13273 (N_13273,N_12929,N_12687);
nand U13274 (N_13274,N_12694,N_12882);
or U13275 (N_13275,N_12926,N_12779);
nor U13276 (N_13276,N_12725,N_12763);
and U13277 (N_13277,N_13106,N_13052);
nand U13278 (N_13278,N_12727,N_13062);
or U13279 (N_13279,N_12673,N_13129);
xnor U13280 (N_13280,N_13080,N_13111);
or U13281 (N_13281,N_12823,N_13142);
xor U13282 (N_13282,N_12657,N_13189);
or U13283 (N_13283,N_12991,N_12815);
nand U13284 (N_13284,N_12615,N_13055);
and U13285 (N_13285,N_12968,N_12724);
nor U13286 (N_13286,N_13198,N_12731);
and U13287 (N_13287,N_12744,N_12677);
xor U13288 (N_13288,N_12739,N_13123);
nand U13289 (N_13289,N_12752,N_12754);
and U13290 (N_13290,N_12661,N_12875);
nor U13291 (N_13291,N_13097,N_12961);
and U13292 (N_13292,N_12901,N_12722);
nor U13293 (N_13293,N_12790,N_12632);
and U13294 (N_13294,N_12649,N_12666);
nor U13295 (N_13295,N_12989,N_12607);
or U13296 (N_13296,N_12861,N_13134);
nor U13297 (N_13297,N_13050,N_12954);
nand U13298 (N_13298,N_13171,N_12817);
nor U13299 (N_13299,N_12772,N_12634);
and U13300 (N_13300,N_13150,N_13186);
and U13301 (N_13301,N_12704,N_13051);
and U13302 (N_13302,N_13184,N_12910);
nor U13303 (N_13303,N_12807,N_13118);
nand U13304 (N_13304,N_12953,N_12733);
nand U13305 (N_13305,N_12783,N_13047);
xnor U13306 (N_13306,N_12775,N_12757);
nand U13307 (N_13307,N_13014,N_12718);
xnor U13308 (N_13308,N_12711,N_13018);
and U13309 (N_13309,N_13072,N_13135);
or U13310 (N_13310,N_12609,N_12635);
nor U13311 (N_13311,N_13140,N_13120);
or U13312 (N_13312,N_12851,N_12928);
and U13313 (N_13313,N_13117,N_12760);
xor U13314 (N_13314,N_12737,N_12869);
nand U13315 (N_13315,N_12637,N_12735);
xor U13316 (N_13316,N_12845,N_13044);
and U13317 (N_13317,N_12781,N_12726);
xor U13318 (N_13318,N_12919,N_12655);
or U13319 (N_13319,N_13030,N_12917);
or U13320 (N_13320,N_12818,N_12913);
and U13321 (N_13321,N_13107,N_12692);
or U13322 (N_13322,N_12784,N_13119);
nand U13323 (N_13323,N_12728,N_12825);
nand U13324 (N_13324,N_12977,N_12619);
and U13325 (N_13325,N_12611,N_13082);
and U13326 (N_13326,N_12923,N_12604);
nor U13327 (N_13327,N_12710,N_12895);
and U13328 (N_13328,N_13146,N_12925);
nor U13329 (N_13329,N_12906,N_12874);
and U13330 (N_13330,N_12667,N_12730);
or U13331 (N_13331,N_13040,N_12723);
nand U13332 (N_13332,N_12931,N_12793);
nor U13333 (N_13333,N_13036,N_13164);
or U13334 (N_13334,N_12803,N_13157);
or U13335 (N_13335,N_12713,N_13159);
nor U13336 (N_13336,N_12888,N_13104);
nand U13337 (N_13337,N_13075,N_12940);
nand U13338 (N_13338,N_12603,N_13170);
nand U13339 (N_13339,N_13138,N_12900);
nor U13340 (N_13340,N_13116,N_12912);
and U13341 (N_13341,N_12962,N_12700);
nor U13342 (N_13342,N_13112,N_12663);
and U13343 (N_13343,N_12871,N_12801);
nand U13344 (N_13344,N_13090,N_13089);
and U13345 (N_13345,N_13008,N_12708);
nand U13346 (N_13346,N_13169,N_12646);
nor U13347 (N_13347,N_12914,N_12771);
nor U13348 (N_13348,N_12865,N_13173);
and U13349 (N_13349,N_12835,N_12955);
and U13350 (N_13350,N_13068,N_12786);
xnor U13351 (N_13351,N_12773,N_12664);
or U13352 (N_13352,N_12935,N_12650);
or U13353 (N_13353,N_12742,N_13028);
or U13354 (N_13354,N_12746,N_13139);
nand U13355 (N_13355,N_13045,N_12791);
and U13356 (N_13356,N_12610,N_12870);
nand U13357 (N_13357,N_13092,N_12831);
xnor U13358 (N_13358,N_13023,N_12660);
nand U13359 (N_13359,N_12800,N_12948);
or U13360 (N_13360,N_13127,N_13187);
and U13361 (N_13361,N_13069,N_12652);
nand U13362 (N_13362,N_12904,N_12764);
nand U13363 (N_13363,N_12893,N_12822);
or U13364 (N_13364,N_12683,N_12613);
or U13365 (N_13365,N_13162,N_12877);
and U13366 (N_13366,N_12608,N_12809);
or U13367 (N_13367,N_12682,N_12636);
nand U13368 (N_13368,N_12684,N_12770);
or U13369 (N_13369,N_13087,N_13003);
and U13370 (N_13370,N_12768,N_12988);
nor U13371 (N_13371,N_12885,N_12645);
nor U13372 (N_13372,N_13046,N_13042);
or U13373 (N_13373,N_12816,N_12819);
nor U13374 (N_13374,N_13060,N_12998);
and U13375 (N_13375,N_12685,N_12921);
nor U13376 (N_13376,N_12976,N_13126);
nor U13377 (N_13377,N_12936,N_13099);
and U13378 (N_13378,N_12872,N_13031);
and U13379 (N_13379,N_12905,N_12686);
nand U13380 (N_13380,N_13026,N_13061);
nand U13381 (N_13381,N_12621,N_13181);
nor U13382 (N_13382,N_12617,N_12691);
or U13383 (N_13383,N_12756,N_13058);
nor U13384 (N_13384,N_13194,N_12867);
nor U13385 (N_13385,N_12808,N_12985);
or U13386 (N_13386,N_12924,N_13172);
or U13387 (N_13387,N_12972,N_13137);
nor U13388 (N_13388,N_12612,N_13010);
xnor U13389 (N_13389,N_12761,N_13193);
or U13390 (N_13390,N_12741,N_12986);
and U13391 (N_13391,N_13048,N_12769);
nand U13392 (N_13392,N_12780,N_12837);
nor U13393 (N_13393,N_13190,N_12938);
nor U13394 (N_13394,N_12676,N_12707);
nor U13395 (N_13395,N_12994,N_12767);
or U13396 (N_13396,N_12907,N_12876);
xnor U13397 (N_13397,N_12844,N_12852);
and U13398 (N_13398,N_12841,N_13178);
nor U13399 (N_13399,N_12622,N_12894);
nor U13400 (N_13400,N_12631,N_12980);
nor U13401 (N_13401,N_13168,N_12947);
nand U13402 (N_13402,N_12679,N_12641);
and U13403 (N_13403,N_13195,N_12849);
or U13404 (N_13404,N_12618,N_13065);
and U13405 (N_13405,N_12978,N_12665);
nor U13406 (N_13406,N_12814,N_13079);
xor U13407 (N_13407,N_12689,N_12824);
or U13408 (N_13408,N_13017,N_12966);
nand U13409 (N_13409,N_13143,N_13076);
nand U13410 (N_13410,N_12678,N_12898);
nand U13411 (N_13411,N_12838,N_12602);
nor U13412 (N_13412,N_13191,N_12973);
and U13413 (N_13413,N_12777,N_13019);
nor U13414 (N_13414,N_12706,N_13059);
xnor U13415 (N_13415,N_12827,N_12640);
or U13416 (N_13416,N_13163,N_13103);
or U13417 (N_13417,N_12605,N_13001);
or U13418 (N_13418,N_12633,N_12860);
nor U13419 (N_13419,N_12889,N_12951);
or U13420 (N_13420,N_12759,N_13020);
nand U13421 (N_13421,N_12941,N_13152);
and U13422 (N_13422,N_12840,N_13066);
nand U13423 (N_13423,N_13011,N_12690);
nor U13424 (N_13424,N_12944,N_12949);
xnor U13425 (N_13425,N_13158,N_12794);
or U13426 (N_13426,N_13101,N_13021);
and U13427 (N_13427,N_12669,N_12751);
or U13428 (N_13428,N_12624,N_12758);
nor U13429 (N_13429,N_12719,N_12826);
nor U13430 (N_13430,N_13093,N_12647);
and U13431 (N_13431,N_13077,N_12648);
or U13432 (N_13432,N_12969,N_12785);
nor U13433 (N_13433,N_12915,N_12696);
nand U13434 (N_13434,N_13078,N_13177);
and U13435 (N_13435,N_12716,N_12732);
nand U13436 (N_13436,N_13121,N_13109);
xor U13437 (N_13437,N_12638,N_12821);
nand U13438 (N_13438,N_12620,N_13182);
nand U13439 (N_13439,N_12749,N_12774);
nand U13440 (N_13440,N_12688,N_13174);
and U13441 (N_13441,N_12628,N_12886);
and U13442 (N_13442,N_13166,N_12950);
or U13443 (N_13443,N_13144,N_13149);
and U13444 (N_13444,N_12712,N_12903);
nor U13445 (N_13445,N_12830,N_12896);
nand U13446 (N_13446,N_13124,N_12623);
or U13447 (N_13447,N_12887,N_12820);
nand U13448 (N_13448,N_12681,N_12802);
or U13449 (N_13449,N_13161,N_12729);
nand U13450 (N_13450,N_12766,N_13167);
nor U13451 (N_13451,N_12883,N_12625);
nor U13452 (N_13452,N_12748,N_12997);
nand U13453 (N_13453,N_13154,N_13102);
or U13454 (N_13454,N_12644,N_12979);
or U13455 (N_13455,N_12833,N_12629);
xor U13456 (N_13456,N_12743,N_13084);
xor U13457 (N_13457,N_13160,N_12932);
or U13458 (N_13458,N_12703,N_12747);
and U13459 (N_13459,N_13053,N_12854);
and U13460 (N_13460,N_12717,N_13038);
nor U13461 (N_13461,N_13179,N_12937);
or U13462 (N_13462,N_12699,N_12983);
xor U13463 (N_13463,N_12943,N_12654);
or U13464 (N_13464,N_13085,N_12671);
or U13465 (N_13465,N_12829,N_12798);
nand U13466 (N_13466,N_13133,N_13185);
nor U13467 (N_13467,N_13029,N_13071);
nand U13468 (N_13468,N_13091,N_12974);
or U13469 (N_13469,N_12828,N_13063);
xnor U13470 (N_13470,N_12651,N_12740);
nor U13471 (N_13471,N_12971,N_13130);
or U13472 (N_13472,N_12810,N_13192);
or U13473 (N_13473,N_12642,N_12705);
nor U13474 (N_13474,N_12967,N_12787);
nor U13475 (N_13475,N_12959,N_12999);
and U13476 (N_13476,N_12736,N_13000);
or U13477 (N_13477,N_13073,N_12778);
nand U13478 (N_13478,N_12804,N_12697);
xor U13479 (N_13479,N_12992,N_12750);
nor U13480 (N_13480,N_13002,N_12834);
nor U13481 (N_13481,N_12879,N_12945);
xnor U13482 (N_13482,N_12714,N_12843);
nand U13483 (N_13483,N_13180,N_13114);
or U13484 (N_13484,N_13175,N_12930);
and U13485 (N_13485,N_12796,N_12639);
xnor U13486 (N_13486,N_13145,N_12892);
nor U13487 (N_13487,N_12765,N_12799);
and U13488 (N_13488,N_12848,N_13081);
or U13489 (N_13489,N_12653,N_12963);
nand U13490 (N_13490,N_13035,N_12762);
nand U13491 (N_13491,N_12805,N_12776);
nand U13492 (N_13492,N_12995,N_12942);
nand U13493 (N_13493,N_12873,N_12662);
nand U13494 (N_13494,N_12956,N_13032);
or U13495 (N_13495,N_12670,N_13005);
or U13496 (N_13496,N_13151,N_12789);
and U13497 (N_13497,N_12734,N_12927);
and U13498 (N_13498,N_13013,N_12970);
nand U13499 (N_13499,N_13113,N_13125);
or U13500 (N_13500,N_12914,N_12876);
xnor U13501 (N_13501,N_12661,N_12991);
xnor U13502 (N_13502,N_12969,N_12662);
nand U13503 (N_13503,N_13036,N_13018);
nand U13504 (N_13504,N_13127,N_12674);
or U13505 (N_13505,N_12812,N_12926);
and U13506 (N_13506,N_12907,N_13181);
and U13507 (N_13507,N_12627,N_13121);
nor U13508 (N_13508,N_12683,N_12952);
or U13509 (N_13509,N_12752,N_12629);
or U13510 (N_13510,N_12943,N_13074);
and U13511 (N_13511,N_12950,N_12683);
nor U13512 (N_13512,N_12766,N_13133);
nor U13513 (N_13513,N_12677,N_13047);
nor U13514 (N_13514,N_12696,N_12650);
and U13515 (N_13515,N_13141,N_12659);
and U13516 (N_13516,N_12736,N_12767);
nand U13517 (N_13517,N_12820,N_12663);
or U13518 (N_13518,N_13068,N_12762);
or U13519 (N_13519,N_13067,N_13084);
nor U13520 (N_13520,N_12824,N_13045);
xor U13521 (N_13521,N_12800,N_13092);
or U13522 (N_13522,N_12962,N_13014);
nand U13523 (N_13523,N_13183,N_12717);
or U13524 (N_13524,N_13138,N_12675);
or U13525 (N_13525,N_12854,N_12830);
and U13526 (N_13526,N_12838,N_13174);
nor U13527 (N_13527,N_12924,N_13136);
xor U13528 (N_13528,N_13048,N_12647);
or U13529 (N_13529,N_12848,N_12709);
nor U13530 (N_13530,N_13178,N_12782);
and U13531 (N_13531,N_12699,N_12929);
nand U13532 (N_13532,N_13013,N_12815);
xor U13533 (N_13533,N_13160,N_12603);
nand U13534 (N_13534,N_12856,N_13041);
xor U13535 (N_13535,N_13024,N_12831);
or U13536 (N_13536,N_12956,N_13190);
nor U13537 (N_13537,N_12632,N_12798);
xor U13538 (N_13538,N_12972,N_12763);
nor U13539 (N_13539,N_13187,N_12771);
nand U13540 (N_13540,N_12997,N_13105);
nand U13541 (N_13541,N_12783,N_13006);
or U13542 (N_13542,N_12890,N_12809);
nor U13543 (N_13543,N_12928,N_12815);
nor U13544 (N_13544,N_12813,N_12941);
nor U13545 (N_13545,N_13076,N_13013);
xor U13546 (N_13546,N_13003,N_12932);
or U13547 (N_13547,N_12614,N_13010);
nand U13548 (N_13548,N_12925,N_12762);
nand U13549 (N_13549,N_12656,N_12873);
xnor U13550 (N_13550,N_12834,N_13177);
and U13551 (N_13551,N_12870,N_12829);
nor U13552 (N_13552,N_12813,N_12945);
nor U13553 (N_13553,N_12748,N_12781);
nor U13554 (N_13554,N_12923,N_12780);
nor U13555 (N_13555,N_13046,N_12604);
xnor U13556 (N_13556,N_13060,N_12890);
and U13557 (N_13557,N_13066,N_12929);
nand U13558 (N_13558,N_13062,N_12702);
nand U13559 (N_13559,N_12776,N_12912);
xnor U13560 (N_13560,N_13071,N_13095);
or U13561 (N_13561,N_13053,N_13032);
nor U13562 (N_13562,N_13038,N_12969);
or U13563 (N_13563,N_12757,N_12746);
and U13564 (N_13564,N_13191,N_12809);
nor U13565 (N_13565,N_13146,N_13058);
nor U13566 (N_13566,N_12895,N_12628);
nand U13567 (N_13567,N_12752,N_12774);
nand U13568 (N_13568,N_13075,N_12780);
and U13569 (N_13569,N_12991,N_12755);
nand U13570 (N_13570,N_13032,N_12806);
nand U13571 (N_13571,N_13089,N_12814);
nand U13572 (N_13572,N_13028,N_12839);
nand U13573 (N_13573,N_12977,N_12801);
nor U13574 (N_13574,N_12823,N_13057);
or U13575 (N_13575,N_12730,N_12688);
xnor U13576 (N_13576,N_13135,N_12762);
nor U13577 (N_13577,N_12601,N_12961);
nor U13578 (N_13578,N_12988,N_12850);
and U13579 (N_13579,N_12805,N_12778);
nor U13580 (N_13580,N_13174,N_12912);
and U13581 (N_13581,N_12970,N_12840);
and U13582 (N_13582,N_12707,N_13083);
nor U13583 (N_13583,N_12622,N_12914);
and U13584 (N_13584,N_12705,N_12726);
nand U13585 (N_13585,N_12653,N_12952);
nor U13586 (N_13586,N_12687,N_12767);
nand U13587 (N_13587,N_12610,N_12739);
nand U13588 (N_13588,N_12947,N_13012);
or U13589 (N_13589,N_13148,N_12787);
or U13590 (N_13590,N_12776,N_12777);
or U13591 (N_13591,N_13065,N_12962);
nand U13592 (N_13592,N_12725,N_12743);
or U13593 (N_13593,N_12750,N_12959);
or U13594 (N_13594,N_12622,N_12787);
and U13595 (N_13595,N_12983,N_13062);
nor U13596 (N_13596,N_12696,N_12785);
or U13597 (N_13597,N_12770,N_12812);
nor U13598 (N_13598,N_12614,N_12675);
and U13599 (N_13599,N_12702,N_12637);
nand U13600 (N_13600,N_12925,N_13095);
nand U13601 (N_13601,N_13072,N_12905);
and U13602 (N_13602,N_12947,N_13195);
xnor U13603 (N_13603,N_12902,N_13174);
nor U13604 (N_13604,N_12856,N_12748);
nor U13605 (N_13605,N_12901,N_12871);
and U13606 (N_13606,N_12606,N_13136);
or U13607 (N_13607,N_13119,N_13039);
nor U13608 (N_13608,N_12921,N_12936);
xor U13609 (N_13609,N_12962,N_12846);
or U13610 (N_13610,N_12898,N_12761);
nor U13611 (N_13611,N_12967,N_13188);
and U13612 (N_13612,N_12773,N_12845);
nand U13613 (N_13613,N_12767,N_13019);
nand U13614 (N_13614,N_12839,N_12795);
and U13615 (N_13615,N_12645,N_12787);
nand U13616 (N_13616,N_12673,N_12635);
and U13617 (N_13617,N_12683,N_13015);
nand U13618 (N_13618,N_13045,N_12924);
xor U13619 (N_13619,N_12905,N_13114);
and U13620 (N_13620,N_12644,N_12987);
nand U13621 (N_13621,N_12916,N_12983);
nand U13622 (N_13622,N_13051,N_13090);
xnor U13623 (N_13623,N_12808,N_13071);
nand U13624 (N_13624,N_12697,N_13038);
and U13625 (N_13625,N_12841,N_12930);
xnor U13626 (N_13626,N_13073,N_13006);
nand U13627 (N_13627,N_13110,N_12697);
nor U13628 (N_13628,N_12775,N_12833);
nand U13629 (N_13629,N_13154,N_12776);
nor U13630 (N_13630,N_13056,N_12950);
nor U13631 (N_13631,N_13085,N_12989);
or U13632 (N_13632,N_12792,N_13001);
nand U13633 (N_13633,N_12675,N_12971);
or U13634 (N_13634,N_12708,N_12739);
xnor U13635 (N_13635,N_13161,N_12762);
nand U13636 (N_13636,N_12747,N_12736);
nor U13637 (N_13637,N_13071,N_12816);
nor U13638 (N_13638,N_12842,N_13194);
nand U13639 (N_13639,N_12931,N_12842);
or U13640 (N_13640,N_12758,N_12889);
nor U13641 (N_13641,N_12625,N_12952);
nor U13642 (N_13642,N_13196,N_12946);
or U13643 (N_13643,N_13183,N_12816);
and U13644 (N_13644,N_13138,N_13192);
nand U13645 (N_13645,N_12642,N_12748);
or U13646 (N_13646,N_12821,N_12710);
or U13647 (N_13647,N_13032,N_12786);
or U13648 (N_13648,N_12735,N_12699);
and U13649 (N_13649,N_12701,N_13062);
or U13650 (N_13650,N_12668,N_12767);
and U13651 (N_13651,N_12771,N_12687);
nand U13652 (N_13652,N_12728,N_12965);
nor U13653 (N_13653,N_13070,N_13085);
nand U13654 (N_13654,N_13042,N_13023);
and U13655 (N_13655,N_12989,N_13167);
nand U13656 (N_13656,N_12659,N_12696);
xnor U13657 (N_13657,N_12962,N_13060);
or U13658 (N_13658,N_12871,N_12765);
nor U13659 (N_13659,N_12626,N_12832);
nand U13660 (N_13660,N_12629,N_12724);
nor U13661 (N_13661,N_12997,N_12733);
xor U13662 (N_13662,N_13029,N_12774);
nor U13663 (N_13663,N_13053,N_13193);
nand U13664 (N_13664,N_12931,N_13086);
xor U13665 (N_13665,N_12875,N_12876);
xor U13666 (N_13666,N_12672,N_12820);
nand U13667 (N_13667,N_13103,N_12783);
nand U13668 (N_13668,N_12972,N_13070);
xnor U13669 (N_13669,N_13133,N_13043);
nand U13670 (N_13670,N_12617,N_13089);
nor U13671 (N_13671,N_12603,N_13195);
nor U13672 (N_13672,N_12642,N_12696);
xnor U13673 (N_13673,N_12860,N_12684);
xnor U13674 (N_13674,N_13179,N_12798);
nor U13675 (N_13675,N_12653,N_13171);
xor U13676 (N_13676,N_13092,N_13143);
nor U13677 (N_13677,N_12739,N_12690);
nor U13678 (N_13678,N_13098,N_12786);
nor U13679 (N_13679,N_12639,N_13035);
nand U13680 (N_13680,N_12930,N_12958);
and U13681 (N_13681,N_12937,N_12987);
or U13682 (N_13682,N_12942,N_13122);
and U13683 (N_13683,N_13188,N_12663);
xor U13684 (N_13684,N_12741,N_13163);
nand U13685 (N_13685,N_13079,N_12734);
nand U13686 (N_13686,N_12661,N_12809);
or U13687 (N_13687,N_12728,N_12824);
or U13688 (N_13688,N_12633,N_13147);
nand U13689 (N_13689,N_13102,N_12921);
or U13690 (N_13690,N_13039,N_12895);
nand U13691 (N_13691,N_12740,N_12619);
nor U13692 (N_13692,N_12824,N_12823);
nand U13693 (N_13693,N_12876,N_13176);
nor U13694 (N_13694,N_13112,N_12921);
or U13695 (N_13695,N_13154,N_13119);
xor U13696 (N_13696,N_13179,N_12910);
and U13697 (N_13697,N_13038,N_12701);
and U13698 (N_13698,N_12820,N_12970);
nand U13699 (N_13699,N_12634,N_13080);
xor U13700 (N_13700,N_12891,N_12769);
nand U13701 (N_13701,N_13002,N_12649);
nand U13702 (N_13702,N_12720,N_12932);
nand U13703 (N_13703,N_12640,N_12881);
or U13704 (N_13704,N_13010,N_13004);
xor U13705 (N_13705,N_12912,N_12820);
nand U13706 (N_13706,N_12714,N_12985);
xor U13707 (N_13707,N_12915,N_12839);
xor U13708 (N_13708,N_13159,N_12733);
nor U13709 (N_13709,N_12823,N_12909);
nor U13710 (N_13710,N_13021,N_13178);
and U13711 (N_13711,N_12870,N_13035);
nor U13712 (N_13712,N_13114,N_12991);
or U13713 (N_13713,N_13045,N_13160);
and U13714 (N_13714,N_12937,N_12698);
nand U13715 (N_13715,N_12967,N_12620);
and U13716 (N_13716,N_12828,N_12875);
nor U13717 (N_13717,N_12608,N_12695);
nand U13718 (N_13718,N_12890,N_13108);
and U13719 (N_13719,N_12675,N_12722);
nor U13720 (N_13720,N_12628,N_12964);
nor U13721 (N_13721,N_12928,N_12806);
or U13722 (N_13722,N_12629,N_12856);
nand U13723 (N_13723,N_13026,N_13126);
nand U13724 (N_13724,N_12668,N_12940);
and U13725 (N_13725,N_12952,N_13003);
or U13726 (N_13726,N_13154,N_12841);
or U13727 (N_13727,N_12636,N_13105);
xnor U13728 (N_13728,N_12940,N_12697);
xor U13729 (N_13729,N_12617,N_12799);
and U13730 (N_13730,N_12638,N_12964);
nor U13731 (N_13731,N_12711,N_12938);
xor U13732 (N_13732,N_12934,N_12760);
or U13733 (N_13733,N_12779,N_12624);
and U13734 (N_13734,N_12611,N_12759);
nand U13735 (N_13735,N_12801,N_12990);
or U13736 (N_13736,N_12968,N_12676);
nor U13737 (N_13737,N_12883,N_12647);
and U13738 (N_13738,N_12961,N_12922);
nor U13739 (N_13739,N_12709,N_12660);
or U13740 (N_13740,N_13013,N_12877);
xnor U13741 (N_13741,N_12786,N_12666);
nand U13742 (N_13742,N_12733,N_12730);
and U13743 (N_13743,N_12986,N_13026);
or U13744 (N_13744,N_13047,N_12919);
or U13745 (N_13745,N_12772,N_13036);
nor U13746 (N_13746,N_12715,N_12888);
nand U13747 (N_13747,N_13058,N_12632);
or U13748 (N_13748,N_13162,N_12747);
or U13749 (N_13749,N_13012,N_12799);
and U13750 (N_13750,N_12684,N_12645);
and U13751 (N_13751,N_12998,N_12948);
and U13752 (N_13752,N_12796,N_12953);
nor U13753 (N_13753,N_12990,N_12961);
xnor U13754 (N_13754,N_12675,N_13188);
nand U13755 (N_13755,N_12634,N_12628);
or U13756 (N_13756,N_12834,N_13163);
xor U13757 (N_13757,N_12747,N_12910);
and U13758 (N_13758,N_13079,N_12933);
xnor U13759 (N_13759,N_12854,N_12711);
nand U13760 (N_13760,N_12743,N_13060);
or U13761 (N_13761,N_12758,N_13023);
or U13762 (N_13762,N_12700,N_12668);
xor U13763 (N_13763,N_12680,N_12739);
and U13764 (N_13764,N_12666,N_12698);
xor U13765 (N_13765,N_13002,N_13114);
nor U13766 (N_13766,N_13017,N_13068);
nand U13767 (N_13767,N_12706,N_13070);
or U13768 (N_13768,N_13031,N_13002);
or U13769 (N_13769,N_12738,N_13180);
and U13770 (N_13770,N_12834,N_13127);
or U13771 (N_13771,N_12852,N_13104);
nand U13772 (N_13772,N_12943,N_12967);
nor U13773 (N_13773,N_12780,N_12995);
and U13774 (N_13774,N_13011,N_13068);
nand U13775 (N_13775,N_13149,N_12964);
or U13776 (N_13776,N_12782,N_12715);
xnor U13777 (N_13777,N_12984,N_13085);
nor U13778 (N_13778,N_13101,N_12986);
xnor U13779 (N_13779,N_13085,N_12856);
and U13780 (N_13780,N_12786,N_12878);
nand U13781 (N_13781,N_12854,N_12940);
or U13782 (N_13782,N_12718,N_12940);
or U13783 (N_13783,N_12959,N_12925);
or U13784 (N_13784,N_13048,N_12976);
and U13785 (N_13785,N_12958,N_12713);
and U13786 (N_13786,N_12680,N_12726);
or U13787 (N_13787,N_13024,N_13011);
nand U13788 (N_13788,N_13124,N_13191);
or U13789 (N_13789,N_13023,N_12905);
and U13790 (N_13790,N_12981,N_13104);
and U13791 (N_13791,N_12944,N_12893);
or U13792 (N_13792,N_13027,N_12625);
nor U13793 (N_13793,N_13006,N_12710);
and U13794 (N_13794,N_13024,N_12842);
and U13795 (N_13795,N_13097,N_12708);
nand U13796 (N_13796,N_13153,N_12654);
nand U13797 (N_13797,N_13172,N_12689);
and U13798 (N_13798,N_12805,N_13167);
nand U13799 (N_13799,N_12838,N_12630);
nand U13800 (N_13800,N_13744,N_13276);
and U13801 (N_13801,N_13631,N_13421);
nor U13802 (N_13802,N_13608,N_13642);
xor U13803 (N_13803,N_13410,N_13296);
and U13804 (N_13804,N_13533,N_13738);
xnor U13805 (N_13805,N_13303,N_13329);
or U13806 (N_13806,N_13536,N_13574);
nor U13807 (N_13807,N_13321,N_13212);
nand U13808 (N_13808,N_13473,N_13632);
or U13809 (N_13809,N_13542,N_13688);
and U13810 (N_13810,N_13352,N_13598);
and U13811 (N_13811,N_13736,N_13555);
nor U13812 (N_13812,N_13780,N_13375);
nand U13813 (N_13813,N_13672,N_13201);
and U13814 (N_13814,N_13205,N_13518);
nand U13815 (N_13815,N_13488,N_13583);
nand U13816 (N_13816,N_13553,N_13753);
nand U13817 (N_13817,N_13378,N_13634);
nor U13818 (N_13818,N_13412,N_13554);
and U13819 (N_13819,N_13589,N_13235);
nor U13820 (N_13820,N_13479,N_13633);
and U13821 (N_13821,N_13575,N_13224);
and U13822 (N_13822,N_13314,N_13728);
xnor U13823 (N_13823,N_13601,N_13717);
nand U13824 (N_13824,N_13743,N_13616);
xnor U13825 (N_13825,N_13415,N_13787);
xnor U13826 (N_13826,N_13770,N_13245);
or U13827 (N_13827,N_13292,N_13648);
or U13828 (N_13828,N_13420,N_13336);
nor U13829 (N_13829,N_13641,N_13316);
nand U13830 (N_13830,N_13539,N_13456);
nand U13831 (N_13831,N_13323,N_13610);
or U13832 (N_13832,N_13541,N_13315);
nand U13833 (N_13833,N_13714,N_13746);
and U13834 (N_13834,N_13291,N_13495);
nor U13835 (N_13835,N_13516,N_13273);
and U13836 (N_13836,N_13401,N_13602);
nand U13837 (N_13837,N_13706,N_13687);
nand U13838 (N_13838,N_13546,N_13644);
xor U13839 (N_13839,N_13763,N_13218);
nor U13840 (N_13840,N_13667,N_13399);
or U13841 (N_13841,N_13288,N_13522);
or U13842 (N_13842,N_13293,N_13766);
and U13843 (N_13843,N_13241,N_13370);
or U13844 (N_13844,N_13573,N_13244);
nor U13845 (N_13845,N_13397,N_13453);
and U13846 (N_13846,N_13376,N_13747);
nor U13847 (N_13847,N_13382,N_13297);
nand U13848 (N_13848,N_13505,N_13446);
and U13849 (N_13849,N_13407,N_13729);
nand U13850 (N_13850,N_13640,N_13263);
or U13851 (N_13851,N_13662,N_13441);
nand U13852 (N_13852,N_13768,N_13423);
and U13853 (N_13853,N_13353,N_13701);
and U13854 (N_13854,N_13210,N_13734);
and U13855 (N_13855,N_13681,N_13796);
or U13856 (N_13856,N_13341,N_13506);
nor U13857 (N_13857,N_13470,N_13585);
nor U13858 (N_13858,N_13285,N_13475);
nor U13859 (N_13859,N_13710,N_13300);
nand U13860 (N_13860,N_13491,N_13777);
nor U13861 (N_13861,N_13481,N_13732);
nor U13862 (N_13862,N_13383,N_13381);
or U13863 (N_13863,N_13695,N_13402);
and U13864 (N_13864,N_13675,N_13607);
nand U13865 (N_13865,N_13236,N_13527);
nor U13866 (N_13866,N_13389,N_13229);
xnor U13867 (N_13867,N_13671,N_13774);
xnor U13868 (N_13868,N_13411,N_13656);
xnor U13869 (N_13869,N_13250,N_13414);
nand U13870 (N_13870,N_13647,N_13448);
nand U13871 (N_13871,N_13689,N_13289);
or U13872 (N_13872,N_13255,N_13438);
or U13873 (N_13873,N_13219,N_13715);
and U13874 (N_13874,N_13424,N_13437);
and U13875 (N_13875,N_13716,N_13617);
or U13876 (N_13876,N_13764,N_13231);
nor U13877 (N_13877,N_13779,N_13708);
and U13878 (N_13878,N_13232,N_13709);
and U13879 (N_13879,N_13760,N_13242);
or U13880 (N_13880,N_13639,N_13317);
xor U13881 (N_13881,N_13624,N_13623);
and U13882 (N_13882,N_13535,N_13545);
nor U13883 (N_13883,N_13429,N_13781);
or U13884 (N_13884,N_13540,N_13347);
and U13885 (N_13885,N_13200,N_13344);
xor U13886 (N_13886,N_13508,N_13304);
xnor U13887 (N_13887,N_13576,N_13691);
nand U13888 (N_13888,N_13275,N_13393);
nand U13889 (N_13889,N_13213,N_13451);
and U13890 (N_13890,N_13579,N_13340);
nor U13891 (N_13891,N_13223,N_13711);
and U13892 (N_13892,N_13374,N_13311);
or U13893 (N_13893,N_13369,N_13472);
and U13894 (N_13894,N_13557,N_13455);
xor U13895 (N_13895,N_13713,N_13512);
and U13896 (N_13896,N_13609,N_13625);
nor U13897 (N_13897,N_13773,N_13400);
or U13898 (N_13898,N_13221,N_13725);
or U13899 (N_13899,N_13595,N_13363);
or U13900 (N_13900,N_13798,N_13325);
nand U13901 (N_13901,N_13504,N_13334);
nand U13902 (N_13902,N_13458,N_13684);
xnor U13903 (N_13903,N_13511,N_13758);
nand U13904 (N_13904,N_13705,N_13605);
or U13905 (N_13905,N_13364,N_13694);
nand U13906 (N_13906,N_13270,N_13570);
and U13907 (N_13907,N_13343,N_13733);
and U13908 (N_13908,N_13251,N_13324);
and U13909 (N_13909,N_13440,N_13449);
and U13910 (N_13910,N_13253,N_13645);
nand U13911 (N_13911,N_13322,N_13745);
nor U13912 (N_13912,N_13700,N_13490);
nor U13913 (N_13913,N_13699,N_13207);
nand U13914 (N_13914,N_13457,N_13281);
nand U13915 (N_13915,N_13597,N_13599);
or U13916 (N_13916,N_13452,N_13749);
and U13917 (N_13917,N_13227,N_13724);
and U13918 (N_13918,N_13283,N_13698);
nor U13919 (N_13919,N_13668,N_13619);
or U13920 (N_13920,N_13445,N_13272);
and U13921 (N_13921,N_13208,N_13404);
or U13922 (N_13922,N_13643,N_13703);
nor U13923 (N_13923,N_13249,N_13372);
nand U13924 (N_13924,N_13433,N_13789);
xor U13925 (N_13925,N_13704,N_13478);
nand U13926 (N_13926,N_13439,N_13266);
nor U13927 (N_13927,N_13556,N_13502);
nor U13928 (N_13928,N_13528,N_13262);
and U13929 (N_13929,N_13564,N_13592);
xnor U13930 (N_13930,N_13509,N_13305);
and U13931 (N_13931,N_13428,N_13767);
nor U13932 (N_13932,N_13307,N_13611);
and U13933 (N_13933,N_13361,N_13447);
nand U13934 (N_13934,N_13791,N_13417);
and U13935 (N_13935,N_13571,N_13216);
or U13936 (N_13936,N_13674,N_13240);
and U13937 (N_13937,N_13515,N_13377);
nand U13938 (N_13938,N_13615,N_13260);
or U13939 (N_13939,N_13566,N_13702);
nor U13940 (N_13940,N_13259,N_13271);
nand U13941 (N_13941,N_13769,N_13351);
nor U13942 (N_13942,N_13718,N_13265);
or U13943 (N_13943,N_13467,N_13432);
and U13944 (N_13944,N_13339,N_13581);
nand U13945 (N_13945,N_13268,N_13604);
and U13946 (N_13946,N_13327,N_13243);
xor U13947 (N_13947,N_13436,N_13355);
nand U13948 (N_13948,N_13471,N_13759);
and U13949 (N_13949,N_13514,N_13477);
xnor U13950 (N_13950,N_13468,N_13345);
or U13951 (N_13951,N_13614,N_13225);
nor U13952 (N_13952,N_13739,N_13434);
nor U13953 (N_13953,N_13299,N_13313);
nor U13954 (N_13954,N_13756,N_13593);
or U13955 (N_13955,N_13498,N_13612);
nor U13956 (N_13956,N_13649,N_13342);
nand U13957 (N_13957,N_13580,N_13572);
nor U13958 (N_13958,N_13679,N_13549);
xor U13959 (N_13959,N_13636,N_13588);
xor U13960 (N_13960,N_13237,N_13408);
or U13961 (N_13961,N_13544,N_13776);
nand U13962 (N_13962,N_13594,N_13652);
and U13963 (N_13963,N_13543,N_13786);
nor U13964 (N_13964,N_13680,N_13395);
xnor U13965 (N_13965,N_13751,N_13409);
or U13966 (N_13966,N_13396,N_13613);
nand U13967 (N_13967,N_13462,N_13220);
nand U13968 (N_13968,N_13469,N_13560);
and U13969 (N_13969,N_13257,N_13228);
nor U13970 (N_13970,N_13525,N_13301);
and U13971 (N_13971,N_13256,N_13782);
or U13972 (N_13972,N_13258,N_13269);
or U13973 (N_13973,N_13627,N_13203);
and U13974 (N_13974,N_13365,N_13772);
nand U13975 (N_13975,N_13577,N_13630);
or U13976 (N_13976,N_13406,N_13320);
or U13977 (N_13977,N_13264,N_13635);
and U13978 (N_13978,N_13444,N_13752);
and U13979 (N_13979,N_13246,N_13394);
or U13980 (N_13980,N_13720,N_13418);
and U13981 (N_13981,N_13480,N_13356);
and U13982 (N_13982,N_13306,N_13357);
nand U13983 (N_13983,N_13463,N_13483);
and U13984 (N_13984,N_13578,N_13510);
nor U13985 (N_13985,N_13214,N_13496);
xnor U13986 (N_13986,N_13665,N_13328);
and U13987 (N_13987,N_13460,N_13657);
nand U13988 (N_13988,N_13308,N_13530);
nand U13989 (N_13989,N_13379,N_13719);
nor U13990 (N_13990,N_13354,N_13692);
or U13991 (N_13991,N_13497,N_13664);
nand U13992 (N_13992,N_13284,N_13559);
nor U13993 (N_13993,N_13712,N_13248);
or U13994 (N_13994,N_13793,N_13425);
nor U13995 (N_13995,N_13792,N_13563);
and U13996 (N_13996,N_13366,N_13215);
nor U13997 (N_13997,N_13252,N_13459);
and U13998 (N_13998,N_13696,N_13678);
nand U13999 (N_13999,N_13443,N_13385);
or U14000 (N_14000,N_13638,N_13690);
and U14001 (N_14001,N_13286,N_13565);
xor U14002 (N_14002,N_13591,N_13280);
or U14003 (N_14003,N_13485,N_13261);
nor U14004 (N_14004,N_13797,N_13517);
xor U14005 (N_14005,N_13741,N_13332);
and U14006 (N_14006,N_13683,N_13750);
nor U14007 (N_14007,N_13360,N_13464);
nand U14008 (N_14008,N_13654,N_13373);
nand U14009 (N_14009,N_13217,N_13621);
nand U14010 (N_14010,N_13461,N_13338);
nand U14011 (N_14011,N_13537,N_13682);
and U14012 (N_14012,N_13333,N_13538);
nor U14013 (N_14013,N_13606,N_13391);
and U14014 (N_14014,N_13465,N_13282);
and U14015 (N_14015,N_13552,N_13788);
nor U14016 (N_14016,N_13659,N_13771);
or U14017 (N_14017,N_13757,N_13513);
xor U14018 (N_14018,N_13666,N_13230);
nor U14019 (N_14019,N_13427,N_13600);
nor U14020 (N_14020,N_13422,N_13287);
xnor U14021 (N_14021,N_13487,N_13474);
nor U14022 (N_14022,N_13295,N_13693);
nand U14023 (N_14023,N_13795,N_13278);
or U14024 (N_14024,N_13646,N_13419);
nand U14025 (N_14025,N_13660,N_13785);
nand U14026 (N_14026,N_13398,N_13524);
or U14027 (N_14027,N_13519,N_13492);
nor U14028 (N_14028,N_13254,N_13442);
and U14029 (N_14029,N_13685,N_13239);
nor U14030 (N_14030,N_13234,N_13661);
or U14031 (N_14031,N_13686,N_13348);
xnor U14032 (N_14032,N_13620,N_13493);
xor U14033 (N_14033,N_13596,N_13392);
or U14034 (N_14034,N_13550,N_13359);
nor U14035 (N_14035,N_13731,N_13310);
or U14036 (N_14036,N_13274,N_13790);
or U14037 (N_14037,N_13318,N_13730);
and U14038 (N_14038,N_13349,N_13558);
nand U14039 (N_14039,N_13294,N_13346);
nand U14040 (N_14040,N_13489,N_13405);
xor U14041 (N_14041,N_13761,N_13722);
nor U14042 (N_14042,N_13486,N_13454);
or U14043 (N_14043,N_13335,N_13551);
nor U14044 (N_14044,N_13426,N_13735);
and U14045 (N_14045,N_13466,N_13450);
or U14046 (N_14046,N_13431,N_13367);
xor U14047 (N_14047,N_13337,N_13507);
nand U14048 (N_14048,N_13529,N_13590);
nor U14049 (N_14049,N_13742,N_13358);
or U14050 (N_14050,N_13204,N_13784);
or U14051 (N_14051,N_13211,N_13775);
nor U14052 (N_14052,N_13721,N_13547);
nand U14053 (N_14053,N_13309,N_13387);
nor U14054 (N_14054,N_13603,N_13503);
nor U14055 (N_14055,N_13302,N_13628);
nor U14056 (N_14056,N_13290,N_13723);
or U14057 (N_14057,N_13676,N_13584);
nor U14058 (N_14058,N_13416,N_13435);
nor U14059 (N_14059,N_13319,N_13568);
or U14060 (N_14060,N_13482,N_13569);
or U14061 (N_14061,N_13655,N_13561);
nor U14062 (N_14062,N_13587,N_13726);
nand U14063 (N_14063,N_13238,N_13388);
nor U14064 (N_14064,N_13567,N_13484);
or U14065 (N_14065,N_13737,N_13520);
xnor U14066 (N_14066,N_13476,N_13740);
nor U14067 (N_14067,N_13362,N_13390);
or U14068 (N_14068,N_13673,N_13765);
nor U14069 (N_14069,N_13755,N_13622);
nand U14070 (N_14070,N_13626,N_13298);
and U14071 (N_14071,N_13526,N_13748);
nand U14072 (N_14072,N_13586,N_13233);
or U14073 (N_14073,N_13658,N_13430);
nand U14074 (N_14074,N_13279,N_13380);
and U14075 (N_14075,N_13629,N_13618);
nor U14076 (N_14076,N_13697,N_13209);
nor U14077 (N_14077,N_13727,N_13521);
or U14078 (N_14078,N_13562,N_13371);
nand U14079 (N_14079,N_13670,N_13226);
xnor U14080 (N_14080,N_13202,N_13330);
or U14081 (N_14081,N_13794,N_13762);
and U14082 (N_14082,N_13501,N_13206);
or U14083 (N_14083,N_13582,N_13386);
or U14084 (N_14084,N_13267,N_13783);
nand U14085 (N_14085,N_13778,N_13494);
and U14086 (N_14086,N_13222,N_13413);
nor U14087 (N_14087,N_13277,N_13653);
nand U14088 (N_14088,N_13523,N_13663);
or U14089 (N_14089,N_13499,N_13531);
nor U14090 (N_14090,N_13500,N_13650);
xor U14091 (N_14091,N_13754,N_13707);
or U14092 (N_14092,N_13331,N_13651);
nand U14093 (N_14093,N_13534,N_13350);
and U14094 (N_14094,N_13548,N_13247);
or U14095 (N_14095,N_13799,N_13669);
nand U14096 (N_14096,N_13637,N_13368);
and U14097 (N_14097,N_13326,N_13677);
nand U14098 (N_14098,N_13403,N_13384);
xor U14099 (N_14099,N_13312,N_13532);
xnor U14100 (N_14100,N_13729,N_13210);
nor U14101 (N_14101,N_13247,N_13682);
or U14102 (N_14102,N_13576,N_13253);
xor U14103 (N_14103,N_13321,N_13439);
or U14104 (N_14104,N_13566,N_13710);
or U14105 (N_14105,N_13676,N_13402);
xnor U14106 (N_14106,N_13563,N_13326);
or U14107 (N_14107,N_13640,N_13428);
nor U14108 (N_14108,N_13243,N_13385);
and U14109 (N_14109,N_13291,N_13776);
nor U14110 (N_14110,N_13236,N_13625);
nand U14111 (N_14111,N_13220,N_13612);
nor U14112 (N_14112,N_13702,N_13309);
nor U14113 (N_14113,N_13400,N_13675);
nor U14114 (N_14114,N_13360,N_13791);
nor U14115 (N_14115,N_13546,N_13589);
or U14116 (N_14116,N_13715,N_13557);
nor U14117 (N_14117,N_13794,N_13248);
nand U14118 (N_14118,N_13678,N_13679);
nand U14119 (N_14119,N_13580,N_13449);
and U14120 (N_14120,N_13727,N_13347);
and U14121 (N_14121,N_13515,N_13593);
nor U14122 (N_14122,N_13618,N_13413);
and U14123 (N_14123,N_13348,N_13557);
nand U14124 (N_14124,N_13323,N_13603);
xnor U14125 (N_14125,N_13575,N_13674);
and U14126 (N_14126,N_13711,N_13289);
or U14127 (N_14127,N_13544,N_13374);
nand U14128 (N_14128,N_13454,N_13605);
and U14129 (N_14129,N_13604,N_13776);
and U14130 (N_14130,N_13610,N_13434);
and U14131 (N_14131,N_13392,N_13316);
nand U14132 (N_14132,N_13418,N_13646);
or U14133 (N_14133,N_13226,N_13580);
nand U14134 (N_14134,N_13290,N_13355);
xnor U14135 (N_14135,N_13543,N_13752);
nand U14136 (N_14136,N_13685,N_13494);
and U14137 (N_14137,N_13796,N_13693);
nor U14138 (N_14138,N_13298,N_13268);
and U14139 (N_14139,N_13551,N_13487);
and U14140 (N_14140,N_13350,N_13207);
nor U14141 (N_14141,N_13461,N_13382);
and U14142 (N_14142,N_13701,N_13237);
xor U14143 (N_14143,N_13432,N_13374);
nand U14144 (N_14144,N_13367,N_13292);
nand U14145 (N_14145,N_13431,N_13525);
nand U14146 (N_14146,N_13693,N_13218);
nand U14147 (N_14147,N_13567,N_13681);
nor U14148 (N_14148,N_13732,N_13574);
nor U14149 (N_14149,N_13538,N_13246);
nor U14150 (N_14150,N_13749,N_13355);
nand U14151 (N_14151,N_13236,N_13461);
nor U14152 (N_14152,N_13372,N_13291);
and U14153 (N_14153,N_13423,N_13721);
and U14154 (N_14154,N_13750,N_13588);
or U14155 (N_14155,N_13311,N_13781);
nor U14156 (N_14156,N_13671,N_13553);
nor U14157 (N_14157,N_13227,N_13424);
nor U14158 (N_14158,N_13599,N_13769);
nor U14159 (N_14159,N_13494,N_13385);
nand U14160 (N_14160,N_13681,N_13725);
or U14161 (N_14161,N_13201,N_13771);
nand U14162 (N_14162,N_13781,N_13631);
nor U14163 (N_14163,N_13744,N_13618);
xnor U14164 (N_14164,N_13797,N_13583);
nand U14165 (N_14165,N_13589,N_13507);
xnor U14166 (N_14166,N_13250,N_13321);
nor U14167 (N_14167,N_13780,N_13677);
and U14168 (N_14168,N_13437,N_13400);
nor U14169 (N_14169,N_13244,N_13206);
nor U14170 (N_14170,N_13738,N_13264);
or U14171 (N_14171,N_13234,N_13725);
nand U14172 (N_14172,N_13617,N_13593);
nand U14173 (N_14173,N_13325,N_13529);
xnor U14174 (N_14174,N_13536,N_13449);
nor U14175 (N_14175,N_13439,N_13437);
nand U14176 (N_14176,N_13792,N_13476);
or U14177 (N_14177,N_13762,N_13657);
and U14178 (N_14178,N_13696,N_13646);
nor U14179 (N_14179,N_13242,N_13243);
or U14180 (N_14180,N_13223,N_13650);
nand U14181 (N_14181,N_13567,N_13640);
xor U14182 (N_14182,N_13403,N_13291);
and U14183 (N_14183,N_13396,N_13442);
and U14184 (N_14184,N_13566,N_13626);
or U14185 (N_14185,N_13557,N_13223);
and U14186 (N_14186,N_13228,N_13685);
nor U14187 (N_14187,N_13253,N_13506);
and U14188 (N_14188,N_13327,N_13493);
nor U14189 (N_14189,N_13551,N_13323);
and U14190 (N_14190,N_13360,N_13722);
or U14191 (N_14191,N_13410,N_13384);
xnor U14192 (N_14192,N_13593,N_13407);
and U14193 (N_14193,N_13378,N_13338);
or U14194 (N_14194,N_13692,N_13368);
nand U14195 (N_14195,N_13617,N_13773);
nand U14196 (N_14196,N_13335,N_13610);
and U14197 (N_14197,N_13347,N_13402);
nor U14198 (N_14198,N_13756,N_13788);
or U14199 (N_14199,N_13258,N_13389);
nor U14200 (N_14200,N_13708,N_13603);
or U14201 (N_14201,N_13266,N_13282);
nand U14202 (N_14202,N_13768,N_13760);
and U14203 (N_14203,N_13695,N_13361);
or U14204 (N_14204,N_13329,N_13201);
or U14205 (N_14205,N_13250,N_13621);
or U14206 (N_14206,N_13450,N_13420);
and U14207 (N_14207,N_13467,N_13564);
nor U14208 (N_14208,N_13325,N_13691);
xnor U14209 (N_14209,N_13688,N_13519);
and U14210 (N_14210,N_13730,N_13384);
or U14211 (N_14211,N_13529,N_13279);
or U14212 (N_14212,N_13498,N_13394);
or U14213 (N_14213,N_13292,N_13452);
nand U14214 (N_14214,N_13640,N_13269);
nor U14215 (N_14215,N_13735,N_13774);
and U14216 (N_14216,N_13762,N_13635);
or U14217 (N_14217,N_13350,N_13669);
or U14218 (N_14218,N_13517,N_13767);
nand U14219 (N_14219,N_13309,N_13215);
nor U14220 (N_14220,N_13368,N_13259);
or U14221 (N_14221,N_13586,N_13331);
or U14222 (N_14222,N_13556,N_13781);
nor U14223 (N_14223,N_13683,N_13463);
nor U14224 (N_14224,N_13298,N_13639);
or U14225 (N_14225,N_13610,N_13290);
nor U14226 (N_14226,N_13780,N_13399);
or U14227 (N_14227,N_13748,N_13432);
or U14228 (N_14228,N_13417,N_13524);
nor U14229 (N_14229,N_13294,N_13394);
nor U14230 (N_14230,N_13626,N_13232);
or U14231 (N_14231,N_13404,N_13402);
or U14232 (N_14232,N_13606,N_13214);
and U14233 (N_14233,N_13563,N_13534);
xnor U14234 (N_14234,N_13232,N_13419);
or U14235 (N_14235,N_13345,N_13372);
or U14236 (N_14236,N_13354,N_13465);
nor U14237 (N_14237,N_13539,N_13583);
xor U14238 (N_14238,N_13431,N_13601);
and U14239 (N_14239,N_13289,N_13634);
and U14240 (N_14240,N_13355,N_13495);
nand U14241 (N_14241,N_13549,N_13530);
nand U14242 (N_14242,N_13630,N_13721);
nor U14243 (N_14243,N_13607,N_13679);
nand U14244 (N_14244,N_13758,N_13389);
and U14245 (N_14245,N_13340,N_13639);
nand U14246 (N_14246,N_13653,N_13771);
nor U14247 (N_14247,N_13463,N_13711);
or U14248 (N_14248,N_13401,N_13790);
nand U14249 (N_14249,N_13670,N_13332);
nand U14250 (N_14250,N_13619,N_13504);
nor U14251 (N_14251,N_13329,N_13434);
nor U14252 (N_14252,N_13452,N_13647);
and U14253 (N_14253,N_13770,N_13280);
and U14254 (N_14254,N_13515,N_13767);
xor U14255 (N_14255,N_13677,N_13407);
nand U14256 (N_14256,N_13279,N_13500);
nor U14257 (N_14257,N_13511,N_13264);
and U14258 (N_14258,N_13231,N_13322);
or U14259 (N_14259,N_13323,N_13748);
nand U14260 (N_14260,N_13499,N_13474);
nor U14261 (N_14261,N_13206,N_13641);
nand U14262 (N_14262,N_13497,N_13765);
nor U14263 (N_14263,N_13571,N_13253);
or U14264 (N_14264,N_13499,N_13622);
or U14265 (N_14265,N_13407,N_13564);
nor U14266 (N_14266,N_13451,N_13301);
xor U14267 (N_14267,N_13322,N_13763);
xnor U14268 (N_14268,N_13645,N_13515);
and U14269 (N_14269,N_13748,N_13274);
nand U14270 (N_14270,N_13772,N_13418);
xnor U14271 (N_14271,N_13608,N_13385);
nand U14272 (N_14272,N_13793,N_13512);
nand U14273 (N_14273,N_13335,N_13628);
or U14274 (N_14274,N_13594,N_13680);
nand U14275 (N_14275,N_13799,N_13759);
or U14276 (N_14276,N_13436,N_13242);
and U14277 (N_14277,N_13478,N_13451);
or U14278 (N_14278,N_13548,N_13274);
and U14279 (N_14279,N_13281,N_13435);
nand U14280 (N_14280,N_13747,N_13748);
nand U14281 (N_14281,N_13405,N_13544);
or U14282 (N_14282,N_13370,N_13724);
nor U14283 (N_14283,N_13667,N_13461);
nand U14284 (N_14284,N_13675,N_13444);
or U14285 (N_14285,N_13752,N_13428);
or U14286 (N_14286,N_13495,N_13729);
nand U14287 (N_14287,N_13332,N_13596);
and U14288 (N_14288,N_13551,N_13480);
or U14289 (N_14289,N_13594,N_13627);
nand U14290 (N_14290,N_13603,N_13362);
and U14291 (N_14291,N_13333,N_13417);
xnor U14292 (N_14292,N_13328,N_13584);
or U14293 (N_14293,N_13409,N_13509);
or U14294 (N_14294,N_13368,N_13649);
nor U14295 (N_14295,N_13652,N_13568);
or U14296 (N_14296,N_13279,N_13503);
nand U14297 (N_14297,N_13391,N_13464);
nand U14298 (N_14298,N_13588,N_13468);
nor U14299 (N_14299,N_13493,N_13711);
nand U14300 (N_14300,N_13333,N_13640);
and U14301 (N_14301,N_13605,N_13336);
and U14302 (N_14302,N_13667,N_13385);
nor U14303 (N_14303,N_13352,N_13524);
or U14304 (N_14304,N_13287,N_13318);
nor U14305 (N_14305,N_13667,N_13589);
and U14306 (N_14306,N_13583,N_13573);
or U14307 (N_14307,N_13237,N_13227);
and U14308 (N_14308,N_13630,N_13239);
and U14309 (N_14309,N_13364,N_13478);
or U14310 (N_14310,N_13512,N_13474);
nand U14311 (N_14311,N_13222,N_13519);
nand U14312 (N_14312,N_13335,N_13580);
nor U14313 (N_14313,N_13746,N_13260);
or U14314 (N_14314,N_13543,N_13411);
nor U14315 (N_14315,N_13748,N_13452);
nand U14316 (N_14316,N_13587,N_13688);
and U14317 (N_14317,N_13487,N_13320);
or U14318 (N_14318,N_13566,N_13784);
nand U14319 (N_14319,N_13695,N_13375);
xnor U14320 (N_14320,N_13625,N_13493);
nor U14321 (N_14321,N_13454,N_13495);
or U14322 (N_14322,N_13255,N_13563);
nand U14323 (N_14323,N_13517,N_13330);
or U14324 (N_14324,N_13397,N_13556);
or U14325 (N_14325,N_13510,N_13343);
or U14326 (N_14326,N_13358,N_13628);
or U14327 (N_14327,N_13549,N_13738);
nor U14328 (N_14328,N_13405,N_13412);
or U14329 (N_14329,N_13547,N_13743);
or U14330 (N_14330,N_13271,N_13737);
nand U14331 (N_14331,N_13470,N_13245);
nor U14332 (N_14332,N_13222,N_13383);
nand U14333 (N_14333,N_13368,N_13223);
or U14334 (N_14334,N_13339,N_13243);
or U14335 (N_14335,N_13762,N_13391);
and U14336 (N_14336,N_13442,N_13506);
or U14337 (N_14337,N_13714,N_13627);
and U14338 (N_14338,N_13220,N_13490);
nand U14339 (N_14339,N_13591,N_13631);
or U14340 (N_14340,N_13613,N_13379);
or U14341 (N_14341,N_13224,N_13556);
or U14342 (N_14342,N_13291,N_13762);
nor U14343 (N_14343,N_13509,N_13783);
nor U14344 (N_14344,N_13224,N_13436);
or U14345 (N_14345,N_13770,N_13688);
nor U14346 (N_14346,N_13738,N_13510);
or U14347 (N_14347,N_13406,N_13208);
nand U14348 (N_14348,N_13566,N_13214);
nand U14349 (N_14349,N_13439,N_13765);
nor U14350 (N_14350,N_13430,N_13660);
nand U14351 (N_14351,N_13306,N_13734);
nand U14352 (N_14352,N_13445,N_13252);
or U14353 (N_14353,N_13469,N_13571);
xor U14354 (N_14354,N_13729,N_13459);
and U14355 (N_14355,N_13206,N_13496);
and U14356 (N_14356,N_13327,N_13299);
nand U14357 (N_14357,N_13381,N_13352);
nand U14358 (N_14358,N_13412,N_13625);
and U14359 (N_14359,N_13795,N_13285);
xor U14360 (N_14360,N_13676,N_13564);
nand U14361 (N_14361,N_13647,N_13544);
and U14362 (N_14362,N_13418,N_13243);
or U14363 (N_14363,N_13652,N_13431);
nand U14364 (N_14364,N_13360,N_13723);
and U14365 (N_14365,N_13710,N_13532);
and U14366 (N_14366,N_13354,N_13458);
nand U14367 (N_14367,N_13619,N_13696);
or U14368 (N_14368,N_13783,N_13690);
nor U14369 (N_14369,N_13215,N_13754);
nor U14370 (N_14370,N_13404,N_13345);
nor U14371 (N_14371,N_13321,N_13672);
or U14372 (N_14372,N_13350,N_13662);
or U14373 (N_14373,N_13485,N_13305);
and U14374 (N_14374,N_13423,N_13661);
and U14375 (N_14375,N_13212,N_13369);
xnor U14376 (N_14376,N_13307,N_13767);
and U14377 (N_14377,N_13586,N_13228);
or U14378 (N_14378,N_13238,N_13417);
or U14379 (N_14379,N_13444,N_13332);
nand U14380 (N_14380,N_13454,N_13479);
nand U14381 (N_14381,N_13226,N_13560);
nand U14382 (N_14382,N_13613,N_13731);
and U14383 (N_14383,N_13773,N_13770);
nand U14384 (N_14384,N_13679,N_13478);
or U14385 (N_14385,N_13591,N_13744);
nand U14386 (N_14386,N_13714,N_13282);
nand U14387 (N_14387,N_13411,N_13377);
xor U14388 (N_14388,N_13750,N_13715);
and U14389 (N_14389,N_13718,N_13732);
nor U14390 (N_14390,N_13418,N_13316);
and U14391 (N_14391,N_13796,N_13341);
nand U14392 (N_14392,N_13462,N_13293);
xor U14393 (N_14393,N_13718,N_13539);
or U14394 (N_14394,N_13410,N_13766);
and U14395 (N_14395,N_13716,N_13634);
and U14396 (N_14396,N_13661,N_13644);
or U14397 (N_14397,N_13260,N_13412);
nor U14398 (N_14398,N_13744,N_13297);
nor U14399 (N_14399,N_13590,N_13640);
nand U14400 (N_14400,N_14054,N_14347);
and U14401 (N_14401,N_14046,N_14114);
or U14402 (N_14402,N_13979,N_13974);
nand U14403 (N_14403,N_14154,N_14051);
nand U14404 (N_14404,N_14183,N_14366);
nand U14405 (N_14405,N_14181,N_14277);
and U14406 (N_14406,N_13839,N_14136);
nand U14407 (N_14407,N_14061,N_13928);
and U14408 (N_14408,N_13814,N_13978);
and U14409 (N_14409,N_14396,N_13903);
or U14410 (N_14410,N_14392,N_14036);
nor U14411 (N_14411,N_13827,N_13890);
nand U14412 (N_14412,N_14211,N_14335);
and U14413 (N_14413,N_14151,N_14263);
and U14414 (N_14414,N_14291,N_14297);
and U14415 (N_14415,N_14340,N_13894);
nand U14416 (N_14416,N_14397,N_14106);
or U14417 (N_14417,N_14039,N_13817);
nor U14418 (N_14418,N_14125,N_13924);
nor U14419 (N_14419,N_13962,N_13819);
nand U14420 (N_14420,N_14091,N_14180);
or U14421 (N_14421,N_14315,N_14285);
xnor U14422 (N_14422,N_14187,N_13923);
nor U14423 (N_14423,N_14327,N_14073);
nand U14424 (N_14424,N_14049,N_14065);
nor U14425 (N_14425,N_14165,N_14213);
and U14426 (N_14426,N_14113,N_14306);
nand U14427 (N_14427,N_13981,N_14055);
xnor U14428 (N_14428,N_14273,N_14123);
nand U14429 (N_14429,N_14178,N_14354);
nor U14430 (N_14430,N_13970,N_14115);
nor U14431 (N_14431,N_14122,N_14271);
nor U14432 (N_14432,N_14393,N_13805);
xnor U14433 (N_14433,N_14184,N_13977);
nor U14434 (N_14434,N_14008,N_14153);
nor U14435 (N_14435,N_14117,N_14133);
and U14436 (N_14436,N_13893,N_14339);
and U14437 (N_14437,N_14244,N_14171);
nand U14438 (N_14438,N_13946,N_14363);
xnor U14439 (N_14439,N_13874,N_13991);
xor U14440 (N_14440,N_14386,N_13863);
nor U14441 (N_14441,N_14215,N_14032);
and U14442 (N_14442,N_13919,N_14116);
or U14443 (N_14443,N_14163,N_14224);
or U14444 (N_14444,N_14161,N_13899);
nand U14445 (N_14445,N_13889,N_13994);
nand U14446 (N_14446,N_13956,N_14089);
and U14447 (N_14447,N_14290,N_14103);
and U14448 (N_14448,N_13950,N_14302);
or U14449 (N_14449,N_13948,N_14310);
or U14450 (N_14450,N_14127,N_14236);
or U14451 (N_14451,N_14353,N_14390);
and U14452 (N_14452,N_13824,N_13808);
or U14453 (N_14453,N_14398,N_14084);
xnor U14454 (N_14454,N_14012,N_13968);
nor U14455 (N_14455,N_14167,N_14110);
xor U14456 (N_14456,N_13828,N_14368);
nand U14457 (N_14457,N_14026,N_14319);
nor U14458 (N_14458,N_14331,N_14197);
xor U14459 (N_14459,N_14194,N_14275);
xnor U14460 (N_14460,N_14253,N_14289);
and U14461 (N_14461,N_14262,N_14040);
nand U14462 (N_14462,N_13897,N_14121);
nor U14463 (N_14463,N_14160,N_14070);
nand U14464 (N_14464,N_14268,N_13856);
nor U14465 (N_14465,N_14332,N_14030);
xnor U14466 (N_14466,N_14149,N_14225);
or U14467 (N_14467,N_14217,N_14349);
or U14468 (N_14468,N_14048,N_14204);
nand U14469 (N_14469,N_13915,N_13975);
or U14470 (N_14470,N_14371,N_14013);
and U14471 (N_14471,N_13826,N_14296);
nor U14472 (N_14472,N_13912,N_13884);
and U14473 (N_14473,N_14345,N_14308);
and U14474 (N_14474,N_14240,N_14232);
or U14475 (N_14475,N_13848,N_14090);
or U14476 (N_14476,N_14237,N_14083);
nand U14477 (N_14477,N_13957,N_14248);
nand U14478 (N_14478,N_13810,N_14064);
and U14479 (N_14479,N_14017,N_13988);
nor U14480 (N_14480,N_13803,N_13844);
and U14481 (N_14481,N_13896,N_13905);
xor U14482 (N_14482,N_14269,N_13875);
nor U14483 (N_14483,N_14135,N_13845);
or U14484 (N_14484,N_14042,N_13992);
nor U14485 (N_14485,N_13886,N_13870);
nand U14486 (N_14486,N_14259,N_14157);
and U14487 (N_14487,N_14364,N_14071);
or U14488 (N_14488,N_13813,N_14260);
or U14489 (N_14489,N_14313,N_13971);
xnor U14490 (N_14490,N_14148,N_13842);
xor U14491 (N_14491,N_14112,N_14241);
nand U14492 (N_14492,N_14309,N_14074);
nor U14493 (N_14493,N_14022,N_14399);
nand U14494 (N_14494,N_14311,N_14384);
or U14495 (N_14495,N_13857,N_14230);
nand U14496 (N_14496,N_13840,N_14214);
nand U14497 (N_14497,N_14174,N_14261);
nand U14498 (N_14498,N_14068,N_13822);
nand U14499 (N_14499,N_13949,N_14201);
or U14500 (N_14500,N_13829,N_14119);
and U14501 (N_14501,N_14179,N_14147);
and U14502 (N_14502,N_14283,N_14281);
and U14503 (N_14503,N_14189,N_13902);
xnor U14504 (N_14504,N_14028,N_14050);
nand U14505 (N_14505,N_14303,N_13849);
nand U14506 (N_14506,N_14295,N_14362);
and U14507 (N_14507,N_13885,N_14239);
or U14508 (N_14508,N_14218,N_14359);
or U14509 (N_14509,N_14190,N_14338);
nor U14510 (N_14510,N_13914,N_14058);
or U14511 (N_14511,N_13821,N_13843);
xnor U14512 (N_14512,N_14124,N_13997);
nor U14513 (N_14513,N_14120,N_13982);
nand U14514 (N_14514,N_13831,N_14280);
or U14515 (N_14515,N_14342,N_14382);
or U14516 (N_14516,N_14229,N_14082);
xor U14517 (N_14517,N_13910,N_13804);
nand U14518 (N_14518,N_14041,N_14069);
nand U14519 (N_14519,N_14209,N_14254);
and U14520 (N_14520,N_14235,N_14100);
nand U14521 (N_14521,N_13887,N_14249);
and U14522 (N_14522,N_14140,N_14192);
nor U14523 (N_14523,N_14238,N_13920);
or U14524 (N_14524,N_13969,N_14387);
nand U14525 (N_14525,N_13999,N_14044);
or U14526 (N_14526,N_13963,N_14144);
nand U14527 (N_14527,N_14098,N_14333);
nor U14528 (N_14528,N_13942,N_14219);
nand U14529 (N_14529,N_14316,N_14169);
and U14530 (N_14530,N_14250,N_13904);
nor U14531 (N_14531,N_14267,N_14326);
or U14532 (N_14532,N_14029,N_13906);
or U14533 (N_14533,N_14001,N_13941);
nor U14534 (N_14534,N_13983,N_14128);
or U14535 (N_14535,N_13931,N_13867);
or U14536 (N_14536,N_14337,N_14130);
nand U14537 (N_14537,N_13864,N_13871);
xnor U14538 (N_14538,N_14199,N_14270);
nand U14539 (N_14539,N_13945,N_14168);
and U14540 (N_14540,N_14023,N_14137);
or U14541 (N_14541,N_14216,N_14314);
and U14542 (N_14542,N_14057,N_14279);
nand U14543 (N_14543,N_13823,N_13850);
or U14544 (N_14544,N_14099,N_13913);
xor U14545 (N_14545,N_13800,N_14336);
xnor U14546 (N_14546,N_14186,N_14019);
and U14547 (N_14547,N_14195,N_13891);
and U14548 (N_14548,N_14207,N_14198);
or U14549 (N_14549,N_14079,N_14107);
and U14550 (N_14550,N_13820,N_14380);
or U14551 (N_14551,N_14294,N_14377);
nand U14552 (N_14552,N_14258,N_14334);
and U14553 (N_14553,N_13853,N_14143);
nand U14554 (N_14554,N_14251,N_14274);
nand U14555 (N_14555,N_14378,N_13955);
nand U14556 (N_14556,N_13985,N_14206);
nand U14557 (N_14557,N_14227,N_13812);
and U14558 (N_14558,N_13989,N_14093);
nor U14559 (N_14559,N_13938,N_14104);
or U14560 (N_14560,N_14142,N_13926);
and U14561 (N_14561,N_14220,N_13818);
xnor U14562 (N_14562,N_13900,N_13965);
or U14563 (N_14563,N_13837,N_13862);
xor U14564 (N_14564,N_14231,N_14286);
or U14565 (N_14565,N_14328,N_13901);
and U14566 (N_14566,N_14150,N_14101);
or U14567 (N_14567,N_13860,N_14242);
and U14568 (N_14568,N_14323,N_14222);
or U14569 (N_14569,N_14221,N_14329);
nor U14570 (N_14570,N_14395,N_14006);
xor U14571 (N_14571,N_14004,N_14086);
xor U14572 (N_14572,N_14246,N_14139);
and U14573 (N_14573,N_14360,N_13881);
or U14574 (N_14574,N_14045,N_14072);
nand U14575 (N_14575,N_14027,N_14391);
nor U14576 (N_14576,N_14374,N_13882);
or U14577 (N_14577,N_14191,N_13951);
nor U14578 (N_14578,N_13972,N_13833);
or U14579 (N_14579,N_14053,N_14155);
nand U14580 (N_14580,N_14379,N_13939);
or U14581 (N_14581,N_14292,N_14376);
xnor U14582 (N_14582,N_14322,N_14152);
or U14583 (N_14583,N_14358,N_13876);
xor U14584 (N_14584,N_14059,N_14385);
and U14585 (N_14585,N_13940,N_14164);
nand U14586 (N_14586,N_14208,N_14000);
xnor U14587 (N_14587,N_13967,N_14272);
nor U14588 (N_14588,N_14043,N_14188);
and U14589 (N_14589,N_14011,N_13835);
nor U14590 (N_14590,N_13851,N_13916);
nor U14591 (N_14591,N_13838,N_13855);
and U14592 (N_14592,N_14038,N_13937);
xor U14593 (N_14593,N_13934,N_14252);
nor U14594 (N_14594,N_14005,N_14346);
nor U14595 (N_14595,N_14202,N_14034);
or U14596 (N_14596,N_14076,N_14126);
xnor U14597 (N_14597,N_14365,N_14330);
or U14598 (N_14598,N_14352,N_14146);
or U14599 (N_14599,N_14276,N_14300);
nor U14600 (N_14600,N_13976,N_14344);
nor U14601 (N_14601,N_13952,N_14243);
or U14602 (N_14602,N_13869,N_13861);
or U14603 (N_14603,N_13960,N_14020);
or U14604 (N_14604,N_13866,N_14321);
nand U14605 (N_14605,N_13917,N_13815);
nand U14606 (N_14606,N_13879,N_13868);
nand U14607 (N_14607,N_14324,N_14356);
or U14608 (N_14608,N_14037,N_14348);
nor U14609 (N_14609,N_14373,N_14255);
or U14610 (N_14610,N_13947,N_14095);
and U14611 (N_14611,N_14233,N_14318);
nand U14612 (N_14612,N_14088,N_13880);
or U14613 (N_14613,N_14031,N_14185);
nor U14614 (N_14614,N_14293,N_14307);
and U14615 (N_14615,N_14381,N_13841);
and U14616 (N_14616,N_13898,N_14355);
or U14617 (N_14617,N_13921,N_13980);
nand U14618 (N_14618,N_14228,N_14375);
and U14619 (N_14619,N_14284,N_14035);
nor U14620 (N_14620,N_14141,N_14021);
nor U14621 (N_14621,N_14193,N_13966);
xor U14622 (N_14622,N_14096,N_14247);
nor U14623 (N_14623,N_13959,N_13933);
and U14624 (N_14624,N_14223,N_13922);
nand U14625 (N_14625,N_13801,N_14305);
nand U14626 (N_14626,N_13892,N_13908);
nor U14627 (N_14627,N_14265,N_13935);
nor U14628 (N_14628,N_14003,N_14389);
nand U14629 (N_14629,N_14172,N_14092);
nand U14630 (N_14630,N_13936,N_13929);
nand U14631 (N_14631,N_14010,N_13825);
and U14632 (N_14632,N_14009,N_14288);
xor U14633 (N_14633,N_13809,N_14094);
or U14634 (N_14634,N_13859,N_14033);
nor U14635 (N_14635,N_14075,N_14388);
or U14636 (N_14636,N_13984,N_13953);
xor U14637 (N_14637,N_13807,N_14234);
nand U14638 (N_14638,N_14138,N_14298);
nor U14639 (N_14639,N_14081,N_14047);
and U14640 (N_14640,N_14087,N_14097);
nor U14641 (N_14641,N_14361,N_14085);
nor U14642 (N_14642,N_13932,N_14024);
xor U14643 (N_14643,N_13990,N_13996);
or U14644 (N_14644,N_14018,N_14257);
nor U14645 (N_14645,N_13943,N_13944);
and U14646 (N_14646,N_14016,N_14299);
nor U14647 (N_14647,N_14205,N_13973);
or U14648 (N_14648,N_14301,N_14109);
or U14649 (N_14649,N_14166,N_14264);
or U14650 (N_14650,N_14156,N_14182);
xnor U14651 (N_14651,N_14025,N_14370);
nand U14652 (N_14652,N_14266,N_13909);
and U14653 (N_14653,N_13873,N_13986);
nand U14654 (N_14654,N_13918,N_14304);
nor U14655 (N_14655,N_14367,N_13888);
xor U14656 (N_14656,N_14325,N_14350);
nor U14657 (N_14657,N_14200,N_13927);
or U14658 (N_14658,N_14278,N_14317);
nand U14659 (N_14659,N_14145,N_13836);
nand U14660 (N_14660,N_14063,N_14177);
nand U14661 (N_14661,N_14210,N_14014);
xor U14662 (N_14662,N_14256,N_14056);
and U14663 (N_14663,N_14062,N_13964);
and U14664 (N_14664,N_14357,N_14312);
nand U14665 (N_14665,N_13907,N_14102);
or U14666 (N_14666,N_13834,N_14111);
and U14667 (N_14667,N_13878,N_13847);
and U14668 (N_14668,N_14078,N_14052);
xor U14669 (N_14669,N_13895,N_14077);
and U14670 (N_14670,N_14196,N_13911);
nor U14671 (N_14671,N_13954,N_14343);
xor U14672 (N_14672,N_13806,N_14170);
nand U14673 (N_14673,N_14060,N_13930);
and U14674 (N_14674,N_14067,N_14383);
nor U14675 (N_14675,N_13858,N_14212);
nand U14676 (N_14676,N_13802,N_14129);
xnor U14677 (N_14677,N_14176,N_14320);
nor U14678 (N_14678,N_13998,N_14341);
nor U14679 (N_14679,N_14282,N_14351);
and U14680 (N_14680,N_13811,N_14203);
nor U14681 (N_14681,N_13993,N_14369);
and U14682 (N_14682,N_13987,N_14162);
or U14683 (N_14683,N_14287,N_13832);
nor U14684 (N_14684,N_14173,N_13877);
and U14685 (N_14685,N_13846,N_13925);
nand U14686 (N_14686,N_14394,N_14245);
nor U14687 (N_14687,N_14105,N_14132);
nor U14688 (N_14688,N_14226,N_14158);
and U14689 (N_14689,N_14007,N_14159);
and U14690 (N_14690,N_14108,N_13830);
or U14691 (N_14691,N_13883,N_14175);
and U14692 (N_14692,N_13816,N_14066);
or U14693 (N_14693,N_14015,N_13854);
nand U14694 (N_14694,N_13852,N_14134);
xor U14695 (N_14695,N_13961,N_14118);
or U14696 (N_14696,N_13872,N_14002);
nor U14697 (N_14697,N_13958,N_13865);
and U14698 (N_14698,N_13995,N_14131);
or U14699 (N_14699,N_14080,N_14372);
or U14700 (N_14700,N_13861,N_13939);
xor U14701 (N_14701,N_14358,N_14323);
or U14702 (N_14702,N_14293,N_14256);
nor U14703 (N_14703,N_13817,N_13997);
and U14704 (N_14704,N_14339,N_13890);
nand U14705 (N_14705,N_14280,N_14252);
xor U14706 (N_14706,N_13956,N_14183);
and U14707 (N_14707,N_14271,N_14184);
or U14708 (N_14708,N_14354,N_13853);
or U14709 (N_14709,N_13850,N_13948);
nor U14710 (N_14710,N_13877,N_13933);
or U14711 (N_14711,N_13831,N_14191);
and U14712 (N_14712,N_13847,N_14102);
and U14713 (N_14713,N_14256,N_14040);
and U14714 (N_14714,N_14044,N_14202);
and U14715 (N_14715,N_13930,N_14231);
and U14716 (N_14716,N_14089,N_14263);
nand U14717 (N_14717,N_13873,N_14314);
nor U14718 (N_14718,N_14191,N_14063);
xnor U14719 (N_14719,N_13867,N_14336);
xnor U14720 (N_14720,N_13968,N_14265);
nand U14721 (N_14721,N_14214,N_14089);
or U14722 (N_14722,N_14131,N_14056);
or U14723 (N_14723,N_14162,N_14252);
and U14724 (N_14724,N_14339,N_14118);
and U14725 (N_14725,N_13891,N_14243);
and U14726 (N_14726,N_14361,N_13946);
and U14727 (N_14727,N_13844,N_13954);
and U14728 (N_14728,N_14138,N_14059);
nor U14729 (N_14729,N_14140,N_14256);
nor U14730 (N_14730,N_13817,N_14062);
nor U14731 (N_14731,N_14299,N_14171);
nor U14732 (N_14732,N_13980,N_14127);
nand U14733 (N_14733,N_13890,N_14301);
and U14734 (N_14734,N_13997,N_13822);
and U14735 (N_14735,N_14070,N_14132);
and U14736 (N_14736,N_13876,N_14110);
and U14737 (N_14737,N_14144,N_14035);
and U14738 (N_14738,N_14099,N_14176);
nor U14739 (N_14739,N_14359,N_14347);
nand U14740 (N_14740,N_14130,N_13949);
and U14741 (N_14741,N_14395,N_14223);
nand U14742 (N_14742,N_14384,N_13947);
or U14743 (N_14743,N_14399,N_14130);
xnor U14744 (N_14744,N_14175,N_13978);
xnor U14745 (N_14745,N_13992,N_13894);
or U14746 (N_14746,N_14151,N_14328);
nand U14747 (N_14747,N_13957,N_14066);
or U14748 (N_14748,N_14281,N_14321);
or U14749 (N_14749,N_13880,N_14106);
xnor U14750 (N_14750,N_14241,N_14362);
or U14751 (N_14751,N_13833,N_14032);
nor U14752 (N_14752,N_14300,N_13862);
nand U14753 (N_14753,N_14239,N_13902);
and U14754 (N_14754,N_14095,N_14105);
and U14755 (N_14755,N_13848,N_13993);
or U14756 (N_14756,N_13987,N_14172);
nand U14757 (N_14757,N_13905,N_14282);
nand U14758 (N_14758,N_14030,N_14217);
and U14759 (N_14759,N_14308,N_14129);
and U14760 (N_14760,N_14138,N_14194);
nor U14761 (N_14761,N_14120,N_14212);
nand U14762 (N_14762,N_14042,N_14351);
and U14763 (N_14763,N_13916,N_14101);
nor U14764 (N_14764,N_14223,N_13975);
nand U14765 (N_14765,N_14361,N_14283);
xor U14766 (N_14766,N_14281,N_14170);
nand U14767 (N_14767,N_13923,N_14102);
nor U14768 (N_14768,N_14193,N_14009);
nor U14769 (N_14769,N_13915,N_14387);
nand U14770 (N_14770,N_13976,N_14146);
or U14771 (N_14771,N_13887,N_14158);
or U14772 (N_14772,N_13966,N_14256);
or U14773 (N_14773,N_13863,N_13884);
nor U14774 (N_14774,N_14250,N_14358);
and U14775 (N_14775,N_14071,N_14304);
nor U14776 (N_14776,N_14077,N_14030);
nand U14777 (N_14777,N_14113,N_14099);
or U14778 (N_14778,N_14333,N_14108);
or U14779 (N_14779,N_14127,N_14372);
nand U14780 (N_14780,N_13956,N_14374);
and U14781 (N_14781,N_14117,N_14036);
or U14782 (N_14782,N_14297,N_14278);
nand U14783 (N_14783,N_14010,N_14121);
nor U14784 (N_14784,N_14320,N_14014);
nand U14785 (N_14785,N_13817,N_13809);
nor U14786 (N_14786,N_13858,N_14173);
nand U14787 (N_14787,N_14195,N_14264);
and U14788 (N_14788,N_14263,N_14200);
xor U14789 (N_14789,N_14055,N_13959);
nor U14790 (N_14790,N_13994,N_14323);
nor U14791 (N_14791,N_14167,N_14091);
or U14792 (N_14792,N_14002,N_13829);
xnor U14793 (N_14793,N_14024,N_14348);
nor U14794 (N_14794,N_13963,N_14069);
nor U14795 (N_14795,N_13879,N_13914);
nor U14796 (N_14796,N_14265,N_13928);
or U14797 (N_14797,N_14259,N_14358);
xor U14798 (N_14798,N_13941,N_13828);
nor U14799 (N_14799,N_13865,N_14166);
nor U14800 (N_14800,N_14336,N_14149);
xor U14801 (N_14801,N_14243,N_13893);
and U14802 (N_14802,N_14336,N_14294);
nor U14803 (N_14803,N_14185,N_14187);
nor U14804 (N_14804,N_14100,N_13883);
and U14805 (N_14805,N_14349,N_14088);
nand U14806 (N_14806,N_13901,N_13909);
nand U14807 (N_14807,N_14134,N_14206);
nand U14808 (N_14808,N_13930,N_13987);
and U14809 (N_14809,N_14379,N_14305);
nand U14810 (N_14810,N_13886,N_13995);
nand U14811 (N_14811,N_13926,N_14156);
and U14812 (N_14812,N_14344,N_13989);
and U14813 (N_14813,N_14031,N_14385);
and U14814 (N_14814,N_14012,N_13879);
and U14815 (N_14815,N_13994,N_14271);
and U14816 (N_14816,N_14118,N_14114);
or U14817 (N_14817,N_14267,N_14017);
xor U14818 (N_14818,N_14239,N_13807);
or U14819 (N_14819,N_14120,N_14251);
and U14820 (N_14820,N_13803,N_14034);
nand U14821 (N_14821,N_13800,N_13876);
nand U14822 (N_14822,N_14282,N_13881);
or U14823 (N_14823,N_14045,N_14263);
nor U14824 (N_14824,N_14296,N_14096);
or U14825 (N_14825,N_14194,N_14350);
nand U14826 (N_14826,N_14347,N_13845);
nor U14827 (N_14827,N_14233,N_13842);
nand U14828 (N_14828,N_13831,N_14236);
and U14829 (N_14829,N_14162,N_14136);
nand U14830 (N_14830,N_14022,N_14260);
and U14831 (N_14831,N_13955,N_14032);
or U14832 (N_14832,N_14058,N_14152);
or U14833 (N_14833,N_14360,N_14370);
nand U14834 (N_14834,N_14102,N_14246);
or U14835 (N_14835,N_14128,N_14133);
xnor U14836 (N_14836,N_14190,N_13801);
nand U14837 (N_14837,N_13998,N_14156);
xnor U14838 (N_14838,N_14038,N_13898);
and U14839 (N_14839,N_14332,N_14072);
nand U14840 (N_14840,N_14258,N_13893);
and U14841 (N_14841,N_14209,N_13889);
or U14842 (N_14842,N_13873,N_14207);
and U14843 (N_14843,N_13846,N_13946);
xor U14844 (N_14844,N_13854,N_14193);
nand U14845 (N_14845,N_14238,N_13843);
or U14846 (N_14846,N_14344,N_14300);
xor U14847 (N_14847,N_14073,N_13922);
and U14848 (N_14848,N_14208,N_14053);
nand U14849 (N_14849,N_14243,N_14106);
and U14850 (N_14850,N_14298,N_14372);
and U14851 (N_14851,N_14355,N_14006);
nor U14852 (N_14852,N_14142,N_14389);
and U14853 (N_14853,N_13807,N_14191);
nor U14854 (N_14854,N_14041,N_13976);
or U14855 (N_14855,N_14257,N_13848);
nand U14856 (N_14856,N_14161,N_14128);
and U14857 (N_14857,N_14310,N_13831);
and U14858 (N_14858,N_14118,N_14377);
nand U14859 (N_14859,N_14205,N_14017);
or U14860 (N_14860,N_14031,N_13977);
or U14861 (N_14861,N_14374,N_13985);
nand U14862 (N_14862,N_14377,N_14305);
and U14863 (N_14863,N_14042,N_14003);
and U14864 (N_14864,N_14056,N_14116);
nor U14865 (N_14865,N_14156,N_13875);
nor U14866 (N_14866,N_14330,N_13958);
and U14867 (N_14867,N_14237,N_14327);
and U14868 (N_14868,N_14346,N_14034);
nand U14869 (N_14869,N_14166,N_14134);
and U14870 (N_14870,N_14179,N_13913);
nor U14871 (N_14871,N_14159,N_14110);
nand U14872 (N_14872,N_14060,N_14371);
nor U14873 (N_14873,N_13961,N_14316);
or U14874 (N_14874,N_13919,N_13860);
nor U14875 (N_14875,N_14391,N_14051);
nor U14876 (N_14876,N_13803,N_14113);
or U14877 (N_14877,N_14368,N_14288);
nor U14878 (N_14878,N_14051,N_13933);
or U14879 (N_14879,N_13831,N_13836);
xor U14880 (N_14880,N_14398,N_14012);
nor U14881 (N_14881,N_14355,N_13949);
nand U14882 (N_14882,N_13887,N_13808);
nand U14883 (N_14883,N_14300,N_13883);
nand U14884 (N_14884,N_14192,N_13999);
or U14885 (N_14885,N_13859,N_14024);
xnor U14886 (N_14886,N_14268,N_14029);
nand U14887 (N_14887,N_14388,N_14073);
nand U14888 (N_14888,N_14023,N_14262);
xnor U14889 (N_14889,N_13825,N_14393);
nand U14890 (N_14890,N_14319,N_13974);
and U14891 (N_14891,N_13862,N_13819);
or U14892 (N_14892,N_14105,N_14192);
nand U14893 (N_14893,N_14353,N_13889);
and U14894 (N_14894,N_13904,N_14161);
xnor U14895 (N_14895,N_13832,N_14244);
xor U14896 (N_14896,N_14392,N_14137);
nor U14897 (N_14897,N_13878,N_13939);
xnor U14898 (N_14898,N_13894,N_13914);
or U14899 (N_14899,N_13801,N_14349);
or U14900 (N_14900,N_14077,N_13958);
nor U14901 (N_14901,N_14290,N_13808);
nor U14902 (N_14902,N_13884,N_14126);
nor U14903 (N_14903,N_14317,N_14337);
nor U14904 (N_14904,N_13989,N_13835);
or U14905 (N_14905,N_13880,N_14046);
nand U14906 (N_14906,N_13995,N_13921);
nor U14907 (N_14907,N_13987,N_14085);
and U14908 (N_14908,N_13904,N_14232);
xor U14909 (N_14909,N_14115,N_14153);
nor U14910 (N_14910,N_13910,N_14392);
and U14911 (N_14911,N_14019,N_14237);
or U14912 (N_14912,N_14215,N_13947);
and U14913 (N_14913,N_14043,N_14126);
and U14914 (N_14914,N_14229,N_14213);
and U14915 (N_14915,N_14243,N_14220);
and U14916 (N_14916,N_13956,N_14326);
nor U14917 (N_14917,N_14023,N_14328);
or U14918 (N_14918,N_14052,N_14274);
xor U14919 (N_14919,N_13938,N_13818);
or U14920 (N_14920,N_14260,N_14017);
and U14921 (N_14921,N_14180,N_14356);
nor U14922 (N_14922,N_13941,N_14104);
nand U14923 (N_14923,N_13856,N_14184);
nand U14924 (N_14924,N_13807,N_13915);
nand U14925 (N_14925,N_14155,N_14184);
nor U14926 (N_14926,N_14050,N_14223);
nand U14927 (N_14927,N_14388,N_14354);
nor U14928 (N_14928,N_13897,N_14029);
xnor U14929 (N_14929,N_14054,N_14373);
nand U14930 (N_14930,N_13837,N_14196);
or U14931 (N_14931,N_14399,N_14217);
nor U14932 (N_14932,N_13856,N_14070);
nor U14933 (N_14933,N_14309,N_14002);
or U14934 (N_14934,N_14067,N_14156);
or U14935 (N_14935,N_13802,N_14264);
nor U14936 (N_14936,N_14063,N_14152);
xor U14937 (N_14937,N_14137,N_14110);
or U14938 (N_14938,N_13869,N_14312);
or U14939 (N_14939,N_14250,N_14277);
nor U14940 (N_14940,N_14223,N_13854);
and U14941 (N_14941,N_14139,N_14309);
and U14942 (N_14942,N_13841,N_14378);
nor U14943 (N_14943,N_14000,N_14095);
and U14944 (N_14944,N_14138,N_14131);
nor U14945 (N_14945,N_14132,N_13887);
nand U14946 (N_14946,N_14386,N_14336);
or U14947 (N_14947,N_13841,N_13953);
xor U14948 (N_14948,N_14162,N_14371);
nor U14949 (N_14949,N_14366,N_13954);
nor U14950 (N_14950,N_14311,N_13959);
nand U14951 (N_14951,N_13911,N_14119);
nor U14952 (N_14952,N_14103,N_14150);
nand U14953 (N_14953,N_13950,N_14357);
nor U14954 (N_14954,N_14196,N_13989);
nor U14955 (N_14955,N_13813,N_13830);
nor U14956 (N_14956,N_14367,N_14364);
nand U14957 (N_14957,N_13806,N_14083);
and U14958 (N_14958,N_13891,N_13942);
nor U14959 (N_14959,N_14319,N_14286);
nor U14960 (N_14960,N_14280,N_13802);
and U14961 (N_14961,N_14256,N_14323);
nor U14962 (N_14962,N_13996,N_14166);
nand U14963 (N_14963,N_13855,N_14248);
nor U14964 (N_14964,N_13902,N_14377);
and U14965 (N_14965,N_14299,N_14370);
nor U14966 (N_14966,N_13884,N_14289);
xor U14967 (N_14967,N_13922,N_14002);
nand U14968 (N_14968,N_14080,N_14091);
nor U14969 (N_14969,N_14080,N_14161);
nand U14970 (N_14970,N_14214,N_13968);
or U14971 (N_14971,N_14137,N_14341);
and U14972 (N_14972,N_14349,N_14134);
or U14973 (N_14973,N_14344,N_14377);
and U14974 (N_14974,N_13864,N_14146);
nor U14975 (N_14975,N_14371,N_14106);
or U14976 (N_14976,N_14154,N_14388);
nand U14977 (N_14977,N_13868,N_14035);
nor U14978 (N_14978,N_14042,N_14244);
or U14979 (N_14979,N_14350,N_14354);
nand U14980 (N_14980,N_14291,N_14223);
nand U14981 (N_14981,N_14391,N_14103);
or U14982 (N_14982,N_14135,N_13941);
or U14983 (N_14983,N_13831,N_13916);
and U14984 (N_14984,N_13882,N_13908);
nor U14985 (N_14985,N_14093,N_14377);
nor U14986 (N_14986,N_14172,N_14230);
and U14987 (N_14987,N_13969,N_14092);
or U14988 (N_14988,N_14043,N_13849);
or U14989 (N_14989,N_14338,N_13833);
and U14990 (N_14990,N_14221,N_14284);
nand U14991 (N_14991,N_14250,N_14115);
and U14992 (N_14992,N_14202,N_13818);
or U14993 (N_14993,N_14023,N_14392);
nor U14994 (N_14994,N_13975,N_14362);
and U14995 (N_14995,N_13848,N_13841);
or U14996 (N_14996,N_14160,N_13886);
and U14997 (N_14997,N_13893,N_14156);
or U14998 (N_14998,N_13848,N_14128);
nand U14999 (N_14999,N_14111,N_13804);
or U15000 (N_15000,N_14740,N_14519);
xnor U15001 (N_15001,N_14703,N_14418);
or U15002 (N_15002,N_14761,N_14553);
nor U15003 (N_15003,N_14438,N_14685);
and U15004 (N_15004,N_14829,N_14623);
and U15005 (N_15005,N_14506,N_14694);
and U15006 (N_15006,N_14733,N_14901);
and U15007 (N_15007,N_14680,N_14862);
nand U15008 (N_15008,N_14711,N_14905);
or U15009 (N_15009,N_14824,N_14976);
nand U15010 (N_15010,N_14531,N_14550);
nor U15011 (N_15011,N_14657,N_14948);
nand U15012 (N_15012,N_14422,N_14458);
and U15013 (N_15013,N_14470,N_14594);
nand U15014 (N_15014,N_14975,N_14805);
xor U15015 (N_15015,N_14760,N_14863);
or U15016 (N_15016,N_14649,N_14897);
nand U15017 (N_15017,N_14993,N_14622);
nor U15018 (N_15018,N_14450,N_14719);
or U15019 (N_15019,N_14745,N_14474);
nor U15020 (N_15020,N_14838,N_14919);
and U15021 (N_15021,N_14826,N_14491);
nor U15022 (N_15022,N_14679,N_14638);
and U15023 (N_15023,N_14442,N_14578);
or U15024 (N_15024,N_14624,N_14788);
nor U15025 (N_15025,N_14634,N_14849);
nand U15026 (N_15026,N_14747,N_14645);
or U15027 (N_15027,N_14423,N_14970);
nor U15028 (N_15028,N_14444,N_14575);
or U15029 (N_15029,N_14419,N_14658);
and U15030 (N_15030,N_14887,N_14405);
nand U15031 (N_15031,N_14425,N_14465);
nor U15032 (N_15032,N_14430,N_14771);
or U15033 (N_15033,N_14522,N_14833);
nor U15034 (N_15034,N_14731,N_14414);
and U15035 (N_15035,N_14844,N_14562);
nor U15036 (N_15036,N_14648,N_14811);
and U15037 (N_15037,N_14873,N_14835);
or U15038 (N_15038,N_14525,N_14670);
and U15039 (N_15039,N_14803,N_14915);
nand U15040 (N_15040,N_14504,N_14674);
nand U15041 (N_15041,N_14582,N_14520);
nor U15042 (N_15042,N_14952,N_14876);
or U15043 (N_15043,N_14896,N_14701);
xor U15044 (N_15044,N_14768,N_14620);
nor U15045 (N_15045,N_14487,N_14951);
or U15046 (N_15046,N_14484,N_14515);
or U15047 (N_15047,N_14945,N_14615);
and U15048 (N_15048,N_14870,N_14936);
xor U15049 (N_15049,N_14696,N_14539);
and U15050 (N_15050,N_14514,N_14435);
xor U15051 (N_15051,N_14930,N_14995);
or U15052 (N_15052,N_14677,N_14523);
and U15053 (N_15053,N_14777,N_14557);
xor U15054 (N_15054,N_14953,N_14804);
xnor U15055 (N_15055,N_14627,N_14505);
or U15056 (N_15056,N_14939,N_14473);
or U15057 (N_15057,N_14791,N_14920);
and U15058 (N_15058,N_14739,N_14810);
or U15059 (N_15059,N_14654,N_14913);
or U15060 (N_15060,N_14601,N_14439);
or U15061 (N_15061,N_14969,N_14540);
or U15062 (N_15062,N_14481,N_14851);
or U15063 (N_15063,N_14538,N_14890);
xnor U15064 (N_15064,N_14786,N_14604);
and U15065 (N_15065,N_14690,N_14571);
xor U15066 (N_15066,N_14613,N_14543);
nand U15067 (N_15067,N_14528,N_14839);
or U15068 (N_15068,N_14879,N_14765);
nand U15069 (N_15069,N_14902,N_14456);
and U15070 (N_15070,N_14569,N_14452);
nand U15071 (N_15071,N_14883,N_14713);
and U15072 (N_15072,N_14854,N_14734);
or U15073 (N_15073,N_14618,N_14885);
xnor U15074 (N_15074,N_14709,N_14981);
or U15075 (N_15075,N_14784,N_14941);
xor U15076 (N_15076,N_14478,N_14437);
and U15077 (N_15077,N_14996,N_14746);
nand U15078 (N_15078,N_14526,N_14860);
xnor U15079 (N_15079,N_14950,N_14779);
or U15080 (N_15080,N_14708,N_14977);
or U15081 (N_15081,N_14721,N_14560);
nand U15082 (N_15082,N_14949,N_14958);
nand U15083 (N_15083,N_14683,N_14602);
nand U15084 (N_15084,N_14954,N_14912);
or U15085 (N_15085,N_14928,N_14937);
or U15086 (N_15086,N_14567,N_14831);
and U15087 (N_15087,N_14732,N_14451);
nor U15088 (N_15088,N_14472,N_14587);
nand U15089 (N_15089,N_14518,N_14922);
xor U15090 (N_15090,N_14960,N_14573);
xor U15091 (N_15091,N_14637,N_14798);
nor U15092 (N_15092,N_14426,N_14632);
and U15093 (N_15093,N_14606,N_14722);
and U15094 (N_15094,N_14743,N_14628);
nand U15095 (N_15095,N_14884,N_14635);
nand U15096 (N_15096,N_14755,N_14455);
nor U15097 (N_15097,N_14845,N_14462);
and U15098 (N_15098,N_14855,N_14880);
nand U15099 (N_15099,N_14821,N_14819);
nand U15100 (N_15100,N_14625,N_14687);
and U15101 (N_15101,N_14772,N_14454);
nand U15102 (N_15102,N_14940,N_14621);
nand U15103 (N_15103,N_14681,N_14642);
xnor U15104 (N_15104,N_14770,N_14999);
nor U15105 (N_15105,N_14978,N_14583);
nor U15106 (N_15106,N_14866,N_14617);
nand U15107 (N_15107,N_14433,N_14527);
or U15108 (N_15108,N_14673,N_14983);
and U15109 (N_15109,N_14700,N_14555);
or U15110 (N_15110,N_14875,N_14877);
nor U15111 (N_15111,N_14840,N_14512);
nor U15112 (N_15112,N_14443,N_14544);
and U15113 (N_15113,N_14900,N_14510);
or U15114 (N_15114,N_14407,N_14497);
nor U15115 (N_15115,N_14809,N_14918);
nand U15116 (N_15116,N_14967,N_14495);
xnor U15117 (N_15117,N_14516,N_14479);
nand U15118 (N_15118,N_14492,N_14769);
or U15119 (N_15119,N_14774,N_14758);
and U15120 (N_15120,N_14785,N_14614);
or U15121 (N_15121,N_14593,N_14716);
nand U15122 (N_15122,N_14572,N_14947);
nor U15123 (N_15123,N_14532,N_14684);
nor U15124 (N_15124,N_14661,N_14790);
and U15125 (N_15125,N_14644,N_14720);
nor U15126 (N_15126,N_14998,N_14545);
or U15127 (N_15127,N_14957,N_14712);
xnor U15128 (N_15128,N_14869,N_14580);
nor U15129 (N_15129,N_14942,N_14974);
nand U15130 (N_15130,N_14453,N_14501);
nand U15131 (N_15131,N_14546,N_14994);
or U15132 (N_15132,N_14726,N_14865);
or U15133 (N_15133,N_14564,N_14850);
nor U15134 (N_15134,N_14989,N_14581);
nand U15135 (N_15135,N_14608,N_14689);
or U15136 (N_15136,N_14893,N_14554);
and U15137 (N_15137,N_14697,N_14535);
nor U15138 (N_15138,N_14923,N_14671);
or U15139 (N_15139,N_14585,N_14801);
xnor U15140 (N_15140,N_14598,N_14600);
nor U15141 (N_15141,N_14933,N_14749);
nand U15142 (N_15142,N_14416,N_14944);
nand U15143 (N_15143,N_14982,N_14822);
nand U15144 (N_15144,N_14886,N_14530);
nand U15145 (N_15145,N_14447,N_14836);
and U15146 (N_15146,N_14847,N_14643);
and U15147 (N_15147,N_14792,N_14925);
or U15148 (N_15148,N_14921,N_14843);
or U15149 (N_15149,N_14841,N_14888);
nor U15150 (N_15150,N_14931,N_14924);
and U15151 (N_15151,N_14903,N_14759);
xor U15152 (N_15152,N_14744,N_14698);
or U15153 (N_15153,N_14415,N_14793);
and U15154 (N_15154,N_14894,N_14757);
nand U15155 (N_15155,N_14971,N_14984);
nor U15156 (N_15156,N_14986,N_14664);
nand U15157 (N_15157,N_14589,N_14429);
nand U15158 (N_15158,N_14424,N_14448);
and U15159 (N_15159,N_14513,N_14874);
nor U15160 (N_15160,N_14653,N_14646);
or U15161 (N_15161,N_14494,N_14586);
xnor U15162 (N_15162,N_14660,N_14872);
and U15163 (N_15163,N_14579,N_14599);
and U15164 (N_15164,N_14682,N_14825);
xor U15165 (N_15165,N_14402,N_14783);
nand U15166 (N_15166,N_14727,N_14688);
or U15167 (N_15167,N_14475,N_14917);
nor U15168 (N_15168,N_14964,N_14480);
or U15169 (N_15169,N_14702,N_14551);
nand U15170 (N_15170,N_14834,N_14899);
nand U15171 (N_15171,N_14817,N_14807);
nand U15172 (N_15172,N_14409,N_14882);
and U15173 (N_15173,N_14493,N_14904);
or U15174 (N_15174,N_14431,N_14440);
and U15175 (N_15175,N_14867,N_14881);
and U15176 (N_15176,N_14932,N_14536);
and U15177 (N_15177,N_14828,N_14837);
nand U15178 (N_15178,N_14542,N_14962);
xnor U15179 (N_15179,N_14421,N_14762);
xnor U15180 (N_15180,N_14662,N_14655);
and U15181 (N_15181,N_14725,N_14449);
nand U15182 (N_15182,N_14509,N_14728);
and U15183 (N_15183,N_14729,N_14754);
and U15184 (N_15184,N_14789,N_14695);
and U15185 (N_15185,N_14891,N_14895);
nor U15186 (N_15186,N_14413,N_14676);
and U15187 (N_15187,N_14730,N_14548);
nand U15188 (N_15188,N_14780,N_14574);
nor U15189 (N_15189,N_14750,N_14609);
nand U15190 (N_15190,N_14503,N_14588);
nand U15191 (N_15191,N_14549,N_14476);
nand U15192 (N_15192,N_14864,N_14767);
nand U15193 (N_15193,N_14558,N_14724);
and U15194 (N_15194,N_14878,N_14929);
nor U15195 (N_15195,N_14537,N_14778);
nand U15196 (N_15196,N_14665,N_14868);
or U15197 (N_15197,N_14796,N_14675);
or U15198 (N_15198,N_14486,N_14692);
nor U15199 (N_15199,N_14595,N_14955);
nor U15200 (N_15200,N_14764,N_14766);
nand U15201 (N_15201,N_14699,N_14577);
nand U15202 (N_15202,N_14799,N_14763);
nor U15203 (N_15203,N_14910,N_14842);
and U15204 (N_15204,N_14496,N_14616);
or U15205 (N_15205,N_14927,N_14943);
xnor U15206 (N_15206,N_14631,N_14808);
and U15207 (N_15207,N_14596,N_14909);
nand U15208 (N_15208,N_14966,N_14477);
and U15209 (N_15209,N_14467,N_14482);
or U15210 (N_15210,N_14650,N_14723);
nor U15211 (N_15211,N_14830,N_14591);
nand U15212 (N_15212,N_14892,N_14411);
nand U15213 (N_15213,N_14773,N_14502);
xor U15214 (N_15214,N_14605,N_14889);
and U15215 (N_15215,N_14959,N_14916);
and U15216 (N_15216,N_14797,N_14633);
or U15217 (N_15217,N_14570,N_14707);
or U15218 (N_15218,N_14787,N_14816);
or U15219 (N_15219,N_14446,N_14432);
and U15220 (N_15220,N_14907,N_14961);
nand U15221 (N_15221,N_14818,N_14814);
xnor U15222 (N_15222,N_14718,N_14956);
and U15223 (N_15223,N_14704,N_14640);
and U15224 (N_15224,N_14693,N_14483);
nor U15225 (N_15225,N_14935,N_14686);
and U15226 (N_15226,N_14946,N_14584);
or U15227 (N_15227,N_14590,N_14517);
or U15228 (N_15228,N_14485,N_14706);
or U15229 (N_15229,N_14667,N_14511);
nand U15230 (N_15230,N_14906,N_14812);
nor U15231 (N_15231,N_14736,N_14813);
nor U15232 (N_15232,N_14802,N_14815);
nand U15233 (N_15233,N_14781,N_14859);
xnor U15234 (N_15234,N_14406,N_14827);
xor U15235 (N_15235,N_14934,N_14498);
and U15236 (N_15236,N_14499,N_14565);
nor U15237 (N_15237,N_14636,N_14412);
or U15238 (N_15238,N_14508,N_14898);
or U15239 (N_15239,N_14612,N_14669);
nor U15240 (N_15240,N_14459,N_14547);
nand U15241 (N_15241,N_14672,N_14710);
nand U15242 (N_15242,N_14991,N_14576);
or U15243 (N_15243,N_14666,N_14436);
and U15244 (N_15244,N_14489,N_14507);
nand U15245 (N_15245,N_14434,N_14820);
nand U15246 (N_15246,N_14806,N_14639);
and U15247 (N_15247,N_14534,N_14782);
nor U15248 (N_15248,N_14592,N_14795);
nor U15249 (N_15249,N_14529,N_14408);
or U15250 (N_15250,N_14552,N_14979);
nand U15251 (N_15251,N_14404,N_14461);
nor U15252 (N_15252,N_14717,N_14742);
and U15253 (N_15253,N_14705,N_14965);
and U15254 (N_15254,N_14626,N_14541);
and U15255 (N_15255,N_14988,N_14656);
nor U15256 (N_15256,N_14775,N_14561);
and U15257 (N_15257,N_14533,N_14990);
or U15258 (N_15258,N_14500,N_14629);
nand U15259 (N_15259,N_14417,N_14464);
or U15260 (N_15260,N_14619,N_14568);
or U15261 (N_15261,N_14972,N_14748);
nand U15262 (N_15262,N_14460,N_14471);
nor U15263 (N_15263,N_14753,N_14427);
and U15264 (N_15264,N_14715,N_14794);
or U15265 (N_15265,N_14914,N_14857);
nor U15266 (N_15266,N_14973,N_14823);
and U15267 (N_15267,N_14490,N_14992);
nor U15268 (N_15268,N_14651,N_14630);
xor U15269 (N_15269,N_14852,N_14563);
nor U15270 (N_15270,N_14756,N_14997);
xnor U15271 (N_15271,N_14400,N_14469);
nand U15272 (N_15272,N_14611,N_14963);
nor U15273 (N_15273,N_14926,N_14911);
and U15274 (N_15274,N_14980,N_14441);
or U15275 (N_15275,N_14908,N_14985);
xor U15276 (N_15276,N_14652,N_14597);
xor U15277 (N_15277,N_14714,N_14800);
or U15278 (N_15278,N_14556,N_14861);
and U15279 (N_15279,N_14603,N_14776);
or U15280 (N_15280,N_14521,N_14466);
nor U15281 (N_15281,N_14832,N_14403);
and U15282 (N_15282,N_14668,N_14987);
and U15283 (N_15283,N_14610,N_14641);
xnor U15284 (N_15284,N_14737,N_14938);
xor U15285 (N_15285,N_14678,N_14663);
or U15286 (N_15286,N_14468,N_14607);
and U15287 (N_15287,N_14858,N_14752);
and U15288 (N_15288,N_14463,N_14401);
or U15289 (N_15289,N_14457,N_14445);
nand U15290 (N_15290,N_14566,N_14647);
nand U15291 (N_15291,N_14488,N_14410);
nor U15292 (N_15292,N_14848,N_14420);
and U15293 (N_15293,N_14738,N_14559);
or U15294 (N_15294,N_14735,N_14871);
and U15295 (N_15295,N_14853,N_14691);
nor U15296 (N_15296,N_14968,N_14659);
and U15297 (N_15297,N_14524,N_14856);
nor U15298 (N_15298,N_14751,N_14428);
and U15299 (N_15299,N_14741,N_14846);
and U15300 (N_15300,N_14432,N_14722);
or U15301 (N_15301,N_14440,N_14830);
nand U15302 (N_15302,N_14491,N_14415);
or U15303 (N_15303,N_14837,N_14886);
nor U15304 (N_15304,N_14811,N_14557);
and U15305 (N_15305,N_14887,N_14468);
nand U15306 (N_15306,N_14517,N_14946);
or U15307 (N_15307,N_14853,N_14816);
nor U15308 (N_15308,N_14628,N_14724);
nand U15309 (N_15309,N_14813,N_14567);
nor U15310 (N_15310,N_14976,N_14996);
nand U15311 (N_15311,N_14911,N_14751);
xor U15312 (N_15312,N_14467,N_14564);
and U15313 (N_15313,N_14487,N_14676);
or U15314 (N_15314,N_14496,N_14494);
nor U15315 (N_15315,N_14452,N_14830);
or U15316 (N_15316,N_14503,N_14973);
and U15317 (N_15317,N_14818,N_14672);
or U15318 (N_15318,N_14831,N_14650);
or U15319 (N_15319,N_14593,N_14840);
or U15320 (N_15320,N_14543,N_14771);
nor U15321 (N_15321,N_14464,N_14741);
and U15322 (N_15322,N_14636,N_14435);
and U15323 (N_15323,N_14613,N_14900);
xor U15324 (N_15324,N_14957,N_14502);
nand U15325 (N_15325,N_14493,N_14813);
and U15326 (N_15326,N_14933,N_14785);
or U15327 (N_15327,N_14550,N_14413);
or U15328 (N_15328,N_14803,N_14720);
or U15329 (N_15329,N_14666,N_14991);
and U15330 (N_15330,N_14565,N_14505);
and U15331 (N_15331,N_14769,N_14872);
or U15332 (N_15332,N_14823,N_14853);
and U15333 (N_15333,N_14995,N_14950);
nor U15334 (N_15334,N_14784,N_14642);
xor U15335 (N_15335,N_14405,N_14603);
or U15336 (N_15336,N_14798,N_14749);
and U15337 (N_15337,N_14419,N_14529);
nor U15338 (N_15338,N_14528,N_14922);
nand U15339 (N_15339,N_14642,N_14866);
and U15340 (N_15340,N_14939,N_14553);
nor U15341 (N_15341,N_14424,N_14923);
nor U15342 (N_15342,N_14877,N_14478);
or U15343 (N_15343,N_14718,N_14988);
and U15344 (N_15344,N_14406,N_14947);
xnor U15345 (N_15345,N_14500,N_14693);
nor U15346 (N_15346,N_14943,N_14644);
and U15347 (N_15347,N_14946,N_14607);
nor U15348 (N_15348,N_14508,N_14635);
nor U15349 (N_15349,N_14843,N_14638);
or U15350 (N_15350,N_14860,N_14467);
or U15351 (N_15351,N_14411,N_14804);
nand U15352 (N_15352,N_14831,N_14767);
and U15353 (N_15353,N_14666,N_14554);
nor U15354 (N_15354,N_14609,N_14453);
or U15355 (N_15355,N_14799,N_14462);
xnor U15356 (N_15356,N_14443,N_14564);
nand U15357 (N_15357,N_14897,N_14507);
nand U15358 (N_15358,N_14801,N_14573);
or U15359 (N_15359,N_14945,N_14482);
nand U15360 (N_15360,N_14601,N_14504);
or U15361 (N_15361,N_14911,N_14544);
or U15362 (N_15362,N_14744,N_14843);
and U15363 (N_15363,N_14744,N_14481);
nand U15364 (N_15364,N_14906,N_14571);
nand U15365 (N_15365,N_14571,N_14859);
nor U15366 (N_15366,N_14594,N_14729);
or U15367 (N_15367,N_14703,N_14701);
and U15368 (N_15368,N_14916,N_14766);
or U15369 (N_15369,N_14484,N_14977);
nor U15370 (N_15370,N_14642,N_14877);
or U15371 (N_15371,N_14738,N_14494);
or U15372 (N_15372,N_14824,N_14883);
nand U15373 (N_15373,N_14704,N_14478);
or U15374 (N_15374,N_14999,N_14921);
xor U15375 (N_15375,N_14755,N_14691);
nor U15376 (N_15376,N_14468,N_14729);
nor U15377 (N_15377,N_14819,N_14927);
or U15378 (N_15378,N_14617,N_14823);
nand U15379 (N_15379,N_14710,N_14975);
nand U15380 (N_15380,N_14416,N_14722);
and U15381 (N_15381,N_14868,N_14789);
or U15382 (N_15382,N_14493,N_14740);
nor U15383 (N_15383,N_14757,N_14878);
or U15384 (N_15384,N_14467,N_14668);
nor U15385 (N_15385,N_14728,N_14442);
or U15386 (N_15386,N_14752,N_14583);
or U15387 (N_15387,N_14503,N_14713);
nand U15388 (N_15388,N_14502,N_14920);
or U15389 (N_15389,N_14689,N_14899);
xnor U15390 (N_15390,N_14649,N_14890);
nor U15391 (N_15391,N_14622,N_14891);
or U15392 (N_15392,N_14743,N_14988);
and U15393 (N_15393,N_14871,N_14695);
nand U15394 (N_15394,N_14717,N_14451);
and U15395 (N_15395,N_14747,N_14876);
nor U15396 (N_15396,N_14666,N_14810);
and U15397 (N_15397,N_14466,N_14718);
xnor U15398 (N_15398,N_14695,N_14447);
and U15399 (N_15399,N_14703,N_14967);
and U15400 (N_15400,N_14705,N_14759);
and U15401 (N_15401,N_14517,N_14562);
xnor U15402 (N_15402,N_14971,N_14808);
or U15403 (N_15403,N_14921,N_14502);
nand U15404 (N_15404,N_14972,N_14873);
nor U15405 (N_15405,N_14972,N_14937);
nor U15406 (N_15406,N_14440,N_14887);
nor U15407 (N_15407,N_14626,N_14991);
xor U15408 (N_15408,N_14778,N_14858);
xor U15409 (N_15409,N_14537,N_14686);
nor U15410 (N_15410,N_14998,N_14630);
or U15411 (N_15411,N_14645,N_14478);
and U15412 (N_15412,N_14477,N_14880);
nand U15413 (N_15413,N_14945,N_14628);
nand U15414 (N_15414,N_14567,N_14599);
nor U15415 (N_15415,N_14842,N_14816);
xnor U15416 (N_15416,N_14910,N_14719);
xor U15417 (N_15417,N_14632,N_14998);
and U15418 (N_15418,N_14506,N_14671);
or U15419 (N_15419,N_14476,N_14505);
or U15420 (N_15420,N_14810,N_14846);
or U15421 (N_15421,N_14437,N_14920);
nand U15422 (N_15422,N_14780,N_14531);
and U15423 (N_15423,N_14435,N_14704);
nor U15424 (N_15424,N_14811,N_14677);
and U15425 (N_15425,N_14676,N_14898);
nand U15426 (N_15426,N_14428,N_14944);
and U15427 (N_15427,N_14731,N_14743);
nand U15428 (N_15428,N_14916,N_14587);
nand U15429 (N_15429,N_14604,N_14850);
nand U15430 (N_15430,N_14740,N_14850);
nand U15431 (N_15431,N_14528,N_14880);
nand U15432 (N_15432,N_14421,N_14793);
nand U15433 (N_15433,N_14754,N_14826);
xor U15434 (N_15434,N_14509,N_14828);
xnor U15435 (N_15435,N_14537,N_14972);
xor U15436 (N_15436,N_14748,N_14534);
nor U15437 (N_15437,N_14644,N_14554);
nand U15438 (N_15438,N_14413,N_14446);
nand U15439 (N_15439,N_14475,N_14868);
or U15440 (N_15440,N_14871,N_14474);
and U15441 (N_15441,N_14554,N_14885);
nand U15442 (N_15442,N_14974,N_14424);
and U15443 (N_15443,N_14722,N_14548);
nand U15444 (N_15444,N_14475,N_14736);
nand U15445 (N_15445,N_14495,N_14534);
and U15446 (N_15446,N_14456,N_14755);
xor U15447 (N_15447,N_14470,N_14769);
xor U15448 (N_15448,N_14644,N_14608);
or U15449 (N_15449,N_14930,N_14973);
and U15450 (N_15450,N_14483,N_14529);
and U15451 (N_15451,N_14775,N_14908);
nor U15452 (N_15452,N_14445,N_14463);
nor U15453 (N_15453,N_14643,N_14483);
or U15454 (N_15454,N_14625,N_14411);
and U15455 (N_15455,N_14924,N_14856);
or U15456 (N_15456,N_14889,N_14560);
nand U15457 (N_15457,N_14734,N_14651);
nor U15458 (N_15458,N_14837,N_14815);
xnor U15459 (N_15459,N_14928,N_14505);
or U15460 (N_15460,N_14537,N_14756);
nor U15461 (N_15461,N_14899,N_14554);
nand U15462 (N_15462,N_14996,N_14720);
and U15463 (N_15463,N_14441,N_14874);
or U15464 (N_15464,N_14522,N_14997);
nor U15465 (N_15465,N_14640,N_14498);
nand U15466 (N_15466,N_14955,N_14488);
nor U15467 (N_15467,N_14773,N_14609);
or U15468 (N_15468,N_14440,N_14893);
or U15469 (N_15469,N_14407,N_14605);
nor U15470 (N_15470,N_14984,N_14965);
and U15471 (N_15471,N_14809,N_14425);
and U15472 (N_15472,N_14935,N_14687);
nor U15473 (N_15473,N_14954,N_14680);
or U15474 (N_15474,N_14857,N_14717);
nor U15475 (N_15475,N_14400,N_14733);
and U15476 (N_15476,N_14675,N_14893);
and U15477 (N_15477,N_14825,N_14655);
and U15478 (N_15478,N_14509,N_14493);
or U15479 (N_15479,N_14551,N_14904);
or U15480 (N_15480,N_14679,N_14595);
xnor U15481 (N_15481,N_14751,N_14464);
nand U15482 (N_15482,N_14915,N_14482);
nand U15483 (N_15483,N_14809,N_14862);
and U15484 (N_15484,N_14419,N_14631);
or U15485 (N_15485,N_14516,N_14689);
nor U15486 (N_15486,N_14700,N_14493);
or U15487 (N_15487,N_14489,N_14699);
nor U15488 (N_15488,N_14552,N_14417);
nand U15489 (N_15489,N_14646,N_14830);
nand U15490 (N_15490,N_14922,N_14761);
or U15491 (N_15491,N_14970,N_14538);
and U15492 (N_15492,N_14669,N_14979);
nor U15493 (N_15493,N_14838,N_14485);
nor U15494 (N_15494,N_14965,N_14661);
nand U15495 (N_15495,N_14941,N_14585);
nor U15496 (N_15496,N_14939,N_14886);
nor U15497 (N_15497,N_14974,N_14903);
nand U15498 (N_15498,N_14921,N_14428);
nor U15499 (N_15499,N_14960,N_14962);
and U15500 (N_15500,N_14729,N_14687);
nor U15501 (N_15501,N_14513,N_14599);
and U15502 (N_15502,N_14765,N_14825);
or U15503 (N_15503,N_14964,N_14582);
nand U15504 (N_15504,N_14419,N_14951);
nand U15505 (N_15505,N_14539,N_14742);
nor U15506 (N_15506,N_14949,N_14732);
or U15507 (N_15507,N_14901,N_14852);
xnor U15508 (N_15508,N_14729,N_14565);
nand U15509 (N_15509,N_14782,N_14641);
or U15510 (N_15510,N_14806,N_14461);
xor U15511 (N_15511,N_14634,N_14917);
nand U15512 (N_15512,N_14970,N_14447);
nor U15513 (N_15513,N_14429,N_14962);
nor U15514 (N_15514,N_14719,N_14714);
nand U15515 (N_15515,N_14899,N_14946);
xnor U15516 (N_15516,N_14406,N_14763);
nand U15517 (N_15517,N_14451,N_14968);
nor U15518 (N_15518,N_14714,N_14827);
and U15519 (N_15519,N_14723,N_14412);
or U15520 (N_15520,N_14791,N_14658);
or U15521 (N_15521,N_14884,N_14978);
or U15522 (N_15522,N_14746,N_14509);
or U15523 (N_15523,N_14633,N_14755);
nand U15524 (N_15524,N_14757,N_14407);
or U15525 (N_15525,N_14435,N_14540);
nor U15526 (N_15526,N_14975,N_14733);
or U15527 (N_15527,N_14723,N_14875);
xnor U15528 (N_15528,N_14810,N_14414);
or U15529 (N_15529,N_14458,N_14661);
and U15530 (N_15530,N_14568,N_14888);
and U15531 (N_15531,N_14850,N_14877);
xnor U15532 (N_15532,N_14749,N_14605);
nand U15533 (N_15533,N_14905,N_14633);
and U15534 (N_15534,N_14562,N_14634);
nor U15535 (N_15535,N_14755,N_14641);
or U15536 (N_15536,N_14539,N_14907);
nand U15537 (N_15537,N_14827,N_14470);
or U15538 (N_15538,N_14408,N_14737);
and U15539 (N_15539,N_14948,N_14627);
nor U15540 (N_15540,N_14916,N_14606);
nor U15541 (N_15541,N_14488,N_14625);
and U15542 (N_15542,N_14803,N_14499);
or U15543 (N_15543,N_14593,N_14872);
and U15544 (N_15544,N_14480,N_14551);
nand U15545 (N_15545,N_14828,N_14489);
xor U15546 (N_15546,N_14725,N_14882);
nor U15547 (N_15547,N_14808,N_14950);
nand U15548 (N_15548,N_14983,N_14497);
and U15549 (N_15549,N_14778,N_14879);
nor U15550 (N_15550,N_14771,N_14741);
nor U15551 (N_15551,N_14413,N_14574);
and U15552 (N_15552,N_14951,N_14779);
or U15553 (N_15553,N_14453,N_14646);
nor U15554 (N_15554,N_14988,N_14648);
and U15555 (N_15555,N_14931,N_14714);
and U15556 (N_15556,N_14958,N_14699);
nor U15557 (N_15557,N_14874,N_14861);
and U15558 (N_15558,N_14610,N_14591);
and U15559 (N_15559,N_14692,N_14673);
nor U15560 (N_15560,N_14924,N_14730);
xor U15561 (N_15561,N_14925,N_14549);
and U15562 (N_15562,N_14862,N_14670);
nor U15563 (N_15563,N_14692,N_14813);
and U15564 (N_15564,N_14548,N_14798);
nand U15565 (N_15565,N_14668,N_14604);
xnor U15566 (N_15566,N_14638,N_14501);
and U15567 (N_15567,N_14961,N_14905);
nand U15568 (N_15568,N_14419,N_14651);
or U15569 (N_15569,N_14893,N_14895);
nor U15570 (N_15570,N_14821,N_14893);
xnor U15571 (N_15571,N_14967,N_14913);
and U15572 (N_15572,N_14497,N_14802);
nor U15573 (N_15573,N_14524,N_14504);
nand U15574 (N_15574,N_14882,N_14608);
and U15575 (N_15575,N_14814,N_14548);
and U15576 (N_15576,N_14819,N_14917);
and U15577 (N_15577,N_14590,N_14439);
and U15578 (N_15578,N_14541,N_14550);
or U15579 (N_15579,N_14710,N_14729);
nor U15580 (N_15580,N_14958,N_14889);
and U15581 (N_15581,N_14918,N_14989);
or U15582 (N_15582,N_14443,N_14956);
and U15583 (N_15583,N_14820,N_14887);
xor U15584 (N_15584,N_14642,N_14492);
nand U15585 (N_15585,N_14724,N_14772);
xnor U15586 (N_15586,N_14807,N_14618);
nand U15587 (N_15587,N_14694,N_14411);
xnor U15588 (N_15588,N_14777,N_14783);
nor U15589 (N_15589,N_14598,N_14920);
nor U15590 (N_15590,N_14519,N_14717);
nand U15591 (N_15591,N_14518,N_14806);
nor U15592 (N_15592,N_14540,N_14699);
nand U15593 (N_15593,N_14724,N_14840);
or U15594 (N_15594,N_14938,N_14569);
xnor U15595 (N_15595,N_14745,N_14824);
nor U15596 (N_15596,N_14634,N_14598);
or U15597 (N_15597,N_14539,N_14702);
and U15598 (N_15598,N_14998,N_14898);
and U15599 (N_15599,N_14411,N_14540);
nand U15600 (N_15600,N_15066,N_15555);
nand U15601 (N_15601,N_15593,N_15298);
or U15602 (N_15602,N_15320,N_15273);
and U15603 (N_15603,N_15245,N_15220);
or U15604 (N_15604,N_15553,N_15057);
nor U15605 (N_15605,N_15041,N_15590);
nand U15606 (N_15606,N_15424,N_15284);
nor U15607 (N_15607,N_15122,N_15489);
nor U15608 (N_15608,N_15543,N_15014);
nand U15609 (N_15609,N_15049,N_15221);
nand U15610 (N_15610,N_15161,N_15462);
nor U15611 (N_15611,N_15060,N_15180);
nor U15612 (N_15612,N_15587,N_15370);
or U15613 (N_15613,N_15451,N_15585);
nor U15614 (N_15614,N_15427,N_15281);
xnor U15615 (N_15615,N_15234,N_15296);
or U15616 (N_15616,N_15052,N_15080);
and U15617 (N_15617,N_15567,N_15056);
nor U15618 (N_15618,N_15279,N_15238);
or U15619 (N_15619,N_15414,N_15045);
and U15620 (N_15620,N_15196,N_15438);
xnor U15621 (N_15621,N_15417,N_15382);
and U15622 (N_15622,N_15218,N_15127);
or U15623 (N_15623,N_15235,N_15465);
and U15624 (N_15624,N_15561,N_15401);
or U15625 (N_15625,N_15065,N_15541);
or U15626 (N_15626,N_15252,N_15483);
nor U15627 (N_15627,N_15446,N_15338);
xor U15628 (N_15628,N_15450,N_15395);
xnor U15629 (N_15629,N_15242,N_15477);
or U15630 (N_15630,N_15393,N_15399);
xor U15631 (N_15631,N_15062,N_15449);
nand U15632 (N_15632,N_15016,N_15211);
nor U15633 (N_15633,N_15519,N_15368);
nor U15634 (N_15634,N_15171,N_15227);
and U15635 (N_15635,N_15311,N_15157);
nor U15636 (N_15636,N_15346,N_15082);
nor U15637 (N_15637,N_15149,N_15093);
and U15638 (N_15638,N_15113,N_15352);
or U15639 (N_15639,N_15473,N_15594);
or U15640 (N_15640,N_15170,N_15323);
or U15641 (N_15641,N_15566,N_15403);
and U15642 (N_15642,N_15570,N_15186);
and U15643 (N_15643,N_15430,N_15431);
nor U15644 (N_15644,N_15268,N_15255);
nor U15645 (N_15645,N_15231,N_15042);
and U15646 (N_15646,N_15520,N_15367);
xnor U15647 (N_15647,N_15074,N_15288);
xor U15648 (N_15648,N_15069,N_15456);
and U15649 (N_15649,N_15175,N_15249);
nand U15650 (N_15650,N_15105,N_15257);
or U15651 (N_15651,N_15592,N_15190);
nand U15652 (N_15652,N_15025,N_15397);
nand U15653 (N_15653,N_15205,N_15275);
and U15654 (N_15654,N_15110,N_15260);
nand U15655 (N_15655,N_15130,N_15419);
nor U15656 (N_15656,N_15484,N_15474);
or U15657 (N_15657,N_15054,N_15534);
nand U15658 (N_15658,N_15576,N_15286);
xnor U15659 (N_15659,N_15387,N_15330);
or U15660 (N_15660,N_15011,N_15126);
nor U15661 (N_15661,N_15578,N_15121);
nand U15662 (N_15662,N_15266,N_15361);
or U15663 (N_15663,N_15481,N_15136);
or U15664 (N_15664,N_15202,N_15568);
nand U15665 (N_15665,N_15537,N_15280);
and U15666 (N_15666,N_15219,N_15172);
and U15667 (N_15667,N_15479,N_15125);
nor U15668 (N_15668,N_15415,N_15454);
and U15669 (N_15669,N_15564,N_15455);
nand U15670 (N_15670,N_15572,N_15335);
or U15671 (N_15671,N_15591,N_15264);
or U15672 (N_15672,N_15114,N_15597);
nand U15673 (N_15673,N_15144,N_15307);
nor U15674 (N_15674,N_15106,N_15493);
and U15675 (N_15675,N_15523,N_15466);
xnor U15676 (N_15676,N_15013,N_15326);
nor U15677 (N_15677,N_15141,N_15118);
or U15678 (N_15678,N_15504,N_15117);
or U15679 (N_15679,N_15253,N_15324);
nor U15680 (N_15680,N_15058,N_15254);
nand U15681 (N_15681,N_15596,N_15471);
nor U15682 (N_15682,N_15285,N_15292);
or U15683 (N_15683,N_15535,N_15169);
nor U15684 (N_15684,N_15001,N_15295);
xnor U15685 (N_15685,N_15162,N_15073);
xnor U15686 (N_15686,N_15050,N_15499);
nor U15687 (N_15687,N_15072,N_15502);
nand U15688 (N_15688,N_15077,N_15487);
and U15689 (N_15689,N_15148,N_15023);
or U15690 (N_15690,N_15312,N_15478);
or U15691 (N_15691,N_15391,N_15491);
or U15692 (N_15692,N_15012,N_15232);
or U15693 (N_15693,N_15021,N_15457);
or U15694 (N_15694,N_15354,N_15133);
or U15695 (N_15695,N_15189,N_15433);
and U15696 (N_15696,N_15165,N_15303);
xor U15697 (N_15697,N_15034,N_15434);
or U15698 (N_15698,N_15159,N_15138);
and U15699 (N_15699,N_15182,N_15586);
nor U15700 (N_15700,N_15293,N_15263);
and U15701 (N_15701,N_15097,N_15026);
and U15702 (N_15702,N_15297,N_15174);
nand U15703 (N_15703,N_15579,N_15142);
or U15704 (N_15704,N_15055,N_15557);
or U15705 (N_15705,N_15542,N_15380);
nand U15706 (N_15706,N_15256,N_15194);
nand U15707 (N_15707,N_15460,N_15091);
or U15708 (N_15708,N_15267,N_15360);
or U15709 (N_15709,N_15135,N_15463);
nand U15710 (N_15710,N_15507,N_15467);
or U15711 (N_15711,N_15505,N_15191);
or U15712 (N_15712,N_15095,N_15390);
nand U15713 (N_15713,N_15398,N_15005);
nand U15714 (N_15714,N_15129,N_15316);
and U15715 (N_15715,N_15468,N_15143);
or U15716 (N_15716,N_15480,N_15540);
and U15717 (N_15717,N_15098,N_15506);
nor U15718 (N_15718,N_15299,N_15007);
and U15719 (N_15719,N_15582,N_15377);
nor U15720 (N_15720,N_15134,N_15269);
or U15721 (N_15721,N_15246,N_15146);
or U15722 (N_15722,N_15495,N_15321);
xnor U15723 (N_15723,N_15508,N_15119);
xnor U15724 (N_15724,N_15469,N_15533);
xnor U15725 (N_15725,N_15396,N_15558);
and U15726 (N_15726,N_15379,N_15029);
nor U15727 (N_15727,N_15214,N_15075);
nand U15728 (N_15728,N_15006,N_15552);
or U15729 (N_15729,N_15109,N_15063);
nand U15730 (N_15730,N_15038,N_15203);
nor U15731 (N_15731,N_15306,N_15490);
nand U15732 (N_15732,N_15375,N_15559);
or U15733 (N_15733,N_15244,N_15532);
or U15734 (N_15734,N_15128,N_15332);
and U15735 (N_15735,N_15429,N_15027);
or U15736 (N_15736,N_15373,N_15197);
nor U15737 (N_15737,N_15522,N_15201);
and U15738 (N_15738,N_15047,N_15158);
xnor U15739 (N_15739,N_15341,N_15061);
and U15740 (N_15740,N_15327,N_15283);
nor U15741 (N_15741,N_15239,N_15363);
nor U15742 (N_15742,N_15309,N_15453);
and U15743 (N_15743,N_15008,N_15563);
nor U15744 (N_15744,N_15193,N_15147);
and U15745 (N_15745,N_15388,N_15413);
and U15746 (N_15746,N_15371,N_15376);
and U15747 (N_15747,N_15319,N_15177);
and U15748 (N_15748,N_15215,N_15521);
or U15749 (N_15749,N_15529,N_15096);
nor U15750 (N_15750,N_15035,N_15347);
xor U15751 (N_15751,N_15536,N_15271);
nand U15752 (N_15752,N_15584,N_15575);
xnor U15753 (N_15753,N_15085,N_15369);
nor U15754 (N_15754,N_15140,N_15204);
nand U15755 (N_15755,N_15084,N_15120);
nand U15756 (N_15756,N_15435,N_15086);
nor U15757 (N_15757,N_15528,N_15313);
and U15758 (N_15758,N_15359,N_15131);
xnor U15759 (N_15759,N_15067,N_15348);
nor U15760 (N_15760,N_15087,N_15545);
or U15761 (N_15761,N_15043,N_15544);
xnor U15762 (N_15762,N_15032,N_15099);
or U15763 (N_15763,N_15046,N_15274);
and U15764 (N_15764,N_15112,N_15291);
nand U15765 (N_15765,N_15198,N_15525);
or U15766 (N_15766,N_15019,N_15531);
nor U15767 (N_15767,N_15418,N_15524);
xor U15768 (N_15768,N_15224,N_15294);
or U15769 (N_15769,N_15183,N_15207);
nor U15770 (N_15770,N_15222,N_15331);
and U15771 (N_15771,N_15514,N_15164);
xnor U15772 (N_15772,N_15248,N_15437);
xor U15773 (N_15773,N_15223,N_15325);
nor U15774 (N_15774,N_15031,N_15150);
nand U15775 (N_15775,N_15365,N_15384);
and U15776 (N_15776,N_15447,N_15459);
nor U15777 (N_15777,N_15314,N_15394);
nor U15778 (N_15778,N_15233,N_15503);
or U15779 (N_15779,N_15343,N_15378);
nor U15780 (N_15780,N_15448,N_15372);
nor U15781 (N_15781,N_15560,N_15250);
nor U15782 (N_15782,N_15265,N_15036);
or U15783 (N_15783,N_15059,N_15156);
nor U15784 (N_15784,N_15276,N_15440);
nand U15785 (N_15785,N_15512,N_15290);
or U15786 (N_15786,N_15188,N_15152);
and U15787 (N_15787,N_15168,N_15580);
or U15788 (N_15788,N_15339,N_15226);
and U15789 (N_15789,N_15199,N_15470);
or U15790 (N_15790,N_15179,N_15442);
xor U15791 (N_15791,N_15488,N_15565);
nor U15792 (N_15792,N_15002,N_15079);
xnor U15793 (N_15793,N_15089,N_15108);
nor U15794 (N_15794,N_15076,N_15476);
or U15795 (N_15795,N_15184,N_15259);
nand U15796 (N_15796,N_15443,N_15538);
and U15797 (N_15797,N_15322,N_15102);
xor U15798 (N_15798,N_15349,N_15334);
nor U15799 (N_15799,N_15464,N_15210);
nor U15800 (N_15800,N_15185,N_15022);
or U15801 (N_15801,N_15145,N_15546);
nand U15802 (N_15802,N_15406,N_15425);
nand U15803 (N_15803,N_15216,N_15333);
xnor U15804 (N_15804,N_15385,N_15598);
nand U15805 (N_15805,N_15383,N_15556);
nand U15806 (N_15806,N_15444,N_15494);
nand U15807 (N_15807,N_15208,N_15048);
nor U15808 (N_15808,N_15195,N_15004);
and U15809 (N_15809,N_15236,N_15404);
or U15810 (N_15810,N_15258,N_15501);
nand U15811 (N_15811,N_15017,N_15412);
and U15812 (N_15812,N_15081,N_15588);
xor U15813 (N_15813,N_15277,N_15517);
nand U15814 (N_15814,N_15229,N_15083);
nor U15815 (N_15815,N_15569,N_15426);
nor U15816 (N_15816,N_15577,N_15270);
nor U15817 (N_15817,N_15305,N_15599);
or U15818 (N_15818,N_15100,N_15356);
and U15819 (N_15819,N_15304,N_15030);
nor U15820 (N_15820,N_15410,N_15228);
and U15821 (N_15821,N_15044,N_15358);
nor U15822 (N_15822,N_15439,N_15436);
and U15823 (N_15823,N_15340,N_15581);
or U15824 (N_15824,N_15513,N_15511);
nand U15825 (N_15825,N_15241,N_15486);
nand U15826 (N_15826,N_15237,N_15589);
nor U15827 (N_15827,N_15153,N_15166);
or U15828 (N_15828,N_15261,N_15010);
or U15829 (N_15829,N_15282,N_15040);
nor U15830 (N_15830,N_15139,N_15287);
nand U15831 (N_15831,N_15498,N_15516);
or U15832 (N_15832,N_15111,N_15357);
nor U15833 (N_15833,N_15344,N_15416);
or U15834 (N_15834,N_15116,N_15289);
or U15835 (N_15835,N_15432,N_15317);
or U15836 (N_15836,N_15018,N_15173);
nand U15837 (N_15837,N_15247,N_15115);
and U15838 (N_15838,N_15003,N_15230);
or U15839 (N_15839,N_15315,N_15064);
or U15840 (N_15840,N_15217,N_15518);
or U15841 (N_15841,N_15137,N_15068);
xor U15842 (N_15842,N_15548,N_15104);
and U15843 (N_15843,N_15527,N_15485);
nor U15844 (N_15844,N_15020,N_15039);
nor U15845 (N_15845,N_15381,N_15408);
and U15846 (N_15846,N_15472,N_15213);
nand U15847 (N_15847,N_15300,N_15251);
or U15848 (N_15848,N_15402,N_15051);
or U15849 (N_15849,N_15337,N_15526);
nor U15850 (N_15850,N_15178,N_15103);
nor U15851 (N_15851,N_15530,N_15094);
or U15852 (N_15852,N_15272,N_15240);
or U15853 (N_15853,N_15124,N_15132);
and U15854 (N_15854,N_15310,N_15458);
or U15855 (N_15855,N_15510,N_15024);
and U15856 (N_15856,N_15151,N_15088);
nand U15857 (N_15857,N_15009,N_15409);
and U15858 (N_15858,N_15421,N_15350);
xor U15859 (N_15859,N_15411,N_15386);
nand U15860 (N_15860,N_15345,N_15187);
nor U15861 (N_15861,N_15496,N_15033);
and U15862 (N_15862,N_15200,N_15209);
nor U15863 (N_15863,N_15037,N_15176);
nor U15864 (N_15864,N_15028,N_15243);
nand U15865 (N_15865,N_15342,N_15452);
xor U15866 (N_15866,N_15329,N_15492);
and U15867 (N_15867,N_15583,N_15071);
nand U15868 (N_15868,N_15154,N_15571);
or U15869 (N_15869,N_15192,N_15461);
nor U15870 (N_15870,N_15475,N_15423);
nor U15871 (N_15871,N_15181,N_15550);
or U15872 (N_15872,N_15509,N_15573);
nand U15873 (N_15873,N_15405,N_15155);
or U15874 (N_15874,N_15053,N_15015);
and U15875 (N_15875,N_15482,N_15262);
nand U15876 (N_15876,N_15539,N_15078);
nor U15877 (N_15877,N_15422,N_15500);
xnor U15878 (N_15878,N_15355,N_15364);
xnor U15879 (N_15879,N_15107,N_15389);
or U15880 (N_15880,N_15308,N_15318);
and U15881 (N_15881,N_15206,N_15090);
or U15882 (N_15882,N_15595,N_15302);
and U15883 (N_15883,N_15441,N_15167);
and U15884 (N_15884,N_15362,N_15160);
or U15885 (N_15885,N_15101,N_15562);
and U15886 (N_15886,N_15551,N_15353);
xnor U15887 (N_15887,N_15547,N_15225);
nor U15888 (N_15888,N_15497,N_15070);
and U15889 (N_15889,N_15163,N_15123);
and U15890 (N_15890,N_15092,N_15328);
xnor U15891 (N_15891,N_15336,N_15428);
xor U15892 (N_15892,N_15407,N_15366);
nand U15893 (N_15893,N_15420,N_15278);
or U15894 (N_15894,N_15392,N_15515);
nor U15895 (N_15895,N_15574,N_15549);
nor U15896 (N_15896,N_15554,N_15212);
and U15897 (N_15897,N_15351,N_15445);
or U15898 (N_15898,N_15374,N_15400);
nand U15899 (N_15899,N_15000,N_15301);
or U15900 (N_15900,N_15098,N_15012);
nand U15901 (N_15901,N_15162,N_15197);
and U15902 (N_15902,N_15458,N_15361);
and U15903 (N_15903,N_15185,N_15309);
or U15904 (N_15904,N_15180,N_15554);
or U15905 (N_15905,N_15340,N_15561);
nor U15906 (N_15906,N_15576,N_15417);
and U15907 (N_15907,N_15012,N_15471);
nand U15908 (N_15908,N_15147,N_15549);
nand U15909 (N_15909,N_15554,N_15351);
nor U15910 (N_15910,N_15380,N_15120);
nand U15911 (N_15911,N_15503,N_15557);
and U15912 (N_15912,N_15352,N_15594);
and U15913 (N_15913,N_15496,N_15060);
nand U15914 (N_15914,N_15023,N_15257);
or U15915 (N_15915,N_15031,N_15566);
and U15916 (N_15916,N_15236,N_15379);
xnor U15917 (N_15917,N_15237,N_15082);
nor U15918 (N_15918,N_15195,N_15469);
nand U15919 (N_15919,N_15519,N_15582);
and U15920 (N_15920,N_15049,N_15084);
and U15921 (N_15921,N_15213,N_15253);
or U15922 (N_15922,N_15105,N_15283);
or U15923 (N_15923,N_15405,N_15593);
nor U15924 (N_15924,N_15348,N_15337);
nor U15925 (N_15925,N_15043,N_15552);
nand U15926 (N_15926,N_15044,N_15070);
nand U15927 (N_15927,N_15536,N_15472);
nor U15928 (N_15928,N_15495,N_15416);
nand U15929 (N_15929,N_15569,N_15256);
nand U15930 (N_15930,N_15577,N_15399);
and U15931 (N_15931,N_15248,N_15514);
and U15932 (N_15932,N_15420,N_15217);
nand U15933 (N_15933,N_15345,N_15070);
nor U15934 (N_15934,N_15574,N_15374);
or U15935 (N_15935,N_15145,N_15262);
xor U15936 (N_15936,N_15223,N_15396);
and U15937 (N_15937,N_15486,N_15316);
nand U15938 (N_15938,N_15232,N_15489);
nand U15939 (N_15939,N_15074,N_15385);
nand U15940 (N_15940,N_15014,N_15327);
or U15941 (N_15941,N_15091,N_15406);
nor U15942 (N_15942,N_15401,N_15488);
nand U15943 (N_15943,N_15226,N_15343);
nand U15944 (N_15944,N_15084,N_15401);
or U15945 (N_15945,N_15486,N_15472);
nand U15946 (N_15946,N_15394,N_15342);
or U15947 (N_15947,N_15068,N_15342);
nor U15948 (N_15948,N_15102,N_15015);
nand U15949 (N_15949,N_15337,N_15293);
and U15950 (N_15950,N_15224,N_15017);
nand U15951 (N_15951,N_15347,N_15271);
and U15952 (N_15952,N_15013,N_15473);
and U15953 (N_15953,N_15023,N_15376);
nand U15954 (N_15954,N_15410,N_15592);
or U15955 (N_15955,N_15472,N_15336);
and U15956 (N_15956,N_15265,N_15079);
nand U15957 (N_15957,N_15397,N_15226);
xnor U15958 (N_15958,N_15115,N_15215);
or U15959 (N_15959,N_15324,N_15320);
nand U15960 (N_15960,N_15028,N_15214);
nor U15961 (N_15961,N_15542,N_15428);
nand U15962 (N_15962,N_15013,N_15275);
nor U15963 (N_15963,N_15593,N_15375);
nor U15964 (N_15964,N_15222,N_15546);
or U15965 (N_15965,N_15257,N_15321);
or U15966 (N_15966,N_15021,N_15069);
and U15967 (N_15967,N_15338,N_15017);
xnor U15968 (N_15968,N_15387,N_15568);
and U15969 (N_15969,N_15203,N_15239);
and U15970 (N_15970,N_15411,N_15093);
nand U15971 (N_15971,N_15380,N_15177);
xor U15972 (N_15972,N_15332,N_15238);
xnor U15973 (N_15973,N_15137,N_15474);
nor U15974 (N_15974,N_15487,N_15169);
nor U15975 (N_15975,N_15392,N_15099);
nand U15976 (N_15976,N_15011,N_15534);
and U15977 (N_15977,N_15138,N_15364);
nor U15978 (N_15978,N_15512,N_15288);
and U15979 (N_15979,N_15117,N_15007);
or U15980 (N_15980,N_15340,N_15466);
or U15981 (N_15981,N_15107,N_15438);
nor U15982 (N_15982,N_15296,N_15081);
or U15983 (N_15983,N_15087,N_15255);
and U15984 (N_15984,N_15140,N_15459);
or U15985 (N_15985,N_15119,N_15539);
nand U15986 (N_15986,N_15228,N_15240);
nor U15987 (N_15987,N_15065,N_15219);
and U15988 (N_15988,N_15220,N_15256);
nor U15989 (N_15989,N_15089,N_15310);
nand U15990 (N_15990,N_15423,N_15104);
and U15991 (N_15991,N_15004,N_15079);
and U15992 (N_15992,N_15426,N_15259);
or U15993 (N_15993,N_15003,N_15410);
xor U15994 (N_15994,N_15052,N_15155);
nand U15995 (N_15995,N_15300,N_15408);
or U15996 (N_15996,N_15126,N_15120);
nand U15997 (N_15997,N_15018,N_15403);
and U15998 (N_15998,N_15423,N_15028);
or U15999 (N_15999,N_15382,N_15001);
and U16000 (N_16000,N_15043,N_15360);
nand U16001 (N_16001,N_15525,N_15376);
nand U16002 (N_16002,N_15091,N_15242);
nor U16003 (N_16003,N_15097,N_15241);
and U16004 (N_16004,N_15015,N_15573);
or U16005 (N_16005,N_15496,N_15415);
nor U16006 (N_16006,N_15477,N_15348);
or U16007 (N_16007,N_15370,N_15535);
and U16008 (N_16008,N_15059,N_15391);
and U16009 (N_16009,N_15465,N_15172);
nor U16010 (N_16010,N_15068,N_15198);
nand U16011 (N_16011,N_15084,N_15416);
and U16012 (N_16012,N_15319,N_15492);
nand U16013 (N_16013,N_15555,N_15185);
xor U16014 (N_16014,N_15331,N_15190);
nand U16015 (N_16015,N_15109,N_15017);
nand U16016 (N_16016,N_15031,N_15090);
or U16017 (N_16017,N_15258,N_15480);
nor U16018 (N_16018,N_15390,N_15027);
nand U16019 (N_16019,N_15189,N_15340);
or U16020 (N_16020,N_15328,N_15340);
nand U16021 (N_16021,N_15514,N_15105);
nand U16022 (N_16022,N_15380,N_15088);
or U16023 (N_16023,N_15351,N_15461);
and U16024 (N_16024,N_15241,N_15599);
or U16025 (N_16025,N_15317,N_15440);
or U16026 (N_16026,N_15309,N_15478);
and U16027 (N_16027,N_15150,N_15019);
nor U16028 (N_16028,N_15421,N_15189);
nand U16029 (N_16029,N_15366,N_15401);
or U16030 (N_16030,N_15490,N_15295);
or U16031 (N_16031,N_15038,N_15404);
and U16032 (N_16032,N_15145,N_15163);
and U16033 (N_16033,N_15177,N_15019);
nor U16034 (N_16034,N_15002,N_15493);
nand U16035 (N_16035,N_15301,N_15546);
or U16036 (N_16036,N_15397,N_15216);
or U16037 (N_16037,N_15485,N_15453);
or U16038 (N_16038,N_15046,N_15523);
or U16039 (N_16039,N_15226,N_15410);
nand U16040 (N_16040,N_15197,N_15142);
xnor U16041 (N_16041,N_15233,N_15398);
or U16042 (N_16042,N_15405,N_15016);
nand U16043 (N_16043,N_15140,N_15554);
nand U16044 (N_16044,N_15391,N_15156);
or U16045 (N_16045,N_15131,N_15421);
and U16046 (N_16046,N_15543,N_15067);
and U16047 (N_16047,N_15565,N_15281);
or U16048 (N_16048,N_15438,N_15345);
and U16049 (N_16049,N_15453,N_15414);
and U16050 (N_16050,N_15170,N_15197);
or U16051 (N_16051,N_15151,N_15156);
nor U16052 (N_16052,N_15516,N_15272);
nand U16053 (N_16053,N_15471,N_15193);
or U16054 (N_16054,N_15206,N_15030);
nor U16055 (N_16055,N_15359,N_15124);
and U16056 (N_16056,N_15016,N_15121);
nand U16057 (N_16057,N_15097,N_15260);
nor U16058 (N_16058,N_15008,N_15579);
nand U16059 (N_16059,N_15291,N_15511);
nand U16060 (N_16060,N_15030,N_15102);
and U16061 (N_16061,N_15063,N_15467);
nand U16062 (N_16062,N_15155,N_15519);
nor U16063 (N_16063,N_15365,N_15430);
or U16064 (N_16064,N_15151,N_15465);
xor U16065 (N_16065,N_15508,N_15171);
nand U16066 (N_16066,N_15359,N_15460);
and U16067 (N_16067,N_15488,N_15336);
xor U16068 (N_16068,N_15240,N_15229);
nand U16069 (N_16069,N_15041,N_15576);
and U16070 (N_16070,N_15291,N_15266);
nor U16071 (N_16071,N_15560,N_15160);
nand U16072 (N_16072,N_15080,N_15411);
nand U16073 (N_16073,N_15591,N_15057);
and U16074 (N_16074,N_15204,N_15075);
or U16075 (N_16075,N_15116,N_15474);
nand U16076 (N_16076,N_15450,N_15318);
nor U16077 (N_16077,N_15279,N_15355);
nand U16078 (N_16078,N_15323,N_15321);
nand U16079 (N_16079,N_15485,N_15537);
or U16080 (N_16080,N_15583,N_15047);
nor U16081 (N_16081,N_15583,N_15043);
nor U16082 (N_16082,N_15210,N_15058);
nor U16083 (N_16083,N_15307,N_15491);
nor U16084 (N_16084,N_15354,N_15434);
nand U16085 (N_16085,N_15505,N_15349);
or U16086 (N_16086,N_15059,N_15332);
and U16087 (N_16087,N_15465,N_15065);
and U16088 (N_16088,N_15298,N_15199);
or U16089 (N_16089,N_15040,N_15019);
nor U16090 (N_16090,N_15126,N_15079);
nand U16091 (N_16091,N_15017,N_15582);
and U16092 (N_16092,N_15584,N_15446);
nor U16093 (N_16093,N_15431,N_15120);
nand U16094 (N_16094,N_15304,N_15135);
nor U16095 (N_16095,N_15438,N_15045);
nor U16096 (N_16096,N_15254,N_15086);
nand U16097 (N_16097,N_15386,N_15253);
xnor U16098 (N_16098,N_15058,N_15498);
and U16099 (N_16099,N_15384,N_15285);
nand U16100 (N_16100,N_15409,N_15051);
nor U16101 (N_16101,N_15031,N_15077);
or U16102 (N_16102,N_15535,N_15479);
nand U16103 (N_16103,N_15517,N_15140);
nand U16104 (N_16104,N_15593,N_15040);
nor U16105 (N_16105,N_15053,N_15305);
nor U16106 (N_16106,N_15598,N_15511);
nor U16107 (N_16107,N_15209,N_15050);
xnor U16108 (N_16108,N_15082,N_15038);
xor U16109 (N_16109,N_15119,N_15310);
and U16110 (N_16110,N_15176,N_15565);
nand U16111 (N_16111,N_15216,N_15029);
nand U16112 (N_16112,N_15418,N_15180);
nand U16113 (N_16113,N_15228,N_15261);
nor U16114 (N_16114,N_15197,N_15369);
xnor U16115 (N_16115,N_15571,N_15194);
nand U16116 (N_16116,N_15146,N_15287);
xnor U16117 (N_16117,N_15137,N_15249);
and U16118 (N_16118,N_15228,N_15043);
nand U16119 (N_16119,N_15573,N_15485);
and U16120 (N_16120,N_15276,N_15427);
or U16121 (N_16121,N_15189,N_15079);
or U16122 (N_16122,N_15514,N_15221);
nand U16123 (N_16123,N_15357,N_15439);
nor U16124 (N_16124,N_15342,N_15266);
or U16125 (N_16125,N_15028,N_15137);
or U16126 (N_16126,N_15030,N_15559);
and U16127 (N_16127,N_15549,N_15584);
nand U16128 (N_16128,N_15075,N_15574);
and U16129 (N_16129,N_15233,N_15087);
xor U16130 (N_16130,N_15409,N_15329);
or U16131 (N_16131,N_15511,N_15162);
nand U16132 (N_16132,N_15113,N_15402);
or U16133 (N_16133,N_15497,N_15086);
nor U16134 (N_16134,N_15295,N_15502);
and U16135 (N_16135,N_15279,N_15359);
and U16136 (N_16136,N_15410,N_15166);
or U16137 (N_16137,N_15353,N_15299);
nor U16138 (N_16138,N_15425,N_15574);
nand U16139 (N_16139,N_15059,N_15303);
or U16140 (N_16140,N_15593,N_15051);
nor U16141 (N_16141,N_15193,N_15544);
or U16142 (N_16142,N_15396,N_15240);
nor U16143 (N_16143,N_15147,N_15009);
nor U16144 (N_16144,N_15478,N_15028);
and U16145 (N_16145,N_15391,N_15347);
nor U16146 (N_16146,N_15134,N_15205);
nor U16147 (N_16147,N_15162,N_15040);
nand U16148 (N_16148,N_15193,N_15474);
and U16149 (N_16149,N_15056,N_15333);
or U16150 (N_16150,N_15404,N_15118);
or U16151 (N_16151,N_15533,N_15332);
xor U16152 (N_16152,N_15115,N_15179);
or U16153 (N_16153,N_15144,N_15089);
xnor U16154 (N_16154,N_15358,N_15423);
and U16155 (N_16155,N_15361,N_15327);
xnor U16156 (N_16156,N_15372,N_15353);
nor U16157 (N_16157,N_15492,N_15386);
or U16158 (N_16158,N_15358,N_15563);
and U16159 (N_16159,N_15201,N_15318);
xnor U16160 (N_16160,N_15406,N_15127);
or U16161 (N_16161,N_15365,N_15394);
and U16162 (N_16162,N_15576,N_15116);
or U16163 (N_16163,N_15353,N_15367);
and U16164 (N_16164,N_15426,N_15538);
and U16165 (N_16165,N_15167,N_15465);
nor U16166 (N_16166,N_15048,N_15101);
nand U16167 (N_16167,N_15369,N_15509);
xnor U16168 (N_16168,N_15506,N_15080);
nor U16169 (N_16169,N_15454,N_15040);
nor U16170 (N_16170,N_15518,N_15078);
and U16171 (N_16171,N_15135,N_15439);
or U16172 (N_16172,N_15155,N_15041);
nor U16173 (N_16173,N_15196,N_15274);
nor U16174 (N_16174,N_15151,N_15344);
and U16175 (N_16175,N_15165,N_15472);
xor U16176 (N_16176,N_15019,N_15329);
and U16177 (N_16177,N_15218,N_15050);
nor U16178 (N_16178,N_15368,N_15318);
or U16179 (N_16179,N_15529,N_15485);
and U16180 (N_16180,N_15345,N_15481);
and U16181 (N_16181,N_15341,N_15527);
and U16182 (N_16182,N_15319,N_15567);
xor U16183 (N_16183,N_15534,N_15252);
nor U16184 (N_16184,N_15350,N_15319);
and U16185 (N_16185,N_15189,N_15344);
or U16186 (N_16186,N_15595,N_15545);
nor U16187 (N_16187,N_15261,N_15569);
nor U16188 (N_16188,N_15413,N_15078);
or U16189 (N_16189,N_15131,N_15498);
nand U16190 (N_16190,N_15534,N_15130);
or U16191 (N_16191,N_15280,N_15041);
nand U16192 (N_16192,N_15444,N_15417);
nor U16193 (N_16193,N_15258,N_15023);
or U16194 (N_16194,N_15567,N_15478);
and U16195 (N_16195,N_15313,N_15471);
or U16196 (N_16196,N_15137,N_15292);
nand U16197 (N_16197,N_15297,N_15590);
nand U16198 (N_16198,N_15483,N_15150);
or U16199 (N_16199,N_15346,N_15107);
xnor U16200 (N_16200,N_15733,N_15808);
nor U16201 (N_16201,N_15947,N_15757);
or U16202 (N_16202,N_15886,N_15637);
nand U16203 (N_16203,N_16019,N_16104);
or U16204 (N_16204,N_16015,N_16073);
or U16205 (N_16205,N_15866,N_15657);
nand U16206 (N_16206,N_16017,N_15704);
xor U16207 (N_16207,N_15964,N_15694);
nand U16208 (N_16208,N_15600,N_15770);
and U16209 (N_16209,N_15801,N_15812);
or U16210 (N_16210,N_15735,N_15689);
and U16211 (N_16211,N_15822,N_16131);
xnor U16212 (N_16212,N_15613,N_16086);
nand U16213 (N_16213,N_15781,N_15897);
or U16214 (N_16214,N_16167,N_15677);
or U16215 (N_16215,N_15805,N_15713);
nand U16216 (N_16216,N_16063,N_15789);
nor U16217 (N_16217,N_16119,N_16084);
nand U16218 (N_16218,N_16060,N_15797);
and U16219 (N_16219,N_16128,N_16079);
nor U16220 (N_16220,N_15852,N_15776);
nand U16221 (N_16221,N_16046,N_15666);
nor U16222 (N_16222,N_15693,N_15909);
and U16223 (N_16223,N_16016,N_15944);
and U16224 (N_16224,N_16145,N_15878);
nand U16225 (N_16225,N_15876,N_16132);
or U16226 (N_16226,N_15896,N_15857);
xor U16227 (N_16227,N_15739,N_15708);
nor U16228 (N_16228,N_15740,N_15912);
xor U16229 (N_16229,N_15969,N_15627);
nor U16230 (N_16230,N_15711,N_16149);
nand U16231 (N_16231,N_15706,N_15678);
or U16232 (N_16232,N_15721,N_15731);
and U16233 (N_16233,N_15763,N_15691);
nor U16234 (N_16234,N_15916,N_16138);
nand U16235 (N_16235,N_15765,N_15843);
or U16236 (N_16236,N_15961,N_15648);
and U16237 (N_16237,N_16035,N_15617);
or U16238 (N_16238,N_15681,N_16069);
nor U16239 (N_16239,N_15943,N_15714);
and U16240 (N_16240,N_15883,N_15702);
nor U16241 (N_16241,N_15755,N_15933);
or U16242 (N_16242,N_16133,N_16198);
nor U16243 (N_16243,N_15874,N_16142);
nand U16244 (N_16244,N_15889,N_15747);
nand U16245 (N_16245,N_15963,N_15919);
nor U16246 (N_16246,N_16177,N_15995);
and U16247 (N_16247,N_15638,N_15937);
nand U16248 (N_16248,N_15982,N_15975);
or U16249 (N_16249,N_15880,N_15741);
nand U16250 (N_16250,N_16162,N_16098);
nor U16251 (N_16251,N_15957,N_15922);
and U16252 (N_16252,N_15705,N_16173);
and U16253 (N_16253,N_16150,N_16110);
nor U16254 (N_16254,N_15811,N_15864);
and U16255 (N_16255,N_16095,N_15728);
or U16256 (N_16256,N_16169,N_15630);
xnor U16257 (N_16257,N_16179,N_15913);
and U16258 (N_16258,N_15855,N_15701);
nor U16259 (N_16259,N_16004,N_15690);
xnor U16260 (N_16260,N_15629,N_15836);
or U16261 (N_16261,N_15951,N_15831);
nor U16262 (N_16262,N_15750,N_16197);
or U16263 (N_16263,N_15732,N_15815);
nand U16264 (N_16264,N_16127,N_15625);
nor U16265 (N_16265,N_15712,N_16076);
or U16266 (N_16266,N_15980,N_15830);
or U16267 (N_16267,N_15610,N_16103);
xor U16268 (N_16268,N_16129,N_16116);
and U16269 (N_16269,N_16148,N_15838);
xor U16270 (N_16270,N_15709,N_15659);
and U16271 (N_16271,N_16165,N_16096);
and U16272 (N_16272,N_15744,N_16108);
nand U16273 (N_16273,N_16011,N_15758);
nand U16274 (N_16274,N_16092,N_15924);
and U16275 (N_16275,N_15804,N_16042);
and U16276 (N_16276,N_15954,N_15832);
nand U16277 (N_16277,N_15819,N_15968);
xor U16278 (N_16278,N_15761,N_15795);
or U16279 (N_16279,N_16083,N_16033);
and U16280 (N_16280,N_16038,N_15844);
or U16281 (N_16281,N_15906,N_15994);
or U16282 (N_16282,N_15923,N_15672);
or U16283 (N_16283,N_16176,N_16008);
nand U16284 (N_16284,N_15614,N_16171);
nor U16285 (N_16285,N_16026,N_15700);
nor U16286 (N_16286,N_15842,N_15865);
nor U16287 (N_16287,N_16022,N_15955);
or U16288 (N_16288,N_15759,N_15680);
and U16289 (N_16289,N_15620,N_16178);
and U16290 (N_16290,N_15885,N_15798);
and U16291 (N_16291,N_15940,N_16153);
and U16292 (N_16292,N_15749,N_16139);
or U16293 (N_16293,N_16041,N_16057);
nor U16294 (N_16294,N_15814,N_15766);
xor U16295 (N_16295,N_16031,N_16101);
nor U16296 (N_16296,N_16045,N_15891);
or U16297 (N_16297,N_15609,N_16053);
nand U16298 (N_16298,N_15978,N_15817);
or U16299 (N_16299,N_16075,N_16037);
or U16300 (N_16300,N_16009,N_15692);
or U16301 (N_16301,N_15958,N_16183);
nor U16302 (N_16302,N_15683,N_15626);
nor U16303 (N_16303,N_16034,N_15664);
nand U16304 (N_16304,N_15979,N_15834);
nand U16305 (N_16305,N_15942,N_15783);
or U16306 (N_16306,N_15604,N_16143);
nor U16307 (N_16307,N_16196,N_15651);
nand U16308 (N_16308,N_15742,N_15738);
or U16309 (N_16309,N_15768,N_15986);
and U16310 (N_16310,N_16146,N_15703);
and U16311 (N_16311,N_16114,N_15818);
or U16312 (N_16312,N_15729,N_16055);
and U16313 (N_16313,N_16036,N_15619);
nand U16314 (N_16314,N_15974,N_15790);
nand U16315 (N_16315,N_15697,N_16054);
nand U16316 (N_16316,N_15959,N_15917);
nor U16317 (N_16317,N_15778,N_16077);
or U16318 (N_16318,N_15928,N_15725);
or U16319 (N_16319,N_15962,N_15977);
or U16320 (N_16320,N_16126,N_15650);
and U16321 (N_16321,N_15737,N_16068);
or U16322 (N_16322,N_16005,N_15950);
or U16323 (N_16323,N_16155,N_15635);
xnor U16324 (N_16324,N_15821,N_15837);
nor U16325 (N_16325,N_16040,N_15860);
or U16326 (N_16326,N_16065,N_15948);
nand U16327 (N_16327,N_15902,N_16089);
and U16328 (N_16328,N_16074,N_15907);
nand U16329 (N_16329,N_16023,N_15661);
or U16330 (N_16330,N_15862,N_15884);
and U16331 (N_16331,N_15688,N_15859);
and U16332 (N_16332,N_15773,N_16051);
xnor U16333 (N_16333,N_16093,N_15901);
or U16334 (N_16334,N_16013,N_15956);
nand U16335 (N_16335,N_16059,N_15810);
nor U16336 (N_16336,N_15871,N_15722);
or U16337 (N_16337,N_16050,N_15935);
nor U16338 (N_16338,N_15772,N_15621);
and U16339 (N_16339,N_15800,N_15899);
and U16340 (N_16340,N_16090,N_16078);
xor U16341 (N_16341,N_15936,N_15726);
nor U16342 (N_16342,N_16071,N_15654);
nor U16343 (N_16343,N_15840,N_16062);
xnor U16344 (N_16344,N_16121,N_15828);
nand U16345 (N_16345,N_16091,N_15807);
xnor U16346 (N_16346,N_15981,N_15892);
nor U16347 (N_16347,N_16181,N_16172);
nor U16348 (N_16348,N_15816,N_15720);
nand U16349 (N_16349,N_16117,N_16120);
or U16350 (N_16350,N_16124,N_16190);
or U16351 (N_16351,N_16028,N_15839);
nand U16352 (N_16352,N_15813,N_16125);
nand U16353 (N_16353,N_15802,N_15868);
nor U16354 (N_16354,N_15825,N_15752);
nand U16355 (N_16355,N_16160,N_15983);
or U16356 (N_16356,N_16010,N_16184);
and U16357 (N_16357,N_15893,N_15673);
and U16358 (N_16358,N_15927,N_15631);
and U16359 (N_16359,N_15762,N_15753);
or U16360 (N_16360,N_15660,N_16020);
nor U16361 (N_16361,N_16175,N_15612);
nor U16362 (N_16362,N_16056,N_15925);
or U16363 (N_16363,N_16140,N_16107);
nand U16364 (N_16364,N_15966,N_15926);
and U16365 (N_16365,N_16161,N_16085);
nor U16366 (N_16366,N_16194,N_15835);
nor U16367 (N_16367,N_16122,N_15652);
nor U16368 (N_16368,N_16049,N_16134);
or U16369 (N_16369,N_15847,N_15989);
nor U16370 (N_16370,N_15777,N_15888);
and U16371 (N_16371,N_15990,N_15791);
and U16372 (N_16372,N_15973,N_16018);
and U16373 (N_16373,N_15827,N_16087);
and U16374 (N_16374,N_16152,N_15856);
nand U16375 (N_16375,N_16001,N_15931);
nor U16376 (N_16376,N_15754,N_15743);
xor U16377 (N_16377,N_15603,N_15786);
or U16378 (N_16378,N_16137,N_15915);
or U16379 (N_16379,N_15881,N_16007);
nor U16380 (N_16380,N_15696,N_16030);
nand U16381 (N_16381,N_15605,N_15751);
or U16382 (N_16382,N_16047,N_16082);
xor U16383 (N_16383,N_15903,N_15684);
and U16384 (N_16384,N_15760,N_15602);
nand U16385 (N_16385,N_15796,N_15686);
and U16386 (N_16386,N_16029,N_15939);
nor U16387 (N_16387,N_16141,N_15787);
or U16388 (N_16388,N_15767,N_15873);
nand U16389 (N_16389,N_15792,N_15829);
nand U16390 (N_16390,N_15769,N_15997);
xor U16391 (N_16391,N_16151,N_15715);
nor U16392 (N_16392,N_16163,N_15952);
and U16393 (N_16393,N_15890,N_15646);
xor U16394 (N_16394,N_15782,N_16102);
nand U16395 (N_16395,N_15938,N_15809);
nand U16396 (N_16396,N_15675,N_16100);
nand U16397 (N_16397,N_15685,N_15622);
nand U16398 (N_16398,N_15639,N_15601);
nor U16399 (N_16399,N_16058,N_15932);
nand U16400 (N_16400,N_16012,N_15988);
nand U16401 (N_16401,N_16043,N_15845);
or U16402 (N_16402,N_16106,N_16193);
nor U16403 (N_16403,N_15823,N_16072);
and U16404 (N_16404,N_15756,N_16191);
xor U16405 (N_16405,N_15820,N_16135);
or U16406 (N_16406,N_15717,N_16080);
xnor U16407 (N_16407,N_15879,N_16088);
nand U16408 (N_16408,N_16032,N_15987);
nand U16409 (N_16409,N_16111,N_15698);
nor U16410 (N_16410,N_15775,N_15846);
nor U16411 (N_16411,N_15929,N_16014);
nand U16412 (N_16412,N_15719,N_15649);
and U16413 (N_16413,N_16003,N_15920);
and U16414 (N_16414,N_16157,N_15616);
xnor U16415 (N_16415,N_16070,N_15803);
or U16416 (N_16416,N_15788,N_15953);
or U16417 (N_16417,N_15985,N_15667);
and U16418 (N_16418,N_15734,N_16025);
and U16419 (N_16419,N_15999,N_15858);
nor U16420 (N_16420,N_15628,N_15921);
nor U16421 (N_16421,N_15965,N_15679);
xor U16422 (N_16422,N_15695,N_15996);
and U16423 (N_16423,N_16048,N_15875);
nor U16424 (N_16424,N_15861,N_15647);
or U16425 (N_16425,N_15736,N_16027);
xnor U16426 (N_16426,N_15870,N_15992);
xor U16427 (N_16427,N_16192,N_16130);
and U16428 (N_16428,N_15615,N_15653);
nor U16429 (N_16429,N_16105,N_16081);
nor U16430 (N_16430,N_16168,N_16061);
nor U16431 (N_16431,N_15972,N_15641);
nor U16432 (N_16432,N_15946,N_16097);
or U16433 (N_16433,N_16052,N_15911);
and U16434 (N_16434,N_15799,N_15877);
and U16435 (N_16435,N_15779,N_15894);
xor U16436 (N_16436,N_16002,N_15707);
nor U16437 (N_16437,N_15655,N_15960);
or U16438 (N_16438,N_16144,N_16158);
nand U16439 (N_16439,N_15668,N_15748);
or U16440 (N_16440,N_16188,N_15914);
or U16441 (N_16441,N_15633,N_15716);
and U16442 (N_16442,N_15849,N_15934);
nand U16443 (N_16443,N_15687,N_16021);
xor U16444 (N_16444,N_15611,N_15918);
and U16445 (N_16445,N_15941,N_16006);
and U16446 (N_16446,N_15806,N_15841);
nor U16447 (N_16447,N_15971,N_15645);
and U16448 (N_16448,N_16099,N_15662);
nor U16449 (N_16449,N_15785,N_15710);
and U16450 (N_16450,N_15606,N_15764);
and U16451 (N_16451,N_15671,N_16195);
or U16452 (N_16452,N_16109,N_15780);
or U16453 (N_16453,N_16000,N_15624);
nand U16454 (N_16454,N_15640,N_15984);
nor U16455 (N_16455,N_16159,N_16154);
or U16456 (N_16456,N_16064,N_15970);
and U16457 (N_16457,N_16123,N_15850);
nand U16458 (N_16458,N_15900,N_15967);
xnor U16459 (N_16459,N_16136,N_15674);
or U16460 (N_16460,N_15699,N_16185);
nand U16461 (N_16461,N_16115,N_15869);
nand U16462 (N_16462,N_15993,N_15663);
or U16463 (N_16463,N_15887,N_15898);
nor U16464 (N_16464,N_15771,N_15658);
or U16465 (N_16465,N_15867,N_15682);
nor U16466 (N_16466,N_15895,N_15998);
nor U16467 (N_16467,N_15976,N_15774);
nand U16468 (N_16468,N_15793,N_16166);
or U16469 (N_16469,N_15730,N_16186);
nor U16470 (N_16470,N_15833,N_15643);
nor U16471 (N_16471,N_15669,N_15636);
nand U16472 (N_16472,N_15794,N_15945);
nand U16473 (N_16473,N_15608,N_15905);
or U16474 (N_16474,N_15618,N_15854);
nor U16475 (N_16475,N_15644,N_16187);
nand U16476 (N_16476,N_15882,N_15863);
and U16477 (N_16477,N_15745,N_15949);
xor U16478 (N_16478,N_16066,N_15904);
or U16479 (N_16479,N_16112,N_15826);
or U16480 (N_16480,N_16147,N_16182);
nand U16481 (N_16481,N_15676,N_15910);
nor U16482 (N_16482,N_15632,N_15665);
nand U16483 (N_16483,N_15670,N_16174);
nor U16484 (N_16484,N_15724,N_15853);
or U16485 (N_16485,N_15634,N_15930);
nor U16486 (N_16486,N_15908,N_16118);
or U16487 (N_16487,N_16180,N_15727);
xnor U16488 (N_16488,N_16039,N_16189);
or U16489 (N_16489,N_15848,N_16024);
nor U16490 (N_16490,N_16094,N_16156);
xnor U16491 (N_16491,N_16199,N_15623);
nor U16492 (N_16492,N_15824,N_15607);
and U16493 (N_16493,N_15718,N_15872);
or U16494 (N_16494,N_16067,N_15746);
or U16495 (N_16495,N_16044,N_15991);
or U16496 (N_16496,N_15851,N_15656);
and U16497 (N_16497,N_16113,N_16164);
xnor U16498 (N_16498,N_15784,N_16170);
nor U16499 (N_16499,N_15723,N_15642);
or U16500 (N_16500,N_16082,N_16077);
or U16501 (N_16501,N_16035,N_15607);
xor U16502 (N_16502,N_16180,N_16020);
nor U16503 (N_16503,N_16068,N_15959);
nor U16504 (N_16504,N_15863,N_15807);
or U16505 (N_16505,N_16114,N_15810);
or U16506 (N_16506,N_16106,N_15905);
nand U16507 (N_16507,N_15873,N_16170);
or U16508 (N_16508,N_15886,N_15747);
and U16509 (N_16509,N_15963,N_15988);
or U16510 (N_16510,N_15898,N_16132);
or U16511 (N_16511,N_15817,N_16134);
nor U16512 (N_16512,N_15884,N_15826);
nand U16513 (N_16513,N_16167,N_16098);
nand U16514 (N_16514,N_15918,N_15800);
nor U16515 (N_16515,N_15740,N_15940);
nor U16516 (N_16516,N_16110,N_15779);
and U16517 (N_16517,N_15948,N_16140);
and U16518 (N_16518,N_15760,N_15658);
nand U16519 (N_16519,N_15851,N_16190);
nand U16520 (N_16520,N_15801,N_15726);
or U16521 (N_16521,N_15799,N_15867);
nand U16522 (N_16522,N_15914,N_16092);
or U16523 (N_16523,N_16109,N_15669);
or U16524 (N_16524,N_15720,N_16033);
nor U16525 (N_16525,N_15615,N_15663);
or U16526 (N_16526,N_15709,N_15805);
nand U16527 (N_16527,N_15734,N_15878);
or U16528 (N_16528,N_16042,N_16051);
and U16529 (N_16529,N_15980,N_15793);
xnor U16530 (N_16530,N_15785,N_15955);
nor U16531 (N_16531,N_16150,N_15657);
nand U16532 (N_16532,N_15841,N_15752);
or U16533 (N_16533,N_15661,N_15837);
nand U16534 (N_16534,N_16024,N_16114);
nand U16535 (N_16535,N_15657,N_15641);
or U16536 (N_16536,N_16020,N_15672);
nor U16537 (N_16537,N_15642,N_16162);
xnor U16538 (N_16538,N_15971,N_16066);
xor U16539 (N_16539,N_15616,N_16084);
nor U16540 (N_16540,N_15951,N_15730);
xor U16541 (N_16541,N_15654,N_15776);
nor U16542 (N_16542,N_15721,N_15714);
and U16543 (N_16543,N_16099,N_16085);
and U16544 (N_16544,N_16159,N_15615);
nand U16545 (N_16545,N_15638,N_15863);
or U16546 (N_16546,N_15841,N_15633);
or U16547 (N_16547,N_16001,N_16032);
and U16548 (N_16548,N_15875,N_15717);
or U16549 (N_16549,N_16059,N_16100);
or U16550 (N_16550,N_15605,N_15816);
nor U16551 (N_16551,N_15729,N_15627);
or U16552 (N_16552,N_16088,N_15655);
nand U16553 (N_16553,N_15945,N_16188);
or U16554 (N_16554,N_15979,N_15982);
nand U16555 (N_16555,N_15750,N_15680);
xor U16556 (N_16556,N_15926,N_15700);
xor U16557 (N_16557,N_15766,N_15748);
or U16558 (N_16558,N_15864,N_16106);
nor U16559 (N_16559,N_15766,N_15861);
and U16560 (N_16560,N_15990,N_15900);
nor U16561 (N_16561,N_15672,N_15989);
xor U16562 (N_16562,N_15796,N_16137);
and U16563 (N_16563,N_16060,N_15841);
or U16564 (N_16564,N_15995,N_16188);
and U16565 (N_16565,N_15715,N_15753);
or U16566 (N_16566,N_16099,N_15854);
and U16567 (N_16567,N_15871,N_15761);
and U16568 (N_16568,N_16117,N_15748);
nand U16569 (N_16569,N_16129,N_16175);
nor U16570 (N_16570,N_15934,N_15678);
nand U16571 (N_16571,N_16199,N_16171);
and U16572 (N_16572,N_15777,N_15706);
nand U16573 (N_16573,N_15883,N_16020);
or U16574 (N_16574,N_16142,N_16170);
and U16575 (N_16575,N_16065,N_15923);
or U16576 (N_16576,N_15601,N_16054);
nand U16577 (N_16577,N_15837,N_15723);
and U16578 (N_16578,N_15901,N_16187);
or U16579 (N_16579,N_15668,N_16002);
and U16580 (N_16580,N_16155,N_15886);
or U16581 (N_16581,N_15913,N_15898);
nor U16582 (N_16582,N_15966,N_15973);
nor U16583 (N_16583,N_16078,N_15784);
and U16584 (N_16584,N_15951,N_16079);
or U16585 (N_16585,N_15998,N_15665);
or U16586 (N_16586,N_15898,N_15873);
and U16587 (N_16587,N_16024,N_16070);
or U16588 (N_16588,N_15842,N_15638);
nand U16589 (N_16589,N_15793,N_16150);
nor U16590 (N_16590,N_16146,N_15875);
or U16591 (N_16591,N_16053,N_16047);
or U16592 (N_16592,N_15978,N_15625);
and U16593 (N_16593,N_16058,N_15641);
or U16594 (N_16594,N_15931,N_16116);
nand U16595 (N_16595,N_15679,N_15621);
nand U16596 (N_16596,N_15600,N_15738);
nor U16597 (N_16597,N_15980,N_15765);
and U16598 (N_16598,N_15722,N_16087);
xnor U16599 (N_16599,N_15733,N_15774);
nor U16600 (N_16600,N_15674,N_15800);
nor U16601 (N_16601,N_15812,N_15745);
nor U16602 (N_16602,N_15886,N_15640);
xor U16603 (N_16603,N_15864,N_15852);
or U16604 (N_16604,N_15601,N_15870);
nor U16605 (N_16605,N_15862,N_15914);
and U16606 (N_16606,N_15795,N_15887);
and U16607 (N_16607,N_15920,N_15665);
and U16608 (N_16608,N_16060,N_15719);
nand U16609 (N_16609,N_15755,N_15858);
nor U16610 (N_16610,N_15884,N_16049);
nor U16611 (N_16611,N_15641,N_15658);
nor U16612 (N_16612,N_15757,N_15708);
nor U16613 (N_16613,N_16037,N_15864);
or U16614 (N_16614,N_15968,N_16042);
and U16615 (N_16615,N_15869,N_15850);
or U16616 (N_16616,N_16007,N_16102);
and U16617 (N_16617,N_15621,N_16148);
nand U16618 (N_16618,N_16003,N_16180);
or U16619 (N_16619,N_15918,N_15906);
xor U16620 (N_16620,N_15872,N_15672);
nand U16621 (N_16621,N_15834,N_15754);
nor U16622 (N_16622,N_15763,N_15777);
nand U16623 (N_16623,N_15961,N_16005);
and U16624 (N_16624,N_15916,N_15868);
and U16625 (N_16625,N_15685,N_15893);
nor U16626 (N_16626,N_15764,N_16067);
and U16627 (N_16627,N_16137,N_16099);
nor U16628 (N_16628,N_15649,N_15695);
nor U16629 (N_16629,N_16018,N_16196);
or U16630 (N_16630,N_16154,N_15840);
or U16631 (N_16631,N_15844,N_15911);
or U16632 (N_16632,N_15741,N_16114);
or U16633 (N_16633,N_15987,N_15810);
nand U16634 (N_16634,N_15643,N_16046);
nand U16635 (N_16635,N_15973,N_15964);
and U16636 (N_16636,N_15618,N_15893);
or U16637 (N_16637,N_15859,N_15751);
or U16638 (N_16638,N_15612,N_15799);
nand U16639 (N_16639,N_16102,N_15954);
nor U16640 (N_16640,N_15666,N_16074);
or U16641 (N_16641,N_16170,N_16159);
nor U16642 (N_16642,N_16180,N_15819);
or U16643 (N_16643,N_16054,N_15681);
nor U16644 (N_16644,N_15948,N_15841);
nor U16645 (N_16645,N_15609,N_16033);
or U16646 (N_16646,N_16156,N_16150);
nor U16647 (N_16647,N_16176,N_16161);
nor U16648 (N_16648,N_16131,N_15926);
or U16649 (N_16649,N_15660,N_15618);
or U16650 (N_16650,N_15873,N_15815);
nor U16651 (N_16651,N_16076,N_16124);
or U16652 (N_16652,N_15991,N_16003);
nor U16653 (N_16653,N_15755,N_15720);
nor U16654 (N_16654,N_16127,N_16115);
nor U16655 (N_16655,N_15787,N_16022);
or U16656 (N_16656,N_15603,N_16110);
xor U16657 (N_16657,N_16010,N_15996);
and U16658 (N_16658,N_15981,N_16084);
and U16659 (N_16659,N_15905,N_15776);
nor U16660 (N_16660,N_15929,N_15678);
or U16661 (N_16661,N_15747,N_15862);
nand U16662 (N_16662,N_15661,N_16050);
or U16663 (N_16663,N_16045,N_15740);
and U16664 (N_16664,N_15645,N_15917);
xnor U16665 (N_16665,N_15903,N_15783);
and U16666 (N_16666,N_15920,N_15605);
xnor U16667 (N_16667,N_15620,N_15851);
nor U16668 (N_16668,N_16197,N_15865);
nor U16669 (N_16669,N_16092,N_15775);
and U16670 (N_16670,N_15848,N_15629);
nand U16671 (N_16671,N_16133,N_15936);
and U16672 (N_16672,N_15762,N_15988);
xor U16673 (N_16673,N_16006,N_15857);
and U16674 (N_16674,N_15806,N_15849);
and U16675 (N_16675,N_15660,N_16100);
xor U16676 (N_16676,N_15679,N_15901);
nor U16677 (N_16677,N_16152,N_15616);
and U16678 (N_16678,N_15916,N_15664);
or U16679 (N_16679,N_15622,N_15620);
or U16680 (N_16680,N_15673,N_15788);
or U16681 (N_16681,N_16103,N_15814);
nor U16682 (N_16682,N_15607,N_15806);
and U16683 (N_16683,N_16006,N_16058);
or U16684 (N_16684,N_16111,N_15770);
or U16685 (N_16685,N_16194,N_15898);
and U16686 (N_16686,N_15724,N_15979);
or U16687 (N_16687,N_15718,N_16183);
xor U16688 (N_16688,N_15999,N_15602);
nand U16689 (N_16689,N_16085,N_15838);
and U16690 (N_16690,N_15994,N_15814);
nand U16691 (N_16691,N_16184,N_15644);
or U16692 (N_16692,N_15745,N_15680);
nand U16693 (N_16693,N_15653,N_15988);
xnor U16694 (N_16694,N_15772,N_16067);
nor U16695 (N_16695,N_16178,N_16180);
nor U16696 (N_16696,N_15834,N_15658);
and U16697 (N_16697,N_15840,N_15633);
or U16698 (N_16698,N_15805,N_15918);
nor U16699 (N_16699,N_16170,N_16161);
nand U16700 (N_16700,N_16151,N_15732);
and U16701 (N_16701,N_15802,N_15770);
and U16702 (N_16702,N_15901,N_16062);
nand U16703 (N_16703,N_15828,N_16163);
nand U16704 (N_16704,N_16196,N_16117);
and U16705 (N_16705,N_16111,N_16089);
nand U16706 (N_16706,N_15789,N_15878);
nand U16707 (N_16707,N_15899,N_16186);
and U16708 (N_16708,N_15667,N_16051);
xnor U16709 (N_16709,N_16141,N_16132);
nand U16710 (N_16710,N_16061,N_16021);
and U16711 (N_16711,N_15967,N_15936);
xor U16712 (N_16712,N_15680,N_16025);
xnor U16713 (N_16713,N_15870,N_15750);
nand U16714 (N_16714,N_15705,N_16081);
and U16715 (N_16715,N_16180,N_16111);
and U16716 (N_16716,N_15810,N_15948);
nor U16717 (N_16717,N_15851,N_15759);
nand U16718 (N_16718,N_16151,N_16082);
nand U16719 (N_16719,N_16120,N_16144);
and U16720 (N_16720,N_15823,N_16063);
or U16721 (N_16721,N_15765,N_15885);
nor U16722 (N_16722,N_15637,N_15693);
and U16723 (N_16723,N_15645,N_16081);
nand U16724 (N_16724,N_15942,N_15710);
and U16725 (N_16725,N_15780,N_15718);
xor U16726 (N_16726,N_16088,N_15639);
nor U16727 (N_16727,N_16060,N_15873);
nand U16728 (N_16728,N_15683,N_15916);
nand U16729 (N_16729,N_15932,N_16154);
and U16730 (N_16730,N_15617,N_15833);
or U16731 (N_16731,N_15616,N_16195);
nand U16732 (N_16732,N_15815,N_15828);
nor U16733 (N_16733,N_15713,N_16153);
nand U16734 (N_16734,N_15941,N_15757);
or U16735 (N_16735,N_15773,N_16027);
nand U16736 (N_16736,N_16061,N_16067);
nand U16737 (N_16737,N_15603,N_15938);
xor U16738 (N_16738,N_15767,N_15779);
nand U16739 (N_16739,N_16098,N_15843);
nor U16740 (N_16740,N_15901,N_15866);
xor U16741 (N_16741,N_15711,N_15789);
nor U16742 (N_16742,N_15712,N_16023);
or U16743 (N_16743,N_15829,N_15944);
or U16744 (N_16744,N_16141,N_16030);
nor U16745 (N_16745,N_15617,N_16044);
and U16746 (N_16746,N_16127,N_15857);
xor U16747 (N_16747,N_15957,N_15723);
nand U16748 (N_16748,N_16071,N_16165);
nand U16749 (N_16749,N_16167,N_16078);
and U16750 (N_16750,N_15735,N_15661);
and U16751 (N_16751,N_16069,N_15844);
nor U16752 (N_16752,N_15750,N_16178);
or U16753 (N_16753,N_15659,N_15676);
or U16754 (N_16754,N_15900,N_15779);
and U16755 (N_16755,N_15648,N_16184);
nor U16756 (N_16756,N_15645,N_16084);
and U16757 (N_16757,N_15705,N_15802);
nor U16758 (N_16758,N_15619,N_15752);
and U16759 (N_16759,N_15993,N_15764);
nand U16760 (N_16760,N_15703,N_16113);
nand U16761 (N_16761,N_15798,N_15693);
or U16762 (N_16762,N_15698,N_15802);
nor U16763 (N_16763,N_15683,N_15855);
nand U16764 (N_16764,N_16196,N_16033);
nand U16765 (N_16765,N_15782,N_15944);
nand U16766 (N_16766,N_15765,N_15792);
nor U16767 (N_16767,N_15667,N_16054);
nand U16768 (N_16768,N_15987,N_16198);
or U16769 (N_16769,N_15990,N_15642);
nand U16770 (N_16770,N_15689,N_15913);
or U16771 (N_16771,N_16030,N_16027);
nand U16772 (N_16772,N_15748,N_15828);
nor U16773 (N_16773,N_16053,N_15815);
xor U16774 (N_16774,N_16096,N_15869);
nand U16775 (N_16775,N_15620,N_15806);
or U16776 (N_16776,N_15982,N_15848);
nand U16777 (N_16777,N_15616,N_15937);
nor U16778 (N_16778,N_15810,N_15774);
nand U16779 (N_16779,N_16008,N_15917);
or U16780 (N_16780,N_15721,N_15605);
nand U16781 (N_16781,N_16058,N_16179);
and U16782 (N_16782,N_15805,N_15909);
or U16783 (N_16783,N_16066,N_15953);
and U16784 (N_16784,N_16074,N_15998);
nor U16785 (N_16785,N_15648,N_16043);
and U16786 (N_16786,N_16041,N_15745);
nor U16787 (N_16787,N_15932,N_15900);
or U16788 (N_16788,N_15679,N_15781);
nand U16789 (N_16789,N_15663,N_16056);
and U16790 (N_16790,N_16054,N_15862);
nand U16791 (N_16791,N_15854,N_15825);
or U16792 (N_16792,N_16121,N_15654);
xnor U16793 (N_16793,N_15864,N_15655);
nor U16794 (N_16794,N_15713,N_15615);
and U16795 (N_16795,N_15943,N_15947);
nand U16796 (N_16796,N_16165,N_15973);
nor U16797 (N_16797,N_16023,N_15837);
and U16798 (N_16798,N_15939,N_16192);
nand U16799 (N_16799,N_15856,N_15792);
nand U16800 (N_16800,N_16474,N_16745);
nor U16801 (N_16801,N_16464,N_16536);
nor U16802 (N_16802,N_16544,N_16327);
nand U16803 (N_16803,N_16755,N_16654);
or U16804 (N_16804,N_16270,N_16606);
nand U16805 (N_16805,N_16597,N_16260);
and U16806 (N_16806,N_16568,N_16400);
nand U16807 (N_16807,N_16674,N_16567);
nor U16808 (N_16808,N_16493,N_16283);
and U16809 (N_16809,N_16616,N_16459);
and U16810 (N_16810,N_16476,N_16300);
or U16811 (N_16811,N_16249,N_16794);
or U16812 (N_16812,N_16598,N_16697);
nand U16813 (N_16813,N_16246,N_16262);
xor U16814 (N_16814,N_16391,N_16271);
xor U16815 (N_16815,N_16741,N_16698);
xor U16816 (N_16816,N_16671,N_16381);
and U16817 (N_16817,N_16768,N_16710);
or U16818 (N_16818,N_16314,N_16565);
or U16819 (N_16819,N_16240,N_16204);
and U16820 (N_16820,N_16345,N_16526);
nor U16821 (N_16821,N_16328,N_16591);
nor U16822 (N_16822,N_16511,N_16492);
nand U16823 (N_16823,N_16286,N_16285);
or U16824 (N_16824,N_16469,N_16625);
nand U16825 (N_16825,N_16666,N_16217);
nand U16826 (N_16826,N_16607,N_16415);
and U16827 (N_16827,N_16471,N_16417);
nand U16828 (N_16828,N_16779,N_16570);
and U16829 (N_16829,N_16257,N_16495);
xnor U16830 (N_16830,N_16422,N_16447);
nor U16831 (N_16831,N_16349,N_16263);
and U16832 (N_16832,N_16432,N_16772);
or U16833 (N_16833,N_16449,N_16221);
nand U16834 (N_16834,N_16399,N_16727);
xnor U16835 (N_16835,N_16456,N_16206);
or U16836 (N_16836,N_16572,N_16346);
xor U16837 (N_16837,N_16664,N_16272);
or U16838 (N_16838,N_16477,N_16594);
nand U16839 (N_16839,N_16467,N_16580);
or U16840 (N_16840,N_16208,N_16401);
and U16841 (N_16841,N_16684,N_16478);
nor U16842 (N_16842,N_16281,N_16546);
xor U16843 (N_16843,N_16481,N_16627);
nor U16844 (N_16844,N_16379,N_16797);
nand U16845 (N_16845,N_16344,N_16538);
nor U16846 (N_16846,N_16776,N_16268);
nand U16847 (N_16847,N_16259,N_16309);
xor U16848 (N_16848,N_16293,N_16408);
and U16849 (N_16849,N_16239,N_16365);
xor U16850 (N_16850,N_16316,N_16515);
nand U16851 (N_16851,N_16446,N_16396);
nor U16852 (N_16852,N_16731,N_16382);
nor U16853 (N_16853,N_16795,N_16235);
nand U16854 (N_16854,N_16215,N_16641);
xor U16855 (N_16855,N_16735,N_16250);
nor U16856 (N_16856,N_16395,N_16788);
nand U16857 (N_16857,N_16413,N_16426);
or U16858 (N_16858,N_16348,N_16763);
nor U16859 (N_16859,N_16343,N_16317);
xnor U16860 (N_16860,N_16553,N_16750);
xnor U16861 (N_16861,N_16609,N_16722);
nor U16862 (N_16862,N_16740,N_16247);
and U16863 (N_16863,N_16789,N_16738);
or U16864 (N_16864,N_16587,N_16605);
nand U16865 (N_16865,N_16678,N_16751);
or U16866 (N_16866,N_16237,N_16700);
xor U16867 (N_16867,N_16455,N_16265);
and U16868 (N_16868,N_16732,N_16454);
or U16869 (N_16869,N_16528,N_16251);
xor U16870 (N_16870,N_16747,N_16397);
nor U16871 (N_16871,N_16551,N_16593);
or U16872 (N_16872,N_16611,N_16313);
or U16873 (N_16873,N_16496,N_16241);
xnor U16874 (N_16874,N_16442,N_16354);
nor U16875 (N_16875,N_16518,N_16321);
and U16876 (N_16876,N_16762,N_16424);
and U16877 (N_16877,N_16216,N_16427);
or U16878 (N_16878,N_16603,N_16554);
nor U16879 (N_16879,N_16758,N_16406);
nand U16880 (N_16880,N_16734,N_16200);
and U16881 (N_16881,N_16367,N_16621);
xnor U16882 (N_16882,N_16589,N_16307);
nand U16883 (N_16883,N_16361,N_16629);
or U16884 (N_16884,N_16729,N_16255);
nor U16885 (N_16885,N_16540,N_16383);
and U16886 (N_16886,N_16563,N_16403);
and U16887 (N_16887,N_16303,N_16480);
nor U16888 (N_16888,N_16416,N_16226);
xor U16889 (N_16889,N_16448,N_16358);
and U16890 (N_16890,N_16760,N_16227);
or U16891 (N_16891,N_16340,N_16637);
or U16892 (N_16892,N_16232,N_16347);
nor U16893 (N_16893,N_16549,N_16709);
and U16894 (N_16894,N_16503,N_16402);
nand U16895 (N_16895,N_16642,N_16213);
xnor U16896 (N_16896,N_16752,N_16470);
nand U16897 (N_16897,N_16608,N_16547);
and U16898 (N_16898,N_16244,N_16541);
and U16899 (N_16899,N_16436,N_16278);
xnor U16900 (N_16900,N_16639,N_16363);
nor U16901 (N_16901,N_16466,N_16749);
nand U16902 (N_16902,N_16502,N_16714);
and U16903 (N_16903,N_16323,N_16368);
and U16904 (N_16904,N_16438,N_16663);
nor U16905 (N_16905,N_16632,N_16719);
or U16906 (N_16906,N_16218,N_16388);
xnor U16907 (N_16907,N_16211,N_16748);
nor U16908 (N_16908,N_16421,N_16634);
or U16909 (N_16909,N_16573,N_16791);
nand U16910 (N_16910,N_16560,N_16407);
and U16911 (N_16911,N_16695,N_16592);
xor U16912 (N_16912,N_16430,N_16585);
or U16913 (N_16913,N_16444,N_16269);
nor U16914 (N_16914,N_16686,N_16513);
nand U16915 (N_16915,N_16506,N_16564);
or U16916 (N_16916,N_16356,N_16633);
and U16917 (N_16917,N_16445,N_16387);
and U16918 (N_16918,N_16780,N_16225);
or U16919 (N_16919,N_16562,N_16504);
and U16920 (N_16920,N_16394,N_16527);
nand U16921 (N_16921,N_16452,N_16352);
or U16922 (N_16922,N_16484,N_16693);
nor U16923 (N_16923,N_16312,N_16337);
nor U16924 (N_16924,N_16242,N_16766);
and U16925 (N_16925,N_16266,N_16332);
nand U16926 (N_16926,N_16465,N_16487);
nand U16927 (N_16927,N_16739,N_16588);
nor U16928 (N_16928,N_16561,N_16673);
nor U16929 (N_16929,N_16304,N_16692);
nor U16930 (N_16930,N_16708,N_16782);
and U16931 (N_16931,N_16725,N_16302);
nand U16932 (N_16932,N_16617,N_16764);
or U16933 (N_16933,N_16556,N_16482);
nand U16934 (N_16934,N_16677,N_16657);
and U16935 (N_16935,N_16569,N_16669);
or U16936 (N_16936,N_16362,N_16203);
or U16937 (N_16937,N_16428,N_16799);
or U16938 (N_16938,N_16509,N_16704);
nor U16939 (N_16939,N_16489,N_16461);
or U16940 (N_16940,N_16201,N_16559);
or U16941 (N_16941,N_16433,N_16355);
nand U16942 (N_16942,N_16679,N_16550);
nand U16943 (N_16943,N_16584,N_16214);
and U16944 (N_16944,N_16728,N_16295);
and U16945 (N_16945,N_16419,N_16276);
xor U16946 (N_16946,N_16523,N_16212);
nor U16947 (N_16947,N_16690,N_16599);
xor U16948 (N_16948,N_16586,N_16299);
nand U16949 (N_16949,N_16277,N_16298);
nor U16950 (N_16950,N_16631,N_16253);
nor U16951 (N_16951,N_16280,N_16656);
nor U16952 (N_16952,N_16672,N_16530);
nor U16953 (N_16953,N_16372,N_16434);
or U16954 (N_16954,N_16202,N_16787);
nor U16955 (N_16955,N_16648,N_16624);
nor U16956 (N_16956,N_16707,N_16575);
nand U16957 (N_16957,N_16736,N_16753);
nand U16958 (N_16958,N_16287,N_16267);
nor U16959 (N_16959,N_16770,N_16498);
or U16960 (N_16960,N_16364,N_16420);
and U16961 (N_16961,N_16497,N_16290);
and U16962 (N_16962,N_16514,N_16219);
nand U16963 (N_16963,N_16775,N_16243);
xor U16964 (N_16964,N_16310,N_16437);
xor U16965 (N_16965,N_16653,N_16668);
nor U16966 (N_16966,N_16721,N_16744);
or U16967 (N_16967,N_16357,N_16222);
or U16968 (N_16968,N_16341,N_16236);
nor U16969 (N_16969,N_16525,N_16715);
or U16970 (N_16970,N_16646,N_16404);
nand U16971 (N_16971,N_16636,N_16441);
and U16972 (N_16972,N_16712,N_16761);
and U16973 (N_16973,N_16228,N_16595);
or U16974 (N_16974,N_16360,N_16409);
and U16975 (N_16975,N_16508,N_16558);
nor U16976 (N_16976,N_16730,N_16661);
nand U16977 (N_16977,N_16548,N_16473);
nor U16978 (N_16978,N_16757,N_16618);
or U16979 (N_16979,N_16458,N_16667);
or U16980 (N_16980,N_16305,N_16398);
nor U16981 (N_16981,N_16326,N_16333);
and U16982 (N_16982,N_16318,N_16769);
nor U16983 (N_16983,N_16571,N_16539);
nor U16984 (N_16984,N_16353,N_16576);
nor U16985 (N_16985,N_16682,N_16512);
nand U16986 (N_16986,N_16288,N_16429);
nor U16987 (N_16987,N_16643,N_16702);
nand U16988 (N_16988,N_16613,N_16790);
xnor U16989 (N_16989,N_16325,N_16322);
or U16990 (N_16990,N_16291,N_16338);
or U16991 (N_16991,N_16623,N_16756);
nand U16992 (N_16992,N_16628,N_16359);
and U16993 (N_16993,N_16425,N_16462);
nor U16994 (N_16994,N_16282,N_16329);
xnor U16995 (N_16995,N_16590,N_16505);
nor U16996 (N_16996,N_16687,N_16334);
nor U16997 (N_16997,N_16274,N_16258);
nand U16998 (N_16998,N_16542,N_16742);
nand U16999 (N_16999,N_16688,N_16600);
or U17000 (N_17000,N_16670,N_16501);
or U17001 (N_17001,N_16207,N_16275);
nand U17002 (N_17002,N_16792,N_16535);
and U17003 (N_17003,N_16294,N_16414);
xnor U17004 (N_17004,N_16410,N_16431);
nor U17005 (N_17005,N_16582,N_16331);
and U17006 (N_17006,N_16650,N_16261);
xnor U17007 (N_17007,N_16279,N_16320);
or U17008 (N_17008,N_16351,N_16366);
and U17009 (N_17009,N_16231,N_16324);
nor U17010 (N_17010,N_16490,N_16578);
or U17011 (N_17011,N_16552,N_16443);
xnor U17012 (N_17012,N_16615,N_16315);
nand U17013 (N_17013,N_16308,N_16635);
nand U17014 (N_17014,N_16660,N_16798);
or U17015 (N_17015,N_16209,N_16507);
or U17016 (N_17016,N_16284,N_16596);
and U17017 (N_17017,N_16223,N_16533);
nand U17018 (N_17018,N_16785,N_16405);
or U17019 (N_17019,N_16703,N_16389);
nand U17020 (N_17020,N_16574,N_16264);
and U17021 (N_17021,N_16374,N_16524);
nand U17022 (N_17022,N_16330,N_16485);
nor U17023 (N_17023,N_16499,N_16500);
nor U17024 (N_17024,N_16786,N_16384);
nand U17025 (N_17025,N_16696,N_16460);
nor U17026 (N_17026,N_16494,N_16774);
nor U17027 (N_17027,N_16342,N_16645);
or U17028 (N_17028,N_16683,N_16457);
nand U17029 (N_17029,N_16306,N_16652);
nor U17030 (N_17030,N_16612,N_16754);
nand U17031 (N_17031,N_16675,N_16238);
or U17032 (N_17032,N_16252,N_16537);
nand U17033 (N_17033,N_16386,N_16706);
nand U17034 (N_17034,N_16411,N_16610);
xnor U17035 (N_17035,N_16651,N_16737);
nor U17036 (N_17036,N_16390,N_16665);
nand U17037 (N_17037,N_16371,N_16640);
nor U17038 (N_17038,N_16311,N_16423);
nor U17039 (N_17039,N_16453,N_16705);
nor U17040 (N_17040,N_16783,N_16681);
or U17041 (N_17041,N_16296,N_16647);
nor U17042 (N_17042,N_16450,N_16602);
and U17043 (N_17043,N_16543,N_16746);
xnor U17044 (N_17044,N_16531,N_16759);
and U17045 (N_17045,N_16796,N_16644);
and U17046 (N_17046,N_16463,N_16655);
or U17047 (N_17047,N_16604,N_16777);
xor U17048 (N_17048,N_16743,N_16778);
nor U17049 (N_17049,N_16370,N_16723);
nand U17050 (N_17050,N_16557,N_16205);
nor U17051 (N_17051,N_16614,N_16583);
nand U17052 (N_17052,N_16517,N_16676);
or U17053 (N_17053,N_16694,N_16510);
nand U17054 (N_17054,N_16577,N_16685);
or U17055 (N_17055,N_16620,N_16773);
or U17056 (N_17056,N_16724,N_16555);
and U17057 (N_17057,N_16581,N_16380);
nor U17058 (N_17058,N_16579,N_16767);
and U17059 (N_17059,N_16210,N_16335);
nand U17060 (N_17060,N_16658,N_16516);
xnor U17061 (N_17061,N_16601,N_16522);
nand U17062 (N_17062,N_16479,N_16440);
or U17063 (N_17063,N_16256,N_16234);
xor U17064 (N_17064,N_16472,N_16289);
nor U17065 (N_17065,N_16248,N_16376);
nor U17066 (N_17066,N_16626,N_16486);
and U17067 (N_17067,N_16273,N_16717);
or U17068 (N_17068,N_16720,N_16771);
or U17069 (N_17069,N_16520,N_16662);
nor U17070 (N_17070,N_16292,N_16716);
nor U17071 (N_17071,N_16319,N_16488);
or U17072 (N_17072,N_16491,N_16373);
nor U17073 (N_17073,N_16619,N_16519);
or U17074 (N_17074,N_16784,N_16726);
and U17075 (N_17075,N_16392,N_16220);
nand U17076 (N_17076,N_16393,N_16229);
or U17077 (N_17077,N_16691,N_16375);
nand U17078 (N_17078,N_16733,N_16439);
nor U17079 (N_17079,N_16301,N_16622);
and U17080 (N_17080,N_16781,N_16534);
and U17081 (N_17081,N_16468,N_16254);
nand U17082 (N_17082,N_16649,N_16701);
xor U17083 (N_17083,N_16545,N_16689);
and U17084 (N_17084,N_16233,N_16297);
and U17085 (N_17085,N_16483,N_16711);
nor U17086 (N_17086,N_16378,N_16336);
and U17087 (N_17087,N_16793,N_16475);
and U17088 (N_17088,N_16350,N_16566);
and U17089 (N_17089,N_16435,N_16659);
or U17090 (N_17090,N_16412,N_16451);
nor U17091 (N_17091,N_16699,N_16521);
nor U17092 (N_17092,N_16377,N_16529);
or U17093 (N_17093,N_16224,N_16765);
nor U17094 (N_17094,N_16230,N_16385);
and U17095 (N_17095,N_16630,N_16713);
or U17096 (N_17096,N_16680,N_16718);
or U17097 (N_17097,N_16532,N_16339);
nor U17098 (N_17098,N_16245,N_16418);
nand U17099 (N_17099,N_16638,N_16369);
and U17100 (N_17100,N_16570,N_16227);
nand U17101 (N_17101,N_16688,N_16415);
nor U17102 (N_17102,N_16785,N_16481);
nand U17103 (N_17103,N_16334,N_16463);
xor U17104 (N_17104,N_16479,N_16689);
nand U17105 (N_17105,N_16574,N_16618);
or U17106 (N_17106,N_16555,N_16637);
nand U17107 (N_17107,N_16645,N_16586);
and U17108 (N_17108,N_16799,N_16486);
nor U17109 (N_17109,N_16303,N_16649);
xor U17110 (N_17110,N_16206,N_16766);
xor U17111 (N_17111,N_16613,N_16727);
and U17112 (N_17112,N_16309,N_16595);
nor U17113 (N_17113,N_16510,N_16493);
nand U17114 (N_17114,N_16637,N_16571);
and U17115 (N_17115,N_16387,N_16474);
and U17116 (N_17116,N_16358,N_16378);
and U17117 (N_17117,N_16526,N_16594);
and U17118 (N_17118,N_16221,N_16452);
and U17119 (N_17119,N_16512,N_16422);
and U17120 (N_17120,N_16508,N_16788);
nor U17121 (N_17121,N_16677,N_16344);
and U17122 (N_17122,N_16681,N_16482);
nand U17123 (N_17123,N_16207,N_16388);
xor U17124 (N_17124,N_16718,N_16403);
nand U17125 (N_17125,N_16577,N_16513);
nand U17126 (N_17126,N_16558,N_16315);
nand U17127 (N_17127,N_16353,N_16536);
and U17128 (N_17128,N_16283,N_16796);
and U17129 (N_17129,N_16773,N_16426);
xor U17130 (N_17130,N_16305,N_16245);
and U17131 (N_17131,N_16739,N_16479);
and U17132 (N_17132,N_16609,N_16561);
nand U17133 (N_17133,N_16655,N_16279);
nor U17134 (N_17134,N_16783,N_16254);
xnor U17135 (N_17135,N_16541,N_16648);
nor U17136 (N_17136,N_16491,N_16646);
nand U17137 (N_17137,N_16724,N_16437);
and U17138 (N_17138,N_16551,N_16771);
or U17139 (N_17139,N_16728,N_16587);
nor U17140 (N_17140,N_16490,N_16389);
xnor U17141 (N_17141,N_16770,N_16634);
xor U17142 (N_17142,N_16798,N_16282);
and U17143 (N_17143,N_16778,N_16688);
or U17144 (N_17144,N_16661,N_16709);
or U17145 (N_17145,N_16291,N_16506);
xor U17146 (N_17146,N_16711,N_16634);
or U17147 (N_17147,N_16459,N_16710);
xnor U17148 (N_17148,N_16421,N_16797);
nand U17149 (N_17149,N_16264,N_16631);
and U17150 (N_17150,N_16453,N_16680);
nand U17151 (N_17151,N_16526,N_16713);
and U17152 (N_17152,N_16450,N_16459);
and U17153 (N_17153,N_16759,N_16253);
xor U17154 (N_17154,N_16567,N_16606);
and U17155 (N_17155,N_16592,N_16264);
and U17156 (N_17156,N_16204,N_16485);
xnor U17157 (N_17157,N_16362,N_16419);
nand U17158 (N_17158,N_16273,N_16539);
and U17159 (N_17159,N_16773,N_16439);
nand U17160 (N_17160,N_16582,N_16370);
nor U17161 (N_17161,N_16421,N_16208);
xor U17162 (N_17162,N_16646,N_16591);
or U17163 (N_17163,N_16633,N_16719);
nand U17164 (N_17164,N_16358,N_16563);
nand U17165 (N_17165,N_16598,N_16428);
nor U17166 (N_17166,N_16543,N_16776);
nor U17167 (N_17167,N_16390,N_16433);
nor U17168 (N_17168,N_16309,N_16438);
nand U17169 (N_17169,N_16243,N_16559);
or U17170 (N_17170,N_16332,N_16240);
nand U17171 (N_17171,N_16503,N_16661);
nor U17172 (N_17172,N_16717,N_16469);
and U17173 (N_17173,N_16492,N_16737);
nor U17174 (N_17174,N_16646,N_16219);
nand U17175 (N_17175,N_16604,N_16415);
nor U17176 (N_17176,N_16464,N_16221);
and U17177 (N_17177,N_16440,N_16699);
nand U17178 (N_17178,N_16697,N_16501);
and U17179 (N_17179,N_16688,N_16389);
nor U17180 (N_17180,N_16663,N_16298);
nand U17181 (N_17181,N_16748,N_16377);
nor U17182 (N_17182,N_16351,N_16735);
or U17183 (N_17183,N_16505,N_16796);
or U17184 (N_17184,N_16299,N_16723);
or U17185 (N_17185,N_16742,N_16609);
nor U17186 (N_17186,N_16460,N_16395);
or U17187 (N_17187,N_16746,N_16587);
and U17188 (N_17188,N_16394,N_16519);
nor U17189 (N_17189,N_16646,N_16446);
nor U17190 (N_17190,N_16450,N_16550);
and U17191 (N_17191,N_16244,N_16375);
nand U17192 (N_17192,N_16359,N_16416);
nor U17193 (N_17193,N_16678,N_16608);
nor U17194 (N_17194,N_16592,N_16790);
or U17195 (N_17195,N_16358,N_16721);
nor U17196 (N_17196,N_16491,N_16246);
nand U17197 (N_17197,N_16380,N_16667);
and U17198 (N_17198,N_16315,N_16220);
and U17199 (N_17199,N_16344,N_16626);
nand U17200 (N_17200,N_16262,N_16355);
and U17201 (N_17201,N_16281,N_16751);
nor U17202 (N_17202,N_16501,N_16793);
and U17203 (N_17203,N_16598,N_16637);
xnor U17204 (N_17204,N_16433,N_16267);
or U17205 (N_17205,N_16517,N_16540);
and U17206 (N_17206,N_16671,N_16780);
nand U17207 (N_17207,N_16735,N_16498);
nor U17208 (N_17208,N_16536,N_16206);
nor U17209 (N_17209,N_16490,N_16200);
and U17210 (N_17210,N_16252,N_16418);
or U17211 (N_17211,N_16674,N_16746);
and U17212 (N_17212,N_16404,N_16451);
or U17213 (N_17213,N_16390,N_16612);
nor U17214 (N_17214,N_16435,N_16645);
or U17215 (N_17215,N_16256,N_16716);
or U17216 (N_17216,N_16455,N_16373);
and U17217 (N_17217,N_16561,N_16302);
nand U17218 (N_17218,N_16472,N_16768);
and U17219 (N_17219,N_16776,N_16417);
nand U17220 (N_17220,N_16548,N_16719);
nand U17221 (N_17221,N_16506,N_16544);
and U17222 (N_17222,N_16624,N_16685);
nor U17223 (N_17223,N_16341,N_16448);
nand U17224 (N_17224,N_16408,N_16372);
and U17225 (N_17225,N_16278,N_16732);
nand U17226 (N_17226,N_16374,N_16655);
and U17227 (N_17227,N_16581,N_16283);
nor U17228 (N_17228,N_16657,N_16464);
and U17229 (N_17229,N_16390,N_16342);
and U17230 (N_17230,N_16486,N_16429);
or U17231 (N_17231,N_16235,N_16780);
nand U17232 (N_17232,N_16304,N_16283);
nand U17233 (N_17233,N_16330,N_16731);
nand U17234 (N_17234,N_16773,N_16770);
or U17235 (N_17235,N_16386,N_16219);
nand U17236 (N_17236,N_16229,N_16459);
and U17237 (N_17237,N_16754,N_16755);
nor U17238 (N_17238,N_16458,N_16383);
xnor U17239 (N_17239,N_16608,N_16211);
nor U17240 (N_17240,N_16351,N_16208);
and U17241 (N_17241,N_16335,N_16237);
and U17242 (N_17242,N_16266,N_16498);
xor U17243 (N_17243,N_16775,N_16317);
and U17244 (N_17244,N_16299,N_16396);
or U17245 (N_17245,N_16606,N_16482);
or U17246 (N_17246,N_16227,N_16394);
and U17247 (N_17247,N_16794,N_16338);
nand U17248 (N_17248,N_16613,N_16796);
or U17249 (N_17249,N_16731,N_16536);
or U17250 (N_17250,N_16753,N_16614);
xor U17251 (N_17251,N_16372,N_16429);
or U17252 (N_17252,N_16787,N_16301);
nand U17253 (N_17253,N_16478,N_16559);
or U17254 (N_17254,N_16399,N_16352);
or U17255 (N_17255,N_16705,N_16342);
or U17256 (N_17256,N_16792,N_16755);
xnor U17257 (N_17257,N_16263,N_16202);
and U17258 (N_17258,N_16362,N_16359);
nor U17259 (N_17259,N_16701,N_16777);
nor U17260 (N_17260,N_16519,N_16464);
or U17261 (N_17261,N_16499,N_16666);
and U17262 (N_17262,N_16347,N_16700);
nand U17263 (N_17263,N_16653,N_16771);
and U17264 (N_17264,N_16274,N_16488);
xnor U17265 (N_17265,N_16717,N_16716);
and U17266 (N_17266,N_16615,N_16277);
or U17267 (N_17267,N_16433,N_16374);
and U17268 (N_17268,N_16389,N_16732);
and U17269 (N_17269,N_16671,N_16612);
or U17270 (N_17270,N_16605,N_16631);
or U17271 (N_17271,N_16737,N_16671);
nand U17272 (N_17272,N_16796,N_16675);
and U17273 (N_17273,N_16598,N_16772);
nor U17274 (N_17274,N_16654,N_16215);
and U17275 (N_17275,N_16291,N_16500);
and U17276 (N_17276,N_16395,N_16280);
nor U17277 (N_17277,N_16302,N_16475);
nor U17278 (N_17278,N_16367,N_16544);
xnor U17279 (N_17279,N_16616,N_16771);
nor U17280 (N_17280,N_16758,N_16452);
and U17281 (N_17281,N_16289,N_16463);
nor U17282 (N_17282,N_16545,N_16475);
xor U17283 (N_17283,N_16256,N_16720);
nor U17284 (N_17284,N_16310,N_16393);
and U17285 (N_17285,N_16229,N_16622);
nand U17286 (N_17286,N_16556,N_16550);
xnor U17287 (N_17287,N_16268,N_16309);
nor U17288 (N_17288,N_16387,N_16642);
nor U17289 (N_17289,N_16350,N_16355);
and U17290 (N_17290,N_16353,N_16445);
nand U17291 (N_17291,N_16543,N_16785);
xor U17292 (N_17292,N_16793,N_16339);
and U17293 (N_17293,N_16677,N_16235);
or U17294 (N_17294,N_16794,N_16632);
xnor U17295 (N_17295,N_16244,N_16616);
nand U17296 (N_17296,N_16692,N_16646);
xnor U17297 (N_17297,N_16775,N_16263);
nand U17298 (N_17298,N_16776,N_16745);
and U17299 (N_17299,N_16448,N_16390);
and U17300 (N_17300,N_16462,N_16237);
xnor U17301 (N_17301,N_16482,N_16599);
nand U17302 (N_17302,N_16294,N_16343);
nand U17303 (N_17303,N_16298,N_16424);
or U17304 (N_17304,N_16549,N_16617);
or U17305 (N_17305,N_16217,N_16324);
nand U17306 (N_17306,N_16572,N_16456);
xnor U17307 (N_17307,N_16747,N_16428);
and U17308 (N_17308,N_16237,N_16331);
or U17309 (N_17309,N_16650,N_16537);
nor U17310 (N_17310,N_16253,N_16494);
nor U17311 (N_17311,N_16483,N_16730);
nor U17312 (N_17312,N_16480,N_16616);
and U17313 (N_17313,N_16410,N_16622);
or U17314 (N_17314,N_16722,N_16792);
nand U17315 (N_17315,N_16251,N_16236);
xor U17316 (N_17316,N_16282,N_16476);
nand U17317 (N_17317,N_16389,N_16438);
or U17318 (N_17318,N_16652,N_16339);
nand U17319 (N_17319,N_16225,N_16652);
nand U17320 (N_17320,N_16261,N_16750);
nor U17321 (N_17321,N_16301,N_16405);
or U17322 (N_17322,N_16766,N_16316);
nand U17323 (N_17323,N_16361,N_16220);
or U17324 (N_17324,N_16336,N_16318);
nor U17325 (N_17325,N_16380,N_16250);
and U17326 (N_17326,N_16223,N_16620);
nand U17327 (N_17327,N_16793,N_16465);
nor U17328 (N_17328,N_16557,N_16256);
nand U17329 (N_17329,N_16778,N_16251);
and U17330 (N_17330,N_16676,N_16279);
xnor U17331 (N_17331,N_16387,N_16213);
xor U17332 (N_17332,N_16234,N_16203);
or U17333 (N_17333,N_16560,N_16431);
nand U17334 (N_17334,N_16283,N_16469);
or U17335 (N_17335,N_16632,N_16444);
nor U17336 (N_17336,N_16644,N_16735);
xnor U17337 (N_17337,N_16396,N_16571);
and U17338 (N_17338,N_16754,N_16752);
or U17339 (N_17339,N_16689,N_16522);
nand U17340 (N_17340,N_16703,N_16543);
or U17341 (N_17341,N_16463,N_16472);
nand U17342 (N_17342,N_16292,N_16330);
nand U17343 (N_17343,N_16509,N_16732);
xnor U17344 (N_17344,N_16516,N_16287);
xor U17345 (N_17345,N_16551,N_16625);
and U17346 (N_17346,N_16205,N_16758);
xnor U17347 (N_17347,N_16569,N_16274);
xor U17348 (N_17348,N_16244,N_16360);
nand U17349 (N_17349,N_16704,N_16785);
nor U17350 (N_17350,N_16300,N_16781);
nand U17351 (N_17351,N_16623,N_16408);
nor U17352 (N_17352,N_16385,N_16358);
and U17353 (N_17353,N_16434,N_16490);
nand U17354 (N_17354,N_16236,N_16436);
nor U17355 (N_17355,N_16268,N_16784);
and U17356 (N_17356,N_16635,N_16622);
nor U17357 (N_17357,N_16510,N_16627);
or U17358 (N_17358,N_16243,N_16761);
nor U17359 (N_17359,N_16615,N_16214);
nand U17360 (N_17360,N_16607,N_16600);
nor U17361 (N_17361,N_16734,N_16414);
nand U17362 (N_17362,N_16471,N_16558);
nand U17363 (N_17363,N_16619,N_16716);
xnor U17364 (N_17364,N_16605,N_16424);
xor U17365 (N_17365,N_16617,N_16618);
or U17366 (N_17366,N_16302,N_16338);
nand U17367 (N_17367,N_16518,N_16535);
xnor U17368 (N_17368,N_16753,N_16327);
or U17369 (N_17369,N_16260,N_16616);
nand U17370 (N_17370,N_16678,N_16510);
xor U17371 (N_17371,N_16737,N_16260);
or U17372 (N_17372,N_16754,N_16718);
nor U17373 (N_17373,N_16636,N_16546);
nor U17374 (N_17374,N_16387,N_16425);
nand U17375 (N_17375,N_16432,N_16494);
and U17376 (N_17376,N_16780,N_16693);
nor U17377 (N_17377,N_16632,N_16426);
nor U17378 (N_17378,N_16333,N_16465);
or U17379 (N_17379,N_16644,N_16765);
or U17380 (N_17380,N_16339,N_16395);
nor U17381 (N_17381,N_16439,N_16230);
and U17382 (N_17382,N_16706,N_16220);
nand U17383 (N_17383,N_16412,N_16309);
and U17384 (N_17384,N_16618,N_16511);
and U17385 (N_17385,N_16311,N_16211);
nand U17386 (N_17386,N_16263,N_16394);
and U17387 (N_17387,N_16361,N_16506);
or U17388 (N_17388,N_16291,N_16406);
nor U17389 (N_17389,N_16700,N_16391);
nand U17390 (N_17390,N_16487,N_16703);
and U17391 (N_17391,N_16246,N_16274);
nor U17392 (N_17392,N_16583,N_16646);
and U17393 (N_17393,N_16267,N_16721);
or U17394 (N_17394,N_16742,N_16726);
and U17395 (N_17395,N_16353,N_16529);
nor U17396 (N_17396,N_16372,N_16764);
nor U17397 (N_17397,N_16519,N_16439);
nand U17398 (N_17398,N_16380,N_16221);
and U17399 (N_17399,N_16351,N_16491);
or U17400 (N_17400,N_17244,N_17315);
nor U17401 (N_17401,N_17106,N_17299);
xnor U17402 (N_17402,N_17004,N_17263);
xor U17403 (N_17403,N_17364,N_16839);
or U17404 (N_17404,N_16994,N_17352);
nor U17405 (N_17405,N_17143,N_17129);
or U17406 (N_17406,N_17121,N_16989);
and U17407 (N_17407,N_16905,N_17387);
nor U17408 (N_17408,N_16842,N_17309);
and U17409 (N_17409,N_16931,N_16964);
or U17410 (N_17410,N_17250,N_17378);
nor U17411 (N_17411,N_17183,N_16906);
or U17412 (N_17412,N_17031,N_16975);
or U17413 (N_17413,N_16932,N_17395);
nor U17414 (N_17414,N_16849,N_16820);
or U17415 (N_17415,N_17115,N_16901);
and U17416 (N_17416,N_17032,N_17148);
xnor U17417 (N_17417,N_16904,N_17009);
and U17418 (N_17418,N_17014,N_17365);
or U17419 (N_17419,N_16859,N_17288);
or U17420 (N_17420,N_16899,N_16982);
or U17421 (N_17421,N_16995,N_16981);
nor U17422 (N_17422,N_16879,N_16959);
or U17423 (N_17423,N_16967,N_17030);
nor U17424 (N_17424,N_16850,N_17381);
or U17425 (N_17425,N_16869,N_16985);
nand U17426 (N_17426,N_17164,N_17191);
and U17427 (N_17427,N_16854,N_17310);
nor U17428 (N_17428,N_17307,N_16939);
nand U17429 (N_17429,N_16993,N_17260);
and U17430 (N_17430,N_17220,N_16917);
nor U17431 (N_17431,N_16963,N_17169);
and U17432 (N_17432,N_16808,N_17335);
nand U17433 (N_17433,N_17186,N_16862);
nand U17434 (N_17434,N_17253,N_16857);
nand U17435 (N_17435,N_17372,N_17005);
xor U17436 (N_17436,N_17059,N_17218);
nor U17437 (N_17437,N_16937,N_17157);
or U17438 (N_17438,N_16884,N_16867);
nand U17439 (N_17439,N_16809,N_17092);
nand U17440 (N_17440,N_17391,N_17346);
and U17441 (N_17441,N_16980,N_17015);
nor U17442 (N_17442,N_16916,N_16825);
and U17443 (N_17443,N_17073,N_17242);
nand U17444 (N_17444,N_16840,N_17010);
nand U17445 (N_17445,N_16816,N_17347);
xnor U17446 (N_17446,N_17227,N_16903);
or U17447 (N_17447,N_16837,N_17167);
nand U17448 (N_17448,N_17174,N_16900);
or U17449 (N_17449,N_16977,N_17246);
and U17450 (N_17450,N_17131,N_17377);
nand U17451 (N_17451,N_17130,N_17057);
and U17452 (N_17452,N_16944,N_17285);
nand U17453 (N_17453,N_17081,N_16845);
and U17454 (N_17454,N_17256,N_17234);
nor U17455 (N_17455,N_16946,N_17105);
xnor U17456 (N_17456,N_17308,N_16934);
or U17457 (N_17457,N_17279,N_16970);
and U17458 (N_17458,N_16880,N_16999);
nand U17459 (N_17459,N_17240,N_16924);
xor U17460 (N_17460,N_17125,N_16908);
and U17461 (N_17461,N_17063,N_16914);
nand U17462 (N_17462,N_17089,N_16812);
xor U17463 (N_17463,N_17231,N_16827);
nor U17464 (N_17464,N_17075,N_17209);
and U17465 (N_17465,N_17257,N_17385);
and U17466 (N_17466,N_17193,N_17120);
and U17467 (N_17467,N_17393,N_16915);
or U17468 (N_17468,N_17002,N_16962);
nand U17469 (N_17469,N_17271,N_17196);
or U17470 (N_17470,N_17275,N_16887);
and U17471 (N_17471,N_17181,N_16949);
nand U17472 (N_17472,N_17062,N_17079);
nand U17473 (N_17473,N_17017,N_16966);
or U17474 (N_17474,N_17328,N_17388);
xor U17475 (N_17475,N_17025,N_17287);
xnor U17476 (N_17476,N_17190,N_17095);
nand U17477 (N_17477,N_17291,N_17053);
nor U17478 (N_17478,N_17072,N_17083);
nor U17479 (N_17479,N_17138,N_17333);
nand U17480 (N_17480,N_16955,N_17329);
nand U17481 (N_17481,N_17068,N_17286);
nor U17482 (N_17482,N_17172,N_17213);
or U17483 (N_17483,N_17300,N_17272);
and U17484 (N_17484,N_17319,N_17156);
and U17485 (N_17485,N_17036,N_17166);
and U17486 (N_17486,N_17254,N_17026);
or U17487 (N_17487,N_16953,N_16947);
or U17488 (N_17488,N_17290,N_16886);
nor U17489 (N_17489,N_16978,N_17197);
nand U17490 (N_17490,N_17248,N_17019);
and U17491 (N_17491,N_17216,N_16851);
or U17492 (N_17492,N_17187,N_17249);
nand U17493 (N_17493,N_17200,N_17359);
nand U17494 (N_17494,N_17219,N_17282);
or U17495 (N_17495,N_17070,N_17323);
and U17496 (N_17496,N_17080,N_17204);
or U17497 (N_17497,N_17350,N_17112);
or U17498 (N_17498,N_17135,N_16984);
nand U17499 (N_17499,N_16865,N_16818);
and U17500 (N_17500,N_17016,N_16822);
xor U17501 (N_17501,N_17238,N_17382);
nand U17502 (N_17502,N_16821,N_17389);
xor U17503 (N_17503,N_17397,N_17304);
or U17504 (N_17504,N_16873,N_16918);
nor U17505 (N_17505,N_17383,N_17332);
nand U17506 (N_17506,N_17044,N_16803);
nor U17507 (N_17507,N_17047,N_17008);
or U17508 (N_17508,N_17178,N_17142);
xor U17509 (N_17509,N_16942,N_17306);
and U17510 (N_17510,N_17163,N_17154);
or U17511 (N_17511,N_16891,N_17192);
and U17512 (N_17512,N_16909,N_16872);
xor U17513 (N_17513,N_17399,N_17311);
nor U17514 (N_17514,N_16968,N_17007);
xor U17515 (N_17515,N_17087,N_17093);
xnor U17516 (N_17516,N_16958,N_17338);
and U17517 (N_17517,N_16890,N_16875);
and U17518 (N_17518,N_17066,N_17180);
and U17519 (N_17519,N_17233,N_17039);
and U17520 (N_17520,N_17085,N_16921);
and U17521 (N_17521,N_17340,N_16801);
and U17522 (N_17522,N_16894,N_16888);
nand U17523 (N_17523,N_17045,N_16861);
and U17524 (N_17524,N_17114,N_17262);
and U17525 (N_17525,N_17111,N_16852);
xnor U17526 (N_17526,N_17296,N_16834);
or U17527 (N_17527,N_17124,N_17176);
and U17528 (N_17528,N_17274,N_17221);
or U17529 (N_17529,N_17116,N_16961);
or U17530 (N_17530,N_17123,N_17302);
nor U17531 (N_17531,N_17363,N_16826);
or U17532 (N_17532,N_17273,N_17358);
nand U17533 (N_17533,N_17136,N_16895);
nand U17534 (N_17534,N_17202,N_17342);
nand U17535 (N_17535,N_16907,N_17050);
nand U17536 (N_17536,N_17327,N_16844);
nor U17537 (N_17537,N_17368,N_17021);
or U17538 (N_17538,N_17100,N_17398);
and U17539 (N_17539,N_17098,N_17033);
xor U17540 (N_17540,N_16829,N_16863);
and U17541 (N_17541,N_17108,N_17203);
nor U17542 (N_17542,N_17243,N_16965);
nand U17543 (N_17543,N_17259,N_17185);
xnor U17544 (N_17544,N_17184,N_17366);
and U17545 (N_17545,N_17305,N_17146);
xor U17546 (N_17546,N_17149,N_16878);
and U17547 (N_17547,N_17023,N_17265);
nand U17548 (N_17548,N_17226,N_17090);
or U17549 (N_17549,N_17054,N_17224);
nor U17550 (N_17550,N_17386,N_16979);
xor U17551 (N_17551,N_17295,N_17225);
nor U17552 (N_17552,N_16853,N_17069);
and U17553 (N_17553,N_17316,N_16896);
or U17554 (N_17554,N_16929,N_17228);
and U17555 (N_17555,N_17109,N_16838);
and U17556 (N_17556,N_17049,N_17268);
nor U17557 (N_17557,N_17162,N_17006);
nand U17558 (N_17558,N_17147,N_17312);
or U17559 (N_17559,N_17195,N_17289);
and U17560 (N_17560,N_17153,N_17040);
and U17561 (N_17561,N_16988,N_17003);
nand U17562 (N_17562,N_17020,N_17188);
nand U17563 (N_17563,N_17237,N_16972);
nor U17564 (N_17564,N_16828,N_17038);
nand U17565 (N_17565,N_17326,N_17379);
and U17566 (N_17566,N_17322,N_17133);
nor U17567 (N_17567,N_17127,N_16856);
and U17568 (N_17568,N_17351,N_17370);
nor U17569 (N_17569,N_16866,N_17018);
or U17570 (N_17570,N_16974,N_16928);
and U17571 (N_17571,N_17277,N_17064);
or U17572 (N_17572,N_17082,N_16943);
and U17573 (N_17573,N_17284,N_16912);
or U17574 (N_17574,N_16902,N_16831);
nor U17575 (N_17575,N_16833,N_16933);
and U17576 (N_17576,N_17171,N_17076);
nor U17577 (N_17577,N_16941,N_17028);
nor U17578 (N_17578,N_17141,N_17128);
xor U17579 (N_17579,N_16889,N_16990);
and U17580 (N_17580,N_16973,N_17074);
and U17581 (N_17581,N_16986,N_17303);
nand U17582 (N_17582,N_17217,N_16960);
or U17583 (N_17583,N_16956,N_16885);
or U17584 (N_17584,N_16874,N_17375);
nor U17585 (N_17585,N_17232,N_16800);
and U17586 (N_17586,N_17107,N_17339);
nor U17587 (N_17587,N_17235,N_16835);
nand U17588 (N_17588,N_16860,N_16807);
and U17589 (N_17589,N_17276,N_17205);
and U17590 (N_17590,N_17215,N_16938);
nand U17591 (N_17591,N_17252,N_16814);
nor U17592 (N_17592,N_17345,N_16892);
nor U17593 (N_17593,N_17035,N_17318);
and U17594 (N_17594,N_16935,N_17043);
nor U17595 (N_17595,N_16925,N_16971);
and U17596 (N_17596,N_17000,N_17103);
nor U17597 (N_17597,N_17159,N_17170);
and U17598 (N_17598,N_16987,N_17251);
nand U17599 (N_17599,N_16951,N_16893);
or U17600 (N_17600,N_17281,N_17241);
or U17601 (N_17601,N_17126,N_17118);
nand U17602 (N_17602,N_17024,N_16832);
or U17603 (N_17603,N_17336,N_17194);
nor U17604 (N_17604,N_17236,N_17212);
and U17605 (N_17605,N_17201,N_17320);
or U17606 (N_17606,N_16824,N_17354);
xor U17607 (N_17607,N_16898,N_17152);
or U17608 (N_17608,N_16913,N_17280);
nor U17609 (N_17609,N_17042,N_16868);
or U17610 (N_17610,N_17060,N_17283);
or U17611 (N_17611,N_17099,N_17230);
or U17612 (N_17612,N_17222,N_16848);
and U17613 (N_17613,N_17071,N_17097);
xor U17614 (N_17614,N_17065,N_17353);
and U17615 (N_17615,N_16940,N_17261);
xor U17616 (N_17616,N_16805,N_17369);
or U17617 (N_17617,N_17058,N_17094);
nor U17618 (N_17618,N_17078,N_17376);
nor U17619 (N_17619,N_16920,N_17361);
xnor U17620 (N_17620,N_17046,N_16811);
and U17621 (N_17621,N_17314,N_16911);
or U17622 (N_17622,N_16817,N_16883);
or U17623 (N_17623,N_17210,N_16952);
and U17624 (N_17624,N_17037,N_17343);
or U17625 (N_17625,N_17144,N_16922);
and U17626 (N_17626,N_17177,N_17384);
nand U17627 (N_17627,N_16876,N_17104);
nand U17628 (N_17628,N_17012,N_17145);
nand U17629 (N_17629,N_17313,N_17301);
nand U17630 (N_17630,N_17168,N_17214);
nor U17631 (N_17631,N_17294,N_17396);
nor U17632 (N_17632,N_17110,N_17349);
nor U17633 (N_17633,N_17119,N_16998);
and U17634 (N_17634,N_17264,N_16813);
and U17635 (N_17635,N_17206,N_16926);
or U17636 (N_17636,N_17086,N_17122);
nand U17637 (N_17637,N_17077,N_16983);
and U17638 (N_17638,N_17132,N_16877);
or U17639 (N_17639,N_17330,N_17139);
xnor U17640 (N_17640,N_17334,N_17325);
and U17641 (N_17641,N_17380,N_16806);
and U17642 (N_17642,N_17298,N_17362);
or U17643 (N_17643,N_17140,N_16910);
and U17644 (N_17644,N_17392,N_16969);
and U17645 (N_17645,N_17293,N_17113);
nand U17646 (N_17646,N_17344,N_17048);
nand U17647 (N_17647,N_17067,N_16919);
xnor U17648 (N_17648,N_16815,N_16855);
nor U17649 (N_17649,N_16802,N_17374);
nand U17650 (N_17650,N_17101,N_16991);
nor U17651 (N_17651,N_17245,N_16847);
or U17652 (N_17652,N_16870,N_17255);
nand U17653 (N_17653,N_16858,N_16823);
nor U17654 (N_17654,N_16819,N_17189);
nand U17655 (N_17655,N_17013,N_17223);
and U17656 (N_17656,N_17034,N_17137);
nor U17657 (N_17657,N_16976,N_17151);
and U17658 (N_17658,N_17348,N_16927);
and U17659 (N_17659,N_17102,N_17292);
and U17660 (N_17660,N_17158,N_17199);
nor U17661 (N_17661,N_17160,N_17084);
or U17662 (N_17662,N_16864,N_17390);
or U17663 (N_17663,N_16846,N_17229);
nand U17664 (N_17664,N_16992,N_17051);
nand U17665 (N_17665,N_17207,N_17096);
xor U17666 (N_17666,N_17337,N_17371);
and U17667 (N_17667,N_16945,N_17258);
nor U17668 (N_17668,N_17341,N_17357);
nor U17669 (N_17669,N_17270,N_16923);
or U17670 (N_17670,N_16810,N_17055);
nand U17671 (N_17671,N_16871,N_16830);
nor U17672 (N_17672,N_17027,N_17029);
xnor U17673 (N_17673,N_17267,N_17324);
or U17674 (N_17674,N_17022,N_17278);
and U17675 (N_17675,N_17041,N_16804);
xnor U17676 (N_17676,N_17394,N_17247);
nand U17677 (N_17677,N_16836,N_17134);
or U17678 (N_17678,N_16957,N_16997);
or U17679 (N_17679,N_16881,N_16948);
xnor U17680 (N_17680,N_17001,N_16843);
and U17681 (N_17681,N_17211,N_17165);
and U17682 (N_17682,N_17179,N_17155);
nand U17683 (N_17683,N_17088,N_17356);
nor U17684 (N_17684,N_16954,N_17161);
or U17685 (N_17685,N_17208,N_17269);
and U17686 (N_17686,N_17321,N_17373);
and U17687 (N_17687,N_17360,N_16996);
nor U17688 (N_17688,N_17331,N_17117);
nor U17689 (N_17689,N_17266,N_16841);
nor U17690 (N_17690,N_17091,N_17175);
and U17691 (N_17691,N_17355,N_16930);
nand U17692 (N_17692,N_17061,N_17052);
and U17693 (N_17693,N_17317,N_17173);
nor U17694 (N_17694,N_16950,N_17198);
or U17695 (N_17695,N_17056,N_17297);
nor U17696 (N_17696,N_16882,N_16936);
or U17697 (N_17697,N_17182,N_16897);
nand U17698 (N_17698,N_17011,N_17150);
or U17699 (N_17699,N_17239,N_17367);
and U17700 (N_17700,N_16971,N_17371);
nand U17701 (N_17701,N_17122,N_17397);
nor U17702 (N_17702,N_16840,N_17036);
and U17703 (N_17703,N_17125,N_17109);
or U17704 (N_17704,N_17227,N_16964);
and U17705 (N_17705,N_17141,N_16883);
nor U17706 (N_17706,N_16804,N_16825);
and U17707 (N_17707,N_16922,N_17068);
and U17708 (N_17708,N_16950,N_17383);
nor U17709 (N_17709,N_17020,N_16854);
and U17710 (N_17710,N_16948,N_17266);
nand U17711 (N_17711,N_16926,N_16997);
nor U17712 (N_17712,N_17018,N_17068);
nand U17713 (N_17713,N_17278,N_16932);
xor U17714 (N_17714,N_17177,N_17013);
nor U17715 (N_17715,N_16986,N_16830);
or U17716 (N_17716,N_17239,N_17179);
or U17717 (N_17717,N_17350,N_17126);
or U17718 (N_17718,N_16842,N_16826);
and U17719 (N_17719,N_17273,N_17030);
xor U17720 (N_17720,N_17080,N_17343);
and U17721 (N_17721,N_17215,N_16845);
nor U17722 (N_17722,N_16943,N_16844);
nor U17723 (N_17723,N_17005,N_16932);
or U17724 (N_17724,N_17199,N_17064);
nand U17725 (N_17725,N_16913,N_17287);
or U17726 (N_17726,N_17381,N_17196);
nor U17727 (N_17727,N_17395,N_16892);
nand U17728 (N_17728,N_17396,N_17341);
nor U17729 (N_17729,N_17269,N_17308);
or U17730 (N_17730,N_17270,N_16826);
xor U17731 (N_17731,N_17138,N_16958);
or U17732 (N_17732,N_17251,N_17287);
or U17733 (N_17733,N_16893,N_17265);
nand U17734 (N_17734,N_17137,N_17109);
nand U17735 (N_17735,N_17151,N_17314);
and U17736 (N_17736,N_17103,N_17351);
nand U17737 (N_17737,N_16984,N_17113);
nor U17738 (N_17738,N_17141,N_17010);
nand U17739 (N_17739,N_16970,N_16869);
nand U17740 (N_17740,N_17397,N_16934);
nor U17741 (N_17741,N_17139,N_16983);
and U17742 (N_17742,N_17120,N_17334);
and U17743 (N_17743,N_17086,N_16930);
nor U17744 (N_17744,N_17357,N_16890);
or U17745 (N_17745,N_17316,N_16958);
nor U17746 (N_17746,N_17207,N_17228);
or U17747 (N_17747,N_16959,N_16939);
or U17748 (N_17748,N_17073,N_17323);
or U17749 (N_17749,N_16998,N_16904);
nand U17750 (N_17750,N_17000,N_17321);
nor U17751 (N_17751,N_17084,N_17328);
or U17752 (N_17752,N_17206,N_17059);
and U17753 (N_17753,N_17379,N_17391);
or U17754 (N_17754,N_16882,N_17375);
nor U17755 (N_17755,N_17118,N_17316);
or U17756 (N_17756,N_16970,N_17157);
and U17757 (N_17757,N_17274,N_17298);
nor U17758 (N_17758,N_17118,N_16833);
and U17759 (N_17759,N_16976,N_16949);
nand U17760 (N_17760,N_16900,N_17103);
nor U17761 (N_17761,N_16908,N_17076);
and U17762 (N_17762,N_17263,N_17114);
nand U17763 (N_17763,N_17004,N_17107);
and U17764 (N_17764,N_16844,N_17151);
or U17765 (N_17765,N_17015,N_17088);
and U17766 (N_17766,N_17352,N_17358);
or U17767 (N_17767,N_17126,N_16824);
and U17768 (N_17768,N_16866,N_17306);
nor U17769 (N_17769,N_17121,N_16872);
nand U17770 (N_17770,N_16875,N_16954);
and U17771 (N_17771,N_16899,N_17200);
nor U17772 (N_17772,N_17012,N_17246);
nor U17773 (N_17773,N_17026,N_17098);
nand U17774 (N_17774,N_17253,N_17111);
and U17775 (N_17775,N_17005,N_16894);
nor U17776 (N_17776,N_17096,N_17002);
and U17777 (N_17777,N_16927,N_16902);
nor U17778 (N_17778,N_17037,N_17309);
and U17779 (N_17779,N_16989,N_17119);
or U17780 (N_17780,N_17032,N_16808);
nand U17781 (N_17781,N_16867,N_16853);
nor U17782 (N_17782,N_16887,N_17019);
nor U17783 (N_17783,N_16975,N_17008);
nand U17784 (N_17784,N_16883,N_17175);
nor U17785 (N_17785,N_16803,N_17339);
nor U17786 (N_17786,N_16921,N_16831);
nor U17787 (N_17787,N_16999,N_17295);
nor U17788 (N_17788,N_16854,N_16936);
nor U17789 (N_17789,N_16868,N_17188);
nand U17790 (N_17790,N_17072,N_17354);
or U17791 (N_17791,N_16875,N_16847);
and U17792 (N_17792,N_16971,N_16932);
and U17793 (N_17793,N_17196,N_16927);
or U17794 (N_17794,N_16842,N_17045);
or U17795 (N_17795,N_17327,N_17246);
nor U17796 (N_17796,N_16963,N_16800);
nand U17797 (N_17797,N_16989,N_17118);
and U17798 (N_17798,N_16832,N_16985);
nor U17799 (N_17799,N_17010,N_17246);
or U17800 (N_17800,N_17236,N_16968);
xor U17801 (N_17801,N_16905,N_17258);
xnor U17802 (N_17802,N_17092,N_17372);
and U17803 (N_17803,N_17342,N_17134);
xor U17804 (N_17804,N_17204,N_17229);
and U17805 (N_17805,N_17277,N_17399);
or U17806 (N_17806,N_17290,N_16826);
and U17807 (N_17807,N_16826,N_17201);
or U17808 (N_17808,N_17108,N_17355);
and U17809 (N_17809,N_16943,N_17329);
and U17810 (N_17810,N_17204,N_16968);
nand U17811 (N_17811,N_17056,N_17205);
nor U17812 (N_17812,N_17162,N_17240);
or U17813 (N_17813,N_16931,N_17376);
and U17814 (N_17814,N_17135,N_17011);
nand U17815 (N_17815,N_17001,N_17321);
and U17816 (N_17816,N_17262,N_17238);
nor U17817 (N_17817,N_16802,N_16973);
or U17818 (N_17818,N_17295,N_17215);
or U17819 (N_17819,N_16820,N_17011);
nand U17820 (N_17820,N_16937,N_16909);
and U17821 (N_17821,N_17341,N_17399);
nand U17822 (N_17822,N_17325,N_16959);
and U17823 (N_17823,N_16935,N_17376);
nor U17824 (N_17824,N_16908,N_16865);
nor U17825 (N_17825,N_17188,N_17233);
or U17826 (N_17826,N_17225,N_17361);
xor U17827 (N_17827,N_17274,N_16882);
nand U17828 (N_17828,N_16811,N_16995);
nor U17829 (N_17829,N_17244,N_17175);
xor U17830 (N_17830,N_16936,N_17374);
nor U17831 (N_17831,N_17036,N_17014);
nor U17832 (N_17832,N_17282,N_17267);
or U17833 (N_17833,N_16886,N_17293);
or U17834 (N_17834,N_17027,N_17178);
and U17835 (N_17835,N_17226,N_17059);
xor U17836 (N_17836,N_16998,N_16961);
and U17837 (N_17837,N_17104,N_17261);
or U17838 (N_17838,N_17326,N_17354);
nand U17839 (N_17839,N_17164,N_17009);
nand U17840 (N_17840,N_17056,N_16846);
or U17841 (N_17841,N_16855,N_16833);
nand U17842 (N_17842,N_16971,N_17079);
nor U17843 (N_17843,N_16956,N_17270);
and U17844 (N_17844,N_17363,N_16922);
and U17845 (N_17845,N_16957,N_16924);
and U17846 (N_17846,N_17105,N_17376);
and U17847 (N_17847,N_16806,N_17221);
nor U17848 (N_17848,N_16815,N_16917);
and U17849 (N_17849,N_16846,N_17260);
or U17850 (N_17850,N_17214,N_17245);
nor U17851 (N_17851,N_17380,N_16818);
xor U17852 (N_17852,N_16813,N_17153);
nand U17853 (N_17853,N_16912,N_17184);
xor U17854 (N_17854,N_17169,N_16937);
xor U17855 (N_17855,N_17208,N_17140);
nand U17856 (N_17856,N_17342,N_17072);
and U17857 (N_17857,N_16898,N_17108);
xnor U17858 (N_17858,N_17373,N_16813);
and U17859 (N_17859,N_17180,N_17316);
nor U17860 (N_17860,N_17358,N_17148);
nor U17861 (N_17861,N_17346,N_17141);
nor U17862 (N_17862,N_17170,N_17311);
nand U17863 (N_17863,N_16897,N_17264);
nand U17864 (N_17864,N_17332,N_16904);
and U17865 (N_17865,N_16820,N_17113);
nor U17866 (N_17866,N_17234,N_17308);
nor U17867 (N_17867,N_17398,N_17251);
and U17868 (N_17868,N_17089,N_16880);
nor U17869 (N_17869,N_16803,N_17261);
nand U17870 (N_17870,N_17325,N_17048);
nand U17871 (N_17871,N_16806,N_16855);
or U17872 (N_17872,N_16956,N_17040);
nand U17873 (N_17873,N_17115,N_17399);
nand U17874 (N_17874,N_16948,N_17211);
nor U17875 (N_17875,N_17354,N_17162);
xor U17876 (N_17876,N_17254,N_17044);
nor U17877 (N_17877,N_16870,N_17254);
xnor U17878 (N_17878,N_17322,N_16896);
nor U17879 (N_17879,N_17302,N_17298);
nand U17880 (N_17880,N_17200,N_17179);
nand U17881 (N_17881,N_17351,N_17303);
nand U17882 (N_17882,N_17202,N_16823);
nand U17883 (N_17883,N_17152,N_16969);
and U17884 (N_17884,N_17211,N_16852);
nand U17885 (N_17885,N_16841,N_17206);
nor U17886 (N_17886,N_17080,N_16894);
nor U17887 (N_17887,N_16998,N_16905);
nand U17888 (N_17888,N_17210,N_17355);
or U17889 (N_17889,N_17306,N_17359);
nor U17890 (N_17890,N_16995,N_17099);
or U17891 (N_17891,N_17006,N_17211);
nor U17892 (N_17892,N_17194,N_17307);
and U17893 (N_17893,N_16891,N_16814);
and U17894 (N_17894,N_17376,N_17267);
nor U17895 (N_17895,N_16906,N_17196);
or U17896 (N_17896,N_16883,N_16855);
or U17897 (N_17897,N_16981,N_17178);
and U17898 (N_17898,N_16818,N_16909);
nand U17899 (N_17899,N_17065,N_17077);
xnor U17900 (N_17900,N_17272,N_17321);
or U17901 (N_17901,N_16844,N_16971);
nand U17902 (N_17902,N_17321,N_16830);
nor U17903 (N_17903,N_17219,N_16968);
nor U17904 (N_17904,N_16839,N_17078);
and U17905 (N_17905,N_17261,N_16865);
xor U17906 (N_17906,N_16829,N_16888);
or U17907 (N_17907,N_16933,N_17384);
nor U17908 (N_17908,N_17263,N_17245);
xor U17909 (N_17909,N_17004,N_16921);
or U17910 (N_17910,N_17317,N_16898);
and U17911 (N_17911,N_16924,N_17387);
and U17912 (N_17912,N_17130,N_16900);
nand U17913 (N_17913,N_17239,N_17225);
nor U17914 (N_17914,N_16854,N_17044);
xnor U17915 (N_17915,N_17171,N_17035);
xor U17916 (N_17916,N_17131,N_16901);
nor U17917 (N_17917,N_16911,N_17185);
or U17918 (N_17918,N_16932,N_17028);
or U17919 (N_17919,N_17289,N_17373);
or U17920 (N_17920,N_17128,N_17055);
nand U17921 (N_17921,N_17264,N_16950);
and U17922 (N_17922,N_16934,N_16846);
and U17923 (N_17923,N_16811,N_17324);
and U17924 (N_17924,N_16942,N_16988);
or U17925 (N_17925,N_17345,N_17073);
nor U17926 (N_17926,N_16803,N_16978);
and U17927 (N_17927,N_17328,N_17114);
xor U17928 (N_17928,N_17341,N_17119);
nor U17929 (N_17929,N_17111,N_17172);
xor U17930 (N_17930,N_16824,N_17191);
and U17931 (N_17931,N_17306,N_17007);
nand U17932 (N_17932,N_16824,N_17270);
xnor U17933 (N_17933,N_17280,N_17307);
nand U17934 (N_17934,N_16923,N_16978);
and U17935 (N_17935,N_17202,N_17343);
nand U17936 (N_17936,N_17209,N_16910);
nor U17937 (N_17937,N_17053,N_17329);
or U17938 (N_17938,N_17181,N_17301);
nand U17939 (N_17939,N_17055,N_16800);
or U17940 (N_17940,N_16859,N_16952);
or U17941 (N_17941,N_16831,N_17191);
and U17942 (N_17942,N_17320,N_16884);
nor U17943 (N_17943,N_16858,N_17399);
nor U17944 (N_17944,N_16942,N_17387);
or U17945 (N_17945,N_17242,N_16889);
nand U17946 (N_17946,N_17160,N_17072);
xnor U17947 (N_17947,N_17060,N_17373);
and U17948 (N_17948,N_17107,N_16855);
or U17949 (N_17949,N_16906,N_17124);
and U17950 (N_17950,N_17021,N_16904);
nand U17951 (N_17951,N_16815,N_17334);
nor U17952 (N_17952,N_17050,N_17356);
and U17953 (N_17953,N_17226,N_17260);
nand U17954 (N_17954,N_16803,N_17365);
nand U17955 (N_17955,N_17353,N_17118);
nand U17956 (N_17956,N_17214,N_17063);
nor U17957 (N_17957,N_17034,N_16898);
nor U17958 (N_17958,N_17134,N_17279);
and U17959 (N_17959,N_17030,N_16875);
nor U17960 (N_17960,N_16980,N_16964);
or U17961 (N_17961,N_17368,N_17362);
nand U17962 (N_17962,N_17318,N_17235);
xor U17963 (N_17963,N_16938,N_17348);
or U17964 (N_17964,N_17076,N_16949);
nor U17965 (N_17965,N_16828,N_17018);
or U17966 (N_17966,N_17157,N_17302);
nand U17967 (N_17967,N_17105,N_17283);
nor U17968 (N_17968,N_17088,N_17227);
nor U17969 (N_17969,N_17063,N_16956);
nand U17970 (N_17970,N_16809,N_17037);
xnor U17971 (N_17971,N_16865,N_17081);
xnor U17972 (N_17972,N_17042,N_16801);
nand U17973 (N_17973,N_17186,N_17346);
or U17974 (N_17974,N_17284,N_17087);
nor U17975 (N_17975,N_17104,N_17110);
and U17976 (N_17976,N_17268,N_17099);
and U17977 (N_17977,N_16982,N_16972);
nand U17978 (N_17978,N_17207,N_17263);
and U17979 (N_17979,N_17247,N_17078);
nand U17980 (N_17980,N_17142,N_17201);
or U17981 (N_17981,N_17326,N_17153);
nand U17982 (N_17982,N_17255,N_16968);
and U17983 (N_17983,N_17101,N_17125);
nand U17984 (N_17984,N_16899,N_16915);
nor U17985 (N_17985,N_16811,N_17396);
and U17986 (N_17986,N_17124,N_17212);
nand U17987 (N_17987,N_17006,N_17247);
nand U17988 (N_17988,N_17150,N_17016);
nor U17989 (N_17989,N_16874,N_17140);
and U17990 (N_17990,N_17099,N_16842);
nor U17991 (N_17991,N_17277,N_17008);
nand U17992 (N_17992,N_17311,N_16865);
nand U17993 (N_17993,N_16877,N_17284);
nand U17994 (N_17994,N_16971,N_17351);
nor U17995 (N_17995,N_16916,N_17192);
xnor U17996 (N_17996,N_16999,N_17199);
nand U17997 (N_17997,N_17306,N_17038);
and U17998 (N_17998,N_16873,N_16970);
nand U17999 (N_17999,N_17290,N_16939);
and U18000 (N_18000,N_17404,N_17438);
or U18001 (N_18001,N_17844,N_17929);
and U18002 (N_18002,N_17612,N_17780);
nor U18003 (N_18003,N_17681,N_17426);
and U18004 (N_18004,N_17430,N_17492);
nor U18005 (N_18005,N_17572,N_17767);
or U18006 (N_18006,N_17688,N_17893);
or U18007 (N_18007,N_17978,N_17656);
nor U18008 (N_18008,N_17673,N_17470);
nand U18009 (N_18009,N_17574,N_17678);
and U18010 (N_18010,N_17568,N_17933);
and U18011 (N_18011,N_17659,N_17799);
nor U18012 (N_18012,N_17861,N_17848);
or U18013 (N_18013,N_17997,N_17468);
or U18014 (N_18014,N_17887,N_17976);
or U18015 (N_18015,N_17850,N_17503);
nand U18016 (N_18016,N_17635,N_17880);
nor U18017 (N_18017,N_17734,N_17723);
nand U18018 (N_18018,N_17616,N_17421);
nor U18019 (N_18019,N_17499,N_17602);
and U18020 (N_18020,N_17807,N_17951);
nor U18021 (N_18021,N_17631,N_17630);
or U18022 (N_18022,N_17483,N_17842);
nand U18023 (N_18023,N_17736,N_17774);
and U18024 (N_18024,N_17541,N_17755);
nand U18025 (N_18025,N_17625,N_17790);
xnor U18026 (N_18026,N_17607,N_17984);
and U18027 (N_18027,N_17511,N_17706);
nand U18028 (N_18028,N_17588,N_17944);
nand U18029 (N_18029,N_17999,N_17741);
nor U18030 (N_18030,N_17765,N_17453);
nand U18031 (N_18031,N_17493,N_17866);
nand U18032 (N_18032,N_17760,N_17838);
nand U18033 (N_18033,N_17731,N_17578);
and U18034 (N_18034,N_17583,N_17895);
nor U18035 (N_18035,N_17879,N_17983);
xnor U18036 (N_18036,N_17431,N_17650);
nand U18037 (N_18037,N_17764,N_17486);
nor U18038 (N_18038,N_17686,N_17539);
and U18039 (N_18039,N_17657,N_17894);
nand U18040 (N_18040,N_17559,N_17520);
and U18041 (N_18041,N_17835,N_17752);
nand U18042 (N_18042,N_17803,N_17993);
nand U18043 (N_18043,N_17950,N_17740);
and U18044 (N_18044,N_17669,N_17905);
nor U18045 (N_18045,N_17963,N_17698);
and U18046 (N_18046,N_17676,N_17967);
xnor U18047 (N_18047,N_17833,N_17919);
and U18048 (N_18048,N_17600,N_17476);
or U18049 (N_18049,N_17674,N_17604);
and U18050 (N_18050,N_17550,N_17447);
nand U18051 (N_18051,N_17609,N_17808);
and U18052 (N_18052,N_17981,N_17622);
nor U18053 (N_18053,N_17451,N_17713);
and U18054 (N_18054,N_17407,N_17987);
nand U18055 (N_18055,N_17529,N_17990);
nand U18056 (N_18056,N_17694,N_17813);
nand U18057 (N_18057,N_17584,N_17491);
or U18058 (N_18058,N_17834,N_17974);
and U18059 (N_18059,N_17965,N_17642);
or U18060 (N_18060,N_17514,N_17562);
nand U18061 (N_18061,N_17467,N_17535);
or U18062 (N_18062,N_17563,N_17544);
and U18063 (N_18063,N_17881,N_17860);
nand U18064 (N_18064,N_17943,N_17537);
or U18065 (N_18065,N_17435,N_17524);
nor U18066 (N_18066,N_17518,N_17434);
or U18067 (N_18067,N_17582,N_17662);
nand U18068 (N_18068,N_17772,N_17968);
nor U18069 (N_18069,N_17739,N_17641);
xnor U18070 (N_18070,N_17816,N_17667);
or U18071 (N_18071,N_17809,N_17849);
or U18072 (N_18072,N_17909,N_17664);
and U18073 (N_18073,N_17819,N_17906);
nand U18074 (N_18074,N_17708,N_17536);
or U18075 (N_18075,N_17721,N_17413);
or U18076 (N_18076,N_17558,N_17403);
and U18077 (N_18077,N_17423,N_17654);
and U18078 (N_18078,N_17644,N_17684);
and U18079 (N_18079,N_17628,N_17753);
nor U18080 (N_18080,N_17865,N_17414);
nor U18081 (N_18081,N_17570,N_17437);
and U18082 (N_18082,N_17627,N_17802);
nor U18083 (N_18083,N_17953,N_17454);
xnor U18084 (N_18084,N_17872,N_17797);
and U18085 (N_18085,N_17979,N_17610);
or U18086 (N_18086,N_17846,N_17488);
or U18087 (N_18087,N_17552,N_17847);
and U18088 (N_18088,N_17497,N_17419);
nor U18089 (N_18089,N_17590,N_17702);
and U18090 (N_18090,N_17623,N_17459);
and U18091 (N_18091,N_17885,N_17882);
nor U18092 (N_18092,N_17675,N_17720);
nor U18093 (N_18093,N_17946,N_17500);
nand U18094 (N_18094,N_17508,N_17750);
nand U18095 (N_18095,N_17996,N_17862);
and U18096 (N_18096,N_17932,N_17977);
xor U18097 (N_18097,N_17748,N_17672);
or U18098 (N_18098,N_17804,N_17545);
nand U18099 (N_18099,N_17761,N_17576);
and U18100 (N_18100,N_17589,N_17697);
nand U18101 (N_18101,N_17854,N_17652);
or U18102 (N_18102,N_17569,N_17806);
nor U18103 (N_18103,N_17494,N_17766);
or U18104 (N_18104,N_17921,N_17971);
or U18105 (N_18105,N_17988,N_17811);
and U18106 (N_18106,N_17690,N_17712);
nor U18107 (N_18107,N_17472,N_17747);
nor U18108 (N_18108,N_17964,N_17636);
nor U18109 (N_18109,N_17617,N_17548);
and U18110 (N_18110,N_17925,N_17462);
or U18111 (N_18111,N_17902,N_17917);
or U18112 (N_18112,N_17516,N_17782);
or U18113 (N_18113,N_17465,N_17920);
nor U18114 (N_18114,N_17605,N_17888);
nor U18115 (N_18115,N_17626,N_17892);
and U18116 (N_18116,N_17638,N_17859);
or U18117 (N_18117,N_17471,N_17639);
nand U18118 (N_18118,N_17540,N_17954);
or U18119 (N_18119,N_17863,N_17601);
or U18120 (N_18120,N_17982,N_17480);
nor U18121 (N_18121,N_17441,N_17818);
and U18122 (N_18122,N_17903,N_17598);
nor U18123 (N_18123,N_17969,N_17824);
or U18124 (N_18124,N_17526,N_17770);
and U18125 (N_18125,N_17512,N_17611);
nor U18126 (N_18126,N_17689,N_17519);
nand U18127 (N_18127,N_17776,N_17670);
nor U18128 (N_18128,N_17826,N_17428);
or U18129 (N_18129,N_17904,N_17629);
nor U18130 (N_18130,N_17821,N_17406);
or U18131 (N_18131,N_17416,N_17707);
and U18132 (N_18132,N_17754,N_17561);
nand U18133 (N_18133,N_17915,N_17883);
and U18134 (N_18134,N_17949,N_17411);
nand U18135 (N_18135,N_17495,N_17710);
and U18136 (N_18136,N_17528,N_17763);
nand U18137 (N_18137,N_17691,N_17485);
or U18138 (N_18138,N_17432,N_17730);
or U18139 (N_18139,N_17719,N_17700);
xor U18140 (N_18140,N_17703,N_17778);
and U18141 (N_18141,N_17533,N_17936);
nand U18142 (N_18142,N_17901,N_17693);
nor U18143 (N_18143,N_17448,N_17487);
and U18144 (N_18144,N_17972,N_17900);
and U18145 (N_18145,N_17685,N_17651);
and U18146 (N_18146,N_17787,N_17573);
and U18147 (N_18147,N_17958,N_17556);
nor U18148 (N_18148,N_17458,N_17655);
xnor U18149 (N_18149,N_17597,N_17409);
nand U18150 (N_18150,N_17908,N_17449);
nor U18151 (N_18151,N_17417,N_17425);
and U18152 (N_18152,N_17554,N_17940);
nand U18153 (N_18153,N_17724,N_17939);
nand U18154 (N_18154,N_17852,N_17839);
nand U18155 (N_18155,N_17444,N_17564);
nand U18156 (N_18156,N_17658,N_17907);
and U18157 (N_18157,N_17624,N_17640);
nor U18158 (N_18158,N_17986,N_17768);
or U18159 (N_18159,N_17412,N_17832);
and U18160 (N_18160,N_17837,N_17677);
nand U18161 (N_18161,N_17913,N_17699);
or U18162 (N_18162,N_17942,N_17975);
and U18163 (N_18163,N_17531,N_17567);
or U18164 (N_18164,N_17911,N_17575);
and U18165 (N_18165,N_17725,N_17711);
or U18166 (N_18166,N_17473,N_17898);
nand U18167 (N_18167,N_17542,N_17445);
nor U18168 (N_18168,N_17599,N_17851);
xnor U18169 (N_18169,N_17566,N_17751);
and U18170 (N_18170,N_17402,N_17783);
or U18171 (N_18171,N_17794,N_17941);
nand U18172 (N_18172,N_17771,N_17443);
or U18173 (N_18173,N_17796,N_17424);
and U18174 (N_18174,N_17515,N_17934);
and U18175 (N_18175,N_17916,N_17952);
and U18176 (N_18176,N_17716,N_17727);
nor U18177 (N_18177,N_17595,N_17948);
xor U18178 (N_18178,N_17891,N_17498);
and U18179 (N_18179,N_17709,N_17504);
or U18180 (N_18180,N_17820,N_17618);
nor U18181 (N_18181,N_17433,N_17692);
and U18182 (N_18182,N_17679,N_17801);
or U18183 (N_18183,N_17665,N_17812);
nand U18184 (N_18184,N_17732,N_17621);
nand U18185 (N_18185,N_17643,N_17991);
or U18186 (N_18186,N_17718,N_17671);
nor U18187 (N_18187,N_17980,N_17758);
nor U18188 (N_18188,N_17745,N_17501);
nor U18189 (N_18189,N_17466,N_17683);
nand U18190 (N_18190,N_17507,N_17634);
xor U18191 (N_18191,N_17505,N_17436);
nand U18192 (N_18192,N_17581,N_17696);
xnor U18193 (N_18193,N_17619,N_17510);
or U18194 (N_18194,N_17653,N_17779);
nor U18195 (N_18195,N_17646,N_17912);
and U18196 (N_18196,N_17935,N_17845);
nand U18197 (N_18197,N_17603,N_17452);
or U18198 (N_18198,N_17795,N_17704);
and U18199 (N_18199,N_17647,N_17857);
and U18200 (N_18200,N_17596,N_17496);
nor U18201 (N_18201,N_17961,N_17439);
nor U18202 (N_18202,N_17868,N_17922);
xor U18203 (N_18203,N_17429,N_17910);
nand U18204 (N_18204,N_17571,N_17926);
nor U18205 (N_18205,N_17632,N_17701);
nor U18206 (N_18206,N_17973,N_17586);
nand U18207 (N_18207,N_17521,N_17405);
nand U18208 (N_18208,N_17717,N_17553);
or U18209 (N_18209,N_17867,N_17746);
or U18210 (N_18210,N_17960,N_17923);
nand U18211 (N_18211,N_17479,N_17956);
nor U18212 (N_18212,N_17890,N_17633);
nand U18213 (N_18213,N_17875,N_17549);
nor U18214 (N_18214,N_17793,N_17897);
and U18215 (N_18215,N_17791,N_17843);
nand U18216 (N_18216,N_17775,N_17937);
and U18217 (N_18217,N_17817,N_17557);
or U18218 (N_18218,N_17560,N_17450);
nand U18219 (N_18219,N_17827,N_17660);
nand U18220 (N_18220,N_17995,N_17858);
or U18221 (N_18221,N_17749,N_17482);
and U18222 (N_18222,N_17864,N_17726);
nand U18223 (N_18223,N_17785,N_17959);
nor U18224 (N_18224,N_17970,N_17856);
xnor U18225 (N_18225,N_17615,N_17648);
nand U18226 (N_18226,N_17580,N_17876);
nand U18227 (N_18227,N_17446,N_17884);
nor U18228 (N_18228,N_17608,N_17733);
nor U18229 (N_18229,N_17469,N_17989);
nand U18230 (N_18230,N_17715,N_17786);
and U18231 (N_18231,N_17440,N_17506);
nor U18232 (N_18232,N_17455,N_17889);
or U18233 (N_18233,N_17415,N_17481);
xnor U18234 (N_18234,N_17687,N_17509);
or U18235 (N_18235,N_17728,N_17757);
and U18236 (N_18236,N_17614,N_17877);
or U18237 (N_18237,N_17896,N_17798);
nor U18238 (N_18238,N_17637,N_17871);
or U18239 (N_18239,N_17695,N_17792);
nor U18240 (N_18240,N_17538,N_17408);
nand U18241 (N_18241,N_17743,N_17773);
nand U18242 (N_18242,N_17682,N_17928);
nand U18243 (N_18243,N_17855,N_17853);
nand U18244 (N_18244,N_17442,N_17502);
nand U18245 (N_18245,N_17661,N_17729);
or U18246 (N_18246,N_17594,N_17680);
nand U18247 (N_18247,N_17593,N_17525);
or U18248 (N_18248,N_17985,N_17577);
or U18249 (N_18249,N_17522,N_17784);
nor U18250 (N_18250,N_17955,N_17777);
and U18251 (N_18251,N_17869,N_17555);
nor U18252 (N_18252,N_17463,N_17489);
and U18253 (N_18253,N_17886,N_17828);
and U18254 (N_18254,N_17401,N_17873);
and U18255 (N_18255,N_17924,N_17927);
nand U18256 (N_18256,N_17478,N_17938);
and U18257 (N_18257,N_17464,N_17810);
xor U18258 (N_18258,N_17705,N_17918);
xnor U18259 (N_18259,N_17962,N_17878);
xnor U18260 (N_18260,N_17815,N_17418);
nand U18261 (N_18261,N_17668,N_17585);
and U18262 (N_18262,N_17649,N_17874);
nor U18263 (N_18263,N_17735,N_17756);
nand U18264 (N_18264,N_17822,N_17742);
nor U18265 (N_18265,N_17998,N_17532);
or U18266 (N_18266,N_17587,N_17714);
and U18267 (N_18267,N_17759,N_17899);
xor U18268 (N_18268,N_17841,N_17613);
or U18269 (N_18269,N_17456,N_17477);
or U18270 (N_18270,N_17543,N_17781);
nand U18271 (N_18271,N_17484,N_17966);
and U18272 (N_18272,N_17475,N_17722);
xnor U18273 (N_18273,N_17825,N_17840);
or U18274 (N_18274,N_17546,N_17461);
or U18275 (N_18275,N_17579,N_17565);
nor U18276 (N_18276,N_17737,N_17870);
nor U18277 (N_18277,N_17744,N_17947);
nand U18278 (N_18278,N_17513,N_17823);
or U18279 (N_18279,N_17591,N_17534);
and U18280 (N_18280,N_17547,N_17836);
and U18281 (N_18281,N_17994,N_17620);
and U18282 (N_18282,N_17830,N_17645);
and U18283 (N_18283,N_17769,N_17490);
and U18284 (N_18284,N_17788,N_17931);
or U18285 (N_18285,N_17422,N_17814);
and U18286 (N_18286,N_17789,N_17663);
and U18287 (N_18287,N_17831,N_17606);
xnor U18288 (N_18288,N_17460,N_17762);
and U18289 (N_18289,N_17829,N_17457);
and U18290 (N_18290,N_17592,N_17474);
xor U18291 (N_18291,N_17945,N_17805);
and U18292 (N_18292,N_17800,N_17400);
and U18293 (N_18293,N_17738,N_17957);
xor U18294 (N_18294,N_17523,N_17427);
nand U18295 (N_18295,N_17930,N_17666);
nand U18296 (N_18296,N_17420,N_17410);
or U18297 (N_18297,N_17527,N_17530);
or U18298 (N_18298,N_17517,N_17914);
nor U18299 (N_18299,N_17551,N_17992);
nor U18300 (N_18300,N_17810,N_17457);
nand U18301 (N_18301,N_17897,N_17750);
and U18302 (N_18302,N_17410,N_17820);
and U18303 (N_18303,N_17903,N_17837);
xnor U18304 (N_18304,N_17901,N_17756);
xor U18305 (N_18305,N_17794,N_17428);
nor U18306 (N_18306,N_17713,N_17681);
and U18307 (N_18307,N_17447,N_17697);
nand U18308 (N_18308,N_17860,N_17609);
and U18309 (N_18309,N_17999,N_17882);
nor U18310 (N_18310,N_17741,N_17501);
nand U18311 (N_18311,N_17802,N_17529);
nor U18312 (N_18312,N_17640,N_17580);
nor U18313 (N_18313,N_17481,N_17533);
and U18314 (N_18314,N_17969,N_17415);
and U18315 (N_18315,N_17781,N_17839);
and U18316 (N_18316,N_17596,N_17519);
xor U18317 (N_18317,N_17907,N_17835);
xnor U18318 (N_18318,N_17930,N_17691);
and U18319 (N_18319,N_17846,N_17509);
nand U18320 (N_18320,N_17589,N_17976);
and U18321 (N_18321,N_17972,N_17448);
nand U18322 (N_18322,N_17820,N_17964);
xor U18323 (N_18323,N_17656,N_17555);
xnor U18324 (N_18324,N_17854,N_17498);
nor U18325 (N_18325,N_17822,N_17506);
and U18326 (N_18326,N_17821,N_17717);
nand U18327 (N_18327,N_17775,N_17664);
and U18328 (N_18328,N_17730,N_17870);
nand U18329 (N_18329,N_17624,N_17723);
and U18330 (N_18330,N_17771,N_17794);
nor U18331 (N_18331,N_17952,N_17938);
and U18332 (N_18332,N_17782,N_17841);
or U18333 (N_18333,N_17787,N_17792);
and U18334 (N_18334,N_17581,N_17562);
nand U18335 (N_18335,N_17680,N_17924);
and U18336 (N_18336,N_17671,N_17888);
or U18337 (N_18337,N_17621,N_17632);
or U18338 (N_18338,N_17656,N_17658);
or U18339 (N_18339,N_17845,N_17766);
and U18340 (N_18340,N_17739,N_17899);
nand U18341 (N_18341,N_17427,N_17987);
or U18342 (N_18342,N_17781,N_17442);
nor U18343 (N_18343,N_17459,N_17711);
xnor U18344 (N_18344,N_17902,N_17594);
nand U18345 (N_18345,N_17521,N_17951);
and U18346 (N_18346,N_17796,N_17488);
and U18347 (N_18347,N_17784,N_17593);
nor U18348 (N_18348,N_17546,N_17904);
and U18349 (N_18349,N_17489,N_17993);
xnor U18350 (N_18350,N_17815,N_17989);
xnor U18351 (N_18351,N_17493,N_17706);
nand U18352 (N_18352,N_17775,N_17912);
or U18353 (N_18353,N_17408,N_17687);
nand U18354 (N_18354,N_17627,N_17861);
or U18355 (N_18355,N_17818,N_17683);
nor U18356 (N_18356,N_17856,N_17471);
and U18357 (N_18357,N_17984,N_17941);
and U18358 (N_18358,N_17878,N_17581);
nor U18359 (N_18359,N_17891,N_17851);
nor U18360 (N_18360,N_17479,N_17609);
or U18361 (N_18361,N_17918,N_17665);
and U18362 (N_18362,N_17700,N_17804);
nand U18363 (N_18363,N_17738,N_17416);
nand U18364 (N_18364,N_17781,N_17986);
nand U18365 (N_18365,N_17422,N_17636);
and U18366 (N_18366,N_17650,N_17777);
and U18367 (N_18367,N_17832,N_17515);
nand U18368 (N_18368,N_17532,N_17505);
nand U18369 (N_18369,N_17814,N_17654);
or U18370 (N_18370,N_17481,N_17899);
nor U18371 (N_18371,N_17633,N_17895);
or U18372 (N_18372,N_17522,N_17633);
nand U18373 (N_18373,N_17668,N_17968);
nor U18374 (N_18374,N_17773,N_17708);
or U18375 (N_18375,N_17558,N_17492);
or U18376 (N_18376,N_17838,N_17857);
or U18377 (N_18377,N_17461,N_17869);
and U18378 (N_18378,N_17528,N_17680);
nand U18379 (N_18379,N_17760,N_17951);
nor U18380 (N_18380,N_17747,N_17965);
and U18381 (N_18381,N_17900,N_17422);
nand U18382 (N_18382,N_17483,N_17551);
nor U18383 (N_18383,N_17656,N_17815);
nand U18384 (N_18384,N_17898,N_17584);
or U18385 (N_18385,N_17775,N_17923);
nor U18386 (N_18386,N_17838,N_17879);
nor U18387 (N_18387,N_17815,N_17955);
nand U18388 (N_18388,N_17790,N_17597);
and U18389 (N_18389,N_17813,N_17443);
or U18390 (N_18390,N_17420,N_17403);
nor U18391 (N_18391,N_17519,N_17549);
nor U18392 (N_18392,N_17723,N_17531);
nand U18393 (N_18393,N_17706,N_17859);
nor U18394 (N_18394,N_17752,N_17715);
xnor U18395 (N_18395,N_17767,N_17977);
xnor U18396 (N_18396,N_17802,N_17461);
or U18397 (N_18397,N_17814,N_17495);
nand U18398 (N_18398,N_17959,N_17483);
and U18399 (N_18399,N_17788,N_17837);
nor U18400 (N_18400,N_17419,N_17624);
or U18401 (N_18401,N_17570,N_17543);
nand U18402 (N_18402,N_17859,N_17544);
or U18403 (N_18403,N_17985,N_17676);
nand U18404 (N_18404,N_17475,N_17761);
nor U18405 (N_18405,N_17513,N_17741);
and U18406 (N_18406,N_17548,N_17796);
nor U18407 (N_18407,N_17597,N_17910);
nor U18408 (N_18408,N_17523,N_17706);
xor U18409 (N_18409,N_17907,N_17503);
nor U18410 (N_18410,N_17870,N_17679);
xor U18411 (N_18411,N_17803,N_17730);
nand U18412 (N_18412,N_17872,N_17770);
nand U18413 (N_18413,N_17961,N_17726);
nand U18414 (N_18414,N_17531,N_17681);
nor U18415 (N_18415,N_17493,N_17778);
nor U18416 (N_18416,N_17641,N_17501);
xnor U18417 (N_18417,N_17762,N_17403);
nand U18418 (N_18418,N_17989,N_17838);
and U18419 (N_18419,N_17567,N_17783);
nor U18420 (N_18420,N_17923,N_17593);
and U18421 (N_18421,N_17825,N_17732);
nor U18422 (N_18422,N_17548,N_17851);
or U18423 (N_18423,N_17829,N_17707);
and U18424 (N_18424,N_17678,N_17724);
nand U18425 (N_18425,N_17787,N_17774);
nor U18426 (N_18426,N_17505,N_17846);
and U18427 (N_18427,N_17848,N_17452);
or U18428 (N_18428,N_17773,N_17559);
nor U18429 (N_18429,N_17887,N_17587);
or U18430 (N_18430,N_17660,N_17529);
or U18431 (N_18431,N_17616,N_17818);
xnor U18432 (N_18432,N_17550,N_17544);
and U18433 (N_18433,N_17535,N_17976);
xnor U18434 (N_18434,N_17470,N_17704);
nand U18435 (N_18435,N_17456,N_17661);
and U18436 (N_18436,N_17809,N_17798);
or U18437 (N_18437,N_17771,N_17870);
nor U18438 (N_18438,N_17467,N_17683);
and U18439 (N_18439,N_17531,N_17652);
nor U18440 (N_18440,N_17524,N_17527);
or U18441 (N_18441,N_17609,N_17981);
nor U18442 (N_18442,N_17833,N_17893);
nor U18443 (N_18443,N_17510,N_17960);
xnor U18444 (N_18444,N_17772,N_17444);
or U18445 (N_18445,N_17973,N_17805);
and U18446 (N_18446,N_17565,N_17526);
and U18447 (N_18447,N_17535,N_17711);
or U18448 (N_18448,N_17421,N_17913);
xnor U18449 (N_18449,N_17745,N_17982);
or U18450 (N_18450,N_17570,N_17518);
nor U18451 (N_18451,N_17501,N_17889);
nand U18452 (N_18452,N_17534,N_17832);
nor U18453 (N_18453,N_17866,N_17978);
nand U18454 (N_18454,N_17879,N_17918);
nor U18455 (N_18455,N_17647,N_17904);
nand U18456 (N_18456,N_17800,N_17984);
or U18457 (N_18457,N_17962,N_17776);
or U18458 (N_18458,N_17695,N_17766);
or U18459 (N_18459,N_17694,N_17651);
or U18460 (N_18460,N_17415,N_17869);
and U18461 (N_18461,N_17404,N_17474);
xnor U18462 (N_18462,N_17802,N_17692);
and U18463 (N_18463,N_17842,N_17563);
or U18464 (N_18464,N_17537,N_17944);
xnor U18465 (N_18465,N_17616,N_17725);
and U18466 (N_18466,N_17502,N_17913);
nor U18467 (N_18467,N_17812,N_17988);
nor U18468 (N_18468,N_17742,N_17554);
or U18469 (N_18469,N_17647,N_17739);
or U18470 (N_18470,N_17631,N_17848);
xor U18471 (N_18471,N_17607,N_17510);
nor U18472 (N_18472,N_17436,N_17774);
nand U18473 (N_18473,N_17545,N_17585);
xnor U18474 (N_18474,N_17545,N_17664);
nor U18475 (N_18475,N_17558,N_17797);
and U18476 (N_18476,N_17425,N_17492);
nand U18477 (N_18477,N_17651,N_17797);
xor U18478 (N_18478,N_17812,N_17858);
and U18479 (N_18479,N_17677,N_17511);
nand U18480 (N_18480,N_17847,N_17771);
and U18481 (N_18481,N_17466,N_17716);
and U18482 (N_18482,N_17923,N_17581);
nand U18483 (N_18483,N_17665,N_17816);
nand U18484 (N_18484,N_17801,N_17847);
nand U18485 (N_18485,N_17503,N_17672);
nor U18486 (N_18486,N_17528,N_17571);
and U18487 (N_18487,N_17934,N_17535);
nor U18488 (N_18488,N_17780,N_17569);
nand U18489 (N_18489,N_17946,N_17916);
or U18490 (N_18490,N_17669,N_17524);
and U18491 (N_18491,N_17998,N_17410);
or U18492 (N_18492,N_17869,N_17545);
or U18493 (N_18493,N_17904,N_17954);
and U18494 (N_18494,N_17956,N_17933);
nand U18495 (N_18495,N_17758,N_17983);
xor U18496 (N_18496,N_17430,N_17964);
nand U18497 (N_18497,N_17491,N_17986);
and U18498 (N_18498,N_17548,N_17599);
and U18499 (N_18499,N_17475,N_17492);
nor U18500 (N_18500,N_17501,N_17448);
or U18501 (N_18501,N_17996,N_17919);
xnor U18502 (N_18502,N_17884,N_17887);
or U18503 (N_18503,N_17690,N_17583);
and U18504 (N_18504,N_17805,N_17578);
or U18505 (N_18505,N_17405,N_17801);
nand U18506 (N_18506,N_17462,N_17800);
and U18507 (N_18507,N_17679,N_17840);
nor U18508 (N_18508,N_17968,N_17530);
or U18509 (N_18509,N_17710,N_17990);
or U18510 (N_18510,N_17878,N_17965);
nand U18511 (N_18511,N_17566,N_17821);
nand U18512 (N_18512,N_17681,N_17686);
and U18513 (N_18513,N_17614,N_17983);
or U18514 (N_18514,N_17691,N_17539);
xor U18515 (N_18515,N_17975,N_17936);
xor U18516 (N_18516,N_17716,N_17828);
nand U18517 (N_18517,N_17684,N_17588);
nand U18518 (N_18518,N_17694,N_17796);
nand U18519 (N_18519,N_17774,N_17858);
xor U18520 (N_18520,N_17519,N_17501);
xnor U18521 (N_18521,N_17672,N_17415);
nor U18522 (N_18522,N_17496,N_17520);
nand U18523 (N_18523,N_17817,N_17448);
nor U18524 (N_18524,N_17495,N_17773);
nor U18525 (N_18525,N_17847,N_17930);
nor U18526 (N_18526,N_17962,N_17709);
or U18527 (N_18527,N_17561,N_17910);
nor U18528 (N_18528,N_17690,N_17559);
nand U18529 (N_18529,N_17603,N_17627);
nand U18530 (N_18530,N_17472,N_17710);
nor U18531 (N_18531,N_17723,N_17812);
and U18532 (N_18532,N_17454,N_17828);
and U18533 (N_18533,N_17576,N_17485);
and U18534 (N_18534,N_17595,N_17493);
or U18535 (N_18535,N_17889,N_17719);
or U18536 (N_18536,N_17679,N_17928);
xnor U18537 (N_18537,N_17892,N_17493);
or U18538 (N_18538,N_17635,N_17618);
nand U18539 (N_18539,N_17419,N_17449);
and U18540 (N_18540,N_17831,N_17469);
nand U18541 (N_18541,N_17981,N_17574);
nor U18542 (N_18542,N_17904,N_17948);
nand U18543 (N_18543,N_17629,N_17664);
nand U18544 (N_18544,N_17737,N_17836);
or U18545 (N_18545,N_17796,N_17742);
nand U18546 (N_18546,N_17442,N_17673);
or U18547 (N_18547,N_17477,N_17751);
nand U18548 (N_18548,N_17655,N_17416);
and U18549 (N_18549,N_17658,N_17737);
and U18550 (N_18550,N_17624,N_17920);
and U18551 (N_18551,N_17748,N_17810);
nor U18552 (N_18552,N_17701,N_17826);
and U18553 (N_18553,N_17594,N_17615);
or U18554 (N_18554,N_17954,N_17594);
xor U18555 (N_18555,N_17638,N_17664);
nand U18556 (N_18556,N_17785,N_17980);
nor U18557 (N_18557,N_17965,N_17471);
and U18558 (N_18558,N_17884,N_17464);
and U18559 (N_18559,N_17925,N_17945);
or U18560 (N_18560,N_17521,N_17897);
or U18561 (N_18561,N_17978,N_17853);
and U18562 (N_18562,N_17425,N_17503);
xor U18563 (N_18563,N_17855,N_17506);
or U18564 (N_18564,N_17764,N_17679);
nor U18565 (N_18565,N_17613,N_17492);
and U18566 (N_18566,N_17739,N_17592);
and U18567 (N_18567,N_17742,N_17561);
nor U18568 (N_18568,N_17820,N_17602);
xor U18569 (N_18569,N_17744,N_17713);
or U18570 (N_18570,N_17966,N_17512);
nor U18571 (N_18571,N_17660,N_17733);
or U18572 (N_18572,N_17477,N_17907);
nor U18573 (N_18573,N_17707,N_17413);
nor U18574 (N_18574,N_17992,N_17450);
nand U18575 (N_18575,N_17993,N_17611);
and U18576 (N_18576,N_17865,N_17715);
xnor U18577 (N_18577,N_17685,N_17415);
or U18578 (N_18578,N_17489,N_17945);
xnor U18579 (N_18579,N_17836,N_17846);
xnor U18580 (N_18580,N_17755,N_17603);
or U18581 (N_18581,N_17497,N_17630);
nor U18582 (N_18582,N_17673,N_17406);
and U18583 (N_18583,N_17764,N_17549);
xor U18584 (N_18584,N_17876,N_17802);
and U18585 (N_18585,N_17941,N_17592);
or U18586 (N_18586,N_17875,N_17457);
nor U18587 (N_18587,N_17492,N_17743);
and U18588 (N_18588,N_17933,N_17939);
and U18589 (N_18589,N_17738,N_17989);
nand U18590 (N_18590,N_17776,N_17973);
nand U18591 (N_18591,N_17411,N_17884);
nor U18592 (N_18592,N_17503,N_17542);
and U18593 (N_18593,N_17543,N_17558);
nand U18594 (N_18594,N_17734,N_17401);
nor U18595 (N_18595,N_17895,N_17741);
nand U18596 (N_18596,N_17458,N_17631);
or U18597 (N_18597,N_17896,N_17977);
and U18598 (N_18598,N_17601,N_17864);
nand U18599 (N_18599,N_17832,N_17519);
and U18600 (N_18600,N_18131,N_18372);
nor U18601 (N_18601,N_18179,N_18230);
and U18602 (N_18602,N_18341,N_18461);
or U18603 (N_18603,N_18575,N_18125);
or U18604 (N_18604,N_18497,N_18479);
nand U18605 (N_18605,N_18012,N_18359);
xor U18606 (N_18606,N_18298,N_18543);
and U18607 (N_18607,N_18189,N_18518);
and U18608 (N_18608,N_18314,N_18139);
or U18609 (N_18609,N_18473,N_18019);
and U18610 (N_18610,N_18507,N_18492);
or U18611 (N_18611,N_18467,N_18099);
nand U18612 (N_18612,N_18539,N_18121);
xnor U18613 (N_18613,N_18151,N_18516);
nand U18614 (N_18614,N_18043,N_18077);
nand U18615 (N_18615,N_18385,N_18547);
xnor U18616 (N_18616,N_18297,N_18579);
nor U18617 (N_18617,N_18571,N_18293);
nand U18618 (N_18618,N_18437,N_18347);
or U18619 (N_18619,N_18324,N_18476);
xnor U18620 (N_18620,N_18373,N_18138);
or U18621 (N_18621,N_18219,N_18104);
nor U18622 (N_18622,N_18585,N_18413);
or U18623 (N_18623,N_18350,N_18424);
and U18624 (N_18624,N_18106,N_18134);
and U18625 (N_18625,N_18430,N_18403);
nor U18626 (N_18626,N_18284,N_18107);
and U18627 (N_18627,N_18258,N_18090);
and U18628 (N_18628,N_18025,N_18371);
or U18629 (N_18629,N_18205,N_18378);
and U18630 (N_18630,N_18156,N_18253);
nor U18631 (N_18631,N_18206,N_18029);
nor U18632 (N_18632,N_18448,N_18480);
nor U18633 (N_18633,N_18182,N_18041);
nand U18634 (N_18634,N_18067,N_18436);
nand U18635 (N_18635,N_18320,N_18274);
or U18636 (N_18636,N_18519,N_18277);
nor U18637 (N_18637,N_18429,N_18535);
nand U18638 (N_18638,N_18181,N_18488);
and U18639 (N_18639,N_18425,N_18556);
or U18640 (N_18640,N_18165,N_18392);
nor U18641 (N_18641,N_18559,N_18288);
xor U18642 (N_18642,N_18399,N_18541);
and U18643 (N_18643,N_18015,N_18301);
nand U18644 (N_18644,N_18431,N_18279);
or U18645 (N_18645,N_18587,N_18358);
xor U18646 (N_18646,N_18576,N_18066);
and U18647 (N_18647,N_18318,N_18102);
nand U18648 (N_18648,N_18536,N_18313);
nor U18649 (N_18649,N_18439,N_18051);
nor U18650 (N_18650,N_18552,N_18130);
nand U18651 (N_18651,N_18241,N_18402);
nand U18652 (N_18652,N_18273,N_18335);
nand U18653 (N_18653,N_18417,N_18454);
nor U18654 (N_18654,N_18122,N_18103);
nand U18655 (N_18655,N_18184,N_18081);
and U18656 (N_18656,N_18387,N_18343);
nand U18657 (N_18657,N_18272,N_18033);
and U18658 (N_18658,N_18054,N_18474);
nand U18659 (N_18659,N_18391,N_18554);
and U18660 (N_18660,N_18309,N_18542);
nor U18661 (N_18661,N_18302,N_18079);
nand U18662 (N_18662,N_18491,N_18523);
or U18663 (N_18663,N_18395,N_18545);
and U18664 (N_18664,N_18455,N_18308);
xnor U18665 (N_18665,N_18123,N_18195);
nor U18666 (N_18666,N_18061,N_18060);
and U18667 (N_18667,N_18355,N_18525);
and U18668 (N_18668,N_18404,N_18129);
nand U18669 (N_18669,N_18083,N_18530);
or U18670 (N_18670,N_18349,N_18038);
or U18671 (N_18671,N_18422,N_18572);
nor U18672 (N_18672,N_18558,N_18591);
and U18673 (N_18673,N_18185,N_18319);
nor U18674 (N_18674,N_18146,N_18581);
or U18675 (N_18675,N_18433,N_18194);
nor U18676 (N_18676,N_18231,N_18336);
nand U18677 (N_18677,N_18064,N_18266);
or U18678 (N_18678,N_18311,N_18058);
nor U18679 (N_18679,N_18128,N_18596);
or U18680 (N_18680,N_18237,N_18111);
nor U18681 (N_18681,N_18239,N_18174);
nand U18682 (N_18682,N_18048,N_18057);
nand U18683 (N_18683,N_18026,N_18468);
nand U18684 (N_18684,N_18566,N_18464);
and U18685 (N_18685,N_18487,N_18326);
nor U18686 (N_18686,N_18505,N_18281);
nand U18687 (N_18687,N_18569,N_18268);
and U18688 (N_18688,N_18234,N_18235);
nor U18689 (N_18689,N_18501,N_18290);
or U18690 (N_18690,N_18097,N_18094);
nor U18691 (N_18691,N_18116,N_18504);
or U18692 (N_18692,N_18008,N_18261);
nand U18693 (N_18693,N_18384,N_18285);
nor U18694 (N_18694,N_18549,N_18475);
or U18695 (N_18695,N_18248,N_18332);
or U18696 (N_18696,N_18551,N_18589);
or U18697 (N_18697,N_18289,N_18307);
and U18698 (N_18698,N_18483,N_18257);
and U18699 (N_18699,N_18271,N_18370);
and U18700 (N_18700,N_18380,N_18220);
or U18701 (N_18701,N_18087,N_18527);
nand U18702 (N_18702,N_18137,N_18486);
and U18703 (N_18703,N_18490,N_18023);
nand U18704 (N_18704,N_18457,N_18163);
nand U18705 (N_18705,N_18339,N_18346);
xnor U18706 (N_18706,N_18147,N_18354);
nand U18707 (N_18707,N_18328,N_18100);
xnor U18708 (N_18708,N_18120,N_18440);
nand U18709 (N_18709,N_18331,N_18159);
nor U18710 (N_18710,N_18022,N_18209);
nor U18711 (N_18711,N_18005,N_18187);
xor U18712 (N_18712,N_18095,N_18124);
nand U18713 (N_18713,N_18421,N_18364);
nand U18714 (N_18714,N_18588,N_18191);
xnor U18715 (N_18715,N_18401,N_18397);
and U18716 (N_18716,N_18213,N_18426);
and U18717 (N_18717,N_18306,N_18316);
and U18718 (N_18718,N_18405,N_18250);
nor U18719 (N_18719,N_18072,N_18166);
or U18720 (N_18720,N_18173,N_18118);
or U18721 (N_18721,N_18365,N_18267);
or U18722 (N_18722,N_18126,N_18286);
or U18723 (N_18723,N_18500,N_18442);
or U18724 (N_18724,N_18374,N_18513);
nor U18725 (N_18725,N_18294,N_18478);
or U18726 (N_18726,N_18567,N_18200);
xnor U18727 (N_18727,N_18254,N_18408);
nor U18728 (N_18728,N_18502,N_18410);
and U18729 (N_18729,N_18047,N_18471);
nor U18730 (N_18730,N_18533,N_18445);
nor U18731 (N_18731,N_18484,N_18140);
nor U18732 (N_18732,N_18063,N_18562);
nand U18733 (N_18733,N_18172,N_18056);
nand U18734 (N_18734,N_18030,N_18360);
nand U18735 (N_18735,N_18327,N_18260);
nand U18736 (N_18736,N_18157,N_18546);
xor U18737 (N_18737,N_18199,N_18450);
and U18738 (N_18738,N_18353,N_18197);
xor U18739 (N_18739,N_18003,N_18532);
nand U18740 (N_18740,N_18031,N_18361);
xnor U18741 (N_18741,N_18269,N_18177);
and U18742 (N_18742,N_18561,N_18382);
and U18743 (N_18743,N_18325,N_18245);
nor U18744 (N_18744,N_18007,N_18082);
or U18745 (N_18745,N_18540,N_18210);
nor U18746 (N_18746,N_18334,N_18252);
nor U18747 (N_18747,N_18338,N_18114);
nor U18748 (N_18748,N_18204,N_18428);
nand U18749 (N_18749,N_18086,N_18323);
nand U18750 (N_18750,N_18175,N_18568);
xor U18751 (N_18751,N_18452,N_18078);
nand U18752 (N_18752,N_18158,N_18362);
or U18753 (N_18753,N_18202,N_18228);
nor U18754 (N_18754,N_18409,N_18407);
or U18755 (N_18755,N_18018,N_18014);
xnor U18756 (N_18756,N_18249,N_18183);
nand U18757 (N_18757,N_18553,N_18059);
nand U18758 (N_18758,N_18388,N_18119);
nand U18759 (N_18759,N_18394,N_18435);
and U18760 (N_18760,N_18526,N_18169);
nand U18761 (N_18761,N_18550,N_18162);
or U18762 (N_18762,N_18312,N_18225);
xor U18763 (N_18763,N_18133,N_18141);
and U18764 (N_18764,N_18155,N_18351);
nor U18765 (N_18765,N_18052,N_18053);
nor U18766 (N_18766,N_18510,N_18108);
and U18767 (N_18767,N_18337,N_18506);
nand U18768 (N_18768,N_18367,N_18074);
and U18769 (N_18769,N_18238,N_18201);
nor U18770 (N_18770,N_18389,N_18152);
nand U18771 (N_18771,N_18393,N_18096);
nor U18772 (N_18772,N_18112,N_18348);
or U18773 (N_18773,N_18171,N_18049);
nand U18774 (N_18774,N_18287,N_18570);
nand U18775 (N_18775,N_18154,N_18366);
nor U18776 (N_18776,N_18212,N_18296);
and U18777 (N_18777,N_18071,N_18376);
nand U18778 (N_18778,N_18198,N_18034);
and U18779 (N_18779,N_18075,N_18017);
and U18780 (N_18780,N_18032,N_18040);
nand U18781 (N_18781,N_18098,N_18529);
or U18782 (N_18782,N_18427,N_18406);
and U18783 (N_18783,N_18011,N_18560);
or U18784 (N_18784,N_18275,N_18001);
or U18785 (N_18785,N_18418,N_18584);
and U18786 (N_18786,N_18000,N_18578);
or U18787 (N_18787,N_18565,N_18217);
nand U18788 (N_18788,N_18514,N_18080);
nor U18789 (N_18789,N_18259,N_18292);
nand U18790 (N_18790,N_18363,N_18167);
and U18791 (N_18791,N_18390,N_18160);
or U18792 (N_18792,N_18415,N_18377);
nand U18793 (N_18793,N_18039,N_18042);
nand U18794 (N_18794,N_18224,N_18263);
xnor U18795 (N_18795,N_18511,N_18573);
nand U18796 (N_18796,N_18329,N_18322);
or U18797 (N_18797,N_18356,N_18344);
and U18798 (N_18798,N_18113,N_18414);
nor U18799 (N_18799,N_18145,N_18170);
or U18800 (N_18800,N_18521,N_18396);
nor U18801 (N_18801,N_18044,N_18276);
nand U18802 (N_18802,N_18420,N_18368);
nand U18803 (N_18803,N_18035,N_18024);
and U18804 (N_18804,N_18262,N_18070);
nor U18805 (N_18805,N_18503,N_18548);
or U18806 (N_18806,N_18013,N_18062);
or U18807 (N_18807,N_18465,N_18592);
nand U18808 (N_18808,N_18223,N_18009);
and U18809 (N_18809,N_18161,N_18432);
xor U18810 (N_18810,N_18557,N_18211);
and U18811 (N_18811,N_18528,N_18105);
nor U18812 (N_18812,N_18028,N_18073);
nor U18813 (N_18813,N_18143,N_18564);
nor U18814 (N_18814,N_18463,N_18089);
or U18815 (N_18815,N_18538,N_18317);
or U18816 (N_18816,N_18438,N_18482);
nand U18817 (N_18817,N_18282,N_18188);
nand U18818 (N_18818,N_18381,N_18416);
xor U18819 (N_18819,N_18244,N_18305);
nor U18820 (N_18820,N_18386,N_18330);
or U18821 (N_18821,N_18117,N_18295);
nand U18822 (N_18822,N_18135,N_18577);
nor U18823 (N_18823,N_18423,N_18534);
and U18824 (N_18824,N_18340,N_18150);
nand U18825 (N_18825,N_18522,N_18352);
or U18826 (N_18826,N_18164,N_18006);
and U18827 (N_18827,N_18515,N_18595);
and U18828 (N_18828,N_18069,N_18412);
or U18829 (N_18829,N_18499,N_18509);
and U18830 (N_18830,N_18524,N_18101);
nand U18831 (N_18831,N_18251,N_18027);
or U18832 (N_18832,N_18176,N_18315);
xnor U18833 (N_18833,N_18214,N_18456);
or U18834 (N_18834,N_18419,N_18093);
nand U18835 (N_18835,N_18411,N_18168);
and U18836 (N_18836,N_18180,N_18470);
or U18837 (N_18837,N_18369,N_18531);
and U18838 (N_18838,N_18555,N_18192);
or U18839 (N_18839,N_18495,N_18256);
nor U18840 (N_18840,N_18459,N_18443);
or U18841 (N_18841,N_18481,N_18010);
nand U18842 (N_18842,N_18472,N_18207);
nand U18843 (N_18843,N_18215,N_18283);
nand U18844 (N_18844,N_18597,N_18037);
and U18845 (N_18845,N_18242,N_18398);
and U18846 (N_18846,N_18144,N_18586);
nand U18847 (N_18847,N_18227,N_18084);
nand U18848 (N_18848,N_18441,N_18498);
and U18849 (N_18849,N_18222,N_18593);
nor U18850 (N_18850,N_18280,N_18255);
nor U18851 (N_18851,N_18247,N_18178);
nor U18852 (N_18852,N_18068,N_18446);
and U18853 (N_18853,N_18520,N_18321);
and U18854 (N_18854,N_18091,N_18264);
or U18855 (N_18855,N_18085,N_18512);
nand U18856 (N_18856,N_18537,N_18278);
and U18857 (N_18857,N_18590,N_18132);
or U18858 (N_18858,N_18036,N_18221);
nor U18859 (N_18859,N_18580,N_18208);
nor U18860 (N_18860,N_18046,N_18379);
and U18861 (N_18861,N_18190,N_18115);
and U18862 (N_18862,N_18243,N_18110);
and U18863 (N_18863,N_18299,N_18021);
nand U18864 (N_18864,N_18055,N_18574);
xor U18865 (N_18865,N_18434,N_18583);
nor U18866 (N_18866,N_18216,N_18383);
and U18867 (N_18867,N_18494,N_18196);
and U18868 (N_18868,N_18598,N_18020);
nor U18869 (N_18869,N_18304,N_18270);
or U18870 (N_18870,N_18462,N_18375);
and U18871 (N_18871,N_18203,N_18142);
nor U18872 (N_18872,N_18517,N_18186);
and U18873 (N_18873,N_18002,N_18447);
nor U18874 (N_18874,N_18148,N_18493);
and U18875 (N_18875,N_18016,N_18451);
xor U18876 (N_18876,N_18291,N_18400);
nand U18877 (N_18877,N_18109,N_18127);
and U18878 (N_18878,N_18449,N_18065);
and U18879 (N_18879,N_18149,N_18004);
nand U18880 (N_18880,N_18599,N_18496);
or U18881 (N_18881,N_18303,N_18232);
nand U18882 (N_18882,N_18458,N_18076);
and U18883 (N_18883,N_18582,N_18594);
nand U18884 (N_18884,N_18050,N_18466);
or U18885 (N_18885,N_18246,N_18088);
and U18886 (N_18886,N_18444,N_18460);
xnor U18887 (N_18887,N_18345,N_18226);
nor U18888 (N_18888,N_18544,N_18229);
nor U18889 (N_18889,N_18136,N_18357);
nand U18890 (N_18890,N_18218,N_18333);
nand U18891 (N_18891,N_18193,N_18563);
nand U18892 (N_18892,N_18092,N_18045);
or U18893 (N_18893,N_18310,N_18300);
or U18894 (N_18894,N_18240,N_18485);
nor U18895 (N_18895,N_18236,N_18508);
nor U18896 (N_18896,N_18153,N_18342);
xor U18897 (N_18897,N_18477,N_18453);
nand U18898 (N_18898,N_18469,N_18265);
or U18899 (N_18899,N_18489,N_18233);
nand U18900 (N_18900,N_18374,N_18538);
nor U18901 (N_18901,N_18512,N_18589);
or U18902 (N_18902,N_18597,N_18169);
and U18903 (N_18903,N_18513,N_18019);
nor U18904 (N_18904,N_18108,N_18266);
and U18905 (N_18905,N_18381,N_18119);
nor U18906 (N_18906,N_18061,N_18047);
or U18907 (N_18907,N_18507,N_18554);
nand U18908 (N_18908,N_18196,N_18491);
nand U18909 (N_18909,N_18320,N_18071);
or U18910 (N_18910,N_18449,N_18503);
and U18911 (N_18911,N_18014,N_18107);
nand U18912 (N_18912,N_18442,N_18140);
and U18913 (N_18913,N_18364,N_18580);
and U18914 (N_18914,N_18418,N_18536);
nor U18915 (N_18915,N_18355,N_18469);
and U18916 (N_18916,N_18023,N_18322);
or U18917 (N_18917,N_18113,N_18032);
xor U18918 (N_18918,N_18297,N_18109);
nor U18919 (N_18919,N_18235,N_18282);
nor U18920 (N_18920,N_18171,N_18018);
or U18921 (N_18921,N_18115,N_18161);
xor U18922 (N_18922,N_18233,N_18129);
nand U18923 (N_18923,N_18268,N_18583);
nor U18924 (N_18924,N_18014,N_18097);
nand U18925 (N_18925,N_18410,N_18489);
and U18926 (N_18926,N_18573,N_18380);
nand U18927 (N_18927,N_18374,N_18473);
or U18928 (N_18928,N_18228,N_18454);
and U18929 (N_18929,N_18485,N_18171);
nand U18930 (N_18930,N_18366,N_18147);
nor U18931 (N_18931,N_18502,N_18062);
nor U18932 (N_18932,N_18140,N_18244);
or U18933 (N_18933,N_18438,N_18575);
nand U18934 (N_18934,N_18400,N_18034);
nor U18935 (N_18935,N_18198,N_18014);
and U18936 (N_18936,N_18333,N_18339);
nand U18937 (N_18937,N_18556,N_18132);
and U18938 (N_18938,N_18504,N_18423);
or U18939 (N_18939,N_18383,N_18119);
xor U18940 (N_18940,N_18487,N_18323);
or U18941 (N_18941,N_18429,N_18162);
or U18942 (N_18942,N_18131,N_18117);
or U18943 (N_18943,N_18346,N_18303);
nor U18944 (N_18944,N_18388,N_18205);
or U18945 (N_18945,N_18591,N_18242);
nand U18946 (N_18946,N_18321,N_18006);
nand U18947 (N_18947,N_18119,N_18358);
and U18948 (N_18948,N_18218,N_18146);
or U18949 (N_18949,N_18222,N_18059);
or U18950 (N_18950,N_18014,N_18568);
nand U18951 (N_18951,N_18112,N_18232);
xnor U18952 (N_18952,N_18423,N_18054);
xnor U18953 (N_18953,N_18597,N_18021);
and U18954 (N_18954,N_18087,N_18390);
nor U18955 (N_18955,N_18443,N_18474);
and U18956 (N_18956,N_18255,N_18268);
nand U18957 (N_18957,N_18441,N_18430);
xnor U18958 (N_18958,N_18296,N_18439);
and U18959 (N_18959,N_18255,N_18079);
nor U18960 (N_18960,N_18331,N_18032);
and U18961 (N_18961,N_18175,N_18217);
xor U18962 (N_18962,N_18094,N_18274);
xnor U18963 (N_18963,N_18595,N_18557);
xor U18964 (N_18964,N_18353,N_18062);
nand U18965 (N_18965,N_18170,N_18543);
nand U18966 (N_18966,N_18145,N_18486);
and U18967 (N_18967,N_18187,N_18291);
nand U18968 (N_18968,N_18558,N_18325);
nor U18969 (N_18969,N_18530,N_18557);
or U18970 (N_18970,N_18448,N_18479);
and U18971 (N_18971,N_18038,N_18546);
nor U18972 (N_18972,N_18439,N_18529);
and U18973 (N_18973,N_18010,N_18231);
nor U18974 (N_18974,N_18541,N_18152);
and U18975 (N_18975,N_18130,N_18200);
nand U18976 (N_18976,N_18459,N_18158);
nand U18977 (N_18977,N_18123,N_18067);
and U18978 (N_18978,N_18049,N_18286);
or U18979 (N_18979,N_18017,N_18585);
and U18980 (N_18980,N_18496,N_18432);
nor U18981 (N_18981,N_18488,N_18175);
nand U18982 (N_18982,N_18332,N_18175);
or U18983 (N_18983,N_18036,N_18593);
and U18984 (N_18984,N_18448,N_18275);
or U18985 (N_18985,N_18319,N_18444);
nand U18986 (N_18986,N_18333,N_18009);
or U18987 (N_18987,N_18110,N_18373);
nand U18988 (N_18988,N_18032,N_18189);
nor U18989 (N_18989,N_18013,N_18593);
and U18990 (N_18990,N_18334,N_18158);
or U18991 (N_18991,N_18280,N_18555);
or U18992 (N_18992,N_18038,N_18224);
or U18993 (N_18993,N_18406,N_18182);
and U18994 (N_18994,N_18030,N_18236);
or U18995 (N_18995,N_18108,N_18333);
and U18996 (N_18996,N_18304,N_18235);
nor U18997 (N_18997,N_18203,N_18366);
or U18998 (N_18998,N_18209,N_18566);
nand U18999 (N_18999,N_18388,N_18278);
nor U19000 (N_19000,N_18012,N_18416);
or U19001 (N_19001,N_18127,N_18133);
and U19002 (N_19002,N_18304,N_18237);
xnor U19003 (N_19003,N_18149,N_18226);
nor U19004 (N_19004,N_18208,N_18146);
nor U19005 (N_19005,N_18494,N_18269);
or U19006 (N_19006,N_18196,N_18394);
or U19007 (N_19007,N_18100,N_18213);
nand U19008 (N_19008,N_18144,N_18326);
and U19009 (N_19009,N_18530,N_18421);
nor U19010 (N_19010,N_18190,N_18478);
or U19011 (N_19011,N_18165,N_18434);
or U19012 (N_19012,N_18192,N_18259);
or U19013 (N_19013,N_18234,N_18422);
nand U19014 (N_19014,N_18409,N_18042);
or U19015 (N_19015,N_18281,N_18016);
xor U19016 (N_19016,N_18383,N_18343);
nor U19017 (N_19017,N_18185,N_18454);
nor U19018 (N_19018,N_18478,N_18570);
or U19019 (N_19019,N_18090,N_18348);
nor U19020 (N_19020,N_18026,N_18152);
nor U19021 (N_19021,N_18498,N_18056);
xnor U19022 (N_19022,N_18324,N_18507);
nand U19023 (N_19023,N_18089,N_18383);
or U19024 (N_19024,N_18275,N_18348);
and U19025 (N_19025,N_18489,N_18359);
and U19026 (N_19026,N_18244,N_18397);
or U19027 (N_19027,N_18185,N_18537);
nor U19028 (N_19028,N_18229,N_18211);
and U19029 (N_19029,N_18077,N_18283);
or U19030 (N_19030,N_18261,N_18407);
nand U19031 (N_19031,N_18366,N_18394);
xnor U19032 (N_19032,N_18387,N_18262);
xnor U19033 (N_19033,N_18482,N_18368);
nand U19034 (N_19034,N_18439,N_18512);
nand U19035 (N_19035,N_18498,N_18400);
or U19036 (N_19036,N_18104,N_18026);
and U19037 (N_19037,N_18276,N_18306);
and U19038 (N_19038,N_18053,N_18519);
nand U19039 (N_19039,N_18246,N_18024);
nor U19040 (N_19040,N_18379,N_18529);
nor U19041 (N_19041,N_18578,N_18186);
or U19042 (N_19042,N_18015,N_18044);
and U19043 (N_19043,N_18031,N_18083);
and U19044 (N_19044,N_18200,N_18420);
xor U19045 (N_19045,N_18535,N_18353);
nor U19046 (N_19046,N_18098,N_18433);
or U19047 (N_19047,N_18141,N_18429);
and U19048 (N_19048,N_18247,N_18411);
nor U19049 (N_19049,N_18245,N_18598);
or U19050 (N_19050,N_18028,N_18440);
and U19051 (N_19051,N_18292,N_18487);
nor U19052 (N_19052,N_18471,N_18199);
xor U19053 (N_19053,N_18090,N_18219);
and U19054 (N_19054,N_18372,N_18543);
nand U19055 (N_19055,N_18458,N_18482);
and U19056 (N_19056,N_18522,N_18445);
or U19057 (N_19057,N_18236,N_18567);
and U19058 (N_19058,N_18484,N_18125);
and U19059 (N_19059,N_18293,N_18557);
xor U19060 (N_19060,N_18094,N_18133);
nor U19061 (N_19061,N_18277,N_18189);
nor U19062 (N_19062,N_18533,N_18564);
xor U19063 (N_19063,N_18163,N_18088);
xor U19064 (N_19064,N_18084,N_18085);
nor U19065 (N_19065,N_18386,N_18398);
or U19066 (N_19066,N_18170,N_18093);
and U19067 (N_19067,N_18342,N_18431);
nand U19068 (N_19068,N_18465,N_18455);
nand U19069 (N_19069,N_18492,N_18223);
and U19070 (N_19070,N_18261,N_18333);
nand U19071 (N_19071,N_18247,N_18260);
or U19072 (N_19072,N_18424,N_18363);
nand U19073 (N_19073,N_18187,N_18485);
nor U19074 (N_19074,N_18106,N_18319);
nor U19075 (N_19075,N_18235,N_18548);
and U19076 (N_19076,N_18239,N_18452);
xnor U19077 (N_19077,N_18488,N_18294);
nor U19078 (N_19078,N_18340,N_18524);
nand U19079 (N_19079,N_18553,N_18506);
or U19080 (N_19080,N_18000,N_18554);
or U19081 (N_19081,N_18137,N_18343);
nand U19082 (N_19082,N_18073,N_18096);
nor U19083 (N_19083,N_18017,N_18594);
and U19084 (N_19084,N_18037,N_18235);
nand U19085 (N_19085,N_18238,N_18534);
nand U19086 (N_19086,N_18536,N_18345);
and U19087 (N_19087,N_18454,N_18260);
nand U19088 (N_19088,N_18560,N_18276);
or U19089 (N_19089,N_18442,N_18195);
and U19090 (N_19090,N_18520,N_18273);
nor U19091 (N_19091,N_18192,N_18294);
or U19092 (N_19092,N_18345,N_18544);
or U19093 (N_19093,N_18483,N_18480);
and U19094 (N_19094,N_18251,N_18441);
or U19095 (N_19095,N_18475,N_18224);
xor U19096 (N_19096,N_18148,N_18596);
or U19097 (N_19097,N_18299,N_18011);
nor U19098 (N_19098,N_18230,N_18480);
nand U19099 (N_19099,N_18119,N_18316);
nand U19100 (N_19100,N_18233,N_18338);
and U19101 (N_19101,N_18532,N_18131);
and U19102 (N_19102,N_18476,N_18276);
or U19103 (N_19103,N_18059,N_18195);
nand U19104 (N_19104,N_18138,N_18437);
and U19105 (N_19105,N_18312,N_18045);
and U19106 (N_19106,N_18597,N_18329);
xnor U19107 (N_19107,N_18489,N_18064);
nor U19108 (N_19108,N_18323,N_18382);
or U19109 (N_19109,N_18546,N_18142);
nand U19110 (N_19110,N_18026,N_18064);
nand U19111 (N_19111,N_18250,N_18481);
nand U19112 (N_19112,N_18137,N_18585);
nor U19113 (N_19113,N_18588,N_18125);
or U19114 (N_19114,N_18397,N_18359);
nand U19115 (N_19115,N_18125,N_18422);
xor U19116 (N_19116,N_18325,N_18138);
nor U19117 (N_19117,N_18050,N_18490);
or U19118 (N_19118,N_18105,N_18343);
nor U19119 (N_19119,N_18547,N_18346);
nor U19120 (N_19120,N_18330,N_18526);
xor U19121 (N_19121,N_18246,N_18294);
nor U19122 (N_19122,N_18366,N_18308);
nor U19123 (N_19123,N_18211,N_18580);
xor U19124 (N_19124,N_18044,N_18383);
nor U19125 (N_19125,N_18103,N_18163);
or U19126 (N_19126,N_18059,N_18432);
and U19127 (N_19127,N_18246,N_18032);
or U19128 (N_19128,N_18367,N_18310);
and U19129 (N_19129,N_18133,N_18507);
nand U19130 (N_19130,N_18043,N_18454);
or U19131 (N_19131,N_18444,N_18554);
nor U19132 (N_19132,N_18347,N_18225);
nor U19133 (N_19133,N_18505,N_18337);
or U19134 (N_19134,N_18465,N_18273);
nor U19135 (N_19135,N_18445,N_18291);
nand U19136 (N_19136,N_18075,N_18182);
and U19137 (N_19137,N_18042,N_18024);
and U19138 (N_19138,N_18020,N_18342);
nand U19139 (N_19139,N_18310,N_18368);
nand U19140 (N_19140,N_18083,N_18359);
and U19141 (N_19141,N_18321,N_18575);
or U19142 (N_19142,N_18449,N_18074);
nand U19143 (N_19143,N_18540,N_18255);
or U19144 (N_19144,N_18106,N_18498);
xor U19145 (N_19145,N_18161,N_18194);
nand U19146 (N_19146,N_18411,N_18490);
nand U19147 (N_19147,N_18573,N_18268);
or U19148 (N_19148,N_18426,N_18075);
nand U19149 (N_19149,N_18515,N_18299);
and U19150 (N_19150,N_18257,N_18165);
and U19151 (N_19151,N_18266,N_18122);
nor U19152 (N_19152,N_18222,N_18447);
or U19153 (N_19153,N_18567,N_18178);
nand U19154 (N_19154,N_18450,N_18322);
and U19155 (N_19155,N_18294,N_18465);
or U19156 (N_19156,N_18489,N_18280);
and U19157 (N_19157,N_18256,N_18259);
nor U19158 (N_19158,N_18480,N_18248);
nand U19159 (N_19159,N_18466,N_18532);
nor U19160 (N_19160,N_18094,N_18411);
nand U19161 (N_19161,N_18169,N_18541);
nand U19162 (N_19162,N_18440,N_18297);
nor U19163 (N_19163,N_18230,N_18056);
and U19164 (N_19164,N_18430,N_18211);
or U19165 (N_19165,N_18471,N_18008);
or U19166 (N_19166,N_18347,N_18435);
nand U19167 (N_19167,N_18523,N_18584);
or U19168 (N_19168,N_18579,N_18425);
xnor U19169 (N_19169,N_18448,N_18443);
nor U19170 (N_19170,N_18511,N_18363);
nand U19171 (N_19171,N_18352,N_18519);
nand U19172 (N_19172,N_18284,N_18509);
and U19173 (N_19173,N_18429,N_18554);
nand U19174 (N_19174,N_18355,N_18538);
nor U19175 (N_19175,N_18399,N_18212);
nor U19176 (N_19176,N_18513,N_18323);
nand U19177 (N_19177,N_18002,N_18305);
and U19178 (N_19178,N_18262,N_18084);
nor U19179 (N_19179,N_18322,N_18055);
and U19180 (N_19180,N_18404,N_18055);
nand U19181 (N_19181,N_18187,N_18575);
nand U19182 (N_19182,N_18583,N_18426);
nand U19183 (N_19183,N_18334,N_18389);
nor U19184 (N_19184,N_18228,N_18048);
nor U19185 (N_19185,N_18521,N_18089);
or U19186 (N_19186,N_18513,N_18182);
nand U19187 (N_19187,N_18582,N_18512);
nand U19188 (N_19188,N_18412,N_18302);
nor U19189 (N_19189,N_18412,N_18354);
and U19190 (N_19190,N_18216,N_18104);
and U19191 (N_19191,N_18376,N_18315);
or U19192 (N_19192,N_18254,N_18426);
nand U19193 (N_19193,N_18412,N_18027);
or U19194 (N_19194,N_18527,N_18032);
nor U19195 (N_19195,N_18029,N_18569);
or U19196 (N_19196,N_18468,N_18540);
or U19197 (N_19197,N_18328,N_18115);
and U19198 (N_19198,N_18464,N_18099);
or U19199 (N_19199,N_18132,N_18526);
and U19200 (N_19200,N_19079,N_18980);
nor U19201 (N_19201,N_18947,N_18705);
and U19202 (N_19202,N_18814,N_18925);
or U19203 (N_19203,N_18862,N_18683);
or U19204 (N_19204,N_18630,N_18963);
xnor U19205 (N_19205,N_18620,N_19017);
and U19206 (N_19206,N_19136,N_19052);
nor U19207 (N_19207,N_18791,N_18691);
and U19208 (N_19208,N_18642,N_18832);
nor U19209 (N_19209,N_19139,N_18845);
or U19210 (N_19210,N_18941,N_18917);
xnor U19211 (N_19211,N_18700,N_19120);
nor U19212 (N_19212,N_19169,N_18701);
nand U19213 (N_19213,N_18651,N_18694);
nand U19214 (N_19214,N_18894,N_18776);
and U19215 (N_19215,N_19014,N_18958);
or U19216 (N_19216,N_18680,N_18920);
or U19217 (N_19217,N_18614,N_19173);
or U19218 (N_19218,N_18883,N_19161);
nand U19219 (N_19219,N_19036,N_19135);
nor U19220 (N_19220,N_18924,N_18652);
xor U19221 (N_19221,N_18686,N_18973);
nor U19222 (N_19222,N_18975,N_19033);
or U19223 (N_19223,N_18954,N_18649);
and U19224 (N_19224,N_19064,N_18606);
nand U19225 (N_19225,N_19012,N_18757);
or U19226 (N_19226,N_18794,N_19035);
xnor U19227 (N_19227,N_18644,N_18689);
or U19228 (N_19228,N_19197,N_18626);
and U19229 (N_19229,N_18638,N_18986);
nand U19230 (N_19230,N_18670,N_18887);
or U19231 (N_19231,N_18764,N_18995);
nor U19232 (N_19232,N_19043,N_18840);
and U19233 (N_19233,N_18781,N_18916);
nand U19234 (N_19234,N_19013,N_18628);
or U19235 (N_19235,N_19106,N_19065);
nor U19236 (N_19236,N_18942,N_18714);
or U19237 (N_19237,N_18601,N_19127);
and U19238 (N_19238,N_18682,N_18793);
and U19239 (N_19239,N_19027,N_18868);
xor U19240 (N_19240,N_19148,N_18792);
nor U19241 (N_19241,N_19032,N_19070);
nor U19242 (N_19242,N_19143,N_18658);
nand U19243 (N_19243,N_19011,N_18877);
or U19244 (N_19244,N_19096,N_19095);
and U19245 (N_19245,N_18923,N_19005);
nor U19246 (N_19246,N_19192,N_18822);
nand U19247 (N_19247,N_18910,N_18798);
or U19248 (N_19248,N_18900,N_19111);
or U19249 (N_19249,N_19194,N_19170);
xnor U19250 (N_19250,N_18911,N_18722);
or U19251 (N_19251,N_18835,N_18807);
nor U19252 (N_19252,N_19168,N_18800);
nand U19253 (N_19253,N_18966,N_18931);
or U19254 (N_19254,N_18663,N_18830);
nor U19255 (N_19255,N_18803,N_19023);
xor U19256 (N_19256,N_19056,N_19094);
nand U19257 (N_19257,N_18990,N_18724);
nand U19258 (N_19258,N_19129,N_19091);
and U19259 (N_19259,N_18846,N_19123);
and U19260 (N_19260,N_19188,N_18838);
and U19261 (N_19261,N_18834,N_18801);
or U19262 (N_19262,N_19072,N_19110);
xnor U19263 (N_19263,N_18977,N_19001);
nand U19264 (N_19264,N_18632,N_19089);
nor U19265 (N_19265,N_18640,N_19198);
or U19266 (N_19266,N_18775,N_18677);
and U19267 (N_19267,N_19021,N_18871);
nor U19268 (N_19268,N_18983,N_18841);
xor U19269 (N_19269,N_18988,N_18913);
or U19270 (N_19270,N_18879,N_18981);
nand U19271 (N_19271,N_18602,N_19097);
xnor U19272 (N_19272,N_18656,N_19047);
nand U19273 (N_19273,N_18943,N_18718);
xor U19274 (N_19274,N_18896,N_19116);
and U19275 (N_19275,N_19151,N_18604);
or U19276 (N_19276,N_18654,N_19006);
nand U19277 (N_19277,N_18777,N_19029);
and U19278 (N_19278,N_18839,N_19164);
nor U19279 (N_19279,N_18639,N_19086);
nand U19280 (N_19280,N_19107,N_18789);
and U19281 (N_19281,N_18989,N_18728);
nor U19282 (N_19282,N_19028,N_19051);
nand U19283 (N_19283,N_18637,N_19195);
or U19284 (N_19284,N_18922,N_19025);
nand U19285 (N_19285,N_19121,N_18698);
and U19286 (N_19286,N_18873,N_19158);
nand U19287 (N_19287,N_18813,N_18819);
nor U19288 (N_19288,N_18696,N_18675);
nor U19289 (N_19289,N_18971,N_18874);
nor U19290 (N_19290,N_19142,N_18704);
xnor U19291 (N_19291,N_18809,N_18710);
or U19292 (N_19292,N_19126,N_18880);
and U19293 (N_19293,N_18780,N_19040);
nand U19294 (N_19294,N_18643,N_18876);
nand U19295 (N_19295,N_19069,N_18991);
xor U19296 (N_19296,N_18742,N_18985);
nor U19297 (N_19297,N_19181,N_18771);
or U19298 (N_19298,N_19009,N_18616);
xor U19299 (N_19299,N_18861,N_19048);
and U19300 (N_19300,N_19179,N_18929);
and U19301 (N_19301,N_18851,N_19180);
nor U19302 (N_19302,N_18815,N_18843);
nand U19303 (N_19303,N_18882,N_18812);
nor U19304 (N_19304,N_18859,N_19191);
nor U19305 (N_19305,N_18984,N_18741);
nand U19306 (N_19306,N_19177,N_18892);
nor U19307 (N_19307,N_18946,N_18927);
or U19308 (N_19308,N_19101,N_18994);
and U19309 (N_19309,N_19075,N_19109);
or U19310 (N_19310,N_18674,N_18782);
or U19311 (N_19311,N_18743,N_18816);
nor U19312 (N_19312,N_18831,N_18996);
nor U19313 (N_19313,N_18895,N_18762);
nor U19314 (N_19314,N_18806,N_18901);
or U19315 (N_19315,N_18768,N_19153);
nor U19316 (N_19316,N_19137,N_18865);
and U19317 (N_19317,N_19060,N_18712);
nor U19318 (N_19318,N_18713,N_18703);
and U19319 (N_19319,N_18869,N_18799);
nor U19320 (N_19320,N_18978,N_19030);
nand U19321 (N_19321,N_18657,N_18624);
and U19322 (N_19322,N_18802,N_18863);
and U19323 (N_19323,N_18945,N_18857);
nand U19324 (N_19324,N_19108,N_18884);
nor U19325 (N_19325,N_18804,N_19113);
nor U19326 (N_19326,N_18821,N_18684);
and U19327 (N_19327,N_18660,N_18766);
nor U19328 (N_19328,N_19088,N_18746);
nand U19329 (N_19329,N_19176,N_18908);
or U19330 (N_19330,N_18905,N_18645);
nor U19331 (N_19331,N_18881,N_19103);
nand U19332 (N_19332,N_19077,N_19133);
or U19333 (N_19333,N_18956,N_18957);
and U19334 (N_19334,N_18779,N_18899);
nor U19335 (N_19335,N_18621,N_19000);
and U19336 (N_19336,N_18953,N_19053);
or U19337 (N_19337,N_18933,N_18854);
nor U19338 (N_19338,N_18787,N_19034);
nor U19339 (N_19339,N_18605,N_18661);
nand U19340 (N_19340,N_18750,N_19073);
or U19341 (N_19341,N_18848,N_18875);
xnor U19342 (N_19342,N_18811,N_18730);
and U19343 (N_19343,N_19076,N_18951);
or U19344 (N_19344,N_18810,N_19098);
xnor U19345 (N_19345,N_18999,N_19145);
or U19346 (N_19346,N_18745,N_18940);
and U19347 (N_19347,N_18818,N_18878);
and U19348 (N_19348,N_18790,N_18650);
nand U19349 (N_19349,N_18837,N_19004);
nand U19350 (N_19350,N_18858,N_18955);
or U19351 (N_19351,N_19026,N_19174);
nor U19352 (N_19352,N_19144,N_19132);
nand U19353 (N_19353,N_18627,N_19057);
or U19354 (N_19354,N_18886,N_19157);
and U19355 (N_19355,N_18936,N_18653);
nand U19356 (N_19356,N_19166,N_18736);
nand U19357 (N_19357,N_18753,N_19066);
xor U19358 (N_19358,N_18631,N_19015);
xor U19359 (N_19359,N_18685,N_19182);
and U19360 (N_19360,N_19125,N_18721);
or U19361 (N_19361,N_18968,N_18849);
xnor U19362 (N_19362,N_18890,N_18711);
nor U19363 (N_19363,N_18906,N_18836);
and U19364 (N_19364,N_18824,N_18709);
nand U19365 (N_19365,N_18784,N_18761);
nor U19366 (N_19366,N_19104,N_18754);
or U19367 (N_19367,N_19084,N_19147);
and U19368 (N_19368,N_18921,N_18797);
and U19369 (N_19369,N_18613,N_18949);
and U19370 (N_19370,N_19010,N_19093);
nand U19371 (N_19371,N_19085,N_19124);
or U19372 (N_19372,N_19022,N_19105);
xor U19373 (N_19373,N_19165,N_18786);
nand U19374 (N_19374,N_18679,N_18747);
and U19375 (N_19375,N_19039,N_19037);
nor U19376 (N_19376,N_19187,N_18737);
xor U19377 (N_19377,N_18928,N_18666);
and U19378 (N_19378,N_18636,N_18629);
nand U19379 (N_19379,N_19046,N_18758);
nor U19380 (N_19380,N_18828,N_19141);
or U19381 (N_19381,N_19038,N_18785);
nor U19382 (N_19382,N_19087,N_18646);
or U19383 (N_19383,N_18934,N_19150);
nand U19384 (N_19384,N_18856,N_19059);
or U19385 (N_19385,N_19130,N_18770);
and U19386 (N_19386,N_18778,N_19122);
and U19387 (N_19387,N_19019,N_18706);
or U19388 (N_19388,N_18727,N_19045);
or U19389 (N_19389,N_19190,N_18829);
nor U19390 (N_19390,N_18635,N_19054);
nand U19391 (N_19391,N_19083,N_19131);
xor U19392 (N_19392,N_18805,N_18998);
xnor U19393 (N_19393,N_19063,N_18962);
and U19394 (N_19394,N_18964,N_18618);
nor U19395 (N_19395,N_18982,N_19062);
nor U19396 (N_19396,N_18987,N_18907);
or U19397 (N_19397,N_18938,N_18600);
and U19398 (N_19398,N_18681,N_19186);
or U19399 (N_19399,N_18693,N_19078);
nor U19400 (N_19400,N_18932,N_18668);
nand U19401 (N_19401,N_19146,N_18699);
nor U19402 (N_19402,N_18969,N_18855);
xnor U19403 (N_19403,N_19189,N_19184);
nand U19404 (N_19404,N_18717,N_18853);
xnor U19405 (N_19405,N_18904,N_18808);
and U19406 (N_19406,N_19199,N_18817);
nor U19407 (N_19407,N_18796,N_19074);
or U19408 (N_19408,N_19155,N_18726);
or U19409 (N_19409,N_18950,N_18827);
xor U19410 (N_19410,N_18773,N_18655);
nor U19411 (N_19411,N_19092,N_18847);
or U19412 (N_19412,N_18774,N_19118);
nor U19413 (N_19413,N_19140,N_18669);
and U19414 (N_19414,N_18959,N_18844);
xor U19415 (N_19415,N_19016,N_18708);
and U19416 (N_19416,N_19178,N_18735);
or U19417 (N_19417,N_19050,N_18738);
nor U19418 (N_19418,N_18607,N_18603);
nand U19419 (N_19419,N_18732,N_18972);
nor U19420 (N_19420,N_18944,N_19055);
nor U19421 (N_19421,N_18748,N_19020);
nor U19422 (N_19422,N_18852,N_18976);
and U19423 (N_19423,N_18850,N_18992);
and U19424 (N_19424,N_19172,N_18625);
nand U19425 (N_19425,N_19042,N_19138);
and U19426 (N_19426,N_19090,N_18926);
xnor U19427 (N_19427,N_18667,N_18939);
xor U19428 (N_19428,N_18898,N_18756);
nand U19429 (N_19429,N_19002,N_18885);
or U19430 (N_19430,N_18752,N_19068);
and U19431 (N_19431,N_19080,N_18690);
or U19432 (N_19432,N_18664,N_18731);
nor U19433 (N_19433,N_18997,N_18672);
and U19434 (N_19434,N_18702,N_18914);
or U19435 (N_19435,N_18715,N_18608);
nand U19436 (N_19436,N_19154,N_18609);
or U19437 (N_19437,N_19007,N_18889);
nor U19438 (N_19438,N_18967,N_19058);
nand U19439 (N_19439,N_19159,N_19061);
and U19440 (N_19440,N_18697,N_18930);
nand U19441 (N_19441,N_19156,N_18867);
or U19442 (N_19442,N_18842,N_18695);
and U19443 (N_19443,N_18872,N_19152);
and U19444 (N_19444,N_19163,N_19003);
nor U19445 (N_19445,N_18622,N_18734);
or U19446 (N_19446,N_18909,N_18870);
or U19447 (N_19447,N_19183,N_18974);
and U19448 (N_19448,N_18719,N_19100);
nor U19449 (N_19449,N_18633,N_19024);
nand U19450 (N_19450,N_18788,N_19102);
xnor U19451 (N_19451,N_18749,N_19117);
and U19452 (N_19452,N_19081,N_19162);
nand U19453 (N_19453,N_18733,N_19175);
and U19454 (N_19454,N_18615,N_18634);
and U19455 (N_19455,N_18820,N_19115);
nand U19456 (N_19456,N_18970,N_19134);
and U19457 (N_19457,N_18769,N_18965);
nand U19458 (N_19458,N_19193,N_18759);
nand U19459 (N_19459,N_18648,N_19082);
and U19460 (N_19460,N_19167,N_18888);
or U19461 (N_19461,N_18723,N_19041);
and U19462 (N_19462,N_18961,N_19044);
and U19463 (N_19463,N_18952,N_18897);
and U19464 (N_19464,N_18617,N_18866);
nand U19465 (N_19465,N_19149,N_18716);
nand U19466 (N_19466,N_18767,N_18915);
and U19467 (N_19467,N_18893,N_19160);
nor U19468 (N_19468,N_18948,N_19185);
nor U19469 (N_19469,N_18765,N_18623);
nor U19470 (N_19470,N_18903,N_18833);
nand U19471 (N_19471,N_18826,N_19067);
xor U19472 (N_19472,N_19114,N_18755);
or U19473 (N_19473,N_18707,N_18935);
and U19474 (N_19474,N_19018,N_18611);
nand U19475 (N_19475,N_18610,N_18739);
nor U19476 (N_19476,N_18902,N_18671);
nor U19477 (N_19477,N_19171,N_19128);
and U19478 (N_19478,N_18937,N_19071);
or U19479 (N_19479,N_18772,N_18783);
nor U19480 (N_19480,N_18919,N_19049);
nor U19481 (N_19481,N_19031,N_18960);
or U19482 (N_19482,N_18720,N_19196);
nor U19483 (N_19483,N_18744,N_18864);
or U19484 (N_19484,N_18641,N_18662);
and U19485 (N_19485,N_18891,N_18678);
xnor U19486 (N_19486,N_18912,N_19008);
or U19487 (N_19487,N_18725,N_18763);
or U19488 (N_19488,N_18692,N_18688);
nand U19489 (N_19489,N_18918,N_18740);
or U19490 (N_19490,N_19119,N_19112);
nor U19491 (N_19491,N_18659,N_18825);
and U19492 (N_19492,N_18612,N_18687);
xor U19493 (N_19493,N_18860,N_18823);
or U19494 (N_19494,N_18673,N_19099);
nand U19495 (N_19495,N_18979,N_18647);
nor U19496 (N_19496,N_18676,N_18619);
nor U19497 (N_19497,N_18993,N_18751);
and U19498 (N_19498,N_18665,N_18795);
nor U19499 (N_19499,N_18760,N_18729);
nor U19500 (N_19500,N_19025,N_18837);
nand U19501 (N_19501,N_18833,N_18978);
and U19502 (N_19502,N_19078,N_18777);
or U19503 (N_19503,N_18785,N_19170);
and U19504 (N_19504,N_19056,N_18905);
and U19505 (N_19505,N_18890,N_18823);
or U19506 (N_19506,N_19096,N_19138);
nor U19507 (N_19507,N_18859,N_19156);
and U19508 (N_19508,N_19042,N_19046);
or U19509 (N_19509,N_19076,N_19011);
nand U19510 (N_19510,N_18811,N_18869);
or U19511 (N_19511,N_18824,N_19080);
or U19512 (N_19512,N_18982,N_18723);
and U19513 (N_19513,N_18611,N_19041);
xnor U19514 (N_19514,N_18822,N_19120);
nand U19515 (N_19515,N_18836,N_18799);
and U19516 (N_19516,N_18649,N_19096);
nor U19517 (N_19517,N_18867,N_18942);
and U19518 (N_19518,N_19049,N_18733);
nand U19519 (N_19519,N_18834,N_18710);
or U19520 (N_19520,N_18789,N_19173);
nand U19521 (N_19521,N_18620,N_18977);
or U19522 (N_19522,N_19177,N_18744);
nand U19523 (N_19523,N_18875,N_18986);
nand U19524 (N_19524,N_18953,N_18789);
xor U19525 (N_19525,N_18962,N_19000);
nor U19526 (N_19526,N_19064,N_18792);
and U19527 (N_19527,N_19048,N_19033);
xnor U19528 (N_19528,N_18747,N_18769);
nand U19529 (N_19529,N_18949,N_18887);
xnor U19530 (N_19530,N_18700,N_18969);
or U19531 (N_19531,N_18600,N_19027);
nand U19532 (N_19532,N_19005,N_19138);
nor U19533 (N_19533,N_18904,N_18783);
xnor U19534 (N_19534,N_18699,N_18790);
nor U19535 (N_19535,N_18674,N_19094);
and U19536 (N_19536,N_19196,N_19192);
or U19537 (N_19537,N_18966,N_18636);
nand U19538 (N_19538,N_19164,N_19020);
xnor U19539 (N_19539,N_19123,N_18838);
nor U19540 (N_19540,N_18782,N_18797);
nand U19541 (N_19541,N_18707,N_19198);
or U19542 (N_19542,N_19032,N_18613);
or U19543 (N_19543,N_18775,N_18778);
or U19544 (N_19544,N_18985,N_18921);
xnor U19545 (N_19545,N_18920,N_18771);
or U19546 (N_19546,N_19182,N_18812);
xnor U19547 (N_19547,N_19132,N_18612);
or U19548 (N_19548,N_19119,N_18715);
or U19549 (N_19549,N_18715,N_18686);
xnor U19550 (N_19550,N_18722,N_19178);
nand U19551 (N_19551,N_18801,N_18973);
nor U19552 (N_19552,N_18960,N_18606);
nor U19553 (N_19553,N_18914,N_18705);
and U19554 (N_19554,N_18822,N_18948);
or U19555 (N_19555,N_19089,N_18629);
nor U19556 (N_19556,N_19189,N_19166);
nor U19557 (N_19557,N_19194,N_18797);
nor U19558 (N_19558,N_18973,N_18785);
nand U19559 (N_19559,N_18661,N_18634);
nor U19560 (N_19560,N_18923,N_18977);
or U19561 (N_19561,N_18863,N_18748);
or U19562 (N_19562,N_18722,N_18789);
nand U19563 (N_19563,N_19173,N_18882);
and U19564 (N_19564,N_18910,N_18957);
or U19565 (N_19565,N_19037,N_19075);
nor U19566 (N_19566,N_18945,N_19198);
xor U19567 (N_19567,N_19077,N_18729);
and U19568 (N_19568,N_18734,N_19029);
and U19569 (N_19569,N_18999,N_18809);
nand U19570 (N_19570,N_18641,N_18763);
and U19571 (N_19571,N_18687,N_18946);
xor U19572 (N_19572,N_18955,N_18775);
nor U19573 (N_19573,N_18766,N_18800);
nand U19574 (N_19574,N_18671,N_18964);
or U19575 (N_19575,N_18959,N_19052);
nand U19576 (N_19576,N_19144,N_18994);
or U19577 (N_19577,N_18833,N_18794);
or U19578 (N_19578,N_19162,N_19144);
xor U19579 (N_19579,N_18903,N_19198);
nor U19580 (N_19580,N_19022,N_19072);
or U19581 (N_19581,N_18775,N_18658);
nor U19582 (N_19582,N_18949,N_18993);
nand U19583 (N_19583,N_18773,N_18998);
nor U19584 (N_19584,N_18703,N_19062);
nor U19585 (N_19585,N_18691,N_19167);
nand U19586 (N_19586,N_19133,N_18683);
or U19587 (N_19587,N_18833,N_18829);
nor U19588 (N_19588,N_19088,N_18763);
or U19589 (N_19589,N_18694,N_18755);
nand U19590 (N_19590,N_19199,N_19126);
and U19591 (N_19591,N_18709,N_18763);
nand U19592 (N_19592,N_18720,N_18852);
nand U19593 (N_19593,N_18918,N_18863);
and U19594 (N_19594,N_19184,N_18772);
or U19595 (N_19595,N_18727,N_18789);
and U19596 (N_19596,N_18676,N_18976);
or U19597 (N_19597,N_18990,N_18603);
or U19598 (N_19598,N_18699,N_19022);
xnor U19599 (N_19599,N_18782,N_19044);
or U19600 (N_19600,N_18797,N_18980);
or U19601 (N_19601,N_19101,N_19056);
xor U19602 (N_19602,N_19163,N_18715);
xor U19603 (N_19603,N_18852,N_18889);
nor U19604 (N_19604,N_18717,N_18797);
nor U19605 (N_19605,N_19127,N_18929);
or U19606 (N_19606,N_18698,N_18752);
and U19607 (N_19607,N_18984,N_19086);
or U19608 (N_19608,N_19122,N_18642);
or U19609 (N_19609,N_19180,N_18900);
xor U19610 (N_19610,N_18620,N_18618);
or U19611 (N_19611,N_19069,N_18750);
or U19612 (N_19612,N_19124,N_18754);
nor U19613 (N_19613,N_18806,N_18837);
and U19614 (N_19614,N_18808,N_18866);
or U19615 (N_19615,N_19077,N_19025);
or U19616 (N_19616,N_19032,N_19021);
or U19617 (N_19617,N_18837,N_18697);
and U19618 (N_19618,N_18972,N_18915);
or U19619 (N_19619,N_19084,N_19199);
or U19620 (N_19620,N_18643,N_19076);
and U19621 (N_19621,N_19050,N_19129);
nand U19622 (N_19622,N_19030,N_19022);
and U19623 (N_19623,N_18839,N_18812);
nand U19624 (N_19624,N_18760,N_18877);
and U19625 (N_19625,N_18635,N_19133);
and U19626 (N_19626,N_18836,N_19182);
and U19627 (N_19627,N_18998,N_19007);
nand U19628 (N_19628,N_18606,N_18866);
or U19629 (N_19629,N_18879,N_19157);
and U19630 (N_19630,N_18619,N_18646);
and U19631 (N_19631,N_19149,N_18808);
or U19632 (N_19632,N_18820,N_18739);
nor U19633 (N_19633,N_19016,N_18646);
and U19634 (N_19634,N_19026,N_18669);
or U19635 (N_19635,N_18993,N_19151);
or U19636 (N_19636,N_19140,N_18830);
nor U19637 (N_19637,N_19044,N_18668);
xnor U19638 (N_19638,N_19188,N_18743);
xnor U19639 (N_19639,N_18847,N_19135);
xor U19640 (N_19640,N_18647,N_19103);
nor U19641 (N_19641,N_19063,N_18802);
or U19642 (N_19642,N_18674,N_18717);
xor U19643 (N_19643,N_18670,N_18942);
or U19644 (N_19644,N_18869,N_18933);
nor U19645 (N_19645,N_18831,N_19146);
and U19646 (N_19646,N_18961,N_18932);
or U19647 (N_19647,N_18600,N_18932);
nor U19648 (N_19648,N_18879,N_18719);
or U19649 (N_19649,N_19150,N_18704);
or U19650 (N_19650,N_18800,N_18618);
nor U19651 (N_19651,N_18612,N_18767);
nand U19652 (N_19652,N_19177,N_19155);
xor U19653 (N_19653,N_19010,N_18807);
xnor U19654 (N_19654,N_18755,N_18887);
nor U19655 (N_19655,N_19134,N_18866);
or U19656 (N_19656,N_18688,N_19111);
and U19657 (N_19657,N_18901,N_18721);
or U19658 (N_19658,N_18627,N_19044);
or U19659 (N_19659,N_19039,N_18699);
and U19660 (N_19660,N_19088,N_18854);
or U19661 (N_19661,N_19013,N_19123);
nor U19662 (N_19662,N_18863,N_18917);
xnor U19663 (N_19663,N_19173,N_19056);
and U19664 (N_19664,N_18673,N_18828);
nand U19665 (N_19665,N_18856,N_18695);
nor U19666 (N_19666,N_18608,N_18981);
and U19667 (N_19667,N_18872,N_18646);
nor U19668 (N_19668,N_18720,N_18981);
or U19669 (N_19669,N_19115,N_18624);
nand U19670 (N_19670,N_18812,N_18829);
and U19671 (N_19671,N_18865,N_18728);
nand U19672 (N_19672,N_18622,N_18600);
xor U19673 (N_19673,N_19129,N_18913);
and U19674 (N_19674,N_18988,N_19036);
nand U19675 (N_19675,N_18637,N_18825);
and U19676 (N_19676,N_18796,N_18810);
nor U19677 (N_19677,N_18659,N_19031);
and U19678 (N_19678,N_18703,N_18748);
xor U19679 (N_19679,N_18721,N_19009);
nor U19680 (N_19680,N_18633,N_19001);
or U19681 (N_19681,N_19104,N_18820);
nand U19682 (N_19682,N_18995,N_18758);
or U19683 (N_19683,N_18846,N_19019);
nor U19684 (N_19684,N_18850,N_18994);
and U19685 (N_19685,N_18690,N_18787);
or U19686 (N_19686,N_18747,N_18623);
nor U19687 (N_19687,N_18800,N_19164);
nand U19688 (N_19688,N_18726,N_19084);
nand U19689 (N_19689,N_18892,N_18897);
or U19690 (N_19690,N_18836,N_18893);
nand U19691 (N_19691,N_19130,N_18684);
nand U19692 (N_19692,N_19032,N_19115);
nand U19693 (N_19693,N_18786,N_19173);
nand U19694 (N_19694,N_18629,N_18691);
nor U19695 (N_19695,N_19117,N_18979);
nand U19696 (N_19696,N_18920,N_18876);
nor U19697 (N_19697,N_18988,N_18924);
or U19698 (N_19698,N_19029,N_19178);
and U19699 (N_19699,N_18600,N_18822);
or U19700 (N_19700,N_19008,N_19109);
nand U19701 (N_19701,N_19054,N_18800);
and U19702 (N_19702,N_18714,N_18967);
nand U19703 (N_19703,N_19084,N_18673);
or U19704 (N_19704,N_18912,N_18927);
and U19705 (N_19705,N_19067,N_18766);
nand U19706 (N_19706,N_19076,N_19036);
nand U19707 (N_19707,N_18743,N_19090);
or U19708 (N_19708,N_18710,N_19135);
and U19709 (N_19709,N_19070,N_18763);
nor U19710 (N_19710,N_18883,N_18696);
and U19711 (N_19711,N_18979,N_19165);
or U19712 (N_19712,N_18799,N_19084);
and U19713 (N_19713,N_18924,N_19061);
or U19714 (N_19714,N_19126,N_19189);
xnor U19715 (N_19715,N_18654,N_19148);
or U19716 (N_19716,N_19033,N_19172);
and U19717 (N_19717,N_18804,N_18926);
nor U19718 (N_19718,N_18681,N_18793);
nand U19719 (N_19719,N_18656,N_19191);
nor U19720 (N_19720,N_19169,N_18633);
nand U19721 (N_19721,N_18950,N_18962);
nand U19722 (N_19722,N_18633,N_18970);
xnor U19723 (N_19723,N_18712,N_18770);
and U19724 (N_19724,N_18804,N_18748);
or U19725 (N_19725,N_18602,N_18702);
nor U19726 (N_19726,N_18605,N_19033);
and U19727 (N_19727,N_18613,N_19182);
or U19728 (N_19728,N_18737,N_18907);
nor U19729 (N_19729,N_18709,N_18987);
or U19730 (N_19730,N_18602,N_18644);
or U19731 (N_19731,N_18749,N_18732);
and U19732 (N_19732,N_18831,N_18793);
nand U19733 (N_19733,N_18765,N_18976);
nor U19734 (N_19734,N_18645,N_19190);
nor U19735 (N_19735,N_18690,N_18616);
and U19736 (N_19736,N_18805,N_19150);
xor U19737 (N_19737,N_18779,N_18858);
and U19738 (N_19738,N_19114,N_18878);
and U19739 (N_19739,N_18800,N_19180);
and U19740 (N_19740,N_19178,N_19136);
or U19741 (N_19741,N_19134,N_19078);
nand U19742 (N_19742,N_19164,N_19148);
and U19743 (N_19743,N_18909,N_18930);
nand U19744 (N_19744,N_19185,N_19113);
or U19745 (N_19745,N_18857,N_19034);
and U19746 (N_19746,N_18813,N_19160);
or U19747 (N_19747,N_18670,N_18987);
nand U19748 (N_19748,N_18625,N_18692);
nor U19749 (N_19749,N_18621,N_19066);
nand U19750 (N_19750,N_19097,N_18816);
and U19751 (N_19751,N_18832,N_18785);
nor U19752 (N_19752,N_18806,N_18989);
xnor U19753 (N_19753,N_18849,N_19045);
nor U19754 (N_19754,N_19117,N_19035);
and U19755 (N_19755,N_18747,N_18672);
and U19756 (N_19756,N_18745,N_18694);
or U19757 (N_19757,N_18777,N_19132);
or U19758 (N_19758,N_19139,N_18763);
xor U19759 (N_19759,N_18835,N_19024);
and U19760 (N_19760,N_19174,N_19014);
nor U19761 (N_19761,N_18945,N_19089);
or U19762 (N_19762,N_19165,N_19158);
or U19763 (N_19763,N_18728,N_18850);
xnor U19764 (N_19764,N_18844,N_18883);
or U19765 (N_19765,N_18929,N_19092);
nand U19766 (N_19766,N_18610,N_18974);
or U19767 (N_19767,N_18973,N_19071);
and U19768 (N_19768,N_19119,N_19052);
and U19769 (N_19769,N_18632,N_18600);
nor U19770 (N_19770,N_18629,N_18689);
nand U19771 (N_19771,N_18984,N_18996);
nor U19772 (N_19772,N_18698,N_18706);
nand U19773 (N_19773,N_18885,N_19024);
or U19774 (N_19774,N_18744,N_18972);
nor U19775 (N_19775,N_18652,N_18719);
and U19776 (N_19776,N_19076,N_19177);
and U19777 (N_19777,N_18642,N_19143);
xor U19778 (N_19778,N_18837,N_18675);
nor U19779 (N_19779,N_18675,N_19171);
and U19780 (N_19780,N_18695,N_18893);
xor U19781 (N_19781,N_19045,N_19005);
xnor U19782 (N_19782,N_18831,N_19082);
nand U19783 (N_19783,N_19104,N_18900);
or U19784 (N_19784,N_18972,N_18936);
nor U19785 (N_19785,N_19118,N_18976);
xnor U19786 (N_19786,N_19137,N_18995);
nand U19787 (N_19787,N_18985,N_18734);
nor U19788 (N_19788,N_19034,N_18629);
or U19789 (N_19789,N_19045,N_18657);
nor U19790 (N_19790,N_18778,N_18873);
or U19791 (N_19791,N_18988,N_18952);
nor U19792 (N_19792,N_18697,N_18964);
and U19793 (N_19793,N_19166,N_19047);
xnor U19794 (N_19794,N_19130,N_18938);
and U19795 (N_19795,N_18959,N_18649);
and U19796 (N_19796,N_19005,N_19168);
or U19797 (N_19797,N_18853,N_18957);
xnor U19798 (N_19798,N_18997,N_19043);
nand U19799 (N_19799,N_18875,N_18612);
nor U19800 (N_19800,N_19766,N_19420);
and U19801 (N_19801,N_19749,N_19301);
nor U19802 (N_19802,N_19785,N_19285);
nor U19803 (N_19803,N_19362,N_19610);
nor U19804 (N_19804,N_19747,N_19311);
nand U19805 (N_19805,N_19230,N_19632);
nor U19806 (N_19806,N_19452,N_19375);
nand U19807 (N_19807,N_19517,N_19326);
and U19808 (N_19808,N_19595,N_19503);
xor U19809 (N_19809,N_19553,N_19599);
or U19810 (N_19810,N_19560,N_19337);
or U19811 (N_19811,N_19284,N_19729);
nand U19812 (N_19812,N_19657,N_19573);
nand U19813 (N_19813,N_19367,N_19349);
or U19814 (N_19814,N_19440,N_19688);
nor U19815 (N_19815,N_19226,N_19535);
nor U19816 (N_19816,N_19544,N_19561);
and U19817 (N_19817,N_19667,N_19200);
xnor U19818 (N_19818,N_19246,N_19725);
nor U19819 (N_19819,N_19626,N_19460);
and U19820 (N_19820,N_19295,N_19518);
and U19821 (N_19821,N_19355,N_19788);
nand U19822 (N_19822,N_19777,N_19609);
nand U19823 (N_19823,N_19720,N_19548);
or U19824 (N_19824,N_19536,N_19792);
nand U19825 (N_19825,N_19649,N_19247);
nand U19826 (N_19826,N_19443,N_19273);
xor U19827 (N_19827,N_19652,N_19514);
nor U19828 (N_19828,N_19594,N_19695);
or U19829 (N_19829,N_19335,N_19556);
nor U19830 (N_19830,N_19702,N_19395);
nor U19831 (N_19831,N_19575,N_19414);
or U19832 (N_19832,N_19733,N_19308);
nand U19833 (N_19833,N_19306,N_19451);
nand U19834 (N_19834,N_19428,N_19380);
and U19835 (N_19835,N_19486,N_19494);
nand U19836 (N_19836,N_19669,N_19277);
and U19837 (N_19837,N_19520,N_19681);
nand U19838 (N_19838,N_19557,N_19552);
or U19839 (N_19839,N_19319,N_19341);
and U19840 (N_19840,N_19692,N_19764);
or U19841 (N_19841,N_19411,N_19572);
nand U19842 (N_19842,N_19316,N_19331);
and U19843 (N_19843,N_19423,N_19715);
nor U19844 (N_19844,N_19678,N_19434);
nand U19845 (N_19845,N_19369,N_19631);
nand U19846 (N_19846,N_19404,N_19671);
nor U19847 (N_19847,N_19645,N_19579);
and U19848 (N_19848,N_19526,N_19630);
xnor U19849 (N_19849,N_19728,N_19623);
xnor U19850 (N_19850,N_19505,N_19488);
nor U19851 (N_19851,N_19492,N_19710);
nor U19852 (N_19852,N_19429,N_19482);
nor U19853 (N_19853,N_19281,N_19576);
nor U19854 (N_19854,N_19727,N_19405);
xor U19855 (N_19855,N_19241,N_19356);
nor U19856 (N_19856,N_19577,N_19374);
or U19857 (N_19857,N_19453,N_19547);
or U19858 (N_19858,N_19291,N_19770);
nand U19859 (N_19859,N_19605,N_19613);
and U19860 (N_19860,N_19515,N_19581);
nor U19861 (N_19861,N_19406,N_19251);
and U19862 (N_19862,N_19707,N_19475);
and U19863 (N_19863,N_19229,N_19738);
or U19864 (N_19864,N_19397,N_19446);
nand U19865 (N_19865,N_19361,N_19712);
nor U19866 (N_19866,N_19313,N_19264);
or U19867 (N_19867,N_19736,N_19732);
and U19868 (N_19868,N_19675,N_19336);
and U19869 (N_19869,N_19621,N_19762);
or U19870 (N_19870,N_19789,N_19696);
nand U19871 (N_19871,N_19597,N_19783);
xnor U19872 (N_19872,N_19372,N_19786);
nor U19873 (N_19873,N_19297,N_19215);
xnor U19874 (N_19874,N_19292,N_19296);
nand U19875 (N_19875,N_19484,N_19352);
and U19876 (N_19876,N_19245,N_19776);
xor U19877 (N_19877,N_19370,N_19759);
nand U19878 (N_19878,N_19504,N_19703);
nor U19879 (N_19879,N_19701,N_19426);
nand U19880 (N_19880,N_19268,N_19564);
nand U19881 (N_19881,N_19741,N_19340);
xor U19882 (N_19882,N_19353,N_19691);
and U19883 (N_19883,N_19534,N_19430);
and U19884 (N_19884,N_19622,N_19679);
and U19885 (N_19885,N_19646,N_19210);
nand U19886 (N_19886,N_19207,N_19690);
xnor U19887 (N_19887,N_19476,N_19346);
nand U19888 (N_19888,N_19376,N_19262);
nor U19889 (N_19889,N_19590,N_19493);
nor U19890 (N_19890,N_19233,N_19265);
or U19891 (N_19891,N_19619,N_19473);
nand U19892 (N_19892,N_19470,N_19275);
or U19893 (N_19893,N_19522,N_19267);
and U19894 (N_19894,N_19381,N_19742);
nor U19895 (N_19895,N_19775,N_19465);
and U19896 (N_19896,N_19477,N_19379);
and U19897 (N_19897,N_19419,N_19592);
and U19898 (N_19898,N_19364,N_19709);
and U19899 (N_19899,N_19431,N_19586);
and U19900 (N_19900,N_19474,N_19773);
and U19901 (N_19901,N_19538,N_19793);
and U19902 (N_19902,N_19432,N_19211);
or U19903 (N_19903,N_19511,N_19332);
nand U19904 (N_19904,N_19441,N_19236);
and U19905 (N_19905,N_19680,N_19795);
nand U19906 (N_19906,N_19371,N_19617);
xor U19907 (N_19907,N_19532,N_19794);
and U19908 (N_19908,N_19697,N_19303);
nand U19909 (N_19909,N_19598,N_19574);
nand U19910 (N_19910,N_19607,N_19318);
nor U19911 (N_19911,N_19386,N_19366);
nor U19912 (N_19912,N_19549,N_19286);
and U19913 (N_19913,N_19490,N_19463);
nand U19914 (N_19914,N_19221,N_19323);
or U19915 (N_19915,N_19704,N_19730);
or U19916 (N_19916,N_19449,N_19798);
xor U19917 (N_19917,N_19653,N_19604);
and U19918 (N_19918,N_19334,N_19300);
nand U19919 (N_19919,N_19464,N_19589);
and U19920 (N_19920,N_19700,N_19350);
or U19921 (N_19921,N_19540,N_19252);
or U19922 (N_19922,N_19787,N_19745);
nor U19923 (N_19923,N_19612,N_19363);
nor U19924 (N_19924,N_19771,N_19239);
nand U19925 (N_19925,N_19317,N_19674);
and U19926 (N_19926,N_19243,N_19743);
and U19927 (N_19927,N_19461,N_19748);
nor U19928 (N_19928,N_19791,N_19280);
or U19929 (N_19929,N_19289,N_19706);
nand U19930 (N_19930,N_19708,N_19663);
xnor U19931 (N_19931,N_19261,N_19278);
nor U19932 (N_19932,N_19591,N_19302);
xnor U19933 (N_19933,N_19714,N_19322);
and U19934 (N_19934,N_19389,N_19304);
xnor U19935 (N_19935,N_19769,N_19781);
or U19936 (N_19936,N_19587,N_19378);
and U19937 (N_19937,N_19754,N_19424);
nand U19938 (N_19938,N_19283,N_19227);
and U19939 (N_19939,N_19348,N_19611);
nor U19940 (N_19940,N_19772,N_19676);
nor U19941 (N_19941,N_19501,N_19539);
xnor U19942 (N_19942,N_19249,N_19498);
nand U19943 (N_19943,N_19293,N_19479);
or U19944 (N_19944,N_19385,N_19750);
nand U19945 (N_19945,N_19299,N_19687);
nor U19946 (N_19946,N_19530,N_19433);
or U19947 (N_19947,N_19782,N_19760);
and U19948 (N_19948,N_19571,N_19529);
nand U19949 (N_19949,N_19224,N_19545);
nor U19950 (N_19950,N_19507,N_19537);
nand U19951 (N_19951,N_19602,N_19359);
nand U19952 (N_19952,N_19244,N_19784);
nor U19953 (N_19953,N_19722,N_19478);
or U19954 (N_19954,N_19480,N_19753);
and U19955 (N_19955,N_19796,N_19664);
nor U19956 (N_19956,N_19481,N_19358);
or U19957 (N_19957,N_19439,N_19287);
xnor U19958 (N_19958,N_19391,N_19237);
or U19959 (N_19959,N_19662,N_19528);
and U19960 (N_19960,N_19469,N_19636);
or U19961 (N_19961,N_19368,N_19487);
and U19962 (N_19962,N_19416,N_19606);
or U19963 (N_19963,N_19684,N_19578);
nor U19964 (N_19964,N_19437,N_19740);
nand U19965 (N_19965,N_19248,N_19569);
nor U19966 (N_19966,N_19394,N_19288);
and U19967 (N_19967,N_19214,N_19307);
and U19968 (N_19968,N_19580,N_19731);
or U19969 (N_19969,N_19543,N_19585);
nor U19970 (N_19970,N_19677,N_19392);
and U19971 (N_19971,N_19400,N_19256);
or U19972 (N_19972,N_19527,N_19413);
and U19973 (N_19973,N_19351,N_19459);
xnor U19974 (N_19974,N_19542,N_19330);
nand U19975 (N_19975,N_19567,N_19625);
or U19976 (N_19976,N_19550,N_19628);
nand U19977 (N_19977,N_19765,N_19314);
nor U19978 (N_19978,N_19398,N_19685);
or U19979 (N_19979,N_19618,N_19635);
nor U19980 (N_19980,N_19755,N_19325);
nand U19981 (N_19981,N_19506,N_19235);
or U19982 (N_19982,N_19694,N_19497);
or U19983 (N_19983,N_19240,N_19570);
and U19984 (N_19984,N_19758,N_19468);
and U19985 (N_19985,N_19454,N_19219);
nor U19986 (N_19986,N_19255,N_19661);
nor U19987 (N_19987,N_19670,N_19533);
and U19988 (N_19988,N_19436,N_19205);
nor U19989 (N_19989,N_19382,N_19624);
nor U19990 (N_19990,N_19383,N_19711);
nor U19991 (N_19991,N_19225,N_19583);
and U19992 (N_19992,N_19417,N_19799);
nor U19993 (N_19993,N_19489,N_19726);
nor U19994 (N_19994,N_19387,N_19377);
or U19995 (N_19995,N_19408,N_19551);
or U19996 (N_19996,N_19555,N_19458);
or U19997 (N_19997,N_19354,N_19797);
xor U19998 (N_19998,N_19365,N_19495);
or U19999 (N_19999,N_19310,N_19234);
and U20000 (N_20000,N_19329,N_19541);
nand U20001 (N_20001,N_19209,N_19500);
nor U20002 (N_20002,N_19201,N_19388);
and U20003 (N_20003,N_19683,N_19524);
nand U20004 (N_20004,N_19312,N_19309);
and U20005 (N_20005,N_19202,N_19217);
or U20006 (N_20006,N_19584,N_19735);
nor U20007 (N_20007,N_19223,N_19333);
nand U20008 (N_20008,N_19212,N_19682);
nor U20009 (N_20009,N_19659,N_19568);
nor U20010 (N_20010,N_19620,N_19409);
xor U20011 (N_20011,N_19637,N_19713);
xor U20012 (N_20012,N_19693,N_19525);
nor U20013 (N_20013,N_19327,N_19258);
and U20014 (N_20014,N_19744,N_19401);
nor U20015 (N_20015,N_19641,N_19238);
nand U20016 (N_20016,N_19338,N_19774);
nor U20017 (N_20017,N_19634,N_19588);
nand U20018 (N_20018,N_19644,N_19467);
nand U20019 (N_20019,N_19344,N_19719);
nand U20020 (N_20020,N_19655,N_19686);
or U20021 (N_20021,N_19457,N_19546);
and U20022 (N_20022,N_19448,N_19734);
or U20023 (N_20023,N_19294,N_19425);
nor U20024 (N_20024,N_19629,N_19393);
nand U20025 (N_20025,N_19204,N_19259);
nor U20026 (N_20026,N_19444,N_19271);
and U20027 (N_20027,N_19421,N_19206);
and U20028 (N_20028,N_19757,N_19402);
nand U20029 (N_20029,N_19274,N_19208);
nand U20030 (N_20030,N_19563,N_19603);
and U20031 (N_20031,N_19455,N_19407);
xnor U20032 (N_20032,N_19582,N_19639);
or U20033 (N_20033,N_19608,N_19510);
or U20034 (N_20034,N_19672,N_19345);
nand U20035 (N_20035,N_19650,N_19660);
nor U20036 (N_20036,N_19499,N_19739);
nand U20037 (N_20037,N_19435,N_19324);
nand U20038 (N_20038,N_19254,N_19565);
nor U20039 (N_20039,N_19519,N_19705);
or U20040 (N_20040,N_19559,N_19640);
and U20041 (N_20041,N_19410,N_19509);
or U20042 (N_20042,N_19315,N_19399);
and U20043 (N_20043,N_19718,N_19232);
and U20044 (N_20044,N_19415,N_19462);
nor U20045 (N_20045,N_19778,N_19203);
and U20046 (N_20046,N_19531,N_19767);
nand U20047 (N_20047,N_19768,N_19242);
nor U20048 (N_20048,N_19456,N_19665);
nor U20049 (N_20049,N_19260,N_19347);
and U20050 (N_20050,N_19373,N_19321);
or U20051 (N_20051,N_19566,N_19222);
or U20052 (N_20052,N_19633,N_19647);
nand U20053 (N_20053,N_19554,N_19780);
nor U20054 (N_20054,N_19231,N_19513);
nor U20055 (N_20055,N_19651,N_19716);
nand U20056 (N_20056,N_19658,N_19752);
nand U20057 (N_20057,N_19562,N_19627);
and U20058 (N_20058,N_19218,N_19496);
nand U20059 (N_20059,N_19508,N_19601);
nand U20060 (N_20060,N_19216,N_19220);
nor U20061 (N_20061,N_19269,N_19756);
or U20062 (N_20062,N_19339,N_19523);
nor U20063 (N_20063,N_19442,N_19790);
nand U20064 (N_20064,N_19761,N_19412);
nand U20065 (N_20065,N_19616,N_19521);
or U20066 (N_20066,N_19516,N_19596);
and U20067 (N_20067,N_19512,N_19485);
nor U20068 (N_20068,N_19638,N_19253);
or U20069 (N_20069,N_19422,N_19558);
and U20070 (N_20070,N_19746,N_19384);
nand U20071 (N_20071,N_19698,N_19257);
and U20072 (N_20072,N_19357,N_19290);
xor U20073 (N_20073,N_19491,N_19343);
nor U20074 (N_20074,N_19279,N_19614);
nand U20075 (N_20075,N_19445,N_19418);
nor U20076 (N_20076,N_19250,N_19751);
nand U20077 (N_20077,N_19648,N_19656);
nand U20078 (N_20078,N_19593,N_19483);
nand U20079 (N_20079,N_19471,N_19390);
nand U20080 (N_20080,N_19320,N_19450);
nor U20081 (N_20081,N_19228,N_19342);
and U20082 (N_20082,N_19666,N_19763);
or U20083 (N_20083,N_19403,N_19723);
and U20084 (N_20084,N_19266,N_19270);
nor U20085 (N_20085,N_19276,N_19615);
nor U20086 (N_20086,N_19654,N_19673);
nor U20087 (N_20087,N_19779,N_19643);
nand U20088 (N_20088,N_19298,N_19396);
or U20089 (N_20089,N_19272,N_19263);
or U20090 (N_20090,N_19472,N_19213);
nand U20091 (N_20091,N_19360,N_19724);
xnor U20092 (N_20092,N_19689,N_19668);
nand U20093 (N_20093,N_19699,N_19438);
and U20094 (N_20094,N_19466,N_19642);
nand U20095 (N_20095,N_19305,N_19721);
or U20096 (N_20096,N_19328,N_19717);
nor U20097 (N_20097,N_19737,N_19600);
or U20098 (N_20098,N_19427,N_19502);
or U20099 (N_20099,N_19282,N_19447);
nand U20100 (N_20100,N_19393,N_19543);
nand U20101 (N_20101,N_19590,N_19392);
and U20102 (N_20102,N_19389,N_19545);
or U20103 (N_20103,N_19595,N_19387);
nor U20104 (N_20104,N_19228,N_19221);
xor U20105 (N_20105,N_19511,N_19214);
nand U20106 (N_20106,N_19643,N_19210);
nand U20107 (N_20107,N_19416,N_19518);
and U20108 (N_20108,N_19239,N_19405);
or U20109 (N_20109,N_19391,N_19246);
nand U20110 (N_20110,N_19726,N_19647);
or U20111 (N_20111,N_19672,N_19780);
nand U20112 (N_20112,N_19496,N_19662);
nor U20113 (N_20113,N_19696,N_19644);
xor U20114 (N_20114,N_19627,N_19766);
xor U20115 (N_20115,N_19733,N_19413);
nor U20116 (N_20116,N_19368,N_19309);
or U20117 (N_20117,N_19515,N_19486);
nand U20118 (N_20118,N_19483,N_19282);
and U20119 (N_20119,N_19672,N_19475);
nand U20120 (N_20120,N_19440,N_19490);
or U20121 (N_20121,N_19485,N_19617);
nand U20122 (N_20122,N_19384,N_19321);
and U20123 (N_20123,N_19238,N_19588);
or U20124 (N_20124,N_19268,N_19626);
nand U20125 (N_20125,N_19561,N_19530);
nor U20126 (N_20126,N_19570,N_19263);
and U20127 (N_20127,N_19286,N_19439);
or U20128 (N_20128,N_19288,N_19232);
and U20129 (N_20129,N_19213,N_19467);
xor U20130 (N_20130,N_19753,N_19734);
nand U20131 (N_20131,N_19793,N_19726);
and U20132 (N_20132,N_19353,N_19378);
and U20133 (N_20133,N_19614,N_19693);
or U20134 (N_20134,N_19562,N_19757);
nor U20135 (N_20135,N_19260,N_19321);
and U20136 (N_20136,N_19435,N_19205);
nand U20137 (N_20137,N_19308,N_19794);
nor U20138 (N_20138,N_19467,N_19711);
and U20139 (N_20139,N_19304,N_19553);
nand U20140 (N_20140,N_19676,N_19205);
nand U20141 (N_20141,N_19770,N_19491);
or U20142 (N_20142,N_19220,N_19748);
and U20143 (N_20143,N_19555,N_19444);
nor U20144 (N_20144,N_19550,N_19349);
nand U20145 (N_20145,N_19419,N_19577);
nor U20146 (N_20146,N_19713,N_19583);
and U20147 (N_20147,N_19615,N_19692);
and U20148 (N_20148,N_19540,N_19355);
nor U20149 (N_20149,N_19671,N_19678);
xnor U20150 (N_20150,N_19665,N_19707);
or U20151 (N_20151,N_19450,N_19268);
or U20152 (N_20152,N_19386,N_19451);
nand U20153 (N_20153,N_19316,N_19690);
and U20154 (N_20154,N_19632,N_19281);
nor U20155 (N_20155,N_19659,N_19645);
nand U20156 (N_20156,N_19656,N_19409);
or U20157 (N_20157,N_19751,N_19712);
and U20158 (N_20158,N_19570,N_19558);
or U20159 (N_20159,N_19700,N_19571);
nor U20160 (N_20160,N_19477,N_19473);
nor U20161 (N_20161,N_19715,N_19385);
nor U20162 (N_20162,N_19319,N_19567);
and U20163 (N_20163,N_19419,N_19616);
nand U20164 (N_20164,N_19723,N_19249);
or U20165 (N_20165,N_19567,N_19797);
and U20166 (N_20166,N_19271,N_19204);
or U20167 (N_20167,N_19503,N_19233);
and U20168 (N_20168,N_19670,N_19531);
or U20169 (N_20169,N_19420,N_19549);
xor U20170 (N_20170,N_19238,N_19704);
nor U20171 (N_20171,N_19299,N_19612);
or U20172 (N_20172,N_19670,N_19339);
xor U20173 (N_20173,N_19604,N_19799);
nand U20174 (N_20174,N_19280,N_19339);
and U20175 (N_20175,N_19320,N_19687);
or U20176 (N_20176,N_19658,N_19726);
nor U20177 (N_20177,N_19575,N_19554);
xor U20178 (N_20178,N_19626,N_19220);
nor U20179 (N_20179,N_19409,N_19222);
and U20180 (N_20180,N_19750,N_19451);
nor U20181 (N_20181,N_19554,N_19309);
nor U20182 (N_20182,N_19752,N_19400);
and U20183 (N_20183,N_19413,N_19269);
or U20184 (N_20184,N_19308,N_19691);
or U20185 (N_20185,N_19233,N_19674);
or U20186 (N_20186,N_19332,N_19400);
nand U20187 (N_20187,N_19719,N_19511);
nor U20188 (N_20188,N_19504,N_19621);
and U20189 (N_20189,N_19402,N_19433);
and U20190 (N_20190,N_19472,N_19411);
nor U20191 (N_20191,N_19302,N_19430);
and U20192 (N_20192,N_19488,N_19600);
nand U20193 (N_20193,N_19379,N_19463);
xor U20194 (N_20194,N_19566,N_19397);
nor U20195 (N_20195,N_19673,N_19705);
xor U20196 (N_20196,N_19593,N_19516);
nor U20197 (N_20197,N_19258,N_19578);
or U20198 (N_20198,N_19368,N_19461);
and U20199 (N_20199,N_19302,N_19346);
nor U20200 (N_20200,N_19326,N_19658);
nand U20201 (N_20201,N_19544,N_19602);
nand U20202 (N_20202,N_19349,N_19721);
or U20203 (N_20203,N_19457,N_19269);
or U20204 (N_20204,N_19551,N_19488);
or U20205 (N_20205,N_19615,N_19380);
nor U20206 (N_20206,N_19354,N_19773);
nor U20207 (N_20207,N_19524,N_19225);
nand U20208 (N_20208,N_19739,N_19635);
nand U20209 (N_20209,N_19678,N_19422);
nor U20210 (N_20210,N_19726,N_19796);
and U20211 (N_20211,N_19526,N_19678);
or U20212 (N_20212,N_19262,N_19651);
nand U20213 (N_20213,N_19654,N_19265);
and U20214 (N_20214,N_19655,N_19741);
nor U20215 (N_20215,N_19686,N_19660);
nand U20216 (N_20216,N_19225,N_19350);
xnor U20217 (N_20217,N_19296,N_19322);
nand U20218 (N_20218,N_19314,N_19641);
and U20219 (N_20219,N_19642,N_19392);
or U20220 (N_20220,N_19215,N_19298);
and U20221 (N_20221,N_19352,N_19520);
xnor U20222 (N_20222,N_19326,N_19374);
nand U20223 (N_20223,N_19614,N_19645);
nor U20224 (N_20224,N_19721,N_19662);
nor U20225 (N_20225,N_19267,N_19775);
nand U20226 (N_20226,N_19589,N_19765);
or U20227 (N_20227,N_19799,N_19455);
nand U20228 (N_20228,N_19308,N_19321);
and U20229 (N_20229,N_19290,N_19431);
or U20230 (N_20230,N_19422,N_19559);
nand U20231 (N_20231,N_19599,N_19469);
xnor U20232 (N_20232,N_19679,N_19353);
or U20233 (N_20233,N_19478,N_19630);
and U20234 (N_20234,N_19354,N_19788);
nand U20235 (N_20235,N_19261,N_19275);
or U20236 (N_20236,N_19678,N_19493);
and U20237 (N_20237,N_19381,N_19427);
and U20238 (N_20238,N_19758,N_19477);
nand U20239 (N_20239,N_19211,N_19676);
nor U20240 (N_20240,N_19410,N_19587);
and U20241 (N_20241,N_19328,N_19469);
nor U20242 (N_20242,N_19345,N_19389);
and U20243 (N_20243,N_19451,N_19738);
or U20244 (N_20244,N_19404,N_19563);
nand U20245 (N_20245,N_19775,N_19734);
nor U20246 (N_20246,N_19455,N_19386);
nor U20247 (N_20247,N_19484,N_19670);
and U20248 (N_20248,N_19406,N_19761);
xor U20249 (N_20249,N_19312,N_19253);
nor U20250 (N_20250,N_19226,N_19621);
and U20251 (N_20251,N_19766,N_19235);
xor U20252 (N_20252,N_19343,N_19330);
or U20253 (N_20253,N_19435,N_19672);
and U20254 (N_20254,N_19591,N_19441);
and U20255 (N_20255,N_19645,N_19456);
and U20256 (N_20256,N_19762,N_19612);
or U20257 (N_20257,N_19709,N_19314);
nand U20258 (N_20258,N_19783,N_19771);
and U20259 (N_20259,N_19459,N_19737);
or U20260 (N_20260,N_19326,N_19562);
or U20261 (N_20261,N_19302,N_19445);
or U20262 (N_20262,N_19651,N_19453);
nor U20263 (N_20263,N_19305,N_19590);
or U20264 (N_20264,N_19752,N_19720);
or U20265 (N_20265,N_19252,N_19539);
nand U20266 (N_20266,N_19541,N_19446);
nand U20267 (N_20267,N_19277,N_19470);
nor U20268 (N_20268,N_19306,N_19739);
and U20269 (N_20269,N_19392,N_19726);
nor U20270 (N_20270,N_19678,N_19347);
nor U20271 (N_20271,N_19695,N_19576);
and U20272 (N_20272,N_19607,N_19680);
nand U20273 (N_20273,N_19515,N_19407);
nand U20274 (N_20274,N_19696,N_19242);
nand U20275 (N_20275,N_19225,N_19472);
or U20276 (N_20276,N_19353,N_19478);
nor U20277 (N_20277,N_19631,N_19427);
and U20278 (N_20278,N_19636,N_19474);
nor U20279 (N_20279,N_19379,N_19660);
xor U20280 (N_20280,N_19652,N_19269);
nand U20281 (N_20281,N_19430,N_19285);
nor U20282 (N_20282,N_19507,N_19710);
nand U20283 (N_20283,N_19798,N_19641);
and U20284 (N_20284,N_19665,N_19701);
and U20285 (N_20285,N_19574,N_19729);
nor U20286 (N_20286,N_19612,N_19312);
and U20287 (N_20287,N_19207,N_19706);
nor U20288 (N_20288,N_19368,N_19202);
or U20289 (N_20289,N_19348,N_19379);
nand U20290 (N_20290,N_19357,N_19224);
nand U20291 (N_20291,N_19706,N_19470);
and U20292 (N_20292,N_19344,N_19569);
nand U20293 (N_20293,N_19317,N_19230);
or U20294 (N_20294,N_19647,N_19632);
nor U20295 (N_20295,N_19440,N_19375);
nand U20296 (N_20296,N_19777,N_19311);
xor U20297 (N_20297,N_19709,N_19698);
nor U20298 (N_20298,N_19412,N_19642);
nor U20299 (N_20299,N_19714,N_19702);
and U20300 (N_20300,N_19411,N_19770);
and U20301 (N_20301,N_19651,N_19275);
nand U20302 (N_20302,N_19530,N_19352);
xor U20303 (N_20303,N_19371,N_19708);
nor U20304 (N_20304,N_19582,N_19216);
and U20305 (N_20305,N_19763,N_19578);
nor U20306 (N_20306,N_19249,N_19245);
nand U20307 (N_20307,N_19395,N_19570);
nor U20308 (N_20308,N_19300,N_19438);
nand U20309 (N_20309,N_19728,N_19304);
and U20310 (N_20310,N_19245,N_19561);
xnor U20311 (N_20311,N_19340,N_19682);
or U20312 (N_20312,N_19725,N_19215);
nand U20313 (N_20313,N_19218,N_19604);
and U20314 (N_20314,N_19626,N_19261);
nor U20315 (N_20315,N_19503,N_19576);
nor U20316 (N_20316,N_19494,N_19639);
nand U20317 (N_20317,N_19254,N_19429);
nand U20318 (N_20318,N_19513,N_19219);
nor U20319 (N_20319,N_19643,N_19740);
and U20320 (N_20320,N_19550,N_19257);
or U20321 (N_20321,N_19423,N_19556);
nand U20322 (N_20322,N_19457,N_19498);
nand U20323 (N_20323,N_19410,N_19372);
nand U20324 (N_20324,N_19431,N_19227);
or U20325 (N_20325,N_19329,N_19343);
and U20326 (N_20326,N_19775,N_19288);
or U20327 (N_20327,N_19251,N_19677);
and U20328 (N_20328,N_19259,N_19584);
nand U20329 (N_20329,N_19676,N_19572);
or U20330 (N_20330,N_19571,N_19696);
or U20331 (N_20331,N_19695,N_19593);
xor U20332 (N_20332,N_19446,N_19721);
xor U20333 (N_20333,N_19639,N_19728);
nand U20334 (N_20334,N_19660,N_19585);
and U20335 (N_20335,N_19674,N_19537);
or U20336 (N_20336,N_19759,N_19702);
or U20337 (N_20337,N_19623,N_19532);
and U20338 (N_20338,N_19783,N_19488);
nor U20339 (N_20339,N_19395,N_19541);
nor U20340 (N_20340,N_19588,N_19234);
and U20341 (N_20341,N_19214,N_19200);
and U20342 (N_20342,N_19694,N_19634);
or U20343 (N_20343,N_19229,N_19288);
and U20344 (N_20344,N_19375,N_19675);
and U20345 (N_20345,N_19365,N_19545);
or U20346 (N_20346,N_19303,N_19377);
or U20347 (N_20347,N_19700,N_19570);
nor U20348 (N_20348,N_19403,N_19676);
or U20349 (N_20349,N_19426,N_19497);
xnor U20350 (N_20350,N_19765,N_19459);
nand U20351 (N_20351,N_19482,N_19215);
and U20352 (N_20352,N_19667,N_19528);
nand U20353 (N_20353,N_19236,N_19707);
nand U20354 (N_20354,N_19486,N_19655);
or U20355 (N_20355,N_19743,N_19797);
nor U20356 (N_20356,N_19498,N_19646);
nand U20357 (N_20357,N_19759,N_19780);
and U20358 (N_20358,N_19345,N_19218);
nor U20359 (N_20359,N_19331,N_19619);
and U20360 (N_20360,N_19708,N_19367);
nand U20361 (N_20361,N_19522,N_19653);
or U20362 (N_20362,N_19366,N_19541);
or U20363 (N_20363,N_19747,N_19236);
nor U20364 (N_20364,N_19222,N_19338);
nand U20365 (N_20365,N_19787,N_19646);
or U20366 (N_20366,N_19265,N_19603);
or U20367 (N_20367,N_19235,N_19341);
nand U20368 (N_20368,N_19494,N_19439);
nand U20369 (N_20369,N_19240,N_19600);
nand U20370 (N_20370,N_19349,N_19725);
nor U20371 (N_20371,N_19371,N_19268);
nand U20372 (N_20372,N_19784,N_19627);
nand U20373 (N_20373,N_19401,N_19233);
nand U20374 (N_20374,N_19343,N_19544);
nand U20375 (N_20375,N_19494,N_19690);
nor U20376 (N_20376,N_19662,N_19285);
or U20377 (N_20377,N_19577,N_19716);
or U20378 (N_20378,N_19418,N_19246);
and U20379 (N_20379,N_19316,N_19768);
and U20380 (N_20380,N_19253,N_19339);
nor U20381 (N_20381,N_19797,N_19687);
or U20382 (N_20382,N_19268,N_19546);
and U20383 (N_20383,N_19791,N_19792);
or U20384 (N_20384,N_19522,N_19464);
nor U20385 (N_20385,N_19676,N_19368);
and U20386 (N_20386,N_19412,N_19680);
and U20387 (N_20387,N_19430,N_19486);
or U20388 (N_20388,N_19281,N_19581);
or U20389 (N_20389,N_19210,N_19593);
or U20390 (N_20390,N_19783,N_19519);
or U20391 (N_20391,N_19266,N_19250);
nand U20392 (N_20392,N_19640,N_19343);
xor U20393 (N_20393,N_19284,N_19762);
and U20394 (N_20394,N_19309,N_19750);
and U20395 (N_20395,N_19529,N_19339);
xor U20396 (N_20396,N_19390,N_19797);
xnor U20397 (N_20397,N_19650,N_19687);
nand U20398 (N_20398,N_19666,N_19363);
or U20399 (N_20399,N_19325,N_19240);
or U20400 (N_20400,N_20197,N_19887);
and U20401 (N_20401,N_19934,N_19865);
xnor U20402 (N_20402,N_20387,N_20179);
and U20403 (N_20403,N_20101,N_19949);
nor U20404 (N_20404,N_20004,N_20284);
nor U20405 (N_20405,N_19946,N_20134);
and U20406 (N_20406,N_20354,N_19855);
xnor U20407 (N_20407,N_20085,N_19896);
xnor U20408 (N_20408,N_20056,N_20224);
nand U20409 (N_20409,N_20283,N_19931);
and U20410 (N_20410,N_20306,N_19952);
nand U20411 (N_20411,N_20291,N_20045);
xor U20412 (N_20412,N_20279,N_20285);
nand U20413 (N_20413,N_20329,N_19820);
nor U20414 (N_20414,N_20181,N_20390);
and U20415 (N_20415,N_20064,N_20212);
and U20416 (N_20416,N_20346,N_20046);
and U20417 (N_20417,N_19812,N_20153);
and U20418 (N_20418,N_20298,N_20376);
or U20419 (N_20419,N_20108,N_20361);
nor U20420 (N_20420,N_20099,N_20371);
nand U20421 (N_20421,N_19907,N_20245);
nand U20422 (N_20422,N_20066,N_19961);
and U20423 (N_20423,N_20198,N_19885);
nand U20424 (N_20424,N_20318,N_19954);
or U20425 (N_20425,N_20143,N_20276);
or U20426 (N_20426,N_19884,N_20208);
or U20427 (N_20427,N_19800,N_19994);
or U20428 (N_20428,N_20128,N_20297);
and U20429 (N_20429,N_20089,N_20104);
and U20430 (N_20430,N_20021,N_19971);
nor U20431 (N_20431,N_20093,N_20012);
nor U20432 (N_20432,N_20055,N_19891);
nor U20433 (N_20433,N_20249,N_20049);
nand U20434 (N_20434,N_20009,N_20278);
or U20435 (N_20435,N_20362,N_19851);
and U20436 (N_20436,N_20023,N_20020);
and U20437 (N_20437,N_19909,N_20203);
or U20438 (N_20438,N_19916,N_20087);
or U20439 (N_20439,N_20303,N_20264);
and U20440 (N_20440,N_20184,N_20137);
nor U20441 (N_20441,N_20215,N_19968);
xor U20442 (N_20442,N_19930,N_19823);
and U20443 (N_20443,N_20373,N_20247);
and U20444 (N_20444,N_20384,N_20206);
and U20445 (N_20445,N_19809,N_19978);
and U20446 (N_20446,N_20383,N_20214);
nand U20447 (N_20447,N_19806,N_20006);
nor U20448 (N_20448,N_20209,N_20251);
and U20449 (N_20449,N_20075,N_20292);
and U20450 (N_20450,N_19827,N_19977);
and U20451 (N_20451,N_20230,N_19955);
and U20452 (N_20452,N_20051,N_20252);
or U20453 (N_20453,N_20146,N_19863);
and U20454 (N_20454,N_20142,N_20183);
nand U20455 (N_20455,N_20368,N_19811);
or U20456 (N_20456,N_20310,N_20242);
xnor U20457 (N_20457,N_20335,N_19849);
or U20458 (N_20458,N_20352,N_20217);
and U20459 (N_20459,N_20305,N_20240);
and U20460 (N_20460,N_20364,N_19973);
and U20461 (N_20461,N_20162,N_20052);
nor U20462 (N_20462,N_20321,N_19964);
or U20463 (N_20463,N_20059,N_19861);
and U20464 (N_20464,N_20271,N_20088);
xnor U20465 (N_20465,N_20355,N_19999);
nor U20466 (N_20466,N_19997,N_20380);
or U20467 (N_20467,N_19804,N_20370);
nand U20468 (N_20468,N_20084,N_19830);
and U20469 (N_20469,N_20317,N_20047);
nand U20470 (N_20470,N_19810,N_19938);
nor U20471 (N_20471,N_20136,N_19932);
and U20472 (N_20472,N_19988,N_20116);
xnor U20473 (N_20473,N_19879,N_19859);
or U20474 (N_20474,N_20316,N_19877);
or U20475 (N_20475,N_20145,N_19819);
and U20476 (N_20476,N_19857,N_20113);
nand U20477 (N_20477,N_20304,N_20274);
and U20478 (N_20478,N_20107,N_19948);
nand U20479 (N_20479,N_19917,N_20094);
nand U20480 (N_20480,N_20092,N_20349);
or U20481 (N_20481,N_20031,N_19981);
nand U20482 (N_20482,N_20180,N_20097);
or U20483 (N_20483,N_20071,N_20398);
nand U20484 (N_20484,N_19963,N_20253);
nor U20485 (N_20485,N_20381,N_19922);
nand U20486 (N_20486,N_20313,N_19956);
nand U20487 (N_20487,N_20225,N_20201);
nand U20488 (N_20488,N_20369,N_20336);
nand U20489 (N_20489,N_20044,N_20377);
nand U20490 (N_20490,N_19870,N_20156);
nor U20491 (N_20491,N_20098,N_20234);
or U20492 (N_20492,N_20299,N_20102);
nand U20493 (N_20493,N_20365,N_20266);
and U20494 (N_20494,N_19921,N_20168);
nor U20495 (N_20495,N_20110,N_20348);
nor U20496 (N_20496,N_20152,N_19803);
or U20497 (N_20497,N_19892,N_20123);
and U20498 (N_20498,N_19894,N_20360);
or U20499 (N_20499,N_20175,N_20246);
or U20500 (N_20500,N_19805,N_19966);
xor U20501 (N_20501,N_19841,N_20219);
nor U20502 (N_20502,N_20058,N_20312);
nor U20503 (N_20503,N_19957,N_19869);
nor U20504 (N_20504,N_20353,N_19993);
nand U20505 (N_20505,N_20151,N_19985);
nor U20506 (N_20506,N_20204,N_19889);
nand U20507 (N_20507,N_20005,N_20135);
nor U20508 (N_20508,N_19846,N_20273);
nor U20509 (N_20509,N_20386,N_20391);
and U20510 (N_20510,N_20029,N_19911);
nand U20511 (N_20511,N_20163,N_20030);
xor U20512 (N_20512,N_20257,N_20345);
nor U20513 (N_20513,N_19888,N_19817);
or U20514 (N_20514,N_20149,N_19845);
and U20515 (N_20515,N_20248,N_20038);
nor U20516 (N_20516,N_20037,N_19920);
nand U20517 (N_20517,N_20119,N_20262);
or U20518 (N_20518,N_20300,N_20309);
and U20519 (N_20519,N_19871,N_20091);
nand U20520 (N_20520,N_20339,N_20036);
or U20521 (N_20521,N_20269,N_19893);
or U20522 (N_20522,N_20019,N_19953);
or U20523 (N_20523,N_19942,N_20025);
and U20524 (N_20524,N_20060,N_20379);
and U20525 (N_20525,N_20182,N_20120);
or U20526 (N_20526,N_19915,N_20256);
and U20527 (N_20527,N_20158,N_19959);
or U20528 (N_20528,N_20086,N_20307);
nor U20529 (N_20529,N_19814,N_19912);
or U20530 (N_20530,N_19828,N_20069);
nor U20531 (N_20531,N_20039,N_20280);
nand U20532 (N_20532,N_19832,N_19943);
nand U20533 (N_20533,N_20199,N_20311);
and U20534 (N_20534,N_20260,N_20125);
nor U20535 (N_20535,N_20105,N_20067);
nand U20536 (N_20536,N_20337,N_20043);
nor U20537 (N_20537,N_20079,N_20357);
or U20538 (N_20538,N_20032,N_20026);
and U20539 (N_20539,N_20147,N_20121);
nor U20540 (N_20540,N_19883,N_20063);
and U20541 (N_20541,N_20027,N_19940);
nand U20542 (N_20542,N_19902,N_19808);
or U20543 (N_20543,N_19886,N_20267);
nor U20544 (N_20544,N_19867,N_19880);
nand U20545 (N_20545,N_20083,N_20341);
and U20546 (N_20546,N_19908,N_19876);
or U20547 (N_20547,N_20195,N_19937);
or U20548 (N_20548,N_20127,N_20315);
or U20549 (N_20549,N_20001,N_20392);
nor U20550 (N_20550,N_20344,N_20161);
and U20551 (N_20551,N_20040,N_20073);
nor U20552 (N_20552,N_20275,N_20374);
and U20553 (N_20553,N_20057,N_20293);
nor U20554 (N_20554,N_20103,N_20393);
and U20555 (N_20555,N_19825,N_19935);
nor U20556 (N_20556,N_20114,N_20078);
and U20557 (N_20557,N_20241,N_20395);
nand U20558 (N_20558,N_19882,N_20216);
and U20559 (N_20559,N_20016,N_19853);
nor U20560 (N_20560,N_20272,N_20132);
nand U20561 (N_20561,N_20333,N_19897);
nand U20562 (N_20562,N_20124,N_19833);
or U20563 (N_20563,N_20160,N_19898);
and U20564 (N_20564,N_19941,N_19858);
nor U20565 (N_20565,N_20263,N_19982);
xor U20566 (N_20566,N_20000,N_20011);
or U20567 (N_20567,N_19962,N_19992);
nor U20568 (N_20568,N_19998,N_20328);
and U20569 (N_20569,N_20254,N_20196);
nor U20570 (N_20570,N_19844,N_20129);
and U20571 (N_20571,N_19950,N_20141);
nand U20572 (N_20572,N_20080,N_20375);
or U20573 (N_20573,N_20324,N_20062);
nor U20574 (N_20574,N_19824,N_20167);
nand U20575 (N_20575,N_20268,N_20111);
nand U20576 (N_20576,N_20191,N_19947);
or U20577 (N_20577,N_20202,N_20399);
or U20578 (N_20578,N_19980,N_20061);
nand U20579 (N_20579,N_19802,N_19856);
nand U20580 (N_20580,N_20385,N_19913);
and U20581 (N_20581,N_20155,N_20322);
nand U20582 (N_20582,N_20082,N_19840);
or U20583 (N_20583,N_20233,N_19875);
or U20584 (N_20584,N_19929,N_20176);
and U20585 (N_20585,N_20048,N_20363);
or U20586 (N_20586,N_20074,N_20223);
nand U20587 (N_20587,N_19995,N_20228);
nor U20588 (N_20588,N_19813,N_19989);
or U20589 (N_20589,N_19834,N_20235);
nor U20590 (N_20590,N_19924,N_20200);
nor U20591 (N_20591,N_19860,N_20286);
or U20592 (N_20592,N_20334,N_20068);
and U20593 (N_20593,N_20090,N_20072);
nor U20594 (N_20594,N_20015,N_20193);
or U20595 (N_20595,N_20347,N_20188);
nor U20596 (N_20596,N_20154,N_19890);
xor U20597 (N_20597,N_19972,N_19951);
and U20598 (N_20598,N_20372,N_20194);
and U20599 (N_20599,N_20243,N_20139);
nor U20600 (N_20600,N_20229,N_20308);
and U20601 (N_20601,N_20095,N_20022);
nor U20602 (N_20602,N_20227,N_20138);
and U20603 (N_20603,N_20014,N_20189);
or U20604 (N_20604,N_19975,N_20319);
nand U20605 (N_20605,N_20250,N_19838);
and U20606 (N_20606,N_19826,N_20294);
xor U20607 (N_20607,N_19958,N_20258);
and U20608 (N_20608,N_19926,N_20077);
or U20609 (N_20609,N_20288,N_20003);
nand U20610 (N_20610,N_20115,N_19835);
or U20611 (N_20611,N_20178,N_19923);
or U20612 (N_20612,N_20332,N_20221);
xor U20613 (N_20613,N_19928,N_20366);
and U20614 (N_20614,N_20244,N_20171);
or U20615 (N_20615,N_19852,N_19987);
or U20616 (N_20616,N_20169,N_19842);
and U20617 (N_20617,N_20338,N_19874);
or U20618 (N_20618,N_20382,N_19905);
and U20619 (N_20619,N_20207,N_20218);
nor U20620 (N_20620,N_20232,N_20255);
and U20621 (N_20621,N_20076,N_19919);
nor U20622 (N_20622,N_19866,N_20261);
nor U20623 (N_20623,N_20290,N_20351);
or U20624 (N_20624,N_20295,N_19847);
nor U20625 (N_20625,N_20222,N_20133);
nand U20626 (N_20626,N_20282,N_19821);
or U20627 (N_20627,N_20320,N_19818);
and U20628 (N_20628,N_19801,N_20157);
or U20629 (N_20629,N_20265,N_20050);
nand U20630 (N_20630,N_20236,N_19839);
or U20631 (N_20631,N_20356,N_19974);
nand U20632 (N_20632,N_20002,N_20106);
nand U20633 (N_20633,N_20388,N_20166);
nand U20634 (N_20634,N_19976,N_19944);
or U20635 (N_20635,N_19816,N_20126);
nand U20636 (N_20636,N_20007,N_20231);
xnor U20637 (N_20637,N_20238,N_20122);
and U20638 (N_20638,N_19986,N_20192);
nor U20639 (N_20639,N_20170,N_20148);
nor U20640 (N_20640,N_20033,N_20187);
nor U20641 (N_20641,N_20367,N_20042);
and U20642 (N_20642,N_19970,N_20340);
and U20643 (N_20643,N_20237,N_19906);
and U20644 (N_20644,N_20131,N_20186);
nand U20645 (N_20645,N_20378,N_19967);
and U20646 (N_20646,N_20314,N_19979);
or U20647 (N_20647,N_20177,N_19990);
and U20648 (N_20648,N_20081,N_20150);
or U20649 (N_20649,N_20034,N_20213);
and U20650 (N_20650,N_20325,N_20185);
or U20651 (N_20651,N_20118,N_19837);
and U20652 (N_20652,N_20017,N_19965);
nor U20653 (N_20653,N_19895,N_20277);
or U20654 (N_20654,N_19983,N_20359);
or U20655 (N_20655,N_19960,N_19901);
nor U20656 (N_20656,N_20112,N_20018);
and U20657 (N_20657,N_19910,N_19848);
nand U20658 (N_20658,N_19900,N_20024);
and U20659 (N_20659,N_20159,N_20096);
nor U20660 (N_20660,N_20397,N_19927);
and U20661 (N_20661,N_19843,N_20013);
and U20662 (N_20662,N_20035,N_19945);
xnor U20663 (N_20663,N_20210,N_20220);
or U20664 (N_20664,N_20165,N_19904);
nor U20665 (N_20665,N_19850,N_19829);
and U20666 (N_20666,N_20054,N_20130);
nand U20667 (N_20667,N_20326,N_20396);
and U20668 (N_20668,N_20259,N_19899);
nand U20669 (N_20669,N_19881,N_19991);
nor U20670 (N_20670,N_20010,N_19878);
nor U20671 (N_20671,N_20100,N_20323);
nand U20672 (N_20672,N_19873,N_20173);
nor U20673 (N_20673,N_20226,N_19836);
nand U20674 (N_20674,N_20211,N_20270);
or U20675 (N_20675,N_20358,N_19862);
nor U20676 (N_20676,N_19918,N_19936);
nor U20677 (N_20677,N_20053,N_19831);
nand U20678 (N_20678,N_20301,N_20041);
nor U20679 (N_20679,N_20343,N_20109);
nor U20680 (N_20680,N_20394,N_19969);
xor U20681 (N_20681,N_20205,N_19854);
nor U20682 (N_20682,N_20190,N_20174);
or U20683 (N_20683,N_20287,N_19868);
or U20684 (N_20684,N_20327,N_20302);
and U20685 (N_20685,N_20164,N_20065);
and U20686 (N_20686,N_20289,N_19864);
nand U20687 (N_20687,N_20296,N_20350);
or U20688 (N_20688,N_20331,N_20008);
nor U20689 (N_20689,N_19914,N_20330);
and U20690 (N_20690,N_19933,N_19815);
nor U20691 (N_20691,N_19903,N_20389);
or U20692 (N_20692,N_20028,N_19822);
or U20693 (N_20693,N_19872,N_19807);
nand U20694 (N_20694,N_20140,N_20144);
nand U20695 (N_20695,N_19984,N_20239);
nand U20696 (N_20696,N_20281,N_19939);
nor U20697 (N_20697,N_20342,N_20172);
nor U20698 (N_20698,N_19996,N_19925);
nor U20699 (N_20699,N_20117,N_20070);
nor U20700 (N_20700,N_20344,N_20216);
and U20701 (N_20701,N_20192,N_19939);
or U20702 (N_20702,N_20240,N_20133);
nand U20703 (N_20703,N_20150,N_19870);
nand U20704 (N_20704,N_19976,N_20090);
and U20705 (N_20705,N_20140,N_20118);
nor U20706 (N_20706,N_19985,N_20283);
and U20707 (N_20707,N_20037,N_19997);
nor U20708 (N_20708,N_20196,N_20040);
or U20709 (N_20709,N_20353,N_20055);
or U20710 (N_20710,N_20332,N_19955);
or U20711 (N_20711,N_20153,N_19811);
nor U20712 (N_20712,N_20167,N_20098);
and U20713 (N_20713,N_19834,N_20108);
and U20714 (N_20714,N_20318,N_20205);
or U20715 (N_20715,N_19905,N_20311);
and U20716 (N_20716,N_20135,N_19902);
nor U20717 (N_20717,N_20236,N_20104);
nor U20718 (N_20718,N_19887,N_20062);
nor U20719 (N_20719,N_19911,N_20255);
nor U20720 (N_20720,N_19965,N_20024);
nor U20721 (N_20721,N_20181,N_19980);
xor U20722 (N_20722,N_19823,N_20031);
xor U20723 (N_20723,N_20311,N_19906);
xnor U20724 (N_20724,N_20394,N_19835);
nand U20725 (N_20725,N_19965,N_19871);
nor U20726 (N_20726,N_20017,N_19969);
or U20727 (N_20727,N_20282,N_20325);
nand U20728 (N_20728,N_20127,N_20241);
nor U20729 (N_20729,N_20099,N_20106);
or U20730 (N_20730,N_20148,N_19996);
nand U20731 (N_20731,N_20223,N_20258);
nand U20732 (N_20732,N_19896,N_19987);
and U20733 (N_20733,N_20019,N_20243);
nand U20734 (N_20734,N_20125,N_20123);
or U20735 (N_20735,N_19847,N_19924);
nor U20736 (N_20736,N_20218,N_19846);
nand U20737 (N_20737,N_19948,N_20146);
nand U20738 (N_20738,N_19995,N_19914);
nand U20739 (N_20739,N_20106,N_20143);
nand U20740 (N_20740,N_20273,N_19957);
or U20741 (N_20741,N_20041,N_19906);
or U20742 (N_20742,N_20395,N_20324);
nand U20743 (N_20743,N_19893,N_20231);
or U20744 (N_20744,N_19945,N_20295);
or U20745 (N_20745,N_19869,N_19824);
nand U20746 (N_20746,N_19849,N_20208);
or U20747 (N_20747,N_20029,N_20093);
nor U20748 (N_20748,N_19879,N_19914);
and U20749 (N_20749,N_19990,N_20193);
nor U20750 (N_20750,N_20015,N_19958);
nor U20751 (N_20751,N_20317,N_19819);
or U20752 (N_20752,N_19901,N_19882);
or U20753 (N_20753,N_19814,N_19974);
or U20754 (N_20754,N_20277,N_19988);
or U20755 (N_20755,N_20304,N_20371);
xor U20756 (N_20756,N_20301,N_20352);
nand U20757 (N_20757,N_20160,N_19889);
or U20758 (N_20758,N_20314,N_19868);
and U20759 (N_20759,N_20045,N_19828);
nand U20760 (N_20760,N_20271,N_20296);
xor U20761 (N_20761,N_19869,N_20109);
nand U20762 (N_20762,N_19974,N_20319);
nand U20763 (N_20763,N_20258,N_20236);
and U20764 (N_20764,N_19844,N_19872);
and U20765 (N_20765,N_20244,N_19893);
or U20766 (N_20766,N_20212,N_20015);
nand U20767 (N_20767,N_19886,N_20060);
nand U20768 (N_20768,N_19990,N_20380);
and U20769 (N_20769,N_20227,N_20062);
nand U20770 (N_20770,N_20188,N_20125);
and U20771 (N_20771,N_20165,N_20014);
nand U20772 (N_20772,N_20200,N_20188);
or U20773 (N_20773,N_20116,N_20318);
nand U20774 (N_20774,N_20136,N_20209);
nor U20775 (N_20775,N_19907,N_20128);
or U20776 (N_20776,N_20355,N_20162);
nand U20777 (N_20777,N_19922,N_20127);
and U20778 (N_20778,N_19904,N_20327);
and U20779 (N_20779,N_20353,N_19817);
nor U20780 (N_20780,N_19891,N_19999);
or U20781 (N_20781,N_20252,N_20274);
nor U20782 (N_20782,N_20337,N_19875);
nand U20783 (N_20783,N_20343,N_19841);
or U20784 (N_20784,N_20355,N_20022);
or U20785 (N_20785,N_20132,N_19983);
and U20786 (N_20786,N_20072,N_20240);
xnor U20787 (N_20787,N_20355,N_20178);
and U20788 (N_20788,N_19936,N_20290);
xnor U20789 (N_20789,N_20022,N_19864);
and U20790 (N_20790,N_20227,N_19872);
and U20791 (N_20791,N_20122,N_19965);
or U20792 (N_20792,N_19905,N_19981);
or U20793 (N_20793,N_20143,N_20362);
and U20794 (N_20794,N_20058,N_20390);
or U20795 (N_20795,N_20143,N_19838);
and U20796 (N_20796,N_19832,N_19882);
nor U20797 (N_20797,N_20300,N_19965);
and U20798 (N_20798,N_20092,N_19915);
or U20799 (N_20799,N_20171,N_20106);
xnor U20800 (N_20800,N_19899,N_20264);
nand U20801 (N_20801,N_20076,N_20303);
nand U20802 (N_20802,N_19903,N_20200);
or U20803 (N_20803,N_20339,N_19986);
xor U20804 (N_20804,N_20094,N_19872);
or U20805 (N_20805,N_20374,N_20352);
nor U20806 (N_20806,N_19852,N_20346);
and U20807 (N_20807,N_19940,N_20211);
or U20808 (N_20808,N_19849,N_20240);
or U20809 (N_20809,N_20358,N_20154);
or U20810 (N_20810,N_20079,N_19991);
nor U20811 (N_20811,N_19955,N_19995);
nand U20812 (N_20812,N_19967,N_19849);
nor U20813 (N_20813,N_20349,N_20237);
nand U20814 (N_20814,N_19935,N_20172);
and U20815 (N_20815,N_20051,N_20181);
nand U20816 (N_20816,N_20389,N_20238);
xnor U20817 (N_20817,N_19861,N_20265);
and U20818 (N_20818,N_20056,N_20231);
or U20819 (N_20819,N_20049,N_20304);
or U20820 (N_20820,N_20260,N_20096);
or U20821 (N_20821,N_20195,N_20369);
nor U20822 (N_20822,N_20061,N_20248);
and U20823 (N_20823,N_19858,N_20347);
or U20824 (N_20824,N_19822,N_19946);
nand U20825 (N_20825,N_19870,N_20359);
nor U20826 (N_20826,N_20010,N_19858);
xnor U20827 (N_20827,N_20330,N_20283);
and U20828 (N_20828,N_20154,N_20335);
xnor U20829 (N_20829,N_19845,N_19940);
or U20830 (N_20830,N_19952,N_19810);
nor U20831 (N_20831,N_20245,N_20186);
nand U20832 (N_20832,N_19939,N_20223);
nand U20833 (N_20833,N_20348,N_20351);
nor U20834 (N_20834,N_20082,N_19922);
xnor U20835 (N_20835,N_19822,N_19889);
nand U20836 (N_20836,N_20393,N_20069);
and U20837 (N_20837,N_19935,N_19804);
and U20838 (N_20838,N_19988,N_20347);
or U20839 (N_20839,N_20027,N_19855);
nor U20840 (N_20840,N_19855,N_20399);
or U20841 (N_20841,N_20377,N_20352);
nor U20842 (N_20842,N_20137,N_20099);
nand U20843 (N_20843,N_20188,N_20012);
or U20844 (N_20844,N_19988,N_20005);
nor U20845 (N_20845,N_20392,N_20224);
and U20846 (N_20846,N_19979,N_20131);
nand U20847 (N_20847,N_20129,N_20367);
and U20848 (N_20848,N_19968,N_20055);
nand U20849 (N_20849,N_19952,N_19826);
nand U20850 (N_20850,N_20031,N_19800);
nor U20851 (N_20851,N_20046,N_20165);
or U20852 (N_20852,N_20088,N_20162);
and U20853 (N_20853,N_19801,N_20031);
nor U20854 (N_20854,N_19844,N_19895);
nand U20855 (N_20855,N_20394,N_19937);
nor U20856 (N_20856,N_20298,N_20114);
nand U20857 (N_20857,N_19944,N_20310);
nor U20858 (N_20858,N_20324,N_20368);
nor U20859 (N_20859,N_20012,N_20277);
and U20860 (N_20860,N_19974,N_19820);
or U20861 (N_20861,N_19934,N_19995);
and U20862 (N_20862,N_19847,N_20242);
nor U20863 (N_20863,N_20090,N_20238);
or U20864 (N_20864,N_20275,N_20136);
nand U20865 (N_20865,N_20090,N_20252);
nand U20866 (N_20866,N_19897,N_20162);
or U20867 (N_20867,N_20044,N_19935);
nand U20868 (N_20868,N_20388,N_19801);
or U20869 (N_20869,N_20279,N_20010);
or U20870 (N_20870,N_20167,N_20124);
and U20871 (N_20871,N_20050,N_20074);
and U20872 (N_20872,N_19912,N_20286);
nor U20873 (N_20873,N_20326,N_19977);
nand U20874 (N_20874,N_19931,N_20161);
nand U20875 (N_20875,N_20124,N_19802);
and U20876 (N_20876,N_19852,N_20041);
or U20877 (N_20877,N_20361,N_20220);
or U20878 (N_20878,N_20279,N_19841);
xnor U20879 (N_20879,N_20342,N_19985);
nand U20880 (N_20880,N_20286,N_19983);
and U20881 (N_20881,N_20256,N_19924);
or U20882 (N_20882,N_20050,N_19807);
nand U20883 (N_20883,N_20146,N_19812);
nor U20884 (N_20884,N_20300,N_20108);
nand U20885 (N_20885,N_20016,N_19829);
nor U20886 (N_20886,N_20137,N_19978);
nand U20887 (N_20887,N_20308,N_20118);
or U20888 (N_20888,N_20185,N_19947);
nor U20889 (N_20889,N_20361,N_20157);
nand U20890 (N_20890,N_20245,N_20116);
or U20891 (N_20891,N_20330,N_20359);
nor U20892 (N_20892,N_20076,N_20236);
or U20893 (N_20893,N_20294,N_19926);
nor U20894 (N_20894,N_20331,N_20125);
xor U20895 (N_20895,N_19925,N_20317);
xor U20896 (N_20896,N_20309,N_20185);
or U20897 (N_20897,N_20094,N_20293);
nand U20898 (N_20898,N_19842,N_20392);
nand U20899 (N_20899,N_20119,N_20003);
nor U20900 (N_20900,N_19824,N_20399);
xor U20901 (N_20901,N_19889,N_20075);
xor U20902 (N_20902,N_20084,N_20040);
and U20903 (N_20903,N_20212,N_19815);
nand U20904 (N_20904,N_20355,N_20313);
or U20905 (N_20905,N_19956,N_19918);
or U20906 (N_20906,N_19949,N_19938);
or U20907 (N_20907,N_20299,N_20035);
nand U20908 (N_20908,N_20347,N_20133);
nand U20909 (N_20909,N_20173,N_20220);
and U20910 (N_20910,N_19830,N_20042);
nor U20911 (N_20911,N_20333,N_20207);
nand U20912 (N_20912,N_20229,N_20358);
or U20913 (N_20913,N_20115,N_19868);
nor U20914 (N_20914,N_19952,N_20203);
and U20915 (N_20915,N_20319,N_20342);
nor U20916 (N_20916,N_20246,N_19964);
nor U20917 (N_20917,N_19880,N_19816);
and U20918 (N_20918,N_20200,N_20083);
nor U20919 (N_20919,N_20030,N_20170);
xnor U20920 (N_20920,N_20209,N_20244);
nor U20921 (N_20921,N_19850,N_20153);
nand U20922 (N_20922,N_19803,N_20005);
nor U20923 (N_20923,N_20134,N_20213);
and U20924 (N_20924,N_20162,N_19948);
and U20925 (N_20925,N_20193,N_20291);
or U20926 (N_20926,N_20148,N_19928);
nand U20927 (N_20927,N_20062,N_20302);
or U20928 (N_20928,N_20095,N_20306);
nand U20929 (N_20929,N_20305,N_19904);
nor U20930 (N_20930,N_20158,N_20356);
nor U20931 (N_20931,N_20127,N_20099);
or U20932 (N_20932,N_19942,N_20052);
xnor U20933 (N_20933,N_20324,N_20263);
or U20934 (N_20934,N_19982,N_19895);
nand U20935 (N_20935,N_20231,N_19967);
nand U20936 (N_20936,N_20108,N_20221);
nand U20937 (N_20937,N_19917,N_20254);
and U20938 (N_20938,N_20130,N_20026);
or U20939 (N_20939,N_20312,N_20148);
and U20940 (N_20940,N_20266,N_19912);
and U20941 (N_20941,N_20012,N_19911);
or U20942 (N_20942,N_19999,N_20135);
nor U20943 (N_20943,N_20357,N_20383);
or U20944 (N_20944,N_19915,N_19921);
nand U20945 (N_20945,N_20035,N_20098);
nor U20946 (N_20946,N_20027,N_19808);
nor U20947 (N_20947,N_20180,N_19944);
or U20948 (N_20948,N_19982,N_19856);
nor U20949 (N_20949,N_20169,N_20266);
and U20950 (N_20950,N_20344,N_20059);
nand U20951 (N_20951,N_20021,N_20078);
nand U20952 (N_20952,N_20080,N_20277);
or U20953 (N_20953,N_20216,N_20127);
and U20954 (N_20954,N_20048,N_20196);
nand U20955 (N_20955,N_20335,N_19907);
or U20956 (N_20956,N_19861,N_20236);
nand U20957 (N_20957,N_19858,N_20142);
and U20958 (N_20958,N_20355,N_20005);
or U20959 (N_20959,N_20161,N_20329);
or U20960 (N_20960,N_20029,N_20282);
nor U20961 (N_20961,N_19853,N_19822);
or U20962 (N_20962,N_19914,N_20308);
nor U20963 (N_20963,N_20227,N_20347);
or U20964 (N_20964,N_20304,N_19992);
nor U20965 (N_20965,N_19872,N_20278);
and U20966 (N_20966,N_20008,N_20171);
nand U20967 (N_20967,N_19879,N_20028);
and U20968 (N_20968,N_20320,N_20390);
nand U20969 (N_20969,N_20024,N_19932);
and U20970 (N_20970,N_20349,N_19870);
and U20971 (N_20971,N_20190,N_20178);
or U20972 (N_20972,N_19912,N_19857);
nor U20973 (N_20973,N_20091,N_19926);
nor U20974 (N_20974,N_19878,N_20161);
nor U20975 (N_20975,N_20244,N_20081);
or U20976 (N_20976,N_19831,N_20282);
or U20977 (N_20977,N_19935,N_19969);
nor U20978 (N_20978,N_19922,N_20212);
or U20979 (N_20979,N_20387,N_20099);
nor U20980 (N_20980,N_20045,N_20150);
xor U20981 (N_20981,N_19885,N_20352);
xnor U20982 (N_20982,N_20328,N_20145);
and U20983 (N_20983,N_20236,N_20124);
nand U20984 (N_20984,N_20063,N_19936);
nand U20985 (N_20985,N_20012,N_20112);
or U20986 (N_20986,N_20055,N_20163);
or U20987 (N_20987,N_19894,N_20398);
and U20988 (N_20988,N_20137,N_20214);
xnor U20989 (N_20989,N_20087,N_19801);
and U20990 (N_20990,N_19913,N_20002);
nand U20991 (N_20991,N_19849,N_20004);
nor U20992 (N_20992,N_20115,N_20288);
and U20993 (N_20993,N_20312,N_20157);
nor U20994 (N_20994,N_19908,N_20269);
and U20995 (N_20995,N_19878,N_20061);
or U20996 (N_20996,N_20353,N_19942);
and U20997 (N_20997,N_20198,N_20003);
and U20998 (N_20998,N_19810,N_20171);
and U20999 (N_20999,N_20198,N_20177);
and U21000 (N_21000,N_20747,N_20662);
xnor U21001 (N_21001,N_20986,N_20442);
nand U21002 (N_21002,N_20431,N_20456);
nand U21003 (N_21003,N_20851,N_20952);
and U21004 (N_21004,N_20542,N_20424);
and U21005 (N_21005,N_20945,N_20719);
and U21006 (N_21006,N_20489,N_20811);
nand U21007 (N_21007,N_20509,N_20537);
or U21008 (N_21008,N_20436,N_20650);
or U21009 (N_21009,N_20631,N_20990);
and U21010 (N_21010,N_20755,N_20754);
nor U21011 (N_21011,N_20702,N_20464);
nand U21012 (N_21012,N_20477,N_20948);
nor U21013 (N_21013,N_20902,N_20828);
and U21014 (N_21014,N_20482,N_20421);
or U21015 (N_21015,N_20790,N_20830);
nor U21016 (N_21016,N_20739,N_20705);
or U21017 (N_21017,N_20645,N_20784);
xor U21018 (N_21018,N_20471,N_20582);
nor U21019 (N_21019,N_20565,N_20765);
nor U21020 (N_21020,N_20411,N_20614);
nor U21021 (N_21021,N_20865,N_20561);
or U21022 (N_21022,N_20776,N_20629);
or U21023 (N_21023,N_20655,N_20801);
nand U21024 (N_21024,N_20647,N_20571);
and U21025 (N_21025,N_20736,N_20906);
or U21026 (N_21026,N_20832,N_20467);
nor U21027 (N_21027,N_20932,N_20954);
or U21028 (N_21028,N_20416,N_20665);
and U21029 (N_21029,N_20810,N_20951);
or U21030 (N_21030,N_20453,N_20463);
nor U21031 (N_21031,N_20995,N_20429);
nor U21032 (N_21032,N_20921,N_20827);
nor U21033 (N_21033,N_20993,N_20982);
and U21034 (N_21034,N_20568,N_20533);
and U21035 (N_21035,N_20481,N_20679);
or U21036 (N_21036,N_20891,N_20675);
nand U21037 (N_21037,N_20888,N_20532);
and U21038 (N_21038,N_20751,N_20806);
nand U21039 (N_21039,N_20446,N_20953);
nand U21040 (N_21040,N_20732,N_20998);
or U21041 (N_21041,N_20819,N_20860);
nand U21042 (N_21042,N_20435,N_20441);
nand U21043 (N_21043,N_20781,N_20761);
nor U21044 (N_21044,N_20600,N_20404);
or U21045 (N_21045,N_20630,N_20844);
nor U21046 (N_21046,N_20486,N_20749);
and U21047 (N_21047,N_20558,N_20717);
xnor U21048 (N_21048,N_20454,N_20997);
nor U21049 (N_21049,N_20974,N_20822);
and U21050 (N_21050,N_20449,N_20625);
and U21051 (N_21051,N_20835,N_20624);
and U21052 (N_21052,N_20651,N_20556);
xnor U21053 (N_21053,N_20599,N_20996);
nor U21054 (N_21054,N_20636,N_20417);
xnor U21055 (N_21055,N_20957,N_20856);
nand U21056 (N_21056,N_20593,N_20607);
or U21057 (N_21057,N_20913,N_20892);
or U21058 (N_21058,N_20712,N_20681);
and U21059 (N_21059,N_20465,N_20748);
nor U21060 (N_21060,N_20545,N_20949);
and U21061 (N_21061,N_20973,N_20531);
xor U21062 (N_21062,N_20871,N_20422);
nor U21063 (N_21063,N_20583,N_20713);
nor U21064 (N_21064,N_20783,N_20491);
or U21065 (N_21065,N_20563,N_20846);
and U21066 (N_21066,N_20508,N_20552);
nor U21067 (N_21067,N_20518,N_20799);
nand U21068 (N_21068,N_20878,N_20672);
and U21069 (N_21069,N_20883,N_20723);
or U21070 (N_21070,N_20470,N_20769);
and U21071 (N_21071,N_20406,N_20578);
nand U21072 (N_21072,N_20512,N_20743);
and U21073 (N_21073,N_20646,N_20648);
nand U21074 (N_21074,N_20617,N_20428);
nand U21075 (N_21075,N_20787,N_20847);
nor U21076 (N_21076,N_20956,N_20658);
nand U21077 (N_21077,N_20480,N_20613);
nor U21078 (N_21078,N_20849,N_20757);
nand U21079 (N_21079,N_20548,N_20495);
and U21080 (N_21080,N_20938,N_20912);
and U21081 (N_21081,N_20425,N_20698);
nand U21082 (N_21082,N_20929,N_20966);
xor U21083 (N_21083,N_20895,N_20668);
xnor U21084 (N_21084,N_20696,N_20426);
or U21085 (N_21085,N_20772,N_20598);
nor U21086 (N_21086,N_20610,N_20553);
or U21087 (N_21087,N_20848,N_20701);
xor U21088 (N_21088,N_20971,N_20451);
nor U21089 (N_21089,N_20573,N_20700);
or U21090 (N_21090,N_20487,N_20958);
nand U21091 (N_21091,N_20817,N_20760);
or U21092 (N_21092,N_20695,N_20460);
nand U21093 (N_21093,N_20643,N_20918);
nor U21094 (N_21094,N_20969,N_20816);
or U21095 (N_21095,N_20709,N_20619);
or U21096 (N_21096,N_20408,N_20722);
nor U21097 (N_21097,N_20814,N_20965);
and U21098 (N_21098,N_20959,N_20853);
nor U21099 (N_21099,N_20526,N_20850);
nor U21100 (N_21100,N_20889,N_20666);
nor U21101 (N_21101,N_20885,N_20445);
nor U21102 (N_21102,N_20841,N_20621);
xnor U21103 (N_21103,N_20922,N_20462);
and U21104 (N_21104,N_20649,N_20942);
nor U21105 (N_21105,N_20882,N_20720);
and U21106 (N_21106,N_20673,N_20551);
xor U21107 (N_21107,N_20438,N_20502);
xor U21108 (N_21108,N_20916,N_20862);
nand U21109 (N_21109,N_20443,N_20601);
or U21110 (N_21110,N_20768,N_20724);
nor U21111 (N_21111,N_20901,N_20867);
or U21112 (N_21112,N_20911,N_20575);
nor U21113 (N_21113,N_20522,N_20845);
or U21114 (N_21114,N_20415,N_20880);
nor U21115 (N_21115,N_20762,N_20633);
and U21116 (N_21116,N_20729,N_20444);
nand U21117 (N_21117,N_20763,N_20523);
nor U21118 (N_21118,N_20457,N_20881);
and U21119 (N_21119,N_20690,N_20989);
or U21120 (N_21120,N_20511,N_20710);
nor U21121 (N_21121,N_20670,N_20984);
or U21122 (N_21122,N_20602,N_20715);
nor U21123 (N_21123,N_20500,N_20574);
or U21124 (N_21124,N_20992,N_20669);
nand U21125 (N_21125,N_20854,N_20788);
and U21126 (N_21126,N_20838,N_20976);
xor U21127 (N_21127,N_20584,N_20725);
or U21128 (N_21128,N_20866,N_20678);
and U21129 (N_21129,N_20595,N_20940);
or U21130 (N_21130,N_20872,N_20525);
nand U21131 (N_21131,N_20664,N_20490);
nand U21132 (N_21132,N_20773,N_20660);
or U21133 (N_21133,N_20927,N_20461);
or U21134 (N_21134,N_20592,N_20766);
xor U21135 (N_21135,N_20753,N_20496);
xor U21136 (N_21136,N_20661,N_20475);
xor U21137 (N_21137,N_20873,N_20430);
nor U21138 (N_21138,N_20688,N_20855);
and U21139 (N_21139,N_20492,N_20620);
nor U21140 (N_21140,N_20612,N_20737);
xor U21141 (N_21141,N_20652,N_20469);
nor U21142 (N_21142,N_20962,N_20896);
nand U21143 (N_21143,N_20586,N_20797);
xnor U21144 (N_21144,N_20994,N_20964);
nand U21145 (N_21145,N_20777,N_20857);
or U21146 (N_21146,N_20539,N_20405);
nand U21147 (N_21147,N_20978,N_20697);
nor U21148 (N_21148,N_20423,N_20946);
nand U21149 (N_21149,N_20779,N_20653);
nand U21150 (N_21150,N_20980,N_20899);
and U21151 (N_21151,N_20618,N_20909);
or U21152 (N_21152,N_20473,N_20514);
or U21153 (N_21153,N_20409,N_20778);
and U21154 (N_21154,N_20884,N_20711);
and U21155 (N_21155,N_20528,N_20597);
and U21156 (N_21156,N_20517,N_20904);
nand U21157 (N_21157,N_20917,N_20616);
and U21158 (N_21158,N_20581,N_20930);
nand U21159 (N_21159,N_20770,N_20876);
xor U21160 (N_21160,N_20824,N_20432);
and U21161 (N_21161,N_20931,N_20924);
and U21162 (N_21162,N_20691,N_20935);
nor U21163 (N_21163,N_20628,N_20606);
nor U21164 (N_21164,N_20401,N_20434);
nor U21165 (N_21165,N_20740,N_20547);
and U21166 (N_21166,N_20983,N_20928);
and U21167 (N_21167,N_20452,N_20756);
nor U21168 (N_21168,N_20676,N_20639);
nor U21169 (N_21169,N_20572,N_20659);
and U21170 (N_21170,N_20791,N_20546);
nor U21171 (N_21171,N_20923,N_20991);
nand U21172 (N_21172,N_20507,N_20569);
or U21173 (N_21173,N_20903,N_20437);
nor U21174 (N_21174,N_20900,N_20591);
or U21175 (N_21175,N_20728,N_20905);
xnor U21176 (N_21176,N_20577,N_20708);
nor U21177 (N_21177,N_20550,N_20513);
or U21178 (N_21178,N_20963,N_20663);
and U21179 (N_21179,N_20609,N_20837);
nand U21180 (N_21180,N_20447,N_20590);
xnor U21181 (N_21181,N_20742,N_20979);
and U21182 (N_21182,N_20735,N_20967);
nand U21183 (N_21183,N_20466,N_20680);
nand U21184 (N_21184,N_20887,N_20535);
nand U21185 (N_21185,N_20524,N_20479);
xor U21186 (N_21186,N_20975,N_20716);
or U21187 (N_21187,N_20472,N_20782);
or U21188 (N_21188,N_20414,N_20746);
and U21189 (N_21189,N_20557,N_20641);
xor U21190 (N_21190,N_20834,N_20852);
nand U21191 (N_21191,N_20585,N_20530);
nand U21192 (N_21192,N_20950,N_20455);
nand U21193 (N_21193,N_20527,N_20807);
nand U21194 (N_21194,N_20407,N_20603);
or U21195 (N_21195,N_20505,N_20412);
or U21196 (N_21196,N_20506,N_20587);
nand U21197 (N_21197,N_20792,N_20682);
nand U21198 (N_21198,N_20886,N_20985);
nor U21199 (N_21199,N_20877,N_20693);
and U21200 (N_21200,N_20501,N_20632);
nand U21201 (N_21201,N_20879,N_20622);
nand U21202 (N_21202,N_20972,N_20638);
or U21203 (N_21203,N_20934,N_20448);
nor U21204 (N_21204,N_20427,N_20555);
nor U21205 (N_21205,N_20543,N_20780);
or U21206 (N_21206,N_20988,N_20786);
or U21207 (N_21207,N_20968,N_20483);
nor U21208 (N_21208,N_20821,N_20744);
nand U21209 (N_21209,N_20499,N_20589);
or U21210 (N_21210,N_20802,N_20920);
and U21211 (N_21211,N_20840,N_20440);
nor U21212 (N_21212,N_20775,N_20741);
nor U21213 (N_21213,N_20726,N_20861);
or U21214 (N_21214,N_20604,N_20800);
and U21215 (N_21215,N_20692,N_20510);
and U21216 (N_21216,N_20529,N_20468);
or U21217 (N_21217,N_20833,N_20699);
nor U21218 (N_21218,N_20497,N_20541);
nor U21219 (N_21219,N_20594,N_20981);
nor U21220 (N_21220,N_20567,N_20640);
nor U21221 (N_21221,N_20794,N_20493);
and U21222 (N_21222,N_20798,N_20635);
or U21223 (N_21223,N_20733,N_20667);
and U21224 (N_21224,N_20826,N_20829);
nand U21225 (N_21225,N_20890,N_20521);
and U21226 (N_21226,N_20403,N_20562);
and U21227 (N_21227,N_20897,N_20674);
xor U21228 (N_21228,N_20818,N_20752);
nor U21229 (N_21229,N_20485,N_20869);
and U21230 (N_21230,N_20413,N_20843);
nand U21231 (N_21231,N_20605,N_20987);
xor U21232 (N_21232,N_20842,N_20559);
or U21233 (N_21233,N_20694,N_20925);
nor U21234 (N_21234,N_20803,N_20704);
or U21235 (N_21235,N_20870,N_20868);
or U21236 (N_21236,N_20795,N_20433);
nor U21237 (N_21237,N_20671,N_20476);
or U21238 (N_21238,N_20936,N_20478);
nand U21239 (N_21239,N_20734,N_20402);
or U21240 (N_21240,N_20893,N_20623);
nor U21241 (N_21241,N_20937,N_20683);
nor U21242 (N_21242,N_20961,N_20588);
and U21243 (N_21243,N_20805,N_20596);
nand U21244 (N_21244,N_20774,N_20793);
and U21245 (N_21245,N_20544,N_20439);
nor U21246 (N_21246,N_20566,N_20560);
or U21247 (N_21247,N_20789,N_20764);
nor U21248 (N_21248,N_20767,N_20474);
or U21249 (N_21249,N_20960,N_20808);
and U21250 (N_21250,N_20536,N_20504);
and U21251 (N_21251,N_20898,N_20919);
nand U21252 (N_21252,N_20944,N_20874);
nand U21253 (N_21253,N_20970,N_20564);
and U21254 (N_21254,N_20684,N_20771);
nand U21255 (N_21255,N_20947,N_20656);
nor U21256 (N_21256,N_20745,N_20540);
and U21257 (N_21257,N_20707,N_20627);
nor U21258 (N_21258,N_20731,N_20579);
and U21259 (N_21259,N_20894,N_20863);
nor U21260 (N_21260,N_20907,N_20815);
and U21261 (N_21261,N_20644,N_20450);
nor U21262 (N_21262,N_20812,N_20459);
nor U21263 (N_21263,N_20839,N_20941);
nand U21264 (N_21264,N_20516,N_20858);
and U21265 (N_21265,N_20910,N_20831);
nor U21266 (N_21266,N_20418,N_20915);
nor U21267 (N_21267,N_20519,N_20549);
nor U21268 (N_21268,N_20820,N_20538);
or U21269 (N_21269,N_20706,N_20657);
or U21270 (N_21270,N_20750,N_20685);
nand U21271 (N_21271,N_20554,N_20721);
nor U21272 (N_21272,N_20933,N_20943);
nand U21273 (N_21273,N_20634,N_20498);
or U21274 (N_21274,N_20836,N_20914);
or U21275 (N_21275,N_20759,N_20611);
nor U21276 (N_21276,N_20703,N_20615);
nor U21277 (N_21277,N_20400,N_20608);
or U21278 (N_21278,N_20730,N_20520);
nor U21279 (N_21279,N_20687,N_20727);
nor U21280 (N_21280,N_20570,N_20738);
and U21281 (N_21281,N_20809,N_20458);
nor U21282 (N_21282,N_20823,N_20908);
nand U21283 (N_21283,N_20939,N_20686);
or U21284 (N_21284,N_20714,N_20875);
and U21285 (N_21285,N_20503,N_20642);
nand U21286 (N_21286,N_20813,N_20419);
nor U21287 (N_21287,N_20955,N_20410);
nand U21288 (N_21288,N_20977,N_20864);
nor U21289 (N_21289,N_20758,N_20677);
or U21290 (N_21290,N_20488,N_20926);
nand U21291 (N_21291,N_20580,N_20804);
or U21292 (N_21292,N_20637,N_20796);
nor U21293 (N_21293,N_20999,N_20515);
nor U21294 (N_21294,N_20718,N_20825);
nor U21295 (N_21295,N_20420,N_20576);
nand U21296 (N_21296,N_20626,N_20689);
nand U21297 (N_21297,N_20859,N_20654);
xor U21298 (N_21298,N_20484,N_20494);
nand U21299 (N_21299,N_20534,N_20785);
nand U21300 (N_21300,N_20708,N_20975);
or U21301 (N_21301,N_20898,N_20593);
and U21302 (N_21302,N_20852,N_20987);
nor U21303 (N_21303,N_20741,N_20932);
nor U21304 (N_21304,N_20721,N_20419);
and U21305 (N_21305,N_20875,N_20705);
and U21306 (N_21306,N_20623,N_20632);
nand U21307 (N_21307,N_20855,N_20802);
nand U21308 (N_21308,N_20421,N_20828);
nand U21309 (N_21309,N_20612,N_20492);
and U21310 (N_21310,N_20630,N_20763);
or U21311 (N_21311,N_20813,N_20727);
and U21312 (N_21312,N_20750,N_20746);
nor U21313 (N_21313,N_20694,N_20832);
nand U21314 (N_21314,N_20424,N_20622);
nor U21315 (N_21315,N_20454,N_20400);
nand U21316 (N_21316,N_20616,N_20625);
nand U21317 (N_21317,N_20802,N_20799);
nand U21318 (N_21318,N_20871,N_20469);
nand U21319 (N_21319,N_20586,N_20444);
and U21320 (N_21320,N_20516,N_20771);
or U21321 (N_21321,N_20963,N_20893);
nor U21322 (N_21322,N_20485,N_20949);
and U21323 (N_21323,N_20502,N_20607);
or U21324 (N_21324,N_20607,N_20880);
xnor U21325 (N_21325,N_20948,N_20674);
xor U21326 (N_21326,N_20810,N_20559);
and U21327 (N_21327,N_20721,N_20804);
xnor U21328 (N_21328,N_20620,N_20438);
nand U21329 (N_21329,N_20707,N_20613);
xnor U21330 (N_21330,N_20975,N_20450);
nand U21331 (N_21331,N_20916,N_20713);
or U21332 (N_21332,N_20929,N_20824);
nor U21333 (N_21333,N_20858,N_20662);
and U21334 (N_21334,N_20538,N_20683);
and U21335 (N_21335,N_20831,N_20606);
nand U21336 (N_21336,N_20830,N_20938);
xnor U21337 (N_21337,N_20814,N_20894);
xnor U21338 (N_21338,N_20530,N_20626);
nand U21339 (N_21339,N_20408,N_20997);
nor U21340 (N_21340,N_20690,N_20646);
xnor U21341 (N_21341,N_20581,N_20427);
or U21342 (N_21342,N_20553,N_20745);
and U21343 (N_21343,N_20702,N_20790);
or U21344 (N_21344,N_20918,N_20499);
or U21345 (N_21345,N_20822,N_20944);
nor U21346 (N_21346,N_20790,N_20951);
and U21347 (N_21347,N_20649,N_20789);
or U21348 (N_21348,N_20456,N_20657);
nor U21349 (N_21349,N_20566,N_20775);
or U21350 (N_21350,N_20690,N_20743);
nand U21351 (N_21351,N_20607,N_20925);
xnor U21352 (N_21352,N_20915,N_20545);
nand U21353 (N_21353,N_20847,N_20915);
or U21354 (N_21354,N_20562,N_20849);
nor U21355 (N_21355,N_20836,N_20695);
and U21356 (N_21356,N_20581,N_20548);
and U21357 (N_21357,N_20710,N_20844);
nand U21358 (N_21358,N_20971,N_20692);
and U21359 (N_21359,N_20727,N_20415);
nor U21360 (N_21360,N_20971,N_20645);
nor U21361 (N_21361,N_20427,N_20965);
and U21362 (N_21362,N_20946,N_20440);
or U21363 (N_21363,N_20429,N_20528);
and U21364 (N_21364,N_20783,N_20567);
or U21365 (N_21365,N_20791,N_20410);
nand U21366 (N_21366,N_20456,N_20723);
nor U21367 (N_21367,N_20659,N_20753);
or U21368 (N_21368,N_20698,N_20615);
nand U21369 (N_21369,N_20771,N_20606);
and U21370 (N_21370,N_20756,N_20741);
or U21371 (N_21371,N_20423,N_20400);
or U21372 (N_21372,N_20742,N_20847);
and U21373 (N_21373,N_20781,N_20656);
xor U21374 (N_21374,N_20683,N_20770);
nor U21375 (N_21375,N_20446,N_20501);
nand U21376 (N_21376,N_20866,N_20562);
nor U21377 (N_21377,N_20587,N_20681);
xnor U21378 (N_21378,N_20730,N_20553);
and U21379 (N_21379,N_20509,N_20616);
or U21380 (N_21380,N_20429,N_20758);
nand U21381 (N_21381,N_20706,N_20585);
or U21382 (N_21382,N_20879,N_20988);
nor U21383 (N_21383,N_20813,N_20671);
xor U21384 (N_21384,N_20487,N_20580);
nor U21385 (N_21385,N_20548,N_20865);
nor U21386 (N_21386,N_20682,N_20911);
nand U21387 (N_21387,N_20645,N_20738);
xor U21388 (N_21388,N_20939,N_20929);
nand U21389 (N_21389,N_20760,N_20442);
or U21390 (N_21390,N_20954,N_20664);
and U21391 (N_21391,N_20750,N_20569);
nand U21392 (N_21392,N_20706,N_20566);
and U21393 (N_21393,N_20725,N_20988);
or U21394 (N_21394,N_20481,N_20623);
nor U21395 (N_21395,N_20592,N_20432);
nor U21396 (N_21396,N_20467,N_20535);
nor U21397 (N_21397,N_20732,N_20686);
xor U21398 (N_21398,N_20956,N_20431);
or U21399 (N_21399,N_20680,N_20646);
nand U21400 (N_21400,N_20796,N_20727);
nand U21401 (N_21401,N_20890,N_20535);
xor U21402 (N_21402,N_20820,N_20516);
xor U21403 (N_21403,N_20926,N_20757);
nor U21404 (N_21404,N_20890,N_20534);
nor U21405 (N_21405,N_20527,N_20925);
xnor U21406 (N_21406,N_20795,N_20536);
nand U21407 (N_21407,N_20614,N_20535);
or U21408 (N_21408,N_20452,N_20939);
nor U21409 (N_21409,N_20775,N_20935);
or U21410 (N_21410,N_20610,N_20992);
nor U21411 (N_21411,N_20930,N_20956);
nand U21412 (N_21412,N_20674,N_20782);
nand U21413 (N_21413,N_20629,N_20943);
nor U21414 (N_21414,N_20621,N_20426);
and U21415 (N_21415,N_20586,N_20874);
nor U21416 (N_21416,N_20423,N_20454);
or U21417 (N_21417,N_20975,N_20955);
and U21418 (N_21418,N_20426,N_20688);
nand U21419 (N_21419,N_20696,N_20574);
nand U21420 (N_21420,N_20808,N_20615);
xor U21421 (N_21421,N_20453,N_20920);
xnor U21422 (N_21422,N_20676,N_20918);
and U21423 (N_21423,N_20569,N_20403);
or U21424 (N_21424,N_20597,N_20659);
or U21425 (N_21425,N_20736,N_20800);
and U21426 (N_21426,N_20870,N_20476);
nand U21427 (N_21427,N_20972,N_20891);
nor U21428 (N_21428,N_20774,N_20457);
or U21429 (N_21429,N_20637,N_20456);
or U21430 (N_21430,N_20980,N_20907);
xnor U21431 (N_21431,N_20501,N_20684);
nand U21432 (N_21432,N_20687,N_20814);
nor U21433 (N_21433,N_20447,N_20704);
nor U21434 (N_21434,N_20698,N_20765);
or U21435 (N_21435,N_20566,N_20725);
and U21436 (N_21436,N_20400,N_20926);
nor U21437 (N_21437,N_20975,N_20707);
nor U21438 (N_21438,N_20946,N_20542);
and U21439 (N_21439,N_20868,N_20866);
nand U21440 (N_21440,N_20436,N_20610);
or U21441 (N_21441,N_20411,N_20493);
or U21442 (N_21442,N_20882,N_20523);
nand U21443 (N_21443,N_20403,N_20677);
xor U21444 (N_21444,N_20463,N_20862);
nand U21445 (N_21445,N_20988,N_20983);
xnor U21446 (N_21446,N_20670,N_20488);
xor U21447 (N_21447,N_20822,N_20416);
nand U21448 (N_21448,N_20643,N_20814);
nor U21449 (N_21449,N_20653,N_20588);
or U21450 (N_21450,N_20537,N_20868);
nand U21451 (N_21451,N_20562,N_20437);
nand U21452 (N_21452,N_20469,N_20485);
and U21453 (N_21453,N_20738,N_20940);
or U21454 (N_21454,N_20792,N_20584);
nor U21455 (N_21455,N_20861,N_20945);
nand U21456 (N_21456,N_20802,N_20803);
and U21457 (N_21457,N_20899,N_20435);
nor U21458 (N_21458,N_20812,N_20883);
and U21459 (N_21459,N_20615,N_20512);
nand U21460 (N_21460,N_20896,N_20907);
or U21461 (N_21461,N_20739,N_20485);
xor U21462 (N_21462,N_20625,N_20706);
nand U21463 (N_21463,N_20450,N_20481);
and U21464 (N_21464,N_20636,N_20935);
nor U21465 (N_21465,N_20921,N_20966);
or U21466 (N_21466,N_20904,N_20827);
and U21467 (N_21467,N_20837,N_20664);
or U21468 (N_21468,N_20579,N_20625);
and U21469 (N_21469,N_20526,N_20921);
nand U21470 (N_21470,N_20761,N_20633);
nand U21471 (N_21471,N_20524,N_20939);
and U21472 (N_21472,N_20546,N_20801);
nand U21473 (N_21473,N_20958,N_20426);
xor U21474 (N_21474,N_20903,N_20996);
nor U21475 (N_21475,N_20633,N_20538);
and U21476 (N_21476,N_20614,N_20542);
nand U21477 (N_21477,N_20703,N_20572);
xnor U21478 (N_21478,N_20497,N_20824);
nand U21479 (N_21479,N_20403,N_20735);
or U21480 (N_21480,N_20594,N_20974);
and U21481 (N_21481,N_20675,N_20517);
nand U21482 (N_21482,N_20732,N_20951);
and U21483 (N_21483,N_20889,N_20771);
nor U21484 (N_21484,N_20664,N_20504);
nor U21485 (N_21485,N_20627,N_20700);
or U21486 (N_21486,N_20986,N_20815);
nor U21487 (N_21487,N_20510,N_20823);
or U21488 (N_21488,N_20473,N_20616);
or U21489 (N_21489,N_20499,N_20567);
nor U21490 (N_21490,N_20956,N_20879);
or U21491 (N_21491,N_20511,N_20768);
and U21492 (N_21492,N_20924,N_20927);
nor U21493 (N_21493,N_20481,N_20527);
nand U21494 (N_21494,N_20756,N_20739);
xor U21495 (N_21495,N_20468,N_20970);
and U21496 (N_21496,N_20605,N_20527);
nand U21497 (N_21497,N_20417,N_20870);
nand U21498 (N_21498,N_20451,N_20654);
xnor U21499 (N_21499,N_20901,N_20702);
nor U21500 (N_21500,N_20984,N_20405);
nor U21501 (N_21501,N_20935,N_20951);
nand U21502 (N_21502,N_20993,N_20574);
nand U21503 (N_21503,N_20904,N_20826);
and U21504 (N_21504,N_20807,N_20415);
nand U21505 (N_21505,N_20895,N_20481);
nand U21506 (N_21506,N_20696,N_20500);
and U21507 (N_21507,N_20739,N_20777);
or U21508 (N_21508,N_20794,N_20533);
nand U21509 (N_21509,N_20969,N_20433);
nor U21510 (N_21510,N_20763,N_20898);
xnor U21511 (N_21511,N_20778,N_20736);
nand U21512 (N_21512,N_20629,N_20568);
or U21513 (N_21513,N_20561,N_20698);
nor U21514 (N_21514,N_20667,N_20659);
or U21515 (N_21515,N_20519,N_20722);
nor U21516 (N_21516,N_20405,N_20418);
nor U21517 (N_21517,N_20667,N_20462);
nand U21518 (N_21518,N_20889,N_20922);
nand U21519 (N_21519,N_20902,N_20481);
or U21520 (N_21520,N_20616,N_20717);
or U21521 (N_21521,N_20936,N_20923);
or U21522 (N_21522,N_20839,N_20447);
nand U21523 (N_21523,N_20442,N_20936);
nor U21524 (N_21524,N_20768,N_20671);
or U21525 (N_21525,N_20890,N_20915);
or U21526 (N_21526,N_20638,N_20518);
nor U21527 (N_21527,N_20657,N_20840);
or U21528 (N_21528,N_20802,N_20767);
nand U21529 (N_21529,N_20761,N_20963);
nor U21530 (N_21530,N_20955,N_20884);
and U21531 (N_21531,N_20516,N_20674);
nand U21532 (N_21532,N_20975,N_20558);
nor U21533 (N_21533,N_20407,N_20932);
and U21534 (N_21534,N_20421,N_20936);
or U21535 (N_21535,N_20823,N_20825);
nor U21536 (N_21536,N_20951,N_20515);
xor U21537 (N_21537,N_20552,N_20611);
nand U21538 (N_21538,N_20416,N_20547);
nor U21539 (N_21539,N_20873,N_20906);
nor U21540 (N_21540,N_20880,N_20727);
or U21541 (N_21541,N_20872,N_20909);
xor U21542 (N_21542,N_20936,N_20614);
nand U21543 (N_21543,N_20725,N_20699);
and U21544 (N_21544,N_20953,N_20630);
or U21545 (N_21545,N_20632,N_20744);
nand U21546 (N_21546,N_20897,N_20850);
and U21547 (N_21547,N_20711,N_20956);
and U21548 (N_21548,N_20900,N_20800);
nand U21549 (N_21549,N_20558,N_20467);
or U21550 (N_21550,N_20722,N_20490);
or U21551 (N_21551,N_20705,N_20827);
or U21552 (N_21552,N_20994,N_20730);
or U21553 (N_21553,N_20945,N_20478);
and U21554 (N_21554,N_20636,N_20460);
nand U21555 (N_21555,N_20883,N_20764);
nor U21556 (N_21556,N_20982,N_20432);
or U21557 (N_21557,N_20712,N_20657);
nand U21558 (N_21558,N_20742,N_20946);
or U21559 (N_21559,N_20777,N_20794);
xor U21560 (N_21560,N_20676,N_20725);
nor U21561 (N_21561,N_20430,N_20480);
nand U21562 (N_21562,N_20448,N_20901);
or U21563 (N_21563,N_20555,N_20480);
or U21564 (N_21564,N_20922,N_20687);
or U21565 (N_21565,N_20499,N_20948);
nand U21566 (N_21566,N_20963,N_20970);
or U21567 (N_21567,N_20492,N_20934);
nand U21568 (N_21568,N_20926,N_20706);
nor U21569 (N_21569,N_20631,N_20674);
and U21570 (N_21570,N_20406,N_20580);
nand U21571 (N_21571,N_20528,N_20773);
nor U21572 (N_21572,N_20694,N_20780);
or U21573 (N_21573,N_20558,N_20626);
and U21574 (N_21574,N_20879,N_20418);
nor U21575 (N_21575,N_20589,N_20758);
or U21576 (N_21576,N_20883,N_20679);
nand U21577 (N_21577,N_20654,N_20831);
nand U21578 (N_21578,N_20849,N_20775);
nand U21579 (N_21579,N_20523,N_20679);
nor U21580 (N_21580,N_20563,N_20725);
or U21581 (N_21581,N_20573,N_20601);
or U21582 (N_21582,N_20487,N_20957);
nand U21583 (N_21583,N_20491,N_20910);
and U21584 (N_21584,N_20441,N_20877);
xnor U21585 (N_21585,N_20402,N_20705);
or U21586 (N_21586,N_20638,N_20845);
xnor U21587 (N_21587,N_20511,N_20717);
xnor U21588 (N_21588,N_20504,N_20780);
nor U21589 (N_21589,N_20908,N_20541);
nor U21590 (N_21590,N_20643,N_20732);
nor U21591 (N_21591,N_20609,N_20709);
and U21592 (N_21592,N_20751,N_20728);
nand U21593 (N_21593,N_20908,N_20509);
nand U21594 (N_21594,N_20957,N_20767);
and U21595 (N_21595,N_20992,N_20884);
or U21596 (N_21596,N_20615,N_20820);
or U21597 (N_21597,N_20672,N_20802);
nor U21598 (N_21598,N_20995,N_20710);
nand U21599 (N_21599,N_20502,N_20727);
or U21600 (N_21600,N_21238,N_21073);
and U21601 (N_21601,N_21273,N_21028);
or U21602 (N_21602,N_21218,N_21467);
or U21603 (N_21603,N_21215,N_21111);
nor U21604 (N_21604,N_21227,N_21569);
xor U21605 (N_21605,N_21145,N_21189);
and U21606 (N_21606,N_21208,N_21517);
xor U21607 (N_21607,N_21287,N_21272);
nand U21608 (N_21608,N_21586,N_21091);
xnor U21609 (N_21609,N_21580,N_21367);
nand U21610 (N_21610,N_21480,N_21550);
and U21611 (N_21611,N_21071,N_21489);
or U21612 (N_21612,N_21088,N_21035);
xnor U21613 (N_21613,N_21519,N_21102);
or U21614 (N_21614,N_21545,N_21572);
and U21615 (N_21615,N_21255,N_21532);
nor U21616 (N_21616,N_21282,N_21042);
or U21617 (N_21617,N_21058,N_21495);
or U21618 (N_21618,N_21149,N_21261);
and U21619 (N_21619,N_21103,N_21194);
nor U21620 (N_21620,N_21222,N_21106);
xnor U21621 (N_21621,N_21464,N_21076);
nand U21622 (N_21622,N_21055,N_21114);
or U21623 (N_21623,N_21119,N_21033);
xor U21624 (N_21624,N_21191,N_21473);
nor U21625 (N_21625,N_21270,N_21478);
and U21626 (N_21626,N_21414,N_21515);
and U21627 (N_21627,N_21306,N_21178);
and U21628 (N_21628,N_21576,N_21059);
and U21629 (N_21629,N_21159,N_21000);
and U21630 (N_21630,N_21300,N_21117);
and U21631 (N_21631,N_21499,N_21556);
nand U21632 (N_21632,N_21253,N_21125);
nand U21633 (N_21633,N_21368,N_21157);
nor U21634 (N_21634,N_21199,N_21390);
xor U21635 (N_21635,N_21265,N_21074);
and U21636 (N_21636,N_21002,N_21320);
nor U21637 (N_21637,N_21493,N_21160);
nor U21638 (N_21638,N_21234,N_21298);
and U21639 (N_21639,N_21455,N_21446);
nor U21640 (N_21640,N_21024,N_21409);
nand U21641 (N_21641,N_21064,N_21213);
and U21642 (N_21642,N_21264,N_21482);
nor U21643 (N_21643,N_21423,N_21010);
xnor U21644 (N_21644,N_21245,N_21528);
nand U21645 (N_21645,N_21297,N_21562);
or U21646 (N_21646,N_21520,N_21483);
nor U21647 (N_21647,N_21439,N_21434);
nor U21648 (N_21648,N_21574,N_21563);
nand U21649 (N_21649,N_21456,N_21212);
and U21650 (N_21650,N_21179,N_21501);
or U21651 (N_21651,N_21382,N_21118);
nor U21652 (N_21652,N_21284,N_21260);
nor U21653 (N_21653,N_21132,N_21012);
and U21654 (N_21654,N_21396,N_21214);
and U21655 (N_21655,N_21588,N_21559);
nor U21656 (N_21656,N_21551,N_21384);
nand U21657 (N_21657,N_21051,N_21529);
nand U21658 (N_21658,N_21344,N_21204);
nor U21659 (N_21659,N_21475,N_21417);
and U21660 (N_21660,N_21343,N_21141);
nand U21661 (N_21661,N_21110,N_21124);
nand U21662 (N_21662,N_21504,N_21155);
nor U21663 (N_21663,N_21121,N_21197);
nand U21664 (N_21664,N_21430,N_21415);
nand U21665 (N_21665,N_21162,N_21100);
nand U21666 (N_21666,N_21196,N_21548);
xor U21667 (N_21667,N_21301,N_21358);
nand U21668 (N_21668,N_21257,N_21275);
nor U21669 (N_21669,N_21011,N_21463);
nand U21670 (N_21670,N_21144,N_21554);
xor U21671 (N_21671,N_21007,N_21205);
or U21672 (N_21672,N_21575,N_21509);
nor U21673 (N_21673,N_21505,N_21249);
and U21674 (N_21674,N_21408,N_21078);
and U21675 (N_21675,N_21046,N_21583);
and U21676 (N_21676,N_21017,N_21349);
nand U21677 (N_21677,N_21377,N_21435);
or U21678 (N_21678,N_21597,N_21416);
nor U21679 (N_21679,N_21246,N_21324);
and U21680 (N_21680,N_21019,N_21190);
and U21681 (N_21681,N_21266,N_21457);
nor U21682 (N_21682,N_21471,N_21412);
or U21683 (N_21683,N_21090,N_21268);
or U21684 (N_21684,N_21128,N_21161);
nor U21685 (N_21685,N_21485,N_21198);
nand U21686 (N_21686,N_21443,N_21444);
nor U21687 (N_21687,N_21406,N_21447);
xnor U21688 (N_21688,N_21437,N_21165);
nand U21689 (N_21689,N_21330,N_21135);
xnor U21690 (N_21690,N_21267,N_21307);
nand U21691 (N_21691,N_21587,N_21543);
nor U21692 (N_21692,N_21129,N_21278);
nor U21693 (N_21693,N_21040,N_21027);
nand U21694 (N_21694,N_21316,N_21022);
and U21695 (N_21695,N_21171,N_21168);
and U21696 (N_21696,N_21549,N_21147);
nand U21697 (N_21697,N_21235,N_21228);
nand U21698 (N_21698,N_21462,N_21403);
nand U21699 (N_21699,N_21351,N_21440);
nand U21700 (N_21700,N_21585,N_21236);
nand U21701 (N_21701,N_21080,N_21321);
and U21702 (N_21702,N_21363,N_21518);
or U21703 (N_21703,N_21522,N_21188);
or U21704 (N_21704,N_21295,N_21389);
and U21705 (N_21705,N_21146,N_21225);
nor U21706 (N_21706,N_21345,N_21036);
or U21707 (N_21707,N_21565,N_21594);
xor U21708 (N_21708,N_21038,N_21421);
nor U21709 (N_21709,N_21507,N_21052);
or U21710 (N_21710,N_21387,N_21131);
xor U21711 (N_21711,N_21281,N_21258);
xor U21712 (N_21712,N_21448,N_21442);
or U21713 (N_21713,N_21026,N_21169);
xor U21714 (N_21714,N_21248,N_21481);
and U21715 (N_21715,N_21573,N_21394);
nor U21716 (N_21716,N_21053,N_21180);
nor U21717 (N_21717,N_21101,N_21288);
nand U21718 (N_21718,N_21104,N_21513);
nand U21719 (N_21719,N_21438,N_21049);
xnor U21720 (N_21720,N_21379,N_21044);
nor U21721 (N_21721,N_21057,N_21337);
nor U21722 (N_21722,N_21458,N_21230);
nor U21723 (N_21723,N_21018,N_21364);
nand U21724 (N_21724,N_21325,N_21450);
and U21725 (N_21725,N_21244,N_21174);
nor U21726 (N_21726,N_21151,N_21233);
nor U21727 (N_21727,N_21431,N_21558);
nand U21728 (N_21728,N_21085,N_21309);
and U21729 (N_21729,N_21291,N_21063);
nand U21730 (N_21730,N_21166,N_21259);
or U21731 (N_21731,N_21185,N_21348);
nor U21732 (N_21732,N_21339,N_21461);
nor U21733 (N_21733,N_21034,N_21087);
nor U21734 (N_21734,N_21383,N_21193);
or U21735 (N_21735,N_21332,N_21491);
or U21736 (N_21736,N_21508,N_21203);
nor U21737 (N_21737,N_21177,N_21219);
nor U21738 (N_21738,N_21240,N_21361);
and U21739 (N_21739,N_21136,N_21561);
nand U21740 (N_21740,N_21003,N_21294);
nor U21741 (N_21741,N_21237,N_21590);
or U21742 (N_21742,N_21187,N_21153);
and U21743 (N_21743,N_21164,N_21474);
and U21744 (N_21744,N_21454,N_21163);
nand U21745 (N_21745,N_21410,N_21452);
or U21746 (N_21746,N_21451,N_21534);
nor U21747 (N_21747,N_21560,N_21109);
nand U21748 (N_21748,N_21362,N_21308);
or U21749 (N_21749,N_21502,N_21015);
nor U21750 (N_21750,N_21072,N_21032);
xnor U21751 (N_21751,N_21356,N_21317);
nor U21752 (N_21752,N_21292,N_21388);
and U21753 (N_21753,N_21154,N_21108);
and U21754 (N_21754,N_21150,N_21223);
nand U21755 (N_21755,N_21593,N_21395);
or U21756 (N_21756,N_21577,N_21582);
or U21757 (N_21757,N_21542,N_21503);
xor U21758 (N_21758,N_21279,N_21182);
and U21759 (N_21759,N_21056,N_21274);
and U21760 (N_21760,N_21599,N_21122);
or U21761 (N_21761,N_21391,N_21436);
xnor U21762 (N_21762,N_21054,N_21354);
nand U21763 (N_21763,N_21449,N_21070);
or U21764 (N_21764,N_21239,N_21526);
nand U21765 (N_21765,N_21202,N_21397);
nor U21766 (N_21766,N_21252,N_21302);
nor U21767 (N_21767,N_21142,N_21570);
and U21768 (N_21768,N_21584,N_21369);
and U21769 (N_21769,N_21422,N_21067);
nor U21770 (N_21770,N_21538,N_21004);
or U21771 (N_21771,N_21350,N_21280);
nor U21772 (N_21772,N_21373,N_21381);
or U21773 (N_21773,N_21095,N_21595);
nor U21774 (N_21774,N_21220,N_21544);
nor U21775 (N_21775,N_21120,N_21041);
nor U21776 (N_21776,N_21009,N_21315);
and U21777 (N_21777,N_21566,N_21031);
and U21778 (N_21778,N_21143,N_21494);
nand U21779 (N_21779,N_21312,N_21285);
nand U21780 (N_21780,N_21472,N_21598);
nand U21781 (N_21781,N_21200,N_21310);
and U21782 (N_21782,N_21083,N_21283);
xor U21783 (N_21783,N_21466,N_21357);
nor U21784 (N_21784,N_21360,N_21243);
or U21785 (N_21785,N_21148,N_21097);
xor U21786 (N_21786,N_21401,N_21293);
xor U21787 (N_21787,N_21271,N_21465);
and U21788 (N_21788,N_21335,N_21427);
nand U21789 (N_21789,N_21242,N_21066);
nand U21790 (N_21790,N_21426,N_21299);
and U21791 (N_21791,N_21130,N_21123);
nand U21792 (N_21792,N_21186,N_21127);
and U21793 (N_21793,N_21393,N_21173);
nand U21794 (N_21794,N_21411,N_21082);
and U21795 (N_21795,N_21428,N_21210);
or U21796 (N_21796,N_21392,N_21578);
or U21797 (N_21797,N_21016,N_21328);
nor U21798 (N_21798,N_21013,N_21536);
nor U21799 (N_21799,N_21581,N_21404);
and U21800 (N_21800,N_21183,N_21366);
nor U21801 (N_21801,N_21487,N_21371);
xor U21802 (N_21802,N_21175,N_21579);
nor U21803 (N_21803,N_21081,N_21029);
nand U21804 (N_21804,N_21341,N_21025);
and U21805 (N_21805,N_21476,N_21453);
or U21806 (N_21806,N_21492,N_21069);
nor U21807 (N_21807,N_21079,N_21318);
nor U21808 (N_21808,N_21303,N_21030);
nand U21809 (N_21809,N_21568,N_21506);
nor U21810 (N_21810,N_21094,N_21195);
and U21811 (N_21811,N_21206,N_21247);
and U21812 (N_21812,N_21425,N_21486);
and U21813 (N_21813,N_21353,N_21112);
or U21814 (N_21814,N_21596,N_21068);
xnor U21815 (N_21815,N_21048,N_21232);
nor U21816 (N_21816,N_21207,N_21510);
xnor U21817 (N_21817,N_21342,N_21217);
nand U21818 (N_21818,N_21322,N_21469);
and U21819 (N_21819,N_21241,N_21224);
nor U21820 (N_21820,N_21209,N_21262);
xnor U21821 (N_21821,N_21296,N_21553);
and U21822 (N_21822,N_21540,N_21184);
and U21823 (N_21823,N_21511,N_21201);
and U21824 (N_21824,N_21311,N_21512);
nor U21825 (N_21825,N_21370,N_21398);
nand U21826 (N_21826,N_21564,N_21347);
nor U21827 (N_21827,N_21375,N_21552);
nor U21828 (N_21828,N_21290,N_21571);
xnor U21829 (N_21829,N_21152,N_21005);
and U21830 (N_21830,N_21400,N_21352);
and U21831 (N_21831,N_21385,N_21374);
nor U21832 (N_21832,N_21591,N_21359);
nor U21833 (N_21833,N_21014,N_21331);
xnor U21834 (N_21834,N_21158,N_21329);
nor U21835 (N_21835,N_21589,N_21250);
nor U21836 (N_21836,N_21105,N_21432);
nor U21837 (N_21837,N_21460,N_21170);
and U21838 (N_21838,N_21211,N_21413);
nand U21839 (N_21839,N_21138,N_21497);
or U21840 (N_21840,N_21045,N_21433);
nand U21841 (N_21841,N_21075,N_21365);
and U21842 (N_21842,N_21405,N_21525);
nand U21843 (N_21843,N_21524,N_21407);
or U21844 (N_21844,N_21541,N_21372);
and U21845 (N_21845,N_21077,N_21336);
or U21846 (N_21846,N_21399,N_21484);
xor U21847 (N_21847,N_21289,N_21139);
nor U21848 (N_21848,N_21319,N_21346);
nand U21849 (N_21849,N_21116,N_21023);
xnor U21850 (N_21850,N_21172,N_21424);
nand U21851 (N_21851,N_21084,N_21133);
xnor U21852 (N_21852,N_21313,N_21380);
nor U21853 (N_21853,N_21065,N_21496);
nor U21854 (N_21854,N_21269,N_21555);
or U21855 (N_21855,N_21402,N_21192);
and U21856 (N_21856,N_21176,N_21470);
xor U21857 (N_21857,N_21021,N_21429);
nand U21858 (N_21858,N_21326,N_21156);
nor U21859 (N_21859,N_21305,N_21323);
xor U21860 (N_21860,N_21468,N_21477);
nand U21861 (N_21861,N_21304,N_21231);
xnor U21862 (N_21862,N_21099,N_21251);
nand U21863 (N_21863,N_21086,N_21592);
nand U21864 (N_21864,N_21539,N_21254);
or U21865 (N_21865,N_21226,N_21498);
and U21866 (N_21866,N_21386,N_21340);
and U21867 (N_21867,N_21546,N_21126);
nor U21868 (N_21868,N_21167,N_21216);
nand U21869 (N_21869,N_21256,N_21376);
or U21870 (N_21870,N_21459,N_21089);
xor U21871 (N_21871,N_21327,N_21527);
xor U21872 (N_21872,N_21530,N_21479);
nand U21873 (N_21873,N_21418,N_21557);
and U21874 (N_21874,N_21338,N_21221);
nor U21875 (N_21875,N_21445,N_21181);
nand U21876 (N_21876,N_21137,N_21276);
nor U21877 (N_21877,N_21277,N_21140);
xor U21878 (N_21878,N_21521,N_21062);
and U21879 (N_21879,N_21008,N_21060);
nor U21880 (N_21880,N_21107,N_21050);
nor U21881 (N_21881,N_21039,N_21488);
nand U21882 (N_21882,N_21334,N_21263);
and U21883 (N_21883,N_21514,N_21537);
xnor U21884 (N_21884,N_21113,N_21333);
nor U21885 (N_21885,N_21531,N_21134);
xor U21886 (N_21886,N_21043,N_21096);
nand U21887 (N_21887,N_21490,N_21378);
and U21888 (N_21888,N_21355,N_21535);
or U21889 (N_21889,N_21115,N_21229);
xnor U21890 (N_21890,N_21314,N_21037);
nand U21891 (N_21891,N_21441,N_21567);
or U21892 (N_21892,N_21061,N_21523);
nor U21893 (N_21893,N_21006,N_21092);
nand U21894 (N_21894,N_21286,N_21020);
or U21895 (N_21895,N_21047,N_21419);
and U21896 (N_21896,N_21547,N_21533);
nand U21897 (N_21897,N_21001,N_21516);
xor U21898 (N_21898,N_21098,N_21093);
and U21899 (N_21899,N_21420,N_21500);
xnor U21900 (N_21900,N_21387,N_21327);
nor U21901 (N_21901,N_21484,N_21590);
xnor U21902 (N_21902,N_21466,N_21526);
or U21903 (N_21903,N_21571,N_21339);
nor U21904 (N_21904,N_21423,N_21307);
nand U21905 (N_21905,N_21505,N_21467);
xor U21906 (N_21906,N_21572,N_21316);
nor U21907 (N_21907,N_21410,N_21253);
or U21908 (N_21908,N_21469,N_21499);
nand U21909 (N_21909,N_21553,N_21281);
nor U21910 (N_21910,N_21055,N_21407);
nand U21911 (N_21911,N_21482,N_21119);
nor U21912 (N_21912,N_21105,N_21330);
and U21913 (N_21913,N_21235,N_21365);
nor U21914 (N_21914,N_21373,N_21253);
nand U21915 (N_21915,N_21172,N_21221);
and U21916 (N_21916,N_21053,N_21283);
nor U21917 (N_21917,N_21394,N_21510);
nand U21918 (N_21918,N_21254,N_21337);
and U21919 (N_21919,N_21499,N_21189);
or U21920 (N_21920,N_21249,N_21022);
nand U21921 (N_21921,N_21503,N_21591);
nand U21922 (N_21922,N_21338,N_21403);
nor U21923 (N_21923,N_21233,N_21364);
and U21924 (N_21924,N_21555,N_21436);
or U21925 (N_21925,N_21345,N_21308);
xnor U21926 (N_21926,N_21405,N_21158);
nor U21927 (N_21927,N_21322,N_21174);
and U21928 (N_21928,N_21219,N_21367);
nand U21929 (N_21929,N_21467,N_21283);
or U21930 (N_21930,N_21243,N_21348);
or U21931 (N_21931,N_21554,N_21222);
and U21932 (N_21932,N_21349,N_21193);
and U21933 (N_21933,N_21144,N_21497);
nor U21934 (N_21934,N_21193,N_21471);
nand U21935 (N_21935,N_21270,N_21346);
or U21936 (N_21936,N_21273,N_21190);
nor U21937 (N_21937,N_21564,N_21312);
nand U21938 (N_21938,N_21331,N_21209);
or U21939 (N_21939,N_21224,N_21478);
and U21940 (N_21940,N_21516,N_21391);
nand U21941 (N_21941,N_21433,N_21283);
nand U21942 (N_21942,N_21504,N_21206);
nand U21943 (N_21943,N_21011,N_21014);
and U21944 (N_21944,N_21040,N_21542);
or U21945 (N_21945,N_21346,N_21476);
and U21946 (N_21946,N_21306,N_21436);
or U21947 (N_21947,N_21192,N_21155);
nand U21948 (N_21948,N_21013,N_21522);
or U21949 (N_21949,N_21566,N_21067);
xnor U21950 (N_21950,N_21315,N_21019);
nor U21951 (N_21951,N_21546,N_21421);
nor U21952 (N_21952,N_21425,N_21278);
nand U21953 (N_21953,N_21358,N_21455);
or U21954 (N_21954,N_21134,N_21483);
or U21955 (N_21955,N_21426,N_21275);
or U21956 (N_21956,N_21378,N_21554);
and U21957 (N_21957,N_21407,N_21099);
and U21958 (N_21958,N_21556,N_21408);
nand U21959 (N_21959,N_21538,N_21531);
nor U21960 (N_21960,N_21161,N_21028);
or U21961 (N_21961,N_21479,N_21580);
xnor U21962 (N_21962,N_21511,N_21579);
nor U21963 (N_21963,N_21573,N_21332);
xor U21964 (N_21964,N_21219,N_21304);
nor U21965 (N_21965,N_21381,N_21455);
and U21966 (N_21966,N_21121,N_21015);
nor U21967 (N_21967,N_21381,N_21122);
and U21968 (N_21968,N_21178,N_21024);
or U21969 (N_21969,N_21546,N_21535);
nor U21970 (N_21970,N_21538,N_21595);
nor U21971 (N_21971,N_21314,N_21299);
and U21972 (N_21972,N_21504,N_21161);
nor U21973 (N_21973,N_21425,N_21344);
nand U21974 (N_21974,N_21485,N_21336);
nand U21975 (N_21975,N_21462,N_21334);
and U21976 (N_21976,N_21228,N_21538);
nor U21977 (N_21977,N_21311,N_21464);
nand U21978 (N_21978,N_21029,N_21531);
nand U21979 (N_21979,N_21195,N_21287);
or U21980 (N_21980,N_21192,N_21503);
and U21981 (N_21981,N_21108,N_21169);
or U21982 (N_21982,N_21310,N_21296);
or U21983 (N_21983,N_21053,N_21287);
nor U21984 (N_21984,N_21033,N_21086);
nand U21985 (N_21985,N_21089,N_21521);
nor U21986 (N_21986,N_21344,N_21315);
or U21987 (N_21987,N_21429,N_21302);
nor U21988 (N_21988,N_21495,N_21133);
nor U21989 (N_21989,N_21572,N_21196);
nand U21990 (N_21990,N_21354,N_21262);
or U21991 (N_21991,N_21438,N_21566);
and U21992 (N_21992,N_21506,N_21447);
and U21993 (N_21993,N_21370,N_21331);
nor U21994 (N_21994,N_21242,N_21320);
and U21995 (N_21995,N_21084,N_21599);
nor U21996 (N_21996,N_21003,N_21184);
or U21997 (N_21997,N_21582,N_21422);
or U21998 (N_21998,N_21390,N_21319);
nand U21999 (N_21999,N_21466,N_21145);
and U22000 (N_22000,N_21459,N_21440);
and U22001 (N_22001,N_21376,N_21255);
or U22002 (N_22002,N_21139,N_21278);
and U22003 (N_22003,N_21364,N_21087);
nor U22004 (N_22004,N_21097,N_21573);
xor U22005 (N_22005,N_21329,N_21050);
or U22006 (N_22006,N_21237,N_21319);
xnor U22007 (N_22007,N_21408,N_21134);
and U22008 (N_22008,N_21343,N_21443);
nand U22009 (N_22009,N_21323,N_21219);
nand U22010 (N_22010,N_21418,N_21124);
nand U22011 (N_22011,N_21241,N_21196);
nor U22012 (N_22012,N_21527,N_21431);
or U22013 (N_22013,N_21098,N_21043);
nand U22014 (N_22014,N_21599,N_21371);
nor U22015 (N_22015,N_21317,N_21340);
nand U22016 (N_22016,N_21439,N_21383);
or U22017 (N_22017,N_21467,N_21148);
xnor U22018 (N_22018,N_21043,N_21440);
and U22019 (N_22019,N_21518,N_21230);
nand U22020 (N_22020,N_21131,N_21162);
nor U22021 (N_22021,N_21332,N_21237);
nor U22022 (N_22022,N_21031,N_21329);
or U22023 (N_22023,N_21454,N_21154);
xor U22024 (N_22024,N_21122,N_21034);
or U22025 (N_22025,N_21595,N_21121);
xor U22026 (N_22026,N_21230,N_21140);
or U22027 (N_22027,N_21570,N_21590);
nand U22028 (N_22028,N_21103,N_21164);
or U22029 (N_22029,N_21279,N_21547);
or U22030 (N_22030,N_21276,N_21098);
nor U22031 (N_22031,N_21195,N_21160);
nor U22032 (N_22032,N_21204,N_21254);
and U22033 (N_22033,N_21378,N_21169);
and U22034 (N_22034,N_21389,N_21589);
xor U22035 (N_22035,N_21372,N_21444);
nand U22036 (N_22036,N_21293,N_21426);
and U22037 (N_22037,N_21509,N_21558);
or U22038 (N_22038,N_21181,N_21044);
or U22039 (N_22039,N_21257,N_21152);
or U22040 (N_22040,N_21440,N_21192);
nand U22041 (N_22041,N_21147,N_21300);
and U22042 (N_22042,N_21410,N_21542);
or U22043 (N_22043,N_21170,N_21461);
or U22044 (N_22044,N_21171,N_21231);
nor U22045 (N_22045,N_21037,N_21578);
nor U22046 (N_22046,N_21304,N_21117);
and U22047 (N_22047,N_21227,N_21390);
nand U22048 (N_22048,N_21152,N_21030);
and U22049 (N_22049,N_21320,N_21245);
nor U22050 (N_22050,N_21422,N_21307);
nor U22051 (N_22051,N_21108,N_21460);
and U22052 (N_22052,N_21090,N_21050);
and U22053 (N_22053,N_21260,N_21508);
xor U22054 (N_22054,N_21554,N_21118);
and U22055 (N_22055,N_21545,N_21578);
or U22056 (N_22056,N_21347,N_21276);
and U22057 (N_22057,N_21583,N_21125);
or U22058 (N_22058,N_21021,N_21092);
xnor U22059 (N_22059,N_21422,N_21384);
or U22060 (N_22060,N_21308,N_21105);
or U22061 (N_22061,N_21263,N_21446);
nand U22062 (N_22062,N_21234,N_21207);
and U22063 (N_22063,N_21466,N_21568);
and U22064 (N_22064,N_21226,N_21070);
nand U22065 (N_22065,N_21593,N_21516);
or U22066 (N_22066,N_21371,N_21506);
or U22067 (N_22067,N_21546,N_21118);
xor U22068 (N_22068,N_21208,N_21224);
and U22069 (N_22069,N_21109,N_21384);
nand U22070 (N_22070,N_21327,N_21418);
nor U22071 (N_22071,N_21376,N_21330);
nand U22072 (N_22072,N_21187,N_21004);
nand U22073 (N_22073,N_21494,N_21155);
nand U22074 (N_22074,N_21526,N_21213);
nor U22075 (N_22075,N_21107,N_21116);
and U22076 (N_22076,N_21565,N_21488);
nand U22077 (N_22077,N_21418,N_21363);
xnor U22078 (N_22078,N_21032,N_21137);
and U22079 (N_22079,N_21260,N_21446);
or U22080 (N_22080,N_21473,N_21556);
or U22081 (N_22081,N_21326,N_21433);
or U22082 (N_22082,N_21158,N_21270);
and U22083 (N_22083,N_21132,N_21573);
and U22084 (N_22084,N_21029,N_21328);
nor U22085 (N_22085,N_21138,N_21139);
nand U22086 (N_22086,N_21439,N_21529);
nor U22087 (N_22087,N_21108,N_21144);
nor U22088 (N_22088,N_21162,N_21210);
xnor U22089 (N_22089,N_21238,N_21583);
nand U22090 (N_22090,N_21481,N_21552);
nand U22091 (N_22091,N_21073,N_21476);
and U22092 (N_22092,N_21140,N_21468);
and U22093 (N_22093,N_21445,N_21106);
nor U22094 (N_22094,N_21191,N_21139);
nor U22095 (N_22095,N_21417,N_21195);
or U22096 (N_22096,N_21565,N_21077);
and U22097 (N_22097,N_21409,N_21230);
and U22098 (N_22098,N_21351,N_21129);
nand U22099 (N_22099,N_21408,N_21462);
nand U22100 (N_22100,N_21394,N_21040);
and U22101 (N_22101,N_21090,N_21260);
nand U22102 (N_22102,N_21100,N_21283);
and U22103 (N_22103,N_21563,N_21511);
nor U22104 (N_22104,N_21433,N_21160);
or U22105 (N_22105,N_21465,N_21406);
or U22106 (N_22106,N_21235,N_21578);
or U22107 (N_22107,N_21329,N_21431);
nand U22108 (N_22108,N_21104,N_21403);
and U22109 (N_22109,N_21003,N_21367);
or U22110 (N_22110,N_21491,N_21584);
or U22111 (N_22111,N_21047,N_21229);
nand U22112 (N_22112,N_21268,N_21538);
and U22113 (N_22113,N_21077,N_21316);
nor U22114 (N_22114,N_21248,N_21172);
or U22115 (N_22115,N_21025,N_21583);
nor U22116 (N_22116,N_21045,N_21115);
nor U22117 (N_22117,N_21155,N_21459);
nor U22118 (N_22118,N_21356,N_21125);
xor U22119 (N_22119,N_21559,N_21594);
or U22120 (N_22120,N_21143,N_21570);
nor U22121 (N_22121,N_21371,N_21548);
nor U22122 (N_22122,N_21461,N_21358);
and U22123 (N_22123,N_21027,N_21293);
and U22124 (N_22124,N_21589,N_21269);
nand U22125 (N_22125,N_21555,N_21363);
nand U22126 (N_22126,N_21237,N_21003);
or U22127 (N_22127,N_21321,N_21241);
and U22128 (N_22128,N_21090,N_21466);
nor U22129 (N_22129,N_21543,N_21492);
or U22130 (N_22130,N_21236,N_21071);
or U22131 (N_22131,N_21264,N_21250);
nand U22132 (N_22132,N_21429,N_21199);
and U22133 (N_22133,N_21068,N_21357);
nor U22134 (N_22134,N_21287,N_21028);
and U22135 (N_22135,N_21024,N_21597);
and U22136 (N_22136,N_21226,N_21062);
or U22137 (N_22137,N_21403,N_21384);
xnor U22138 (N_22138,N_21454,N_21160);
nor U22139 (N_22139,N_21169,N_21183);
or U22140 (N_22140,N_21142,N_21322);
and U22141 (N_22141,N_21352,N_21226);
nand U22142 (N_22142,N_21328,N_21035);
or U22143 (N_22143,N_21147,N_21545);
nor U22144 (N_22144,N_21532,N_21478);
and U22145 (N_22145,N_21583,N_21457);
nor U22146 (N_22146,N_21126,N_21457);
xor U22147 (N_22147,N_21240,N_21151);
or U22148 (N_22148,N_21440,N_21421);
nand U22149 (N_22149,N_21031,N_21168);
xnor U22150 (N_22150,N_21437,N_21050);
xor U22151 (N_22151,N_21291,N_21065);
nand U22152 (N_22152,N_21370,N_21383);
nor U22153 (N_22153,N_21209,N_21484);
and U22154 (N_22154,N_21373,N_21060);
and U22155 (N_22155,N_21218,N_21011);
xor U22156 (N_22156,N_21058,N_21193);
xor U22157 (N_22157,N_21049,N_21075);
nor U22158 (N_22158,N_21373,N_21384);
and U22159 (N_22159,N_21585,N_21591);
or U22160 (N_22160,N_21020,N_21009);
and U22161 (N_22161,N_21398,N_21291);
nand U22162 (N_22162,N_21089,N_21479);
nor U22163 (N_22163,N_21047,N_21458);
and U22164 (N_22164,N_21356,N_21054);
nand U22165 (N_22165,N_21397,N_21369);
nor U22166 (N_22166,N_21277,N_21434);
xor U22167 (N_22167,N_21542,N_21473);
or U22168 (N_22168,N_21399,N_21596);
or U22169 (N_22169,N_21338,N_21048);
or U22170 (N_22170,N_21463,N_21515);
and U22171 (N_22171,N_21054,N_21431);
nor U22172 (N_22172,N_21134,N_21331);
nor U22173 (N_22173,N_21334,N_21505);
nor U22174 (N_22174,N_21444,N_21594);
and U22175 (N_22175,N_21583,N_21075);
nor U22176 (N_22176,N_21523,N_21511);
and U22177 (N_22177,N_21499,N_21301);
nand U22178 (N_22178,N_21408,N_21125);
nor U22179 (N_22179,N_21498,N_21249);
and U22180 (N_22180,N_21486,N_21278);
xor U22181 (N_22181,N_21054,N_21043);
and U22182 (N_22182,N_21370,N_21435);
nand U22183 (N_22183,N_21248,N_21020);
nand U22184 (N_22184,N_21060,N_21124);
nor U22185 (N_22185,N_21322,N_21537);
nand U22186 (N_22186,N_21541,N_21297);
and U22187 (N_22187,N_21368,N_21500);
and U22188 (N_22188,N_21065,N_21321);
or U22189 (N_22189,N_21149,N_21405);
nor U22190 (N_22190,N_21563,N_21541);
nor U22191 (N_22191,N_21511,N_21595);
nor U22192 (N_22192,N_21143,N_21417);
or U22193 (N_22193,N_21038,N_21451);
and U22194 (N_22194,N_21521,N_21106);
nor U22195 (N_22195,N_21491,N_21153);
nand U22196 (N_22196,N_21397,N_21428);
and U22197 (N_22197,N_21016,N_21535);
nor U22198 (N_22198,N_21439,N_21262);
or U22199 (N_22199,N_21493,N_21282);
or U22200 (N_22200,N_22030,N_21908);
or U22201 (N_22201,N_21697,N_22069);
nor U22202 (N_22202,N_21974,N_22133);
and U22203 (N_22203,N_21986,N_21676);
nor U22204 (N_22204,N_21721,N_21724);
or U22205 (N_22205,N_22059,N_21686);
or U22206 (N_22206,N_21819,N_21913);
and U22207 (N_22207,N_21649,N_22074);
nor U22208 (N_22208,N_22114,N_22000);
and U22209 (N_22209,N_22019,N_21678);
or U22210 (N_22210,N_21743,N_21995);
and U22211 (N_22211,N_21934,N_21831);
nor U22212 (N_22212,N_21618,N_21951);
xnor U22213 (N_22213,N_21834,N_21758);
nand U22214 (N_22214,N_21882,N_22130);
nand U22215 (N_22215,N_22186,N_21639);
nor U22216 (N_22216,N_21863,N_21768);
nor U22217 (N_22217,N_21693,N_21806);
xor U22218 (N_22218,N_21792,N_21738);
or U22219 (N_22219,N_22189,N_22141);
nor U22220 (N_22220,N_21750,N_22092);
nor U22221 (N_22221,N_21628,N_21999);
or U22222 (N_22222,N_22024,N_22159);
nand U22223 (N_22223,N_21720,N_22048);
xnor U22224 (N_22224,N_21810,N_22004);
nand U22225 (N_22225,N_21947,N_21993);
and U22226 (N_22226,N_22055,N_21958);
nor U22227 (N_22227,N_21983,N_22009);
nor U22228 (N_22228,N_21621,N_21856);
or U22229 (N_22229,N_21719,N_22149);
nor U22230 (N_22230,N_21898,N_21836);
or U22231 (N_22231,N_22148,N_21645);
or U22232 (N_22232,N_21790,N_21729);
nand U22233 (N_22233,N_21840,N_21795);
nor U22234 (N_22234,N_21804,N_21896);
nor U22235 (N_22235,N_21927,N_22120);
nand U22236 (N_22236,N_21933,N_22010);
xor U22237 (N_22237,N_21734,N_21873);
and U22238 (N_22238,N_21937,N_21679);
nor U22239 (N_22239,N_22080,N_22053);
nor U22240 (N_22240,N_21919,N_21793);
nand U22241 (N_22241,N_21845,N_21814);
nand U22242 (N_22242,N_21888,N_21765);
nor U22243 (N_22243,N_22140,N_21626);
nor U22244 (N_22244,N_21813,N_22040);
xor U22245 (N_22245,N_21877,N_21635);
nor U22246 (N_22246,N_21981,N_22005);
xnor U22247 (N_22247,N_21783,N_21699);
nand U22248 (N_22248,N_21610,N_21891);
nand U22249 (N_22249,N_21970,N_21668);
or U22250 (N_22250,N_22191,N_21672);
nand U22251 (N_22251,N_21713,N_21736);
nor U22252 (N_22252,N_21885,N_21656);
and U22253 (N_22253,N_21786,N_21922);
and U22254 (N_22254,N_21715,N_21828);
and U22255 (N_22255,N_22104,N_21780);
or U22256 (N_22256,N_21952,N_22015);
xor U22257 (N_22257,N_22129,N_22071);
nand U22258 (N_22258,N_21769,N_21853);
or U22259 (N_22259,N_21906,N_21777);
or U22260 (N_22260,N_21946,N_21627);
and U22261 (N_22261,N_22115,N_21704);
or U22262 (N_22262,N_21924,N_21812);
and U22263 (N_22263,N_21601,N_22042);
nand U22264 (N_22264,N_22135,N_21954);
nor U22265 (N_22265,N_21962,N_21920);
nor U22266 (N_22266,N_21789,N_22100);
xor U22267 (N_22267,N_21778,N_21918);
nand U22268 (N_22268,N_22028,N_21982);
and U22269 (N_22269,N_21605,N_21817);
or U22270 (N_22270,N_21915,N_21741);
xnor U22271 (N_22271,N_21646,N_21772);
and U22272 (N_22272,N_21904,N_21648);
nand U22273 (N_22273,N_21994,N_22188);
xor U22274 (N_22274,N_21722,N_21859);
and U22275 (N_22275,N_21881,N_21643);
or U22276 (N_22276,N_21655,N_21797);
or U22277 (N_22277,N_22112,N_22187);
nor U22278 (N_22278,N_21886,N_21826);
nand U22279 (N_22279,N_22142,N_21718);
nor U22280 (N_22280,N_21811,N_21953);
xor U22281 (N_22281,N_21996,N_22056);
and U22282 (N_22282,N_22164,N_21868);
nand U22283 (N_22283,N_21726,N_21916);
nor U22284 (N_22284,N_22105,N_22096);
or U22285 (N_22285,N_21884,N_21689);
xnor U22286 (N_22286,N_21696,N_21972);
and U22287 (N_22287,N_21692,N_21880);
nand U22288 (N_22288,N_22116,N_21802);
nand U22289 (N_22289,N_21740,N_21932);
xor U22290 (N_22290,N_22183,N_21712);
nor U22291 (N_22291,N_22083,N_22051);
xor U22292 (N_22292,N_21682,N_22097);
nand U22293 (N_22293,N_22160,N_22124);
and U22294 (N_22294,N_21754,N_21869);
and U22295 (N_22295,N_21889,N_22122);
nor U22296 (N_22296,N_21905,N_21979);
nand U22297 (N_22297,N_22166,N_21787);
or U22298 (N_22298,N_21847,N_21878);
nand U22299 (N_22299,N_21807,N_22151);
and U22300 (N_22300,N_21690,N_21710);
nand U22301 (N_22301,N_21717,N_21631);
nor U22302 (N_22302,N_21921,N_22084);
nand U22303 (N_22303,N_22144,N_21669);
and U22304 (N_22304,N_22006,N_21989);
and U22305 (N_22305,N_22063,N_22134);
and U22306 (N_22306,N_21911,N_22181);
or U22307 (N_22307,N_22075,N_21650);
and U22308 (N_22308,N_21624,N_21688);
and U22309 (N_22309,N_21727,N_21959);
xor U22310 (N_22310,N_22155,N_21956);
nand U22311 (N_22311,N_22008,N_21684);
and U22312 (N_22312,N_21865,N_21773);
xor U22313 (N_22313,N_22038,N_22003);
xnor U22314 (N_22314,N_22065,N_22177);
nand U22315 (N_22315,N_22190,N_21653);
and U22316 (N_22316,N_21964,N_22067);
nor U22317 (N_22317,N_21666,N_22027);
nand U22318 (N_22318,N_21914,N_21879);
and U22319 (N_22319,N_22108,N_22046);
nand U22320 (N_22320,N_21867,N_21785);
nand U22321 (N_22321,N_21667,N_21900);
nor U22322 (N_22322,N_21917,N_22193);
or U22323 (N_22323,N_21971,N_21941);
nor U22324 (N_22324,N_22026,N_21788);
nor U22325 (N_22325,N_21706,N_21809);
nand U22326 (N_22326,N_22079,N_22111);
nor U22327 (N_22327,N_21665,N_22125);
or U22328 (N_22328,N_21730,N_21830);
nor U22329 (N_22329,N_22171,N_21857);
nand U22330 (N_22330,N_21829,N_22131);
or U22331 (N_22331,N_21822,N_22179);
and U22332 (N_22332,N_21942,N_21897);
nand U22333 (N_22333,N_22158,N_21851);
xor U22334 (N_22334,N_21808,N_22087);
and U22335 (N_22335,N_22176,N_21861);
nand U22336 (N_22336,N_21600,N_22168);
or U22337 (N_22337,N_21864,N_22045);
and U22338 (N_22338,N_21770,N_22066);
or U22339 (N_22339,N_21659,N_22049);
nor U22340 (N_22340,N_22013,N_21936);
or U22341 (N_22341,N_21733,N_21620);
and U22342 (N_22342,N_21703,N_22002);
or U22343 (N_22343,N_22021,N_21849);
nor U22344 (N_22344,N_21671,N_22077);
nand U22345 (N_22345,N_21776,N_21931);
and U22346 (N_22346,N_21670,N_21943);
and U22347 (N_22347,N_21640,N_21606);
nor U22348 (N_22348,N_22172,N_22139);
nand U22349 (N_22349,N_21850,N_21700);
nand U22350 (N_22350,N_22039,N_21641);
nand U22351 (N_22351,N_22043,N_22011);
xor U22352 (N_22352,N_21798,N_21766);
nand U22353 (N_22353,N_21816,N_22025);
or U22354 (N_22354,N_22060,N_22192);
nand U22355 (N_22355,N_22072,N_22194);
xnor U22356 (N_22356,N_21732,N_21815);
nor U22357 (N_22357,N_21841,N_21955);
nor U22358 (N_22358,N_21756,N_21779);
and U22359 (N_22359,N_21698,N_22161);
nand U22360 (N_22360,N_22090,N_21607);
xnor U22361 (N_22361,N_22001,N_22031);
and U22362 (N_22362,N_22052,N_22153);
xnor U22363 (N_22363,N_21753,N_21866);
nand U22364 (N_22364,N_21794,N_22016);
nand U22365 (N_22365,N_21782,N_21848);
nor U22366 (N_22366,N_21895,N_22170);
or U22367 (N_22367,N_21912,N_21883);
or U22368 (N_22368,N_22036,N_22126);
nor U22369 (N_22369,N_22068,N_21761);
or U22370 (N_22370,N_21680,N_22118);
xor U22371 (N_22371,N_21751,N_21839);
nor U22372 (N_22372,N_21949,N_21760);
and U22373 (N_22373,N_21661,N_22091);
and U22374 (N_22374,N_21651,N_21695);
and U22375 (N_22375,N_21854,N_21691);
or U22376 (N_22376,N_21616,N_21612);
nor U22377 (N_22377,N_22101,N_22098);
nand U22378 (N_22378,N_21745,N_22123);
and U22379 (N_22379,N_22197,N_22064);
and U22380 (N_22380,N_21764,N_22081);
nor U22381 (N_22381,N_22119,N_21614);
and U22382 (N_22382,N_22157,N_22089);
nor U22383 (N_22383,N_22106,N_21892);
nand U22384 (N_22384,N_21967,N_21910);
nand U22385 (N_22385,N_21664,N_21843);
or U22386 (N_22386,N_21928,N_21742);
nand U22387 (N_22387,N_21821,N_21630);
and U22388 (N_22388,N_21976,N_21615);
and U22389 (N_22389,N_21781,N_21683);
and U22390 (N_22390,N_21835,N_21739);
or U22391 (N_22391,N_21784,N_22137);
and U22392 (N_22392,N_22033,N_22154);
and U22393 (N_22393,N_21998,N_22162);
nor U22394 (N_22394,N_21948,N_21842);
or U22395 (N_22395,N_22014,N_21632);
xnor U22396 (N_22396,N_22032,N_22095);
xor U22397 (N_22397,N_21702,N_21987);
nand U22398 (N_22398,N_21992,N_21746);
and U22399 (N_22399,N_22184,N_21709);
nand U22400 (N_22400,N_21929,N_22070);
nand U22401 (N_22401,N_22062,N_21663);
nand U22402 (N_22402,N_22165,N_22061);
nand U22403 (N_22403,N_22195,N_21611);
xnor U22404 (N_22404,N_21613,N_21716);
nand U22405 (N_22405,N_21930,N_21938);
nor U22406 (N_22406,N_22086,N_21731);
nand U22407 (N_22407,N_22037,N_22110);
and U22408 (N_22408,N_21893,N_21796);
and U22409 (N_22409,N_22174,N_21852);
and U22410 (N_22410,N_22107,N_21625);
nand U22411 (N_22411,N_22128,N_21755);
or U22412 (N_22412,N_21735,N_22182);
and U22413 (N_22413,N_22073,N_21875);
or U22414 (N_22414,N_21708,N_22023);
or U22415 (N_22415,N_22088,N_21660);
or U22416 (N_22416,N_22198,N_21838);
or U22417 (N_22417,N_21874,N_21681);
xor U22418 (N_22418,N_21894,N_22121);
nor U22419 (N_22419,N_22143,N_21837);
and U22420 (N_22420,N_22169,N_22029);
nor U22421 (N_22421,N_21961,N_21673);
and U22422 (N_22422,N_22173,N_21991);
or U22423 (N_22423,N_21677,N_21890);
nor U22424 (N_22424,N_22099,N_21871);
nand U22425 (N_22425,N_22034,N_21767);
nor U22426 (N_22426,N_21633,N_22175);
and U22427 (N_22427,N_21820,N_21622);
or U22428 (N_22428,N_21824,N_21602);
and U22429 (N_22429,N_22094,N_21675);
nand U22430 (N_22430,N_21623,N_21763);
nor U22431 (N_22431,N_21714,N_22007);
and U22432 (N_22432,N_22103,N_21725);
nand U22433 (N_22433,N_21926,N_21757);
and U22434 (N_22434,N_22057,N_21858);
nand U22435 (N_22435,N_22117,N_22138);
or U22436 (N_22436,N_21771,N_21711);
nor U22437 (N_22437,N_21907,N_22196);
nor U22438 (N_22438,N_21748,N_21872);
nor U22439 (N_22439,N_22163,N_21844);
and U22440 (N_22440,N_22132,N_21899);
or U22441 (N_22441,N_21965,N_21980);
nand U22442 (N_22442,N_21985,N_21801);
or U22443 (N_22443,N_21657,N_21800);
nor U22444 (N_22444,N_21966,N_22058);
and U22445 (N_22445,N_21634,N_22136);
xnor U22446 (N_22446,N_21990,N_21774);
nor U22447 (N_22447,N_21876,N_21723);
nand U22448 (N_22448,N_21957,N_21644);
or U22449 (N_22449,N_21997,N_21638);
and U22450 (N_22450,N_21799,N_22044);
nor U22451 (N_22451,N_21827,N_22109);
or U22452 (N_22452,N_21687,N_21860);
nand U22453 (N_22453,N_21870,N_21940);
nand U22454 (N_22454,N_21609,N_21744);
and U22455 (N_22455,N_22041,N_22035);
nor U22456 (N_22456,N_22180,N_21969);
nand U22457 (N_22457,N_21832,N_21749);
xnor U22458 (N_22458,N_21747,N_21846);
and U22459 (N_22459,N_22150,N_21674);
and U22460 (N_22460,N_21707,N_21775);
nand U22461 (N_22461,N_21909,N_21728);
nand U22462 (N_22462,N_21608,N_21662);
or U22463 (N_22463,N_21603,N_21803);
xor U22464 (N_22464,N_22082,N_21737);
nand U22465 (N_22465,N_21752,N_21945);
nand U22466 (N_22466,N_22047,N_22102);
or U22467 (N_22467,N_21825,N_21944);
nand U22468 (N_22468,N_21984,N_22178);
or U22469 (N_22469,N_22050,N_21617);
nand U22470 (N_22470,N_22167,N_22127);
nand U22471 (N_22471,N_21818,N_21939);
nand U22472 (N_22472,N_21963,N_21855);
and U22473 (N_22473,N_22076,N_21977);
or U22474 (N_22474,N_22012,N_21629);
xnor U22475 (N_22475,N_21759,N_21762);
nand U22476 (N_22476,N_21887,N_22017);
xor U22477 (N_22477,N_21968,N_21805);
and U22478 (N_22478,N_22147,N_21862);
nor U22479 (N_22479,N_21658,N_21925);
nand U22480 (N_22480,N_21901,N_22199);
nor U22481 (N_22481,N_21652,N_22078);
and U22482 (N_22482,N_21619,N_21701);
xnor U22483 (N_22483,N_21923,N_21637);
nor U22484 (N_22484,N_22093,N_22145);
or U22485 (N_22485,N_21694,N_21604);
nor U22486 (N_22486,N_21833,N_21823);
xnor U22487 (N_22487,N_21902,N_22156);
nor U22488 (N_22488,N_21988,N_22152);
xnor U22489 (N_22489,N_21960,N_21654);
nand U22490 (N_22490,N_22146,N_22054);
nor U22491 (N_22491,N_21685,N_21636);
nor U22492 (N_22492,N_22185,N_21705);
and U22493 (N_22493,N_22022,N_21978);
nand U22494 (N_22494,N_22085,N_21647);
xnor U22495 (N_22495,N_21950,N_22113);
xnor U22496 (N_22496,N_22020,N_21935);
nor U22497 (N_22497,N_21903,N_21975);
xor U22498 (N_22498,N_21791,N_22018);
xor U22499 (N_22499,N_21973,N_21642);
nand U22500 (N_22500,N_21844,N_22127);
and U22501 (N_22501,N_21707,N_21947);
nand U22502 (N_22502,N_21744,N_22024);
nand U22503 (N_22503,N_21840,N_21642);
nor U22504 (N_22504,N_22045,N_21829);
nor U22505 (N_22505,N_21950,N_22111);
nand U22506 (N_22506,N_21677,N_22050);
nand U22507 (N_22507,N_22044,N_22178);
or U22508 (N_22508,N_22157,N_21713);
nand U22509 (N_22509,N_22102,N_22015);
or U22510 (N_22510,N_21931,N_21778);
or U22511 (N_22511,N_21604,N_22184);
and U22512 (N_22512,N_22051,N_22127);
and U22513 (N_22513,N_21928,N_21937);
nor U22514 (N_22514,N_21888,N_22045);
or U22515 (N_22515,N_22116,N_22021);
nand U22516 (N_22516,N_21610,N_21649);
and U22517 (N_22517,N_21826,N_21765);
nor U22518 (N_22518,N_21712,N_22016);
or U22519 (N_22519,N_21851,N_22134);
and U22520 (N_22520,N_21607,N_21712);
nor U22521 (N_22521,N_21608,N_22152);
nor U22522 (N_22522,N_21816,N_21675);
and U22523 (N_22523,N_21774,N_21657);
nor U22524 (N_22524,N_21703,N_21654);
and U22525 (N_22525,N_21920,N_21634);
nor U22526 (N_22526,N_21673,N_22076);
nor U22527 (N_22527,N_21617,N_22018);
or U22528 (N_22528,N_22073,N_21829);
nand U22529 (N_22529,N_21643,N_22150);
nor U22530 (N_22530,N_22088,N_21765);
and U22531 (N_22531,N_21628,N_21879);
or U22532 (N_22532,N_21949,N_22017);
nand U22533 (N_22533,N_21835,N_21687);
or U22534 (N_22534,N_22053,N_21847);
or U22535 (N_22535,N_22193,N_21925);
and U22536 (N_22536,N_21976,N_21630);
nand U22537 (N_22537,N_22192,N_21832);
nor U22538 (N_22538,N_21606,N_21961);
and U22539 (N_22539,N_21783,N_22039);
or U22540 (N_22540,N_21899,N_21911);
xnor U22541 (N_22541,N_22042,N_21708);
and U22542 (N_22542,N_21601,N_21625);
nor U22543 (N_22543,N_21659,N_21603);
nand U22544 (N_22544,N_21958,N_21976);
and U22545 (N_22545,N_21748,N_22042);
and U22546 (N_22546,N_22168,N_21956);
and U22547 (N_22547,N_21947,N_22024);
nand U22548 (N_22548,N_22032,N_21799);
or U22549 (N_22549,N_21600,N_22007);
nand U22550 (N_22550,N_22029,N_21988);
nor U22551 (N_22551,N_22154,N_21759);
and U22552 (N_22552,N_22010,N_21927);
or U22553 (N_22553,N_22046,N_21764);
nor U22554 (N_22554,N_21766,N_21656);
and U22555 (N_22555,N_22111,N_22164);
nand U22556 (N_22556,N_21997,N_22118);
and U22557 (N_22557,N_22084,N_21781);
nor U22558 (N_22558,N_21648,N_22114);
nand U22559 (N_22559,N_22049,N_21910);
nor U22560 (N_22560,N_22061,N_21963);
and U22561 (N_22561,N_22131,N_22056);
or U22562 (N_22562,N_22010,N_21945);
nor U22563 (N_22563,N_22150,N_22120);
or U22564 (N_22564,N_22191,N_21855);
or U22565 (N_22565,N_21947,N_21976);
and U22566 (N_22566,N_22178,N_22017);
or U22567 (N_22567,N_21974,N_21765);
nand U22568 (N_22568,N_22149,N_21650);
or U22569 (N_22569,N_21895,N_22110);
and U22570 (N_22570,N_21891,N_21915);
and U22571 (N_22571,N_22045,N_21837);
nand U22572 (N_22572,N_22086,N_22074);
nor U22573 (N_22573,N_21842,N_21941);
nor U22574 (N_22574,N_21868,N_21741);
and U22575 (N_22575,N_21842,N_21616);
or U22576 (N_22576,N_21760,N_21758);
and U22577 (N_22577,N_21664,N_22080);
nand U22578 (N_22578,N_21676,N_22110);
and U22579 (N_22579,N_22097,N_22198);
or U22580 (N_22580,N_22168,N_21935);
nand U22581 (N_22581,N_22112,N_22058);
nand U22582 (N_22582,N_21861,N_22158);
nand U22583 (N_22583,N_22190,N_21953);
or U22584 (N_22584,N_21998,N_21992);
nand U22585 (N_22585,N_22073,N_21667);
and U22586 (N_22586,N_21946,N_21841);
nor U22587 (N_22587,N_21783,N_21809);
nor U22588 (N_22588,N_21841,N_21622);
or U22589 (N_22589,N_21903,N_22032);
nand U22590 (N_22590,N_21627,N_21757);
or U22591 (N_22591,N_22033,N_21631);
and U22592 (N_22592,N_21739,N_21701);
or U22593 (N_22593,N_21713,N_21699);
nor U22594 (N_22594,N_21872,N_21903);
and U22595 (N_22595,N_21862,N_21904);
nand U22596 (N_22596,N_22138,N_21921);
nand U22597 (N_22597,N_22176,N_22002);
nor U22598 (N_22598,N_21639,N_21743);
or U22599 (N_22599,N_21641,N_21639);
nor U22600 (N_22600,N_21957,N_21761);
nor U22601 (N_22601,N_21915,N_21983);
or U22602 (N_22602,N_22026,N_22162);
or U22603 (N_22603,N_21765,N_21755);
xnor U22604 (N_22604,N_22068,N_21790);
nor U22605 (N_22605,N_21703,N_21856);
or U22606 (N_22606,N_22088,N_21613);
and U22607 (N_22607,N_22045,N_21645);
nand U22608 (N_22608,N_21843,N_21822);
or U22609 (N_22609,N_22063,N_21899);
nand U22610 (N_22610,N_21814,N_21802);
nor U22611 (N_22611,N_21845,N_21685);
and U22612 (N_22612,N_21970,N_22199);
xnor U22613 (N_22613,N_22118,N_22126);
xnor U22614 (N_22614,N_22005,N_21759);
nand U22615 (N_22615,N_21670,N_21621);
nor U22616 (N_22616,N_21613,N_22167);
and U22617 (N_22617,N_21809,N_21626);
nor U22618 (N_22618,N_21780,N_21769);
xor U22619 (N_22619,N_21830,N_21934);
nand U22620 (N_22620,N_21956,N_22072);
nand U22621 (N_22621,N_21719,N_21948);
nor U22622 (N_22622,N_22114,N_21798);
and U22623 (N_22623,N_22039,N_22191);
xnor U22624 (N_22624,N_22141,N_21635);
and U22625 (N_22625,N_22137,N_22143);
nor U22626 (N_22626,N_21768,N_22111);
or U22627 (N_22627,N_22059,N_21930);
or U22628 (N_22628,N_22126,N_21676);
or U22629 (N_22629,N_21881,N_21886);
nor U22630 (N_22630,N_21823,N_21650);
and U22631 (N_22631,N_22156,N_22017);
nand U22632 (N_22632,N_22033,N_21804);
and U22633 (N_22633,N_22171,N_22033);
nor U22634 (N_22634,N_21781,N_22098);
and U22635 (N_22635,N_22106,N_22082);
nor U22636 (N_22636,N_21804,N_21910);
and U22637 (N_22637,N_21627,N_21895);
nor U22638 (N_22638,N_21842,N_21900);
nand U22639 (N_22639,N_21889,N_21993);
and U22640 (N_22640,N_21729,N_22156);
nand U22641 (N_22641,N_22119,N_22126);
and U22642 (N_22642,N_21623,N_22130);
and U22643 (N_22643,N_21890,N_21812);
nor U22644 (N_22644,N_22142,N_21653);
nor U22645 (N_22645,N_21650,N_22023);
or U22646 (N_22646,N_21622,N_21864);
nand U22647 (N_22647,N_21733,N_21899);
xnor U22648 (N_22648,N_22198,N_21666);
or U22649 (N_22649,N_22043,N_21845);
nand U22650 (N_22650,N_21987,N_21935);
nor U22651 (N_22651,N_21892,N_21779);
xor U22652 (N_22652,N_21725,N_21685);
or U22653 (N_22653,N_22135,N_22062);
nor U22654 (N_22654,N_21762,N_21800);
or U22655 (N_22655,N_21637,N_22098);
nor U22656 (N_22656,N_22002,N_21729);
and U22657 (N_22657,N_22021,N_21690);
xor U22658 (N_22658,N_21655,N_21906);
nor U22659 (N_22659,N_22190,N_21603);
or U22660 (N_22660,N_22017,N_21765);
and U22661 (N_22661,N_21630,N_22024);
and U22662 (N_22662,N_22101,N_21827);
xnor U22663 (N_22663,N_21771,N_21649);
xor U22664 (N_22664,N_21678,N_21687);
xnor U22665 (N_22665,N_22159,N_22064);
and U22666 (N_22666,N_21802,N_21875);
nand U22667 (N_22667,N_21750,N_21732);
or U22668 (N_22668,N_21836,N_21778);
or U22669 (N_22669,N_21931,N_21824);
and U22670 (N_22670,N_21993,N_22104);
nor U22671 (N_22671,N_21964,N_21837);
nor U22672 (N_22672,N_21666,N_21816);
nand U22673 (N_22673,N_21924,N_21889);
nor U22674 (N_22674,N_21810,N_21790);
and U22675 (N_22675,N_22187,N_22030);
or U22676 (N_22676,N_21957,N_21929);
nand U22677 (N_22677,N_21638,N_21678);
or U22678 (N_22678,N_22095,N_22181);
nor U22679 (N_22679,N_22059,N_21740);
xnor U22680 (N_22680,N_21776,N_21618);
nor U22681 (N_22681,N_21747,N_21948);
nand U22682 (N_22682,N_22180,N_21885);
or U22683 (N_22683,N_21770,N_21675);
or U22684 (N_22684,N_21631,N_21741);
or U22685 (N_22685,N_22024,N_22157);
nor U22686 (N_22686,N_21849,N_22176);
or U22687 (N_22687,N_21650,N_21887);
or U22688 (N_22688,N_21955,N_21676);
nand U22689 (N_22689,N_21765,N_21893);
nand U22690 (N_22690,N_21946,N_22159);
or U22691 (N_22691,N_22197,N_22003);
nand U22692 (N_22692,N_22020,N_21885);
and U22693 (N_22693,N_22149,N_22090);
xnor U22694 (N_22694,N_21746,N_21788);
and U22695 (N_22695,N_21717,N_21696);
nor U22696 (N_22696,N_21610,N_21828);
nand U22697 (N_22697,N_21768,N_21757);
and U22698 (N_22698,N_21853,N_21665);
xnor U22699 (N_22699,N_21826,N_22167);
and U22700 (N_22700,N_21618,N_21809);
nand U22701 (N_22701,N_21688,N_21621);
and U22702 (N_22702,N_21780,N_21969);
or U22703 (N_22703,N_21607,N_21699);
nand U22704 (N_22704,N_22104,N_22128);
nor U22705 (N_22705,N_21631,N_21876);
nand U22706 (N_22706,N_21836,N_21660);
nor U22707 (N_22707,N_21790,N_21693);
and U22708 (N_22708,N_22149,N_21818);
or U22709 (N_22709,N_21733,N_22138);
nor U22710 (N_22710,N_21771,N_21961);
or U22711 (N_22711,N_22051,N_21805);
and U22712 (N_22712,N_21779,N_21898);
or U22713 (N_22713,N_21684,N_21872);
and U22714 (N_22714,N_21881,N_22120);
or U22715 (N_22715,N_21903,N_21822);
and U22716 (N_22716,N_22041,N_21718);
nor U22717 (N_22717,N_22165,N_21986);
xnor U22718 (N_22718,N_21974,N_22046);
nor U22719 (N_22719,N_22018,N_21975);
nand U22720 (N_22720,N_22118,N_22038);
and U22721 (N_22721,N_21662,N_21720);
or U22722 (N_22722,N_21777,N_21856);
nor U22723 (N_22723,N_21810,N_21745);
nand U22724 (N_22724,N_21746,N_21615);
nor U22725 (N_22725,N_21708,N_21843);
and U22726 (N_22726,N_21964,N_21757);
and U22727 (N_22727,N_21987,N_21712);
and U22728 (N_22728,N_21690,N_21954);
nand U22729 (N_22729,N_22170,N_22193);
nand U22730 (N_22730,N_21984,N_21677);
nand U22731 (N_22731,N_22158,N_21723);
nand U22732 (N_22732,N_21625,N_21886);
nand U22733 (N_22733,N_21946,N_22041);
or U22734 (N_22734,N_21630,N_21744);
xor U22735 (N_22735,N_21605,N_21900);
and U22736 (N_22736,N_21636,N_21628);
and U22737 (N_22737,N_21627,N_21614);
and U22738 (N_22738,N_21657,N_22185);
xor U22739 (N_22739,N_22015,N_21745);
and U22740 (N_22740,N_21855,N_21872);
nor U22741 (N_22741,N_21867,N_22105);
nor U22742 (N_22742,N_21670,N_22040);
or U22743 (N_22743,N_22004,N_22086);
nand U22744 (N_22744,N_22123,N_21715);
nand U22745 (N_22745,N_22024,N_22195);
and U22746 (N_22746,N_22138,N_21628);
nand U22747 (N_22747,N_21750,N_21919);
or U22748 (N_22748,N_21605,N_22010);
nor U22749 (N_22749,N_21982,N_22182);
or U22750 (N_22750,N_21677,N_21628);
xnor U22751 (N_22751,N_22037,N_21743);
nand U22752 (N_22752,N_22018,N_21795);
nor U22753 (N_22753,N_21637,N_21898);
or U22754 (N_22754,N_21629,N_21857);
or U22755 (N_22755,N_21686,N_21761);
xor U22756 (N_22756,N_22061,N_21634);
nand U22757 (N_22757,N_21740,N_22118);
xnor U22758 (N_22758,N_21646,N_21945);
xor U22759 (N_22759,N_22133,N_21835);
nand U22760 (N_22760,N_21669,N_22124);
nand U22761 (N_22761,N_21978,N_21979);
and U22762 (N_22762,N_22063,N_21650);
nand U22763 (N_22763,N_21965,N_21934);
xnor U22764 (N_22764,N_21814,N_21726);
or U22765 (N_22765,N_22129,N_21914);
and U22766 (N_22766,N_22166,N_22052);
or U22767 (N_22767,N_22157,N_22055);
and U22768 (N_22768,N_22181,N_22035);
or U22769 (N_22769,N_21863,N_21961);
nor U22770 (N_22770,N_21779,N_21910);
or U22771 (N_22771,N_21790,N_22087);
xor U22772 (N_22772,N_21740,N_22193);
nand U22773 (N_22773,N_21912,N_21908);
nor U22774 (N_22774,N_21979,N_22092);
nor U22775 (N_22775,N_21800,N_21789);
nand U22776 (N_22776,N_21866,N_22179);
nor U22777 (N_22777,N_21897,N_21762);
nor U22778 (N_22778,N_21810,N_21789);
or U22779 (N_22779,N_21638,N_21761);
nor U22780 (N_22780,N_22076,N_22175);
and U22781 (N_22781,N_22136,N_21704);
nor U22782 (N_22782,N_21807,N_21737);
or U22783 (N_22783,N_21626,N_21988);
nor U22784 (N_22784,N_21999,N_21800);
nand U22785 (N_22785,N_21707,N_22017);
nor U22786 (N_22786,N_22154,N_21691);
nor U22787 (N_22787,N_22056,N_22168);
xor U22788 (N_22788,N_22075,N_21931);
or U22789 (N_22789,N_21976,N_21769);
nor U22790 (N_22790,N_21806,N_22179);
nor U22791 (N_22791,N_22151,N_22026);
nor U22792 (N_22792,N_21652,N_21678);
and U22793 (N_22793,N_21798,N_22050);
and U22794 (N_22794,N_21916,N_21803);
nand U22795 (N_22795,N_21680,N_21646);
nand U22796 (N_22796,N_21980,N_22069);
and U22797 (N_22797,N_21922,N_21625);
nand U22798 (N_22798,N_21652,N_21693);
and U22799 (N_22799,N_22007,N_22155);
nor U22800 (N_22800,N_22575,N_22652);
or U22801 (N_22801,N_22689,N_22214);
or U22802 (N_22802,N_22283,N_22375);
and U22803 (N_22803,N_22626,N_22237);
nor U22804 (N_22804,N_22667,N_22372);
and U22805 (N_22805,N_22329,N_22202);
and U22806 (N_22806,N_22728,N_22712);
xnor U22807 (N_22807,N_22785,N_22479);
nand U22808 (N_22808,N_22755,N_22619);
nand U22809 (N_22809,N_22484,N_22752);
nand U22810 (N_22810,N_22271,N_22680);
xor U22811 (N_22811,N_22360,N_22552);
or U22812 (N_22812,N_22522,N_22673);
nand U22813 (N_22813,N_22705,N_22394);
nor U22814 (N_22814,N_22393,N_22465);
nor U22815 (N_22815,N_22747,N_22316);
nor U22816 (N_22816,N_22299,N_22563);
or U22817 (N_22817,N_22562,N_22649);
and U22818 (N_22818,N_22604,N_22226);
or U22819 (N_22819,N_22487,N_22711);
nor U22820 (N_22820,N_22401,N_22606);
and U22821 (N_22821,N_22352,N_22421);
or U22822 (N_22822,N_22249,N_22732);
and U22823 (N_22823,N_22654,N_22751);
and U22824 (N_22824,N_22485,N_22456);
or U22825 (N_22825,N_22742,N_22405);
xor U22826 (N_22826,N_22235,N_22684);
nand U22827 (N_22827,N_22764,N_22605);
nor U22828 (N_22828,N_22277,N_22679);
or U22829 (N_22829,N_22592,N_22525);
nand U22830 (N_22830,N_22453,N_22433);
nor U22831 (N_22831,N_22641,N_22313);
nand U22832 (N_22832,N_22560,N_22501);
or U22833 (N_22833,N_22591,N_22681);
nand U22834 (N_22834,N_22507,N_22767);
and U22835 (N_22835,N_22784,N_22266);
nand U22836 (N_22836,N_22726,N_22279);
nand U22837 (N_22837,N_22451,N_22642);
or U22838 (N_22838,N_22746,N_22765);
and U22839 (N_22839,N_22454,N_22725);
nor U22840 (N_22840,N_22416,N_22212);
nand U22841 (N_22841,N_22207,N_22583);
and U22842 (N_22842,N_22596,N_22607);
xor U22843 (N_22843,N_22611,N_22753);
and U22844 (N_22844,N_22512,N_22386);
or U22845 (N_22845,N_22276,N_22253);
or U22846 (N_22846,N_22661,N_22568);
nor U22847 (N_22847,N_22263,N_22796);
and U22848 (N_22848,N_22458,N_22448);
nor U22849 (N_22849,N_22534,N_22584);
and U22850 (N_22850,N_22308,N_22520);
and U22851 (N_22851,N_22398,N_22208);
nor U22852 (N_22852,N_22224,N_22788);
or U22853 (N_22853,N_22213,N_22422);
nand U22854 (N_22854,N_22706,N_22380);
nand U22855 (N_22855,N_22444,N_22466);
and U22856 (N_22856,N_22566,N_22757);
nor U22857 (N_22857,N_22221,N_22690);
nor U22858 (N_22858,N_22797,N_22325);
and U22859 (N_22859,N_22735,N_22531);
or U22860 (N_22860,N_22762,N_22406);
nand U22861 (N_22861,N_22232,N_22574);
or U22862 (N_22862,N_22216,N_22546);
or U22863 (N_22863,N_22709,N_22290);
and U22864 (N_22864,N_22419,N_22505);
nor U22865 (N_22865,N_22662,N_22715);
nand U22866 (N_22866,N_22252,N_22514);
or U22867 (N_22867,N_22340,N_22473);
or U22868 (N_22868,N_22353,N_22238);
nor U22869 (N_22869,N_22675,N_22723);
xnor U22870 (N_22870,N_22257,N_22532);
nand U22871 (N_22871,N_22341,N_22286);
nand U22872 (N_22872,N_22663,N_22293);
nor U22873 (N_22873,N_22786,N_22287);
nand U22874 (N_22874,N_22339,N_22550);
nor U22875 (N_22875,N_22326,N_22586);
or U22876 (N_22876,N_22389,N_22270);
xnor U22877 (N_22877,N_22506,N_22775);
or U22878 (N_22878,N_22612,N_22660);
nand U22879 (N_22879,N_22200,N_22640);
xor U22880 (N_22880,N_22536,N_22687);
nor U22881 (N_22881,N_22542,N_22518);
nor U22882 (N_22882,N_22646,N_22510);
nor U22883 (N_22883,N_22582,N_22631);
or U22884 (N_22884,N_22248,N_22215);
nand U22885 (N_22885,N_22634,N_22436);
and U22886 (N_22886,N_22678,N_22616);
nand U22887 (N_22887,N_22384,N_22537);
nand U22888 (N_22888,N_22504,N_22256);
xor U22889 (N_22889,N_22599,N_22557);
or U22890 (N_22890,N_22332,N_22624);
nand U22891 (N_22891,N_22328,N_22378);
nor U22892 (N_22892,N_22264,N_22201);
and U22893 (N_22893,N_22637,N_22701);
nand U22894 (N_22894,N_22603,N_22269);
nand U22895 (N_22895,N_22569,N_22744);
nand U22896 (N_22896,N_22553,N_22615);
and U22897 (N_22897,N_22338,N_22704);
nand U22898 (N_22898,N_22243,N_22296);
and U22899 (N_22899,N_22478,N_22435);
or U22900 (N_22900,N_22301,N_22486);
nor U22901 (N_22901,N_22399,N_22390);
or U22902 (N_22902,N_22239,N_22539);
nand U22903 (N_22903,N_22260,N_22364);
nor U22904 (N_22904,N_22502,N_22674);
or U22905 (N_22905,N_22609,N_22628);
and U22906 (N_22906,N_22209,N_22242);
or U22907 (N_22907,N_22524,N_22585);
and U22908 (N_22908,N_22227,N_22648);
and U22909 (N_22909,N_22424,N_22490);
nor U22910 (N_22910,N_22371,N_22432);
xor U22911 (N_22911,N_22570,N_22408);
nor U22912 (N_22912,N_22695,N_22685);
nor U22913 (N_22913,N_22217,N_22736);
nand U22914 (N_22914,N_22267,N_22545);
nand U22915 (N_22915,N_22666,N_22298);
or U22916 (N_22916,N_22733,N_22443);
nand U22917 (N_22917,N_22468,N_22403);
and U22918 (N_22918,N_22288,N_22638);
nor U22919 (N_22919,N_22431,N_22556);
and U22920 (N_22920,N_22770,N_22409);
nor U22921 (N_22921,N_22282,N_22356);
and U22922 (N_22922,N_22411,N_22551);
nor U22923 (N_22923,N_22791,N_22750);
or U22924 (N_22924,N_22668,N_22721);
or U22925 (N_22925,N_22348,N_22359);
nor U22926 (N_22926,N_22320,N_22349);
or U22927 (N_22927,N_22740,N_22460);
nor U22928 (N_22928,N_22598,N_22608);
or U22929 (N_22929,N_22315,N_22295);
nand U22930 (N_22930,N_22474,N_22677);
nand U22931 (N_22931,N_22657,N_22331);
nor U22932 (N_22932,N_22759,N_22676);
nand U22933 (N_22933,N_22776,N_22400);
nand U22934 (N_22934,N_22392,N_22697);
and U22935 (N_22935,N_22768,N_22467);
nand U22936 (N_22936,N_22610,N_22795);
nand U22937 (N_22937,N_22577,N_22730);
or U22938 (N_22938,N_22481,N_22529);
nor U22939 (N_22939,N_22727,N_22255);
nand U22940 (N_22940,N_22643,N_22494);
nand U22941 (N_22941,N_22731,N_22368);
or U22942 (N_22942,N_22622,N_22787);
nor U22943 (N_22943,N_22285,N_22700);
and U22944 (N_22944,N_22457,N_22312);
nand U22945 (N_22945,N_22639,N_22627);
nand U22946 (N_22946,N_22449,N_22655);
nand U22947 (N_22947,N_22554,N_22330);
nand U22948 (N_22948,N_22720,N_22523);
and U22949 (N_22949,N_22541,N_22683);
nand U22950 (N_22950,N_22305,N_22410);
or U22951 (N_22951,N_22650,N_22691);
or U22952 (N_22952,N_22749,N_22345);
xnor U22953 (N_22953,N_22278,N_22722);
nor U22954 (N_22954,N_22636,N_22475);
or U22955 (N_22955,N_22304,N_22713);
or U22956 (N_22956,N_22373,N_22220);
or U22957 (N_22957,N_22420,N_22632);
or U22958 (N_22958,N_22576,N_22588);
or U22959 (N_22959,N_22223,N_22633);
and U22960 (N_22960,N_22777,N_22397);
nor U22961 (N_22961,N_22710,N_22236);
nand U22962 (N_22962,N_22635,N_22307);
nor U22963 (N_22963,N_22404,N_22210);
or U22964 (N_22964,N_22580,N_22280);
or U22965 (N_22965,N_22365,N_22517);
nand U22966 (N_22966,N_22273,N_22387);
or U22967 (N_22967,N_22707,N_22488);
or U22968 (N_22968,N_22528,N_22559);
or U22969 (N_22969,N_22565,N_22760);
xor U22970 (N_22970,N_22461,N_22464);
nor U22971 (N_22971,N_22672,N_22245);
nand U22972 (N_22972,N_22521,N_22388);
or U22973 (N_22973,N_22363,N_22427);
nor U22974 (N_22974,N_22761,N_22218);
nand U22975 (N_22975,N_22737,N_22367);
nand U22976 (N_22976,N_22254,N_22423);
and U22977 (N_22977,N_22347,N_22602);
nor U22978 (N_22978,N_22743,N_22780);
xnor U22979 (N_22979,N_22434,N_22548);
nand U22980 (N_22980,N_22513,N_22319);
and U22981 (N_22981,N_22440,N_22342);
xnor U22982 (N_22982,N_22503,N_22758);
or U22983 (N_22983,N_22555,N_22211);
nor U22984 (N_22984,N_22450,N_22284);
xor U22985 (N_22985,N_22272,N_22561);
nor U22986 (N_22986,N_22206,N_22527);
or U22987 (N_22987,N_22385,N_22739);
nor U22988 (N_22988,N_22425,N_22274);
and U22989 (N_22989,N_22333,N_22578);
xor U22990 (N_22990,N_22600,N_22265);
nor U22991 (N_22991,N_22754,N_22703);
or U22992 (N_22992,N_22289,N_22601);
or U22993 (N_22993,N_22292,N_22799);
or U22994 (N_22994,N_22439,N_22794);
or U22995 (N_22995,N_22516,N_22558);
nor U22996 (N_22996,N_22446,N_22669);
xor U22997 (N_22997,N_22623,N_22294);
nand U22998 (N_22998,N_22708,N_22509);
nor U22999 (N_22999,N_22590,N_22366);
and U23000 (N_23000,N_22250,N_22477);
or U23001 (N_23001,N_22480,N_22745);
or U23002 (N_23002,N_22225,N_22718);
or U23003 (N_23003,N_22682,N_22738);
nand U23004 (N_23004,N_22204,N_22258);
nand U23005 (N_23005,N_22547,N_22515);
and U23006 (N_23006,N_22716,N_22589);
or U23007 (N_23007,N_22219,N_22724);
or U23008 (N_23008,N_22205,N_22476);
xor U23009 (N_23009,N_22381,N_22459);
xor U23010 (N_23010,N_22396,N_22593);
and U23011 (N_23011,N_22694,N_22350);
xnor U23012 (N_23012,N_22595,N_22262);
nand U23013 (N_23013,N_22617,N_22658);
nor U23014 (N_23014,N_22698,N_22798);
xor U23015 (N_23015,N_22621,N_22361);
nand U23016 (N_23016,N_22463,N_22544);
or U23017 (N_23017,N_22748,N_22259);
nor U23018 (N_23018,N_22343,N_22418);
or U23019 (N_23019,N_22229,N_22354);
and U23020 (N_23020,N_22246,N_22355);
and U23021 (N_23021,N_22664,N_22358);
or U23022 (N_23022,N_22379,N_22630);
nand U23023 (N_23023,N_22414,N_22251);
and U23024 (N_23024,N_22572,N_22491);
or U23025 (N_23025,N_22769,N_22686);
or U23026 (N_23026,N_22564,N_22344);
or U23027 (N_23027,N_22702,N_22793);
nand U23028 (N_23028,N_22659,N_22581);
or U23029 (N_23029,N_22651,N_22222);
nor U23030 (N_23030,N_22370,N_22543);
xnor U23031 (N_23031,N_22377,N_22309);
nor U23032 (N_23032,N_22773,N_22645);
and U23033 (N_23033,N_22442,N_22228);
nand U23034 (N_23034,N_22597,N_22782);
nand U23035 (N_23035,N_22535,N_22644);
nor U23036 (N_23036,N_22383,N_22779);
or U23037 (N_23037,N_22496,N_22625);
and U23038 (N_23038,N_22571,N_22376);
xor U23039 (N_23039,N_22268,N_22734);
or U23040 (N_23040,N_22653,N_22241);
and U23041 (N_23041,N_22323,N_22493);
nor U23042 (N_23042,N_22362,N_22500);
nand U23043 (N_23043,N_22346,N_22321);
nor U23044 (N_23044,N_22311,N_22413);
and U23045 (N_23045,N_22692,N_22511);
nor U23046 (N_23046,N_22526,N_22412);
or U23047 (N_23047,N_22324,N_22756);
and U23048 (N_23048,N_22437,N_22233);
nand U23049 (N_23049,N_22447,N_22567);
nand U23050 (N_23050,N_22303,N_22291);
and U23051 (N_23051,N_22441,N_22771);
and U23052 (N_23052,N_22471,N_22455);
and U23053 (N_23053,N_22497,N_22470);
and U23054 (N_23054,N_22402,N_22337);
nand U23055 (N_23055,N_22766,N_22300);
nand U23056 (N_23056,N_22335,N_22774);
and U23057 (N_23057,N_22573,N_22391);
or U23058 (N_23058,N_22415,N_22462);
nand U23059 (N_23059,N_22314,N_22763);
and U23060 (N_23060,N_22789,N_22445);
nand U23061 (N_23061,N_22336,N_22696);
nor U23062 (N_23062,N_22613,N_22483);
and U23063 (N_23063,N_22719,N_22647);
and U23064 (N_23064,N_22428,N_22469);
and U23065 (N_23065,N_22247,N_22489);
and U23066 (N_23066,N_22374,N_22369);
or U23067 (N_23067,N_22318,N_22203);
nor U23068 (N_23068,N_22549,N_22540);
and U23069 (N_23069,N_22482,N_22614);
nand U23070 (N_23070,N_22281,N_22620);
and U23071 (N_23071,N_22519,N_22327);
or U23072 (N_23072,N_22357,N_22472);
or U23073 (N_23073,N_22240,N_22729);
and U23074 (N_23074,N_22790,N_22688);
nand U23075 (N_23075,N_22230,N_22275);
or U23076 (N_23076,N_22231,N_22438);
and U23077 (N_23077,N_22302,N_22498);
nor U23078 (N_23078,N_22407,N_22430);
nor U23079 (N_23079,N_22426,N_22317);
nand U23080 (N_23080,N_22656,N_22310);
or U23081 (N_23081,N_22693,N_22417);
and U23082 (N_23082,N_22778,N_22772);
nor U23083 (N_23083,N_22334,N_22781);
nand U23084 (N_23084,N_22508,N_22714);
nor U23085 (N_23085,N_22261,N_22618);
or U23086 (N_23086,N_22395,N_22579);
and U23087 (N_23087,N_22306,N_22499);
or U23088 (N_23088,N_22538,N_22670);
nand U23089 (N_23089,N_22665,N_22244);
xor U23090 (N_23090,N_22587,N_22234);
nor U23091 (N_23091,N_22629,N_22322);
or U23092 (N_23092,N_22492,N_22594);
nor U23093 (N_23093,N_22382,N_22495);
xnor U23094 (N_23094,N_22533,N_22783);
and U23095 (N_23095,N_22530,N_22792);
xor U23096 (N_23096,N_22671,N_22429);
and U23097 (N_23097,N_22297,N_22452);
nor U23098 (N_23098,N_22741,N_22351);
nor U23099 (N_23099,N_22717,N_22699);
or U23100 (N_23100,N_22403,N_22755);
or U23101 (N_23101,N_22726,N_22238);
nor U23102 (N_23102,N_22493,N_22479);
nor U23103 (N_23103,N_22343,N_22550);
xor U23104 (N_23104,N_22517,N_22695);
or U23105 (N_23105,N_22265,N_22421);
or U23106 (N_23106,N_22730,N_22792);
and U23107 (N_23107,N_22312,N_22559);
or U23108 (N_23108,N_22547,N_22569);
or U23109 (N_23109,N_22365,N_22341);
nor U23110 (N_23110,N_22372,N_22683);
or U23111 (N_23111,N_22205,N_22366);
nand U23112 (N_23112,N_22515,N_22461);
or U23113 (N_23113,N_22377,N_22267);
nor U23114 (N_23114,N_22703,N_22336);
xnor U23115 (N_23115,N_22754,N_22788);
and U23116 (N_23116,N_22202,N_22225);
or U23117 (N_23117,N_22705,N_22282);
nand U23118 (N_23118,N_22757,N_22598);
or U23119 (N_23119,N_22482,N_22789);
nor U23120 (N_23120,N_22650,N_22516);
or U23121 (N_23121,N_22675,N_22651);
and U23122 (N_23122,N_22660,N_22520);
xor U23123 (N_23123,N_22223,N_22277);
nand U23124 (N_23124,N_22354,N_22761);
nor U23125 (N_23125,N_22281,N_22697);
nand U23126 (N_23126,N_22329,N_22669);
nand U23127 (N_23127,N_22650,N_22565);
nand U23128 (N_23128,N_22523,N_22556);
nand U23129 (N_23129,N_22237,N_22542);
nand U23130 (N_23130,N_22772,N_22525);
or U23131 (N_23131,N_22566,N_22379);
and U23132 (N_23132,N_22769,N_22681);
or U23133 (N_23133,N_22377,N_22667);
nand U23134 (N_23134,N_22674,N_22408);
nor U23135 (N_23135,N_22642,N_22799);
nor U23136 (N_23136,N_22251,N_22362);
nand U23137 (N_23137,N_22614,N_22275);
and U23138 (N_23138,N_22406,N_22537);
nand U23139 (N_23139,N_22417,N_22513);
or U23140 (N_23140,N_22241,N_22288);
xor U23141 (N_23141,N_22333,N_22743);
nor U23142 (N_23142,N_22408,N_22416);
or U23143 (N_23143,N_22384,N_22672);
xnor U23144 (N_23144,N_22634,N_22788);
and U23145 (N_23145,N_22670,N_22471);
nand U23146 (N_23146,N_22514,N_22691);
or U23147 (N_23147,N_22248,N_22672);
nand U23148 (N_23148,N_22403,N_22421);
nor U23149 (N_23149,N_22478,N_22419);
or U23150 (N_23150,N_22370,N_22493);
and U23151 (N_23151,N_22367,N_22594);
and U23152 (N_23152,N_22585,N_22780);
nor U23153 (N_23153,N_22320,N_22331);
xnor U23154 (N_23154,N_22575,N_22202);
nand U23155 (N_23155,N_22747,N_22710);
nand U23156 (N_23156,N_22441,N_22489);
and U23157 (N_23157,N_22765,N_22757);
nor U23158 (N_23158,N_22428,N_22541);
and U23159 (N_23159,N_22380,N_22223);
or U23160 (N_23160,N_22269,N_22503);
nand U23161 (N_23161,N_22566,N_22763);
and U23162 (N_23162,N_22298,N_22228);
or U23163 (N_23163,N_22706,N_22404);
or U23164 (N_23164,N_22693,N_22705);
nor U23165 (N_23165,N_22515,N_22235);
nor U23166 (N_23166,N_22626,N_22787);
xor U23167 (N_23167,N_22659,N_22643);
xor U23168 (N_23168,N_22417,N_22432);
nand U23169 (N_23169,N_22716,N_22564);
nand U23170 (N_23170,N_22349,N_22302);
or U23171 (N_23171,N_22340,N_22660);
nand U23172 (N_23172,N_22254,N_22683);
xnor U23173 (N_23173,N_22677,N_22263);
nand U23174 (N_23174,N_22414,N_22515);
and U23175 (N_23175,N_22779,N_22295);
nand U23176 (N_23176,N_22393,N_22640);
nor U23177 (N_23177,N_22283,N_22360);
nor U23178 (N_23178,N_22634,N_22459);
nor U23179 (N_23179,N_22421,N_22511);
nand U23180 (N_23180,N_22383,N_22625);
or U23181 (N_23181,N_22636,N_22502);
and U23182 (N_23182,N_22606,N_22223);
xor U23183 (N_23183,N_22206,N_22777);
nor U23184 (N_23184,N_22436,N_22728);
nor U23185 (N_23185,N_22257,N_22715);
nand U23186 (N_23186,N_22799,N_22490);
nand U23187 (N_23187,N_22705,N_22254);
or U23188 (N_23188,N_22633,N_22661);
or U23189 (N_23189,N_22355,N_22740);
xnor U23190 (N_23190,N_22751,N_22463);
xor U23191 (N_23191,N_22271,N_22718);
nand U23192 (N_23192,N_22693,N_22315);
nand U23193 (N_23193,N_22735,N_22264);
or U23194 (N_23194,N_22580,N_22346);
nor U23195 (N_23195,N_22612,N_22375);
nand U23196 (N_23196,N_22633,N_22250);
nor U23197 (N_23197,N_22695,N_22623);
and U23198 (N_23198,N_22710,N_22322);
xor U23199 (N_23199,N_22368,N_22535);
or U23200 (N_23200,N_22438,N_22400);
nor U23201 (N_23201,N_22521,N_22706);
nor U23202 (N_23202,N_22241,N_22385);
nor U23203 (N_23203,N_22631,N_22336);
xor U23204 (N_23204,N_22481,N_22466);
nor U23205 (N_23205,N_22318,N_22290);
and U23206 (N_23206,N_22603,N_22220);
nor U23207 (N_23207,N_22711,N_22289);
nand U23208 (N_23208,N_22773,N_22663);
nor U23209 (N_23209,N_22782,N_22659);
or U23210 (N_23210,N_22321,N_22705);
and U23211 (N_23211,N_22440,N_22708);
or U23212 (N_23212,N_22241,N_22327);
or U23213 (N_23213,N_22241,N_22767);
and U23214 (N_23214,N_22403,N_22395);
xor U23215 (N_23215,N_22756,N_22769);
or U23216 (N_23216,N_22461,N_22254);
nand U23217 (N_23217,N_22485,N_22368);
nor U23218 (N_23218,N_22241,N_22599);
or U23219 (N_23219,N_22223,N_22783);
nor U23220 (N_23220,N_22229,N_22723);
and U23221 (N_23221,N_22586,N_22696);
xnor U23222 (N_23222,N_22639,N_22473);
and U23223 (N_23223,N_22536,N_22601);
or U23224 (N_23224,N_22784,N_22524);
or U23225 (N_23225,N_22673,N_22237);
nor U23226 (N_23226,N_22587,N_22586);
nand U23227 (N_23227,N_22706,N_22774);
or U23228 (N_23228,N_22707,N_22501);
nand U23229 (N_23229,N_22350,N_22477);
and U23230 (N_23230,N_22733,N_22519);
nor U23231 (N_23231,N_22632,N_22261);
and U23232 (N_23232,N_22653,N_22488);
and U23233 (N_23233,N_22225,N_22771);
nand U23234 (N_23234,N_22209,N_22222);
and U23235 (N_23235,N_22752,N_22368);
xnor U23236 (N_23236,N_22710,N_22677);
and U23237 (N_23237,N_22527,N_22394);
and U23238 (N_23238,N_22761,N_22608);
xor U23239 (N_23239,N_22237,N_22319);
or U23240 (N_23240,N_22750,N_22637);
nand U23241 (N_23241,N_22435,N_22503);
nor U23242 (N_23242,N_22667,N_22696);
nand U23243 (N_23243,N_22515,N_22718);
nand U23244 (N_23244,N_22362,N_22314);
nand U23245 (N_23245,N_22349,N_22734);
nor U23246 (N_23246,N_22775,N_22342);
or U23247 (N_23247,N_22699,N_22457);
xor U23248 (N_23248,N_22426,N_22241);
or U23249 (N_23249,N_22714,N_22780);
nor U23250 (N_23250,N_22208,N_22707);
and U23251 (N_23251,N_22549,N_22672);
nand U23252 (N_23252,N_22722,N_22653);
xnor U23253 (N_23253,N_22601,N_22605);
and U23254 (N_23254,N_22313,N_22627);
or U23255 (N_23255,N_22538,N_22368);
nand U23256 (N_23256,N_22354,N_22765);
nand U23257 (N_23257,N_22304,N_22523);
or U23258 (N_23258,N_22624,N_22619);
or U23259 (N_23259,N_22684,N_22600);
nor U23260 (N_23260,N_22475,N_22304);
nor U23261 (N_23261,N_22205,N_22540);
nor U23262 (N_23262,N_22792,N_22782);
or U23263 (N_23263,N_22487,N_22331);
nand U23264 (N_23264,N_22354,N_22386);
nor U23265 (N_23265,N_22372,N_22609);
nor U23266 (N_23266,N_22521,N_22571);
xnor U23267 (N_23267,N_22738,N_22371);
nand U23268 (N_23268,N_22367,N_22728);
or U23269 (N_23269,N_22483,N_22358);
nand U23270 (N_23270,N_22305,N_22277);
nor U23271 (N_23271,N_22789,N_22494);
nor U23272 (N_23272,N_22662,N_22380);
and U23273 (N_23273,N_22289,N_22210);
nor U23274 (N_23274,N_22203,N_22748);
xor U23275 (N_23275,N_22432,N_22363);
nor U23276 (N_23276,N_22706,N_22264);
and U23277 (N_23277,N_22408,N_22794);
nor U23278 (N_23278,N_22270,N_22268);
and U23279 (N_23279,N_22647,N_22323);
or U23280 (N_23280,N_22271,N_22482);
nor U23281 (N_23281,N_22506,N_22534);
and U23282 (N_23282,N_22608,N_22314);
or U23283 (N_23283,N_22780,N_22475);
xor U23284 (N_23284,N_22730,N_22510);
or U23285 (N_23285,N_22550,N_22769);
and U23286 (N_23286,N_22470,N_22208);
nor U23287 (N_23287,N_22507,N_22413);
and U23288 (N_23288,N_22668,N_22342);
and U23289 (N_23289,N_22713,N_22229);
nor U23290 (N_23290,N_22683,N_22654);
and U23291 (N_23291,N_22482,N_22569);
nand U23292 (N_23292,N_22287,N_22609);
nand U23293 (N_23293,N_22794,N_22587);
or U23294 (N_23294,N_22306,N_22309);
and U23295 (N_23295,N_22511,N_22526);
nor U23296 (N_23296,N_22569,N_22554);
and U23297 (N_23297,N_22672,N_22774);
and U23298 (N_23298,N_22287,N_22258);
or U23299 (N_23299,N_22536,N_22533);
and U23300 (N_23300,N_22218,N_22220);
or U23301 (N_23301,N_22527,N_22583);
nand U23302 (N_23302,N_22514,N_22323);
or U23303 (N_23303,N_22525,N_22312);
and U23304 (N_23304,N_22756,N_22356);
and U23305 (N_23305,N_22662,N_22589);
nand U23306 (N_23306,N_22662,N_22455);
nand U23307 (N_23307,N_22704,N_22459);
and U23308 (N_23308,N_22540,N_22612);
xor U23309 (N_23309,N_22249,N_22406);
and U23310 (N_23310,N_22473,N_22692);
nor U23311 (N_23311,N_22764,N_22627);
and U23312 (N_23312,N_22789,N_22757);
xnor U23313 (N_23313,N_22733,N_22258);
nor U23314 (N_23314,N_22586,N_22714);
and U23315 (N_23315,N_22482,N_22572);
nand U23316 (N_23316,N_22606,N_22643);
nand U23317 (N_23317,N_22621,N_22752);
or U23318 (N_23318,N_22203,N_22693);
or U23319 (N_23319,N_22333,N_22232);
or U23320 (N_23320,N_22703,N_22359);
nor U23321 (N_23321,N_22246,N_22215);
and U23322 (N_23322,N_22587,N_22380);
nand U23323 (N_23323,N_22748,N_22357);
nor U23324 (N_23324,N_22785,N_22263);
nor U23325 (N_23325,N_22663,N_22665);
xor U23326 (N_23326,N_22215,N_22521);
xor U23327 (N_23327,N_22533,N_22461);
or U23328 (N_23328,N_22725,N_22653);
and U23329 (N_23329,N_22558,N_22746);
or U23330 (N_23330,N_22727,N_22309);
nor U23331 (N_23331,N_22765,N_22614);
and U23332 (N_23332,N_22496,N_22594);
or U23333 (N_23333,N_22336,N_22345);
nand U23334 (N_23334,N_22372,N_22531);
or U23335 (N_23335,N_22482,N_22627);
and U23336 (N_23336,N_22277,N_22693);
and U23337 (N_23337,N_22279,N_22401);
and U23338 (N_23338,N_22750,N_22579);
and U23339 (N_23339,N_22727,N_22308);
xnor U23340 (N_23340,N_22628,N_22789);
xor U23341 (N_23341,N_22537,N_22586);
nor U23342 (N_23342,N_22727,N_22564);
and U23343 (N_23343,N_22767,N_22563);
xnor U23344 (N_23344,N_22451,N_22467);
and U23345 (N_23345,N_22332,N_22287);
and U23346 (N_23346,N_22633,N_22259);
and U23347 (N_23347,N_22476,N_22217);
nand U23348 (N_23348,N_22428,N_22416);
nor U23349 (N_23349,N_22220,N_22652);
nand U23350 (N_23350,N_22780,N_22210);
xnor U23351 (N_23351,N_22679,N_22634);
nor U23352 (N_23352,N_22752,N_22551);
nand U23353 (N_23353,N_22440,N_22274);
nand U23354 (N_23354,N_22525,N_22517);
or U23355 (N_23355,N_22212,N_22267);
nor U23356 (N_23356,N_22614,N_22401);
nor U23357 (N_23357,N_22306,N_22736);
nor U23358 (N_23358,N_22509,N_22247);
nor U23359 (N_23359,N_22369,N_22242);
nor U23360 (N_23360,N_22311,N_22756);
and U23361 (N_23361,N_22769,N_22492);
nor U23362 (N_23362,N_22263,N_22544);
or U23363 (N_23363,N_22394,N_22422);
nand U23364 (N_23364,N_22682,N_22296);
and U23365 (N_23365,N_22241,N_22443);
nor U23366 (N_23366,N_22415,N_22553);
and U23367 (N_23367,N_22258,N_22662);
xor U23368 (N_23368,N_22543,N_22440);
and U23369 (N_23369,N_22727,N_22415);
nor U23370 (N_23370,N_22757,N_22689);
and U23371 (N_23371,N_22458,N_22521);
nand U23372 (N_23372,N_22242,N_22317);
and U23373 (N_23373,N_22204,N_22449);
or U23374 (N_23374,N_22640,N_22603);
xnor U23375 (N_23375,N_22792,N_22409);
or U23376 (N_23376,N_22337,N_22689);
or U23377 (N_23377,N_22468,N_22610);
or U23378 (N_23378,N_22771,N_22251);
nand U23379 (N_23379,N_22525,N_22636);
nand U23380 (N_23380,N_22726,N_22611);
nand U23381 (N_23381,N_22213,N_22323);
and U23382 (N_23382,N_22264,N_22730);
nand U23383 (N_23383,N_22501,N_22699);
and U23384 (N_23384,N_22458,N_22536);
xor U23385 (N_23385,N_22452,N_22548);
and U23386 (N_23386,N_22402,N_22703);
xor U23387 (N_23387,N_22338,N_22591);
nor U23388 (N_23388,N_22312,N_22350);
or U23389 (N_23389,N_22657,N_22440);
or U23390 (N_23390,N_22661,N_22346);
nor U23391 (N_23391,N_22781,N_22307);
and U23392 (N_23392,N_22682,N_22767);
nor U23393 (N_23393,N_22491,N_22472);
xor U23394 (N_23394,N_22412,N_22609);
xnor U23395 (N_23395,N_22339,N_22697);
nor U23396 (N_23396,N_22756,N_22551);
or U23397 (N_23397,N_22297,N_22298);
nor U23398 (N_23398,N_22461,N_22528);
nor U23399 (N_23399,N_22590,N_22227);
nor U23400 (N_23400,N_22882,N_22936);
or U23401 (N_23401,N_23007,N_23096);
nand U23402 (N_23402,N_23105,N_23274);
and U23403 (N_23403,N_22841,N_23385);
or U23404 (N_23404,N_23263,N_23094);
nor U23405 (N_23405,N_22877,N_22946);
nand U23406 (N_23406,N_22939,N_23093);
nor U23407 (N_23407,N_22923,N_23081);
nor U23408 (N_23408,N_23141,N_23090);
nor U23409 (N_23409,N_23341,N_23085);
nor U23410 (N_23410,N_22926,N_22948);
or U23411 (N_23411,N_23362,N_23117);
nand U23412 (N_23412,N_22959,N_23071);
nor U23413 (N_23413,N_23387,N_23181);
xnor U23414 (N_23414,N_22966,N_23185);
nand U23415 (N_23415,N_23324,N_22894);
nor U23416 (N_23416,N_23111,N_23336);
nor U23417 (N_23417,N_22896,N_22901);
nand U23418 (N_23418,N_23133,N_23041);
nor U23419 (N_23419,N_22871,N_22891);
or U23420 (N_23420,N_23121,N_23220);
nand U23421 (N_23421,N_23310,N_23143);
and U23422 (N_23422,N_23192,N_22952);
and U23423 (N_23423,N_22943,N_23388);
nand U23424 (N_23424,N_23312,N_22953);
xnor U23425 (N_23425,N_23276,N_23011);
xor U23426 (N_23426,N_22869,N_22992);
nand U23427 (N_23427,N_23019,N_22876);
xnor U23428 (N_23428,N_23159,N_23035);
nor U23429 (N_23429,N_23024,N_23307);
nor U23430 (N_23430,N_23199,N_22805);
or U23431 (N_23431,N_23296,N_22941);
or U23432 (N_23432,N_22814,N_22934);
nand U23433 (N_23433,N_22884,N_23206);
xnor U23434 (N_23434,N_23124,N_22879);
and U23435 (N_23435,N_23172,N_23176);
nor U23436 (N_23436,N_23382,N_22824);
or U23437 (N_23437,N_22883,N_23087);
and U23438 (N_23438,N_23345,N_23318);
nand U23439 (N_23439,N_23036,N_23219);
or U23440 (N_23440,N_22956,N_22973);
and U23441 (N_23441,N_23226,N_22813);
and U23442 (N_23442,N_23045,N_22870);
or U23443 (N_23443,N_23150,N_22987);
nand U23444 (N_23444,N_23334,N_22995);
nand U23445 (N_23445,N_22802,N_23251);
or U23446 (N_23446,N_23368,N_23184);
or U23447 (N_23447,N_23142,N_23114);
and U23448 (N_23448,N_22836,N_23287);
or U23449 (N_23449,N_23367,N_22857);
nor U23450 (N_23450,N_22800,N_22861);
and U23451 (N_23451,N_22917,N_23332);
nand U23452 (N_23452,N_23380,N_23005);
or U23453 (N_23453,N_22954,N_23107);
xor U23454 (N_23454,N_22911,N_23315);
nor U23455 (N_23455,N_23089,N_23164);
nor U23456 (N_23456,N_23076,N_23179);
and U23457 (N_23457,N_23155,N_23122);
nor U23458 (N_23458,N_23297,N_22951);
nand U23459 (N_23459,N_23053,N_22895);
nor U23460 (N_23460,N_23062,N_22937);
nor U23461 (N_23461,N_23050,N_23083);
nor U23462 (N_23462,N_23228,N_23342);
and U23463 (N_23463,N_23032,N_23149);
and U23464 (N_23464,N_23357,N_23112);
or U23465 (N_23465,N_23070,N_23046);
and U23466 (N_23466,N_22831,N_23372);
nor U23467 (N_23467,N_22872,N_23059);
nand U23468 (N_23468,N_22867,N_23061);
and U23469 (N_23469,N_23271,N_23077);
or U23470 (N_23470,N_23086,N_22838);
or U23471 (N_23471,N_23370,N_22809);
and U23472 (N_23472,N_22904,N_22958);
xnor U23473 (N_23473,N_23158,N_22881);
nor U23474 (N_23474,N_23069,N_23174);
nor U23475 (N_23475,N_23288,N_23012);
nor U23476 (N_23476,N_23183,N_23091);
nand U23477 (N_23477,N_23033,N_23291);
xor U23478 (N_23478,N_23366,N_23213);
and U23479 (N_23479,N_23000,N_23075);
and U23480 (N_23480,N_22806,N_23097);
nor U23481 (N_23481,N_22807,N_23186);
and U23482 (N_23482,N_23238,N_22910);
or U23483 (N_23483,N_22962,N_23116);
xnor U23484 (N_23484,N_23225,N_23021);
nor U23485 (N_23485,N_23234,N_23146);
nand U23486 (N_23486,N_23148,N_23264);
and U23487 (N_23487,N_23386,N_22845);
or U23488 (N_23488,N_23257,N_23216);
or U23489 (N_23489,N_23048,N_23189);
and U23490 (N_23490,N_23065,N_23020);
nor U23491 (N_23491,N_23335,N_22982);
nor U23492 (N_23492,N_22835,N_22930);
nor U23493 (N_23493,N_23110,N_23308);
nor U23494 (N_23494,N_23329,N_23355);
and U23495 (N_23495,N_23381,N_23130);
or U23496 (N_23496,N_23352,N_23135);
and U23497 (N_23497,N_22975,N_23215);
nand U23498 (N_23498,N_23242,N_23131);
or U23499 (N_23499,N_23322,N_23152);
nand U23500 (N_23500,N_22988,N_22990);
or U23501 (N_23501,N_22864,N_23068);
or U23502 (N_23502,N_23350,N_22850);
nand U23503 (N_23503,N_23361,N_23072);
nand U23504 (N_23504,N_23317,N_23369);
xnor U23505 (N_23505,N_22862,N_23016);
nand U23506 (N_23506,N_23339,N_23222);
and U23507 (N_23507,N_22829,N_22826);
nand U23508 (N_23508,N_22977,N_22944);
xor U23509 (N_23509,N_23349,N_22963);
or U23510 (N_23510,N_23359,N_23134);
and U23511 (N_23511,N_23284,N_23095);
and U23512 (N_23512,N_23205,N_22905);
or U23513 (N_23513,N_22858,N_23175);
and U23514 (N_23514,N_22994,N_22912);
nor U23515 (N_23515,N_23364,N_22929);
nand U23516 (N_23516,N_23119,N_22859);
and U23517 (N_23517,N_22860,N_23260);
or U23518 (N_23518,N_23346,N_22967);
or U23519 (N_23519,N_23080,N_23254);
and U23520 (N_23520,N_22920,N_23259);
nand U23521 (N_23521,N_23229,N_22914);
nor U23522 (N_23522,N_23098,N_23203);
nand U23523 (N_23523,N_23233,N_22866);
nor U23524 (N_23524,N_23275,N_23191);
or U23525 (N_23525,N_22938,N_23003);
or U23526 (N_23526,N_23347,N_23123);
nand U23527 (N_23527,N_22964,N_23197);
nand U23528 (N_23528,N_23280,N_22898);
and U23529 (N_23529,N_23211,N_23290);
xor U23530 (N_23530,N_23207,N_22844);
nand U23531 (N_23531,N_22916,N_23398);
nor U23532 (N_23532,N_22803,N_22822);
or U23533 (N_23533,N_23006,N_23079);
nand U23534 (N_23534,N_22849,N_23025);
and U23535 (N_23535,N_23344,N_22874);
and U23536 (N_23536,N_22837,N_23137);
nor U23537 (N_23537,N_23266,N_23244);
or U23538 (N_23538,N_23161,N_22834);
nor U23539 (N_23539,N_23375,N_23316);
and U23540 (N_23540,N_23210,N_23034);
nand U23541 (N_23541,N_23343,N_23049);
or U23542 (N_23542,N_23147,N_22940);
and U23543 (N_23543,N_22945,N_22842);
nand U23544 (N_23544,N_23304,N_23017);
xor U23545 (N_23545,N_22928,N_23196);
nor U23546 (N_23546,N_23051,N_23374);
and U23547 (N_23547,N_23074,N_23294);
and U23548 (N_23548,N_23323,N_22906);
nand U23549 (N_23549,N_23232,N_22918);
and U23550 (N_23550,N_23397,N_22972);
or U23551 (N_23551,N_23391,N_22865);
nand U23552 (N_23552,N_23273,N_23394);
nor U23553 (N_23553,N_23258,N_22801);
or U23554 (N_23554,N_22919,N_22878);
and U23555 (N_23555,N_23384,N_23188);
or U23556 (N_23556,N_22932,N_23262);
nor U23557 (N_23557,N_23039,N_22961);
nor U23558 (N_23558,N_22991,N_23201);
xnor U23559 (N_23559,N_22893,N_23088);
nor U23560 (N_23560,N_23328,N_22888);
or U23561 (N_23561,N_22812,N_23333);
or U23562 (N_23562,N_22974,N_23340);
nor U23563 (N_23563,N_23099,N_23371);
or U23564 (N_23564,N_23283,N_22947);
nor U23565 (N_23565,N_22965,N_23157);
nand U23566 (N_23566,N_23057,N_23047);
nand U23567 (N_23567,N_23389,N_23305);
nand U23568 (N_23568,N_23113,N_22984);
nor U23569 (N_23569,N_22828,N_23253);
nand U23570 (N_23570,N_23127,N_23212);
nand U23571 (N_23571,N_23351,N_23010);
nand U23572 (N_23572,N_23100,N_22855);
or U23573 (N_23573,N_23331,N_22983);
or U23574 (N_23574,N_22892,N_23353);
nand U23575 (N_23575,N_23128,N_23311);
or U23576 (N_23576,N_22889,N_23092);
nand U23577 (N_23577,N_23289,N_23390);
and U23578 (N_23578,N_22942,N_23140);
and U23579 (N_23579,N_23395,N_22847);
or U23580 (N_23580,N_23145,N_22897);
or U23581 (N_23581,N_23177,N_23023);
and U23582 (N_23582,N_23103,N_23246);
and U23583 (N_23583,N_23376,N_23230);
or U23584 (N_23584,N_22804,N_22825);
and U23585 (N_23585,N_22955,N_23354);
and U23586 (N_23586,N_23139,N_23073);
xor U23587 (N_23587,N_23237,N_23378);
and U23588 (N_23588,N_23306,N_23162);
nor U23589 (N_23589,N_23292,N_23043);
xnor U23590 (N_23590,N_23365,N_22908);
xnor U23591 (N_23591,N_22854,N_23055);
and U23592 (N_23592,N_23102,N_23144);
and U23593 (N_23593,N_22880,N_23187);
and U23594 (N_23594,N_23293,N_23223);
and U23595 (N_23595,N_23221,N_22853);
nand U23596 (N_23596,N_23125,N_22873);
or U23597 (N_23597,N_22968,N_23373);
nor U23598 (N_23598,N_23214,N_23261);
and U23599 (N_23599,N_23272,N_23321);
nand U23600 (N_23600,N_23240,N_22852);
and U23601 (N_23601,N_23247,N_22821);
and U23602 (N_23602,N_23115,N_22997);
nand U23603 (N_23603,N_23363,N_23396);
and U23604 (N_23604,N_22935,N_22887);
and U23605 (N_23605,N_22971,N_23154);
xnor U23606 (N_23606,N_23030,N_22863);
and U23607 (N_23607,N_23042,N_22833);
or U23608 (N_23608,N_23004,N_23153);
or U23609 (N_23609,N_23082,N_23178);
and U23610 (N_23610,N_23279,N_23319);
and U23611 (N_23611,N_22996,N_23109);
or U23612 (N_23612,N_22999,N_23008);
nand U23613 (N_23613,N_23399,N_22950);
nor U23614 (N_23614,N_23227,N_22810);
nand U23615 (N_23615,N_23132,N_23248);
nor U23616 (N_23616,N_22993,N_23204);
and U23617 (N_23617,N_23166,N_23392);
and U23618 (N_23618,N_22915,N_22979);
nand U23619 (N_23619,N_22986,N_22981);
nor U23620 (N_23620,N_23235,N_22960);
or U23621 (N_23621,N_23326,N_23108);
and U23622 (N_23622,N_22816,N_23151);
nor U23623 (N_23623,N_23194,N_23029);
and U23624 (N_23624,N_23001,N_23193);
nand U23625 (N_23625,N_22899,N_23106);
and U23626 (N_23626,N_22856,N_23038);
and U23627 (N_23627,N_23224,N_22875);
nor U23628 (N_23628,N_23267,N_23180);
or U23629 (N_23629,N_22830,N_23066);
and U23630 (N_23630,N_23241,N_23136);
nand U23631 (N_23631,N_23327,N_23270);
nand U23632 (N_23632,N_22832,N_23052);
or U23633 (N_23633,N_22815,N_23250);
nand U23634 (N_23634,N_22868,N_23190);
nand U23635 (N_23635,N_23078,N_23298);
nand U23636 (N_23636,N_23202,N_22900);
and U23637 (N_23637,N_23383,N_23054);
nor U23638 (N_23638,N_23256,N_22924);
nor U23639 (N_23639,N_23299,N_23168);
and U23640 (N_23640,N_22818,N_22820);
nor U23641 (N_23641,N_22890,N_23026);
nand U23642 (N_23642,N_23377,N_23301);
or U23643 (N_23643,N_22903,N_23195);
and U23644 (N_23644,N_22921,N_22817);
nand U23645 (N_23645,N_23027,N_23058);
and U23646 (N_23646,N_23064,N_22931);
and U23647 (N_23647,N_22902,N_23218);
nand U23648 (N_23648,N_23356,N_23170);
or U23649 (N_23649,N_23013,N_23084);
nor U23650 (N_23650,N_23120,N_23269);
nor U23651 (N_23651,N_23163,N_23282);
xnor U23652 (N_23652,N_22927,N_23031);
nand U23653 (N_23653,N_23277,N_23015);
xor U23654 (N_23654,N_22976,N_23330);
or U23655 (N_23655,N_23138,N_22957);
nor U23656 (N_23656,N_22969,N_23243);
nand U23657 (N_23657,N_23236,N_23165);
nand U23658 (N_23658,N_23379,N_23360);
nor U23659 (N_23659,N_23002,N_23009);
nor U23660 (N_23660,N_23067,N_22819);
or U23661 (N_23661,N_23217,N_23126);
nor U23662 (N_23662,N_23265,N_23245);
nand U23663 (N_23663,N_23118,N_23056);
xor U23664 (N_23664,N_23104,N_23295);
nand U23665 (N_23665,N_23198,N_22907);
nand U23666 (N_23666,N_22885,N_23200);
and U23667 (N_23667,N_22808,N_23338);
and U23668 (N_23668,N_22949,N_23182);
and U23669 (N_23669,N_23101,N_23314);
nor U23670 (N_23670,N_22909,N_23022);
or U23671 (N_23671,N_23063,N_23040);
or U23672 (N_23672,N_23044,N_22922);
nor U23673 (N_23673,N_23300,N_22851);
nand U23674 (N_23674,N_23239,N_23156);
nor U23675 (N_23675,N_23208,N_23303);
nand U23676 (N_23676,N_23281,N_22840);
nand U23677 (N_23677,N_22886,N_23286);
nand U23678 (N_23678,N_22811,N_23209);
or U23679 (N_23679,N_22989,N_23171);
and U23680 (N_23680,N_23358,N_23014);
and U23681 (N_23681,N_22823,N_23302);
or U23682 (N_23682,N_23285,N_23231);
nor U23683 (N_23683,N_23268,N_23309);
nand U23684 (N_23684,N_23037,N_23060);
nor U23685 (N_23685,N_23129,N_23252);
and U23686 (N_23686,N_22913,N_22985);
and U23687 (N_23687,N_22998,N_23325);
nor U23688 (N_23688,N_22846,N_23337);
and U23689 (N_23689,N_22827,N_22848);
xnor U23690 (N_23690,N_23249,N_23320);
nor U23691 (N_23691,N_23169,N_23173);
or U23692 (N_23692,N_23160,N_23028);
nor U23693 (N_23693,N_22839,N_23348);
nor U23694 (N_23694,N_23167,N_23313);
nor U23695 (N_23695,N_22933,N_23393);
xor U23696 (N_23696,N_23018,N_23255);
nand U23697 (N_23697,N_22980,N_22925);
nand U23698 (N_23698,N_22978,N_22843);
nand U23699 (N_23699,N_23278,N_22970);
and U23700 (N_23700,N_23314,N_23102);
nor U23701 (N_23701,N_22845,N_23251);
and U23702 (N_23702,N_23100,N_22981);
nand U23703 (N_23703,N_23287,N_23025);
or U23704 (N_23704,N_22847,N_23277);
nor U23705 (N_23705,N_23050,N_23072);
nand U23706 (N_23706,N_22822,N_23129);
nand U23707 (N_23707,N_22838,N_23207);
nor U23708 (N_23708,N_23249,N_23377);
nor U23709 (N_23709,N_22840,N_23374);
nor U23710 (N_23710,N_22888,N_23305);
or U23711 (N_23711,N_23036,N_23193);
nor U23712 (N_23712,N_22945,N_23320);
xor U23713 (N_23713,N_23330,N_23159);
or U23714 (N_23714,N_23236,N_23185);
nand U23715 (N_23715,N_23069,N_22855);
nand U23716 (N_23716,N_22845,N_22993);
nand U23717 (N_23717,N_23384,N_23023);
nand U23718 (N_23718,N_23177,N_22852);
nor U23719 (N_23719,N_23182,N_22996);
or U23720 (N_23720,N_22904,N_23244);
nor U23721 (N_23721,N_22930,N_22958);
nor U23722 (N_23722,N_22925,N_23317);
nand U23723 (N_23723,N_23115,N_22803);
nand U23724 (N_23724,N_23001,N_23349);
nor U23725 (N_23725,N_23077,N_23156);
or U23726 (N_23726,N_23109,N_23113);
nor U23727 (N_23727,N_22988,N_22838);
nor U23728 (N_23728,N_23071,N_22939);
xor U23729 (N_23729,N_22819,N_23301);
or U23730 (N_23730,N_22905,N_22827);
nand U23731 (N_23731,N_23309,N_23337);
or U23732 (N_23732,N_23270,N_23069);
and U23733 (N_23733,N_22913,N_22933);
xor U23734 (N_23734,N_22812,N_23334);
nand U23735 (N_23735,N_23047,N_22863);
or U23736 (N_23736,N_23274,N_23157);
nor U23737 (N_23737,N_23374,N_23383);
and U23738 (N_23738,N_23011,N_22994);
or U23739 (N_23739,N_23258,N_23044);
or U23740 (N_23740,N_22800,N_22974);
nor U23741 (N_23741,N_23358,N_23013);
and U23742 (N_23742,N_23182,N_22902);
nand U23743 (N_23743,N_22838,N_23358);
or U23744 (N_23744,N_23397,N_23222);
and U23745 (N_23745,N_23133,N_23254);
nand U23746 (N_23746,N_23204,N_23050);
nor U23747 (N_23747,N_23242,N_23135);
or U23748 (N_23748,N_22821,N_23005);
nand U23749 (N_23749,N_23270,N_23193);
nor U23750 (N_23750,N_22969,N_23200);
and U23751 (N_23751,N_23358,N_23287);
nand U23752 (N_23752,N_23049,N_23260);
or U23753 (N_23753,N_23309,N_22937);
nand U23754 (N_23754,N_23205,N_23320);
or U23755 (N_23755,N_22874,N_23299);
or U23756 (N_23756,N_22994,N_22973);
or U23757 (N_23757,N_22884,N_23138);
nor U23758 (N_23758,N_23231,N_22869);
xor U23759 (N_23759,N_23289,N_22933);
nand U23760 (N_23760,N_23253,N_23291);
nor U23761 (N_23761,N_22815,N_23177);
nand U23762 (N_23762,N_22917,N_23211);
nor U23763 (N_23763,N_23085,N_23041);
and U23764 (N_23764,N_22958,N_23020);
nor U23765 (N_23765,N_23111,N_23235);
nand U23766 (N_23766,N_23041,N_23390);
nand U23767 (N_23767,N_23184,N_23099);
or U23768 (N_23768,N_23011,N_23026);
and U23769 (N_23769,N_22951,N_23141);
nand U23770 (N_23770,N_23044,N_23021);
xor U23771 (N_23771,N_23397,N_23220);
or U23772 (N_23772,N_23152,N_22907);
xnor U23773 (N_23773,N_22964,N_23053);
or U23774 (N_23774,N_22860,N_23345);
nor U23775 (N_23775,N_22940,N_22942);
or U23776 (N_23776,N_22896,N_23306);
nor U23777 (N_23777,N_23266,N_23209);
nand U23778 (N_23778,N_23256,N_23340);
nand U23779 (N_23779,N_23334,N_23093);
or U23780 (N_23780,N_22951,N_22924);
xor U23781 (N_23781,N_23333,N_22908);
xnor U23782 (N_23782,N_23201,N_22936);
nor U23783 (N_23783,N_23142,N_23239);
xor U23784 (N_23784,N_23353,N_22968);
nand U23785 (N_23785,N_23153,N_23241);
and U23786 (N_23786,N_22817,N_23190);
xor U23787 (N_23787,N_22997,N_22894);
or U23788 (N_23788,N_22877,N_22827);
and U23789 (N_23789,N_22851,N_22979);
and U23790 (N_23790,N_23107,N_22857);
nor U23791 (N_23791,N_23337,N_23174);
or U23792 (N_23792,N_23264,N_22825);
nor U23793 (N_23793,N_22883,N_23205);
and U23794 (N_23794,N_23389,N_23135);
nand U23795 (N_23795,N_23220,N_23350);
nand U23796 (N_23796,N_23218,N_22914);
nand U23797 (N_23797,N_22968,N_22867);
or U23798 (N_23798,N_22807,N_23294);
nor U23799 (N_23799,N_23182,N_22927);
or U23800 (N_23800,N_23355,N_22833);
xor U23801 (N_23801,N_22809,N_22956);
nor U23802 (N_23802,N_22868,N_23287);
or U23803 (N_23803,N_22827,N_23026);
nand U23804 (N_23804,N_23095,N_23187);
or U23805 (N_23805,N_22843,N_23273);
nand U23806 (N_23806,N_22840,N_23145);
xor U23807 (N_23807,N_23188,N_22981);
or U23808 (N_23808,N_22923,N_22838);
or U23809 (N_23809,N_23063,N_23103);
or U23810 (N_23810,N_23028,N_23378);
or U23811 (N_23811,N_22919,N_23265);
nor U23812 (N_23812,N_23197,N_23270);
xor U23813 (N_23813,N_22876,N_22945);
nor U23814 (N_23814,N_22881,N_23027);
and U23815 (N_23815,N_22834,N_23031);
nand U23816 (N_23816,N_22871,N_23363);
or U23817 (N_23817,N_23048,N_23000);
nor U23818 (N_23818,N_23214,N_23118);
or U23819 (N_23819,N_23010,N_23331);
nor U23820 (N_23820,N_23388,N_22814);
xor U23821 (N_23821,N_23299,N_23352);
nand U23822 (N_23822,N_23386,N_23088);
nand U23823 (N_23823,N_22864,N_23304);
xnor U23824 (N_23824,N_23276,N_23146);
or U23825 (N_23825,N_22903,N_22833);
nor U23826 (N_23826,N_23264,N_22811);
xor U23827 (N_23827,N_23101,N_23373);
xor U23828 (N_23828,N_22828,N_23075);
nor U23829 (N_23829,N_22875,N_23108);
nand U23830 (N_23830,N_23314,N_22934);
nor U23831 (N_23831,N_23297,N_23143);
xor U23832 (N_23832,N_23204,N_22945);
nand U23833 (N_23833,N_22850,N_23196);
nand U23834 (N_23834,N_23354,N_23197);
xnor U23835 (N_23835,N_22920,N_23052);
nor U23836 (N_23836,N_22867,N_23252);
or U23837 (N_23837,N_23120,N_23367);
or U23838 (N_23838,N_23073,N_23303);
and U23839 (N_23839,N_23335,N_23132);
nand U23840 (N_23840,N_22912,N_23265);
and U23841 (N_23841,N_23192,N_22820);
xor U23842 (N_23842,N_22998,N_22854);
or U23843 (N_23843,N_23352,N_23080);
and U23844 (N_23844,N_22897,N_23347);
xor U23845 (N_23845,N_22951,N_22890);
xnor U23846 (N_23846,N_23064,N_22955);
or U23847 (N_23847,N_23210,N_22890);
nand U23848 (N_23848,N_23246,N_23232);
and U23849 (N_23849,N_23279,N_23313);
or U23850 (N_23850,N_23336,N_22961);
and U23851 (N_23851,N_23104,N_23058);
and U23852 (N_23852,N_22984,N_23348);
nand U23853 (N_23853,N_22857,N_23391);
xnor U23854 (N_23854,N_23385,N_23391);
or U23855 (N_23855,N_23113,N_23174);
and U23856 (N_23856,N_23131,N_23284);
and U23857 (N_23857,N_22920,N_22838);
nand U23858 (N_23858,N_23071,N_22940);
xor U23859 (N_23859,N_23204,N_22941);
xor U23860 (N_23860,N_23060,N_23227);
and U23861 (N_23861,N_23107,N_22885);
or U23862 (N_23862,N_22920,N_22846);
nor U23863 (N_23863,N_23362,N_23064);
nand U23864 (N_23864,N_22911,N_22878);
or U23865 (N_23865,N_23266,N_22867);
nor U23866 (N_23866,N_23135,N_23114);
and U23867 (N_23867,N_22898,N_23091);
nor U23868 (N_23868,N_22819,N_22961);
nor U23869 (N_23869,N_23181,N_23131);
and U23870 (N_23870,N_23397,N_23346);
nor U23871 (N_23871,N_23141,N_23084);
nor U23872 (N_23872,N_22853,N_23146);
nand U23873 (N_23873,N_22897,N_23124);
xor U23874 (N_23874,N_23097,N_23207);
nor U23875 (N_23875,N_22819,N_23175);
xor U23876 (N_23876,N_23316,N_23119);
nand U23877 (N_23877,N_22904,N_22815);
nand U23878 (N_23878,N_23209,N_23172);
or U23879 (N_23879,N_22918,N_23285);
nand U23880 (N_23880,N_22926,N_23292);
and U23881 (N_23881,N_22999,N_22967);
nand U23882 (N_23882,N_22984,N_23044);
nor U23883 (N_23883,N_23015,N_23171);
or U23884 (N_23884,N_22967,N_23382);
nand U23885 (N_23885,N_23170,N_22865);
nand U23886 (N_23886,N_22990,N_22983);
nor U23887 (N_23887,N_22831,N_23262);
and U23888 (N_23888,N_23067,N_22948);
nand U23889 (N_23889,N_23328,N_23062);
and U23890 (N_23890,N_23206,N_22952);
nor U23891 (N_23891,N_22973,N_23229);
nor U23892 (N_23892,N_23190,N_23031);
nand U23893 (N_23893,N_23149,N_23146);
nand U23894 (N_23894,N_23132,N_23370);
or U23895 (N_23895,N_22922,N_22935);
xnor U23896 (N_23896,N_23183,N_23173);
xor U23897 (N_23897,N_23260,N_23057);
and U23898 (N_23898,N_23162,N_22937);
nor U23899 (N_23899,N_22928,N_22918);
nor U23900 (N_23900,N_23056,N_23126);
or U23901 (N_23901,N_23042,N_23201);
xnor U23902 (N_23902,N_23314,N_23203);
nand U23903 (N_23903,N_23354,N_22855);
nand U23904 (N_23904,N_23333,N_23116);
nand U23905 (N_23905,N_23146,N_23331);
and U23906 (N_23906,N_23373,N_23035);
and U23907 (N_23907,N_22931,N_23275);
nor U23908 (N_23908,N_22994,N_22935);
and U23909 (N_23909,N_23094,N_23104);
and U23910 (N_23910,N_23246,N_22997);
xor U23911 (N_23911,N_22960,N_23378);
xnor U23912 (N_23912,N_23286,N_22947);
nor U23913 (N_23913,N_22999,N_22907);
or U23914 (N_23914,N_22879,N_23217);
and U23915 (N_23915,N_23276,N_23382);
nor U23916 (N_23916,N_23148,N_23201);
or U23917 (N_23917,N_23113,N_22979);
nor U23918 (N_23918,N_23027,N_23006);
nand U23919 (N_23919,N_22870,N_23254);
nand U23920 (N_23920,N_23247,N_22924);
xor U23921 (N_23921,N_22959,N_23138);
xor U23922 (N_23922,N_22838,N_23007);
nor U23923 (N_23923,N_23060,N_23298);
and U23924 (N_23924,N_23035,N_23093);
nor U23925 (N_23925,N_23134,N_23004);
nand U23926 (N_23926,N_23034,N_23266);
xnor U23927 (N_23927,N_23023,N_22826);
nand U23928 (N_23928,N_23039,N_22897);
xnor U23929 (N_23929,N_23399,N_22921);
and U23930 (N_23930,N_22935,N_22872);
xnor U23931 (N_23931,N_22825,N_23008);
or U23932 (N_23932,N_22918,N_22960);
nand U23933 (N_23933,N_22822,N_22960);
or U23934 (N_23934,N_22865,N_22941);
nand U23935 (N_23935,N_22926,N_22904);
nor U23936 (N_23936,N_23008,N_23046);
xor U23937 (N_23937,N_23071,N_23078);
nand U23938 (N_23938,N_23208,N_23225);
xor U23939 (N_23939,N_23207,N_22925);
nor U23940 (N_23940,N_23340,N_22846);
nand U23941 (N_23941,N_23167,N_23310);
nand U23942 (N_23942,N_22873,N_22966);
and U23943 (N_23943,N_23097,N_22862);
xor U23944 (N_23944,N_23391,N_23133);
or U23945 (N_23945,N_23232,N_23163);
nor U23946 (N_23946,N_22909,N_23252);
and U23947 (N_23947,N_22872,N_23248);
and U23948 (N_23948,N_23252,N_23391);
nand U23949 (N_23949,N_22831,N_23008);
nand U23950 (N_23950,N_22937,N_23305);
nand U23951 (N_23951,N_22902,N_23360);
xnor U23952 (N_23952,N_23266,N_22851);
or U23953 (N_23953,N_23328,N_23065);
or U23954 (N_23954,N_23212,N_23204);
nand U23955 (N_23955,N_23217,N_23083);
xnor U23956 (N_23956,N_23033,N_23039);
and U23957 (N_23957,N_23244,N_23167);
or U23958 (N_23958,N_22877,N_22843);
nor U23959 (N_23959,N_23001,N_22975);
or U23960 (N_23960,N_23022,N_22848);
nor U23961 (N_23961,N_23109,N_23215);
or U23962 (N_23962,N_23101,N_23242);
or U23963 (N_23963,N_23323,N_23263);
nand U23964 (N_23964,N_23318,N_23038);
nor U23965 (N_23965,N_23124,N_23099);
and U23966 (N_23966,N_23387,N_23192);
xnor U23967 (N_23967,N_23302,N_22877);
xnor U23968 (N_23968,N_22993,N_22864);
and U23969 (N_23969,N_23227,N_23392);
and U23970 (N_23970,N_23132,N_23356);
nand U23971 (N_23971,N_22948,N_23310);
nand U23972 (N_23972,N_23237,N_23038);
xnor U23973 (N_23973,N_23377,N_23172);
nand U23974 (N_23974,N_23328,N_23245);
or U23975 (N_23975,N_23265,N_23389);
and U23976 (N_23976,N_22905,N_23324);
or U23977 (N_23977,N_22983,N_23241);
and U23978 (N_23978,N_23268,N_22852);
nor U23979 (N_23979,N_23379,N_22867);
or U23980 (N_23980,N_23322,N_22860);
or U23981 (N_23981,N_22805,N_22978);
and U23982 (N_23982,N_23069,N_23191);
nor U23983 (N_23983,N_22879,N_23305);
or U23984 (N_23984,N_23149,N_22901);
nand U23985 (N_23985,N_23349,N_23108);
and U23986 (N_23986,N_23197,N_23310);
nand U23987 (N_23987,N_23087,N_23192);
and U23988 (N_23988,N_22970,N_23023);
or U23989 (N_23989,N_23064,N_23036);
nor U23990 (N_23990,N_23368,N_23307);
nor U23991 (N_23991,N_23115,N_23399);
and U23992 (N_23992,N_22910,N_23121);
and U23993 (N_23993,N_23272,N_22967);
and U23994 (N_23994,N_23018,N_22826);
xor U23995 (N_23995,N_22912,N_23317);
and U23996 (N_23996,N_23384,N_23002);
nor U23997 (N_23997,N_23058,N_23311);
nand U23998 (N_23998,N_22884,N_23020);
nor U23999 (N_23999,N_23358,N_23183);
nand U24000 (N_24000,N_23751,N_23816);
nand U24001 (N_24001,N_23828,N_23552);
nor U24002 (N_24002,N_23892,N_23404);
and U24003 (N_24003,N_23633,N_23506);
xnor U24004 (N_24004,N_23851,N_23693);
nand U24005 (N_24005,N_23403,N_23960);
and U24006 (N_24006,N_23544,N_23972);
or U24007 (N_24007,N_23997,N_23658);
xnor U24008 (N_24008,N_23792,N_23976);
nand U24009 (N_24009,N_23598,N_23743);
or U24010 (N_24010,N_23984,N_23660);
or U24011 (N_24011,N_23454,N_23741);
or U24012 (N_24012,N_23737,N_23464);
xnor U24013 (N_24013,N_23535,N_23745);
nand U24014 (N_24014,N_23837,N_23589);
xnor U24015 (N_24015,N_23523,N_23424);
nand U24016 (N_24016,N_23441,N_23877);
nor U24017 (N_24017,N_23527,N_23492);
nand U24018 (N_24018,N_23964,N_23482);
nand U24019 (N_24019,N_23754,N_23744);
nand U24020 (N_24020,N_23966,N_23635);
xor U24021 (N_24021,N_23847,N_23762);
and U24022 (N_24022,N_23409,N_23873);
or U24023 (N_24023,N_23659,N_23592);
or U24024 (N_24024,N_23508,N_23583);
or U24025 (N_24025,N_23996,N_23759);
and U24026 (N_24026,N_23553,N_23462);
nor U24027 (N_24027,N_23685,N_23600);
xor U24028 (N_24028,N_23823,N_23785);
nor U24029 (N_24029,N_23747,N_23879);
or U24030 (N_24030,N_23712,N_23477);
or U24031 (N_24031,N_23532,N_23418);
or U24032 (N_24032,N_23510,N_23574);
nand U24033 (N_24033,N_23728,N_23449);
nor U24034 (N_24034,N_23905,N_23849);
and U24035 (N_24035,N_23834,N_23983);
nor U24036 (N_24036,N_23804,N_23585);
nand U24037 (N_24037,N_23439,N_23611);
nor U24038 (N_24038,N_23886,N_23698);
nand U24039 (N_24039,N_23739,N_23519);
nand U24040 (N_24040,N_23433,N_23749);
or U24041 (N_24041,N_23881,N_23594);
or U24042 (N_24042,N_23723,N_23421);
nor U24043 (N_24043,N_23802,N_23461);
nand U24044 (N_24044,N_23995,N_23599);
or U24045 (N_24045,N_23734,N_23683);
nand U24046 (N_24046,N_23790,N_23573);
or U24047 (N_24047,N_23590,N_23758);
or U24048 (N_24048,N_23929,N_23530);
or U24049 (N_24049,N_23575,N_23624);
and U24050 (N_24050,N_23752,N_23703);
nand U24051 (N_24051,N_23761,N_23609);
nand U24052 (N_24052,N_23870,N_23806);
and U24053 (N_24053,N_23755,N_23437);
or U24054 (N_24054,N_23911,N_23496);
nand U24055 (N_24055,N_23676,N_23612);
nand U24056 (N_24056,N_23490,N_23940);
nor U24057 (N_24057,N_23444,N_23643);
or U24058 (N_24058,N_23625,N_23824);
and U24059 (N_24059,N_23414,N_23571);
and U24060 (N_24060,N_23738,N_23945);
nand U24061 (N_24061,N_23668,N_23783);
and U24062 (N_24062,N_23467,N_23674);
and U24063 (N_24063,N_23710,N_23460);
and U24064 (N_24064,N_23662,N_23914);
and U24065 (N_24065,N_23500,N_23998);
nor U24066 (N_24066,N_23434,N_23430);
nor U24067 (N_24067,N_23807,N_23503);
and U24068 (N_24068,N_23864,N_23717);
or U24069 (N_24069,N_23623,N_23488);
nor U24070 (N_24070,N_23420,N_23858);
and U24071 (N_24071,N_23440,N_23551);
nand U24072 (N_24072,N_23910,N_23988);
xor U24073 (N_24073,N_23595,N_23796);
nor U24074 (N_24074,N_23493,N_23567);
nand U24075 (N_24075,N_23400,N_23821);
and U24076 (N_24076,N_23419,N_23713);
and U24077 (N_24077,N_23686,N_23608);
or U24078 (N_24078,N_23657,N_23813);
nand U24079 (N_24079,N_23669,N_23426);
xnor U24080 (N_24080,N_23512,N_23974);
xnor U24081 (N_24081,N_23913,N_23915);
and U24082 (N_24082,N_23774,N_23570);
nand U24083 (N_24083,N_23541,N_23616);
nor U24084 (N_24084,N_23401,N_23885);
xnor U24085 (N_24085,N_23748,N_23920);
and U24086 (N_24086,N_23750,N_23619);
xor U24087 (N_24087,N_23793,N_23861);
or U24088 (N_24088,N_23696,N_23466);
nor U24089 (N_24089,N_23952,N_23602);
or U24090 (N_24090,N_23800,N_23591);
nor U24091 (N_24091,N_23631,N_23706);
nand U24092 (N_24092,N_23465,N_23990);
nand U24093 (N_24093,N_23639,N_23724);
nand U24094 (N_24094,N_23642,N_23561);
nand U24095 (N_24095,N_23498,N_23636);
or U24096 (N_24096,N_23582,N_23961);
or U24097 (N_24097,N_23903,N_23880);
and U24098 (N_24098,N_23967,N_23630);
nor U24099 (N_24099,N_23581,N_23540);
nand U24100 (N_24100,N_23432,N_23515);
and U24101 (N_24101,N_23661,N_23822);
or U24102 (N_24102,N_23843,N_23832);
and U24103 (N_24103,N_23842,N_23451);
nand U24104 (N_24104,N_23875,N_23850);
or U24105 (N_24105,N_23692,N_23664);
nand U24106 (N_24106,N_23939,N_23415);
nand U24107 (N_24107,N_23691,N_23704);
or U24108 (N_24108,N_23714,N_23931);
nor U24109 (N_24109,N_23766,N_23829);
and U24110 (N_24110,N_23924,N_23884);
nor U24111 (N_24111,N_23546,N_23999);
nor U24112 (N_24112,N_23618,N_23406);
or U24113 (N_24113,N_23564,N_23840);
nor U24114 (N_24114,N_23771,N_23562);
nand U24115 (N_24115,N_23978,N_23930);
or U24116 (N_24116,N_23673,N_23912);
or U24117 (N_24117,N_23678,N_23448);
nand U24118 (N_24118,N_23483,N_23620);
nor U24119 (N_24119,N_23601,N_23906);
nor U24120 (N_24120,N_23878,N_23932);
and U24121 (N_24121,N_23969,N_23736);
nand U24122 (N_24122,N_23679,N_23809);
nor U24123 (N_24123,N_23525,N_23962);
nor U24124 (N_24124,N_23777,N_23632);
nand U24125 (N_24125,N_23947,N_23982);
and U24126 (N_24126,N_23726,N_23648);
or U24127 (N_24127,N_23533,N_23442);
or U24128 (N_24128,N_23672,N_23764);
or U24129 (N_24129,N_23702,N_23455);
nor U24130 (N_24130,N_23933,N_23993);
and U24131 (N_24131,N_23528,N_23645);
or U24132 (N_24132,N_23588,N_23946);
or U24133 (N_24133,N_23471,N_23563);
nand U24134 (N_24134,N_23656,N_23789);
and U24135 (N_24135,N_23919,N_23787);
or U24136 (N_24136,N_23480,N_23487);
xor U24137 (N_24137,N_23705,N_23470);
or U24138 (N_24138,N_23943,N_23841);
nor U24139 (N_24139,N_23408,N_23959);
or U24140 (N_24140,N_23894,N_23887);
or U24141 (N_24141,N_23497,N_23604);
xor U24142 (N_24142,N_23901,N_23992);
or U24143 (N_24143,N_23667,N_23935);
nor U24144 (N_24144,N_23463,N_23446);
or U24145 (N_24145,N_23778,N_23922);
and U24146 (N_24146,N_23942,N_23413);
and U24147 (N_24147,N_23457,N_23797);
or U24148 (N_24148,N_23486,N_23957);
or U24149 (N_24149,N_23476,N_23916);
and U24150 (N_24150,N_23665,N_23890);
nor U24151 (N_24151,N_23504,N_23513);
nand U24152 (N_24152,N_23534,N_23980);
xnor U24153 (N_24153,N_23836,N_23615);
and U24154 (N_24154,N_23977,N_23740);
and U24155 (N_24155,N_23495,N_23555);
and U24156 (N_24156,N_23556,N_23794);
xnor U24157 (N_24157,N_23819,N_23926);
nor U24158 (N_24158,N_23720,N_23474);
or U24159 (N_24159,N_23469,N_23863);
and U24160 (N_24160,N_23955,N_23989);
or U24161 (N_24161,N_23803,N_23820);
nand U24162 (N_24162,N_23481,N_23459);
nand U24163 (N_24163,N_23954,N_23407);
nor U24164 (N_24164,N_23908,N_23893);
nand U24165 (N_24165,N_23427,N_23904);
or U24166 (N_24166,N_23772,N_23429);
xor U24167 (N_24167,N_23514,N_23860);
xnor U24168 (N_24168,N_23944,N_23422);
nand U24169 (N_24169,N_23622,N_23666);
nand U24170 (N_24170,N_23991,N_23447);
or U24171 (N_24171,N_23979,N_23502);
and U24172 (N_24172,N_23688,N_23613);
nand U24173 (N_24173,N_23681,N_23950);
nand U24174 (N_24174,N_23545,N_23918);
and U24175 (N_24175,N_23499,N_23557);
nor U24176 (N_24176,N_23788,N_23452);
and U24177 (N_24177,N_23485,N_23647);
or U24178 (N_24178,N_23605,N_23652);
and U24179 (N_24179,N_23644,N_23610);
nand U24180 (N_24180,N_23938,N_23867);
and U24181 (N_24181,N_23517,N_23554);
nand U24182 (N_24182,N_23453,N_23852);
or U24183 (N_24183,N_23770,N_23786);
nand U24184 (N_24184,N_23970,N_23687);
and U24185 (N_24185,N_23951,N_23649);
nand U24186 (N_24186,N_23833,N_23853);
nand U24187 (N_24187,N_23765,N_23577);
nand U24188 (N_24188,N_23509,N_23732);
nor U24189 (N_24189,N_23529,N_23963);
or U24190 (N_24190,N_23902,N_23937);
xor U24191 (N_24191,N_23646,N_23614);
nand U24192 (N_24192,N_23768,N_23539);
and U24193 (N_24193,N_23671,N_23568);
and U24194 (N_24194,N_23869,N_23458);
or U24195 (N_24195,N_23580,N_23578);
nor U24196 (N_24196,N_23559,N_23923);
xor U24197 (N_24197,N_23838,N_23675);
or U24198 (N_24198,N_23773,N_23735);
xor U24199 (N_24199,N_23928,N_23891);
nand U24200 (N_24200,N_23505,N_23965);
nor U24201 (N_24201,N_23727,N_23538);
nand U24202 (N_24202,N_23986,N_23412);
and U24203 (N_24203,N_23862,N_23569);
or U24204 (N_24204,N_23700,N_23697);
nor U24205 (N_24205,N_23572,N_23898);
nand U24206 (N_24206,N_23814,N_23815);
nor U24207 (N_24207,N_23634,N_23468);
nor U24208 (N_24208,N_23699,N_23973);
or U24209 (N_24209,N_23994,N_23417);
and U24210 (N_24210,N_23524,N_23817);
nor U24211 (N_24211,N_23907,N_23956);
or U24212 (N_24212,N_23731,N_23876);
and U24213 (N_24213,N_23981,N_23895);
nor U24214 (N_24214,N_23767,N_23596);
xor U24215 (N_24215,N_23684,N_23948);
and U24216 (N_24216,N_23402,N_23711);
nand U24217 (N_24217,N_23936,N_23899);
or U24218 (N_24218,N_23690,N_23709);
nand U24219 (N_24219,N_23542,N_23521);
and U24220 (N_24220,N_23775,N_23653);
and U24221 (N_24221,N_23694,N_23549);
nand U24222 (N_24222,N_23576,N_23810);
xnor U24223 (N_24223,N_23416,N_23801);
nor U24224 (N_24224,N_23719,N_23827);
or U24225 (N_24225,N_23606,N_23655);
nand U24226 (N_24226,N_23680,N_23730);
nand U24227 (N_24227,N_23949,N_23494);
and U24228 (N_24228,N_23479,N_23971);
xor U24229 (N_24229,N_23707,N_23757);
xor U24230 (N_24230,N_23511,N_23799);
or U24231 (N_24231,N_23587,N_23987);
nor U24232 (N_24232,N_23866,N_23882);
xnor U24233 (N_24233,N_23701,N_23543);
nand U24234 (N_24234,N_23968,N_23909);
nand U24235 (N_24235,N_23782,N_23626);
and U24236 (N_24236,N_23868,N_23900);
nand U24237 (N_24237,N_23586,N_23769);
nor U24238 (N_24238,N_23760,N_23566);
nor U24239 (N_24239,N_23670,N_23725);
or U24240 (N_24240,N_23795,N_23507);
nor U24241 (N_24241,N_23818,N_23518);
nand U24242 (N_24242,N_23742,N_23560);
nand U24243 (N_24243,N_23548,N_23830);
nor U24244 (N_24244,N_23791,N_23531);
nor U24245 (N_24245,N_23445,N_23663);
or U24246 (N_24246,N_23854,N_23689);
or U24247 (N_24247,N_23856,N_23537);
nand U24248 (N_24248,N_23859,N_23784);
nand U24249 (N_24249,N_23925,N_23756);
nand U24250 (N_24250,N_23410,N_23934);
xor U24251 (N_24251,N_23826,N_23593);
or U24252 (N_24252,N_23522,N_23550);
nor U24253 (N_24253,N_23845,N_23516);
xnor U24254 (N_24254,N_23654,N_23855);
nor U24255 (N_24255,N_23921,N_23889);
and U24256 (N_24256,N_23597,N_23637);
nor U24257 (N_24257,N_23491,N_23733);
nor U24258 (N_24258,N_23489,N_23721);
nor U24259 (N_24259,N_23953,N_23780);
and U24260 (N_24260,N_23846,N_23848);
nand U24261 (N_24261,N_23917,N_23718);
nor U24262 (N_24262,N_23781,N_23865);
nand U24263 (N_24263,N_23547,N_23708);
nand U24264 (N_24264,N_23638,N_23779);
xnor U24265 (N_24265,N_23425,N_23475);
nor U24266 (N_24266,N_23844,N_23520);
nand U24267 (N_24267,N_23411,N_23438);
nor U24268 (N_24268,N_23565,N_23558);
or U24269 (N_24269,N_23677,N_23473);
nor U24270 (N_24270,N_23857,N_23888);
nand U24271 (N_24271,N_23798,N_23872);
nand U24272 (N_24272,N_23484,N_23436);
xor U24273 (N_24273,N_23456,N_23423);
nand U24274 (N_24274,N_23941,N_23958);
nand U24275 (N_24275,N_23975,N_23682);
or U24276 (N_24276,N_23450,N_23428);
and U24277 (N_24277,N_23627,N_23443);
nand U24278 (N_24278,N_23603,N_23835);
nand U24279 (N_24279,N_23722,N_23501);
or U24280 (N_24280,N_23716,N_23825);
or U24281 (N_24281,N_23812,N_23871);
nor U24282 (N_24282,N_23628,N_23715);
or U24283 (N_24283,N_23874,N_23831);
and U24284 (N_24284,N_23763,N_23478);
nand U24285 (N_24285,N_23695,N_23985);
and U24286 (N_24286,N_23526,N_23776);
and U24287 (N_24287,N_23927,N_23650);
nor U24288 (N_24288,N_23897,N_23472);
and U24289 (N_24289,N_23536,N_23805);
or U24290 (N_24290,N_23640,N_23629);
or U24291 (N_24291,N_23811,N_23641);
nand U24292 (N_24292,N_23431,N_23651);
or U24293 (N_24293,N_23883,N_23753);
nor U24294 (N_24294,N_23896,N_23621);
xor U24295 (N_24295,N_23746,N_23808);
nor U24296 (N_24296,N_23729,N_23579);
nor U24297 (N_24297,N_23839,N_23405);
and U24298 (N_24298,N_23607,N_23584);
nand U24299 (N_24299,N_23617,N_23435);
nand U24300 (N_24300,N_23540,N_23898);
or U24301 (N_24301,N_23610,N_23607);
xor U24302 (N_24302,N_23606,N_23860);
and U24303 (N_24303,N_23988,N_23448);
nand U24304 (N_24304,N_23658,N_23513);
xnor U24305 (N_24305,N_23722,N_23743);
or U24306 (N_24306,N_23463,N_23424);
and U24307 (N_24307,N_23911,N_23553);
or U24308 (N_24308,N_23853,N_23531);
nand U24309 (N_24309,N_23841,N_23488);
or U24310 (N_24310,N_23473,N_23657);
and U24311 (N_24311,N_23885,N_23752);
or U24312 (N_24312,N_23524,N_23897);
xor U24313 (N_24313,N_23577,N_23405);
and U24314 (N_24314,N_23505,N_23404);
and U24315 (N_24315,N_23945,N_23936);
and U24316 (N_24316,N_23975,N_23884);
nand U24317 (N_24317,N_23535,N_23881);
and U24318 (N_24318,N_23779,N_23423);
and U24319 (N_24319,N_23951,N_23928);
and U24320 (N_24320,N_23834,N_23825);
nand U24321 (N_24321,N_23939,N_23696);
nand U24322 (N_24322,N_23937,N_23893);
or U24323 (N_24323,N_23863,N_23848);
or U24324 (N_24324,N_23752,N_23974);
nor U24325 (N_24325,N_23408,N_23956);
nor U24326 (N_24326,N_23563,N_23596);
nand U24327 (N_24327,N_23477,N_23776);
nand U24328 (N_24328,N_23507,N_23731);
and U24329 (N_24329,N_23736,N_23436);
nor U24330 (N_24330,N_23466,N_23718);
nor U24331 (N_24331,N_23595,N_23846);
xnor U24332 (N_24332,N_23748,N_23840);
and U24333 (N_24333,N_23676,N_23908);
nor U24334 (N_24334,N_23941,N_23610);
nand U24335 (N_24335,N_23626,N_23677);
nand U24336 (N_24336,N_23611,N_23554);
nor U24337 (N_24337,N_23785,N_23666);
and U24338 (N_24338,N_23575,N_23849);
or U24339 (N_24339,N_23826,N_23712);
and U24340 (N_24340,N_23621,N_23805);
and U24341 (N_24341,N_23573,N_23825);
nand U24342 (N_24342,N_23944,N_23708);
nor U24343 (N_24343,N_23507,N_23852);
or U24344 (N_24344,N_23954,N_23791);
nand U24345 (N_24345,N_23953,N_23892);
or U24346 (N_24346,N_23986,N_23839);
nor U24347 (N_24347,N_23623,N_23925);
nor U24348 (N_24348,N_23456,N_23652);
and U24349 (N_24349,N_23688,N_23905);
nor U24350 (N_24350,N_23454,N_23907);
or U24351 (N_24351,N_23693,N_23413);
nor U24352 (N_24352,N_23935,N_23468);
or U24353 (N_24353,N_23814,N_23433);
and U24354 (N_24354,N_23669,N_23935);
nand U24355 (N_24355,N_23618,N_23757);
nand U24356 (N_24356,N_23861,N_23757);
nor U24357 (N_24357,N_23511,N_23951);
nor U24358 (N_24358,N_23710,N_23762);
or U24359 (N_24359,N_23804,N_23857);
nand U24360 (N_24360,N_23918,N_23843);
nand U24361 (N_24361,N_23954,N_23803);
or U24362 (N_24362,N_23895,N_23912);
and U24363 (N_24363,N_23787,N_23690);
and U24364 (N_24364,N_23663,N_23521);
or U24365 (N_24365,N_23680,N_23435);
or U24366 (N_24366,N_23896,N_23963);
or U24367 (N_24367,N_23809,N_23741);
xnor U24368 (N_24368,N_23471,N_23693);
nor U24369 (N_24369,N_23552,N_23700);
xor U24370 (N_24370,N_23687,N_23628);
nand U24371 (N_24371,N_23839,N_23894);
nor U24372 (N_24372,N_23862,N_23516);
and U24373 (N_24373,N_23748,N_23719);
nor U24374 (N_24374,N_23652,N_23956);
nand U24375 (N_24375,N_23521,N_23585);
xnor U24376 (N_24376,N_23958,N_23765);
xor U24377 (N_24377,N_23692,N_23983);
nand U24378 (N_24378,N_23825,N_23654);
and U24379 (N_24379,N_23787,N_23959);
or U24380 (N_24380,N_23751,N_23447);
nor U24381 (N_24381,N_23657,N_23665);
nor U24382 (N_24382,N_23814,N_23843);
and U24383 (N_24383,N_23919,N_23784);
nor U24384 (N_24384,N_23629,N_23487);
or U24385 (N_24385,N_23700,N_23400);
and U24386 (N_24386,N_23485,N_23624);
nand U24387 (N_24387,N_23905,N_23428);
nand U24388 (N_24388,N_23507,N_23862);
nand U24389 (N_24389,N_23975,N_23962);
nand U24390 (N_24390,N_23543,N_23742);
nand U24391 (N_24391,N_23596,N_23715);
nand U24392 (N_24392,N_23720,N_23949);
and U24393 (N_24393,N_23661,N_23461);
nor U24394 (N_24394,N_23624,N_23459);
nand U24395 (N_24395,N_23515,N_23743);
or U24396 (N_24396,N_23713,N_23639);
and U24397 (N_24397,N_23457,N_23406);
nand U24398 (N_24398,N_23753,N_23896);
or U24399 (N_24399,N_23520,N_23940);
and U24400 (N_24400,N_23530,N_23705);
or U24401 (N_24401,N_23495,N_23656);
or U24402 (N_24402,N_23777,N_23925);
and U24403 (N_24403,N_23877,N_23484);
or U24404 (N_24404,N_23950,N_23943);
and U24405 (N_24405,N_23682,N_23712);
and U24406 (N_24406,N_23563,N_23758);
or U24407 (N_24407,N_23792,N_23901);
xor U24408 (N_24408,N_23446,N_23788);
nand U24409 (N_24409,N_23729,N_23508);
nand U24410 (N_24410,N_23562,N_23602);
or U24411 (N_24411,N_23751,N_23426);
nor U24412 (N_24412,N_23864,N_23522);
nand U24413 (N_24413,N_23541,N_23860);
xnor U24414 (N_24414,N_23672,N_23640);
nand U24415 (N_24415,N_23702,N_23534);
nor U24416 (N_24416,N_23959,N_23475);
nand U24417 (N_24417,N_23674,N_23729);
nor U24418 (N_24418,N_23726,N_23664);
and U24419 (N_24419,N_23904,N_23652);
nor U24420 (N_24420,N_23656,N_23542);
xor U24421 (N_24421,N_23917,N_23867);
or U24422 (N_24422,N_23817,N_23920);
nand U24423 (N_24423,N_23709,N_23855);
or U24424 (N_24424,N_23856,N_23878);
or U24425 (N_24425,N_23853,N_23540);
nand U24426 (N_24426,N_23942,N_23875);
nor U24427 (N_24427,N_23952,N_23498);
or U24428 (N_24428,N_23653,N_23596);
or U24429 (N_24429,N_23862,N_23859);
xnor U24430 (N_24430,N_23851,N_23442);
xor U24431 (N_24431,N_23783,N_23875);
and U24432 (N_24432,N_23560,N_23605);
xnor U24433 (N_24433,N_23411,N_23836);
and U24434 (N_24434,N_23624,N_23730);
xnor U24435 (N_24435,N_23428,N_23812);
or U24436 (N_24436,N_23926,N_23842);
xnor U24437 (N_24437,N_23824,N_23924);
or U24438 (N_24438,N_23489,N_23628);
nor U24439 (N_24439,N_23523,N_23417);
or U24440 (N_24440,N_23942,N_23898);
nor U24441 (N_24441,N_23858,N_23624);
and U24442 (N_24442,N_23850,N_23716);
nand U24443 (N_24443,N_23737,N_23564);
nor U24444 (N_24444,N_23871,N_23673);
and U24445 (N_24445,N_23893,N_23775);
nand U24446 (N_24446,N_23596,N_23753);
nor U24447 (N_24447,N_23991,N_23683);
nor U24448 (N_24448,N_23520,N_23949);
nand U24449 (N_24449,N_23956,N_23932);
or U24450 (N_24450,N_23650,N_23719);
nor U24451 (N_24451,N_23563,N_23604);
nor U24452 (N_24452,N_23593,N_23920);
nor U24453 (N_24453,N_23670,N_23883);
and U24454 (N_24454,N_23565,N_23492);
nand U24455 (N_24455,N_23993,N_23558);
xnor U24456 (N_24456,N_23581,N_23787);
nor U24457 (N_24457,N_23795,N_23837);
and U24458 (N_24458,N_23883,N_23642);
nor U24459 (N_24459,N_23525,N_23847);
nand U24460 (N_24460,N_23749,N_23867);
nor U24461 (N_24461,N_23428,N_23437);
nor U24462 (N_24462,N_23451,N_23748);
xnor U24463 (N_24463,N_23787,N_23526);
nand U24464 (N_24464,N_23515,N_23684);
or U24465 (N_24465,N_23858,N_23620);
nor U24466 (N_24466,N_23859,N_23960);
or U24467 (N_24467,N_23580,N_23980);
or U24468 (N_24468,N_23997,N_23703);
or U24469 (N_24469,N_23714,N_23697);
and U24470 (N_24470,N_23837,N_23764);
or U24471 (N_24471,N_23831,N_23833);
and U24472 (N_24472,N_23614,N_23872);
and U24473 (N_24473,N_23582,N_23647);
xnor U24474 (N_24474,N_23894,N_23540);
and U24475 (N_24475,N_23947,N_23693);
or U24476 (N_24476,N_23564,N_23919);
nand U24477 (N_24477,N_23574,N_23697);
nor U24478 (N_24478,N_23847,N_23987);
nor U24479 (N_24479,N_23554,N_23929);
and U24480 (N_24480,N_23471,N_23975);
nand U24481 (N_24481,N_23749,N_23979);
and U24482 (N_24482,N_23472,N_23986);
nand U24483 (N_24483,N_23587,N_23704);
nor U24484 (N_24484,N_23821,N_23799);
or U24485 (N_24485,N_23978,N_23882);
xnor U24486 (N_24486,N_23666,N_23767);
nor U24487 (N_24487,N_23597,N_23629);
or U24488 (N_24488,N_23971,N_23557);
xnor U24489 (N_24489,N_23943,N_23954);
and U24490 (N_24490,N_23729,N_23741);
xnor U24491 (N_24491,N_23762,N_23911);
xnor U24492 (N_24492,N_23642,N_23675);
and U24493 (N_24493,N_23764,N_23667);
or U24494 (N_24494,N_23826,N_23939);
nand U24495 (N_24495,N_23625,N_23487);
and U24496 (N_24496,N_23550,N_23736);
xor U24497 (N_24497,N_23632,N_23559);
or U24498 (N_24498,N_23680,N_23611);
xnor U24499 (N_24499,N_23626,N_23438);
or U24500 (N_24500,N_23729,N_23934);
xor U24501 (N_24501,N_23703,N_23816);
or U24502 (N_24502,N_23401,N_23472);
nand U24503 (N_24503,N_23440,N_23831);
nand U24504 (N_24504,N_23886,N_23418);
or U24505 (N_24505,N_23573,N_23696);
nor U24506 (N_24506,N_23532,N_23744);
or U24507 (N_24507,N_23423,N_23946);
nor U24508 (N_24508,N_23881,N_23949);
and U24509 (N_24509,N_23753,N_23641);
nand U24510 (N_24510,N_23454,N_23877);
or U24511 (N_24511,N_23849,N_23644);
nand U24512 (N_24512,N_23492,N_23590);
and U24513 (N_24513,N_23832,N_23702);
xnor U24514 (N_24514,N_23824,N_23651);
nor U24515 (N_24515,N_23849,N_23695);
xnor U24516 (N_24516,N_23400,N_23679);
and U24517 (N_24517,N_23557,N_23612);
and U24518 (N_24518,N_23613,N_23415);
and U24519 (N_24519,N_23777,N_23875);
xor U24520 (N_24520,N_23985,N_23461);
nor U24521 (N_24521,N_23499,N_23800);
nor U24522 (N_24522,N_23982,N_23778);
nor U24523 (N_24523,N_23696,N_23913);
or U24524 (N_24524,N_23916,N_23982);
or U24525 (N_24525,N_23601,N_23753);
nor U24526 (N_24526,N_23438,N_23970);
and U24527 (N_24527,N_23689,N_23580);
or U24528 (N_24528,N_23646,N_23427);
or U24529 (N_24529,N_23583,N_23850);
nor U24530 (N_24530,N_23795,N_23735);
or U24531 (N_24531,N_23420,N_23601);
nor U24532 (N_24532,N_23928,N_23813);
or U24533 (N_24533,N_23970,N_23512);
nand U24534 (N_24534,N_23566,N_23665);
xor U24535 (N_24535,N_23927,N_23653);
or U24536 (N_24536,N_23636,N_23892);
and U24537 (N_24537,N_23675,N_23807);
nor U24538 (N_24538,N_23769,N_23771);
nand U24539 (N_24539,N_23734,N_23776);
nor U24540 (N_24540,N_23560,N_23958);
or U24541 (N_24541,N_23906,N_23888);
nand U24542 (N_24542,N_23637,N_23475);
and U24543 (N_24543,N_23414,N_23549);
or U24544 (N_24544,N_23956,N_23705);
nor U24545 (N_24545,N_23759,N_23721);
nor U24546 (N_24546,N_23843,N_23846);
and U24547 (N_24547,N_23472,N_23697);
or U24548 (N_24548,N_23533,N_23848);
nand U24549 (N_24549,N_23449,N_23532);
nor U24550 (N_24550,N_23920,N_23523);
nor U24551 (N_24551,N_23931,N_23824);
nand U24552 (N_24552,N_23520,N_23661);
and U24553 (N_24553,N_23457,N_23847);
or U24554 (N_24554,N_23565,N_23673);
nor U24555 (N_24555,N_23612,N_23722);
and U24556 (N_24556,N_23955,N_23868);
and U24557 (N_24557,N_23940,N_23576);
or U24558 (N_24558,N_23738,N_23642);
or U24559 (N_24559,N_23961,N_23404);
nor U24560 (N_24560,N_23984,N_23774);
or U24561 (N_24561,N_23970,N_23773);
nand U24562 (N_24562,N_23676,N_23996);
nor U24563 (N_24563,N_23795,N_23578);
xor U24564 (N_24564,N_23699,N_23928);
or U24565 (N_24565,N_23646,N_23744);
or U24566 (N_24566,N_23461,N_23829);
and U24567 (N_24567,N_23803,N_23686);
nor U24568 (N_24568,N_23704,N_23770);
xnor U24569 (N_24569,N_23504,N_23736);
nor U24570 (N_24570,N_23906,N_23962);
nor U24571 (N_24571,N_23779,N_23829);
xor U24572 (N_24572,N_23972,N_23568);
nor U24573 (N_24573,N_23887,N_23741);
and U24574 (N_24574,N_23890,N_23757);
or U24575 (N_24575,N_23974,N_23791);
nor U24576 (N_24576,N_23410,N_23554);
and U24577 (N_24577,N_23421,N_23740);
and U24578 (N_24578,N_23582,N_23416);
nand U24579 (N_24579,N_23895,N_23892);
xor U24580 (N_24580,N_23864,N_23662);
and U24581 (N_24581,N_23836,N_23726);
and U24582 (N_24582,N_23809,N_23632);
nand U24583 (N_24583,N_23895,N_23631);
or U24584 (N_24584,N_23559,N_23854);
or U24585 (N_24585,N_23995,N_23932);
xnor U24586 (N_24586,N_23432,N_23544);
or U24587 (N_24587,N_23818,N_23452);
nor U24588 (N_24588,N_23587,N_23604);
or U24589 (N_24589,N_23873,N_23753);
nand U24590 (N_24590,N_23607,N_23994);
and U24591 (N_24591,N_23828,N_23865);
nand U24592 (N_24592,N_23679,N_23812);
nand U24593 (N_24593,N_23791,N_23735);
xnor U24594 (N_24594,N_23823,N_23632);
nor U24595 (N_24595,N_23958,N_23425);
or U24596 (N_24596,N_23537,N_23421);
and U24597 (N_24597,N_23448,N_23669);
or U24598 (N_24598,N_23910,N_23680);
xor U24599 (N_24599,N_23914,N_23794);
and U24600 (N_24600,N_24582,N_24214);
nor U24601 (N_24601,N_24161,N_24276);
xnor U24602 (N_24602,N_24425,N_24576);
and U24603 (N_24603,N_24448,N_24092);
or U24604 (N_24604,N_24527,N_24479);
xnor U24605 (N_24605,N_24159,N_24472);
and U24606 (N_24606,N_24247,N_24340);
and U24607 (N_24607,N_24360,N_24329);
and U24608 (N_24608,N_24100,N_24200);
xor U24609 (N_24609,N_24441,N_24573);
nor U24610 (N_24610,N_24241,N_24244);
or U24611 (N_24611,N_24580,N_24506);
nand U24612 (N_24612,N_24139,N_24566);
and U24613 (N_24613,N_24378,N_24598);
and U24614 (N_24614,N_24445,N_24381);
nor U24615 (N_24615,N_24373,N_24518);
xor U24616 (N_24616,N_24228,N_24267);
and U24617 (N_24617,N_24177,N_24334);
nand U24618 (N_24618,N_24254,N_24306);
nand U24619 (N_24619,N_24450,N_24534);
or U24620 (N_24620,N_24204,N_24412);
and U24621 (N_24621,N_24237,N_24415);
nand U24622 (N_24622,N_24560,N_24289);
nand U24623 (N_24623,N_24300,N_24030);
nor U24624 (N_24624,N_24286,N_24122);
nor U24625 (N_24625,N_24256,N_24565);
and U24626 (N_24626,N_24364,N_24368);
or U24627 (N_24627,N_24240,N_24149);
and U24628 (N_24628,N_24206,N_24567);
nand U24629 (N_24629,N_24380,N_24581);
nand U24630 (N_24630,N_24008,N_24321);
and U24631 (N_24631,N_24062,N_24554);
nand U24632 (N_24632,N_24452,N_24317);
or U24633 (N_24633,N_24271,N_24231);
and U24634 (N_24634,N_24191,N_24385);
and U24635 (N_24635,N_24562,N_24355);
or U24636 (N_24636,N_24436,N_24586);
and U24637 (N_24637,N_24398,N_24134);
or U24638 (N_24638,N_24165,N_24215);
or U24639 (N_24639,N_24339,N_24502);
xnor U24640 (N_24640,N_24377,N_24085);
nor U24641 (N_24641,N_24151,N_24195);
nor U24642 (N_24642,N_24496,N_24524);
and U24643 (N_24643,N_24468,N_24067);
and U24644 (N_24644,N_24014,N_24136);
or U24645 (N_24645,N_24293,N_24145);
xnor U24646 (N_24646,N_24235,N_24033);
and U24647 (N_24647,N_24087,N_24375);
nand U24648 (N_24648,N_24034,N_24457);
and U24649 (N_24649,N_24402,N_24279);
or U24650 (N_24650,N_24261,N_24587);
and U24651 (N_24651,N_24048,N_24444);
or U24652 (N_24652,N_24089,N_24113);
nand U24653 (N_24653,N_24110,N_24023);
nor U24654 (N_24654,N_24304,N_24309);
xnor U24655 (N_24655,N_24447,N_24007);
nor U24656 (N_24656,N_24127,N_24564);
or U24657 (N_24657,N_24264,N_24394);
nor U24658 (N_24658,N_24411,N_24262);
or U24659 (N_24659,N_24546,N_24515);
nand U24660 (N_24660,N_24574,N_24266);
nor U24661 (N_24661,N_24212,N_24561);
and U24662 (N_24662,N_24181,N_24156);
nor U24663 (N_24663,N_24084,N_24589);
and U24664 (N_24664,N_24164,N_24491);
nand U24665 (N_24665,N_24349,N_24374);
or U24666 (N_24666,N_24188,N_24318);
nand U24667 (N_24667,N_24397,N_24290);
and U24668 (N_24668,N_24541,N_24405);
nor U24669 (N_24669,N_24201,N_24114);
or U24670 (N_24670,N_24162,N_24115);
or U24671 (N_24671,N_24348,N_24578);
nand U24672 (N_24672,N_24492,N_24210);
or U24673 (N_24673,N_24124,N_24166);
and U24674 (N_24674,N_24253,N_24310);
and U24675 (N_24675,N_24004,N_24484);
and U24676 (N_24676,N_24192,N_24336);
xnor U24677 (N_24677,N_24182,N_24096);
nand U24678 (N_24678,N_24171,N_24446);
and U24679 (N_24679,N_24503,N_24260);
nand U24680 (N_24680,N_24167,N_24391);
xor U24681 (N_24681,N_24035,N_24508);
nor U24682 (N_24682,N_24390,N_24054);
or U24683 (N_24683,N_24430,N_24439);
nor U24684 (N_24684,N_24307,N_24073);
or U24685 (N_24685,N_24265,N_24044);
or U24686 (N_24686,N_24345,N_24388);
and U24687 (N_24687,N_24248,N_24314);
nand U24688 (N_24688,N_24011,N_24514);
or U24689 (N_24689,N_24333,N_24093);
and U24690 (N_24690,N_24507,N_24025);
nand U24691 (N_24691,N_24153,N_24505);
nor U24692 (N_24692,N_24571,N_24474);
nor U24693 (N_24693,N_24437,N_24274);
and U24694 (N_24694,N_24395,N_24434);
and U24695 (N_24695,N_24451,N_24331);
or U24696 (N_24696,N_24190,N_24460);
and U24697 (N_24697,N_24072,N_24088);
and U24698 (N_24698,N_24409,N_24109);
nor U24699 (N_24699,N_24453,N_24098);
xnor U24700 (N_24700,N_24022,N_24401);
nor U24701 (N_24701,N_24046,N_24427);
nor U24702 (N_24702,N_24393,N_24358);
nand U24703 (N_24703,N_24268,N_24140);
nand U24704 (N_24704,N_24488,N_24549);
or U24705 (N_24705,N_24456,N_24226);
nor U24706 (N_24706,N_24440,N_24510);
nor U24707 (N_24707,N_24111,N_24594);
nand U24708 (N_24708,N_24026,N_24197);
or U24709 (N_24709,N_24540,N_24074);
nor U24710 (N_24710,N_24399,N_24179);
nor U24711 (N_24711,N_24057,N_24012);
or U24712 (N_24712,N_24220,N_24094);
or U24713 (N_24713,N_24207,N_24335);
nor U24714 (N_24714,N_24234,N_24218);
or U24715 (N_24715,N_24202,N_24327);
and U24716 (N_24716,N_24275,N_24351);
nand U24717 (N_24717,N_24396,N_24548);
nand U24718 (N_24718,N_24371,N_24176);
nand U24719 (N_24719,N_24282,N_24146);
nand U24720 (N_24720,N_24497,N_24407);
nor U24721 (N_24721,N_24051,N_24223);
xnor U24722 (N_24722,N_24435,N_24525);
and U24723 (N_24723,N_24370,N_24168);
and U24724 (N_24724,N_24121,N_24133);
nor U24725 (N_24725,N_24064,N_24287);
or U24726 (N_24726,N_24079,N_24285);
or U24727 (N_24727,N_24086,N_24043);
and U24728 (N_24728,N_24422,N_24238);
nand U24729 (N_24729,N_24591,N_24366);
nor U24730 (N_24730,N_24353,N_24352);
or U24731 (N_24731,N_24119,N_24350);
nor U24732 (N_24732,N_24438,N_24311);
nor U24733 (N_24733,N_24263,N_24211);
and U24734 (N_24734,N_24229,N_24107);
and U24735 (N_24735,N_24015,N_24294);
or U24736 (N_24736,N_24183,N_24498);
or U24737 (N_24737,N_24481,N_24344);
xor U24738 (N_24738,N_24489,N_24077);
or U24739 (N_24739,N_24028,N_24493);
and U24740 (N_24740,N_24059,N_24475);
and U24741 (N_24741,N_24278,N_24143);
nor U24742 (N_24742,N_24213,N_24083);
nand U24743 (N_24743,N_24376,N_24513);
xor U24744 (N_24744,N_24326,N_24225);
and U24745 (N_24745,N_24270,N_24150);
and U24746 (N_24746,N_24593,N_24157);
or U24747 (N_24747,N_24404,N_24521);
or U24748 (N_24748,N_24575,N_24246);
or U24749 (N_24749,N_24512,N_24049);
and U24750 (N_24750,N_24076,N_24346);
and U24751 (N_24751,N_24584,N_24101);
and U24752 (N_24752,N_24420,N_24550);
or U24753 (N_24753,N_24486,N_24347);
nor U24754 (N_24754,N_24509,N_24466);
or U24755 (N_24755,N_24426,N_24198);
nor U24756 (N_24756,N_24495,N_24147);
nand U24757 (N_24757,N_24099,N_24082);
xnor U24758 (N_24758,N_24019,N_24520);
nor U24759 (N_24759,N_24125,N_24002);
and U24760 (N_24760,N_24583,N_24120);
nor U24761 (N_24761,N_24557,N_24280);
and U24762 (N_24762,N_24330,N_24464);
or U24763 (N_24763,N_24416,N_24563);
and U24764 (N_24764,N_24106,N_24209);
nor U24765 (N_24765,N_24245,N_24185);
or U24766 (N_24766,N_24128,N_24005);
nand U24767 (N_24767,N_24478,N_24555);
nor U24768 (N_24768,N_24537,N_24118);
nand U24769 (N_24769,N_24558,N_24538);
nor U24770 (N_24770,N_24227,N_24470);
xnor U24771 (N_24771,N_24367,N_24112);
nor U24772 (N_24772,N_24383,N_24526);
xnor U24773 (N_24773,N_24539,N_24431);
and U24774 (N_24774,N_24455,N_24163);
nor U24775 (N_24775,N_24047,N_24018);
and U24776 (N_24776,N_24467,N_24403);
and U24777 (N_24777,N_24053,N_24522);
nand U24778 (N_24778,N_24090,N_24081);
nand U24779 (N_24779,N_24588,N_24042);
or U24780 (N_24780,N_24001,N_24596);
or U24781 (N_24781,N_24408,N_24230);
nand U24782 (N_24782,N_24559,N_24061);
xnor U24783 (N_24783,N_24239,N_24308);
xnor U24784 (N_24784,N_24418,N_24442);
nor U24785 (N_24785,N_24324,N_24499);
and U24786 (N_24786,N_24013,N_24342);
nor U24787 (N_24787,N_24219,N_24568);
nor U24788 (N_24788,N_24194,N_24462);
nand U24789 (N_24789,N_24116,N_24516);
nand U24790 (N_24790,N_24095,N_24003);
nor U24791 (N_24791,N_24216,N_24531);
nand U24792 (N_24792,N_24320,N_24429);
and U24793 (N_24793,N_24322,N_24363);
xor U24794 (N_24794,N_24424,N_24006);
nand U24795 (N_24795,N_24313,N_24205);
or U24796 (N_24796,N_24052,N_24292);
and U24797 (N_24797,N_24108,N_24528);
and U24798 (N_24798,N_24104,N_24102);
and U24799 (N_24799,N_24536,N_24454);
or U24800 (N_24800,N_24193,N_24433);
and U24801 (N_24801,N_24039,N_24080);
nor U24802 (N_24802,N_24414,N_24458);
nand U24803 (N_24803,N_24585,N_24020);
or U24804 (N_24804,N_24459,N_24511);
and U24805 (N_24805,N_24530,N_24523);
nor U24806 (N_24806,N_24590,N_24301);
and U24807 (N_24807,N_24259,N_24032);
or U24808 (N_24808,N_24251,N_24400);
nand U24809 (N_24809,N_24535,N_24480);
or U24810 (N_24810,N_24010,N_24572);
nor U24811 (N_24811,N_24075,N_24142);
nand U24812 (N_24812,N_24196,N_24545);
or U24813 (N_24813,N_24302,N_24419);
nand U24814 (N_24814,N_24105,N_24490);
nand U24815 (N_24815,N_24174,N_24291);
or U24816 (N_24816,N_24410,N_24131);
nor U24817 (N_24817,N_24471,N_24144);
or U24818 (N_24818,N_24063,N_24386);
nand U24819 (N_24819,N_24553,N_24362);
and U24820 (N_24820,N_24221,N_24135);
or U24821 (N_24821,N_24141,N_24243);
and U24822 (N_24822,N_24504,N_24384);
and U24823 (N_24823,N_24298,N_24357);
and U24824 (N_24824,N_24038,N_24337);
and U24825 (N_24825,N_24570,N_24543);
or U24826 (N_24826,N_24529,N_24041);
or U24827 (N_24827,N_24569,N_24222);
and U24828 (N_24828,N_24060,N_24233);
nand U24829 (N_24829,N_24487,N_24449);
xnor U24830 (N_24830,N_24485,N_24392);
nor U24831 (N_24831,N_24242,N_24186);
nor U24832 (N_24832,N_24117,N_24172);
nand U24833 (N_24833,N_24372,N_24483);
nand U24834 (N_24834,N_24078,N_24597);
nor U24835 (N_24835,N_24066,N_24305);
and U24836 (N_24836,N_24443,N_24379);
and U24837 (N_24837,N_24519,N_24097);
nor U24838 (N_24838,N_24138,N_24547);
and U24839 (N_24839,N_24236,N_24272);
and U24840 (N_24840,N_24056,N_24232);
and U24841 (N_24841,N_24316,N_24417);
nor U24842 (N_24842,N_24199,N_24423);
nor U24843 (N_24843,N_24065,N_24387);
or U24844 (N_24844,N_24130,N_24413);
and U24845 (N_24845,N_24252,N_24432);
nand U24846 (N_24846,N_24169,N_24461);
and U24847 (N_24847,N_24517,N_24189);
nand U24848 (N_24848,N_24354,N_24132);
xnor U24849 (N_24849,N_24017,N_24055);
nand U24850 (N_24850,N_24180,N_24465);
and U24851 (N_24851,N_24250,N_24369);
and U24852 (N_24852,N_24482,N_24269);
nor U24853 (N_24853,N_24069,N_24257);
nor U24854 (N_24854,N_24359,N_24137);
and U24855 (N_24855,N_24071,N_24070);
xor U24856 (N_24856,N_24551,N_24592);
nor U24857 (N_24857,N_24009,N_24152);
xor U24858 (N_24858,N_24361,N_24343);
or U24859 (N_24859,N_24031,N_24338);
or U24860 (N_24860,N_24170,N_24428);
and U24861 (N_24861,N_24068,N_24577);
nand U24862 (N_24862,N_24160,N_24341);
and U24863 (N_24863,N_24158,N_24382);
nand U24864 (N_24864,N_24532,N_24421);
nand U24865 (N_24865,N_24103,N_24303);
nor U24866 (N_24866,N_24389,N_24552);
nor U24867 (N_24867,N_24297,N_24494);
nand U24868 (N_24868,N_24154,N_24365);
nor U24869 (N_24869,N_24277,N_24544);
nor U24870 (N_24870,N_24473,N_24469);
nand U24871 (N_24871,N_24178,N_24024);
and U24872 (N_24872,N_24155,N_24126);
nand U24873 (N_24873,N_24477,N_24000);
and U24874 (N_24874,N_24299,N_24315);
and U24875 (N_24875,N_24045,N_24016);
or U24876 (N_24876,N_24123,N_24021);
or U24877 (N_24877,N_24173,N_24187);
nand U24878 (N_24878,N_24312,N_24281);
nor U24879 (N_24879,N_24050,N_24283);
xor U24880 (N_24880,N_24027,N_24029);
nor U24881 (N_24881,N_24501,N_24476);
or U24882 (N_24882,N_24595,N_24273);
xor U24883 (N_24883,N_24296,N_24203);
nand U24884 (N_24884,N_24323,N_24091);
and U24885 (N_24885,N_24175,N_24258);
nor U24886 (N_24886,N_24224,N_24208);
xnor U24887 (N_24887,N_24129,N_24406);
nor U24888 (N_24888,N_24037,N_24332);
nand U24889 (N_24889,N_24325,N_24148);
xnor U24890 (N_24890,N_24184,N_24533);
nand U24891 (N_24891,N_24255,N_24319);
nor U24892 (N_24892,N_24500,N_24579);
xnor U24893 (N_24893,N_24288,N_24058);
and U24894 (N_24894,N_24036,N_24249);
or U24895 (N_24895,N_24284,N_24356);
nand U24896 (N_24896,N_24599,N_24556);
nor U24897 (N_24897,N_24463,N_24328);
or U24898 (N_24898,N_24542,N_24295);
or U24899 (N_24899,N_24217,N_24040);
nor U24900 (N_24900,N_24527,N_24082);
and U24901 (N_24901,N_24203,N_24337);
or U24902 (N_24902,N_24079,N_24494);
nor U24903 (N_24903,N_24195,N_24240);
xnor U24904 (N_24904,N_24309,N_24420);
nand U24905 (N_24905,N_24106,N_24323);
and U24906 (N_24906,N_24313,N_24014);
and U24907 (N_24907,N_24330,N_24451);
or U24908 (N_24908,N_24185,N_24459);
and U24909 (N_24909,N_24139,N_24596);
nor U24910 (N_24910,N_24155,N_24136);
nor U24911 (N_24911,N_24277,N_24562);
or U24912 (N_24912,N_24500,N_24263);
and U24913 (N_24913,N_24328,N_24386);
xnor U24914 (N_24914,N_24076,N_24361);
or U24915 (N_24915,N_24393,N_24120);
nand U24916 (N_24916,N_24470,N_24334);
or U24917 (N_24917,N_24222,N_24551);
or U24918 (N_24918,N_24080,N_24127);
and U24919 (N_24919,N_24337,N_24228);
nand U24920 (N_24920,N_24521,N_24143);
nor U24921 (N_24921,N_24340,N_24401);
and U24922 (N_24922,N_24084,N_24456);
or U24923 (N_24923,N_24192,N_24517);
nand U24924 (N_24924,N_24031,N_24262);
nor U24925 (N_24925,N_24187,N_24004);
nor U24926 (N_24926,N_24054,N_24162);
nor U24927 (N_24927,N_24211,N_24248);
and U24928 (N_24928,N_24370,N_24198);
xor U24929 (N_24929,N_24049,N_24454);
and U24930 (N_24930,N_24250,N_24089);
or U24931 (N_24931,N_24362,N_24244);
nand U24932 (N_24932,N_24320,N_24544);
and U24933 (N_24933,N_24586,N_24300);
nor U24934 (N_24934,N_24069,N_24100);
or U24935 (N_24935,N_24338,N_24218);
nand U24936 (N_24936,N_24022,N_24532);
and U24937 (N_24937,N_24282,N_24083);
xor U24938 (N_24938,N_24019,N_24169);
or U24939 (N_24939,N_24367,N_24352);
nor U24940 (N_24940,N_24422,N_24042);
nand U24941 (N_24941,N_24527,N_24118);
and U24942 (N_24942,N_24135,N_24515);
and U24943 (N_24943,N_24467,N_24255);
xnor U24944 (N_24944,N_24004,N_24449);
or U24945 (N_24945,N_24537,N_24362);
or U24946 (N_24946,N_24209,N_24171);
or U24947 (N_24947,N_24056,N_24264);
nand U24948 (N_24948,N_24165,N_24013);
and U24949 (N_24949,N_24272,N_24596);
nor U24950 (N_24950,N_24591,N_24211);
and U24951 (N_24951,N_24052,N_24334);
xor U24952 (N_24952,N_24219,N_24431);
or U24953 (N_24953,N_24355,N_24188);
nand U24954 (N_24954,N_24024,N_24129);
nand U24955 (N_24955,N_24033,N_24259);
nor U24956 (N_24956,N_24132,N_24206);
nand U24957 (N_24957,N_24098,N_24212);
or U24958 (N_24958,N_24463,N_24357);
nor U24959 (N_24959,N_24360,N_24428);
nand U24960 (N_24960,N_24022,N_24129);
nor U24961 (N_24961,N_24281,N_24243);
or U24962 (N_24962,N_24352,N_24106);
nand U24963 (N_24963,N_24210,N_24241);
nand U24964 (N_24964,N_24388,N_24000);
or U24965 (N_24965,N_24070,N_24036);
or U24966 (N_24966,N_24416,N_24225);
and U24967 (N_24967,N_24398,N_24548);
nand U24968 (N_24968,N_24156,N_24145);
nand U24969 (N_24969,N_24307,N_24063);
nand U24970 (N_24970,N_24226,N_24202);
xnor U24971 (N_24971,N_24549,N_24223);
nor U24972 (N_24972,N_24081,N_24589);
nor U24973 (N_24973,N_24443,N_24086);
nand U24974 (N_24974,N_24018,N_24475);
or U24975 (N_24975,N_24399,N_24299);
and U24976 (N_24976,N_24419,N_24274);
xnor U24977 (N_24977,N_24271,N_24326);
xor U24978 (N_24978,N_24155,N_24152);
nand U24979 (N_24979,N_24291,N_24180);
or U24980 (N_24980,N_24321,N_24152);
or U24981 (N_24981,N_24011,N_24010);
nor U24982 (N_24982,N_24144,N_24450);
or U24983 (N_24983,N_24579,N_24055);
or U24984 (N_24984,N_24313,N_24551);
nand U24985 (N_24985,N_24473,N_24072);
or U24986 (N_24986,N_24117,N_24437);
nor U24987 (N_24987,N_24010,N_24545);
nand U24988 (N_24988,N_24523,N_24161);
nor U24989 (N_24989,N_24542,N_24121);
and U24990 (N_24990,N_24463,N_24330);
nor U24991 (N_24991,N_24176,N_24512);
nand U24992 (N_24992,N_24355,N_24456);
nor U24993 (N_24993,N_24170,N_24471);
nor U24994 (N_24994,N_24405,N_24510);
nor U24995 (N_24995,N_24020,N_24281);
and U24996 (N_24996,N_24117,N_24239);
and U24997 (N_24997,N_24438,N_24089);
or U24998 (N_24998,N_24548,N_24422);
nor U24999 (N_24999,N_24070,N_24259);
nand U25000 (N_25000,N_24076,N_24581);
xnor U25001 (N_25001,N_24029,N_24387);
nand U25002 (N_25002,N_24117,N_24328);
and U25003 (N_25003,N_24166,N_24135);
and U25004 (N_25004,N_24506,N_24514);
and U25005 (N_25005,N_24146,N_24341);
nor U25006 (N_25006,N_24383,N_24572);
and U25007 (N_25007,N_24248,N_24032);
or U25008 (N_25008,N_24325,N_24117);
nand U25009 (N_25009,N_24243,N_24180);
and U25010 (N_25010,N_24506,N_24161);
nand U25011 (N_25011,N_24034,N_24124);
nor U25012 (N_25012,N_24100,N_24366);
nor U25013 (N_25013,N_24118,N_24385);
or U25014 (N_25014,N_24498,N_24394);
nor U25015 (N_25015,N_24173,N_24015);
or U25016 (N_25016,N_24263,N_24570);
xor U25017 (N_25017,N_24494,N_24376);
nand U25018 (N_25018,N_24034,N_24430);
nand U25019 (N_25019,N_24135,N_24277);
nor U25020 (N_25020,N_24127,N_24155);
and U25021 (N_25021,N_24449,N_24276);
and U25022 (N_25022,N_24574,N_24282);
nor U25023 (N_25023,N_24582,N_24139);
or U25024 (N_25024,N_24433,N_24569);
and U25025 (N_25025,N_24199,N_24044);
or U25026 (N_25026,N_24310,N_24062);
and U25027 (N_25027,N_24580,N_24437);
and U25028 (N_25028,N_24113,N_24421);
xor U25029 (N_25029,N_24464,N_24016);
or U25030 (N_25030,N_24598,N_24376);
nand U25031 (N_25031,N_24244,N_24318);
nand U25032 (N_25032,N_24465,N_24307);
nor U25033 (N_25033,N_24421,N_24267);
nor U25034 (N_25034,N_24149,N_24473);
nor U25035 (N_25035,N_24478,N_24434);
nand U25036 (N_25036,N_24187,N_24146);
nor U25037 (N_25037,N_24134,N_24457);
nor U25038 (N_25038,N_24394,N_24563);
nor U25039 (N_25039,N_24580,N_24154);
and U25040 (N_25040,N_24076,N_24270);
nand U25041 (N_25041,N_24111,N_24168);
nand U25042 (N_25042,N_24289,N_24471);
nor U25043 (N_25043,N_24128,N_24540);
and U25044 (N_25044,N_24363,N_24237);
nor U25045 (N_25045,N_24001,N_24439);
nor U25046 (N_25046,N_24487,N_24058);
xor U25047 (N_25047,N_24297,N_24484);
xor U25048 (N_25048,N_24035,N_24312);
and U25049 (N_25049,N_24586,N_24202);
or U25050 (N_25050,N_24123,N_24078);
nor U25051 (N_25051,N_24069,N_24078);
and U25052 (N_25052,N_24062,N_24456);
nand U25053 (N_25053,N_24303,N_24546);
nand U25054 (N_25054,N_24323,N_24281);
and U25055 (N_25055,N_24003,N_24464);
nand U25056 (N_25056,N_24309,N_24214);
nand U25057 (N_25057,N_24510,N_24453);
and U25058 (N_25058,N_24090,N_24599);
or U25059 (N_25059,N_24045,N_24435);
nor U25060 (N_25060,N_24464,N_24336);
nor U25061 (N_25061,N_24229,N_24279);
nand U25062 (N_25062,N_24345,N_24391);
nor U25063 (N_25063,N_24182,N_24281);
or U25064 (N_25064,N_24130,N_24204);
and U25065 (N_25065,N_24530,N_24156);
and U25066 (N_25066,N_24020,N_24163);
nor U25067 (N_25067,N_24480,N_24366);
and U25068 (N_25068,N_24367,N_24291);
and U25069 (N_25069,N_24102,N_24059);
or U25070 (N_25070,N_24310,N_24325);
nand U25071 (N_25071,N_24517,N_24495);
xnor U25072 (N_25072,N_24328,N_24151);
or U25073 (N_25073,N_24544,N_24268);
nor U25074 (N_25074,N_24571,N_24153);
and U25075 (N_25075,N_24303,N_24322);
or U25076 (N_25076,N_24436,N_24275);
nor U25077 (N_25077,N_24087,N_24215);
or U25078 (N_25078,N_24516,N_24029);
xnor U25079 (N_25079,N_24283,N_24512);
nor U25080 (N_25080,N_24360,N_24048);
nand U25081 (N_25081,N_24339,N_24247);
xor U25082 (N_25082,N_24169,N_24548);
nor U25083 (N_25083,N_24061,N_24104);
or U25084 (N_25084,N_24387,N_24081);
nand U25085 (N_25085,N_24274,N_24552);
nor U25086 (N_25086,N_24101,N_24120);
nand U25087 (N_25087,N_24394,N_24571);
or U25088 (N_25088,N_24383,N_24481);
and U25089 (N_25089,N_24556,N_24238);
and U25090 (N_25090,N_24097,N_24102);
nand U25091 (N_25091,N_24593,N_24216);
nand U25092 (N_25092,N_24092,N_24031);
nor U25093 (N_25093,N_24358,N_24274);
nand U25094 (N_25094,N_24317,N_24284);
or U25095 (N_25095,N_24268,N_24462);
and U25096 (N_25096,N_24530,N_24147);
and U25097 (N_25097,N_24259,N_24223);
and U25098 (N_25098,N_24402,N_24161);
nor U25099 (N_25099,N_24130,N_24064);
or U25100 (N_25100,N_24232,N_24013);
xor U25101 (N_25101,N_24161,N_24097);
and U25102 (N_25102,N_24108,N_24301);
nand U25103 (N_25103,N_24331,N_24579);
xor U25104 (N_25104,N_24317,N_24363);
and U25105 (N_25105,N_24409,N_24265);
nand U25106 (N_25106,N_24159,N_24543);
or U25107 (N_25107,N_24450,N_24487);
and U25108 (N_25108,N_24224,N_24331);
nand U25109 (N_25109,N_24132,N_24219);
or U25110 (N_25110,N_24042,N_24488);
nand U25111 (N_25111,N_24178,N_24007);
or U25112 (N_25112,N_24076,N_24384);
nand U25113 (N_25113,N_24073,N_24160);
nor U25114 (N_25114,N_24587,N_24209);
or U25115 (N_25115,N_24281,N_24287);
nand U25116 (N_25116,N_24574,N_24072);
and U25117 (N_25117,N_24309,N_24176);
nor U25118 (N_25118,N_24136,N_24455);
nor U25119 (N_25119,N_24172,N_24583);
nand U25120 (N_25120,N_24166,N_24571);
or U25121 (N_25121,N_24594,N_24323);
nor U25122 (N_25122,N_24184,N_24103);
and U25123 (N_25123,N_24593,N_24052);
xor U25124 (N_25124,N_24464,N_24490);
and U25125 (N_25125,N_24330,N_24249);
or U25126 (N_25126,N_24407,N_24047);
or U25127 (N_25127,N_24411,N_24168);
nor U25128 (N_25128,N_24011,N_24133);
nor U25129 (N_25129,N_24146,N_24595);
xnor U25130 (N_25130,N_24354,N_24170);
nand U25131 (N_25131,N_24162,N_24290);
nand U25132 (N_25132,N_24078,N_24384);
and U25133 (N_25133,N_24138,N_24460);
and U25134 (N_25134,N_24362,N_24272);
or U25135 (N_25135,N_24409,N_24453);
nand U25136 (N_25136,N_24212,N_24396);
or U25137 (N_25137,N_24531,N_24417);
and U25138 (N_25138,N_24225,N_24072);
nor U25139 (N_25139,N_24036,N_24089);
and U25140 (N_25140,N_24593,N_24413);
or U25141 (N_25141,N_24410,N_24102);
and U25142 (N_25142,N_24341,N_24403);
or U25143 (N_25143,N_24342,N_24330);
nand U25144 (N_25144,N_24228,N_24029);
and U25145 (N_25145,N_24097,N_24077);
xnor U25146 (N_25146,N_24470,N_24111);
and U25147 (N_25147,N_24144,N_24040);
nor U25148 (N_25148,N_24289,N_24122);
and U25149 (N_25149,N_24106,N_24099);
xnor U25150 (N_25150,N_24434,N_24504);
nor U25151 (N_25151,N_24345,N_24464);
or U25152 (N_25152,N_24330,N_24224);
nand U25153 (N_25153,N_24323,N_24399);
nand U25154 (N_25154,N_24015,N_24078);
and U25155 (N_25155,N_24131,N_24590);
xor U25156 (N_25156,N_24525,N_24233);
and U25157 (N_25157,N_24126,N_24054);
and U25158 (N_25158,N_24493,N_24291);
xor U25159 (N_25159,N_24324,N_24119);
and U25160 (N_25160,N_24083,N_24097);
nor U25161 (N_25161,N_24395,N_24520);
or U25162 (N_25162,N_24469,N_24272);
nand U25163 (N_25163,N_24020,N_24542);
xor U25164 (N_25164,N_24064,N_24173);
nor U25165 (N_25165,N_24050,N_24019);
and U25166 (N_25166,N_24248,N_24427);
and U25167 (N_25167,N_24445,N_24058);
and U25168 (N_25168,N_24279,N_24119);
or U25169 (N_25169,N_24597,N_24100);
or U25170 (N_25170,N_24047,N_24279);
and U25171 (N_25171,N_24179,N_24225);
nand U25172 (N_25172,N_24269,N_24355);
nand U25173 (N_25173,N_24150,N_24576);
xnor U25174 (N_25174,N_24287,N_24525);
or U25175 (N_25175,N_24320,N_24243);
nand U25176 (N_25176,N_24586,N_24031);
and U25177 (N_25177,N_24029,N_24505);
nand U25178 (N_25178,N_24372,N_24110);
or U25179 (N_25179,N_24041,N_24149);
nand U25180 (N_25180,N_24398,N_24359);
xor U25181 (N_25181,N_24083,N_24278);
nor U25182 (N_25182,N_24165,N_24592);
nand U25183 (N_25183,N_24222,N_24022);
nor U25184 (N_25184,N_24549,N_24119);
and U25185 (N_25185,N_24254,N_24341);
or U25186 (N_25186,N_24526,N_24226);
or U25187 (N_25187,N_24412,N_24219);
and U25188 (N_25188,N_24013,N_24178);
nand U25189 (N_25189,N_24209,N_24093);
and U25190 (N_25190,N_24583,N_24209);
and U25191 (N_25191,N_24384,N_24343);
and U25192 (N_25192,N_24422,N_24472);
nand U25193 (N_25193,N_24222,N_24149);
or U25194 (N_25194,N_24436,N_24582);
nand U25195 (N_25195,N_24410,N_24244);
xnor U25196 (N_25196,N_24067,N_24512);
nand U25197 (N_25197,N_24208,N_24598);
nor U25198 (N_25198,N_24410,N_24447);
and U25199 (N_25199,N_24098,N_24127);
nand U25200 (N_25200,N_25196,N_24962);
or U25201 (N_25201,N_25035,N_24773);
nand U25202 (N_25202,N_24879,N_24911);
or U25203 (N_25203,N_24667,N_24774);
or U25204 (N_25204,N_24820,N_25191);
nand U25205 (N_25205,N_24945,N_25033);
and U25206 (N_25206,N_25128,N_25134);
or U25207 (N_25207,N_25030,N_25151);
nand U25208 (N_25208,N_24842,N_24872);
or U25209 (N_25209,N_25192,N_25157);
nor U25210 (N_25210,N_24968,N_24764);
nand U25211 (N_25211,N_25029,N_24873);
or U25212 (N_25212,N_24678,N_25153);
nand U25213 (N_25213,N_24643,N_24955);
or U25214 (N_25214,N_24960,N_24626);
and U25215 (N_25215,N_24659,N_24966);
or U25216 (N_25216,N_25082,N_25154);
or U25217 (N_25217,N_25050,N_25100);
or U25218 (N_25218,N_24909,N_24613);
and U25219 (N_25219,N_25039,N_25062);
or U25220 (N_25220,N_24767,N_24937);
nand U25221 (N_25221,N_25049,N_24699);
or U25222 (N_25222,N_24615,N_24660);
or U25223 (N_25223,N_24923,N_24727);
and U25224 (N_25224,N_24834,N_24738);
nor U25225 (N_25225,N_24681,N_25195);
and U25226 (N_25226,N_24698,N_25112);
nand U25227 (N_25227,N_24928,N_24953);
nand U25228 (N_25228,N_24910,N_25102);
nand U25229 (N_25229,N_24722,N_25105);
xnor U25230 (N_25230,N_25115,N_24694);
nand U25231 (N_25231,N_24841,N_25043);
and U25232 (N_25232,N_25048,N_25013);
or U25233 (N_25233,N_24925,N_25199);
or U25234 (N_25234,N_24724,N_25011);
nand U25235 (N_25235,N_25190,N_24739);
xor U25236 (N_25236,N_25149,N_24623);
and U25237 (N_25237,N_24988,N_24757);
and U25238 (N_25238,N_25012,N_24870);
or U25239 (N_25239,N_25074,N_25131);
or U25240 (N_25240,N_25124,N_24862);
nand U25241 (N_25241,N_24935,N_25120);
and U25242 (N_25242,N_24705,N_24737);
nand U25243 (N_25243,N_24632,N_24712);
nand U25244 (N_25244,N_24624,N_24830);
nor U25245 (N_25245,N_24703,N_24800);
and U25246 (N_25246,N_25023,N_24895);
or U25247 (N_25247,N_24979,N_25066);
and U25248 (N_25248,N_25025,N_24817);
xor U25249 (N_25249,N_24832,N_24642);
nor U25250 (N_25250,N_25000,N_25178);
and U25251 (N_25251,N_24707,N_24798);
nand U25252 (N_25252,N_24686,N_25089);
nand U25253 (N_25253,N_24696,N_25047);
and U25254 (N_25254,N_24889,N_25179);
or U25255 (N_25255,N_24628,N_25129);
nor U25256 (N_25256,N_24813,N_25072);
or U25257 (N_25257,N_24714,N_25180);
and U25258 (N_25258,N_24876,N_24689);
and U25259 (N_25259,N_25093,N_25144);
or U25260 (N_25260,N_24864,N_25171);
and U25261 (N_25261,N_25143,N_25007);
xnor U25262 (N_25262,N_24908,N_25136);
or U25263 (N_25263,N_24922,N_25032);
or U25264 (N_25264,N_25004,N_24904);
nand U25265 (N_25265,N_24947,N_24652);
nand U25266 (N_25266,N_24975,N_24827);
or U25267 (N_25267,N_25160,N_25034);
and U25268 (N_25268,N_24723,N_25140);
or U25269 (N_25269,N_25070,N_24636);
or U25270 (N_25270,N_25064,N_24963);
and U25271 (N_25271,N_25168,N_24846);
nand U25272 (N_25272,N_24944,N_24987);
and U25273 (N_25273,N_25107,N_25158);
and U25274 (N_25274,N_24796,N_24608);
nor U25275 (N_25275,N_24651,N_24679);
and U25276 (N_25276,N_24951,N_24753);
nor U25277 (N_25277,N_24690,N_24666);
and U25278 (N_25278,N_24758,N_24663);
nand U25279 (N_25279,N_25113,N_24620);
nand U25280 (N_25280,N_24989,N_24932);
nor U25281 (N_25281,N_25162,N_24805);
nor U25282 (N_25282,N_24756,N_25078);
nand U25283 (N_25283,N_24957,N_25014);
nand U25284 (N_25284,N_25185,N_25150);
or U25285 (N_25285,N_24625,N_24631);
and U25286 (N_25286,N_25016,N_24985);
xor U25287 (N_25287,N_24638,N_24969);
nand U25288 (N_25288,N_24839,N_24622);
or U25289 (N_25289,N_24728,N_24677);
nand U25290 (N_25290,N_24715,N_24760);
nor U25291 (N_25291,N_25063,N_25044);
and U25292 (N_25292,N_24617,N_25104);
xor U25293 (N_25293,N_24890,N_25197);
and U25294 (N_25294,N_24629,N_24614);
nand U25295 (N_25295,N_24956,N_24888);
and U25296 (N_25296,N_25056,N_24853);
and U25297 (N_25297,N_24995,N_24740);
xor U25298 (N_25298,N_25094,N_24627);
and U25299 (N_25299,N_25036,N_25139);
or U25300 (N_25300,N_24790,N_24648);
and U25301 (N_25301,N_24828,N_24754);
nand U25302 (N_25302,N_24967,N_24885);
and U25303 (N_25303,N_25127,N_24996);
and U25304 (N_25304,N_24831,N_24863);
xnor U25305 (N_25305,N_25132,N_25164);
or U25306 (N_25306,N_24693,N_24902);
nor U25307 (N_25307,N_24609,N_24942);
nand U25308 (N_25308,N_24840,N_24769);
nand U25309 (N_25309,N_24994,N_24915);
and U25310 (N_25310,N_24905,N_24761);
nor U25311 (N_25311,N_24797,N_25075);
or U25312 (N_25312,N_24640,N_25020);
and U25313 (N_25313,N_24893,N_24751);
and U25314 (N_25314,N_24986,N_24752);
or U25315 (N_25315,N_24824,N_25121);
nand U25316 (N_25316,N_24765,N_24946);
or U25317 (N_25317,N_25077,N_24771);
nand U25318 (N_25318,N_24743,N_24772);
or U25319 (N_25319,N_24734,N_24821);
xor U25320 (N_25320,N_24600,N_24822);
nand U25321 (N_25321,N_25015,N_25116);
and U25322 (N_25322,N_24976,N_24793);
or U25323 (N_25323,N_24861,N_24646);
xnor U25324 (N_25324,N_24886,N_24656);
xnor U25325 (N_25325,N_24649,N_24984);
nand U25326 (N_25326,N_24786,N_25040);
nor U25327 (N_25327,N_24692,N_24683);
or U25328 (N_25328,N_24768,N_24662);
nor U25329 (N_25329,N_25123,N_24744);
nor U25330 (N_25330,N_25001,N_24639);
and U25331 (N_25331,N_24949,N_25103);
or U25332 (N_25332,N_24982,N_24924);
nand U25333 (N_25333,N_25084,N_25059);
nor U25334 (N_25334,N_24725,N_24778);
and U25335 (N_25335,N_24784,N_25122);
or U25336 (N_25336,N_24671,N_24837);
nor U25337 (N_25337,N_25182,N_25085);
nor U25338 (N_25338,N_24606,N_25073);
and U25339 (N_25339,N_24981,N_24933);
and U25340 (N_25340,N_24990,N_24763);
or U25341 (N_25341,N_25133,N_24941);
nor U25342 (N_25342,N_24731,N_25163);
and U25343 (N_25343,N_24780,N_24802);
nor U25344 (N_25344,N_24914,N_24602);
and U25345 (N_25345,N_24826,N_24611);
nor U25346 (N_25346,N_24898,N_24920);
xor U25347 (N_25347,N_24630,N_25053);
xnor U25348 (N_25348,N_24973,N_25137);
nor U25349 (N_25349,N_25135,N_24661);
or U25350 (N_25350,N_25096,N_24897);
and U25351 (N_25351,N_25161,N_24672);
nand U25352 (N_25352,N_24717,N_24687);
or U25353 (N_25353,N_24972,N_24647);
or U25354 (N_25354,N_25028,N_24637);
or U25355 (N_25355,N_24791,N_24934);
and U25356 (N_25356,N_24892,N_24847);
or U25357 (N_25357,N_24604,N_24766);
and U25358 (N_25358,N_24799,N_24815);
nand U25359 (N_25359,N_24749,N_24748);
nand U25360 (N_25360,N_24779,N_24977);
nand U25361 (N_25361,N_25106,N_25187);
or U25362 (N_25362,N_24880,N_24843);
xnor U25363 (N_25363,N_24891,N_24788);
nor U25364 (N_25364,N_25099,N_24812);
nor U25365 (N_25365,N_24718,N_24998);
and U25366 (N_25366,N_24811,N_25159);
nor U25367 (N_25367,N_24903,N_24850);
xor U25368 (N_25368,N_25156,N_24869);
or U25369 (N_25369,N_25046,N_24948);
nand U25370 (N_25370,N_24653,N_24709);
or U25371 (N_25371,N_24755,N_25147);
xor U25372 (N_25372,N_25087,N_24776);
nand U25373 (N_25373,N_25008,N_24896);
xnor U25374 (N_25374,N_24710,N_24618);
nor U25375 (N_25375,N_24803,N_24871);
or U25376 (N_25376,N_24697,N_24645);
xor U25377 (N_25377,N_25017,N_25186);
or U25378 (N_25378,N_24838,N_24675);
and U25379 (N_25379,N_24787,N_25010);
nor U25380 (N_25380,N_25022,N_24745);
nor U25381 (N_25381,N_25198,N_25126);
nand U25382 (N_25382,N_25021,N_24736);
nand U25383 (N_25383,N_24999,N_25173);
or U25384 (N_25384,N_25111,N_25145);
xnor U25385 (N_25385,N_24641,N_24921);
and U25386 (N_25386,N_25108,N_24810);
nor U25387 (N_25387,N_24954,N_25086);
or U25388 (N_25388,N_24819,N_24866);
nor U25389 (N_25389,N_24829,N_25042);
or U25390 (N_25390,N_24719,N_25183);
and U25391 (N_25391,N_25076,N_24650);
or U25392 (N_25392,N_24936,N_25055);
nand U25393 (N_25393,N_24877,N_24865);
nand U25394 (N_25394,N_25069,N_24655);
or U25395 (N_25395,N_25189,N_24759);
nor U25396 (N_25396,N_24881,N_24695);
nor U25397 (N_25397,N_25081,N_25117);
xnor U25398 (N_25398,N_24792,N_25091);
or U25399 (N_25399,N_24775,N_25052);
nand U25400 (N_25400,N_24634,N_24906);
nand U25401 (N_25401,N_24742,N_24732);
and U25402 (N_25402,N_24894,N_24711);
nor U25403 (N_25403,N_24916,N_24918);
nor U25404 (N_25404,N_24721,N_24974);
nor U25405 (N_25405,N_25057,N_25167);
nor U25406 (N_25406,N_24852,N_24701);
nand U25407 (N_25407,N_24702,N_24993);
and U25408 (N_25408,N_25027,N_24927);
nor U25409 (N_25409,N_24619,N_24612);
nand U25410 (N_25410,N_24913,N_24929);
xnor U25411 (N_25411,N_24808,N_24868);
xnor U25412 (N_25412,N_25061,N_25002);
nor U25413 (N_25413,N_25009,N_25006);
nand U25414 (N_25414,N_25142,N_25079);
and U25415 (N_25415,N_24807,N_25155);
xor U25416 (N_25416,N_24912,N_25060);
and U25417 (N_25417,N_24919,N_24635);
or U25418 (N_25418,N_24644,N_24726);
nand U25419 (N_25419,N_25037,N_24729);
nor U25420 (N_25420,N_25194,N_24716);
nor U25421 (N_25421,N_25175,N_24848);
or U25422 (N_25422,N_24783,N_25152);
nor U25423 (N_25423,N_25118,N_25071);
and U25424 (N_25424,N_25166,N_25141);
or U25425 (N_25425,N_25114,N_24603);
and U25426 (N_25426,N_24730,N_24669);
and U25427 (N_25427,N_24688,N_24825);
nand U25428 (N_25428,N_24833,N_25024);
or U25429 (N_25429,N_24938,N_24939);
nand U25430 (N_25430,N_24809,N_24605);
or U25431 (N_25431,N_24857,N_25130);
nand U25432 (N_25432,N_24950,N_25058);
xor U25433 (N_25433,N_25045,N_24654);
or U25434 (N_25434,N_24882,N_24735);
nor U25435 (N_25435,N_24964,N_25110);
nand U25436 (N_25436,N_25193,N_25097);
nor U25437 (N_25437,N_24691,N_24849);
nand U25438 (N_25438,N_24610,N_24704);
or U25439 (N_25439,N_25119,N_25031);
xnor U25440 (N_25440,N_24673,N_24854);
or U25441 (N_25441,N_25174,N_24762);
nand U25442 (N_25442,N_24836,N_24991);
nor U25443 (N_25443,N_24875,N_24633);
or U25444 (N_25444,N_25172,N_25101);
xor U25445 (N_25445,N_25184,N_25068);
nor U25446 (N_25446,N_24930,N_24818);
xor U25447 (N_25447,N_24970,N_24794);
nand U25448 (N_25448,N_25067,N_24958);
xnor U25449 (N_25449,N_24607,N_24887);
nor U25450 (N_25450,N_25005,N_25148);
nand U25451 (N_25451,N_24943,N_25095);
nand U25452 (N_25452,N_24601,N_24747);
xor U25453 (N_25453,N_24965,N_24777);
nand U25454 (N_25454,N_24878,N_25065);
nor U25455 (N_25455,N_24884,N_25109);
and U25456 (N_25456,N_25146,N_24845);
or U25457 (N_25457,N_24992,N_24959);
or U25458 (N_25458,N_24785,N_24658);
or U25459 (N_25459,N_25165,N_25018);
nor U25460 (N_25460,N_24961,N_24708);
and U25461 (N_25461,N_24917,N_24816);
nand U25462 (N_25462,N_24668,N_25090);
and U25463 (N_25463,N_24782,N_24746);
nand U25464 (N_25464,N_24971,N_24684);
nor U25465 (N_25465,N_25054,N_25169);
nand U25466 (N_25466,N_24664,N_25098);
and U25467 (N_25467,N_24804,N_24750);
and U25468 (N_25468,N_24940,N_24789);
nand U25469 (N_25469,N_24674,N_24983);
or U25470 (N_25470,N_24676,N_24856);
nor U25471 (N_25471,N_24801,N_25051);
or U25472 (N_25472,N_24657,N_24851);
nand U25473 (N_25473,N_24685,N_24741);
nand U25474 (N_25474,N_24883,N_24795);
and U25475 (N_25475,N_24770,N_24781);
and U25476 (N_25476,N_24814,N_24858);
nor U25477 (N_25477,N_24806,N_24980);
and U25478 (N_25478,N_25181,N_24978);
nand U25479 (N_25479,N_25125,N_25170);
and U25480 (N_25480,N_25026,N_24665);
and U25481 (N_25481,N_25041,N_24713);
nor U25482 (N_25482,N_24901,N_24899);
and U25483 (N_25483,N_25176,N_24860);
nand U25484 (N_25484,N_24952,N_24859);
and U25485 (N_25485,N_25092,N_25088);
and U25486 (N_25486,N_25188,N_25003);
and U25487 (N_25487,N_24835,N_24733);
and U25488 (N_25488,N_24900,N_24670);
xnor U25489 (N_25489,N_24997,N_24867);
or U25490 (N_25490,N_25177,N_24874);
and U25491 (N_25491,N_24680,N_24823);
or U25492 (N_25492,N_24931,N_24926);
and U25493 (N_25493,N_24616,N_24700);
and U25494 (N_25494,N_24682,N_25019);
and U25495 (N_25495,N_25138,N_25080);
or U25496 (N_25496,N_24855,N_24706);
nand U25497 (N_25497,N_25083,N_24621);
or U25498 (N_25498,N_24907,N_24720);
and U25499 (N_25499,N_24844,N_25038);
and U25500 (N_25500,N_25120,N_25020);
xnor U25501 (N_25501,N_24862,N_24984);
xor U25502 (N_25502,N_24818,N_25056);
nand U25503 (N_25503,N_24678,N_25000);
nor U25504 (N_25504,N_25176,N_24697);
and U25505 (N_25505,N_24995,N_24720);
nand U25506 (N_25506,N_24635,N_24917);
nor U25507 (N_25507,N_25017,N_24899);
and U25508 (N_25508,N_24996,N_25121);
nor U25509 (N_25509,N_24968,N_25188);
or U25510 (N_25510,N_25134,N_24833);
xnor U25511 (N_25511,N_24797,N_24695);
or U25512 (N_25512,N_24949,N_25053);
nor U25513 (N_25513,N_25031,N_24628);
and U25514 (N_25514,N_24914,N_24870);
xor U25515 (N_25515,N_24615,N_25106);
xnor U25516 (N_25516,N_24663,N_25020);
nand U25517 (N_25517,N_25197,N_24994);
and U25518 (N_25518,N_24747,N_24706);
nand U25519 (N_25519,N_25198,N_24912);
nand U25520 (N_25520,N_24769,N_24659);
or U25521 (N_25521,N_24707,N_24787);
nor U25522 (N_25522,N_25111,N_24663);
nor U25523 (N_25523,N_25110,N_25043);
and U25524 (N_25524,N_25043,N_25005);
nor U25525 (N_25525,N_25010,N_24886);
and U25526 (N_25526,N_25002,N_25091);
and U25527 (N_25527,N_24687,N_25193);
and U25528 (N_25528,N_24720,N_24847);
or U25529 (N_25529,N_24703,N_24794);
nand U25530 (N_25530,N_24901,N_25153);
nand U25531 (N_25531,N_24814,N_24797);
or U25532 (N_25532,N_25090,N_24750);
xor U25533 (N_25533,N_25197,N_25180);
and U25534 (N_25534,N_24639,N_24852);
and U25535 (N_25535,N_24778,N_24809);
nor U25536 (N_25536,N_24609,N_24708);
xor U25537 (N_25537,N_24787,N_25089);
or U25538 (N_25538,N_25150,N_25194);
xnor U25539 (N_25539,N_25014,N_24977);
and U25540 (N_25540,N_25122,N_25057);
xor U25541 (N_25541,N_25014,N_24943);
xnor U25542 (N_25542,N_24714,N_24634);
and U25543 (N_25543,N_24977,N_25068);
and U25544 (N_25544,N_25121,N_24884);
nand U25545 (N_25545,N_24938,N_24811);
or U25546 (N_25546,N_24604,N_25167);
or U25547 (N_25547,N_25055,N_24686);
and U25548 (N_25548,N_24862,N_25034);
nand U25549 (N_25549,N_24991,N_24907);
nor U25550 (N_25550,N_25197,N_24912);
nor U25551 (N_25551,N_24931,N_25069);
or U25552 (N_25552,N_24808,N_24823);
or U25553 (N_25553,N_24989,N_24923);
nor U25554 (N_25554,N_25069,N_24656);
nand U25555 (N_25555,N_24736,N_25102);
xnor U25556 (N_25556,N_24962,N_24913);
xnor U25557 (N_25557,N_24862,N_24754);
nor U25558 (N_25558,N_25164,N_24740);
or U25559 (N_25559,N_24944,N_24744);
nor U25560 (N_25560,N_24800,N_25076);
nand U25561 (N_25561,N_24963,N_24849);
xnor U25562 (N_25562,N_24619,N_24760);
nand U25563 (N_25563,N_24780,N_25039);
nor U25564 (N_25564,N_24912,N_25167);
nand U25565 (N_25565,N_24984,N_24897);
nand U25566 (N_25566,N_25194,N_24857);
nand U25567 (N_25567,N_24999,N_25033);
or U25568 (N_25568,N_24614,N_25191);
nand U25569 (N_25569,N_24869,N_25194);
nand U25570 (N_25570,N_25161,N_24630);
nand U25571 (N_25571,N_24773,N_24961);
nand U25572 (N_25572,N_25008,N_24606);
nand U25573 (N_25573,N_24661,N_24749);
or U25574 (N_25574,N_24945,N_24839);
nand U25575 (N_25575,N_25123,N_25054);
nand U25576 (N_25576,N_24603,N_24831);
nand U25577 (N_25577,N_25123,N_24929);
nand U25578 (N_25578,N_24914,N_24803);
nand U25579 (N_25579,N_24982,N_24677);
nand U25580 (N_25580,N_24862,N_24969);
and U25581 (N_25581,N_25042,N_24893);
or U25582 (N_25582,N_25088,N_24727);
or U25583 (N_25583,N_25060,N_24883);
or U25584 (N_25584,N_25129,N_24737);
nor U25585 (N_25585,N_25059,N_24834);
nand U25586 (N_25586,N_25181,N_25031);
and U25587 (N_25587,N_24884,N_25197);
nor U25588 (N_25588,N_25131,N_25026);
or U25589 (N_25589,N_25092,N_25127);
nor U25590 (N_25590,N_24662,N_25021);
nor U25591 (N_25591,N_25182,N_25140);
nor U25592 (N_25592,N_25174,N_24814);
and U25593 (N_25593,N_25003,N_24607);
xor U25594 (N_25594,N_24668,N_25071);
and U25595 (N_25595,N_25026,N_24900);
and U25596 (N_25596,N_25195,N_24646);
nand U25597 (N_25597,N_24739,N_24807);
or U25598 (N_25598,N_24771,N_24624);
nand U25599 (N_25599,N_25125,N_25063);
nor U25600 (N_25600,N_24865,N_25148);
and U25601 (N_25601,N_24625,N_24861);
nor U25602 (N_25602,N_25193,N_24819);
xor U25603 (N_25603,N_24680,N_24765);
and U25604 (N_25604,N_24873,N_24829);
or U25605 (N_25605,N_25017,N_25168);
nand U25606 (N_25606,N_24885,N_24782);
nor U25607 (N_25607,N_25033,N_24909);
nor U25608 (N_25608,N_24987,N_25047);
xnor U25609 (N_25609,N_24876,N_25146);
nand U25610 (N_25610,N_24613,N_24922);
and U25611 (N_25611,N_24827,N_25198);
or U25612 (N_25612,N_24907,N_24977);
xor U25613 (N_25613,N_25083,N_24835);
nand U25614 (N_25614,N_24775,N_25007);
and U25615 (N_25615,N_24877,N_24833);
or U25616 (N_25616,N_25026,N_25146);
nand U25617 (N_25617,N_24902,N_24996);
xnor U25618 (N_25618,N_24693,N_25066);
and U25619 (N_25619,N_25064,N_24895);
xnor U25620 (N_25620,N_25158,N_24984);
or U25621 (N_25621,N_25087,N_24990);
and U25622 (N_25622,N_25003,N_24626);
or U25623 (N_25623,N_24710,N_25021);
xnor U25624 (N_25624,N_24904,N_24783);
xor U25625 (N_25625,N_24776,N_24927);
nor U25626 (N_25626,N_24908,N_24928);
nand U25627 (N_25627,N_24845,N_24871);
xnor U25628 (N_25628,N_24923,N_24840);
nand U25629 (N_25629,N_25049,N_24886);
nor U25630 (N_25630,N_24908,N_24914);
nand U25631 (N_25631,N_25196,N_25154);
and U25632 (N_25632,N_25096,N_24662);
nand U25633 (N_25633,N_24897,N_24820);
and U25634 (N_25634,N_25010,N_25064);
nor U25635 (N_25635,N_24990,N_24815);
nand U25636 (N_25636,N_24767,N_25108);
or U25637 (N_25637,N_25146,N_24892);
nor U25638 (N_25638,N_24901,N_24996);
or U25639 (N_25639,N_25188,N_25072);
nor U25640 (N_25640,N_24903,N_25168);
nor U25641 (N_25641,N_25042,N_24791);
and U25642 (N_25642,N_24683,N_24833);
nand U25643 (N_25643,N_24731,N_24876);
and U25644 (N_25644,N_24952,N_24941);
nand U25645 (N_25645,N_24966,N_24684);
or U25646 (N_25646,N_24781,N_24700);
nand U25647 (N_25647,N_25103,N_24699);
and U25648 (N_25648,N_24706,N_24780);
xnor U25649 (N_25649,N_24908,N_24804);
nand U25650 (N_25650,N_24808,N_24801);
or U25651 (N_25651,N_25019,N_24984);
nand U25652 (N_25652,N_24779,N_25189);
nor U25653 (N_25653,N_24686,N_25062);
or U25654 (N_25654,N_24669,N_24934);
and U25655 (N_25655,N_24662,N_24934);
xor U25656 (N_25656,N_24866,N_25036);
and U25657 (N_25657,N_25103,N_24996);
and U25658 (N_25658,N_25028,N_24987);
and U25659 (N_25659,N_25052,N_24947);
nand U25660 (N_25660,N_24730,N_25050);
nor U25661 (N_25661,N_25021,N_25174);
and U25662 (N_25662,N_24742,N_24883);
or U25663 (N_25663,N_24657,N_24866);
nand U25664 (N_25664,N_25123,N_24661);
and U25665 (N_25665,N_25117,N_25064);
nand U25666 (N_25666,N_25090,N_25016);
or U25667 (N_25667,N_24737,N_25052);
nand U25668 (N_25668,N_24896,N_24901);
nor U25669 (N_25669,N_25107,N_24757);
or U25670 (N_25670,N_25000,N_25056);
nor U25671 (N_25671,N_24747,N_24676);
or U25672 (N_25672,N_25104,N_24739);
nand U25673 (N_25673,N_24936,N_24800);
nand U25674 (N_25674,N_25142,N_24819);
or U25675 (N_25675,N_24729,N_24716);
nand U25676 (N_25676,N_24994,N_25182);
or U25677 (N_25677,N_24635,N_24796);
nor U25678 (N_25678,N_25058,N_24851);
nor U25679 (N_25679,N_24701,N_24984);
or U25680 (N_25680,N_24735,N_24983);
and U25681 (N_25681,N_25007,N_24898);
nor U25682 (N_25682,N_25096,N_24706);
and U25683 (N_25683,N_25098,N_25005);
and U25684 (N_25684,N_24972,N_24613);
nor U25685 (N_25685,N_24690,N_25111);
nor U25686 (N_25686,N_24732,N_25145);
nand U25687 (N_25687,N_24951,N_25051);
or U25688 (N_25688,N_25033,N_24980);
nand U25689 (N_25689,N_24787,N_24629);
nor U25690 (N_25690,N_25048,N_24635);
xor U25691 (N_25691,N_24827,N_24748);
xor U25692 (N_25692,N_24690,N_24706);
xnor U25693 (N_25693,N_24650,N_24729);
or U25694 (N_25694,N_24923,N_24716);
nand U25695 (N_25695,N_25015,N_24672);
or U25696 (N_25696,N_24938,N_25154);
and U25697 (N_25697,N_24825,N_25069);
nand U25698 (N_25698,N_25057,N_24870);
or U25699 (N_25699,N_24669,N_25040);
nor U25700 (N_25700,N_24623,N_24768);
xnor U25701 (N_25701,N_24603,N_24962);
or U25702 (N_25702,N_24922,N_24981);
xor U25703 (N_25703,N_24737,N_24706);
nand U25704 (N_25704,N_25049,N_24637);
nand U25705 (N_25705,N_24927,N_24920);
and U25706 (N_25706,N_24806,N_25127);
or U25707 (N_25707,N_24771,N_24721);
or U25708 (N_25708,N_24880,N_24724);
xnor U25709 (N_25709,N_25038,N_24647);
nor U25710 (N_25710,N_24970,N_25098);
and U25711 (N_25711,N_24991,N_25050);
nor U25712 (N_25712,N_24749,N_25083);
xnor U25713 (N_25713,N_24910,N_24887);
and U25714 (N_25714,N_24993,N_24739);
or U25715 (N_25715,N_25026,N_24971);
xnor U25716 (N_25716,N_24723,N_24861);
and U25717 (N_25717,N_24811,N_24723);
or U25718 (N_25718,N_25171,N_25147);
and U25719 (N_25719,N_24705,N_25112);
nor U25720 (N_25720,N_24904,N_25081);
nand U25721 (N_25721,N_24630,N_24844);
and U25722 (N_25722,N_24973,N_24862);
and U25723 (N_25723,N_24673,N_24733);
and U25724 (N_25724,N_24693,N_25126);
and U25725 (N_25725,N_24913,N_24880);
nor U25726 (N_25726,N_24669,N_25034);
nor U25727 (N_25727,N_25127,N_24699);
nor U25728 (N_25728,N_24762,N_24681);
xor U25729 (N_25729,N_25087,N_24620);
and U25730 (N_25730,N_24695,N_24812);
nor U25731 (N_25731,N_25036,N_24647);
nand U25732 (N_25732,N_25048,N_25154);
or U25733 (N_25733,N_24773,N_25034);
nor U25734 (N_25734,N_24621,N_24759);
nor U25735 (N_25735,N_24774,N_24784);
nand U25736 (N_25736,N_24789,N_24846);
and U25737 (N_25737,N_24649,N_24641);
nor U25738 (N_25738,N_25127,N_25028);
and U25739 (N_25739,N_24996,N_25091);
and U25740 (N_25740,N_24992,N_24851);
or U25741 (N_25741,N_24847,N_25035);
xor U25742 (N_25742,N_24657,N_25058);
or U25743 (N_25743,N_24941,N_24693);
nand U25744 (N_25744,N_24819,N_24609);
or U25745 (N_25745,N_25055,N_24926);
or U25746 (N_25746,N_24809,N_25143);
xnor U25747 (N_25747,N_25164,N_25009);
nor U25748 (N_25748,N_24892,N_25001);
or U25749 (N_25749,N_25104,N_25055);
nor U25750 (N_25750,N_24876,N_24649);
nor U25751 (N_25751,N_24916,N_24911);
nor U25752 (N_25752,N_24839,N_24670);
and U25753 (N_25753,N_24605,N_25053);
or U25754 (N_25754,N_24618,N_24676);
nor U25755 (N_25755,N_24821,N_25118);
nor U25756 (N_25756,N_24946,N_25052);
nand U25757 (N_25757,N_25113,N_25137);
or U25758 (N_25758,N_24705,N_24763);
and U25759 (N_25759,N_25092,N_24886);
and U25760 (N_25760,N_25058,N_24611);
or U25761 (N_25761,N_25089,N_24632);
nand U25762 (N_25762,N_24653,N_25180);
or U25763 (N_25763,N_25130,N_25030);
and U25764 (N_25764,N_24657,N_25024);
or U25765 (N_25765,N_24658,N_24601);
and U25766 (N_25766,N_25190,N_25025);
nor U25767 (N_25767,N_24913,N_24614);
nand U25768 (N_25768,N_24614,N_24929);
nand U25769 (N_25769,N_24638,N_24937);
or U25770 (N_25770,N_24691,N_25107);
or U25771 (N_25771,N_24772,N_24697);
and U25772 (N_25772,N_24628,N_24857);
nand U25773 (N_25773,N_24821,N_24680);
xnor U25774 (N_25774,N_25075,N_25042);
nand U25775 (N_25775,N_25184,N_25061);
and U25776 (N_25776,N_24945,N_25007);
nand U25777 (N_25777,N_24872,N_25163);
nor U25778 (N_25778,N_24784,N_25051);
nor U25779 (N_25779,N_24639,N_24739);
nor U25780 (N_25780,N_25063,N_24663);
or U25781 (N_25781,N_24915,N_24781);
and U25782 (N_25782,N_25001,N_24628);
nand U25783 (N_25783,N_24927,N_24950);
nor U25784 (N_25784,N_25082,N_24706);
nand U25785 (N_25785,N_24837,N_25070);
xnor U25786 (N_25786,N_25003,N_25025);
nand U25787 (N_25787,N_24848,N_24976);
xnor U25788 (N_25788,N_24657,N_24629);
nand U25789 (N_25789,N_24894,N_24617);
or U25790 (N_25790,N_24630,N_25108);
and U25791 (N_25791,N_25131,N_24938);
and U25792 (N_25792,N_24640,N_24916);
and U25793 (N_25793,N_25109,N_25124);
nand U25794 (N_25794,N_24829,N_25032);
nor U25795 (N_25795,N_24991,N_24857);
xor U25796 (N_25796,N_25018,N_24790);
and U25797 (N_25797,N_24861,N_24915);
nand U25798 (N_25798,N_24707,N_25060);
or U25799 (N_25799,N_25142,N_24924);
nand U25800 (N_25800,N_25364,N_25635);
and U25801 (N_25801,N_25738,N_25283);
nor U25802 (N_25802,N_25404,N_25717);
nor U25803 (N_25803,N_25634,N_25599);
nor U25804 (N_25804,N_25551,N_25756);
and U25805 (N_25805,N_25236,N_25466);
xor U25806 (N_25806,N_25242,N_25301);
or U25807 (N_25807,N_25358,N_25509);
xnor U25808 (N_25808,N_25694,N_25453);
xor U25809 (N_25809,N_25501,N_25249);
and U25810 (N_25810,N_25472,N_25684);
xnor U25811 (N_25811,N_25674,N_25677);
nor U25812 (N_25812,N_25243,N_25701);
or U25813 (N_25813,N_25467,N_25418);
xor U25814 (N_25814,N_25350,N_25465);
nand U25815 (N_25815,N_25286,N_25444);
or U25816 (N_25816,N_25308,N_25511);
nor U25817 (N_25817,N_25436,N_25517);
and U25818 (N_25818,N_25798,N_25568);
nor U25819 (N_25819,N_25547,N_25700);
and U25820 (N_25820,N_25414,N_25422);
nor U25821 (N_25821,N_25428,N_25312);
nand U25822 (N_25822,N_25720,N_25755);
nand U25823 (N_25823,N_25359,N_25653);
and U25824 (N_25824,N_25267,N_25377);
nor U25825 (N_25825,N_25617,N_25745);
or U25826 (N_25826,N_25485,N_25493);
xnor U25827 (N_25827,N_25697,N_25206);
and U25828 (N_25828,N_25380,N_25619);
nand U25829 (N_25829,N_25222,N_25544);
nor U25830 (N_25830,N_25651,N_25344);
or U25831 (N_25831,N_25354,N_25514);
nor U25832 (N_25832,N_25743,N_25337);
and U25833 (N_25833,N_25785,N_25740);
nor U25834 (N_25834,N_25665,N_25586);
xor U25835 (N_25835,N_25248,N_25282);
nor U25836 (N_25836,N_25250,N_25291);
and U25837 (N_25837,N_25708,N_25468);
or U25838 (N_25838,N_25688,N_25253);
nand U25839 (N_25839,N_25405,N_25706);
nor U25840 (N_25840,N_25481,N_25722);
and U25841 (N_25841,N_25524,N_25461);
and U25842 (N_25842,N_25205,N_25211);
nor U25843 (N_25843,N_25434,N_25378);
nand U25844 (N_25844,N_25754,N_25426);
xor U25845 (N_25845,N_25790,N_25583);
nand U25846 (N_25846,N_25726,N_25556);
nand U25847 (N_25847,N_25505,N_25258);
nor U25848 (N_25848,N_25395,N_25631);
or U25849 (N_25849,N_25503,N_25593);
or U25850 (N_25850,N_25579,N_25229);
nand U25851 (N_25851,N_25686,N_25207);
and U25852 (N_25852,N_25682,N_25399);
or U25853 (N_25853,N_25530,N_25425);
and U25854 (N_25854,N_25273,N_25246);
or U25855 (N_25855,N_25742,N_25478);
and U25856 (N_25856,N_25375,N_25406);
or U25857 (N_25857,N_25462,N_25666);
and U25858 (N_25858,N_25765,N_25690);
and U25859 (N_25859,N_25285,N_25268);
and U25860 (N_25860,N_25794,N_25607);
or U25861 (N_25861,N_25540,N_25214);
or U25862 (N_25862,N_25739,N_25373);
nor U25863 (N_25863,N_25669,N_25681);
or U25864 (N_25864,N_25591,N_25679);
nor U25865 (N_25865,N_25621,N_25241);
xor U25866 (N_25866,N_25314,N_25317);
and U25867 (N_25867,N_25360,N_25353);
nand U25868 (N_25868,N_25624,N_25298);
or U25869 (N_25869,N_25777,N_25332);
nand U25870 (N_25870,N_25367,N_25451);
and U25871 (N_25871,N_25704,N_25259);
or U25872 (N_25872,N_25470,N_25616);
and U25873 (N_25873,N_25459,N_25416);
and U25874 (N_25874,N_25491,N_25334);
nor U25875 (N_25875,N_25333,N_25322);
or U25876 (N_25876,N_25587,N_25512);
or U25877 (N_25877,N_25476,N_25389);
nor U25878 (N_25878,N_25382,N_25786);
xnor U25879 (N_25879,N_25529,N_25490);
and U25880 (N_25880,N_25772,N_25329);
or U25881 (N_25881,N_25254,N_25363);
or U25882 (N_25882,N_25584,N_25369);
or U25883 (N_25883,N_25492,N_25356);
and U25884 (N_25884,N_25637,N_25304);
nand U25885 (N_25885,N_25608,N_25439);
and U25886 (N_25886,N_25237,N_25646);
or U25887 (N_25887,N_25245,N_25753);
or U25888 (N_25888,N_25531,N_25227);
and U25889 (N_25889,N_25603,N_25498);
and U25890 (N_25890,N_25589,N_25230);
nor U25891 (N_25891,N_25252,N_25793);
xor U25892 (N_25892,N_25705,N_25613);
and U25893 (N_25893,N_25394,N_25689);
xnor U25894 (N_25894,N_25600,N_25480);
or U25895 (N_25895,N_25471,N_25667);
xnor U25896 (N_25896,N_25678,N_25327);
and U25897 (N_25897,N_25400,N_25348);
and U25898 (N_25898,N_25733,N_25311);
nor U25899 (N_25899,N_25675,N_25257);
nand U25900 (N_25900,N_25432,N_25219);
or U25901 (N_25901,N_25647,N_25352);
or U25902 (N_25902,N_25645,N_25762);
nor U25903 (N_25903,N_25764,N_25566);
xnor U25904 (N_25904,N_25421,N_25216);
xnor U25905 (N_25905,N_25403,N_25622);
or U25906 (N_25906,N_25374,N_25330);
nand U25907 (N_25907,N_25244,N_25691);
xor U25908 (N_25908,N_25497,N_25397);
and U25909 (N_25909,N_25202,N_25487);
nand U25910 (N_25910,N_25671,N_25567);
xnor U25911 (N_25911,N_25734,N_25393);
or U25912 (N_25912,N_25293,N_25477);
or U25913 (N_25913,N_25661,N_25435);
nand U25914 (N_25914,N_25737,N_25656);
nor U25915 (N_25915,N_25787,N_25758);
nor U25916 (N_25916,N_25309,N_25464);
or U25917 (N_25917,N_25657,N_25396);
nand U25918 (N_25918,N_25446,N_25507);
or U25919 (N_25919,N_25773,N_25528);
nor U25920 (N_25920,N_25592,N_25695);
nor U25921 (N_25921,N_25429,N_25554);
nand U25922 (N_25922,N_25424,N_25506);
nor U25923 (N_25923,N_25571,N_25536);
nor U25924 (N_25924,N_25287,N_25610);
nor U25925 (N_25925,N_25574,N_25225);
and U25926 (N_25926,N_25539,N_25663);
nor U25927 (N_25927,N_25714,N_25636);
nand U25928 (N_25928,N_25321,N_25718);
nor U25929 (N_25929,N_25447,N_25313);
xor U25930 (N_25930,N_25456,N_25233);
and U25931 (N_25931,N_25220,N_25278);
and U25932 (N_25932,N_25792,N_25319);
or U25933 (N_25933,N_25379,N_25759);
nand U25934 (N_25934,N_25711,N_25719);
xor U25935 (N_25935,N_25747,N_25280);
or U25936 (N_25936,N_25768,N_25372);
nor U25937 (N_25937,N_25519,N_25209);
and U25938 (N_25938,N_25411,N_25376);
nor U25939 (N_25939,N_25288,N_25226);
or U25940 (N_25940,N_25510,N_25668);
nand U25941 (N_25941,N_25549,N_25296);
xor U25942 (N_25942,N_25208,N_25781);
nor U25943 (N_25943,N_25455,N_25274);
nand U25944 (N_25944,N_25541,N_25799);
nor U25945 (N_25945,N_25228,N_25552);
and U25946 (N_25946,N_25500,N_25351);
and U25947 (N_25947,N_25407,N_25565);
and U25948 (N_25948,N_25215,N_25537);
or U25949 (N_25949,N_25221,N_25774);
nor U25950 (N_25950,N_25315,N_25670);
and U25951 (N_25951,N_25408,N_25295);
nand U25952 (N_25952,N_25290,N_25335);
or U25953 (N_25953,N_25345,N_25204);
xnor U25954 (N_25954,N_25449,N_25255);
and U25955 (N_25955,N_25732,N_25299);
and U25956 (N_25956,N_25496,N_25275);
and U25957 (N_25957,N_25307,N_25448);
and U25958 (N_25958,N_25757,N_25326);
nand U25959 (N_25959,N_25516,N_25323);
and U25960 (N_25960,N_25489,N_25385);
nand U25961 (N_25961,N_25623,N_25265);
nor U25962 (N_25962,N_25638,N_25523);
nor U25963 (N_25963,N_25650,N_25475);
nand U25964 (N_25964,N_25442,N_25796);
and U25965 (N_25965,N_25402,N_25751);
and U25966 (N_25966,N_25458,N_25595);
and U25967 (N_25967,N_25572,N_25218);
and U25968 (N_25968,N_25618,N_25680);
nand U25969 (N_25969,N_25558,N_25521);
or U25970 (N_25970,N_25370,N_25398);
and U25971 (N_25971,N_25388,N_25783);
or U25972 (N_25972,N_25716,N_25673);
nand U25973 (N_25973,N_25658,N_25576);
or U25974 (N_25974,N_25342,N_25629);
and U25975 (N_25975,N_25550,N_25557);
nor U25976 (N_25976,N_25266,N_25585);
and U25977 (N_25977,N_25609,N_25562);
and U25978 (N_25978,N_25769,N_25349);
and U25979 (N_25979,N_25494,N_25409);
or U25980 (N_25980,N_25692,N_25683);
xor U25981 (N_25981,N_25766,N_25341);
and U25982 (N_25982,N_25502,N_25534);
and U25983 (N_25983,N_25605,N_25748);
or U25984 (N_25984,N_25495,N_25235);
nor U25985 (N_25985,N_25224,N_25284);
nor U25986 (N_25986,N_25546,N_25553);
and U25987 (N_25987,N_25580,N_25386);
and U25988 (N_25988,N_25325,N_25361);
and U25989 (N_25989,N_25542,N_25427);
xnor U25990 (N_25990,N_25563,N_25672);
or U25991 (N_25991,N_25212,N_25597);
nand U25992 (N_25992,N_25729,N_25644);
xnor U25993 (N_25993,N_25770,N_25318);
or U25994 (N_25994,N_25518,N_25577);
nor U25995 (N_25995,N_25336,N_25611);
or U25996 (N_25996,N_25279,N_25417);
xor U25997 (N_25997,N_25676,N_25788);
or U25998 (N_25998,N_25401,N_25355);
nand U25999 (N_25999,N_25483,N_25338);
xnor U26000 (N_26000,N_25201,N_25231);
xnor U26001 (N_26001,N_25693,N_25789);
or U26002 (N_26002,N_25240,N_25302);
nand U26003 (N_26003,N_25620,N_25744);
nand U26004 (N_26004,N_25515,N_25707);
or U26005 (N_26005,N_25604,N_25276);
or U26006 (N_26006,N_25390,N_25431);
xnor U26007 (N_26007,N_25710,N_25270);
nor U26008 (N_26008,N_25251,N_25520);
nand U26009 (N_26009,N_25628,N_25685);
nor U26010 (N_26010,N_25612,N_25564);
or U26011 (N_26011,N_25383,N_25441);
nor U26012 (N_26012,N_25440,N_25731);
or U26013 (N_26013,N_25569,N_25649);
nor U26014 (N_26014,N_25594,N_25239);
nand U26015 (N_26015,N_25713,N_25535);
or U26016 (N_26016,N_25721,N_25749);
nor U26017 (N_26017,N_25238,N_25533);
nor U26018 (N_26018,N_25632,N_25699);
or U26019 (N_26019,N_25504,N_25633);
or U26020 (N_26020,N_25615,N_25423);
nor U26021 (N_26021,N_25445,N_25760);
xnor U26022 (N_26022,N_25545,N_25642);
nand U26023 (N_26023,N_25387,N_25771);
and U26024 (N_26024,N_25570,N_25626);
and U26025 (N_26025,N_25588,N_25532);
nand U26026 (N_26026,N_25601,N_25210);
nand U26027 (N_26027,N_25247,N_25303);
or U26028 (N_26028,N_25277,N_25728);
or U26029 (N_26029,N_25525,N_25602);
nor U26030 (N_26030,N_25508,N_25640);
nand U26031 (N_26031,N_25606,N_25526);
nand U26032 (N_26032,N_25648,N_25347);
and U26033 (N_26033,N_25412,N_25371);
nand U26034 (N_26034,N_25264,N_25746);
and U26035 (N_26035,N_25346,N_25730);
and U26036 (N_26036,N_25763,N_25260);
and U26037 (N_26037,N_25778,N_25659);
nand U26038 (N_26038,N_25482,N_25262);
or U26039 (N_26039,N_25614,N_25784);
or U26040 (N_26040,N_25761,N_25437);
or U26041 (N_26041,N_25513,N_25232);
or U26042 (N_26042,N_25430,N_25297);
or U26043 (N_26043,N_25488,N_25779);
nor U26044 (N_26044,N_25573,N_25339);
nand U26045 (N_26045,N_25664,N_25797);
nand U26046 (N_26046,N_25450,N_25538);
nand U26047 (N_26047,N_25200,N_25340);
and U26048 (N_26048,N_25598,N_25527);
or U26049 (N_26049,N_25310,N_25419);
nand U26050 (N_26050,N_25271,N_25791);
and U26051 (N_26051,N_25559,N_25474);
or U26052 (N_26052,N_25256,N_25343);
or U26053 (N_26053,N_25357,N_25292);
nor U26054 (N_26054,N_25630,N_25365);
nand U26055 (N_26055,N_25715,N_25328);
nand U26056 (N_26056,N_25627,N_25484);
and U26057 (N_26057,N_25281,N_25780);
and U26058 (N_26058,N_25294,N_25223);
nor U26059 (N_26059,N_25331,N_25457);
and U26060 (N_26060,N_25454,N_25641);
nor U26061 (N_26061,N_25499,N_25782);
nor U26062 (N_26062,N_25479,N_25723);
or U26063 (N_26063,N_25702,N_25581);
nand U26064 (N_26064,N_25703,N_25463);
or U26065 (N_26065,N_25776,N_25625);
or U26066 (N_26066,N_25555,N_25696);
xnor U26067 (N_26067,N_25767,N_25655);
nor U26068 (N_26068,N_25443,N_25560);
or U26069 (N_26069,N_25415,N_25639);
and U26070 (N_26070,N_25543,N_25234);
nor U26071 (N_26071,N_25366,N_25561);
nand U26072 (N_26072,N_25420,N_25724);
or U26073 (N_26073,N_25709,N_25750);
or U26074 (N_26074,N_25460,N_25652);
nor U26075 (N_26075,N_25272,N_25741);
xnor U26076 (N_26076,N_25433,N_25410);
and U26077 (N_26077,N_25300,N_25596);
and U26078 (N_26078,N_25213,N_25316);
nand U26079 (N_26079,N_25662,N_25469);
and U26080 (N_26080,N_25712,N_25473);
and U26081 (N_26081,N_25775,N_25548);
nand U26082 (N_26082,N_25203,N_25306);
xnor U26083 (N_26083,N_25486,N_25660);
or U26084 (N_26084,N_25263,N_25217);
nor U26085 (N_26085,N_25269,N_25725);
xor U26086 (N_26086,N_25736,N_25522);
nand U26087 (N_26087,N_25643,N_25582);
or U26088 (N_26088,N_25687,N_25654);
nor U26089 (N_26089,N_25381,N_25261);
and U26090 (N_26090,N_25413,N_25795);
nor U26091 (N_26091,N_25698,N_25362);
and U26092 (N_26092,N_25305,N_25735);
or U26093 (N_26093,N_25324,N_25384);
nor U26094 (N_26094,N_25575,N_25727);
nand U26095 (N_26095,N_25391,N_25590);
or U26096 (N_26096,N_25438,N_25320);
and U26097 (N_26097,N_25752,N_25578);
nor U26098 (N_26098,N_25368,N_25289);
nor U26099 (N_26099,N_25452,N_25392);
nand U26100 (N_26100,N_25555,N_25212);
nor U26101 (N_26101,N_25456,N_25272);
nor U26102 (N_26102,N_25675,N_25632);
xor U26103 (N_26103,N_25796,N_25230);
or U26104 (N_26104,N_25333,N_25324);
and U26105 (N_26105,N_25708,N_25234);
and U26106 (N_26106,N_25569,N_25321);
nand U26107 (N_26107,N_25518,N_25702);
and U26108 (N_26108,N_25365,N_25206);
nor U26109 (N_26109,N_25575,N_25203);
nand U26110 (N_26110,N_25532,N_25778);
or U26111 (N_26111,N_25258,N_25500);
nor U26112 (N_26112,N_25665,N_25678);
or U26113 (N_26113,N_25303,N_25588);
nand U26114 (N_26114,N_25431,N_25609);
xor U26115 (N_26115,N_25529,N_25624);
or U26116 (N_26116,N_25217,N_25592);
and U26117 (N_26117,N_25480,N_25499);
or U26118 (N_26118,N_25234,N_25304);
and U26119 (N_26119,N_25240,N_25371);
nand U26120 (N_26120,N_25463,N_25533);
or U26121 (N_26121,N_25223,N_25210);
nor U26122 (N_26122,N_25327,N_25495);
or U26123 (N_26123,N_25779,N_25448);
nand U26124 (N_26124,N_25730,N_25589);
nor U26125 (N_26125,N_25723,N_25615);
nand U26126 (N_26126,N_25475,N_25618);
nor U26127 (N_26127,N_25307,N_25625);
and U26128 (N_26128,N_25548,N_25218);
or U26129 (N_26129,N_25216,N_25325);
nor U26130 (N_26130,N_25749,N_25292);
nor U26131 (N_26131,N_25609,N_25423);
nor U26132 (N_26132,N_25227,N_25274);
and U26133 (N_26133,N_25521,N_25689);
or U26134 (N_26134,N_25330,N_25472);
or U26135 (N_26135,N_25378,N_25683);
nor U26136 (N_26136,N_25366,N_25698);
and U26137 (N_26137,N_25546,N_25783);
and U26138 (N_26138,N_25355,N_25369);
nor U26139 (N_26139,N_25760,N_25345);
nor U26140 (N_26140,N_25638,N_25354);
nor U26141 (N_26141,N_25460,N_25654);
or U26142 (N_26142,N_25398,N_25733);
and U26143 (N_26143,N_25417,N_25745);
and U26144 (N_26144,N_25251,N_25656);
or U26145 (N_26145,N_25657,N_25329);
xnor U26146 (N_26146,N_25683,N_25327);
nor U26147 (N_26147,N_25249,N_25326);
and U26148 (N_26148,N_25651,N_25675);
nand U26149 (N_26149,N_25457,N_25228);
xnor U26150 (N_26150,N_25283,N_25470);
nor U26151 (N_26151,N_25272,N_25743);
or U26152 (N_26152,N_25409,N_25253);
and U26153 (N_26153,N_25780,N_25310);
nor U26154 (N_26154,N_25558,N_25440);
or U26155 (N_26155,N_25600,N_25388);
nand U26156 (N_26156,N_25322,N_25760);
and U26157 (N_26157,N_25749,N_25338);
or U26158 (N_26158,N_25442,N_25477);
nor U26159 (N_26159,N_25257,N_25281);
xor U26160 (N_26160,N_25691,N_25599);
or U26161 (N_26161,N_25551,N_25436);
or U26162 (N_26162,N_25532,N_25469);
or U26163 (N_26163,N_25636,N_25454);
and U26164 (N_26164,N_25343,N_25489);
nand U26165 (N_26165,N_25792,N_25762);
nor U26166 (N_26166,N_25501,N_25422);
xnor U26167 (N_26167,N_25667,N_25771);
xor U26168 (N_26168,N_25440,N_25216);
or U26169 (N_26169,N_25618,N_25721);
and U26170 (N_26170,N_25607,N_25421);
xor U26171 (N_26171,N_25325,N_25656);
or U26172 (N_26172,N_25512,N_25583);
xnor U26173 (N_26173,N_25376,N_25666);
and U26174 (N_26174,N_25371,N_25702);
nor U26175 (N_26175,N_25491,N_25764);
or U26176 (N_26176,N_25448,N_25432);
nand U26177 (N_26177,N_25480,N_25529);
and U26178 (N_26178,N_25389,N_25400);
nand U26179 (N_26179,N_25322,N_25628);
nand U26180 (N_26180,N_25405,N_25266);
nor U26181 (N_26181,N_25332,N_25386);
and U26182 (N_26182,N_25589,N_25786);
and U26183 (N_26183,N_25235,N_25216);
nor U26184 (N_26184,N_25349,N_25320);
xnor U26185 (N_26185,N_25736,N_25677);
nor U26186 (N_26186,N_25744,N_25341);
xor U26187 (N_26187,N_25756,N_25407);
nand U26188 (N_26188,N_25764,N_25692);
or U26189 (N_26189,N_25795,N_25703);
and U26190 (N_26190,N_25226,N_25675);
and U26191 (N_26191,N_25586,N_25206);
nand U26192 (N_26192,N_25585,N_25791);
or U26193 (N_26193,N_25269,N_25655);
and U26194 (N_26194,N_25276,N_25698);
and U26195 (N_26195,N_25565,N_25270);
and U26196 (N_26196,N_25380,N_25562);
nor U26197 (N_26197,N_25760,N_25455);
nor U26198 (N_26198,N_25360,N_25214);
xnor U26199 (N_26199,N_25593,N_25308);
nand U26200 (N_26200,N_25223,N_25306);
and U26201 (N_26201,N_25369,N_25294);
xnor U26202 (N_26202,N_25479,N_25468);
or U26203 (N_26203,N_25376,N_25724);
nand U26204 (N_26204,N_25367,N_25274);
xor U26205 (N_26205,N_25631,N_25576);
nor U26206 (N_26206,N_25796,N_25621);
and U26207 (N_26207,N_25409,N_25250);
and U26208 (N_26208,N_25332,N_25768);
xnor U26209 (N_26209,N_25760,N_25398);
or U26210 (N_26210,N_25455,N_25221);
xnor U26211 (N_26211,N_25503,N_25385);
and U26212 (N_26212,N_25355,N_25256);
nand U26213 (N_26213,N_25435,N_25756);
nand U26214 (N_26214,N_25356,N_25343);
and U26215 (N_26215,N_25591,N_25347);
and U26216 (N_26216,N_25786,N_25620);
nor U26217 (N_26217,N_25296,N_25443);
and U26218 (N_26218,N_25383,N_25235);
or U26219 (N_26219,N_25409,N_25652);
or U26220 (N_26220,N_25452,N_25635);
and U26221 (N_26221,N_25727,N_25540);
or U26222 (N_26222,N_25437,N_25309);
or U26223 (N_26223,N_25761,N_25528);
nor U26224 (N_26224,N_25414,N_25434);
and U26225 (N_26225,N_25434,N_25639);
or U26226 (N_26226,N_25642,N_25661);
or U26227 (N_26227,N_25401,N_25624);
nand U26228 (N_26228,N_25535,N_25404);
nand U26229 (N_26229,N_25754,N_25652);
or U26230 (N_26230,N_25379,N_25451);
nor U26231 (N_26231,N_25616,N_25666);
or U26232 (N_26232,N_25599,N_25230);
or U26233 (N_26233,N_25767,N_25627);
xor U26234 (N_26234,N_25591,N_25222);
and U26235 (N_26235,N_25442,N_25480);
nand U26236 (N_26236,N_25552,N_25376);
and U26237 (N_26237,N_25693,N_25484);
xor U26238 (N_26238,N_25703,N_25698);
and U26239 (N_26239,N_25610,N_25575);
xor U26240 (N_26240,N_25764,N_25703);
nand U26241 (N_26241,N_25520,N_25586);
and U26242 (N_26242,N_25622,N_25531);
nor U26243 (N_26243,N_25459,N_25483);
nand U26244 (N_26244,N_25220,N_25280);
xnor U26245 (N_26245,N_25464,N_25322);
or U26246 (N_26246,N_25278,N_25638);
nand U26247 (N_26247,N_25321,N_25211);
and U26248 (N_26248,N_25662,N_25722);
nand U26249 (N_26249,N_25555,N_25483);
or U26250 (N_26250,N_25488,N_25697);
nor U26251 (N_26251,N_25345,N_25785);
xor U26252 (N_26252,N_25294,N_25316);
or U26253 (N_26253,N_25216,N_25654);
and U26254 (N_26254,N_25251,N_25548);
or U26255 (N_26255,N_25726,N_25445);
nor U26256 (N_26256,N_25464,N_25225);
and U26257 (N_26257,N_25589,N_25385);
or U26258 (N_26258,N_25343,N_25706);
and U26259 (N_26259,N_25541,N_25447);
nor U26260 (N_26260,N_25442,N_25512);
or U26261 (N_26261,N_25439,N_25473);
and U26262 (N_26262,N_25383,N_25683);
and U26263 (N_26263,N_25248,N_25614);
nand U26264 (N_26264,N_25306,N_25248);
nor U26265 (N_26265,N_25519,N_25708);
nor U26266 (N_26266,N_25280,N_25766);
nand U26267 (N_26267,N_25615,N_25202);
nor U26268 (N_26268,N_25509,N_25420);
or U26269 (N_26269,N_25313,N_25294);
or U26270 (N_26270,N_25373,N_25709);
nor U26271 (N_26271,N_25607,N_25666);
or U26272 (N_26272,N_25658,N_25760);
or U26273 (N_26273,N_25464,N_25289);
nand U26274 (N_26274,N_25455,N_25672);
or U26275 (N_26275,N_25603,N_25255);
or U26276 (N_26276,N_25536,N_25341);
nor U26277 (N_26277,N_25243,N_25798);
nand U26278 (N_26278,N_25457,N_25436);
or U26279 (N_26279,N_25374,N_25600);
or U26280 (N_26280,N_25383,N_25209);
and U26281 (N_26281,N_25412,N_25372);
xor U26282 (N_26282,N_25368,N_25317);
nand U26283 (N_26283,N_25277,N_25672);
nor U26284 (N_26284,N_25501,N_25234);
nor U26285 (N_26285,N_25514,N_25586);
and U26286 (N_26286,N_25669,N_25734);
nor U26287 (N_26287,N_25771,N_25654);
or U26288 (N_26288,N_25387,N_25577);
or U26289 (N_26289,N_25557,N_25370);
or U26290 (N_26290,N_25556,N_25434);
or U26291 (N_26291,N_25227,N_25705);
and U26292 (N_26292,N_25411,N_25204);
xor U26293 (N_26293,N_25743,N_25591);
or U26294 (N_26294,N_25511,N_25316);
and U26295 (N_26295,N_25232,N_25372);
xnor U26296 (N_26296,N_25687,N_25518);
or U26297 (N_26297,N_25458,N_25759);
nor U26298 (N_26298,N_25530,N_25614);
or U26299 (N_26299,N_25793,N_25429);
or U26300 (N_26300,N_25270,N_25454);
nand U26301 (N_26301,N_25342,N_25533);
nand U26302 (N_26302,N_25265,N_25292);
nand U26303 (N_26303,N_25630,N_25728);
nand U26304 (N_26304,N_25603,N_25300);
nand U26305 (N_26305,N_25727,N_25651);
nand U26306 (N_26306,N_25658,N_25593);
nor U26307 (N_26307,N_25557,N_25232);
or U26308 (N_26308,N_25597,N_25750);
nor U26309 (N_26309,N_25221,N_25699);
xnor U26310 (N_26310,N_25696,N_25708);
nor U26311 (N_26311,N_25557,N_25349);
or U26312 (N_26312,N_25410,N_25723);
nand U26313 (N_26313,N_25288,N_25260);
nand U26314 (N_26314,N_25652,N_25217);
and U26315 (N_26315,N_25495,N_25278);
nor U26316 (N_26316,N_25695,N_25769);
xnor U26317 (N_26317,N_25329,N_25599);
nand U26318 (N_26318,N_25443,N_25576);
and U26319 (N_26319,N_25450,N_25673);
or U26320 (N_26320,N_25727,N_25290);
nand U26321 (N_26321,N_25486,N_25460);
nand U26322 (N_26322,N_25208,N_25642);
nand U26323 (N_26323,N_25376,N_25696);
nor U26324 (N_26324,N_25636,N_25717);
or U26325 (N_26325,N_25448,N_25395);
or U26326 (N_26326,N_25284,N_25376);
and U26327 (N_26327,N_25311,N_25675);
or U26328 (N_26328,N_25676,N_25339);
or U26329 (N_26329,N_25351,N_25637);
and U26330 (N_26330,N_25732,N_25344);
and U26331 (N_26331,N_25310,N_25545);
and U26332 (N_26332,N_25267,N_25480);
nor U26333 (N_26333,N_25644,N_25585);
nand U26334 (N_26334,N_25442,N_25532);
and U26335 (N_26335,N_25752,N_25793);
nor U26336 (N_26336,N_25799,N_25226);
nor U26337 (N_26337,N_25326,N_25296);
nor U26338 (N_26338,N_25630,N_25423);
nand U26339 (N_26339,N_25338,N_25401);
or U26340 (N_26340,N_25540,N_25737);
nand U26341 (N_26341,N_25798,N_25796);
nand U26342 (N_26342,N_25787,N_25319);
and U26343 (N_26343,N_25739,N_25276);
nand U26344 (N_26344,N_25663,N_25442);
xor U26345 (N_26345,N_25330,N_25532);
and U26346 (N_26346,N_25734,N_25238);
nand U26347 (N_26347,N_25299,N_25328);
nand U26348 (N_26348,N_25701,N_25347);
nand U26349 (N_26349,N_25792,N_25597);
xor U26350 (N_26350,N_25568,N_25776);
or U26351 (N_26351,N_25425,N_25402);
nor U26352 (N_26352,N_25607,N_25791);
nor U26353 (N_26353,N_25357,N_25488);
nand U26354 (N_26354,N_25649,N_25257);
or U26355 (N_26355,N_25713,N_25573);
nand U26356 (N_26356,N_25566,N_25433);
nor U26357 (N_26357,N_25248,N_25603);
or U26358 (N_26358,N_25239,N_25489);
nand U26359 (N_26359,N_25781,N_25726);
or U26360 (N_26360,N_25716,N_25579);
nand U26361 (N_26361,N_25593,N_25638);
or U26362 (N_26362,N_25698,N_25682);
xnor U26363 (N_26363,N_25492,N_25330);
nor U26364 (N_26364,N_25226,N_25394);
xnor U26365 (N_26365,N_25452,N_25742);
nor U26366 (N_26366,N_25300,N_25385);
and U26367 (N_26367,N_25523,N_25731);
nand U26368 (N_26368,N_25795,N_25622);
xnor U26369 (N_26369,N_25377,N_25512);
xor U26370 (N_26370,N_25737,N_25352);
nor U26371 (N_26371,N_25336,N_25371);
nand U26372 (N_26372,N_25208,N_25617);
and U26373 (N_26373,N_25740,N_25574);
nor U26374 (N_26374,N_25659,N_25477);
nor U26375 (N_26375,N_25318,N_25618);
or U26376 (N_26376,N_25781,N_25319);
and U26377 (N_26377,N_25601,N_25385);
nor U26378 (N_26378,N_25542,N_25405);
and U26379 (N_26379,N_25783,N_25481);
and U26380 (N_26380,N_25360,N_25403);
and U26381 (N_26381,N_25755,N_25665);
or U26382 (N_26382,N_25600,N_25517);
nor U26383 (N_26383,N_25282,N_25441);
nand U26384 (N_26384,N_25299,N_25441);
and U26385 (N_26385,N_25759,N_25563);
xnor U26386 (N_26386,N_25332,N_25211);
xor U26387 (N_26387,N_25678,N_25322);
and U26388 (N_26388,N_25627,N_25647);
or U26389 (N_26389,N_25239,N_25609);
nor U26390 (N_26390,N_25522,N_25255);
nor U26391 (N_26391,N_25524,N_25255);
nand U26392 (N_26392,N_25562,N_25646);
and U26393 (N_26393,N_25782,N_25715);
and U26394 (N_26394,N_25530,N_25605);
and U26395 (N_26395,N_25748,N_25434);
or U26396 (N_26396,N_25252,N_25662);
nand U26397 (N_26397,N_25635,N_25292);
xnor U26398 (N_26398,N_25731,N_25517);
nand U26399 (N_26399,N_25688,N_25240);
nor U26400 (N_26400,N_26299,N_25961);
or U26401 (N_26401,N_25886,N_26366);
nand U26402 (N_26402,N_26039,N_26030);
nor U26403 (N_26403,N_26390,N_26160);
and U26404 (N_26404,N_25848,N_25952);
or U26405 (N_26405,N_26158,N_26290);
nor U26406 (N_26406,N_26057,N_26395);
nor U26407 (N_26407,N_26074,N_26284);
nor U26408 (N_26408,N_26133,N_26287);
xor U26409 (N_26409,N_26154,N_26337);
or U26410 (N_26410,N_26372,N_26345);
nor U26411 (N_26411,N_26286,N_26075);
nand U26412 (N_26412,N_26099,N_25887);
or U26413 (N_26413,N_25822,N_25833);
nand U26414 (N_26414,N_26013,N_25973);
or U26415 (N_26415,N_26378,N_25812);
and U26416 (N_26416,N_26262,N_25817);
nand U26417 (N_26417,N_26233,N_26006);
nand U26418 (N_26418,N_26203,N_25948);
or U26419 (N_26419,N_26276,N_26321);
or U26420 (N_26420,N_26219,N_26236);
nor U26421 (N_26421,N_26015,N_26305);
and U26422 (N_26422,N_26361,N_26298);
xor U26423 (N_26423,N_25946,N_26359);
nor U26424 (N_26424,N_26307,N_26289);
or U26425 (N_26425,N_26352,N_26109);
and U26426 (N_26426,N_25939,N_26318);
and U26427 (N_26427,N_25809,N_26020);
nand U26428 (N_26428,N_26082,N_26027);
nor U26429 (N_26429,N_26253,N_26172);
nand U26430 (N_26430,N_25991,N_26089);
or U26431 (N_26431,N_26358,N_26189);
nor U26432 (N_26432,N_26312,N_25815);
and U26433 (N_26433,N_25898,N_26205);
or U26434 (N_26434,N_25901,N_26269);
nor U26435 (N_26435,N_25857,N_25861);
and U26436 (N_26436,N_25888,N_26068);
xnor U26437 (N_26437,N_25892,N_26041);
nand U26438 (N_26438,N_25947,N_26391);
nor U26439 (N_26439,N_26139,N_25836);
nor U26440 (N_26440,N_26384,N_26070);
or U26441 (N_26441,N_26187,N_26315);
and U26442 (N_26442,N_26373,N_26334);
nor U26443 (N_26443,N_26363,N_26153);
and U26444 (N_26444,N_26227,N_26155);
and U26445 (N_26445,N_26196,N_26170);
nor U26446 (N_26446,N_26338,N_26224);
and U26447 (N_26447,N_25823,N_25907);
or U26448 (N_26448,N_26360,N_25934);
nor U26449 (N_26449,N_25805,N_25839);
and U26450 (N_26450,N_26377,N_25889);
nand U26451 (N_26451,N_25849,N_26145);
nor U26452 (N_26452,N_25858,N_25832);
and U26453 (N_26453,N_26060,N_25814);
or U26454 (N_26454,N_26392,N_26137);
or U26455 (N_26455,N_26353,N_25843);
nor U26456 (N_26456,N_26232,N_26190);
nand U26457 (N_26457,N_26052,N_26201);
xnor U26458 (N_26458,N_25962,N_26072);
and U26459 (N_26459,N_25916,N_26314);
and U26460 (N_26460,N_26215,N_25903);
nand U26461 (N_26461,N_26168,N_25957);
nand U26462 (N_26462,N_26009,N_26240);
nor U26463 (N_26463,N_26382,N_26093);
nand U26464 (N_26464,N_26291,N_26288);
nand U26465 (N_26465,N_25928,N_25841);
and U26466 (N_26466,N_26239,N_26258);
nor U26467 (N_26467,N_26230,N_25831);
nand U26468 (N_26468,N_26306,N_26293);
nand U26469 (N_26469,N_25895,N_26029);
and U26470 (N_26470,N_26113,N_26004);
nand U26471 (N_26471,N_25804,N_26136);
xnor U26472 (N_26472,N_26025,N_25983);
or U26473 (N_26473,N_25874,N_26121);
xnor U26474 (N_26474,N_25918,N_26256);
nor U26475 (N_26475,N_25975,N_26396);
and U26476 (N_26476,N_25913,N_26161);
and U26477 (N_26477,N_26126,N_25820);
nand U26478 (N_26478,N_26175,N_26058);
or U26479 (N_26479,N_26207,N_26105);
nand U26480 (N_26480,N_26177,N_25846);
nor U26481 (N_26481,N_26016,N_25922);
nor U26482 (N_26482,N_26330,N_26194);
nor U26483 (N_26483,N_26134,N_26092);
or U26484 (N_26484,N_26270,N_25968);
xor U26485 (N_26485,N_26302,N_26008);
nand U26486 (N_26486,N_26340,N_26179);
or U26487 (N_26487,N_26255,N_26220);
and U26488 (N_26488,N_26387,N_26350);
or U26489 (N_26489,N_26007,N_25924);
nor U26490 (N_26490,N_26103,N_26244);
nand U26491 (N_26491,N_26341,N_25837);
nand U26492 (N_26492,N_25927,N_25915);
and U26493 (N_26493,N_26308,N_26188);
or U26494 (N_26494,N_26087,N_25875);
xor U26495 (N_26495,N_25908,N_25802);
nor U26496 (N_26496,N_26148,N_26144);
nand U26497 (N_26497,N_26200,N_25919);
nor U26498 (N_26498,N_26296,N_25929);
nand U26499 (N_26499,N_25803,N_26368);
xor U26500 (N_26500,N_26003,N_25932);
or U26501 (N_26501,N_26046,N_26128);
and U26502 (N_26502,N_26049,N_25982);
and U26503 (N_26503,N_26026,N_25865);
nand U26504 (N_26504,N_26309,N_25876);
nand U26505 (N_26505,N_25828,N_26294);
or U26506 (N_26506,N_26333,N_26024);
and U26507 (N_26507,N_25980,N_26169);
or U26508 (N_26508,N_26226,N_26110);
nor U26509 (N_26509,N_25897,N_25869);
nand U26510 (N_26510,N_26117,N_25830);
nand U26511 (N_26511,N_26346,N_26282);
nand U26512 (N_26512,N_26295,N_26059);
xor U26513 (N_26513,N_25998,N_25992);
nor U26514 (N_26514,N_25920,N_26329);
and U26515 (N_26515,N_25891,N_26062);
or U26516 (N_26516,N_25976,N_25978);
and U26517 (N_26517,N_26266,N_25979);
xnor U26518 (N_26518,N_26159,N_25867);
xor U26519 (N_26519,N_26115,N_26311);
or U26520 (N_26520,N_26053,N_25995);
and U26521 (N_26521,N_26037,N_26260);
nand U26522 (N_26522,N_26047,N_26186);
and U26523 (N_26523,N_25813,N_26019);
nor U26524 (N_26524,N_26209,N_25999);
nand U26525 (N_26525,N_26332,N_25956);
nand U26526 (N_26526,N_26324,N_26356);
nand U26527 (N_26527,N_25900,N_25873);
or U26528 (N_26528,N_25997,N_26193);
or U26529 (N_26529,N_26124,N_26261);
or U26530 (N_26530,N_26038,N_26385);
nand U26531 (N_26531,N_26241,N_25994);
or U26532 (N_26532,N_26225,N_25800);
nor U26533 (N_26533,N_26118,N_26376);
and U26534 (N_26534,N_26279,N_26149);
xnor U26535 (N_26535,N_25967,N_25941);
xnor U26536 (N_26536,N_26218,N_25808);
nand U26537 (N_26537,N_26238,N_25878);
and U26538 (N_26538,N_26357,N_25989);
nand U26539 (N_26539,N_26393,N_25827);
xor U26540 (N_26540,N_26073,N_26151);
xnor U26541 (N_26541,N_26397,N_26192);
and U26542 (N_26542,N_26135,N_25951);
and U26543 (N_26543,N_26214,N_25866);
and U26544 (N_26544,N_26132,N_26274);
nor U26545 (N_26545,N_26348,N_25872);
nor U26546 (N_26546,N_26349,N_26303);
nand U26547 (N_26547,N_26246,N_26183);
or U26548 (N_26548,N_26374,N_25883);
and U26549 (N_26549,N_25852,N_26223);
or U26550 (N_26550,N_26138,N_25818);
or U26551 (N_26551,N_26032,N_25933);
and U26552 (N_26552,N_25993,N_25955);
xnor U26553 (N_26553,N_26066,N_26129);
and U26554 (N_26554,N_26206,N_26213);
and U26555 (N_26555,N_25851,N_26166);
xnor U26556 (N_26556,N_26267,N_26304);
nand U26557 (N_26557,N_26095,N_26141);
nor U26558 (N_26558,N_25996,N_26000);
or U26559 (N_26559,N_26331,N_25940);
xnor U26560 (N_26560,N_26280,N_25885);
nor U26561 (N_26561,N_26090,N_25925);
nand U26562 (N_26562,N_26381,N_26056);
nor U26563 (N_26563,N_26259,N_26061);
nor U26564 (N_26564,N_26107,N_25990);
nand U26565 (N_26565,N_26263,N_26388);
and U26566 (N_26566,N_26033,N_26327);
nand U26567 (N_26567,N_26116,N_26222);
or U26568 (N_26568,N_26195,N_26386);
or U26569 (N_26569,N_26085,N_26104);
nor U26570 (N_26570,N_26081,N_25842);
xor U26571 (N_26571,N_25954,N_26322);
and U26572 (N_26572,N_26048,N_25949);
xor U26573 (N_26573,N_26001,N_26229);
nor U26574 (N_26574,N_26002,N_26369);
nand U26575 (N_26575,N_26265,N_25824);
or U26576 (N_26576,N_26180,N_26042);
nand U26577 (N_26577,N_25970,N_25819);
xor U26578 (N_26578,N_25926,N_26018);
nand U26579 (N_26579,N_25893,N_26017);
nor U26580 (N_26580,N_25935,N_26198);
and U26581 (N_26581,N_26143,N_26098);
or U26582 (N_26582,N_26370,N_26108);
nor U26583 (N_26583,N_25972,N_26328);
nor U26584 (N_26584,N_26182,N_25906);
nor U26585 (N_26585,N_26171,N_25930);
or U26586 (N_26586,N_26140,N_26300);
and U26587 (N_26587,N_26122,N_25896);
or U26588 (N_26588,N_25944,N_25937);
or U26589 (N_26589,N_26210,N_26100);
nand U26590 (N_26590,N_25909,N_26045);
and U26591 (N_26591,N_25862,N_25838);
nor U26592 (N_26592,N_25870,N_26086);
nor U26593 (N_26593,N_25881,N_26242);
nand U26594 (N_26594,N_25816,N_26326);
and U26595 (N_26595,N_26375,N_25964);
and U26596 (N_26596,N_25931,N_26181);
or U26597 (N_26597,N_26231,N_25960);
nor U26598 (N_26598,N_26067,N_26063);
or U26599 (N_26599,N_26012,N_26251);
nor U26600 (N_26600,N_25859,N_26273);
nor U26601 (N_26601,N_25902,N_26114);
or U26602 (N_26602,N_26043,N_26344);
or U26603 (N_26603,N_25950,N_25882);
nand U26604 (N_26604,N_25880,N_26123);
and U26605 (N_26605,N_25953,N_26257);
nand U26606 (N_26606,N_26031,N_26130);
or U26607 (N_26607,N_26167,N_25971);
or U26608 (N_26608,N_26005,N_26162);
and U26609 (N_26609,N_26091,N_26221);
xnor U26610 (N_26610,N_26335,N_25904);
and U26611 (N_26611,N_25905,N_25826);
or U26612 (N_26612,N_26010,N_25829);
nor U26613 (N_26613,N_26325,N_26011);
and U26614 (N_26614,N_26150,N_26084);
or U26615 (N_26615,N_25834,N_26083);
or U26616 (N_26616,N_26178,N_26342);
nand U26617 (N_26617,N_26398,N_26364);
nand U26618 (N_26618,N_26365,N_26272);
nor U26619 (N_26619,N_26347,N_26268);
xor U26620 (N_26620,N_25923,N_26237);
or U26621 (N_26621,N_26389,N_25877);
nor U26622 (N_26622,N_26281,N_25853);
or U26623 (N_26623,N_26069,N_26234);
or U26624 (N_26624,N_26080,N_26394);
nand U26625 (N_26625,N_26297,N_26174);
nor U26626 (N_26626,N_26022,N_26142);
nand U26627 (N_26627,N_26147,N_26319);
xor U26628 (N_26628,N_25958,N_26367);
or U26629 (N_26629,N_26096,N_25864);
nand U26630 (N_26630,N_25879,N_26343);
nand U26631 (N_26631,N_26079,N_26354);
nor U26632 (N_26632,N_25985,N_26014);
xor U26633 (N_26633,N_26247,N_26173);
and U26634 (N_26634,N_26278,N_25912);
nor U26635 (N_26635,N_25959,N_25963);
nand U26636 (N_26636,N_25965,N_26264);
xnor U26637 (N_26637,N_26399,N_26034);
or U26638 (N_26638,N_26184,N_26283);
nand U26639 (N_26639,N_26212,N_26097);
or U26640 (N_26640,N_26120,N_25987);
or U26641 (N_26641,N_25981,N_25847);
nand U26642 (N_26642,N_25825,N_26320);
nand U26643 (N_26643,N_25807,N_26152);
nor U26644 (N_26644,N_25806,N_26023);
xnor U26645 (N_26645,N_26076,N_25854);
xnor U26646 (N_26646,N_25821,N_26094);
and U26647 (N_26647,N_25917,N_26035);
nand U26648 (N_26648,N_26292,N_26028);
nor U26649 (N_26649,N_26250,N_26051);
and U26650 (N_26650,N_26044,N_26249);
xor U26651 (N_26651,N_25850,N_26156);
nand U26652 (N_26652,N_26271,N_25986);
nor U26653 (N_26653,N_26275,N_26131);
and U26654 (N_26654,N_26191,N_26285);
nor U26655 (N_26655,N_26248,N_26111);
nand U26656 (N_26656,N_26071,N_26055);
nand U26657 (N_26657,N_26383,N_26380);
xnor U26658 (N_26658,N_26211,N_25938);
and U26659 (N_26659,N_25845,N_26106);
nor U26660 (N_26660,N_25868,N_25855);
and U26661 (N_26661,N_26036,N_26202);
or U26662 (N_26662,N_26146,N_25969);
xnor U26663 (N_26663,N_26351,N_26204);
xor U26664 (N_26664,N_26050,N_25844);
and U26665 (N_26665,N_25894,N_26208);
xor U26666 (N_26666,N_26252,N_25911);
xor U26667 (N_26667,N_26199,N_26112);
and U26668 (N_26668,N_25899,N_26078);
xor U26669 (N_26669,N_25890,N_25977);
nand U26670 (N_26670,N_26064,N_26317);
and U26671 (N_26671,N_26176,N_26243);
and U26672 (N_26672,N_25910,N_26371);
nor U26673 (N_26673,N_26301,N_26101);
or U26674 (N_26674,N_26362,N_26164);
nand U26675 (N_26675,N_25974,N_26021);
xor U26676 (N_26676,N_26077,N_25811);
or U26677 (N_26677,N_26339,N_25856);
nand U26678 (N_26678,N_26310,N_25936);
and U26679 (N_26679,N_26379,N_26336);
and U26680 (N_26680,N_25871,N_26197);
xor U26681 (N_26681,N_26235,N_26228);
or U26682 (N_26682,N_25943,N_26313);
nor U26683 (N_26683,N_25942,N_25945);
and U26684 (N_26684,N_25840,N_26323);
xor U26685 (N_26685,N_26040,N_26163);
or U26686 (N_26686,N_26217,N_26254);
nand U26687 (N_26687,N_25863,N_26054);
nand U26688 (N_26688,N_26355,N_26316);
or U26689 (N_26689,N_26088,N_26125);
nand U26690 (N_26690,N_25801,N_26119);
or U26691 (N_26691,N_25921,N_25988);
xor U26692 (N_26692,N_25835,N_26277);
and U26693 (N_26693,N_25914,N_26065);
and U26694 (N_26694,N_26216,N_26102);
nand U26695 (N_26695,N_26245,N_26157);
or U26696 (N_26696,N_26165,N_26185);
and U26697 (N_26697,N_25884,N_25966);
nor U26698 (N_26698,N_25860,N_26127);
or U26699 (N_26699,N_25984,N_25810);
or U26700 (N_26700,N_26140,N_26349);
nor U26701 (N_26701,N_25862,N_26226);
and U26702 (N_26702,N_26003,N_25879);
nor U26703 (N_26703,N_26349,N_26092);
and U26704 (N_26704,N_26211,N_25969);
or U26705 (N_26705,N_26050,N_26377);
nand U26706 (N_26706,N_26366,N_26203);
xnor U26707 (N_26707,N_26254,N_25932);
and U26708 (N_26708,N_26083,N_25807);
or U26709 (N_26709,N_26147,N_25805);
nor U26710 (N_26710,N_25991,N_26251);
nor U26711 (N_26711,N_25879,N_26140);
and U26712 (N_26712,N_25919,N_25815);
or U26713 (N_26713,N_25998,N_25909);
nor U26714 (N_26714,N_26238,N_25869);
nand U26715 (N_26715,N_26325,N_26028);
or U26716 (N_26716,N_26079,N_26239);
or U26717 (N_26717,N_26292,N_26119);
or U26718 (N_26718,N_26041,N_25862);
nor U26719 (N_26719,N_26380,N_26275);
or U26720 (N_26720,N_26015,N_25935);
xnor U26721 (N_26721,N_25966,N_26363);
or U26722 (N_26722,N_26176,N_26141);
or U26723 (N_26723,N_26010,N_25896);
or U26724 (N_26724,N_26039,N_26233);
or U26725 (N_26725,N_26024,N_25926);
xor U26726 (N_26726,N_25847,N_26295);
nand U26727 (N_26727,N_26280,N_26301);
and U26728 (N_26728,N_26352,N_26367);
and U26729 (N_26729,N_26384,N_26153);
nor U26730 (N_26730,N_26357,N_25887);
xor U26731 (N_26731,N_26035,N_25919);
nor U26732 (N_26732,N_25901,N_26384);
xnor U26733 (N_26733,N_26388,N_26338);
or U26734 (N_26734,N_26085,N_26318);
xnor U26735 (N_26735,N_26026,N_25953);
nor U26736 (N_26736,N_25879,N_26270);
and U26737 (N_26737,N_26338,N_26386);
nor U26738 (N_26738,N_26233,N_26077);
and U26739 (N_26739,N_26135,N_26294);
or U26740 (N_26740,N_26376,N_26338);
or U26741 (N_26741,N_26220,N_26208);
and U26742 (N_26742,N_26142,N_26221);
nand U26743 (N_26743,N_25834,N_25808);
nand U26744 (N_26744,N_25855,N_25937);
nand U26745 (N_26745,N_25980,N_26291);
or U26746 (N_26746,N_25907,N_26149);
xnor U26747 (N_26747,N_25847,N_26315);
and U26748 (N_26748,N_26390,N_26108);
and U26749 (N_26749,N_26148,N_26258);
xnor U26750 (N_26750,N_26064,N_26017);
or U26751 (N_26751,N_26081,N_26161);
nor U26752 (N_26752,N_26056,N_26007);
and U26753 (N_26753,N_26138,N_25819);
nand U26754 (N_26754,N_26260,N_26123);
nand U26755 (N_26755,N_25911,N_25921);
nand U26756 (N_26756,N_26217,N_25906);
nand U26757 (N_26757,N_26308,N_25878);
xor U26758 (N_26758,N_26022,N_25927);
and U26759 (N_26759,N_26033,N_26387);
and U26760 (N_26760,N_25997,N_26226);
or U26761 (N_26761,N_26222,N_25862);
and U26762 (N_26762,N_26373,N_26247);
nand U26763 (N_26763,N_25998,N_25861);
or U26764 (N_26764,N_26336,N_26221);
nor U26765 (N_26765,N_26197,N_26027);
nand U26766 (N_26766,N_26325,N_25835);
nor U26767 (N_26767,N_26349,N_26225);
nor U26768 (N_26768,N_25850,N_26239);
nor U26769 (N_26769,N_25841,N_26207);
or U26770 (N_26770,N_26372,N_26393);
nand U26771 (N_26771,N_25905,N_25934);
nand U26772 (N_26772,N_26381,N_26098);
nor U26773 (N_26773,N_25997,N_25972);
and U26774 (N_26774,N_26168,N_26032);
and U26775 (N_26775,N_26399,N_26211);
xnor U26776 (N_26776,N_25854,N_26102);
nor U26777 (N_26777,N_26079,N_26035);
or U26778 (N_26778,N_26228,N_25956);
or U26779 (N_26779,N_25973,N_26215);
nand U26780 (N_26780,N_26243,N_25842);
xnor U26781 (N_26781,N_26002,N_25929);
xnor U26782 (N_26782,N_25888,N_25862);
or U26783 (N_26783,N_26357,N_26197);
nor U26784 (N_26784,N_26179,N_26183);
xor U26785 (N_26785,N_25875,N_25878);
nand U26786 (N_26786,N_25969,N_26040);
or U26787 (N_26787,N_25936,N_26086);
or U26788 (N_26788,N_25909,N_26040);
and U26789 (N_26789,N_25934,N_26311);
nand U26790 (N_26790,N_26378,N_26161);
nor U26791 (N_26791,N_26215,N_26386);
and U26792 (N_26792,N_26186,N_25960);
nand U26793 (N_26793,N_26157,N_26139);
nand U26794 (N_26794,N_26329,N_26013);
nor U26795 (N_26795,N_26221,N_26291);
or U26796 (N_26796,N_26265,N_26388);
nand U26797 (N_26797,N_25917,N_26390);
xor U26798 (N_26798,N_26073,N_25914);
and U26799 (N_26799,N_26209,N_26066);
nor U26800 (N_26800,N_26057,N_25953);
nand U26801 (N_26801,N_26092,N_26245);
or U26802 (N_26802,N_25878,N_26139);
nand U26803 (N_26803,N_26106,N_26317);
or U26804 (N_26804,N_26346,N_26102);
nand U26805 (N_26805,N_25809,N_26196);
nand U26806 (N_26806,N_26182,N_26030);
or U26807 (N_26807,N_25971,N_26098);
nand U26808 (N_26808,N_26100,N_26378);
or U26809 (N_26809,N_25840,N_26221);
nor U26810 (N_26810,N_25812,N_25980);
nor U26811 (N_26811,N_25920,N_25935);
nand U26812 (N_26812,N_26060,N_26072);
nor U26813 (N_26813,N_25896,N_25832);
xnor U26814 (N_26814,N_25915,N_25826);
and U26815 (N_26815,N_25925,N_25978);
nor U26816 (N_26816,N_26272,N_26185);
nand U26817 (N_26817,N_26178,N_26155);
nor U26818 (N_26818,N_25898,N_26116);
nand U26819 (N_26819,N_26276,N_25875);
nor U26820 (N_26820,N_26349,N_25998);
or U26821 (N_26821,N_26183,N_25892);
and U26822 (N_26822,N_25861,N_26037);
and U26823 (N_26823,N_25857,N_25923);
and U26824 (N_26824,N_26248,N_25957);
xnor U26825 (N_26825,N_26200,N_26195);
nor U26826 (N_26826,N_26357,N_26388);
and U26827 (N_26827,N_26375,N_26119);
and U26828 (N_26828,N_25917,N_26050);
xor U26829 (N_26829,N_25967,N_25934);
xnor U26830 (N_26830,N_26324,N_26395);
xor U26831 (N_26831,N_26244,N_25955);
or U26832 (N_26832,N_25832,N_26257);
and U26833 (N_26833,N_25983,N_26307);
or U26834 (N_26834,N_25829,N_26313);
or U26835 (N_26835,N_26196,N_26153);
xor U26836 (N_26836,N_26328,N_25989);
xnor U26837 (N_26837,N_26059,N_26272);
nand U26838 (N_26838,N_25805,N_26343);
and U26839 (N_26839,N_25923,N_26247);
or U26840 (N_26840,N_25940,N_25981);
nand U26841 (N_26841,N_25875,N_26092);
nand U26842 (N_26842,N_26175,N_26174);
nor U26843 (N_26843,N_25973,N_26303);
nor U26844 (N_26844,N_26146,N_25934);
nor U26845 (N_26845,N_26123,N_26195);
and U26846 (N_26846,N_26269,N_26291);
or U26847 (N_26847,N_25926,N_25848);
or U26848 (N_26848,N_26250,N_25820);
nor U26849 (N_26849,N_26215,N_25875);
nor U26850 (N_26850,N_26176,N_26318);
and U26851 (N_26851,N_25836,N_26124);
nor U26852 (N_26852,N_26143,N_26120);
nand U26853 (N_26853,N_26061,N_26231);
nor U26854 (N_26854,N_26126,N_26314);
and U26855 (N_26855,N_25955,N_26355);
nor U26856 (N_26856,N_26154,N_26113);
nand U26857 (N_26857,N_25894,N_26337);
nand U26858 (N_26858,N_25853,N_26245);
and U26859 (N_26859,N_25914,N_25921);
or U26860 (N_26860,N_26044,N_26041);
nand U26861 (N_26861,N_26042,N_26369);
or U26862 (N_26862,N_26158,N_26129);
or U26863 (N_26863,N_26159,N_26318);
and U26864 (N_26864,N_26185,N_25852);
and U26865 (N_26865,N_26121,N_26128);
nor U26866 (N_26866,N_26039,N_26092);
nor U26867 (N_26867,N_26193,N_25851);
and U26868 (N_26868,N_25987,N_26059);
or U26869 (N_26869,N_25860,N_25934);
xnor U26870 (N_26870,N_26218,N_26094);
nor U26871 (N_26871,N_26326,N_26042);
nand U26872 (N_26872,N_26175,N_26388);
nor U26873 (N_26873,N_26065,N_26140);
nor U26874 (N_26874,N_26030,N_26173);
nand U26875 (N_26875,N_25805,N_26148);
nor U26876 (N_26876,N_25860,N_26162);
and U26877 (N_26877,N_26356,N_26390);
or U26878 (N_26878,N_26041,N_25972);
or U26879 (N_26879,N_26100,N_25825);
nand U26880 (N_26880,N_26199,N_26142);
or U26881 (N_26881,N_26363,N_25804);
and U26882 (N_26882,N_26126,N_26049);
or U26883 (N_26883,N_26389,N_26152);
nor U26884 (N_26884,N_26039,N_26089);
nor U26885 (N_26885,N_26031,N_26280);
and U26886 (N_26886,N_25865,N_26194);
nor U26887 (N_26887,N_26195,N_25825);
nand U26888 (N_26888,N_26058,N_25913);
or U26889 (N_26889,N_25817,N_25858);
nand U26890 (N_26890,N_26248,N_26197);
nor U26891 (N_26891,N_26101,N_26005);
and U26892 (N_26892,N_26184,N_25916);
nor U26893 (N_26893,N_26063,N_26088);
and U26894 (N_26894,N_25846,N_26150);
nor U26895 (N_26895,N_25948,N_26382);
xnor U26896 (N_26896,N_26197,N_25849);
nor U26897 (N_26897,N_26334,N_26166);
or U26898 (N_26898,N_25905,N_26108);
nand U26899 (N_26899,N_26136,N_25871);
nand U26900 (N_26900,N_26219,N_25935);
xnor U26901 (N_26901,N_25903,N_26024);
nand U26902 (N_26902,N_26077,N_25948);
or U26903 (N_26903,N_26118,N_25802);
nand U26904 (N_26904,N_25920,N_25921);
nor U26905 (N_26905,N_26184,N_26374);
nand U26906 (N_26906,N_26343,N_26059);
and U26907 (N_26907,N_26152,N_26368);
and U26908 (N_26908,N_26299,N_25823);
and U26909 (N_26909,N_26113,N_25946);
and U26910 (N_26910,N_26240,N_26323);
nor U26911 (N_26911,N_26030,N_26163);
or U26912 (N_26912,N_26346,N_26112);
or U26913 (N_26913,N_25903,N_26234);
nor U26914 (N_26914,N_26156,N_26382);
nor U26915 (N_26915,N_26258,N_25809);
nor U26916 (N_26916,N_26251,N_26362);
xor U26917 (N_26917,N_25834,N_26296);
nand U26918 (N_26918,N_25889,N_26052);
and U26919 (N_26919,N_26260,N_26381);
or U26920 (N_26920,N_26230,N_25803);
nand U26921 (N_26921,N_26064,N_26045);
nor U26922 (N_26922,N_26265,N_25849);
and U26923 (N_26923,N_25854,N_26217);
and U26924 (N_26924,N_26032,N_25977);
nand U26925 (N_26925,N_26064,N_26351);
and U26926 (N_26926,N_25800,N_25964);
nand U26927 (N_26927,N_25877,N_26298);
nand U26928 (N_26928,N_26281,N_25860);
xor U26929 (N_26929,N_25944,N_25982);
and U26930 (N_26930,N_25926,N_26011);
xor U26931 (N_26931,N_25818,N_26284);
nand U26932 (N_26932,N_26337,N_25955);
xor U26933 (N_26933,N_26109,N_25991);
nand U26934 (N_26934,N_26367,N_26168);
nand U26935 (N_26935,N_26057,N_26238);
nand U26936 (N_26936,N_25817,N_26037);
and U26937 (N_26937,N_26385,N_26068);
or U26938 (N_26938,N_26042,N_26064);
and U26939 (N_26939,N_26036,N_25984);
nor U26940 (N_26940,N_26256,N_26037);
nand U26941 (N_26941,N_26302,N_26268);
and U26942 (N_26942,N_25828,N_26236);
or U26943 (N_26943,N_26261,N_25985);
nand U26944 (N_26944,N_25831,N_25913);
and U26945 (N_26945,N_25912,N_26207);
nor U26946 (N_26946,N_25961,N_25897);
and U26947 (N_26947,N_26374,N_26004);
nand U26948 (N_26948,N_26341,N_25846);
or U26949 (N_26949,N_26299,N_25910);
and U26950 (N_26950,N_25822,N_26101);
and U26951 (N_26951,N_26251,N_26229);
nor U26952 (N_26952,N_26155,N_26373);
nand U26953 (N_26953,N_25990,N_26283);
and U26954 (N_26954,N_26066,N_26326);
nand U26955 (N_26955,N_26297,N_25976);
nor U26956 (N_26956,N_25986,N_25802);
or U26957 (N_26957,N_26142,N_25857);
or U26958 (N_26958,N_26097,N_26084);
nor U26959 (N_26959,N_26025,N_26238);
nand U26960 (N_26960,N_26020,N_25903);
and U26961 (N_26961,N_26253,N_25823);
or U26962 (N_26962,N_25949,N_26343);
or U26963 (N_26963,N_25862,N_26030);
nand U26964 (N_26964,N_26340,N_25869);
and U26965 (N_26965,N_26310,N_26181);
xor U26966 (N_26966,N_26390,N_26204);
xor U26967 (N_26967,N_26374,N_25803);
or U26968 (N_26968,N_26280,N_25921);
xor U26969 (N_26969,N_25998,N_26023);
nand U26970 (N_26970,N_26345,N_26169);
nor U26971 (N_26971,N_26314,N_26193);
xnor U26972 (N_26972,N_26208,N_26165);
nand U26973 (N_26973,N_26398,N_26035);
nor U26974 (N_26974,N_26178,N_26126);
or U26975 (N_26975,N_26189,N_25940);
or U26976 (N_26976,N_26308,N_25834);
nand U26977 (N_26977,N_26392,N_26211);
and U26978 (N_26978,N_26190,N_26392);
nand U26979 (N_26979,N_25996,N_26203);
or U26980 (N_26980,N_25842,N_25975);
or U26981 (N_26981,N_26061,N_26204);
or U26982 (N_26982,N_25934,N_26018);
and U26983 (N_26983,N_26280,N_26164);
nor U26984 (N_26984,N_26122,N_26155);
and U26985 (N_26985,N_26238,N_26032);
xor U26986 (N_26986,N_26059,N_26291);
nand U26987 (N_26987,N_26345,N_26242);
nand U26988 (N_26988,N_26206,N_25939);
or U26989 (N_26989,N_25815,N_26032);
and U26990 (N_26990,N_25846,N_25832);
or U26991 (N_26991,N_26309,N_26161);
and U26992 (N_26992,N_25949,N_26190);
xor U26993 (N_26993,N_26271,N_26150);
nor U26994 (N_26994,N_25924,N_26183);
nor U26995 (N_26995,N_25861,N_26346);
nand U26996 (N_26996,N_25815,N_26107);
xor U26997 (N_26997,N_26158,N_26334);
xor U26998 (N_26998,N_25836,N_25873);
nand U26999 (N_26999,N_26117,N_25948);
nand U27000 (N_27000,N_26626,N_26706);
nor U27001 (N_27001,N_26430,N_26793);
nand U27002 (N_27002,N_26742,N_26577);
and U27003 (N_27003,N_26778,N_26897);
nand U27004 (N_27004,N_26894,N_26705);
nand U27005 (N_27005,N_26614,N_26676);
and U27006 (N_27006,N_26752,N_26491);
nor U27007 (N_27007,N_26966,N_26525);
xor U27008 (N_27008,N_26432,N_26629);
xor U27009 (N_27009,N_26483,N_26587);
or U27010 (N_27010,N_26600,N_26848);
and U27011 (N_27011,N_26630,N_26740);
and U27012 (N_27012,N_26883,N_26866);
nor U27013 (N_27013,N_26790,N_26685);
or U27014 (N_27014,N_26786,N_26610);
nand U27015 (N_27015,N_26689,N_26726);
or U27016 (N_27016,N_26962,N_26604);
xor U27017 (N_27017,N_26990,N_26542);
nand U27018 (N_27018,N_26869,N_26949);
nand U27019 (N_27019,N_26646,N_26903);
and U27020 (N_27020,N_26765,N_26414);
or U27021 (N_27021,N_26932,N_26548);
nand U27022 (N_27022,N_26720,N_26977);
nor U27023 (N_27023,N_26888,N_26423);
and U27024 (N_27024,N_26463,N_26677);
and U27025 (N_27025,N_26519,N_26531);
nor U27026 (N_27026,N_26405,N_26737);
and U27027 (N_27027,N_26582,N_26514);
or U27028 (N_27028,N_26942,N_26656);
nor U27029 (N_27029,N_26798,N_26973);
or U27030 (N_27030,N_26593,N_26540);
and U27031 (N_27031,N_26641,N_26533);
and U27032 (N_27032,N_26708,N_26821);
or U27033 (N_27033,N_26832,N_26671);
and U27034 (N_27034,N_26880,N_26684);
and U27035 (N_27035,N_26748,N_26701);
or U27036 (N_27036,N_26958,N_26484);
nor U27037 (N_27037,N_26722,N_26675);
and U27038 (N_27038,N_26861,N_26657);
or U27039 (N_27039,N_26695,N_26594);
and U27040 (N_27040,N_26851,N_26744);
and U27041 (N_27041,N_26856,N_26743);
xor U27042 (N_27042,N_26444,N_26833);
or U27043 (N_27043,N_26824,N_26855);
or U27044 (N_27044,N_26960,N_26950);
nor U27045 (N_27045,N_26905,N_26565);
nand U27046 (N_27046,N_26835,N_26789);
nor U27047 (N_27047,N_26490,N_26486);
xor U27048 (N_27048,N_26443,N_26546);
or U27049 (N_27049,N_26749,N_26874);
xor U27050 (N_27050,N_26598,N_26899);
nand U27051 (N_27051,N_26710,N_26475);
or U27052 (N_27052,N_26516,N_26415);
or U27053 (N_27053,N_26758,N_26918);
nand U27054 (N_27054,N_26761,N_26434);
nand U27055 (N_27055,N_26844,N_26556);
nor U27056 (N_27056,N_26885,N_26760);
or U27057 (N_27057,N_26550,N_26733);
or U27058 (N_27058,N_26755,N_26800);
nand U27059 (N_27059,N_26609,N_26538);
xnor U27060 (N_27060,N_26995,N_26687);
xor U27061 (N_27061,N_26471,N_26619);
and U27062 (N_27062,N_26402,N_26795);
xor U27063 (N_27063,N_26948,N_26964);
nor U27064 (N_27064,N_26882,N_26602);
nand U27065 (N_27065,N_26834,N_26853);
nor U27066 (N_27066,N_26569,N_26818);
nor U27067 (N_27067,N_26508,N_26728);
or U27068 (N_27068,N_26713,N_26502);
and U27069 (N_27069,N_26469,N_26745);
nor U27070 (N_27070,N_26939,N_26766);
xor U27071 (N_27071,N_26418,N_26972);
nand U27072 (N_27072,N_26771,N_26725);
nand U27073 (N_27073,N_26757,N_26498);
or U27074 (N_27074,N_26764,N_26480);
nand U27075 (N_27075,N_26460,N_26754);
and U27076 (N_27076,N_26476,N_26497);
or U27077 (N_27077,N_26530,N_26524);
nor U27078 (N_27078,N_26830,N_26961);
nand U27079 (N_27079,N_26563,N_26534);
nand U27080 (N_27080,N_26521,N_26920);
nor U27081 (N_27081,N_26731,N_26442);
nand U27082 (N_27082,N_26971,N_26464);
xor U27083 (N_27083,N_26727,N_26479);
xnor U27084 (N_27084,N_26886,N_26583);
and U27085 (N_27085,N_26980,N_26586);
or U27086 (N_27086,N_26819,N_26691);
xnor U27087 (N_27087,N_26455,N_26421);
or U27088 (N_27088,N_26683,N_26408);
nand U27089 (N_27089,N_26867,N_26978);
xor U27090 (N_27090,N_26784,N_26732);
and U27091 (N_27091,N_26906,N_26769);
or U27092 (N_27092,N_26605,N_26924);
and U27093 (N_27093,N_26747,N_26581);
nor U27094 (N_27094,N_26661,N_26511);
and U27095 (N_27095,N_26453,N_26400);
or U27096 (N_27096,N_26631,N_26570);
nand U27097 (N_27097,N_26670,N_26551);
nor U27098 (N_27098,N_26679,N_26810);
or U27099 (N_27099,N_26998,N_26986);
xor U27100 (N_27100,N_26714,N_26893);
nand U27101 (N_27101,N_26527,N_26751);
and U27102 (N_27102,N_26723,N_26428);
and U27103 (N_27103,N_26987,N_26815);
or U27104 (N_27104,N_26739,N_26787);
nand U27105 (N_27105,N_26774,N_26804);
nor U27106 (N_27106,N_26952,N_26997);
nand U27107 (N_27107,N_26823,N_26578);
nor U27108 (N_27108,N_26608,N_26473);
nor U27109 (N_27109,N_26681,N_26857);
nand U27110 (N_27110,N_26493,N_26648);
and U27111 (N_27111,N_26505,N_26572);
and U27112 (N_27112,N_26644,N_26999);
and U27113 (N_27113,N_26518,N_26707);
and U27114 (N_27114,N_26552,N_26775);
nor U27115 (N_27115,N_26612,N_26788);
nor U27116 (N_27116,N_26445,N_26930);
or U27117 (N_27117,N_26425,N_26427);
nand U27118 (N_27118,N_26495,N_26702);
nand U27119 (N_27119,N_26763,N_26811);
nand U27120 (N_27120,N_26864,N_26773);
or U27121 (N_27121,N_26943,N_26965);
nand U27122 (N_27122,N_26913,N_26596);
or U27123 (N_27123,N_26472,N_26808);
nor U27124 (N_27124,N_26543,N_26426);
nor U27125 (N_27125,N_26996,N_26624);
and U27126 (N_27126,N_26412,N_26523);
nor U27127 (N_27127,N_26579,N_26509);
nand U27128 (N_27128,N_26459,N_26450);
nor U27129 (N_27129,N_26500,N_26557);
or U27130 (N_27130,N_26916,N_26532);
nor U27131 (N_27131,N_26481,N_26925);
or U27132 (N_27132,N_26506,N_26709);
nor U27133 (N_27133,N_26911,N_26881);
or U27134 (N_27134,N_26983,N_26663);
and U27135 (N_27135,N_26776,N_26892);
nand U27136 (N_27136,N_26777,N_26416);
and U27137 (N_27137,N_26558,N_26574);
or U27138 (N_27138,N_26877,N_26467);
or U27139 (N_27139,N_26654,N_26576);
and U27140 (N_27140,N_26847,N_26665);
nor U27141 (N_27141,N_26649,N_26896);
nor U27142 (N_27142,N_26741,N_26912);
or U27143 (N_27143,N_26528,N_26780);
nand U27144 (N_27144,N_26955,N_26976);
or U27145 (N_27145,N_26696,N_26822);
nand U27146 (N_27146,N_26994,N_26974);
nand U27147 (N_27147,N_26436,N_26621);
nor U27148 (N_27148,N_26424,N_26831);
nand U27149 (N_27149,N_26828,N_26607);
or U27150 (N_27150,N_26802,N_26501);
nand U27151 (N_27151,N_26940,N_26721);
or U27152 (N_27152,N_26410,N_26870);
xnor U27153 (N_27153,N_26568,N_26711);
nor U27154 (N_27154,N_26917,N_26873);
xor U27155 (N_27155,N_26627,N_26555);
and U27156 (N_27156,N_26461,N_26653);
or U27157 (N_27157,N_26618,N_26719);
nor U27158 (N_27158,N_26597,N_26512);
and U27159 (N_27159,N_26448,N_26541);
nand U27160 (N_27160,N_26813,N_26839);
xor U27161 (N_27161,N_26560,N_26736);
nor U27162 (N_27162,N_26845,N_26431);
nand U27163 (N_27163,N_26573,N_26933);
nor U27164 (N_27164,N_26781,N_26664);
or U27165 (N_27165,N_26536,N_26876);
nand U27166 (N_27166,N_26515,N_26858);
xnor U27167 (N_27167,N_26931,N_26561);
xor U27168 (N_27168,N_26984,N_26606);
and U27169 (N_27169,N_26992,N_26651);
and U27170 (N_27170,N_26553,N_26884);
and U27171 (N_27171,N_26891,N_26829);
nor U27172 (N_27172,N_26470,N_26645);
nand U27173 (N_27173,N_26628,N_26441);
nand U27174 (N_27174,N_26575,N_26796);
nand U27175 (N_27175,N_26915,N_26817);
or U27176 (N_27176,N_26639,N_26989);
or U27177 (N_27177,N_26953,N_26499);
and U27178 (N_27178,N_26636,N_26988);
nand U27179 (N_27179,N_26717,N_26584);
and U27180 (N_27180,N_26993,N_26746);
nand U27181 (N_27181,N_26487,N_26878);
or U27182 (N_27182,N_26836,N_26406);
or U27183 (N_27183,N_26566,N_26941);
and U27184 (N_27184,N_26794,N_26633);
and U27185 (N_27185,N_26951,N_26447);
nand U27186 (N_27186,N_26782,N_26634);
or U27187 (N_27187,N_26843,N_26507);
and U27188 (N_27188,N_26446,N_26504);
nand U27189 (N_27189,N_26682,N_26935);
xnor U27190 (N_27190,N_26826,N_26842);
nor U27191 (N_27191,N_26545,N_26513);
nand U27192 (N_27192,N_26922,N_26623);
nor U27193 (N_27193,N_26729,N_26970);
nor U27194 (N_27194,N_26954,N_26936);
nand U27195 (N_27195,N_26674,N_26975);
xor U27196 (N_27196,N_26738,N_26868);
or U27197 (N_27197,N_26640,N_26693);
nor U27198 (N_27198,N_26890,N_26547);
and U27199 (N_27199,N_26840,N_26872);
or U27200 (N_27200,N_26809,N_26734);
or U27201 (N_27201,N_26452,N_26750);
nor U27202 (N_27202,N_26852,N_26599);
or U27203 (N_27203,N_26680,N_26959);
or U27204 (N_27204,N_26718,N_26946);
xor U27205 (N_27205,N_26712,N_26716);
nor U27206 (N_27206,N_26429,N_26590);
nor U27207 (N_27207,N_26642,N_26660);
nand U27208 (N_27208,N_26699,N_26979);
and U27209 (N_27209,N_26413,N_26482);
or U27210 (N_27210,N_26403,N_26860);
xnor U27211 (N_27211,N_26419,N_26859);
and U27212 (N_27212,N_26704,N_26875);
nor U27213 (N_27213,N_26820,N_26635);
and U27214 (N_27214,N_26549,N_26603);
and U27215 (N_27215,N_26535,N_26567);
or U27216 (N_27216,N_26827,N_26615);
nor U27217 (N_27217,N_26724,N_26417);
and U27218 (N_27218,N_26816,N_26753);
and U27219 (N_27219,N_26929,N_26667);
nor U27220 (N_27220,N_26921,N_26692);
nand U27221 (N_27221,N_26456,N_26458);
or U27222 (N_27222,N_26554,N_26433);
and U27223 (N_27223,N_26411,N_26871);
or U27224 (N_27224,N_26889,N_26901);
nor U27225 (N_27225,N_26956,N_26934);
and U27226 (N_27226,N_26910,N_26601);
nor U27227 (N_27227,N_26814,N_26909);
xnor U27228 (N_27228,N_26647,N_26468);
and U27229 (N_27229,N_26799,N_26902);
and U27230 (N_27230,N_26617,N_26401);
and U27231 (N_27231,N_26474,N_26489);
nor U27232 (N_27232,N_26658,N_26620);
and U27233 (N_27233,N_26659,N_26981);
and U27234 (N_27234,N_26927,N_26779);
or U27235 (N_27235,N_26907,N_26862);
nand U27236 (N_27236,N_26592,N_26564);
nor U27237 (N_27237,N_26985,N_26703);
and U27238 (N_27238,N_26947,N_26967);
nand U27239 (N_27239,N_26544,N_26895);
nor U27240 (N_27240,N_26825,N_26517);
nor U27241 (N_27241,N_26991,N_26887);
or U27242 (N_27242,N_26437,N_26407);
nor U27243 (N_27243,N_26914,N_26422);
nor U27244 (N_27244,N_26923,N_26580);
nor U27245 (N_27245,N_26638,N_26944);
xor U27246 (N_27246,N_26937,N_26632);
nor U27247 (N_27247,N_26477,N_26945);
or U27248 (N_27248,N_26678,N_26457);
or U27249 (N_27249,N_26846,N_26697);
nor U27250 (N_27250,N_26803,N_26462);
nor U27251 (N_27251,N_26919,N_26449);
xor U27252 (N_27252,N_26438,N_26756);
nand U27253 (N_27253,N_26841,N_26439);
nand U27254 (N_27254,N_26662,N_26928);
and U27255 (N_27255,N_26898,N_26494);
nand U27256 (N_27256,N_26957,N_26837);
or U27257 (N_27257,N_26537,N_26772);
and U27258 (N_27258,N_26451,N_26762);
nor U27259 (N_27259,N_26698,N_26938);
and U27260 (N_27260,N_26792,N_26963);
nor U27261 (N_27261,N_26650,N_26672);
and U27262 (N_27262,N_26559,N_26807);
nor U27263 (N_27263,N_26613,N_26510);
or U27264 (N_27264,N_26865,N_26838);
or U27265 (N_27265,N_26770,N_26591);
xnor U27266 (N_27266,N_26503,N_26404);
nand U27267 (N_27267,N_26690,N_26571);
nor U27268 (N_27268,N_26589,N_26688);
nand U27269 (N_27269,N_26622,N_26759);
nor U27270 (N_27270,N_26562,N_26616);
nand U27271 (N_27271,N_26539,N_26435);
nand U27272 (N_27272,N_26655,N_26904);
xnor U27273 (N_27273,N_26496,N_26908);
and U27274 (N_27274,N_26637,N_26879);
xor U27275 (N_27275,N_26767,N_26715);
xnor U27276 (N_27276,N_26783,N_26588);
nand U27277 (N_27277,N_26673,N_26595);
and U27278 (N_27278,N_26968,N_26791);
nor U27279 (N_27279,N_26805,N_26466);
and U27280 (N_27280,N_26900,N_26801);
nor U27281 (N_27281,N_26625,N_26611);
nand U27282 (N_27282,N_26454,N_26668);
xor U27283 (N_27283,N_26694,N_26440);
and U27284 (N_27284,N_26666,N_26850);
nor U27285 (N_27285,N_26585,N_26409);
and U27286 (N_27286,N_26485,N_26982);
xor U27287 (N_27287,N_26488,N_26669);
nor U27288 (N_27288,N_26768,N_26520);
nand U27289 (N_27289,N_26643,N_26849);
nor U27290 (N_27290,N_26526,N_26785);
and U27291 (N_27291,N_26522,N_26806);
or U27292 (N_27292,N_26686,N_26812);
and U27293 (N_27293,N_26797,N_26969);
and U27294 (N_27294,N_26926,N_26652);
xor U27295 (N_27295,N_26854,N_26863);
nand U27296 (N_27296,N_26420,N_26700);
nand U27297 (N_27297,N_26478,N_26730);
or U27298 (N_27298,N_26735,N_26465);
and U27299 (N_27299,N_26529,N_26492);
nor U27300 (N_27300,N_26985,N_26723);
or U27301 (N_27301,N_26833,N_26854);
and U27302 (N_27302,N_26531,N_26504);
nor U27303 (N_27303,N_26882,N_26898);
or U27304 (N_27304,N_26540,N_26690);
nand U27305 (N_27305,N_26834,N_26759);
and U27306 (N_27306,N_26693,N_26968);
nor U27307 (N_27307,N_26502,N_26595);
xor U27308 (N_27308,N_26526,N_26862);
nor U27309 (N_27309,N_26866,N_26498);
nor U27310 (N_27310,N_26761,N_26577);
nand U27311 (N_27311,N_26909,N_26566);
or U27312 (N_27312,N_26689,N_26727);
or U27313 (N_27313,N_26714,N_26502);
nand U27314 (N_27314,N_26493,N_26401);
nand U27315 (N_27315,N_26920,N_26496);
nand U27316 (N_27316,N_26824,N_26812);
xnor U27317 (N_27317,N_26744,N_26675);
and U27318 (N_27318,N_26620,N_26671);
nand U27319 (N_27319,N_26755,N_26974);
and U27320 (N_27320,N_26669,N_26944);
and U27321 (N_27321,N_26894,N_26564);
or U27322 (N_27322,N_26518,N_26713);
or U27323 (N_27323,N_26646,N_26522);
or U27324 (N_27324,N_26597,N_26574);
xnor U27325 (N_27325,N_26468,N_26490);
nor U27326 (N_27326,N_26635,N_26909);
or U27327 (N_27327,N_26612,N_26476);
or U27328 (N_27328,N_26643,N_26553);
nor U27329 (N_27329,N_26835,N_26454);
nor U27330 (N_27330,N_26794,N_26693);
or U27331 (N_27331,N_26674,N_26480);
nand U27332 (N_27332,N_26779,N_26905);
or U27333 (N_27333,N_26978,N_26546);
or U27334 (N_27334,N_26994,N_26562);
or U27335 (N_27335,N_26431,N_26492);
and U27336 (N_27336,N_26809,N_26716);
nor U27337 (N_27337,N_26610,N_26580);
nor U27338 (N_27338,N_26537,N_26843);
and U27339 (N_27339,N_26874,N_26679);
and U27340 (N_27340,N_26980,N_26949);
nand U27341 (N_27341,N_26808,N_26438);
or U27342 (N_27342,N_26466,N_26480);
xnor U27343 (N_27343,N_26766,N_26674);
nor U27344 (N_27344,N_26945,N_26664);
or U27345 (N_27345,N_26493,N_26559);
nor U27346 (N_27346,N_26513,N_26785);
or U27347 (N_27347,N_26553,N_26595);
nor U27348 (N_27348,N_26719,N_26786);
or U27349 (N_27349,N_26728,N_26779);
and U27350 (N_27350,N_26772,N_26463);
nor U27351 (N_27351,N_26819,N_26747);
and U27352 (N_27352,N_26513,N_26988);
nand U27353 (N_27353,N_26918,N_26685);
xor U27354 (N_27354,N_26684,N_26700);
and U27355 (N_27355,N_26451,N_26794);
nand U27356 (N_27356,N_26735,N_26461);
nor U27357 (N_27357,N_26750,N_26893);
or U27358 (N_27358,N_26687,N_26735);
or U27359 (N_27359,N_26856,N_26809);
or U27360 (N_27360,N_26611,N_26935);
or U27361 (N_27361,N_26848,N_26906);
nor U27362 (N_27362,N_26403,N_26588);
nor U27363 (N_27363,N_26557,N_26515);
nand U27364 (N_27364,N_26551,N_26865);
xor U27365 (N_27365,N_26975,N_26628);
and U27366 (N_27366,N_26729,N_26950);
and U27367 (N_27367,N_26909,N_26990);
or U27368 (N_27368,N_26870,N_26580);
or U27369 (N_27369,N_26422,N_26535);
or U27370 (N_27370,N_26530,N_26503);
or U27371 (N_27371,N_26669,N_26457);
and U27372 (N_27372,N_26632,N_26517);
nand U27373 (N_27373,N_26831,N_26689);
or U27374 (N_27374,N_26930,N_26630);
nor U27375 (N_27375,N_26842,N_26724);
nand U27376 (N_27376,N_26892,N_26713);
or U27377 (N_27377,N_26595,N_26453);
nor U27378 (N_27378,N_26591,N_26981);
and U27379 (N_27379,N_26555,N_26776);
or U27380 (N_27380,N_26536,N_26740);
or U27381 (N_27381,N_26993,N_26990);
nor U27382 (N_27382,N_26670,N_26557);
and U27383 (N_27383,N_26499,N_26917);
nor U27384 (N_27384,N_26754,N_26778);
or U27385 (N_27385,N_26807,N_26535);
nor U27386 (N_27386,N_26584,N_26461);
or U27387 (N_27387,N_26835,N_26783);
and U27388 (N_27388,N_26920,N_26434);
and U27389 (N_27389,N_26494,N_26452);
nand U27390 (N_27390,N_26939,N_26914);
xnor U27391 (N_27391,N_26522,N_26504);
nor U27392 (N_27392,N_26584,N_26485);
and U27393 (N_27393,N_26426,N_26911);
nor U27394 (N_27394,N_26658,N_26876);
or U27395 (N_27395,N_26857,N_26984);
nand U27396 (N_27396,N_26990,N_26460);
and U27397 (N_27397,N_26857,N_26992);
nor U27398 (N_27398,N_26433,N_26436);
or U27399 (N_27399,N_26991,N_26735);
nand U27400 (N_27400,N_26683,N_26606);
nand U27401 (N_27401,N_26516,N_26715);
or U27402 (N_27402,N_26621,N_26530);
xnor U27403 (N_27403,N_26848,N_26670);
nor U27404 (N_27404,N_26562,N_26894);
nand U27405 (N_27405,N_26763,N_26949);
or U27406 (N_27406,N_26649,N_26561);
or U27407 (N_27407,N_26601,N_26481);
or U27408 (N_27408,N_26457,N_26506);
or U27409 (N_27409,N_26590,N_26719);
nor U27410 (N_27410,N_26597,N_26969);
nand U27411 (N_27411,N_26750,N_26696);
or U27412 (N_27412,N_26473,N_26642);
nor U27413 (N_27413,N_26455,N_26791);
nand U27414 (N_27414,N_26623,N_26927);
nand U27415 (N_27415,N_26457,N_26805);
nand U27416 (N_27416,N_26805,N_26883);
nand U27417 (N_27417,N_26481,N_26651);
and U27418 (N_27418,N_26511,N_26579);
nand U27419 (N_27419,N_26658,N_26962);
or U27420 (N_27420,N_26614,N_26933);
nand U27421 (N_27421,N_26931,N_26674);
and U27422 (N_27422,N_26413,N_26841);
or U27423 (N_27423,N_26560,N_26844);
nand U27424 (N_27424,N_26487,N_26947);
nand U27425 (N_27425,N_26845,N_26998);
xnor U27426 (N_27426,N_26584,N_26842);
nor U27427 (N_27427,N_26434,N_26799);
or U27428 (N_27428,N_26913,N_26943);
xnor U27429 (N_27429,N_26821,N_26914);
and U27430 (N_27430,N_26900,N_26518);
or U27431 (N_27431,N_26805,N_26747);
nand U27432 (N_27432,N_26697,N_26984);
nor U27433 (N_27433,N_26581,N_26968);
nor U27434 (N_27434,N_26492,N_26584);
xor U27435 (N_27435,N_26565,N_26739);
nor U27436 (N_27436,N_26859,N_26855);
nand U27437 (N_27437,N_26444,N_26807);
or U27438 (N_27438,N_26523,N_26813);
and U27439 (N_27439,N_26919,N_26943);
nand U27440 (N_27440,N_26842,N_26913);
or U27441 (N_27441,N_26923,N_26417);
and U27442 (N_27442,N_26627,N_26599);
and U27443 (N_27443,N_26888,N_26493);
and U27444 (N_27444,N_26718,N_26955);
nor U27445 (N_27445,N_26535,N_26628);
nand U27446 (N_27446,N_26517,N_26523);
or U27447 (N_27447,N_26663,N_26639);
nand U27448 (N_27448,N_26437,N_26733);
xnor U27449 (N_27449,N_26919,N_26896);
or U27450 (N_27450,N_26527,N_26864);
nor U27451 (N_27451,N_26440,N_26454);
or U27452 (N_27452,N_26747,N_26460);
nand U27453 (N_27453,N_26470,N_26767);
and U27454 (N_27454,N_26883,N_26885);
nand U27455 (N_27455,N_26524,N_26531);
and U27456 (N_27456,N_26638,N_26693);
nand U27457 (N_27457,N_26703,N_26907);
nand U27458 (N_27458,N_26766,N_26754);
nor U27459 (N_27459,N_26847,N_26697);
or U27460 (N_27460,N_26907,N_26716);
and U27461 (N_27461,N_26963,N_26797);
and U27462 (N_27462,N_26924,N_26663);
or U27463 (N_27463,N_26765,N_26994);
xnor U27464 (N_27464,N_26479,N_26791);
nor U27465 (N_27465,N_26960,N_26734);
nor U27466 (N_27466,N_26943,N_26929);
or U27467 (N_27467,N_26742,N_26710);
nand U27468 (N_27468,N_26432,N_26590);
and U27469 (N_27469,N_26905,N_26904);
or U27470 (N_27470,N_26798,N_26684);
xor U27471 (N_27471,N_26736,N_26498);
nor U27472 (N_27472,N_26469,N_26611);
or U27473 (N_27473,N_26461,N_26986);
or U27474 (N_27474,N_26583,N_26932);
or U27475 (N_27475,N_26618,N_26643);
and U27476 (N_27476,N_26628,N_26810);
or U27477 (N_27477,N_26662,N_26675);
or U27478 (N_27478,N_26684,N_26531);
nand U27479 (N_27479,N_26907,N_26932);
nand U27480 (N_27480,N_26616,N_26567);
nor U27481 (N_27481,N_26734,N_26627);
or U27482 (N_27482,N_26809,N_26474);
nor U27483 (N_27483,N_26885,N_26416);
and U27484 (N_27484,N_26704,N_26850);
nor U27485 (N_27485,N_26796,N_26697);
or U27486 (N_27486,N_26640,N_26923);
or U27487 (N_27487,N_26410,N_26542);
nand U27488 (N_27488,N_26651,N_26642);
and U27489 (N_27489,N_26941,N_26878);
or U27490 (N_27490,N_26519,N_26458);
nand U27491 (N_27491,N_26696,N_26704);
nand U27492 (N_27492,N_26433,N_26484);
nand U27493 (N_27493,N_26822,N_26649);
nand U27494 (N_27494,N_26656,N_26866);
or U27495 (N_27495,N_26475,N_26601);
and U27496 (N_27496,N_26552,N_26934);
or U27497 (N_27497,N_26971,N_26498);
or U27498 (N_27498,N_26984,N_26930);
nand U27499 (N_27499,N_26457,N_26748);
nand U27500 (N_27500,N_26840,N_26789);
xnor U27501 (N_27501,N_26983,N_26721);
nor U27502 (N_27502,N_26720,N_26515);
xor U27503 (N_27503,N_26812,N_26846);
nor U27504 (N_27504,N_26795,N_26782);
and U27505 (N_27505,N_26716,N_26646);
nor U27506 (N_27506,N_26765,N_26670);
nand U27507 (N_27507,N_26860,N_26521);
or U27508 (N_27508,N_26811,N_26996);
and U27509 (N_27509,N_26904,N_26751);
and U27510 (N_27510,N_26751,N_26697);
and U27511 (N_27511,N_26472,N_26548);
or U27512 (N_27512,N_26483,N_26861);
and U27513 (N_27513,N_26779,N_26706);
and U27514 (N_27514,N_26503,N_26868);
or U27515 (N_27515,N_26950,N_26495);
xor U27516 (N_27516,N_26416,N_26843);
nor U27517 (N_27517,N_26440,N_26546);
nand U27518 (N_27518,N_26489,N_26892);
and U27519 (N_27519,N_26736,N_26597);
nand U27520 (N_27520,N_26467,N_26984);
xor U27521 (N_27521,N_26631,N_26656);
nand U27522 (N_27522,N_26662,N_26641);
xor U27523 (N_27523,N_26713,N_26978);
nor U27524 (N_27524,N_26574,N_26529);
nor U27525 (N_27525,N_26406,N_26796);
and U27526 (N_27526,N_26524,N_26912);
nor U27527 (N_27527,N_26577,N_26583);
nand U27528 (N_27528,N_26698,N_26608);
nand U27529 (N_27529,N_26703,N_26454);
and U27530 (N_27530,N_26784,N_26887);
nand U27531 (N_27531,N_26903,N_26791);
nand U27532 (N_27532,N_26691,N_26884);
nor U27533 (N_27533,N_26430,N_26571);
nor U27534 (N_27534,N_26906,N_26624);
nand U27535 (N_27535,N_26748,N_26912);
nor U27536 (N_27536,N_26422,N_26541);
nor U27537 (N_27537,N_26582,N_26958);
or U27538 (N_27538,N_26507,N_26814);
nand U27539 (N_27539,N_26928,N_26895);
or U27540 (N_27540,N_26411,N_26562);
xnor U27541 (N_27541,N_26524,N_26977);
or U27542 (N_27542,N_26705,N_26548);
nor U27543 (N_27543,N_26983,N_26514);
or U27544 (N_27544,N_26616,N_26795);
nor U27545 (N_27545,N_26604,N_26885);
nand U27546 (N_27546,N_26557,N_26872);
and U27547 (N_27547,N_26939,N_26411);
or U27548 (N_27548,N_26403,N_26423);
nand U27549 (N_27549,N_26975,N_26995);
xor U27550 (N_27550,N_26816,N_26893);
or U27551 (N_27551,N_26640,N_26733);
nor U27552 (N_27552,N_26421,N_26673);
and U27553 (N_27553,N_26674,N_26878);
or U27554 (N_27554,N_26588,N_26684);
nand U27555 (N_27555,N_26650,N_26501);
nand U27556 (N_27556,N_26615,N_26495);
and U27557 (N_27557,N_26465,N_26656);
nand U27558 (N_27558,N_26458,N_26676);
or U27559 (N_27559,N_26552,N_26701);
and U27560 (N_27560,N_26597,N_26573);
or U27561 (N_27561,N_26932,N_26725);
and U27562 (N_27562,N_26519,N_26581);
and U27563 (N_27563,N_26931,N_26836);
or U27564 (N_27564,N_26933,N_26958);
nand U27565 (N_27565,N_26416,N_26785);
nand U27566 (N_27566,N_26807,N_26907);
nor U27567 (N_27567,N_26570,N_26618);
and U27568 (N_27568,N_26479,N_26676);
nand U27569 (N_27569,N_26963,N_26869);
or U27570 (N_27570,N_26769,N_26968);
nand U27571 (N_27571,N_26463,N_26790);
xor U27572 (N_27572,N_26939,N_26833);
nor U27573 (N_27573,N_26582,N_26459);
and U27574 (N_27574,N_26464,N_26920);
and U27575 (N_27575,N_26833,N_26742);
or U27576 (N_27576,N_26949,N_26582);
nand U27577 (N_27577,N_26766,N_26868);
and U27578 (N_27578,N_26924,N_26987);
and U27579 (N_27579,N_26569,N_26657);
or U27580 (N_27580,N_26594,N_26866);
xor U27581 (N_27581,N_26682,N_26661);
or U27582 (N_27582,N_26460,N_26736);
or U27583 (N_27583,N_26641,N_26499);
xor U27584 (N_27584,N_26444,N_26476);
and U27585 (N_27585,N_26808,N_26749);
or U27586 (N_27586,N_26635,N_26872);
and U27587 (N_27587,N_26865,N_26488);
nand U27588 (N_27588,N_26732,N_26893);
nand U27589 (N_27589,N_26913,N_26898);
and U27590 (N_27590,N_26911,N_26753);
or U27591 (N_27591,N_26926,N_26464);
nand U27592 (N_27592,N_26514,N_26511);
xnor U27593 (N_27593,N_26503,N_26635);
and U27594 (N_27594,N_26549,N_26981);
xnor U27595 (N_27595,N_26838,N_26723);
xor U27596 (N_27596,N_26938,N_26648);
and U27597 (N_27597,N_26584,N_26940);
xor U27598 (N_27598,N_26500,N_26548);
and U27599 (N_27599,N_26839,N_26581);
nand U27600 (N_27600,N_27378,N_27434);
nor U27601 (N_27601,N_27126,N_27221);
or U27602 (N_27602,N_27147,N_27492);
or U27603 (N_27603,N_27171,N_27174);
nand U27604 (N_27604,N_27482,N_27183);
nand U27605 (N_27605,N_27359,N_27481);
nor U27606 (N_27606,N_27440,N_27450);
or U27607 (N_27607,N_27494,N_27089);
nor U27608 (N_27608,N_27417,N_27239);
and U27609 (N_27609,N_27069,N_27556);
nor U27610 (N_27610,N_27531,N_27118);
and U27611 (N_27611,N_27389,N_27567);
and U27612 (N_27612,N_27581,N_27051);
and U27613 (N_27613,N_27025,N_27369);
and U27614 (N_27614,N_27011,N_27255);
xnor U27615 (N_27615,N_27114,N_27224);
nand U27616 (N_27616,N_27304,N_27329);
nor U27617 (N_27617,N_27112,N_27148);
and U27618 (N_27618,N_27274,N_27530);
or U27619 (N_27619,N_27280,N_27008);
nand U27620 (N_27620,N_27220,N_27299);
or U27621 (N_27621,N_27105,N_27132);
nor U27622 (N_27622,N_27419,N_27334);
nand U27623 (N_27623,N_27545,N_27431);
nor U27624 (N_27624,N_27548,N_27111);
or U27625 (N_27625,N_27381,N_27117);
nor U27626 (N_27626,N_27475,N_27289);
or U27627 (N_27627,N_27321,N_27598);
nand U27628 (N_27628,N_27091,N_27507);
xor U27629 (N_27629,N_27367,N_27028);
and U27630 (N_27630,N_27133,N_27311);
or U27631 (N_27631,N_27356,N_27511);
and U27632 (N_27632,N_27101,N_27084);
nand U27633 (N_27633,N_27582,N_27045);
xnor U27634 (N_27634,N_27169,N_27570);
and U27635 (N_27635,N_27514,N_27443);
nor U27636 (N_27636,N_27000,N_27563);
and U27637 (N_27637,N_27486,N_27070);
and U27638 (N_27638,N_27216,N_27064);
or U27639 (N_27639,N_27517,N_27022);
and U27640 (N_27640,N_27013,N_27504);
and U27641 (N_27641,N_27577,N_27116);
or U27642 (N_27642,N_27003,N_27516);
nor U27643 (N_27643,N_27525,N_27081);
nor U27644 (N_27644,N_27290,N_27226);
and U27645 (N_27645,N_27241,N_27146);
nor U27646 (N_27646,N_27217,N_27341);
xor U27647 (N_27647,N_27223,N_27250);
or U27648 (N_27648,N_27184,N_27115);
or U27649 (N_27649,N_27319,N_27015);
nor U27650 (N_27650,N_27547,N_27447);
nand U27651 (N_27651,N_27138,N_27455);
nand U27652 (N_27652,N_27100,N_27033);
and U27653 (N_27653,N_27576,N_27420);
or U27654 (N_27654,N_27142,N_27264);
nor U27655 (N_27655,N_27400,N_27303);
or U27656 (N_27656,N_27057,N_27578);
nor U27657 (N_27657,N_27103,N_27230);
and U27658 (N_27658,N_27181,N_27421);
or U27659 (N_27659,N_27054,N_27506);
nand U27660 (N_27660,N_27108,N_27365);
or U27661 (N_27661,N_27353,N_27173);
nand U27662 (N_27662,N_27083,N_27058);
and U27663 (N_27663,N_27266,N_27515);
and U27664 (N_27664,N_27043,N_27235);
nor U27665 (N_27665,N_27408,N_27595);
nor U27666 (N_27666,N_27305,N_27466);
and U27667 (N_27667,N_27096,N_27134);
nand U27668 (N_27668,N_27212,N_27010);
and U27669 (N_27669,N_27277,N_27553);
nor U27670 (N_27670,N_27448,N_27564);
and U27671 (N_27671,N_27491,N_27292);
nor U27672 (N_27672,N_27219,N_27565);
or U27673 (N_27673,N_27210,N_27388);
nand U27674 (N_27674,N_27288,N_27037);
and U27675 (N_27675,N_27035,N_27415);
xor U27676 (N_27676,N_27442,N_27205);
nand U27677 (N_27677,N_27143,N_27071);
nor U27678 (N_27678,N_27554,N_27177);
or U27679 (N_27679,N_27426,N_27179);
nand U27680 (N_27680,N_27485,N_27480);
and U27681 (N_27681,N_27263,N_27055);
nor U27682 (N_27682,N_27123,N_27272);
and U27683 (N_27683,N_27469,N_27549);
nor U27684 (N_27684,N_27049,N_27159);
nor U27685 (N_27685,N_27544,N_27286);
nand U27686 (N_27686,N_27167,N_27537);
nor U27687 (N_27687,N_27457,N_27413);
and U27688 (N_27688,N_27462,N_27453);
or U27689 (N_27689,N_27374,N_27393);
or U27690 (N_27690,N_27436,N_27340);
nor U27691 (N_27691,N_27063,N_27380);
or U27692 (N_27692,N_27501,N_27354);
nor U27693 (N_27693,N_27467,N_27360);
xnor U27694 (N_27694,N_27430,N_27092);
xnor U27695 (N_27695,N_27026,N_27307);
nand U27696 (N_27696,N_27519,N_27158);
or U27697 (N_27697,N_27362,N_27074);
nand U27698 (N_27698,N_27505,N_27327);
and U27699 (N_27699,N_27445,N_27464);
nor U27700 (N_27700,N_27468,N_27558);
and U27701 (N_27701,N_27317,N_27416);
xor U27702 (N_27702,N_27366,N_27594);
nor U27703 (N_27703,N_27247,N_27282);
and U27704 (N_27704,N_27082,N_27301);
nand U27705 (N_27705,N_27076,N_27532);
and U27706 (N_27706,N_27170,N_27093);
xor U27707 (N_27707,N_27333,N_27031);
and U27708 (N_27708,N_27155,N_27522);
nand U27709 (N_27709,N_27489,N_27017);
and U27710 (N_27710,N_27348,N_27561);
xor U27711 (N_27711,N_27542,N_27451);
or U27712 (N_27712,N_27399,N_27568);
nand U27713 (N_27713,N_27509,N_27152);
and U27714 (N_27714,N_27499,N_27056);
xnor U27715 (N_27715,N_27193,N_27271);
and U27716 (N_27716,N_27463,N_27488);
nand U27717 (N_27717,N_27175,N_27345);
nor U27718 (N_27718,N_27386,N_27222);
xor U27719 (N_27719,N_27300,N_27465);
nand U27720 (N_27720,N_27346,N_27551);
or U27721 (N_27721,N_27039,N_27336);
and U27722 (N_27722,N_27127,N_27014);
nor U27723 (N_27723,N_27543,N_27141);
nand U27724 (N_27724,N_27176,N_27232);
or U27725 (N_27725,N_27361,N_27569);
or U27726 (N_27726,N_27145,N_27166);
nand U27727 (N_27727,N_27005,N_27358);
or U27728 (N_27728,N_27429,N_27294);
or U27729 (N_27729,N_27200,N_27207);
nor U27730 (N_27730,N_27363,N_27552);
nand U27731 (N_27731,N_27587,N_27113);
or U27732 (N_27732,N_27061,N_27086);
or U27733 (N_27733,N_27237,N_27298);
or U27734 (N_27734,N_27262,N_27023);
or U27735 (N_27735,N_27187,N_27487);
and U27736 (N_27736,N_27573,N_27376);
nand U27737 (N_27737,N_27036,N_27244);
nor U27738 (N_27738,N_27593,N_27052);
nand U27739 (N_27739,N_27240,N_27483);
and U27740 (N_27740,N_27287,N_27119);
and U27741 (N_27741,N_27323,N_27372);
or U27742 (N_27742,N_27382,N_27371);
or U27743 (N_27743,N_27104,N_27225);
nand U27744 (N_27744,N_27161,N_27414);
nand U27745 (N_27745,N_27208,N_27528);
xnor U27746 (N_27746,N_27477,N_27314);
nand U27747 (N_27747,N_27392,N_27053);
nor U27748 (N_27748,N_27461,N_27197);
nor U27749 (N_27749,N_27163,N_27559);
and U27750 (N_27750,N_27546,N_27202);
nor U27751 (N_27751,N_27107,N_27410);
xor U27752 (N_27752,N_27347,N_27256);
or U27753 (N_27753,N_27047,N_27330);
and U27754 (N_27754,N_27164,N_27490);
nand U27755 (N_27755,N_27030,N_27526);
xnor U27756 (N_27756,N_27059,N_27557);
nand U27757 (N_27757,N_27048,N_27404);
or U27758 (N_27758,N_27018,N_27066);
nand U27759 (N_27759,N_27215,N_27097);
and U27760 (N_27760,N_27131,N_27213);
xnor U27761 (N_27761,N_27186,N_27050);
or U27762 (N_27762,N_27580,N_27398);
nand U27763 (N_27763,N_27099,N_27273);
nor U27764 (N_27764,N_27253,N_27510);
nor U27765 (N_27765,N_27579,N_27407);
xor U27766 (N_27766,N_27065,N_27078);
nor U27767 (N_27767,N_27206,N_27428);
and U27768 (N_27768,N_27342,N_27395);
or U27769 (N_27769,N_27586,N_27021);
xor U27770 (N_27770,N_27332,N_27503);
and U27771 (N_27771,N_27328,N_27007);
nand U27772 (N_27772,N_27373,N_27535);
and U27773 (N_27773,N_27384,N_27150);
nand U27774 (N_27774,N_27474,N_27275);
xnor U27775 (N_27775,N_27269,N_27302);
and U27776 (N_27776,N_27009,N_27585);
nor U27777 (N_27777,N_27427,N_27194);
nand U27778 (N_27778,N_27137,N_27077);
nor U27779 (N_27779,N_27596,N_27315);
nor U27780 (N_27780,N_27479,N_27438);
or U27781 (N_27781,N_27344,N_27460);
or U27782 (N_27782,N_27368,N_27513);
or U27783 (N_27783,N_27153,N_27527);
or U27784 (N_27784,N_27297,N_27204);
nand U27785 (N_27785,N_27533,N_27095);
or U27786 (N_27786,N_27180,N_27238);
nand U27787 (N_27787,N_27029,N_27560);
or U27788 (N_27788,N_27397,N_27004);
nor U27789 (N_27789,N_27182,N_27012);
or U27790 (N_27790,N_27523,N_27080);
nand U27791 (N_27791,N_27521,N_27040);
nand U27792 (N_27792,N_27098,N_27350);
and U27793 (N_27793,N_27377,N_27038);
nor U27794 (N_27794,N_27476,N_27190);
nand U27795 (N_27795,N_27437,N_27245);
and U27796 (N_27796,N_27394,N_27090);
or U27797 (N_27797,N_27572,N_27418);
or U27798 (N_27798,N_27458,N_27518);
and U27799 (N_27799,N_27102,N_27391);
nor U27800 (N_27800,N_27062,N_27188);
and U27801 (N_27801,N_27313,N_27191);
and U27802 (N_27802,N_27067,N_27046);
and U27803 (N_27803,N_27379,N_27075);
nor U27804 (N_27804,N_27144,N_27320);
and U27805 (N_27805,N_27267,N_27259);
nor U27806 (N_27806,N_27343,N_27575);
and U27807 (N_27807,N_27497,N_27122);
or U27808 (N_27808,N_27409,N_27094);
and U27809 (N_27809,N_27540,N_27157);
nand U27810 (N_27810,N_27214,N_27261);
or U27811 (N_27811,N_27441,N_27493);
or U27812 (N_27812,N_27258,N_27162);
and U27813 (N_27813,N_27584,N_27251);
nor U27814 (N_27814,N_27550,N_27411);
xor U27815 (N_27815,N_27425,N_27592);
nand U27816 (N_27816,N_27041,N_27281);
or U27817 (N_27817,N_27452,N_27339);
and U27818 (N_27818,N_27402,N_27234);
xnor U27819 (N_27819,N_27032,N_27423);
and U27820 (N_27820,N_27591,N_27412);
nand U27821 (N_27821,N_27284,N_27308);
and U27822 (N_27822,N_27120,N_27279);
and U27823 (N_27823,N_27165,N_27446);
nand U27824 (N_27824,N_27338,N_27405);
nor U27825 (N_27825,N_27471,N_27472);
xnor U27826 (N_27826,N_27268,N_27079);
and U27827 (N_27827,N_27529,N_27498);
nor U27828 (N_27828,N_27484,N_27020);
and U27829 (N_27829,N_27588,N_27270);
xnor U27830 (N_27830,N_27199,N_27072);
or U27831 (N_27831,N_27473,N_27512);
nand U27832 (N_27832,N_27125,N_27396);
nand U27833 (N_27833,N_27508,N_27589);
xnor U27834 (N_27834,N_27088,N_27265);
nor U27835 (N_27835,N_27424,N_27306);
nor U27836 (N_27836,N_27185,N_27502);
nor U27837 (N_27837,N_27370,N_27016);
or U27838 (N_27838,N_27172,N_27325);
and U27839 (N_27839,N_27326,N_27283);
nor U27840 (N_27840,N_27168,N_27231);
or U27841 (N_27841,N_27324,N_27390);
or U27842 (N_27842,N_27121,N_27406);
or U27843 (N_27843,N_27566,N_27439);
nand U27844 (N_27844,N_27583,N_27139);
or U27845 (N_27845,N_27478,N_27312);
nor U27846 (N_27846,N_27401,N_27236);
xor U27847 (N_27847,N_27495,N_27524);
or U27848 (N_27848,N_27432,N_27500);
and U27849 (N_27849,N_27135,N_27073);
nand U27850 (N_27850,N_27385,N_27001);
or U27851 (N_27851,N_27278,N_27599);
or U27852 (N_27852,N_27110,N_27140);
and U27853 (N_27853,N_27571,N_27192);
and U27854 (N_27854,N_27590,N_27087);
nor U27855 (N_27855,N_27189,N_27019);
nand U27856 (N_27856,N_27209,N_27203);
nor U27857 (N_27857,N_27276,N_27496);
xor U27858 (N_27858,N_27433,N_27296);
or U27859 (N_27859,N_27106,N_27211);
xnor U27860 (N_27860,N_27160,N_27124);
or U27861 (N_27861,N_27309,N_27252);
or U27862 (N_27862,N_27196,N_27316);
and U27863 (N_27863,N_27295,N_27006);
xor U27864 (N_27864,N_27352,N_27539);
nand U27865 (N_27865,N_27002,N_27248);
nor U27866 (N_27866,N_27198,N_27027);
nor U27867 (N_27867,N_27034,N_27291);
nor U27868 (N_27868,N_27470,N_27357);
nor U27869 (N_27869,N_27024,N_27422);
and U27870 (N_27870,N_27154,N_27534);
nand U27871 (N_27871,N_27129,N_27136);
and U27872 (N_27872,N_27536,N_27068);
and U27873 (N_27873,N_27310,N_27227);
nor U27874 (N_27874,N_27156,N_27403);
and U27875 (N_27875,N_27322,N_27337);
nand U27876 (N_27876,N_27257,N_27130);
nand U27877 (N_27877,N_27042,N_27454);
nor U27878 (N_27878,N_27555,N_27254);
xnor U27879 (N_27879,N_27355,N_27201);
nand U27880 (N_27880,N_27318,N_27044);
and U27881 (N_27881,N_27246,N_27538);
nand U27882 (N_27882,N_27597,N_27520);
or U27883 (N_27883,N_27260,N_27085);
nand U27884 (N_27884,N_27149,N_27228);
or U27885 (N_27885,N_27249,N_27229);
nand U27886 (N_27886,N_27335,N_27364);
and U27887 (N_27887,N_27233,N_27151);
or U27888 (N_27888,N_27178,N_27349);
nor U27889 (N_27889,N_27562,N_27218);
and U27890 (N_27890,N_27387,N_27060);
and U27891 (N_27891,N_27242,N_27449);
nand U27892 (N_27892,N_27375,N_27541);
nor U27893 (N_27893,N_27243,N_27351);
or U27894 (N_27894,N_27293,N_27574);
or U27895 (N_27895,N_27285,N_27109);
or U27896 (N_27896,N_27456,N_27383);
nand U27897 (N_27897,N_27128,N_27444);
or U27898 (N_27898,N_27331,N_27195);
nor U27899 (N_27899,N_27435,N_27459);
and U27900 (N_27900,N_27536,N_27599);
and U27901 (N_27901,N_27550,N_27150);
and U27902 (N_27902,N_27068,N_27042);
nor U27903 (N_27903,N_27545,N_27469);
nand U27904 (N_27904,N_27227,N_27518);
nand U27905 (N_27905,N_27015,N_27355);
nor U27906 (N_27906,N_27136,N_27338);
or U27907 (N_27907,N_27227,N_27393);
nand U27908 (N_27908,N_27444,N_27521);
nand U27909 (N_27909,N_27115,N_27596);
nand U27910 (N_27910,N_27101,N_27584);
and U27911 (N_27911,N_27167,N_27081);
nor U27912 (N_27912,N_27460,N_27455);
nor U27913 (N_27913,N_27086,N_27236);
and U27914 (N_27914,N_27072,N_27303);
nor U27915 (N_27915,N_27479,N_27074);
nor U27916 (N_27916,N_27128,N_27271);
nand U27917 (N_27917,N_27278,N_27561);
nor U27918 (N_27918,N_27472,N_27073);
nor U27919 (N_27919,N_27380,N_27530);
and U27920 (N_27920,N_27247,N_27343);
or U27921 (N_27921,N_27531,N_27028);
nor U27922 (N_27922,N_27390,N_27129);
nor U27923 (N_27923,N_27144,N_27329);
and U27924 (N_27924,N_27028,N_27582);
nor U27925 (N_27925,N_27056,N_27528);
and U27926 (N_27926,N_27318,N_27241);
nor U27927 (N_27927,N_27023,N_27502);
or U27928 (N_27928,N_27054,N_27257);
and U27929 (N_27929,N_27532,N_27559);
nor U27930 (N_27930,N_27365,N_27196);
and U27931 (N_27931,N_27345,N_27327);
nor U27932 (N_27932,N_27552,N_27195);
nor U27933 (N_27933,N_27296,N_27122);
nand U27934 (N_27934,N_27390,N_27573);
and U27935 (N_27935,N_27078,N_27449);
nand U27936 (N_27936,N_27478,N_27495);
or U27937 (N_27937,N_27265,N_27060);
nand U27938 (N_27938,N_27100,N_27283);
or U27939 (N_27939,N_27432,N_27391);
xnor U27940 (N_27940,N_27532,N_27299);
nor U27941 (N_27941,N_27190,N_27234);
nand U27942 (N_27942,N_27576,N_27540);
xnor U27943 (N_27943,N_27225,N_27407);
or U27944 (N_27944,N_27054,N_27544);
nor U27945 (N_27945,N_27401,N_27435);
nand U27946 (N_27946,N_27076,N_27349);
and U27947 (N_27947,N_27588,N_27222);
and U27948 (N_27948,N_27452,N_27224);
nand U27949 (N_27949,N_27321,N_27536);
nor U27950 (N_27950,N_27516,N_27503);
and U27951 (N_27951,N_27098,N_27173);
xor U27952 (N_27952,N_27288,N_27570);
nand U27953 (N_27953,N_27430,N_27578);
or U27954 (N_27954,N_27403,N_27351);
and U27955 (N_27955,N_27473,N_27438);
or U27956 (N_27956,N_27492,N_27140);
nor U27957 (N_27957,N_27153,N_27195);
nand U27958 (N_27958,N_27196,N_27164);
nor U27959 (N_27959,N_27578,N_27597);
nor U27960 (N_27960,N_27459,N_27213);
nand U27961 (N_27961,N_27276,N_27597);
or U27962 (N_27962,N_27218,N_27322);
or U27963 (N_27963,N_27029,N_27203);
nor U27964 (N_27964,N_27266,N_27539);
nor U27965 (N_27965,N_27096,N_27570);
nand U27966 (N_27966,N_27573,N_27412);
xor U27967 (N_27967,N_27033,N_27426);
or U27968 (N_27968,N_27046,N_27140);
nand U27969 (N_27969,N_27324,N_27163);
and U27970 (N_27970,N_27133,N_27252);
or U27971 (N_27971,N_27518,N_27530);
and U27972 (N_27972,N_27175,N_27573);
nor U27973 (N_27973,N_27587,N_27512);
or U27974 (N_27974,N_27344,N_27361);
and U27975 (N_27975,N_27215,N_27582);
nand U27976 (N_27976,N_27327,N_27145);
and U27977 (N_27977,N_27132,N_27370);
xnor U27978 (N_27978,N_27221,N_27427);
and U27979 (N_27979,N_27512,N_27506);
nand U27980 (N_27980,N_27536,N_27453);
xor U27981 (N_27981,N_27046,N_27078);
and U27982 (N_27982,N_27456,N_27140);
or U27983 (N_27983,N_27379,N_27024);
nand U27984 (N_27984,N_27291,N_27230);
nand U27985 (N_27985,N_27250,N_27222);
nor U27986 (N_27986,N_27376,N_27265);
and U27987 (N_27987,N_27187,N_27173);
nand U27988 (N_27988,N_27294,N_27185);
nand U27989 (N_27989,N_27115,N_27326);
or U27990 (N_27990,N_27376,N_27294);
nor U27991 (N_27991,N_27017,N_27364);
xor U27992 (N_27992,N_27162,N_27299);
nand U27993 (N_27993,N_27429,N_27374);
and U27994 (N_27994,N_27570,N_27557);
or U27995 (N_27995,N_27169,N_27147);
or U27996 (N_27996,N_27424,N_27282);
nor U27997 (N_27997,N_27535,N_27226);
or U27998 (N_27998,N_27559,N_27136);
nor U27999 (N_27999,N_27499,N_27280);
nand U28000 (N_28000,N_27294,N_27470);
xor U28001 (N_28001,N_27185,N_27211);
xnor U28002 (N_28002,N_27326,N_27537);
nand U28003 (N_28003,N_27209,N_27408);
or U28004 (N_28004,N_27028,N_27322);
nand U28005 (N_28005,N_27466,N_27161);
or U28006 (N_28006,N_27365,N_27040);
nand U28007 (N_28007,N_27242,N_27583);
nor U28008 (N_28008,N_27183,N_27591);
or U28009 (N_28009,N_27332,N_27148);
nand U28010 (N_28010,N_27123,N_27588);
nand U28011 (N_28011,N_27127,N_27346);
nand U28012 (N_28012,N_27430,N_27576);
nor U28013 (N_28013,N_27422,N_27279);
nor U28014 (N_28014,N_27510,N_27236);
nand U28015 (N_28015,N_27289,N_27002);
xor U28016 (N_28016,N_27438,N_27338);
nor U28017 (N_28017,N_27330,N_27108);
and U28018 (N_28018,N_27353,N_27484);
nand U28019 (N_28019,N_27261,N_27302);
and U28020 (N_28020,N_27177,N_27417);
and U28021 (N_28021,N_27036,N_27126);
or U28022 (N_28022,N_27032,N_27287);
nor U28023 (N_28023,N_27264,N_27277);
nand U28024 (N_28024,N_27539,N_27416);
and U28025 (N_28025,N_27095,N_27137);
and U28026 (N_28026,N_27450,N_27148);
nor U28027 (N_28027,N_27566,N_27308);
nor U28028 (N_28028,N_27350,N_27124);
and U28029 (N_28029,N_27583,N_27333);
or U28030 (N_28030,N_27376,N_27263);
nor U28031 (N_28031,N_27311,N_27196);
and U28032 (N_28032,N_27226,N_27547);
nor U28033 (N_28033,N_27216,N_27542);
or U28034 (N_28034,N_27185,N_27511);
and U28035 (N_28035,N_27253,N_27559);
nor U28036 (N_28036,N_27170,N_27353);
and U28037 (N_28037,N_27164,N_27510);
xnor U28038 (N_28038,N_27368,N_27038);
xor U28039 (N_28039,N_27249,N_27152);
nor U28040 (N_28040,N_27432,N_27514);
xnor U28041 (N_28041,N_27512,N_27024);
nor U28042 (N_28042,N_27117,N_27018);
nor U28043 (N_28043,N_27480,N_27181);
and U28044 (N_28044,N_27470,N_27522);
xor U28045 (N_28045,N_27310,N_27078);
nand U28046 (N_28046,N_27172,N_27347);
and U28047 (N_28047,N_27516,N_27099);
and U28048 (N_28048,N_27470,N_27303);
nor U28049 (N_28049,N_27022,N_27562);
nand U28050 (N_28050,N_27544,N_27140);
nor U28051 (N_28051,N_27482,N_27481);
xnor U28052 (N_28052,N_27218,N_27155);
xor U28053 (N_28053,N_27590,N_27091);
or U28054 (N_28054,N_27062,N_27514);
xor U28055 (N_28055,N_27170,N_27486);
or U28056 (N_28056,N_27423,N_27285);
nand U28057 (N_28057,N_27563,N_27434);
xnor U28058 (N_28058,N_27202,N_27182);
nand U28059 (N_28059,N_27416,N_27028);
or U28060 (N_28060,N_27382,N_27445);
or U28061 (N_28061,N_27436,N_27054);
and U28062 (N_28062,N_27021,N_27148);
or U28063 (N_28063,N_27396,N_27499);
xor U28064 (N_28064,N_27543,N_27149);
nand U28065 (N_28065,N_27057,N_27129);
nand U28066 (N_28066,N_27536,N_27003);
nor U28067 (N_28067,N_27333,N_27238);
nand U28068 (N_28068,N_27075,N_27422);
nor U28069 (N_28069,N_27277,N_27065);
or U28070 (N_28070,N_27589,N_27295);
or U28071 (N_28071,N_27118,N_27182);
and U28072 (N_28072,N_27088,N_27364);
nand U28073 (N_28073,N_27520,N_27123);
or U28074 (N_28074,N_27338,N_27560);
and U28075 (N_28075,N_27145,N_27383);
nor U28076 (N_28076,N_27403,N_27166);
nor U28077 (N_28077,N_27013,N_27563);
and U28078 (N_28078,N_27344,N_27472);
or U28079 (N_28079,N_27352,N_27498);
xnor U28080 (N_28080,N_27325,N_27460);
xnor U28081 (N_28081,N_27213,N_27149);
and U28082 (N_28082,N_27448,N_27524);
or U28083 (N_28083,N_27197,N_27326);
nand U28084 (N_28084,N_27082,N_27429);
and U28085 (N_28085,N_27380,N_27120);
nor U28086 (N_28086,N_27530,N_27331);
nor U28087 (N_28087,N_27561,N_27406);
nor U28088 (N_28088,N_27099,N_27160);
or U28089 (N_28089,N_27491,N_27569);
nor U28090 (N_28090,N_27031,N_27364);
nor U28091 (N_28091,N_27429,N_27250);
and U28092 (N_28092,N_27516,N_27091);
nand U28093 (N_28093,N_27067,N_27104);
xor U28094 (N_28094,N_27295,N_27092);
or U28095 (N_28095,N_27564,N_27579);
and U28096 (N_28096,N_27471,N_27534);
nand U28097 (N_28097,N_27486,N_27295);
xnor U28098 (N_28098,N_27432,N_27488);
and U28099 (N_28099,N_27378,N_27555);
nor U28100 (N_28100,N_27499,N_27144);
nand U28101 (N_28101,N_27295,N_27237);
xnor U28102 (N_28102,N_27176,N_27595);
or U28103 (N_28103,N_27254,N_27131);
and U28104 (N_28104,N_27064,N_27581);
nor U28105 (N_28105,N_27241,N_27430);
or U28106 (N_28106,N_27400,N_27584);
nand U28107 (N_28107,N_27247,N_27280);
nor U28108 (N_28108,N_27155,N_27200);
or U28109 (N_28109,N_27239,N_27118);
xnor U28110 (N_28110,N_27462,N_27032);
and U28111 (N_28111,N_27515,N_27420);
and U28112 (N_28112,N_27055,N_27451);
or U28113 (N_28113,N_27227,N_27165);
nor U28114 (N_28114,N_27031,N_27519);
nand U28115 (N_28115,N_27081,N_27507);
nor U28116 (N_28116,N_27516,N_27036);
nor U28117 (N_28117,N_27325,N_27401);
and U28118 (N_28118,N_27449,N_27050);
xor U28119 (N_28119,N_27124,N_27108);
and U28120 (N_28120,N_27243,N_27486);
nand U28121 (N_28121,N_27599,N_27357);
nand U28122 (N_28122,N_27555,N_27128);
xor U28123 (N_28123,N_27446,N_27325);
nand U28124 (N_28124,N_27198,N_27582);
nand U28125 (N_28125,N_27214,N_27003);
nor U28126 (N_28126,N_27026,N_27509);
or U28127 (N_28127,N_27291,N_27257);
xor U28128 (N_28128,N_27411,N_27482);
xnor U28129 (N_28129,N_27486,N_27095);
nor U28130 (N_28130,N_27563,N_27497);
and U28131 (N_28131,N_27264,N_27214);
or U28132 (N_28132,N_27186,N_27012);
or U28133 (N_28133,N_27306,N_27153);
or U28134 (N_28134,N_27288,N_27386);
and U28135 (N_28135,N_27145,N_27517);
xor U28136 (N_28136,N_27189,N_27138);
nor U28137 (N_28137,N_27509,N_27574);
or U28138 (N_28138,N_27587,N_27092);
or U28139 (N_28139,N_27062,N_27549);
and U28140 (N_28140,N_27339,N_27323);
nor U28141 (N_28141,N_27381,N_27169);
nor U28142 (N_28142,N_27307,N_27190);
nor U28143 (N_28143,N_27360,N_27242);
or U28144 (N_28144,N_27473,N_27561);
nor U28145 (N_28145,N_27106,N_27322);
nand U28146 (N_28146,N_27349,N_27042);
nor U28147 (N_28147,N_27219,N_27512);
or U28148 (N_28148,N_27471,N_27429);
and U28149 (N_28149,N_27308,N_27021);
and U28150 (N_28150,N_27171,N_27282);
or U28151 (N_28151,N_27292,N_27405);
nor U28152 (N_28152,N_27254,N_27476);
nand U28153 (N_28153,N_27203,N_27504);
or U28154 (N_28154,N_27336,N_27078);
nor U28155 (N_28155,N_27545,N_27167);
nor U28156 (N_28156,N_27156,N_27462);
nand U28157 (N_28157,N_27402,N_27205);
nor U28158 (N_28158,N_27372,N_27345);
or U28159 (N_28159,N_27589,N_27027);
or U28160 (N_28160,N_27000,N_27234);
or U28161 (N_28161,N_27550,N_27087);
and U28162 (N_28162,N_27555,N_27353);
and U28163 (N_28163,N_27039,N_27324);
nor U28164 (N_28164,N_27093,N_27585);
xor U28165 (N_28165,N_27486,N_27224);
nor U28166 (N_28166,N_27215,N_27259);
nor U28167 (N_28167,N_27302,N_27428);
nand U28168 (N_28168,N_27191,N_27384);
and U28169 (N_28169,N_27068,N_27411);
nand U28170 (N_28170,N_27498,N_27086);
nor U28171 (N_28171,N_27165,N_27342);
nand U28172 (N_28172,N_27147,N_27196);
and U28173 (N_28173,N_27047,N_27521);
xor U28174 (N_28174,N_27520,N_27031);
or U28175 (N_28175,N_27233,N_27468);
or U28176 (N_28176,N_27168,N_27408);
nor U28177 (N_28177,N_27547,N_27249);
and U28178 (N_28178,N_27263,N_27523);
nand U28179 (N_28179,N_27151,N_27495);
nand U28180 (N_28180,N_27216,N_27256);
or U28181 (N_28181,N_27091,N_27376);
nand U28182 (N_28182,N_27219,N_27540);
xnor U28183 (N_28183,N_27183,N_27327);
nor U28184 (N_28184,N_27400,N_27225);
and U28185 (N_28185,N_27449,N_27584);
or U28186 (N_28186,N_27310,N_27098);
or U28187 (N_28187,N_27515,N_27081);
and U28188 (N_28188,N_27329,N_27162);
or U28189 (N_28189,N_27336,N_27197);
nand U28190 (N_28190,N_27125,N_27213);
or U28191 (N_28191,N_27289,N_27075);
or U28192 (N_28192,N_27523,N_27421);
nand U28193 (N_28193,N_27192,N_27202);
nor U28194 (N_28194,N_27154,N_27258);
nor U28195 (N_28195,N_27342,N_27517);
nor U28196 (N_28196,N_27189,N_27541);
or U28197 (N_28197,N_27358,N_27083);
nor U28198 (N_28198,N_27283,N_27567);
nand U28199 (N_28199,N_27066,N_27535);
xor U28200 (N_28200,N_27819,N_27958);
nand U28201 (N_28201,N_28029,N_28125);
and U28202 (N_28202,N_28142,N_27658);
or U28203 (N_28203,N_28134,N_27681);
nor U28204 (N_28204,N_27607,N_27817);
and U28205 (N_28205,N_27999,N_27638);
nand U28206 (N_28206,N_28147,N_27875);
nand U28207 (N_28207,N_27617,N_27651);
nand U28208 (N_28208,N_27858,N_27785);
or U28209 (N_28209,N_28180,N_27720);
nand U28210 (N_28210,N_28126,N_27864);
and U28211 (N_28211,N_27989,N_27622);
nor U28212 (N_28212,N_28038,N_27884);
nand U28213 (N_28213,N_27956,N_27769);
or U28214 (N_28214,N_28163,N_27692);
nor U28215 (N_28215,N_27805,N_27993);
nand U28216 (N_28216,N_27994,N_28064);
and U28217 (N_28217,N_27978,N_27827);
or U28218 (N_28218,N_27948,N_27820);
and U28219 (N_28219,N_27867,N_28085);
and U28220 (N_28220,N_27639,N_28111);
xnor U28221 (N_28221,N_27961,N_28196);
and U28222 (N_28222,N_28004,N_27979);
or U28223 (N_28223,N_28195,N_27871);
nand U28224 (N_28224,N_27739,N_28159);
and U28225 (N_28225,N_27753,N_28103);
nor U28226 (N_28226,N_28054,N_28059);
nor U28227 (N_28227,N_27945,N_28089);
xor U28228 (N_28228,N_28137,N_27756);
and U28229 (N_28229,N_27755,N_27888);
and U28230 (N_28230,N_27667,N_27934);
xnor U28231 (N_28231,N_27759,N_28181);
nand U28232 (N_28232,N_27841,N_27822);
nand U28233 (N_28233,N_27840,N_28068);
or U28234 (N_28234,N_27851,N_27665);
or U28235 (N_28235,N_27828,N_27644);
and U28236 (N_28236,N_27626,N_28176);
nor U28237 (N_28237,N_27904,N_27936);
nor U28238 (N_28238,N_27842,N_27605);
nor U28239 (N_28239,N_27895,N_28003);
nor U28240 (N_28240,N_27923,N_28072);
and U28241 (N_28241,N_28047,N_27619);
xnor U28242 (N_28242,N_27866,N_27992);
nand U28243 (N_28243,N_27959,N_27854);
nor U28244 (N_28244,N_27793,N_28030);
nor U28245 (N_28245,N_27809,N_28182);
nand U28246 (N_28246,N_27621,N_28185);
nor U28247 (N_28247,N_27761,N_28136);
and U28248 (N_28248,N_27786,N_28178);
xnor U28249 (N_28249,N_28024,N_27876);
nor U28250 (N_28250,N_28048,N_27971);
or U28251 (N_28251,N_28110,N_27608);
or U28252 (N_28252,N_27660,N_27729);
or U28253 (N_28253,N_28012,N_27987);
or U28254 (N_28254,N_28148,N_28073);
nand U28255 (N_28255,N_27612,N_27799);
or U28256 (N_28256,N_28013,N_27614);
or U28257 (N_28257,N_27630,N_28162);
nor U28258 (N_28258,N_27661,N_27913);
nor U28259 (N_28259,N_27616,N_27790);
xor U28260 (N_28260,N_28139,N_28133);
and U28261 (N_28261,N_27878,N_28094);
or U28262 (N_28262,N_27779,N_27650);
nand U28263 (N_28263,N_27758,N_27812);
or U28264 (N_28264,N_27816,N_27982);
nor U28265 (N_28265,N_27601,N_27833);
nor U28266 (N_28266,N_27736,N_28143);
and U28267 (N_28267,N_27670,N_28160);
or U28268 (N_28268,N_28018,N_27767);
nor U28269 (N_28269,N_27821,N_28077);
nor U28270 (N_28270,N_28067,N_28005);
and U28271 (N_28271,N_27776,N_28192);
or U28272 (N_28272,N_27922,N_27707);
and U28273 (N_28273,N_27659,N_28141);
nand U28274 (N_28274,N_27764,N_27990);
and U28275 (N_28275,N_27818,N_27929);
nor U28276 (N_28276,N_28023,N_27883);
and U28277 (N_28277,N_27643,N_28131);
nor U28278 (N_28278,N_27868,N_27916);
and U28279 (N_28279,N_27724,N_27698);
or U28280 (N_28280,N_28001,N_27918);
and U28281 (N_28281,N_27957,N_27711);
or U28282 (N_28282,N_27834,N_28198);
or U28283 (N_28283,N_27832,N_27733);
or U28284 (N_28284,N_27708,N_27728);
and U28285 (N_28285,N_28155,N_27852);
nor U28286 (N_28286,N_27632,N_28123);
nor U28287 (N_28287,N_27750,N_27940);
xor U28288 (N_28288,N_28091,N_27985);
and U28289 (N_28289,N_28172,N_28145);
nand U28290 (N_28290,N_27682,N_27705);
xor U28291 (N_28291,N_28154,N_27772);
or U28292 (N_28292,N_28071,N_27843);
nor U28293 (N_28293,N_27977,N_27653);
nand U28294 (N_28294,N_28149,N_27932);
xor U28295 (N_28295,N_28042,N_27810);
or U28296 (N_28296,N_27796,N_28086);
nor U28297 (N_28297,N_27893,N_27966);
or U28298 (N_28298,N_28122,N_27835);
nor U28299 (N_28299,N_27860,N_27901);
nor U28300 (N_28300,N_27873,N_27775);
or U28301 (N_28301,N_27748,N_27732);
nor U28302 (N_28302,N_27807,N_28112);
xor U28303 (N_28303,N_27642,N_27754);
xnor U28304 (N_28304,N_28020,N_27791);
nor U28305 (N_28305,N_28120,N_27611);
or U28306 (N_28306,N_27896,N_27766);
nand U28307 (N_28307,N_27846,N_27986);
nor U28308 (N_28308,N_28044,N_27910);
and U28309 (N_28309,N_27844,N_28039);
nand U28310 (N_28310,N_27744,N_27928);
and U28311 (N_28311,N_28058,N_27801);
xnor U28312 (N_28312,N_27699,N_27964);
nand U28313 (N_28313,N_28109,N_28032);
nand U28314 (N_28314,N_27602,N_28189);
xor U28315 (N_28315,N_27920,N_27675);
nand U28316 (N_28316,N_27944,N_27740);
nor U28317 (N_28317,N_27980,N_28011);
nor U28318 (N_28318,N_27949,N_27898);
and U28319 (N_28319,N_27781,N_27831);
or U28320 (N_28320,N_28078,N_28138);
nor U28321 (N_28321,N_27814,N_27830);
xor U28322 (N_28322,N_27701,N_27770);
nand U28323 (N_28323,N_28046,N_27943);
nor U28324 (N_28324,N_27973,N_27674);
nand U28325 (N_28325,N_28037,N_27710);
and U28326 (N_28326,N_27935,N_28100);
xnor U28327 (N_28327,N_28049,N_27955);
nand U28328 (N_28328,N_28164,N_27806);
and U28329 (N_28329,N_28121,N_28061);
and U28330 (N_28330,N_27773,N_28014);
or U28331 (N_28331,N_27863,N_27631);
nor U28332 (N_28332,N_27921,N_28070);
nor U28333 (N_28333,N_27778,N_28144);
nor U28334 (N_28334,N_27996,N_28127);
or U28335 (N_28335,N_27743,N_27604);
or U28336 (N_28336,N_27782,N_27765);
or U28337 (N_28337,N_27984,N_27908);
nor U28338 (N_28338,N_27856,N_28188);
or U28339 (N_28339,N_28135,N_27919);
nor U28340 (N_28340,N_27677,N_27900);
nand U28341 (N_28341,N_27933,N_28065);
nor U28342 (N_28342,N_27712,N_27862);
or U28343 (N_28343,N_27991,N_27942);
or U28344 (N_28344,N_27633,N_27897);
or U28345 (N_28345,N_27899,N_27686);
or U28346 (N_28346,N_27741,N_28167);
or U28347 (N_28347,N_27972,N_28115);
nor U28348 (N_28348,N_27877,N_27647);
or U28349 (N_28349,N_28177,N_27716);
nand U28350 (N_28350,N_27855,N_27709);
or U28351 (N_28351,N_27967,N_27804);
nand U28352 (N_28352,N_28060,N_27826);
or U28353 (N_28353,N_27946,N_28007);
nand U28354 (N_28354,N_27627,N_28052);
and U28355 (N_28355,N_27727,N_27668);
and U28356 (N_28356,N_27881,N_28080);
xor U28357 (N_28357,N_27894,N_27742);
or U28358 (N_28358,N_27794,N_28084);
and U28359 (N_28359,N_28082,N_27976);
nor U28360 (N_28360,N_27839,N_27706);
nand U28361 (N_28361,N_27671,N_27880);
and U28362 (N_28362,N_28186,N_28193);
and U28363 (N_28363,N_28107,N_27850);
nand U28364 (N_28364,N_27702,N_27718);
or U28365 (N_28365,N_28026,N_27952);
xnor U28366 (N_28366,N_28025,N_28034);
or U28367 (N_28367,N_27823,N_27926);
and U28368 (N_28368,N_28099,N_27879);
xor U28369 (N_28369,N_27669,N_27914);
nand U28370 (N_28370,N_27695,N_27652);
nor U28371 (N_28371,N_27678,N_27998);
and U28372 (N_28372,N_27849,N_27625);
nand U28373 (N_28373,N_27676,N_27800);
or U28374 (N_28374,N_27745,N_27947);
nand U28375 (N_28375,N_28116,N_27609);
nand U28376 (N_28376,N_28170,N_27937);
nand U28377 (N_28377,N_27789,N_27645);
or U28378 (N_28378,N_28016,N_28132);
or U28379 (N_28379,N_28000,N_27751);
nor U28380 (N_28380,N_27837,N_27715);
nand U28381 (N_28381,N_27870,N_28043);
and U28382 (N_28382,N_28033,N_28096);
xor U28383 (N_28383,N_28140,N_28031);
nor U28384 (N_28384,N_27646,N_28150);
or U28385 (N_28385,N_28088,N_28173);
nor U28386 (N_28386,N_28179,N_27906);
or U28387 (N_28387,N_27788,N_28101);
nor U28388 (N_28388,N_28161,N_28128);
nor U28389 (N_28389,N_27845,N_28114);
and U28390 (N_28390,N_27648,N_27963);
nand U28391 (N_28391,N_27815,N_28028);
and U28392 (N_28392,N_27924,N_27666);
or U28393 (N_28393,N_27872,N_27885);
xor U28394 (N_28394,N_27628,N_27606);
or U28395 (N_28395,N_27757,N_28036);
and U28396 (N_28396,N_27915,N_27795);
nor U28397 (N_28397,N_28197,N_27861);
or U28398 (N_28398,N_27685,N_27700);
or U28399 (N_28399,N_27891,N_27637);
or U28400 (N_28400,N_27752,N_28092);
xor U28401 (N_28401,N_27808,N_27763);
nor U28402 (N_28402,N_27687,N_27641);
nand U28403 (N_28403,N_27838,N_27780);
nor U28404 (N_28404,N_27771,N_27760);
and U28405 (N_28405,N_28104,N_27723);
and U28406 (N_28406,N_27655,N_27703);
and U28407 (N_28407,N_27654,N_28008);
and U28408 (N_28408,N_27965,N_27848);
or U28409 (N_28409,N_27774,N_27981);
nand U28410 (N_28410,N_27951,N_27696);
and U28411 (N_28411,N_27731,N_27825);
and U28412 (N_28412,N_27938,N_28009);
or U28413 (N_28413,N_27749,N_27911);
or U28414 (N_28414,N_28184,N_28050);
xnor U28415 (N_28415,N_28051,N_28095);
nor U28416 (N_28416,N_27636,N_27802);
and U28417 (N_28417,N_28053,N_28090);
xnor U28418 (N_28418,N_28019,N_27931);
nand U28419 (N_28419,N_27688,N_27662);
nand U28420 (N_28420,N_28027,N_27912);
nand U28421 (N_28421,N_27634,N_27787);
and U28422 (N_28422,N_27882,N_28108);
and U28423 (N_28423,N_27704,N_28022);
or U28424 (N_28424,N_28063,N_27603);
nand U28425 (N_28425,N_28081,N_28183);
and U28426 (N_28426,N_27777,N_27730);
nand U28427 (N_28427,N_28113,N_27683);
xnor U28428 (N_28428,N_27968,N_28165);
and U28429 (N_28429,N_28117,N_27672);
nand U28430 (N_28430,N_28074,N_27693);
xnor U28431 (N_28431,N_27925,N_27697);
or U28432 (N_28432,N_27684,N_28157);
and U28433 (N_28433,N_27954,N_27624);
xnor U28434 (N_28434,N_28062,N_27974);
and U28435 (N_28435,N_27995,N_28119);
or U28436 (N_28436,N_27890,N_28056);
nor U28437 (N_28437,N_28124,N_27635);
or U28438 (N_28438,N_28158,N_27829);
and U28439 (N_28439,N_27722,N_27738);
or U28440 (N_28440,N_28171,N_27869);
nor U28441 (N_28441,N_27917,N_27783);
and U28442 (N_28442,N_27657,N_27610);
xnor U28443 (N_28443,N_28055,N_27694);
or U28444 (N_28444,N_28045,N_28168);
or U28445 (N_28445,N_28041,N_28146);
nand U28446 (N_28446,N_27813,N_28105);
or U28447 (N_28447,N_28175,N_28166);
and U28448 (N_28448,N_27629,N_27950);
and U28449 (N_28449,N_28040,N_28083);
nand U28450 (N_28450,N_27784,N_27721);
nor U28451 (N_28451,N_27746,N_27735);
nand U28452 (N_28452,N_27734,N_27836);
nor U28453 (N_28453,N_27930,N_28057);
nand U28454 (N_28454,N_28015,N_28097);
nor U28455 (N_28455,N_28118,N_28076);
or U28456 (N_28456,N_27726,N_27725);
nor U28457 (N_28457,N_27859,N_28066);
nor U28458 (N_28458,N_27714,N_27892);
nor U28459 (N_28459,N_28035,N_28106);
nand U28460 (N_28460,N_27623,N_27747);
nor U28461 (N_28461,N_27997,N_28075);
or U28462 (N_28462,N_28130,N_27909);
nand U28463 (N_28463,N_27887,N_27713);
and U28464 (N_28464,N_27620,N_27615);
nor U28465 (N_28465,N_28169,N_27649);
nand U28466 (N_28466,N_27792,N_28153);
nand U28467 (N_28467,N_28093,N_27953);
xor U28468 (N_28468,N_27768,N_27905);
and U28469 (N_28469,N_27960,N_28069);
nor U28470 (N_28470,N_27798,N_27988);
nor U28471 (N_28471,N_28152,N_27970);
nand U28472 (N_28472,N_28199,N_28006);
nor U28473 (N_28473,N_27853,N_27689);
nand U28474 (N_28474,N_27663,N_27618);
nor U28475 (N_28475,N_27983,N_27902);
nor U28476 (N_28476,N_28017,N_27613);
or U28477 (N_28477,N_27824,N_27886);
nand U28478 (N_28478,N_27927,N_27673);
nand U28479 (N_28479,N_28021,N_27797);
or U28480 (N_28480,N_27690,N_28190);
nand U28481 (N_28481,N_27874,N_27656);
or U28482 (N_28482,N_27691,N_28102);
or U28483 (N_28483,N_28151,N_27640);
or U28484 (N_28484,N_28187,N_27803);
and U28485 (N_28485,N_27907,N_28174);
or U28486 (N_28486,N_27865,N_27962);
and U28487 (N_28487,N_27680,N_27679);
nand U28488 (N_28488,N_27737,N_27941);
nand U28489 (N_28489,N_28079,N_28156);
or U28490 (N_28490,N_27889,N_27762);
nand U28491 (N_28491,N_27719,N_27664);
nor U28492 (N_28492,N_27857,N_28087);
or U28493 (N_28493,N_27975,N_28194);
xor U28494 (N_28494,N_27717,N_27939);
nor U28495 (N_28495,N_28129,N_28098);
nor U28496 (N_28496,N_28191,N_28002);
or U28497 (N_28497,N_28010,N_27969);
nor U28498 (N_28498,N_27811,N_27847);
nor U28499 (N_28499,N_27903,N_27600);
nor U28500 (N_28500,N_28173,N_27755);
nor U28501 (N_28501,N_28028,N_27617);
and U28502 (N_28502,N_28090,N_27864);
nand U28503 (N_28503,N_27686,N_27618);
nand U28504 (N_28504,N_28136,N_27639);
and U28505 (N_28505,N_27897,N_28128);
xor U28506 (N_28506,N_27949,N_27720);
nor U28507 (N_28507,N_28003,N_28050);
and U28508 (N_28508,N_27755,N_27994);
and U28509 (N_28509,N_27828,N_27993);
or U28510 (N_28510,N_27745,N_27770);
nand U28511 (N_28511,N_27781,N_27742);
or U28512 (N_28512,N_27811,N_27831);
and U28513 (N_28513,N_27924,N_27778);
or U28514 (N_28514,N_27965,N_27811);
nand U28515 (N_28515,N_27814,N_27837);
nor U28516 (N_28516,N_27801,N_28138);
nand U28517 (N_28517,N_28122,N_27894);
or U28518 (N_28518,N_27701,N_27635);
and U28519 (N_28519,N_27925,N_27904);
nand U28520 (N_28520,N_27813,N_28019);
nand U28521 (N_28521,N_28164,N_28111);
and U28522 (N_28522,N_27733,N_27940);
nor U28523 (N_28523,N_27980,N_27968);
nor U28524 (N_28524,N_27917,N_27801);
nand U28525 (N_28525,N_28182,N_27867);
and U28526 (N_28526,N_27886,N_28075);
nand U28527 (N_28527,N_27649,N_27930);
nand U28528 (N_28528,N_27789,N_27667);
xnor U28529 (N_28529,N_28052,N_27651);
xnor U28530 (N_28530,N_27913,N_28082);
and U28531 (N_28531,N_27905,N_27708);
and U28532 (N_28532,N_27778,N_27827);
nand U28533 (N_28533,N_27827,N_28199);
or U28534 (N_28534,N_27628,N_27855);
or U28535 (N_28535,N_27764,N_28190);
nand U28536 (N_28536,N_27779,N_27688);
nand U28537 (N_28537,N_28198,N_27940);
nand U28538 (N_28538,N_27991,N_27948);
nand U28539 (N_28539,N_27602,N_27848);
xnor U28540 (N_28540,N_27785,N_28199);
and U28541 (N_28541,N_27800,N_28107);
nor U28542 (N_28542,N_28057,N_27964);
nand U28543 (N_28543,N_27722,N_28031);
or U28544 (N_28544,N_27713,N_27881);
nor U28545 (N_28545,N_27937,N_28109);
or U28546 (N_28546,N_27751,N_28059);
and U28547 (N_28547,N_27752,N_27851);
nor U28548 (N_28548,N_28098,N_27900);
and U28549 (N_28549,N_27931,N_27960);
xor U28550 (N_28550,N_27852,N_28100);
or U28551 (N_28551,N_28146,N_27788);
or U28552 (N_28552,N_27711,N_28061);
or U28553 (N_28553,N_28002,N_28186);
or U28554 (N_28554,N_27670,N_27893);
nand U28555 (N_28555,N_28052,N_27614);
and U28556 (N_28556,N_27799,N_28164);
and U28557 (N_28557,N_27923,N_28070);
or U28558 (N_28558,N_27851,N_28119);
xor U28559 (N_28559,N_27945,N_27715);
or U28560 (N_28560,N_28184,N_27616);
or U28561 (N_28561,N_28063,N_27864);
nand U28562 (N_28562,N_27805,N_28062);
or U28563 (N_28563,N_27807,N_28142);
or U28564 (N_28564,N_28136,N_27963);
or U28565 (N_28565,N_27995,N_28017);
and U28566 (N_28566,N_28036,N_27985);
nor U28567 (N_28567,N_28182,N_27787);
xnor U28568 (N_28568,N_27607,N_28150);
nand U28569 (N_28569,N_27849,N_27907);
and U28570 (N_28570,N_27904,N_27706);
xnor U28571 (N_28571,N_27750,N_27912);
or U28572 (N_28572,N_27822,N_28056);
nor U28573 (N_28573,N_28045,N_27820);
nor U28574 (N_28574,N_27985,N_27942);
or U28575 (N_28575,N_27747,N_28174);
nand U28576 (N_28576,N_28158,N_28022);
nand U28577 (N_28577,N_28089,N_27900);
nor U28578 (N_28578,N_27680,N_28012);
nor U28579 (N_28579,N_28159,N_27836);
and U28580 (N_28580,N_28135,N_27687);
xor U28581 (N_28581,N_27672,N_27826);
nor U28582 (N_28582,N_27710,N_27851);
or U28583 (N_28583,N_28180,N_28189);
or U28584 (N_28584,N_28016,N_27639);
nor U28585 (N_28585,N_27968,N_28080);
or U28586 (N_28586,N_27750,N_27958);
nand U28587 (N_28587,N_27894,N_27626);
nor U28588 (N_28588,N_27925,N_27620);
nand U28589 (N_28589,N_27940,N_28003);
nor U28590 (N_28590,N_27610,N_27842);
nand U28591 (N_28591,N_27839,N_28051);
xor U28592 (N_28592,N_28018,N_27930);
or U28593 (N_28593,N_27941,N_28035);
nand U28594 (N_28594,N_28154,N_27825);
nand U28595 (N_28595,N_27627,N_28163);
and U28596 (N_28596,N_28060,N_27764);
nand U28597 (N_28597,N_27830,N_27714);
or U28598 (N_28598,N_27917,N_27843);
nor U28599 (N_28599,N_27769,N_27706);
or U28600 (N_28600,N_27931,N_28048);
nor U28601 (N_28601,N_28000,N_28035);
and U28602 (N_28602,N_27955,N_27839);
nor U28603 (N_28603,N_27734,N_27754);
or U28604 (N_28604,N_27767,N_27741);
nor U28605 (N_28605,N_27928,N_27698);
nand U28606 (N_28606,N_27736,N_27941);
nor U28607 (N_28607,N_27689,N_27980);
xnor U28608 (N_28608,N_28054,N_27834);
or U28609 (N_28609,N_28011,N_28135);
nand U28610 (N_28610,N_28116,N_27987);
and U28611 (N_28611,N_27896,N_27910);
nor U28612 (N_28612,N_28010,N_28072);
nor U28613 (N_28613,N_27625,N_27600);
nand U28614 (N_28614,N_28046,N_27843);
nand U28615 (N_28615,N_28098,N_27868);
xor U28616 (N_28616,N_27625,N_27686);
nor U28617 (N_28617,N_27939,N_28079);
or U28618 (N_28618,N_27802,N_27619);
and U28619 (N_28619,N_28151,N_27975);
nand U28620 (N_28620,N_27773,N_27620);
or U28621 (N_28621,N_27641,N_28063);
nand U28622 (N_28622,N_27961,N_28011);
or U28623 (N_28623,N_27712,N_27878);
and U28624 (N_28624,N_27966,N_28155);
nor U28625 (N_28625,N_27751,N_27894);
and U28626 (N_28626,N_27714,N_27998);
or U28627 (N_28627,N_27737,N_28199);
and U28628 (N_28628,N_27809,N_28157);
nand U28629 (N_28629,N_28130,N_27614);
nor U28630 (N_28630,N_27703,N_28162);
nor U28631 (N_28631,N_28158,N_28190);
nand U28632 (N_28632,N_27960,N_27808);
and U28633 (N_28633,N_27985,N_27655);
nor U28634 (N_28634,N_27657,N_27769);
nand U28635 (N_28635,N_27810,N_27989);
xor U28636 (N_28636,N_28093,N_27617);
xor U28637 (N_28637,N_28017,N_27763);
or U28638 (N_28638,N_28184,N_28185);
xnor U28639 (N_28639,N_27782,N_28132);
and U28640 (N_28640,N_28024,N_28137);
nor U28641 (N_28641,N_28175,N_28189);
nand U28642 (N_28642,N_28130,N_27952);
or U28643 (N_28643,N_27963,N_27830);
nor U28644 (N_28644,N_27660,N_28167);
nor U28645 (N_28645,N_28056,N_28050);
nand U28646 (N_28646,N_28145,N_27945);
or U28647 (N_28647,N_28014,N_27808);
nor U28648 (N_28648,N_28054,N_28030);
nor U28649 (N_28649,N_27661,N_27971);
or U28650 (N_28650,N_28035,N_28100);
and U28651 (N_28651,N_27682,N_27614);
or U28652 (N_28652,N_28007,N_27688);
and U28653 (N_28653,N_27731,N_28014);
nand U28654 (N_28654,N_27865,N_28193);
nor U28655 (N_28655,N_28158,N_28106);
and U28656 (N_28656,N_28089,N_28102);
nand U28657 (N_28657,N_27718,N_27785);
or U28658 (N_28658,N_27633,N_28010);
nand U28659 (N_28659,N_27750,N_27811);
xor U28660 (N_28660,N_27783,N_27616);
or U28661 (N_28661,N_27617,N_27977);
or U28662 (N_28662,N_27874,N_27702);
nand U28663 (N_28663,N_27736,N_27689);
or U28664 (N_28664,N_28014,N_27932);
and U28665 (N_28665,N_28192,N_27936);
and U28666 (N_28666,N_28014,N_28109);
nand U28667 (N_28667,N_28091,N_27764);
or U28668 (N_28668,N_28023,N_27887);
nand U28669 (N_28669,N_28195,N_28160);
or U28670 (N_28670,N_28071,N_28148);
xor U28671 (N_28671,N_27936,N_27801);
and U28672 (N_28672,N_27877,N_28121);
xnor U28673 (N_28673,N_28088,N_28106);
xor U28674 (N_28674,N_27859,N_27871);
or U28675 (N_28675,N_27979,N_27850);
or U28676 (N_28676,N_28042,N_28092);
nand U28677 (N_28677,N_27806,N_27852);
nor U28678 (N_28678,N_27991,N_28118);
nor U28679 (N_28679,N_28181,N_27746);
nor U28680 (N_28680,N_28020,N_27755);
nor U28681 (N_28681,N_27925,N_28153);
nor U28682 (N_28682,N_27744,N_27695);
xor U28683 (N_28683,N_28173,N_27996);
or U28684 (N_28684,N_27841,N_27747);
nand U28685 (N_28685,N_27670,N_28022);
nor U28686 (N_28686,N_28157,N_27708);
nand U28687 (N_28687,N_27879,N_27867);
or U28688 (N_28688,N_27809,N_27905);
nand U28689 (N_28689,N_28197,N_27847);
nand U28690 (N_28690,N_28014,N_28026);
nand U28691 (N_28691,N_28106,N_28022);
nand U28692 (N_28692,N_28035,N_27715);
nand U28693 (N_28693,N_28039,N_27721);
nand U28694 (N_28694,N_27864,N_27909);
or U28695 (N_28695,N_27922,N_27716);
and U28696 (N_28696,N_27683,N_27842);
xnor U28697 (N_28697,N_28001,N_28026);
or U28698 (N_28698,N_28178,N_28164);
nor U28699 (N_28699,N_28000,N_27852);
nand U28700 (N_28700,N_28144,N_28071);
or U28701 (N_28701,N_27928,N_28189);
nand U28702 (N_28702,N_28036,N_27879);
and U28703 (N_28703,N_27982,N_27976);
xor U28704 (N_28704,N_28103,N_28030);
and U28705 (N_28705,N_27854,N_28170);
nor U28706 (N_28706,N_27688,N_28145);
or U28707 (N_28707,N_27869,N_27883);
nor U28708 (N_28708,N_27802,N_28161);
and U28709 (N_28709,N_28128,N_28028);
nor U28710 (N_28710,N_27698,N_28048);
and U28711 (N_28711,N_27623,N_27679);
xnor U28712 (N_28712,N_27819,N_27990);
nor U28713 (N_28713,N_27898,N_27803);
or U28714 (N_28714,N_28178,N_27737);
nand U28715 (N_28715,N_27728,N_27833);
xnor U28716 (N_28716,N_28096,N_27893);
xnor U28717 (N_28717,N_28143,N_27762);
nand U28718 (N_28718,N_28198,N_28050);
xor U28719 (N_28719,N_27974,N_27649);
nand U28720 (N_28720,N_27641,N_28138);
xnor U28721 (N_28721,N_27811,N_28067);
nor U28722 (N_28722,N_28086,N_27845);
and U28723 (N_28723,N_27911,N_28097);
nand U28724 (N_28724,N_27686,N_27959);
xnor U28725 (N_28725,N_27704,N_27837);
nand U28726 (N_28726,N_27615,N_27643);
nor U28727 (N_28727,N_27612,N_27810);
nand U28728 (N_28728,N_27880,N_28148);
nand U28729 (N_28729,N_27920,N_27971);
xnor U28730 (N_28730,N_28137,N_27859);
nor U28731 (N_28731,N_27705,N_27605);
nand U28732 (N_28732,N_27703,N_27867);
and U28733 (N_28733,N_27888,N_27818);
or U28734 (N_28734,N_27602,N_28194);
xnor U28735 (N_28735,N_28149,N_27993);
nand U28736 (N_28736,N_27941,N_27909);
and U28737 (N_28737,N_27743,N_28076);
or U28738 (N_28738,N_27749,N_27608);
nor U28739 (N_28739,N_27722,N_27608);
or U28740 (N_28740,N_27827,N_27759);
or U28741 (N_28741,N_27809,N_28088);
and U28742 (N_28742,N_28190,N_27715);
nor U28743 (N_28743,N_28073,N_28106);
and U28744 (N_28744,N_27653,N_27997);
nor U28745 (N_28745,N_28010,N_28070);
xnor U28746 (N_28746,N_27732,N_27838);
xnor U28747 (N_28747,N_28181,N_28089);
and U28748 (N_28748,N_27950,N_27722);
xnor U28749 (N_28749,N_27953,N_28138);
or U28750 (N_28750,N_27706,N_27966);
or U28751 (N_28751,N_27875,N_27659);
nor U28752 (N_28752,N_27933,N_27856);
and U28753 (N_28753,N_28197,N_27829);
and U28754 (N_28754,N_27952,N_28182);
nand U28755 (N_28755,N_27682,N_28008);
or U28756 (N_28756,N_27671,N_27851);
or U28757 (N_28757,N_27752,N_28056);
nand U28758 (N_28758,N_27961,N_28179);
or U28759 (N_28759,N_27943,N_27795);
xor U28760 (N_28760,N_28144,N_28054);
nand U28761 (N_28761,N_27642,N_27856);
and U28762 (N_28762,N_27986,N_28022);
nor U28763 (N_28763,N_27737,N_27949);
nor U28764 (N_28764,N_27631,N_28166);
nor U28765 (N_28765,N_27754,N_28115);
nor U28766 (N_28766,N_27965,N_28078);
nand U28767 (N_28767,N_27881,N_27611);
nand U28768 (N_28768,N_28032,N_27908);
nor U28769 (N_28769,N_27884,N_27804);
nor U28770 (N_28770,N_27709,N_28128);
nand U28771 (N_28771,N_28042,N_27951);
or U28772 (N_28772,N_27932,N_27761);
nor U28773 (N_28773,N_27608,N_27669);
and U28774 (N_28774,N_27974,N_27627);
or U28775 (N_28775,N_27640,N_28083);
nor U28776 (N_28776,N_28022,N_27616);
nor U28777 (N_28777,N_27866,N_28006);
nor U28778 (N_28778,N_27944,N_28019);
or U28779 (N_28779,N_27853,N_28106);
nor U28780 (N_28780,N_27901,N_28099);
nor U28781 (N_28781,N_27936,N_27748);
or U28782 (N_28782,N_28046,N_27694);
nand U28783 (N_28783,N_27616,N_28009);
nor U28784 (N_28784,N_27780,N_28098);
or U28785 (N_28785,N_27812,N_27628);
nand U28786 (N_28786,N_27796,N_28047);
and U28787 (N_28787,N_27637,N_27929);
nor U28788 (N_28788,N_28015,N_27625);
nand U28789 (N_28789,N_27932,N_28017);
nand U28790 (N_28790,N_27919,N_27979);
nor U28791 (N_28791,N_27927,N_28071);
and U28792 (N_28792,N_27996,N_27877);
nand U28793 (N_28793,N_27655,N_27749);
or U28794 (N_28794,N_27928,N_28128);
or U28795 (N_28795,N_27937,N_27916);
and U28796 (N_28796,N_27751,N_27613);
xnor U28797 (N_28797,N_27797,N_27969);
and U28798 (N_28798,N_27684,N_27961);
nor U28799 (N_28799,N_27893,N_27797);
and U28800 (N_28800,N_28470,N_28236);
and U28801 (N_28801,N_28451,N_28742);
xnor U28802 (N_28802,N_28260,N_28755);
nor U28803 (N_28803,N_28442,N_28384);
nor U28804 (N_28804,N_28393,N_28323);
xnor U28805 (N_28805,N_28539,N_28310);
nand U28806 (N_28806,N_28762,N_28220);
nand U28807 (N_28807,N_28397,N_28471);
and U28808 (N_28808,N_28559,N_28738);
nand U28809 (N_28809,N_28459,N_28322);
and U28810 (N_28810,N_28777,N_28340);
nand U28811 (N_28811,N_28207,N_28720);
and U28812 (N_28812,N_28757,N_28282);
or U28813 (N_28813,N_28558,N_28360);
and U28814 (N_28814,N_28683,N_28756);
nand U28815 (N_28815,N_28784,N_28237);
and U28816 (N_28816,N_28351,N_28350);
nand U28817 (N_28817,N_28484,N_28329);
or U28818 (N_28818,N_28311,N_28209);
nand U28819 (N_28819,N_28366,N_28268);
nor U28820 (N_28820,N_28303,N_28345);
and U28821 (N_28821,N_28555,N_28272);
and U28822 (N_28822,N_28604,N_28599);
nand U28823 (N_28823,N_28563,N_28717);
nand U28824 (N_28824,N_28705,N_28513);
nand U28825 (N_28825,N_28331,N_28505);
xnor U28826 (N_28826,N_28244,N_28709);
and U28827 (N_28827,N_28456,N_28792);
nand U28828 (N_28828,N_28464,N_28702);
nor U28829 (N_28829,N_28579,N_28488);
nand U28830 (N_28830,N_28342,N_28431);
nand U28831 (N_28831,N_28284,N_28361);
or U28832 (N_28832,N_28706,N_28715);
nand U28833 (N_28833,N_28576,N_28733);
and U28834 (N_28834,N_28443,N_28673);
or U28835 (N_28835,N_28634,N_28222);
and U28836 (N_28836,N_28628,N_28518);
nand U28837 (N_28837,N_28496,N_28290);
or U28838 (N_28838,N_28694,N_28573);
nand U28839 (N_28839,N_28250,N_28646);
or U28840 (N_28840,N_28652,N_28789);
and U28841 (N_28841,N_28580,N_28206);
and U28842 (N_28842,N_28453,N_28753);
nand U28843 (N_28843,N_28502,N_28438);
or U28844 (N_28844,N_28759,N_28328);
nor U28845 (N_28845,N_28776,N_28463);
xor U28846 (N_28846,N_28631,N_28658);
nand U28847 (N_28847,N_28202,N_28257);
and U28848 (N_28848,N_28386,N_28280);
nor U28849 (N_28849,N_28743,N_28647);
nor U28850 (N_28850,N_28781,N_28273);
nor U28851 (N_28851,N_28740,N_28294);
nand U28852 (N_28852,N_28668,N_28359);
or U28853 (N_28853,N_28779,N_28653);
nor U28854 (N_28854,N_28548,N_28487);
or U28855 (N_28855,N_28622,N_28427);
or U28856 (N_28856,N_28748,N_28216);
nand U28857 (N_28857,N_28317,N_28557);
nor U28858 (N_28858,N_28379,N_28609);
and U28859 (N_28859,N_28274,N_28400);
and U28860 (N_28860,N_28746,N_28674);
or U28861 (N_28861,N_28507,N_28293);
and U28862 (N_28862,N_28452,N_28461);
nor U28863 (N_28863,N_28474,N_28449);
and U28864 (N_28864,N_28356,N_28565);
or U28865 (N_28865,N_28349,N_28473);
nand U28866 (N_28866,N_28265,N_28786);
nor U28867 (N_28867,N_28335,N_28574);
nand U28868 (N_28868,N_28594,N_28312);
or U28869 (N_28869,N_28319,N_28736);
or U28870 (N_28870,N_28527,N_28681);
and U28871 (N_28871,N_28561,N_28691);
nor U28872 (N_28872,N_28578,N_28223);
nand U28873 (N_28873,N_28430,N_28554);
or U28874 (N_28874,N_28306,N_28568);
or U28875 (N_28875,N_28258,N_28371);
or U28876 (N_28876,N_28607,N_28656);
nor U28877 (N_28877,N_28208,N_28435);
nor U28878 (N_28878,N_28642,N_28663);
nor U28879 (N_28879,N_28670,N_28472);
nor U28880 (N_28880,N_28572,N_28590);
and U28881 (N_28881,N_28367,N_28398);
and U28882 (N_28882,N_28466,N_28725);
nand U28883 (N_28883,N_28585,N_28546);
or U28884 (N_28884,N_28662,N_28440);
and U28885 (N_28885,N_28562,N_28245);
and U28886 (N_28886,N_28637,N_28300);
and U28887 (N_28887,N_28531,N_28751);
nand U28888 (N_28888,N_28327,N_28549);
or U28889 (N_28889,N_28448,N_28763);
nor U28890 (N_28890,N_28541,N_28227);
xnor U28891 (N_28891,N_28688,N_28426);
and U28892 (N_28892,N_28538,N_28299);
or U28893 (N_28893,N_28354,N_28231);
or U28894 (N_28894,N_28352,N_28401);
and U28895 (N_28895,N_28727,N_28644);
or U28896 (N_28896,N_28510,N_28616);
and U28897 (N_28897,N_28512,N_28372);
or U28898 (N_28898,N_28424,N_28376);
nor U28899 (N_28899,N_28246,N_28506);
nand U28900 (N_28900,N_28754,N_28785);
nor U28901 (N_28901,N_28788,N_28229);
nand U28902 (N_28902,N_28730,N_28326);
nor U28903 (N_28903,N_28529,N_28385);
and U28904 (N_28904,N_28591,N_28457);
nor U28905 (N_28905,N_28680,N_28693);
nand U28906 (N_28906,N_28315,N_28467);
nor U28907 (N_28907,N_28783,N_28666);
nand U28908 (N_28908,N_28621,N_28712);
and U28909 (N_28909,N_28469,N_28758);
nor U28910 (N_28910,N_28492,N_28497);
or U28911 (N_28911,N_28339,N_28597);
nand U28912 (N_28912,N_28677,N_28445);
nor U28913 (N_28913,N_28545,N_28460);
or U28914 (N_28914,N_28728,N_28570);
or U28915 (N_28915,N_28796,N_28262);
nand U28916 (N_28916,N_28575,N_28532);
xnor U28917 (N_28917,N_28791,N_28455);
xor U28918 (N_28918,N_28544,N_28203);
nor U28919 (N_28919,N_28217,N_28234);
nor U28920 (N_28920,N_28588,N_28287);
nand U28921 (N_28921,N_28719,N_28291);
nand U28922 (N_28922,N_28407,N_28414);
nand U28923 (N_28923,N_28745,N_28774);
xor U28924 (N_28924,N_28700,N_28556);
xor U28925 (N_28925,N_28675,N_28655);
or U28926 (N_28926,N_28627,N_28269);
nor U28927 (N_28927,N_28213,N_28498);
and U28928 (N_28928,N_28416,N_28739);
nand U28929 (N_28929,N_28794,N_28678);
nor U28930 (N_28930,N_28228,N_28550);
nor U28931 (N_28931,N_28483,N_28699);
and U28932 (N_28932,N_28687,N_28271);
and U28933 (N_28933,N_28664,N_28423);
and U28934 (N_28934,N_28566,N_28251);
and U28935 (N_28935,N_28295,N_28343);
or U28936 (N_28936,N_28241,N_28434);
or U28937 (N_28937,N_28406,N_28204);
nand U28938 (N_28938,N_28704,N_28582);
and U28939 (N_28939,N_28744,N_28635);
nor U28940 (N_28940,N_28615,N_28242);
xor U28941 (N_28941,N_28767,N_28648);
nand U28942 (N_28942,N_28761,N_28309);
nand U28943 (N_28943,N_28316,N_28729);
nor U28944 (N_28944,N_28528,N_28569);
nor U28945 (N_28945,N_28617,N_28252);
nor U28946 (N_28946,N_28358,N_28612);
nand U28947 (N_28947,N_28645,N_28436);
xnor U28948 (N_28948,N_28410,N_28296);
nand U28949 (N_28949,N_28638,N_28418);
xnor U28950 (N_28950,N_28253,N_28347);
xor U28951 (N_28951,N_28679,N_28598);
and U28952 (N_28952,N_28396,N_28490);
nor U28953 (N_28953,N_28649,N_28651);
or U28954 (N_28954,N_28314,N_28288);
nand U28955 (N_28955,N_28551,N_28522);
nor U28956 (N_28956,N_28703,N_28479);
or U28957 (N_28957,N_28749,N_28696);
and U28958 (N_28958,N_28485,N_28281);
and U28959 (N_28959,N_28261,N_28224);
and U28960 (N_28960,N_28491,N_28540);
and U28961 (N_28961,N_28239,N_28526);
nand U28962 (N_28962,N_28307,N_28337);
nand U28963 (N_28963,N_28797,N_28403);
xor U28964 (N_28964,N_28798,N_28643);
xnor U28965 (N_28965,N_28332,N_28458);
or U28966 (N_28966,N_28760,N_28308);
nor U28967 (N_28967,N_28238,N_28489);
nor U28968 (N_28968,N_28773,N_28698);
xnor U28969 (N_28969,N_28793,N_28364);
nand U28970 (N_28970,N_28665,N_28405);
or U28971 (N_28971,N_28475,N_28221);
nand U28972 (N_28972,N_28593,N_28369);
nor U28973 (N_28973,N_28641,N_28583);
nor U28974 (N_28974,N_28377,N_28375);
nor U28975 (N_28975,N_28277,N_28750);
and U28976 (N_28976,N_28571,N_28338);
xor U28977 (N_28977,N_28346,N_28721);
nor U28978 (N_28978,N_28500,N_28795);
nand U28979 (N_28979,N_28420,N_28447);
nand U28980 (N_28980,N_28370,N_28596);
nand U28981 (N_28981,N_28333,N_28595);
nand U28982 (N_28982,N_28639,N_28263);
and U28983 (N_28983,N_28486,N_28632);
nand U28984 (N_28984,N_28536,N_28508);
or U28985 (N_28985,N_28205,N_28765);
or U28986 (N_28986,N_28465,N_28324);
nand U28987 (N_28987,N_28256,N_28504);
nor U28988 (N_28988,N_28605,N_28499);
or U28989 (N_28989,N_28399,N_28610);
or U28990 (N_28990,N_28355,N_28654);
or U28991 (N_28991,N_28279,N_28477);
nor U28992 (N_28992,N_28247,N_28378);
xnor U28993 (N_28993,N_28584,N_28537);
nor U28994 (N_28994,N_28368,N_28259);
xnor U28995 (N_28995,N_28592,N_28685);
nor U28996 (N_28996,N_28425,N_28577);
and U28997 (N_28997,N_28480,N_28707);
or U28998 (N_28998,N_28439,N_28524);
and U28999 (N_28999,N_28567,N_28283);
nor U29000 (N_29000,N_28735,N_28650);
and U29001 (N_29001,N_28408,N_28402);
nor U29002 (N_29002,N_28667,N_28468);
and U29003 (N_29003,N_28240,N_28640);
nand U29004 (N_29004,N_28363,N_28737);
and U29005 (N_29005,N_28422,N_28444);
nand U29006 (N_29006,N_28606,N_28623);
xor U29007 (N_29007,N_28432,N_28501);
nor U29008 (N_29008,N_28629,N_28482);
nor U29009 (N_29009,N_28603,N_28718);
nand U29010 (N_29010,N_28600,N_28374);
nor U29011 (N_29011,N_28441,N_28362);
and U29012 (N_29012,N_28478,N_28417);
or U29013 (N_29013,N_28782,N_28611);
and U29014 (N_29014,N_28454,N_28692);
and U29015 (N_29015,N_28373,N_28768);
nand U29016 (N_29016,N_28318,N_28225);
or U29017 (N_29017,N_28334,N_28534);
xnor U29018 (N_29018,N_28357,N_28676);
or U29019 (N_29019,N_28428,N_28313);
and U29020 (N_29020,N_28613,N_28301);
nand U29021 (N_29021,N_28476,N_28521);
nand U29022 (N_29022,N_28320,N_28519);
nand U29023 (N_29023,N_28330,N_28686);
and U29024 (N_29024,N_28302,N_28726);
nand U29025 (N_29025,N_28429,N_28626);
and U29026 (N_29026,N_28353,N_28219);
xnor U29027 (N_29027,N_28503,N_28747);
and U29028 (N_29028,N_28233,N_28278);
or U29029 (N_29029,N_28415,N_28602);
and U29030 (N_29030,N_28619,N_28481);
and U29031 (N_29031,N_28248,N_28341);
xor U29032 (N_29032,N_28230,N_28382);
and U29033 (N_29033,N_28215,N_28243);
nor U29034 (N_29034,N_28708,N_28542);
xnor U29035 (N_29035,N_28581,N_28625);
and U29036 (N_29036,N_28714,N_28421);
nor U29037 (N_29037,N_28553,N_28620);
and U29038 (N_29038,N_28732,N_28286);
nand U29039 (N_29039,N_28778,N_28601);
nor U29040 (N_29040,N_28344,N_28409);
nor U29041 (N_29041,N_28517,N_28766);
nor U29042 (N_29042,N_28270,N_28516);
xor U29043 (N_29043,N_28495,N_28711);
xnor U29044 (N_29044,N_28547,N_28433);
nand U29045 (N_29045,N_28226,N_28520);
nor U29046 (N_29046,N_28701,N_28235);
nand U29047 (N_29047,N_28201,N_28672);
and U29048 (N_29048,N_28212,N_28365);
nand U29049 (N_29049,N_28775,N_28723);
nor U29050 (N_29050,N_28394,N_28321);
or U29051 (N_29051,N_28325,N_28552);
and U29052 (N_29052,N_28589,N_28276);
and U29053 (N_29053,N_28525,N_28450);
and U29054 (N_29054,N_28210,N_28614);
nand U29055 (N_29055,N_28211,N_28669);
xor U29056 (N_29056,N_28390,N_28298);
nand U29057 (N_29057,N_28413,N_28660);
and U29058 (N_29058,N_28722,N_28404);
and U29059 (N_29059,N_28690,N_28264);
nor U29060 (N_29060,N_28587,N_28695);
nor U29061 (N_29061,N_28618,N_28304);
nor U29062 (N_29062,N_28523,N_28636);
or U29063 (N_29063,N_28764,N_28336);
or U29064 (N_29064,N_28218,N_28586);
nor U29065 (N_29065,N_28535,N_28249);
or U29066 (N_29066,N_28391,N_28383);
nor U29067 (N_29067,N_28543,N_28514);
or U29068 (N_29068,N_28724,N_28689);
or U29069 (N_29069,N_28790,N_28289);
xor U29070 (N_29070,N_28297,N_28285);
nor U29071 (N_29071,N_28266,N_28395);
nor U29072 (N_29072,N_28419,N_28381);
nor U29073 (N_29073,N_28799,N_28741);
or U29074 (N_29074,N_28697,N_28769);
and U29075 (N_29075,N_28684,N_28254);
nand U29076 (N_29076,N_28624,N_28255);
nand U29077 (N_29077,N_28446,N_28437);
and U29078 (N_29078,N_28380,N_28682);
and U29079 (N_29079,N_28633,N_28780);
and U29080 (N_29080,N_28494,N_28659);
and U29081 (N_29081,N_28530,N_28232);
and U29082 (N_29082,N_28509,N_28713);
nor U29083 (N_29083,N_28710,N_28389);
and U29084 (N_29084,N_28392,N_28787);
or U29085 (N_29085,N_28771,N_28772);
and U29086 (N_29086,N_28731,N_28630);
or U29087 (N_29087,N_28275,N_28752);
nand U29088 (N_29088,N_28462,N_28661);
and U29089 (N_29089,N_28770,N_28533);
xor U29090 (N_29090,N_28671,N_28511);
and U29091 (N_29091,N_28734,N_28292);
xor U29092 (N_29092,N_28608,N_28305);
xor U29093 (N_29093,N_28560,N_28267);
nand U29094 (N_29094,N_28412,N_28493);
nand U29095 (N_29095,N_28564,N_28716);
or U29096 (N_29096,N_28657,N_28388);
or U29097 (N_29097,N_28200,N_28515);
and U29098 (N_29098,N_28214,N_28411);
or U29099 (N_29099,N_28348,N_28387);
nand U29100 (N_29100,N_28769,N_28235);
or U29101 (N_29101,N_28268,N_28266);
nor U29102 (N_29102,N_28679,N_28252);
nand U29103 (N_29103,N_28230,N_28754);
nor U29104 (N_29104,N_28570,N_28417);
or U29105 (N_29105,N_28735,N_28787);
nand U29106 (N_29106,N_28351,N_28387);
or U29107 (N_29107,N_28599,N_28287);
or U29108 (N_29108,N_28763,N_28666);
xnor U29109 (N_29109,N_28550,N_28296);
nor U29110 (N_29110,N_28541,N_28591);
nor U29111 (N_29111,N_28559,N_28375);
nor U29112 (N_29112,N_28733,N_28648);
nor U29113 (N_29113,N_28737,N_28663);
nand U29114 (N_29114,N_28591,N_28350);
and U29115 (N_29115,N_28551,N_28381);
nor U29116 (N_29116,N_28330,N_28660);
and U29117 (N_29117,N_28522,N_28345);
xnor U29118 (N_29118,N_28781,N_28507);
or U29119 (N_29119,N_28270,N_28665);
nand U29120 (N_29120,N_28434,N_28683);
or U29121 (N_29121,N_28653,N_28737);
nor U29122 (N_29122,N_28737,N_28398);
xnor U29123 (N_29123,N_28431,N_28623);
nand U29124 (N_29124,N_28607,N_28340);
and U29125 (N_29125,N_28305,N_28738);
nand U29126 (N_29126,N_28526,N_28505);
xor U29127 (N_29127,N_28438,N_28213);
nor U29128 (N_29128,N_28376,N_28768);
nand U29129 (N_29129,N_28626,N_28607);
nand U29130 (N_29130,N_28290,N_28470);
and U29131 (N_29131,N_28338,N_28415);
nor U29132 (N_29132,N_28210,N_28535);
nor U29133 (N_29133,N_28416,N_28394);
nor U29134 (N_29134,N_28314,N_28589);
and U29135 (N_29135,N_28479,N_28528);
nand U29136 (N_29136,N_28746,N_28560);
nand U29137 (N_29137,N_28461,N_28605);
nand U29138 (N_29138,N_28791,N_28504);
or U29139 (N_29139,N_28632,N_28470);
nor U29140 (N_29140,N_28780,N_28731);
nand U29141 (N_29141,N_28353,N_28448);
or U29142 (N_29142,N_28237,N_28671);
nand U29143 (N_29143,N_28432,N_28576);
and U29144 (N_29144,N_28330,N_28264);
and U29145 (N_29145,N_28524,N_28217);
nor U29146 (N_29146,N_28359,N_28767);
and U29147 (N_29147,N_28793,N_28558);
nand U29148 (N_29148,N_28420,N_28557);
nand U29149 (N_29149,N_28478,N_28659);
nor U29150 (N_29150,N_28345,N_28439);
and U29151 (N_29151,N_28308,N_28244);
or U29152 (N_29152,N_28726,N_28578);
nand U29153 (N_29153,N_28309,N_28356);
nor U29154 (N_29154,N_28536,N_28430);
or U29155 (N_29155,N_28340,N_28311);
and U29156 (N_29156,N_28606,N_28586);
nand U29157 (N_29157,N_28223,N_28262);
xnor U29158 (N_29158,N_28752,N_28592);
xor U29159 (N_29159,N_28649,N_28410);
and U29160 (N_29160,N_28488,N_28291);
and U29161 (N_29161,N_28431,N_28415);
and U29162 (N_29162,N_28248,N_28790);
xnor U29163 (N_29163,N_28738,N_28323);
nor U29164 (N_29164,N_28795,N_28685);
xor U29165 (N_29165,N_28622,N_28335);
and U29166 (N_29166,N_28703,N_28307);
nor U29167 (N_29167,N_28607,N_28260);
xnor U29168 (N_29168,N_28599,N_28365);
and U29169 (N_29169,N_28210,N_28691);
nor U29170 (N_29170,N_28651,N_28484);
nand U29171 (N_29171,N_28231,N_28572);
or U29172 (N_29172,N_28554,N_28272);
nand U29173 (N_29173,N_28410,N_28451);
xor U29174 (N_29174,N_28383,N_28609);
xor U29175 (N_29175,N_28720,N_28705);
and U29176 (N_29176,N_28255,N_28769);
xnor U29177 (N_29177,N_28438,N_28733);
nor U29178 (N_29178,N_28711,N_28498);
nor U29179 (N_29179,N_28347,N_28288);
or U29180 (N_29180,N_28624,N_28300);
nor U29181 (N_29181,N_28229,N_28356);
nand U29182 (N_29182,N_28514,N_28720);
or U29183 (N_29183,N_28733,N_28342);
nand U29184 (N_29184,N_28435,N_28582);
nor U29185 (N_29185,N_28454,N_28395);
nand U29186 (N_29186,N_28230,N_28460);
and U29187 (N_29187,N_28714,N_28445);
and U29188 (N_29188,N_28779,N_28335);
xnor U29189 (N_29189,N_28696,N_28725);
or U29190 (N_29190,N_28261,N_28642);
xnor U29191 (N_29191,N_28719,N_28473);
or U29192 (N_29192,N_28317,N_28605);
nor U29193 (N_29193,N_28384,N_28763);
nand U29194 (N_29194,N_28479,N_28359);
nor U29195 (N_29195,N_28343,N_28424);
or U29196 (N_29196,N_28630,N_28463);
and U29197 (N_29197,N_28707,N_28599);
or U29198 (N_29198,N_28387,N_28703);
nand U29199 (N_29199,N_28523,N_28420);
nor U29200 (N_29200,N_28716,N_28533);
and U29201 (N_29201,N_28585,N_28715);
nor U29202 (N_29202,N_28674,N_28528);
nor U29203 (N_29203,N_28709,N_28504);
or U29204 (N_29204,N_28449,N_28488);
nand U29205 (N_29205,N_28613,N_28566);
or U29206 (N_29206,N_28328,N_28783);
nor U29207 (N_29207,N_28238,N_28499);
or U29208 (N_29208,N_28690,N_28331);
or U29209 (N_29209,N_28311,N_28392);
nand U29210 (N_29210,N_28328,N_28435);
nor U29211 (N_29211,N_28597,N_28732);
xor U29212 (N_29212,N_28567,N_28699);
nand U29213 (N_29213,N_28709,N_28673);
nand U29214 (N_29214,N_28792,N_28711);
or U29215 (N_29215,N_28661,N_28490);
xnor U29216 (N_29216,N_28776,N_28561);
xor U29217 (N_29217,N_28205,N_28696);
nor U29218 (N_29218,N_28696,N_28259);
nor U29219 (N_29219,N_28275,N_28715);
or U29220 (N_29220,N_28277,N_28673);
nor U29221 (N_29221,N_28471,N_28648);
nor U29222 (N_29222,N_28342,N_28750);
and U29223 (N_29223,N_28634,N_28219);
xnor U29224 (N_29224,N_28791,N_28594);
nor U29225 (N_29225,N_28379,N_28217);
or U29226 (N_29226,N_28428,N_28664);
and U29227 (N_29227,N_28773,N_28472);
and U29228 (N_29228,N_28776,N_28283);
and U29229 (N_29229,N_28714,N_28768);
and U29230 (N_29230,N_28735,N_28335);
or U29231 (N_29231,N_28667,N_28478);
nor U29232 (N_29232,N_28767,N_28565);
nand U29233 (N_29233,N_28524,N_28756);
or U29234 (N_29234,N_28774,N_28759);
nand U29235 (N_29235,N_28577,N_28513);
nor U29236 (N_29236,N_28471,N_28543);
and U29237 (N_29237,N_28586,N_28719);
nor U29238 (N_29238,N_28754,N_28409);
xor U29239 (N_29239,N_28339,N_28502);
nor U29240 (N_29240,N_28252,N_28785);
xnor U29241 (N_29241,N_28236,N_28544);
or U29242 (N_29242,N_28450,N_28508);
and U29243 (N_29243,N_28661,N_28312);
and U29244 (N_29244,N_28609,N_28796);
nand U29245 (N_29245,N_28548,N_28794);
and U29246 (N_29246,N_28296,N_28623);
nor U29247 (N_29247,N_28394,N_28441);
and U29248 (N_29248,N_28500,N_28710);
xnor U29249 (N_29249,N_28500,N_28456);
nand U29250 (N_29250,N_28528,N_28669);
and U29251 (N_29251,N_28503,N_28358);
nand U29252 (N_29252,N_28535,N_28483);
nand U29253 (N_29253,N_28632,N_28527);
nand U29254 (N_29254,N_28737,N_28510);
nor U29255 (N_29255,N_28251,N_28727);
or U29256 (N_29256,N_28442,N_28623);
or U29257 (N_29257,N_28622,N_28316);
and U29258 (N_29258,N_28516,N_28777);
and U29259 (N_29259,N_28502,N_28413);
nand U29260 (N_29260,N_28338,N_28645);
or U29261 (N_29261,N_28281,N_28608);
nand U29262 (N_29262,N_28461,N_28719);
nor U29263 (N_29263,N_28774,N_28230);
and U29264 (N_29264,N_28345,N_28274);
and U29265 (N_29265,N_28582,N_28791);
nand U29266 (N_29266,N_28726,N_28214);
xnor U29267 (N_29267,N_28694,N_28564);
nand U29268 (N_29268,N_28291,N_28345);
and U29269 (N_29269,N_28438,N_28285);
and U29270 (N_29270,N_28475,N_28249);
and U29271 (N_29271,N_28237,N_28662);
nor U29272 (N_29272,N_28305,N_28240);
nor U29273 (N_29273,N_28375,N_28313);
nor U29274 (N_29274,N_28606,N_28356);
and U29275 (N_29275,N_28658,N_28551);
nor U29276 (N_29276,N_28224,N_28244);
nand U29277 (N_29277,N_28786,N_28325);
or U29278 (N_29278,N_28765,N_28733);
or U29279 (N_29279,N_28578,N_28688);
nor U29280 (N_29280,N_28480,N_28226);
nor U29281 (N_29281,N_28754,N_28318);
and U29282 (N_29282,N_28296,N_28462);
xnor U29283 (N_29283,N_28369,N_28762);
nand U29284 (N_29284,N_28600,N_28539);
nand U29285 (N_29285,N_28282,N_28291);
or U29286 (N_29286,N_28363,N_28486);
nand U29287 (N_29287,N_28424,N_28657);
nor U29288 (N_29288,N_28599,N_28222);
nand U29289 (N_29289,N_28398,N_28218);
nand U29290 (N_29290,N_28212,N_28575);
nand U29291 (N_29291,N_28472,N_28561);
nor U29292 (N_29292,N_28423,N_28795);
or U29293 (N_29293,N_28659,N_28277);
or U29294 (N_29294,N_28457,N_28662);
nand U29295 (N_29295,N_28684,N_28406);
nand U29296 (N_29296,N_28216,N_28269);
xnor U29297 (N_29297,N_28755,N_28602);
nor U29298 (N_29298,N_28210,N_28555);
or U29299 (N_29299,N_28760,N_28356);
or U29300 (N_29300,N_28715,N_28672);
xor U29301 (N_29301,N_28773,N_28245);
nor U29302 (N_29302,N_28779,N_28664);
or U29303 (N_29303,N_28571,N_28202);
nor U29304 (N_29304,N_28222,N_28201);
nor U29305 (N_29305,N_28715,N_28432);
nor U29306 (N_29306,N_28295,N_28207);
and U29307 (N_29307,N_28474,N_28664);
nor U29308 (N_29308,N_28738,N_28616);
and U29309 (N_29309,N_28686,N_28571);
and U29310 (N_29310,N_28702,N_28490);
or U29311 (N_29311,N_28630,N_28629);
nand U29312 (N_29312,N_28522,N_28244);
nand U29313 (N_29313,N_28682,N_28324);
or U29314 (N_29314,N_28710,N_28648);
nor U29315 (N_29315,N_28758,N_28762);
nor U29316 (N_29316,N_28328,N_28252);
and U29317 (N_29317,N_28550,N_28210);
nand U29318 (N_29318,N_28293,N_28698);
nor U29319 (N_29319,N_28213,N_28256);
xnor U29320 (N_29320,N_28551,N_28405);
nand U29321 (N_29321,N_28793,N_28292);
nand U29322 (N_29322,N_28446,N_28456);
and U29323 (N_29323,N_28636,N_28541);
and U29324 (N_29324,N_28527,N_28398);
or U29325 (N_29325,N_28519,N_28552);
nor U29326 (N_29326,N_28680,N_28448);
nor U29327 (N_29327,N_28686,N_28706);
nand U29328 (N_29328,N_28599,N_28428);
xor U29329 (N_29329,N_28570,N_28511);
or U29330 (N_29330,N_28299,N_28657);
and U29331 (N_29331,N_28245,N_28574);
nand U29332 (N_29332,N_28261,N_28202);
and U29333 (N_29333,N_28498,N_28600);
nor U29334 (N_29334,N_28630,N_28314);
nor U29335 (N_29335,N_28561,N_28562);
nand U29336 (N_29336,N_28548,N_28686);
nor U29337 (N_29337,N_28210,N_28274);
xnor U29338 (N_29338,N_28486,N_28761);
xor U29339 (N_29339,N_28312,N_28384);
or U29340 (N_29340,N_28225,N_28695);
or U29341 (N_29341,N_28577,N_28572);
nand U29342 (N_29342,N_28594,N_28333);
or U29343 (N_29343,N_28467,N_28507);
or U29344 (N_29344,N_28430,N_28422);
or U29345 (N_29345,N_28678,N_28588);
nor U29346 (N_29346,N_28770,N_28588);
nand U29347 (N_29347,N_28373,N_28325);
nor U29348 (N_29348,N_28412,N_28272);
nor U29349 (N_29349,N_28579,N_28350);
xnor U29350 (N_29350,N_28721,N_28480);
or U29351 (N_29351,N_28218,N_28587);
xnor U29352 (N_29352,N_28760,N_28318);
nand U29353 (N_29353,N_28712,N_28453);
xor U29354 (N_29354,N_28307,N_28673);
nand U29355 (N_29355,N_28715,N_28377);
or U29356 (N_29356,N_28509,N_28711);
and U29357 (N_29357,N_28473,N_28615);
or U29358 (N_29358,N_28704,N_28278);
or U29359 (N_29359,N_28795,N_28369);
nor U29360 (N_29360,N_28300,N_28409);
and U29361 (N_29361,N_28639,N_28723);
xnor U29362 (N_29362,N_28423,N_28648);
nor U29363 (N_29363,N_28594,N_28666);
and U29364 (N_29364,N_28612,N_28204);
or U29365 (N_29365,N_28651,N_28553);
nor U29366 (N_29366,N_28615,N_28783);
xor U29367 (N_29367,N_28764,N_28356);
nor U29368 (N_29368,N_28416,N_28277);
nand U29369 (N_29369,N_28438,N_28745);
xor U29370 (N_29370,N_28488,N_28377);
nand U29371 (N_29371,N_28616,N_28795);
and U29372 (N_29372,N_28598,N_28425);
xnor U29373 (N_29373,N_28449,N_28277);
or U29374 (N_29374,N_28225,N_28539);
nand U29375 (N_29375,N_28506,N_28783);
nor U29376 (N_29376,N_28720,N_28790);
or U29377 (N_29377,N_28381,N_28288);
and U29378 (N_29378,N_28681,N_28321);
nand U29379 (N_29379,N_28762,N_28782);
nor U29380 (N_29380,N_28764,N_28593);
or U29381 (N_29381,N_28510,N_28784);
nand U29382 (N_29382,N_28751,N_28728);
xor U29383 (N_29383,N_28665,N_28770);
xnor U29384 (N_29384,N_28576,N_28663);
xnor U29385 (N_29385,N_28292,N_28661);
nor U29386 (N_29386,N_28300,N_28760);
nand U29387 (N_29387,N_28536,N_28237);
nand U29388 (N_29388,N_28799,N_28237);
or U29389 (N_29389,N_28304,N_28538);
or U29390 (N_29390,N_28387,N_28720);
nor U29391 (N_29391,N_28508,N_28687);
or U29392 (N_29392,N_28415,N_28332);
nand U29393 (N_29393,N_28261,N_28401);
and U29394 (N_29394,N_28362,N_28757);
xor U29395 (N_29395,N_28314,N_28548);
xor U29396 (N_29396,N_28428,N_28620);
or U29397 (N_29397,N_28694,N_28669);
and U29398 (N_29398,N_28725,N_28420);
or U29399 (N_29399,N_28409,N_28623);
and U29400 (N_29400,N_28995,N_29151);
nor U29401 (N_29401,N_29329,N_29333);
nand U29402 (N_29402,N_29399,N_28915);
nor U29403 (N_29403,N_28991,N_28969);
nor U29404 (N_29404,N_28896,N_29222);
xor U29405 (N_29405,N_29350,N_28844);
xor U29406 (N_29406,N_28968,N_29062);
and U29407 (N_29407,N_28858,N_28971);
nor U29408 (N_29408,N_29383,N_29249);
nor U29409 (N_29409,N_29189,N_29215);
and U29410 (N_29410,N_28992,N_29396);
and U29411 (N_29411,N_29261,N_29070);
and U29412 (N_29412,N_28856,N_29086);
nor U29413 (N_29413,N_28930,N_29287);
nand U29414 (N_29414,N_29094,N_28916);
nor U29415 (N_29415,N_28926,N_29243);
nor U29416 (N_29416,N_28867,N_28813);
and U29417 (N_29417,N_29015,N_28944);
or U29418 (N_29418,N_29120,N_29081);
and U29419 (N_29419,N_29105,N_29114);
nand U29420 (N_29420,N_29392,N_28846);
and U29421 (N_29421,N_29080,N_29225);
nand U29422 (N_29422,N_29233,N_29009);
and U29423 (N_29423,N_28809,N_28840);
and U29424 (N_29424,N_28989,N_29038);
nor U29425 (N_29425,N_28895,N_29027);
or U29426 (N_29426,N_28835,N_28909);
nand U29427 (N_29427,N_29369,N_29177);
nor U29428 (N_29428,N_28913,N_29072);
or U29429 (N_29429,N_29194,N_29244);
nand U29430 (N_29430,N_28817,N_29171);
nor U29431 (N_29431,N_29364,N_28990);
nand U29432 (N_29432,N_29276,N_29358);
and U29433 (N_29433,N_29008,N_28843);
nand U29434 (N_29434,N_29365,N_28839);
nand U29435 (N_29435,N_28860,N_28902);
and U29436 (N_29436,N_29272,N_28879);
nor U29437 (N_29437,N_29210,N_29326);
or U29438 (N_29438,N_29263,N_29338);
nor U29439 (N_29439,N_29061,N_28910);
and U29440 (N_29440,N_29058,N_29254);
and U29441 (N_29441,N_29273,N_28975);
nand U29442 (N_29442,N_28954,N_29197);
or U29443 (N_29443,N_29238,N_29096);
nor U29444 (N_29444,N_29057,N_28887);
nand U29445 (N_29445,N_28946,N_28830);
nor U29446 (N_29446,N_29262,N_29380);
nor U29447 (N_29447,N_28802,N_29322);
xnor U29448 (N_29448,N_29285,N_29303);
and U29449 (N_29449,N_28812,N_29306);
nand U29450 (N_29450,N_29325,N_29124);
xor U29451 (N_29451,N_29386,N_29093);
xor U29452 (N_29452,N_29252,N_28826);
nand U29453 (N_29453,N_28899,N_28934);
nor U29454 (N_29454,N_29219,N_29313);
nand U29455 (N_29455,N_29376,N_29024);
and U29456 (N_29456,N_29293,N_29107);
nand U29457 (N_29457,N_29299,N_29271);
nand U29458 (N_29458,N_29052,N_28834);
nor U29459 (N_29459,N_29095,N_28893);
nor U29460 (N_29460,N_28801,N_29394);
nor U29461 (N_29461,N_29355,N_29224);
or U29462 (N_29462,N_29278,N_29112);
xor U29463 (N_29463,N_28937,N_29368);
or U29464 (N_29464,N_28947,N_29054);
or U29465 (N_29465,N_29091,N_28862);
nor U29466 (N_29466,N_28912,N_29140);
nor U29467 (N_29467,N_29384,N_29099);
or U29468 (N_29468,N_29059,N_29314);
and U29469 (N_29469,N_28820,N_28985);
nand U29470 (N_29470,N_29268,N_29126);
and U29471 (N_29471,N_29173,N_29339);
nand U29472 (N_29472,N_28883,N_29361);
nor U29473 (N_29473,N_29362,N_29075);
nor U29474 (N_29474,N_29218,N_28850);
and U29475 (N_29475,N_28927,N_29163);
nor U29476 (N_29476,N_29315,N_29253);
or U29477 (N_29477,N_29133,N_29154);
nor U29478 (N_29478,N_29161,N_29143);
nor U29479 (N_29479,N_29257,N_29076);
and U29480 (N_29480,N_29320,N_29312);
nand U29481 (N_29481,N_29083,N_28961);
nor U29482 (N_29482,N_29235,N_28807);
and U29483 (N_29483,N_29245,N_29087);
or U29484 (N_29484,N_29341,N_29201);
or U29485 (N_29485,N_29319,N_29085);
nor U29486 (N_29486,N_29012,N_28922);
nand U29487 (N_29487,N_29385,N_28924);
nand U29488 (N_29488,N_29242,N_29007);
xnor U29489 (N_29489,N_29138,N_29018);
nand U29490 (N_29490,N_29283,N_28940);
or U29491 (N_29491,N_29296,N_29181);
or U29492 (N_29492,N_28898,N_29348);
or U29493 (N_29493,N_29041,N_29373);
and U29494 (N_29494,N_29198,N_29204);
nor U29495 (N_29495,N_29195,N_29387);
or U29496 (N_29496,N_29145,N_29367);
or U29497 (N_29497,N_29352,N_29001);
and U29498 (N_29498,N_29188,N_29005);
and U29499 (N_29499,N_28849,N_28978);
nor U29500 (N_29500,N_28859,N_29232);
and U29501 (N_29501,N_29183,N_29311);
nor U29502 (N_29502,N_29134,N_28907);
nand U29503 (N_29503,N_28966,N_28963);
and U29504 (N_29504,N_28943,N_29044);
or U29505 (N_29505,N_28806,N_29137);
and U29506 (N_29506,N_28953,N_29381);
or U29507 (N_29507,N_28933,N_28831);
nor U29508 (N_29508,N_29101,N_29020);
nand U29509 (N_29509,N_28804,N_29123);
and U29510 (N_29510,N_29398,N_29056);
nand U29511 (N_29511,N_29340,N_28837);
and U29512 (N_29512,N_28874,N_28816);
or U29513 (N_29513,N_29234,N_29220);
or U29514 (N_29514,N_29042,N_29327);
or U29515 (N_29515,N_29004,N_29088);
and U29516 (N_29516,N_29223,N_28897);
nand U29517 (N_29517,N_28894,N_29308);
or U29518 (N_29518,N_28920,N_29221);
nand U29519 (N_29519,N_28853,N_29354);
nor U29520 (N_29520,N_29184,N_28986);
or U29521 (N_29521,N_28890,N_29351);
and U29522 (N_29522,N_29214,N_28901);
and U29523 (N_29523,N_29193,N_29023);
nor U29524 (N_29524,N_29174,N_29025);
nor U29525 (N_29525,N_29344,N_28911);
or U29526 (N_29526,N_29190,N_28972);
nor U29527 (N_29527,N_29121,N_29275);
or U29528 (N_29528,N_29391,N_29168);
nor U29529 (N_29529,N_29212,N_29157);
nand U29530 (N_29530,N_29270,N_29068);
nor U29531 (N_29531,N_29342,N_28976);
or U29532 (N_29532,N_29046,N_29382);
nor U29533 (N_29533,N_29089,N_29256);
or U29534 (N_29534,N_29304,N_29192);
and U29535 (N_29535,N_29162,N_29000);
nand U29536 (N_29536,N_28960,N_29179);
nor U29537 (N_29537,N_29139,N_29282);
nor U29538 (N_29538,N_29169,N_28871);
nor U29539 (N_29539,N_28942,N_29284);
and U29540 (N_29540,N_29017,N_28983);
xnor U29541 (N_29541,N_28868,N_29251);
or U29542 (N_29542,N_29289,N_29217);
nor U29543 (N_29543,N_29265,N_29301);
and U29544 (N_29544,N_29135,N_29132);
xor U29545 (N_29545,N_29360,N_29334);
xor U29546 (N_29546,N_29090,N_28993);
xor U29547 (N_29547,N_28981,N_29034);
or U29548 (N_29548,N_28982,N_29324);
or U29549 (N_29549,N_28936,N_28938);
and U29550 (N_29550,N_28928,N_29175);
nor U29551 (N_29551,N_28889,N_28842);
nor U29552 (N_29552,N_28965,N_29371);
or U29553 (N_29553,N_28827,N_28823);
nand U29554 (N_29554,N_29337,N_29200);
nand U29555 (N_29555,N_29002,N_29307);
nand U29556 (N_29556,N_28863,N_29335);
or U29557 (N_29557,N_29021,N_28882);
or U29558 (N_29558,N_29241,N_29274);
or U29559 (N_29559,N_29206,N_29055);
or U29560 (N_29560,N_29050,N_29003);
or U29561 (N_29561,N_28908,N_28814);
nand U29562 (N_29562,N_28892,N_28905);
and U29563 (N_29563,N_28866,N_29146);
and U29564 (N_29564,N_29028,N_29259);
nor U29565 (N_29565,N_29113,N_29035);
or U29566 (N_29566,N_29064,N_29288);
and U29567 (N_29567,N_28900,N_29109);
and U29568 (N_29568,N_29202,N_29240);
or U29569 (N_29569,N_29250,N_29014);
and U29570 (N_29570,N_29116,N_29230);
or U29571 (N_29571,N_28811,N_29203);
nand U29572 (N_29572,N_28931,N_28906);
nand U29573 (N_29573,N_28872,N_29309);
xor U29574 (N_29574,N_28815,N_29353);
and U29575 (N_29575,N_28925,N_29084);
and U29576 (N_29576,N_29155,N_29305);
nor U29577 (N_29577,N_28885,N_28848);
nand U29578 (N_29578,N_29037,N_28951);
and U29579 (N_29579,N_28950,N_29049);
nor U29580 (N_29580,N_29102,N_29048);
or U29581 (N_29581,N_29266,N_29264);
or U29582 (N_29582,N_29153,N_29033);
or U29583 (N_29583,N_28855,N_29280);
nor U29584 (N_29584,N_28917,N_29228);
nand U29585 (N_29585,N_29165,N_28980);
or U29586 (N_29586,N_29029,N_29302);
and U29587 (N_29587,N_29104,N_28818);
nor U29588 (N_29588,N_28939,N_29103);
nor U29589 (N_29589,N_29331,N_28829);
or U29590 (N_29590,N_28800,N_29279);
or U29591 (N_29591,N_29281,N_29388);
nand U29592 (N_29592,N_29032,N_29150);
and U29593 (N_29593,N_28869,N_29318);
or U29594 (N_29594,N_28891,N_28956);
xnor U29595 (N_29595,N_28865,N_28870);
and U29596 (N_29596,N_29292,N_29186);
and U29597 (N_29597,N_29310,N_29164);
or U29598 (N_29598,N_29205,N_29156);
nor U29599 (N_29599,N_29073,N_28988);
or U29600 (N_29600,N_29260,N_29129);
nor U29601 (N_29601,N_28854,N_29363);
nand U29602 (N_29602,N_29269,N_28861);
xnor U29603 (N_29603,N_28952,N_29078);
nor U29604 (N_29604,N_28876,N_29239);
nand U29605 (N_29605,N_29255,N_28803);
nor U29606 (N_29606,N_28875,N_28888);
or U29607 (N_29607,N_28998,N_29393);
nor U29608 (N_29608,N_29013,N_29016);
nand U29609 (N_29609,N_29297,N_28880);
nor U29610 (N_29610,N_29097,N_29185);
or U29611 (N_29611,N_29349,N_29092);
nand U29612 (N_29612,N_29026,N_28918);
nor U29613 (N_29613,N_29328,N_28984);
and U29614 (N_29614,N_28929,N_29213);
and U29615 (N_29615,N_28878,N_29006);
nand U29616 (N_29616,N_29321,N_29236);
or U29617 (N_29617,N_29040,N_29065);
and U29618 (N_29618,N_29053,N_28886);
and U29619 (N_29619,N_29118,N_28821);
nor U29620 (N_29620,N_29182,N_28967);
nor U29621 (N_29621,N_28923,N_28949);
or U29622 (N_29622,N_29159,N_29359);
and U29623 (N_29623,N_29160,N_28970);
nand U29624 (N_29624,N_29207,N_29031);
and U29625 (N_29625,N_28999,N_28852);
or U29626 (N_29626,N_28836,N_28974);
or U29627 (N_29627,N_28832,N_28824);
or U29628 (N_29628,N_29142,N_29043);
nor U29629 (N_29629,N_29347,N_29290);
and U29630 (N_29630,N_28921,N_29128);
nor U29631 (N_29631,N_29374,N_29115);
and U29632 (N_29632,N_28945,N_28805);
or U29633 (N_29633,N_28864,N_29237);
nor U29634 (N_29634,N_29343,N_29366);
nand U29635 (N_29635,N_29036,N_29071);
and U29636 (N_29636,N_29216,N_28833);
or U29637 (N_29637,N_28914,N_29267);
and U29638 (N_29638,N_29227,N_29180);
nor U29639 (N_29639,N_29208,N_29379);
and U29640 (N_29640,N_29390,N_28847);
nor U29641 (N_29641,N_28957,N_29176);
nand U29642 (N_29642,N_29147,N_29127);
and U29643 (N_29643,N_29294,N_29247);
nor U29644 (N_29644,N_29051,N_28932);
nor U29645 (N_29645,N_28810,N_28881);
and U29646 (N_29646,N_29125,N_29063);
or U29647 (N_29647,N_29098,N_28838);
and U29648 (N_29648,N_29141,N_29248);
nand U29649 (N_29649,N_29295,N_29323);
nand U29650 (N_29650,N_29286,N_28962);
nor U29651 (N_29651,N_29144,N_29229);
or U29652 (N_29652,N_28845,N_29316);
xor U29653 (N_29653,N_29030,N_29011);
and U29654 (N_29654,N_29336,N_29356);
xnor U29655 (N_29655,N_29082,N_28884);
or U29656 (N_29656,N_29079,N_29346);
nor U29657 (N_29657,N_29231,N_28941);
or U29658 (N_29658,N_29010,N_28822);
xnor U29659 (N_29659,N_29199,N_29022);
nand U29660 (N_29660,N_28935,N_29149);
and U29661 (N_29661,N_28959,N_29166);
nand U29662 (N_29662,N_29019,N_28948);
or U29663 (N_29663,N_29332,N_29246);
nand U29664 (N_29664,N_29067,N_29122);
or U29665 (N_29665,N_28955,N_29074);
and U29666 (N_29666,N_28958,N_28994);
and U29667 (N_29667,N_29045,N_29187);
and U29668 (N_29668,N_29152,N_29209);
and U29669 (N_29669,N_28977,N_29345);
or U29670 (N_29670,N_29357,N_28964);
nand U29671 (N_29671,N_29106,N_28825);
or U29672 (N_29672,N_28997,N_29136);
nand U29673 (N_29673,N_28919,N_29178);
nand U29674 (N_29674,N_29111,N_29148);
and U29675 (N_29675,N_29377,N_28857);
nand U29676 (N_29676,N_29211,N_29378);
nor U29677 (N_29677,N_28851,N_29317);
and U29678 (N_29678,N_29108,N_29130);
nor U29679 (N_29679,N_29300,N_28819);
nor U29680 (N_29680,N_28973,N_28979);
or U29681 (N_29681,N_29131,N_29077);
or U29682 (N_29682,N_29191,N_29389);
and U29683 (N_29683,N_29291,N_29158);
nor U29684 (N_29684,N_28987,N_29370);
or U29685 (N_29685,N_29196,N_29395);
nand U29686 (N_29686,N_29226,N_29170);
and U29687 (N_29687,N_28904,N_29375);
xnor U29688 (N_29688,N_29372,N_28828);
or U29689 (N_29689,N_28873,N_29298);
or U29690 (N_29690,N_28903,N_28841);
and U29691 (N_29691,N_29047,N_29172);
nand U29692 (N_29692,N_29119,N_29277);
nor U29693 (N_29693,N_29100,N_29069);
nand U29694 (N_29694,N_29066,N_29330);
nand U29695 (N_29695,N_29039,N_29167);
or U29696 (N_29696,N_28808,N_28996);
or U29697 (N_29697,N_28877,N_29117);
and U29698 (N_29698,N_29258,N_29110);
nand U29699 (N_29699,N_29060,N_29397);
and U29700 (N_29700,N_29360,N_29062);
nor U29701 (N_29701,N_28869,N_28976);
and U29702 (N_29702,N_29368,N_28908);
nor U29703 (N_29703,N_28832,N_28925);
or U29704 (N_29704,N_28985,N_28994);
nand U29705 (N_29705,N_29014,N_29123);
or U29706 (N_29706,N_29227,N_29347);
xnor U29707 (N_29707,N_29109,N_29198);
nand U29708 (N_29708,N_28951,N_29319);
nor U29709 (N_29709,N_29002,N_29038);
nor U29710 (N_29710,N_29194,N_29218);
xnor U29711 (N_29711,N_29031,N_29161);
xor U29712 (N_29712,N_29363,N_29296);
nor U29713 (N_29713,N_28984,N_29030);
or U29714 (N_29714,N_29153,N_28911);
or U29715 (N_29715,N_29392,N_28840);
nand U29716 (N_29716,N_29371,N_28824);
or U29717 (N_29717,N_29229,N_28882);
and U29718 (N_29718,N_28841,N_29352);
and U29719 (N_29719,N_29255,N_29094);
or U29720 (N_29720,N_29301,N_28832);
xor U29721 (N_29721,N_28866,N_28919);
nor U29722 (N_29722,N_29140,N_29022);
or U29723 (N_29723,N_28947,N_29102);
and U29724 (N_29724,N_29342,N_29119);
and U29725 (N_29725,N_29224,N_28851);
nand U29726 (N_29726,N_28838,N_28818);
nor U29727 (N_29727,N_29334,N_28850);
and U29728 (N_29728,N_29195,N_29263);
nand U29729 (N_29729,N_29366,N_28987);
nand U29730 (N_29730,N_29394,N_29223);
nand U29731 (N_29731,N_29195,N_29323);
or U29732 (N_29732,N_29028,N_29133);
nand U29733 (N_29733,N_29026,N_29242);
nand U29734 (N_29734,N_29059,N_28848);
nor U29735 (N_29735,N_28804,N_29026);
nor U29736 (N_29736,N_29203,N_29230);
and U29737 (N_29737,N_28941,N_29260);
xnor U29738 (N_29738,N_29311,N_28969);
xnor U29739 (N_29739,N_28917,N_29099);
xor U29740 (N_29740,N_28925,N_29110);
nand U29741 (N_29741,N_28858,N_28905);
nor U29742 (N_29742,N_28824,N_29079);
or U29743 (N_29743,N_29346,N_28852);
nor U29744 (N_29744,N_28932,N_28819);
nand U29745 (N_29745,N_28969,N_29206);
or U29746 (N_29746,N_29177,N_28856);
nor U29747 (N_29747,N_29285,N_29009);
xor U29748 (N_29748,N_29191,N_29097);
or U29749 (N_29749,N_29028,N_29267);
and U29750 (N_29750,N_29371,N_28873);
or U29751 (N_29751,N_29009,N_29361);
and U29752 (N_29752,N_29149,N_28876);
and U29753 (N_29753,N_29056,N_29210);
and U29754 (N_29754,N_29082,N_29083);
or U29755 (N_29755,N_28813,N_29102);
and U29756 (N_29756,N_29050,N_29089);
or U29757 (N_29757,N_29020,N_28932);
nand U29758 (N_29758,N_28999,N_29370);
and U29759 (N_29759,N_28991,N_29259);
nor U29760 (N_29760,N_29195,N_29089);
nor U29761 (N_29761,N_28970,N_29261);
nand U29762 (N_29762,N_29360,N_29236);
nand U29763 (N_29763,N_29138,N_28831);
or U29764 (N_29764,N_29179,N_29188);
nor U29765 (N_29765,N_28988,N_29253);
nor U29766 (N_29766,N_28893,N_29284);
nand U29767 (N_29767,N_29236,N_29131);
nand U29768 (N_29768,N_29264,N_29227);
or U29769 (N_29769,N_28868,N_28949);
nor U29770 (N_29770,N_29310,N_29079);
nand U29771 (N_29771,N_28937,N_28823);
nand U29772 (N_29772,N_29145,N_29161);
or U29773 (N_29773,N_29119,N_28921);
nand U29774 (N_29774,N_29227,N_29003);
nand U29775 (N_29775,N_29132,N_29215);
nor U29776 (N_29776,N_28965,N_29344);
nand U29777 (N_29777,N_29398,N_29213);
and U29778 (N_29778,N_29043,N_28890);
nor U29779 (N_29779,N_28948,N_29331);
and U29780 (N_29780,N_28969,N_29319);
xor U29781 (N_29781,N_29020,N_29045);
nor U29782 (N_29782,N_29290,N_29298);
or U29783 (N_29783,N_29390,N_29124);
or U29784 (N_29784,N_29115,N_29399);
nand U29785 (N_29785,N_28929,N_29349);
and U29786 (N_29786,N_28820,N_28916);
xor U29787 (N_29787,N_28838,N_29270);
xor U29788 (N_29788,N_29087,N_29115);
nor U29789 (N_29789,N_29019,N_28865);
or U29790 (N_29790,N_29126,N_29358);
xnor U29791 (N_29791,N_29303,N_28888);
nor U29792 (N_29792,N_29109,N_29245);
nor U29793 (N_29793,N_29327,N_28919);
or U29794 (N_29794,N_29136,N_28850);
xor U29795 (N_29795,N_28871,N_29090);
nor U29796 (N_29796,N_28839,N_29185);
or U29797 (N_29797,N_29311,N_29162);
or U29798 (N_29798,N_29226,N_29335);
nand U29799 (N_29799,N_29262,N_29124);
and U29800 (N_29800,N_29356,N_29319);
or U29801 (N_29801,N_28809,N_29100);
nand U29802 (N_29802,N_29151,N_29320);
and U29803 (N_29803,N_29307,N_28814);
and U29804 (N_29804,N_28995,N_29027);
nand U29805 (N_29805,N_29305,N_28954);
and U29806 (N_29806,N_29003,N_29006);
nand U29807 (N_29807,N_29091,N_28835);
and U29808 (N_29808,N_28919,N_29036);
nor U29809 (N_29809,N_29088,N_28982);
nand U29810 (N_29810,N_29037,N_29215);
nor U29811 (N_29811,N_28813,N_29106);
nand U29812 (N_29812,N_29043,N_28804);
or U29813 (N_29813,N_29044,N_29292);
nand U29814 (N_29814,N_29086,N_29063);
or U29815 (N_29815,N_29258,N_28829);
and U29816 (N_29816,N_29282,N_29079);
nor U29817 (N_29817,N_29050,N_29075);
or U29818 (N_29818,N_29120,N_29381);
nor U29819 (N_29819,N_29171,N_29139);
and U29820 (N_29820,N_28875,N_29340);
nor U29821 (N_29821,N_29282,N_29241);
nand U29822 (N_29822,N_28891,N_28971);
and U29823 (N_29823,N_28930,N_29052);
or U29824 (N_29824,N_29124,N_29379);
nor U29825 (N_29825,N_29289,N_29039);
nand U29826 (N_29826,N_28907,N_29377);
nand U29827 (N_29827,N_29286,N_28882);
and U29828 (N_29828,N_29284,N_29254);
xor U29829 (N_29829,N_28858,N_29384);
and U29830 (N_29830,N_28883,N_29219);
nor U29831 (N_29831,N_29283,N_28844);
nand U29832 (N_29832,N_29181,N_28800);
or U29833 (N_29833,N_29073,N_28882);
and U29834 (N_29834,N_29251,N_29253);
or U29835 (N_29835,N_29271,N_29236);
nand U29836 (N_29836,N_29212,N_29192);
and U29837 (N_29837,N_29122,N_29205);
or U29838 (N_29838,N_28945,N_29101);
xor U29839 (N_29839,N_29296,N_29237);
nand U29840 (N_29840,N_29028,N_29349);
xnor U29841 (N_29841,N_29310,N_29170);
xnor U29842 (N_29842,N_28880,N_29245);
and U29843 (N_29843,N_29295,N_28860);
nand U29844 (N_29844,N_29261,N_29321);
and U29845 (N_29845,N_28945,N_29171);
and U29846 (N_29846,N_28962,N_29234);
or U29847 (N_29847,N_29060,N_28862);
nand U29848 (N_29848,N_29037,N_28948);
nor U29849 (N_29849,N_29079,N_29293);
xnor U29850 (N_29850,N_28912,N_29324);
and U29851 (N_29851,N_29305,N_28998);
or U29852 (N_29852,N_29156,N_28956);
and U29853 (N_29853,N_29263,N_29047);
or U29854 (N_29854,N_29295,N_28910);
nor U29855 (N_29855,N_29381,N_29209);
nor U29856 (N_29856,N_28824,N_29047);
or U29857 (N_29857,N_29062,N_28924);
or U29858 (N_29858,N_28940,N_29053);
or U29859 (N_29859,N_29100,N_28889);
nand U29860 (N_29860,N_28979,N_29298);
and U29861 (N_29861,N_29213,N_29346);
or U29862 (N_29862,N_28889,N_29103);
and U29863 (N_29863,N_28930,N_29279);
nor U29864 (N_29864,N_29009,N_29301);
nor U29865 (N_29865,N_29001,N_29281);
or U29866 (N_29866,N_29199,N_29207);
or U29867 (N_29867,N_29381,N_29002);
nor U29868 (N_29868,N_28896,N_29392);
xor U29869 (N_29869,N_29095,N_28898);
nor U29870 (N_29870,N_29056,N_29028);
xor U29871 (N_29871,N_29076,N_29253);
and U29872 (N_29872,N_28903,N_28942);
nand U29873 (N_29873,N_28937,N_29370);
xnor U29874 (N_29874,N_28924,N_29380);
nand U29875 (N_29875,N_29333,N_28890);
nand U29876 (N_29876,N_29079,N_29185);
nand U29877 (N_29877,N_29198,N_29096);
or U29878 (N_29878,N_29286,N_28862);
xor U29879 (N_29879,N_28904,N_29329);
nand U29880 (N_29880,N_29264,N_28865);
nor U29881 (N_29881,N_29156,N_28827);
nand U29882 (N_29882,N_29092,N_29233);
nor U29883 (N_29883,N_28876,N_29020);
nand U29884 (N_29884,N_29026,N_28984);
and U29885 (N_29885,N_29327,N_29080);
and U29886 (N_29886,N_29298,N_29309);
nor U29887 (N_29887,N_29397,N_28990);
nor U29888 (N_29888,N_29112,N_29153);
and U29889 (N_29889,N_29078,N_28855);
nand U29890 (N_29890,N_29164,N_29017);
nor U29891 (N_29891,N_29147,N_29007);
and U29892 (N_29892,N_29215,N_28874);
and U29893 (N_29893,N_29276,N_28807);
nand U29894 (N_29894,N_29053,N_29353);
xor U29895 (N_29895,N_29192,N_28823);
nand U29896 (N_29896,N_29314,N_28841);
nor U29897 (N_29897,N_28861,N_29054);
and U29898 (N_29898,N_29107,N_29122);
nand U29899 (N_29899,N_28954,N_29136);
or U29900 (N_29900,N_29205,N_29189);
nor U29901 (N_29901,N_28872,N_29057);
nor U29902 (N_29902,N_29376,N_29241);
nand U29903 (N_29903,N_29164,N_29144);
xor U29904 (N_29904,N_28902,N_28889);
and U29905 (N_29905,N_29111,N_29015);
or U29906 (N_29906,N_29335,N_29193);
nand U29907 (N_29907,N_29108,N_28912);
and U29908 (N_29908,N_29392,N_29315);
xor U29909 (N_29909,N_29288,N_28952);
or U29910 (N_29910,N_29023,N_28899);
nand U29911 (N_29911,N_29330,N_29112);
nand U29912 (N_29912,N_29393,N_29058);
and U29913 (N_29913,N_29102,N_28982);
nand U29914 (N_29914,N_29081,N_28878);
nor U29915 (N_29915,N_29214,N_29033);
nor U29916 (N_29916,N_28806,N_28893);
and U29917 (N_29917,N_28910,N_29340);
nor U29918 (N_29918,N_29068,N_29277);
or U29919 (N_29919,N_29169,N_28984);
or U29920 (N_29920,N_29244,N_29318);
nand U29921 (N_29921,N_29205,N_29148);
and U29922 (N_29922,N_28875,N_29151);
nand U29923 (N_29923,N_29194,N_29131);
or U29924 (N_29924,N_28914,N_29273);
nand U29925 (N_29925,N_28881,N_29181);
and U29926 (N_29926,N_29016,N_29025);
and U29927 (N_29927,N_29092,N_29066);
and U29928 (N_29928,N_28945,N_29295);
nor U29929 (N_29929,N_29247,N_29226);
or U29930 (N_29930,N_29370,N_29076);
xnor U29931 (N_29931,N_29245,N_29096);
and U29932 (N_29932,N_28866,N_29097);
or U29933 (N_29933,N_29025,N_29399);
nand U29934 (N_29934,N_28985,N_29196);
nand U29935 (N_29935,N_29089,N_29038);
nand U29936 (N_29936,N_29360,N_28835);
or U29937 (N_29937,N_29256,N_29219);
and U29938 (N_29938,N_29000,N_29261);
nor U29939 (N_29939,N_29218,N_28914);
nor U29940 (N_29940,N_29320,N_28949);
and U29941 (N_29941,N_28996,N_28807);
and U29942 (N_29942,N_28913,N_28984);
or U29943 (N_29943,N_29258,N_29187);
and U29944 (N_29944,N_29132,N_29232);
nor U29945 (N_29945,N_28997,N_28946);
or U29946 (N_29946,N_28964,N_29282);
xor U29947 (N_29947,N_29254,N_28969);
nor U29948 (N_29948,N_29366,N_29091);
nor U29949 (N_29949,N_28938,N_28821);
nor U29950 (N_29950,N_29278,N_29087);
and U29951 (N_29951,N_28881,N_29238);
nand U29952 (N_29952,N_29168,N_29398);
nor U29953 (N_29953,N_29314,N_29216);
nand U29954 (N_29954,N_28992,N_28962);
nor U29955 (N_29955,N_29156,N_29376);
and U29956 (N_29956,N_28970,N_29065);
or U29957 (N_29957,N_29102,N_28892);
and U29958 (N_29958,N_28969,N_29336);
nand U29959 (N_29959,N_29266,N_28961);
and U29960 (N_29960,N_28856,N_29384);
nand U29961 (N_29961,N_28861,N_29245);
nand U29962 (N_29962,N_28938,N_29075);
or U29963 (N_29963,N_29156,N_28811);
and U29964 (N_29964,N_29236,N_29232);
or U29965 (N_29965,N_29307,N_28985);
nand U29966 (N_29966,N_29035,N_28911);
and U29967 (N_29967,N_29288,N_29094);
nor U29968 (N_29968,N_29009,N_28943);
and U29969 (N_29969,N_28819,N_28889);
or U29970 (N_29970,N_29277,N_29157);
nor U29971 (N_29971,N_29237,N_28924);
nand U29972 (N_29972,N_28847,N_29117);
nor U29973 (N_29973,N_28983,N_29049);
and U29974 (N_29974,N_29209,N_29237);
or U29975 (N_29975,N_29399,N_29052);
nor U29976 (N_29976,N_28911,N_29054);
nor U29977 (N_29977,N_29262,N_29074);
nand U29978 (N_29978,N_29316,N_29339);
nand U29979 (N_29979,N_29101,N_29196);
nor U29980 (N_29980,N_29359,N_29005);
and U29981 (N_29981,N_29382,N_29136);
nand U29982 (N_29982,N_29123,N_29290);
xnor U29983 (N_29983,N_29103,N_28930);
and U29984 (N_29984,N_29032,N_29123);
nor U29985 (N_29985,N_29110,N_29103);
nor U29986 (N_29986,N_29347,N_28849);
and U29987 (N_29987,N_28813,N_29236);
nand U29988 (N_29988,N_28838,N_28968);
nor U29989 (N_29989,N_28873,N_29025);
nor U29990 (N_29990,N_29181,N_28880);
nor U29991 (N_29991,N_29331,N_28904);
or U29992 (N_29992,N_29116,N_28804);
or U29993 (N_29993,N_29022,N_28849);
xnor U29994 (N_29994,N_28984,N_29136);
nand U29995 (N_29995,N_28924,N_28891);
nor U29996 (N_29996,N_29381,N_28927);
nand U29997 (N_29997,N_29269,N_29268);
nor U29998 (N_29998,N_28995,N_29075);
nor U29999 (N_29999,N_29360,N_29335);
nor UO_0 (O_0,N_29612,N_29816);
or UO_1 (O_1,N_29731,N_29810);
or UO_2 (O_2,N_29526,N_29765);
or UO_3 (O_3,N_29912,N_29618);
or UO_4 (O_4,N_29668,N_29587);
nor UO_5 (O_5,N_29589,N_29455);
xnor UO_6 (O_6,N_29624,N_29642);
nor UO_7 (O_7,N_29702,N_29517);
and UO_8 (O_8,N_29713,N_29674);
nand UO_9 (O_9,N_29917,N_29960);
or UO_10 (O_10,N_29956,N_29959);
and UO_11 (O_11,N_29644,N_29783);
nor UO_12 (O_12,N_29716,N_29619);
xnor UO_13 (O_13,N_29954,N_29970);
nor UO_14 (O_14,N_29527,N_29724);
nand UO_15 (O_15,N_29550,N_29925);
nand UO_16 (O_16,N_29901,N_29498);
and UO_17 (O_17,N_29452,N_29634);
and UO_18 (O_18,N_29757,N_29523);
or UO_19 (O_19,N_29690,N_29659);
nand UO_20 (O_20,N_29622,N_29820);
or UO_21 (O_21,N_29617,N_29726);
xnor UO_22 (O_22,N_29836,N_29575);
nand UO_23 (O_23,N_29793,N_29483);
nor UO_24 (O_24,N_29633,N_29427);
nor UO_25 (O_25,N_29621,N_29818);
nand UO_26 (O_26,N_29808,N_29802);
and UO_27 (O_27,N_29769,N_29687);
nor UO_28 (O_28,N_29598,N_29817);
and UO_29 (O_29,N_29722,N_29999);
or UO_30 (O_30,N_29932,N_29710);
nand UO_31 (O_31,N_29748,N_29464);
nor UO_32 (O_32,N_29511,N_29800);
and UO_33 (O_33,N_29758,N_29711);
nor UO_34 (O_34,N_29682,N_29902);
nor UO_35 (O_35,N_29964,N_29775);
nor UO_36 (O_36,N_29584,N_29512);
nand UO_37 (O_37,N_29773,N_29468);
xor UO_38 (O_38,N_29777,N_29447);
nand UO_39 (O_39,N_29551,N_29503);
and UO_40 (O_40,N_29924,N_29540);
or UO_41 (O_41,N_29533,N_29840);
xor UO_42 (O_42,N_29554,N_29892);
xnor UO_43 (O_43,N_29896,N_29868);
nor UO_44 (O_44,N_29762,N_29578);
or UO_45 (O_45,N_29437,N_29654);
nand UO_46 (O_46,N_29407,N_29515);
and UO_47 (O_47,N_29418,N_29882);
xor UO_48 (O_48,N_29448,N_29566);
xnor UO_49 (O_49,N_29709,N_29691);
nand UO_50 (O_50,N_29531,N_29506);
or UO_51 (O_51,N_29862,N_29849);
nor UO_52 (O_52,N_29530,N_29522);
and UO_53 (O_53,N_29543,N_29583);
or UO_54 (O_54,N_29827,N_29423);
or UO_55 (O_55,N_29857,N_29438);
nor UO_56 (O_56,N_29978,N_29948);
nor UO_57 (O_57,N_29613,N_29981);
nor UO_58 (O_58,N_29934,N_29411);
and UO_59 (O_59,N_29994,N_29837);
xnor UO_60 (O_60,N_29648,N_29614);
and UO_61 (O_61,N_29676,N_29852);
or UO_62 (O_62,N_29694,N_29957);
nand UO_63 (O_63,N_29939,N_29847);
nand UO_64 (O_64,N_29535,N_29577);
and UO_65 (O_65,N_29927,N_29440);
or UO_66 (O_66,N_29919,N_29997);
and UO_67 (O_67,N_29824,N_29660);
and UO_68 (O_68,N_29652,N_29665);
and UO_69 (O_69,N_29737,N_29579);
nor UO_70 (O_70,N_29476,N_29456);
nor UO_71 (O_71,N_29799,N_29630);
xnor UO_72 (O_72,N_29637,N_29541);
nor UO_73 (O_73,N_29938,N_29524);
and UO_74 (O_74,N_29562,N_29560);
nand UO_75 (O_75,N_29596,N_29569);
or UO_76 (O_76,N_29843,N_29461);
and UO_77 (O_77,N_29525,N_29872);
nor UO_78 (O_78,N_29897,N_29942);
or UO_79 (O_79,N_29510,N_29628);
xor UO_80 (O_80,N_29805,N_29556);
or UO_81 (O_81,N_29558,N_29539);
or UO_82 (O_82,N_29958,N_29814);
xnor UO_83 (O_83,N_29615,N_29460);
and UO_84 (O_84,N_29663,N_29993);
nand UO_85 (O_85,N_29764,N_29638);
or UO_86 (O_86,N_29492,N_29421);
or UO_87 (O_87,N_29830,N_29565);
nand UO_88 (O_88,N_29794,N_29940);
and UO_89 (O_89,N_29721,N_29858);
nand UO_90 (O_90,N_29855,N_29479);
or UO_91 (O_91,N_29878,N_29782);
nor UO_92 (O_92,N_29792,N_29995);
and UO_93 (O_93,N_29497,N_29640);
nand UO_94 (O_94,N_29576,N_29755);
or UO_95 (O_95,N_29985,N_29671);
nand UO_96 (O_96,N_29720,N_29888);
nand UO_97 (O_97,N_29520,N_29605);
nand UO_98 (O_98,N_29428,N_29678);
and UO_99 (O_99,N_29909,N_29555);
and UO_100 (O_100,N_29686,N_29889);
nand UO_101 (O_101,N_29725,N_29867);
and UO_102 (O_102,N_29952,N_29851);
and UO_103 (O_103,N_29759,N_29600);
xnor UO_104 (O_104,N_29723,N_29951);
nor UO_105 (O_105,N_29632,N_29875);
nor UO_106 (O_106,N_29683,N_29883);
and UO_107 (O_107,N_29623,N_29935);
or UO_108 (O_108,N_29458,N_29786);
or UO_109 (O_109,N_29803,N_29705);
nor UO_110 (O_110,N_29698,N_29564);
or UO_111 (O_111,N_29974,N_29747);
nand UO_112 (O_112,N_29546,N_29751);
nand UO_113 (O_113,N_29666,N_29494);
and UO_114 (O_114,N_29839,N_29749);
nor UO_115 (O_115,N_29983,N_29491);
nand UO_116 (O_116,N_29815,N_29672);
nand UO_117 (O_117,N_29922,N_29445);
nor UO_118 (O_118,N_29753,N_29673);
and UO_119 (O_119,N_29500,N_29453);
and UO_120 (O_120,N_29863,N_29548);
nor UO_121 (O_121,N_29697,N_29403);
nand UO_122 (O_122,N_29788,N_29465);
nand UO_123 (O_123,N_29823,N_29832);
and UO_124 (O_124,N_29963,N_29886);
or UO_125 (O_125,N_29661,N_29499);
xnor UO_126 (O_126,N_29439,N_29833);
nand UO_127 (O_127,N_29881,N_29400);
and UO_128 (O_128,N_29534,N_29887);
nor UO_129 (O_129,N_29508,N_29580);
xor UO_130 (O_130,N_29821,N_29984);
nand UO_131 (O_131,N_29610,N_29410);
and UO_132 (O_132,N_29846,N_29706);
nor UO_133 (O_133,N_29923,N_29760);
or UO_134 (O_134,N_29903,N_29908);
xnor UO_135 (O_135,N_29718,N_29419);
nor UO_136 (O_136,N_29462,N_29426);
or UO_137 (O_137,N_29750,N_29544);
or UO_138 (O_138,N_29504,N_29844);
or UO_139 (O_139,N_29475,N_29944);
and UO_140 (O_140,N_29982,N_29996);
and UO_141 (O_141,N_29700,N_29953);
nand UO_142 (O_142,N_29838,N_29943);
and UO_143 (O_143,N_29485,N_29649);
and UO_144 (O_144,N_29514,N_29826);
nand UO_145 (O_145,N_29825,N_29402);
nor UO_146 (O_146,N_29732,N_29891);
and UO_147 (O_147,N_29904,N_29877);
and UO_148 (O_148,N_29568,N_29425);
nor UO_149 (O_149,N_29480,N_29860);
nor UO_150 (O_150,N_29451,N_29651);
and UO_151 (O_151,N_29443,N_29945);
nand UO_152 (O_152,N_29599,N_29928);
nand UO_153 (O_153,N_29501,N_29519);
or UO_154 (O_154,N_29906,N_29469);
and UO_155 (O_155,N_29968,N_29801);
xnor UO_156 (O_156,N_29972,N_29738);
nor UO_157 (O_157,N_29869,N_29653);
and UO_158 (O_158,N_29662,N_29975);
or UO_159 (O_159,N_29756,N_29916);
or UO_160 (O_160,N_29905,N_29433);
nand UO_161 (O_161,N_29603,N_29745);
and UO_162 (O_162,N_29899,N_29482);
nand UO_163 (O_163,N_29442,N_29845);
and UO_164 (O_164,N_29986,N_29781);
nand UO_165 (O_165,N_29717,N_29636);
nand UO_166 (O_166,N_29620,N_29937);
and UO_167 (O_167,N_29629,N_29696);
xnor UO_168 (O_168,N_29449,N_29571);
nor UO_169 (O_169,N_29518,N_29656);
or UO_170 (O_170,N_29557,N_29645);
xnor UO_171 (O_171,N_29429,N_29703);
nor UO_172 (O_172,N_29595,N_29474);
nand UO_173 (O_173,N_29812,N_29992);
nor UO_174 (O_174,N_29414,N_29549);
nor UO_175 (O_175,N_29563,N_29704);
xor UO_176 (O_176,N_29987,N_29627);
or UO_177 (O_177,N_29693,N_29763);
and UO_178 (O_178,N_29488,N_29797);
nand UO_179 (O_179,N_29790,N_29741);
or UO_180 (O_180,N_29733,N_29911);
xnor UO_181 (O_181,N_29424,N_29772);
nand UO_182 (O_182,N_29477,N_29767);
and UO_183 (O_183,N_29873,N_29936);
or UO_184 (O_184,N_29980,N_29695);
or UO_185 (O_185,N_29921,N_29545);
nand UO_186 (O_186,N_29890,N_29798);
and UO_187 (O_187,N_29606,N_29412);
nor UO_188 (O_188,N_29967,N_29454);
or UO_189 (O_189,N_29910,N_29865);
and UO_190 (O_190,N_29719,N_29505);
nand UO_191 (O_191,N_29989,N_29949);
nand UO_192 (O_192,N_29417,N_29728);
or UO_193 (O_193,N_29876,N_29470);
or UO_194 (O_194,N_29626,N_29941);
or UO_195 (O_195,N_29898,N_29708);
or UO_196 (O_196,N_29643,N_29658);
xnor UO_197 (O_197,N_29684,N_29679);
nand UO_198 (O_198,N_29639,N_29692);
and UO_199 (O_199,N_29528,N_29971);
nor UO_200 (O_200,N_29593,N_29813);
nor UO_201 (O_201,N_29574,N_29413);
nand UO_202 (O_202,N_29736,N_29707);
xor UO_203 (O_203,N_29486,N_29879);
xor UO_204 (O_204,N_29408,N_29913);
or UO_205 (O_205,N_29553,N_29570);
nor UO_206 (O_206,N_29436,N_29866);
nand UO_207 (O_207,N_29609,N_29594);
or UO_208 (O_208,N_29406,N_29842);
and UO_209 (O_209,N_29804,N_29730);
nand UO_210 (O_210,N_29536,N_29493);
and UO_211 (O_211,N_29946,N_29787);
nor UO_212 (O_212,N_29415,N_29680);
nand UO_213 (O_213,N_29822,N_29495);
nand UO_214 (O_214,N_29784,N_29516);
nor UO_215 (O_215,N_29715,N_29667);
or UO_216 (O_216,N_29885,N_29586);
or UO_217 (O_217,N_29988,N_29740);
nor UO_218 (O_218,N_29647,N_29914);
nand UO_219 (O_219,N_29870,N_29752);
or UO_220 (O_220,N_29601,N_29743);
or UO_221 (O_221,N_29796,N_29604);
nor UO_222 (O_222,N_29559,N_29547);
nand UO_223 (O_223,N_29607,N_29854);
or UO_224 (O_224,N_29795,N_29831);
nand UO_225 (O_225,N_29920,N_29467);
or UO_226 (O_226,N_29859,N_29807);
nand UO_227 (O_227,N_29509,N_29611);
or UO_228 (O_228,N_29466,N_29727);
or UO_229 (O_229,N_29746,N_29496);
nor UO_230 (O_230,N_29655,N_29789);
and UO_231 (O_231,N_29635,N_29712);
nor UO_232 (O_232,N_29532,N_29699);
nand UO_233 (O_233,N_29616,N_29597);
or UO_234 (O_234,N_29998,N_29701);
xor UO_235 (O_235,N_29809,N_29537);
nand UO_236 (O_236,N_29441,N_29471);
or UO_237 (O_237,N_29864,N_29669);
and UO_238 (O_238,N_29582,N_29489);
nor UO_239 (O_239,N_29894,N_29401);
or UO_240 (O_240,N_29561,N_29538);
or UO_241 (O_241,N_29947,N_29969);
xor UO_242 (O_242,N_29893,N_29856);
and UO_243 (O_243,N_29435,N_29572);
nor UO_244 (O_244,N_29588,N_29965);
nor UO_245 (O_245,N_29729,N_29895);
or UO_246 (O_246,N_29871,N_29472);
or UO_247 (O_247,N_29432,N_29608);
or UO_248 (O_248,N_29675,N_29774);
or UO_249 (O_249,N_29507,N_29689);
nor UO_250 (O_250,N_29734,N_29444);
and UO_251 (O_251,N_29585,N_29819);
and UO_252 (O_252,N_29446,N_29779);
nor UO_253 (O_253,N_29950,N_29677);
xnor UO_254 (O_254,N_29529,N_29918);
nand UO_255 (O_255,N_29513,N_29961);
or UO_256 (O_256,N_29646,N_29834);
and UO_257 (O_257,N_29930,N_29811);
nand UO_258 (O_258,N_29766,N_29739);
nand UO_259 (O_259,N_29434,N_29431);
nand UO_260 (O_260,N_29592,N_29430);
or UO_261 (O_261,N_29552,N_29567);
and UO_262 (O_262,N_29991,N_29478);
nor UO_263 (O_263,N_29776,N_29742);
nand UO_264 (O_264,N_29521,N_29900);
nor UO_265 (O_265,N_29768,N_29602);
nand UO_266 (O_266,N_29581,N_29966);
or UO_267 (O_267,N_29405,N_29990);
nor UO_268 (O_268,N_29778,N_29907);
nand UO_269 (O_269,N_29962,N_29976);
xnor UO_270 (O_270,N_29422,N_29977);
and UO_271 (O_271,N_29487,N_29880);
nand UO_272 (O_272,N_29735,N_29841);
or UO_273 (O_273,N_29484,N_29785);
or UO_274 (O_274,N_29850,N_29463);
nand UO_275 (O_275,N_29473,N_29780);
nand UO_276 (O_276,N_29459,N_29926);
or UO_277 (O_277,N_29641,N_29657);
nand UO_278 (O_278,N_29542,N_29457);
nand UO_279 (O_279,N_29955,N_29979);
nor UO_280 (O_280,N_29861,N_29591);
xor UO_281 (O_281,N_29744,N_29409);
or UO_282 (O_282,N_29502,N_29848);
xor UO_283 (O_283,N_29481,N_29828);
or UO_284 (O_284,N_29931,N_29829);
or UO_285 (O_285,N_29404,N_29973);
xor UO_286 (O_286,N_29416,N_29915);
and UO_287 (O_287,N_29688,N_29685);
or UO_288 (O_288,N_29884,N_29573);
nand UO_289 (O_289,N_29933,N_29874);
nor UO_290 (O_290,N_29625,N_29681);
or UO_291 (O_291,N_29450,N_29791);
nand UO_292 (O_292,N_29761,N_29490);
xnor UO_293 (O_293,N_29770,N_29650);
and UO_294 (O_294,N_29853,N_29664);
nand UO_295 (O_295,N_29631,N_29754);
and UO_296 (O_296,N_29835,N_29670);
nor UO_297 (O_297,N_29929,N_29590);
and UO_298 (O_298,N_29806,N_29714);
nor UO_299 (O_299,N_29771,N_29420);
nand UO_300 (O_300,N_29402,N_29534);
or UO_301 (O_301,N_29640,N_29636);
nor UO_302 (O_302,N_29791,N_29805);
nand UO_303 (O_303,N_29925,N_29735);
nor UO_304 (O_304,N_29400,N_29518);
nand UO_305 (O_305,N_29907,N_29961);
nand UO_306 (O_306,N_29567,N_29669);
nand UO_307 (O_307,N_29889,N_29458);
or UO_308 (O_308,N_29568,N_29854);
and UO_309 (O_309,N_29880,N_29799);
and UO_310 (O_310,N_29543,N_29484);
nor UO_311 (O_311,N_29735,N_29746);
nand UO_312 (O_312,N_29517,N_29646);
or UO_313 (O_313,N_29699,N_29814);
or UO_314 (O_314,N_29712,N_29506);
or UO_315 (O_315,N_29894,N_29546);
or UO_316 (O_316,N_29475,N_29523);
nor UO_317 (O_317,N_29698,N_29413);
nand UO_318 (O_318,N_29889,N_29838);
or UO_319 (O_319,N_29452,N_29839);
nand UO_320 (O_320,N_29963,N_29910);
nor UO_321 (O_321,N_29823,N_29678);
xnor UO_322 (O_322,N_29623,N_29774);
or UO_323 (O_323,N_29813,N_29991);
or UO_324 (O_324,N_29987,N_29637);
nand UO_325 (O_325,N_29452,N_29691);
or UO_326 (O_326,N_29842,N_29555);
nor UO_327 (O_327,N_29932,N_29572);
nor UO_328 (O_328,N_29460,N_29640);
nor UO_329 (O_329,N_29569,N_29869);
and UO_330 (O_330,N_29601,N_29462);
nand UO_331 (O_331,N_29598,N_29420);
nand UO_332 (O_332,N_29413,N_29801);
xnor UO_333 (O_333,N_29423,N_29863);
or UO_334 (O_334,N_29429,N_29799);
nor UO_335 (O_335,N_29686,N_29528);
and UO_336 (O_336,N_29540,N_29987);
nor UO_337 (O_337,N_29478,N_29476);
nor UO_338 (O_338,N_29713,N_29571);
nor UO_339 (O_339,N_29461,N_29480);
nand UO_340 (O_340,N_29710,N_29435);
nand UO_341 (O_341,N_29920,N_29704);
or UO_342 (O_342,N_29706,N_29531);
nor UO_343 (O_343,N_29675,N_29896);
or UO_344 (O_344,N_29645,N_29707);
xor UO_345 (O_345,N_29633,N_29526);
or UO_346 (O_346,N_29582,N_29560);
and UO_347 (O_347,N_29928,N_29959);
or UO_348 (O_348,N_29605,N_29962);
nor UO_349 (O_349,N_29484,N_29877);
nand UO_350 (O_350,N_29919,N_29401);
nand UO_351 (O_351,N_29969,N_29839);
nand UO_352 (O_352,N_29499,N_29683);
nor UO_353 (O_353,N_29650,N_29847);
or UO_354 (O_354,N_29986,N_29977);
nand UO_355 (O_355,N_29991,N_29645);
xor UO_356 (O_356,N_29596,N_29674);
xor UO_357 (O_357,N_29580,N_29797);
nand UO_358 (O_358,N_29864,N_29441);
nand UO_359 (O_359,N_29584,N_29985);
nor UO_360 (O_360,N_29870,N_29861);
nor UO_361 (O_361,N_29435,N_29400);
nand UO_362 (O_362,N_29597,N_29653);
or UO_363 (O_363,N_29882,N_29425);
nand UO_364 (O_364,N_29756,N_29837);
or UO_365 (O_365,N_29404,N_29674);
nor UO_366 (O_366,N_29772,N_29527);
xor UO_367 (O_367,N_29650,N_29659);
nor UO_368 (O_368,N_29623,N_29537);
or UO_369 (O_369,N_29536,N_29734);
nand UO_370 (O_370,N_29969,N_29939);
xor UO_371 (O_371,N_29602,N_29773);
nand UO_372 (O_372,N_29653,N_29847);
or UO_373 (O_373,N_29482,N_29815);
nor UO_374 (O_374,N_29680,N_29405);
nor UO_375 (O_375,N_29935,N_29758);
nand UO_376 (O_376,N_29568,N_29402);
and UO_377 (O_377,N_29691,N_29589);
or UO_378 (O_378,N_29642,N_29764);
or UO_379 (O_379,N_29707,N_29834);
and UO_380 (O_380,N_29906,N_29548);
nor UO_381 (O_381,N_29526,N_29427);
or UO_382 (O_382,N_29955,N_29783);
and UO_383 (O_383,N_29659,N_29530);
nor UO_384 (O_384,N_29561,N_29845);
nand UO_385 (O_385,N_29791,N_29881);
or UO_386 (O_386,N_29576,N_29657);
or UO_387 (O_387,N_29703,N_29584);
or UO_388 (O_388,N_29596,N_29937);
nand UO_389 (O_389,N_29643,N_29947);
nand UO_390 (O_390,N_29850,N_29987);
or UO_391 (O_391,N_29543,N_29499);
nor UO_392 (O_392,N_29711,N_29975);
nor UO_393 (O_393,N_29679,N_29677);
nand UO_394 (O_394,N_29913,N_29676);
or UO_395 (O_395,N_29947,N_29449);
and UO_396 (O_396,N_29815,N_29550);
and UO_397 (O_397,N_29915,N_29536);
or UO_398 (O_398,N_29744,N_29880);
nor UO_399 (O_399,N_29940,N_29968);
nand UO_400 (O_400,N_29865,N_29774);
or UO_401 (O_401,N_29566,N_29635);
nand UO_402 (O_402,N_29755,N_29537);
nor UO_403 (O_403,N_29710,N_29998);
nor UO_404 (O_404,N_29868,N_29955);
nand UO_405 (O_405,N_29850,N_29577);
and UO_406 (O_406,N_29679,N_29932);
nand UO_407 (O_407,N_29477,N_29900);
nand UO_408 (O_408,N_29666,N_29439);
nand UO_409 (O_409,N_29559,N_29555);
and UO_410 (O_410,N_29584,N_29737);
nor UO_411 (O_411,N_29867,N_29976);
or UO_412 (O_412,N_29647,N_29622);
or UO_413 (O_413,N_29404,N_29419);
and UO_414 (O_414,N_29832,N_29461);
and UO_415 (O_415,N_29621,N_29442);
nand UO_416 (O_416,N_29495,N_29522);
and UO_417 (O_417,N_29665,N_29432);
and UO_418 (O_418,N_29677,N_29985);
and UO_419 (O_419,N_29575,N_29672);
and UO_420 (O_420,N_29544,N_29588);
nand UO_421 (O_421,N_29465,N_29829);
xor UO_422 (O_422,N_29411,N_29693);
or UO_423 (O_423,N_29599,N_29963);
nand UO_424 (O_424,N_29506,N_29825);
nand UO_425 (O_425,N_29424,N_29561);
xnor UO_426 (O_426,N_29553,N_29657);
nor UO_427 (O_427,N_29977,N_29616);
nor UO_428 (O_428,N_29748,N_29949);
or UO_429 (O_429,N_29734,N_29701);
or UO_430 (O_430,N_29402,N_29964);
or UO_431 (O_431,N_29604,N_29786);
and UO_432 (O_432,N_29747,N_29923);
xor UO_433 (O_433,N_29760,N_29691);
nand UO_434 (O_434,N_29531,N_29922);
nand UO_435 (O_435,N_29711,N_29743);
and UO_436 (O_436,N_29403,N_29731);
nand UO_437 (O_437,N_29956,N_29451);
nand UO_438 (O_438,N_29830,N_29621);
nand UO_439 (O_439,N_29650,N_29457);
or UO_440 (O_440,N_29717,N_29976);
nor UO_441 (O_441,N_29642,N_29800);
nand UO_442 (O_442,N_29751,N_29808);
nor UO_443 (O_443,N_29678,N_29512);
or UO_444 (O_444,N_29851,N_29961);
nand UO_445 (O_445,N_29606,N_29999);
or UO_446 (O_446,N_29795,N_29817);
and UO_447 (O_447,N_29582,N_29402);
or UO_448 (O_448,N_29592,N_29953);
nor UO_449 (O_449,N_29879,N_29710);
and UO_450 (O_450,N_29886,N_29596);
nand UO_451 (O_451,N_29431,N_29626);
and UO_452 (O_452,N_29680,N_29504);
nand UO_453 (O_453,N_29826,N_29741);
nor UO_454 (O_454,N_29526,N_29541);
nand UO_455 (O_455,N_29589,N_29477);
nand UO_456 (O_456,N_29500,N_29442);
nand UO_457 (O_457,N_29650,N_29517);
xnor UO_458 (O_458,N_29743,N_29881);
nand UO_459 (O_459,N_29621,N_29678);
and UO_460 (O_460,N_29528,N_29448);
nand UO_461 (O_461,N_29545,N_29595);
and UO_462 (O_462,N_29826,N_29495);
or UO_463 (O_463,N_29697,N_29400);
and UO_464 (O_464,N_29978,N_29502);
nand UO_465 (O_465,N_29802,N_29657);
and UO_466 (O_466,N_29748,N_29826);
and UO_467 (O_467,N_29460,N_29534);
or UO_468 (O_468,N_29546,N_29904);
and UO_469 (O_469,N_29866,N_29504);
nand UO_470 (O_470,N_29826,N_29441);
xnor UO_471 (O_471,N_29795,N_29468);
nor UO_472 (O_472,N_29854,N_29497);
and UO_473 (O_473,N_29908,N_29686);
nand UO_474 (O_474,N_29450,N_29897);
or UO_475 (O_475,N_29717,N_29493);
nor UO_476 (O_476,N_29880,N_29899);
nand UO_477 (O_477,N_29713,N_29670);
nor UO_478 (O_478,N_29631,N_29874);
or UO_479 (O_479,N_29993,N_29722);
nor UO_480 (O_480,N_29753,N_29418);
xor UO_481 (O_481,N_29433,N_29925);
nor UO_482 (O_482,N_29887,N_29526);
or UO_483 (O_483,N_29943,N_29682);
nor UO_484 (O_484,N_29616,N_29543);
nor UO_485 (O_485,N_29816,N_29787);
nand UO_486 (O_486,N_29946,N_29429);
and UO_487 (O_487,N_29538,N_29534);
and UO_488 (O_488,N_29539,N_29816);
xnor UO_489 (O_489,N_29421,N_29954);
and UO_490 (O_490,N_29494,N_29865);
or UO_491 (O_491,N_29818,N_29882);
or UO_492 (O_492,N_29552,N_29995);
or UO_493 (O_493,N_29555,N_29725);
xor UO_494 (O_494,N_29467,N_29698);
nand UO_495 (O_495,N_29576,N_29508);
and UO_496 (O_496,N_29981,N_29744);
or UO_497 (O_497,N_29886,N_29988);
or UO_498 (O_498,N_29544,N_29924);
xnor UO_499 (O_499,N_29425,N_29847);
nand UO_500 (O_500,N_29443,N_29786);
nand UO_501 (O_501,N_29463,N_29485);
nand UO_502 (O_502,N_29919,N_29884);
xnor UO_503 (O_503,N_29451,N_29776);
and UO_504 (O_504,N_29684,N_29836);
nand UO_505 (O_505,N_29991,N_29628);
nor UO_506 (O_506,N_29768,N_29656);
xor UO_507 (O_507,N_29510,N_29595);
xnor UO_508 (O_508,N_29471,N_29902);
xor UO_509 (O_509,N_29905,N_29698);
xor UO_510 (O_510,N_29652,N_29868);
and UO_511 (O_511,N_29424,N_29663);
nor UO_512 (O_512,N_29813,N_29899);
or UO_513 (O_513,N_29542,N_29563);
and UO_514 (O_514,N_29791,N_29891);
nor UO_515 (O_515,N_29770,N_29630);
nor UO_516 (O_516,N_29772,N_29874);
nor UO_517 (O_517,N_29401,N_29656);
nand UO_518 (O_518,N_29658,N_29846);
and UO_519 (O_519,N_29472,N_29963);
and UO_520 (O_520,N_29735,N_29877);
or UO_521 (O_521,N_29718,N_29875);
nor UO_522 (O_522,N_29859,N_29604);
nand UO_523 (O_523,N_29805,N_29780);
nand UO_524 (O_524,N_29855,N_29886);
nor UO_525 (O_525,N_29833,N_29815);
nor UO_526 (O_526,N_29530,N_29883);
nor UO_527 (O_527,N_29897,N_29690);
nand UO_528 (O_528,N_29542,N_29897);
nor UO_529 (O_529,N_29533,N_29851);
or UO_530 (O_530,N_29409,N_29674);
nor UO_531 (O_531,N_29580,N_29950);
nand UO_532 (O_532,N_29851,N_29847);
or UO_533 (O_533,N_29592,N_29586);
nor UO_534 (O_534,N_29902,N_29572);
nand UO_535 (O_535,N_29503,N_29960);
xnor UO_536 (O_536,N_29670,N_29744);
and UO_537 (O_537,N_29967,N_29635);
and UO_538 (O_538,N_29682,N_29491);
nor UO_539 (O_539,N_29507,N_29724);
or UO_540 (O_540,N_29468,N_29870);
xnor UO_541 (O_541,N_29400,N_29901);
or UO_542 (O_542,N_29525,N_29519);
xor UO_543 (O_543,N_29467,N_29476);
nand UO_544 (O_544,N_29692,N_29664);
or UO_545 (O_545,N_29992,N_29736);
and UO_546 (O_546,N_29723,N_29823);
nand UO_547 (O_547,N_29978,N_29553);
and UO_548 (O_548,N_29461,N_29415);
nor UO_549 (O_549,N_29555,N_29806);
nor UO_550 (O_550,N_29661,N_29487);
nand UO_551 (O_551,N_29778,N_29667);
or UO_552 (O_552,N_29727,N_29405);
nand UO_553 (O_553,N_29702,N_29801);
or UO_554 (O_554,N_29797,N_29857);
and UO_555 (O_555,N_29810,N_29756);
nand UO_556 (O_556,N_29558,N_29870);
and UO_557 (O_557,N_29895,N_29696);
or UO_558 (O_558,N_29817,N_29850);
nor UO_559 (O_559,N_29974,N_29529);
nand UO_560 (O_560,N_29697,N_29777);
or UO_561 (O_561,N_29567,N_29710);
or UO_562 (O_562,N_29574,N_29448);
nand UO_563 (O_563,N_29643,N_29668);
xor UO_564 (O_564,N_29489,N_29626);
or UO_565 (O_565,N_29742,N_29511);
and UO_566 (O_566,N_29690,N_29650);
and UO_567 (O_567,N_29734,N_29554);
and UO_568 (O_568,N_29819,N_29705);
and UO_569 (O_569,N_29529,N_29712);
nor UO_570 (O_570,N_29968,N_29975);
or UO_571 (O_571,N_29593,N_29843);
or UO_572 (O_572,N_29622,N_29881);
or UO_573 (O_573,N_29828,N_29875);
and UO_574 (O_574,N_29491,N_29938);
nand UO_575 (O_575,N_29924,N_29791);
or UO_576 (O_576,N_29761,N_29725);
nand UO_577 (O_577,N_29476,N_29616);
and UO_578 (O_578,N_29825,N_29944);
and UO_579 (O_579,N_29408,N_29865);
xor UO_580 (O_580,N_29987,N_29807);
and UO_581 (O_581,N_29481,N_29820);
or UO_582 (O_582,N_29556,N_29801);
nor UO_583 (O_583,N_29803,N_29760);
or UO_584 (O_584,N_29621,N_29629);
nand UO_585 (O_585,N_29446,N_29623);
or UO_586 (O_586,N_29979,N_29664);
or UO_587 (O_587,N_29771,N_29700);
and UO_588 (O_588,N_29561,N_29617);
xor UO_589 (O_589,N_29733,N_29491);
nand UO_590 (O_590,N_29978,N_29957);
and UO_591 (O_591,N_29696,N_29554);
nor UO_592 (O_592,N_29872,N_29901);
xor UO_593 (O_593,N_29907,N_29722);
nand UO_594 (O_594,N_29955,N_29563);
nor UO_595 (O_595,N_29734,N_29750);
nor UO_596 (O_596,N_29938,N_29834);
nand UO_597 (O_597,N_29970,N_29801);
nand UO_598 (O_598,N_29976,N_29926);
or UO_599 (O_599,N_29905,N_29975);
and UO_600 (O_600,N_29542,N_29765);
nand UO_601 (O_601,N_29597,N_29855);
or UO_602 (O_602,N_29930,N_29795);
or UO_603 (O_603,N_29572,N_29698);
and UO_604 (O_604,N_29434,N_29641);
xor UO_605 (O_605,N_29572,N_29645);
nand UO_606 (O_606,N_29507,N_29950);
nor UO_607 (O_607,N_29969,N_29694);
or UO_608 (O_608,N_29817,N_29509);
nand UO_609 (O_609,N_29875,N_29806);
nor UO_610 (O_610,N_29902,N_29862);
and UO_611 (O_611,N_29734,N_29546);
nand UO_612 (O_612,N_29861,N_29668);
nor UO_613 (O_613,N_29942,N_29507);
or UO_614 (O_614,N_29749,N_29746);
and UO_615 (O_615,N_29725,N_29926);
nor UO_616 (O_616,N_29626,N_29652);
and UO_617 (O_617,N_29860,N_29527);
nor UO_618 (O_618,N_29603,N_29688);
or UO_619 (O_619,N_29697,N_29607);
nand UO_620 (O_620,N_29492,N_29638);
nand UO_621 (O_621,N_29796,N_29460);
nor UO_622 (O_622,N_29760,N_29489);
and UO_623 (O_623,N_29454,N_29670);
nand UO_624 (O_624,N_29761,N_29704);
or UO_625 (O_625,N_29869,N_29836);
nor UO_626 (O_626,N_29474,N_29721);
xor UO_627 (O_627,N_29986,N_29631);
nor UO_628 (O_628,N_29922,N_29697);
or UO_629 (O_629,N_29930,N_29944);
nor UO_630 (O_630,N_29747,N_29690);
and UO_631 (O_631,N_29884,N_29656);
or UO_632 (O_632,N_29492,N_29956);
or UO_633 (O_633,N_29961,N_29632);
nand UO_634 (O_634,N_29844,N_29935);
nor UO_635 (O_635,N_29467,N_29758);
and UO_636 (O_636,N_29664,N_29925);
nor UO_637 (O_637,N_29425,N_29698);
and UO_638 (O_638,N_29801,N_29520);
xor UO_639 (O_639,N_29713,N_29667);
nand UO_640 (O_640,N_29465,N_29421);
and UO_641 (O_641,N_29756,N_29585);
or UO_642 (O_642,N_29689,N_29550);
nand UO_643 (O_643,N_29755,N_29613);
or UO_644 (O_644,N_29561,N_29625);
nor UO_645 (O_645,N_29741,N_29457);
and UO_646 (O_646,N_29517,N_29487);
and UO_647 (O_647,N_29470,N_29949);
and UO_648 (O_648,N_29425,N_29497);
and UO_649 (O_649,N_29979,N_29427);
nor UO_650 (O_650,N_29637,N_29627);
and UO_651 (O_651,N_29944,N_29875);
nor UO_652 (O_652,N_29889,N_29786);
nand UO_653 (O_653,N_29478,N_29811);
nand UO_654 (O_654,N_29867,N_29449);
and UO_655 (O_655,N_29468,N_29963);
nor UO_656 (O_656,N_29476,N_29427);
and UO_657 (O_657,N_29402,N_29909);
or UO_658 (O_658,N_29515,N_29406);
nor UO_659 (O_659,N_29937,N_29998);
nor UO_660 (O_660,N_29882,N_29617);
or UO_661 (O_661,N_29689,N_29579);
nor UO_662 (O_662,N_29924,N_29424);
and UO_663 (O_663,N_29564,N_29499);
and UO_664 (O_664,N_29578,N_29517);
nor UO_665 (O_665,N_29929,N_29819);
nand UO_666 (O_666,N_29741,N_29918);
and UO_667 (O_667,N_29922,N_29646);
and UO_668 (O_668,N_29560,N_29958);
and UO_669 (O_669,N_29831,N_29815);
and UO_670 (O_670,N_29609,N_29498);
or UO_671 (O_671,N_29402,N_29412);
nand UO_672 (O_672,N_29612,N_29784);
nand UO_673 (O_673,N_29965,N_29925);
or UO_674 (O_674,N_29781,N_29576);
nand UO_675 (O_675,N_29812,N_29973);
and UO_676 (O_676,N_29795,N_29835);
nand UO_677 (O_677,N_29952,N_29899);
xor UO_678 (O_678,N_29900,N_29909);
nor UO_679 (O_679,N_29652,N_29634);
nor UO_680 (O_680,N_29576,N_29902);
nor UO_681 (O_681,N_29681,N_29741);
nor UO_682 (O_682,N_29766,N_29404);
nor UO_683 (O_683,N_29670,N_29456);
nor UO_684 (O_684,N_29400,N_29792);
nor UO_685 (O_685,N_29914,N_29613);
nand UO_686 (O_686,N_29790,N_29964);
or UO_687 (O_687,N_29953,N_29996);
nor UO_688 (O_688,N_29946,N_29880);
nor UO_689 (O_689,N_29597,N_29721);
nand UO_690 (O_690,N_29901,N_29861);
and UO_691 (O_691,N_29882,N_29685);
or UO_692 (O_692,N_29617,N_29773);
or UO_693 (O_693,N_29844,N_29756);
nor UO_694 (O_694,N_29739,N_29573);
and UO_695 (O_695,N_29665,N_29408);
or UO_696 (O_696,N_29574,N_29496);
nor UO_697 (O_697,N_29872,N_29666);
nor UO_698 (O_698,N_29442,N_29420);
xor UO_699 (O_699,N_29629,N_29400);
or UO_700 (O_700,N_29882,N_29605);
and UO_701 (O_701,N_29651,N_29838);
xor UO_702 (O_702,N_29932,N_29866);
nor UO_703 (O_703,N_29574,N_29443);
and UO_704 (O_704,N_29958,N_29713);
nor UO_705 (O_705,N_29403,N_29505);
or UO_706 (O_706,N_29922,N_29682);
and UO_707 (O_707,N_29659,N_29685);
or UO_708 (O_708,N_29476,N_29608);
or UO_709 (O_709,N_29663,N_29742);
or UO_710 (O_710,N_29414,N_29481);
or UO_711 (O_711,N_29499,N_29868);
or UO_712 (O_712,N_29566,N_29815);
xor UO_713 (O_713,N_29996,N_29421);
nand UO_714 (O_714,N_29470,N_29861);
and UO_715 (O_715,N_29687,N_29976);
and UO_716 (O_716,N_29960,N_29535);
xor UO_717 (O_717,N_29849,N_29732);
or UO_718 (O_718,N_29832,N_29463);
nor UO_719 (O_719,N_29470,N_29538);
nor UO_720 (O_720,N_29596,N_29827);
xnor UO_721 (O_721,N_29489,N_29801);
and UO_722 (O_722,N_29454,N_29496);
nor UO_723 (O_723,N_29914,N_29639);
or UO_724 (O_724,N_29560,N_29670);
and UO_725 (O_725,N_29583,N_29892);
xnor UO_726 (O_726,N_29528,N_29867);
and UO_727 (O_727,N_29702,N_29878);
nand UO_728 (O_728,N_29747,N_29836);
or UO_729 (O_729,N_29735,N_29401);
nor UO_730 (O_730,N_29852,N_29933);
or UO_731 (O_731,N_29934,N_29694);
xnor UO_732 (O_732,N_29932,N_29863);
nor UO_733 (O_733,N_29504,N_29877);
and UO_734 (O_734,N_29773,N_29663);
or UO_735 (O_735,N_29576,N_29497);
nand UO_736 (O_736,N_29587,N_29770);
nor UO_737 (O_737,N_29655,N_29935);
or UO_738 (O_738,N_29423,N_29544);
nor UO_739 (O_739,N_29739,N_29507);
or UO_740 (O_740,N_29569,N_29995);
or UO_741 (O_741,N_29629,N_29770);
and UO_742 (O_742,N_29730,N_29820);
xnor UO_743 (O_743,N_29760,N_29742);
nand UO_744 (O_744,N_29744,N_29902);
nand UO_745 (O_745,N_29660,N_29971);
nand UO_746 (O_746,N_29822,N_29407);
nor UO_747 (O_747,N_29597,N_29694);
and UO_748 (O_748,N_29608,N_29455);
nor UO_749 (O_749,N_29697,N_29873);
or UO_750 (O_750,N_29743,N_29501);
or UO_751 (O_751,N_29613,N_29928);
or UO_752 (O_752,N_29526,N_29590);
nor UO_753 (O_753,N_29948,N_29718);
nand UO_754 (O_754,N_29812,N_29722);
nand UO_755 (O_755,N_29543,N_29714);
or UO_756 (O_756,N_29587,N_29848);
nand UO_757 (O_757,N_29510,N_29598);
nand UO_758 (O_758,N_29572,N_29617);
nor UO_759 (O_759,N_29426,N_29758);
and UO_760 (O_760,N_29566,N_29987);
and UO_761 (O_761,N_29851,N_29878);
nand UO_762 (O_762,N_29453,N_29527);
or UO_763 (O_763,N_29962,N_29453);
and UO_764 (O_764,N_29414,N_29724);
or UO_765 (O_765,N_29875,N_29465);
nor UO_766 (O_766,N_29428,N_29760);
nor UO_767 (O_767,N_29697,N_29783);
nand UO_768 (O_768,N_29865,N_29888);
or UO_769 (O_769,N_29418,N_29965);
nor UO_770 (O_770,N_29687,N_29958);
nor UO_771 (O_771,N_29769,N_29721);
and UO_772 (O_772,N_29675,N_29754);
nor UO_773 (O_773,N_29924,N_29768);
nand UO_774 (O_774,N_29592,N_29640);
and UO_775 (O_775,N_29668,N_29898);
nor UO_776 (O_776,N_29831,N_29819);
nand UO_777 (O_777,N_29984,N_29782);
and UO_778 (O_778,N_29720,N_29426);
xor UO_779 (O_779,N_29615,N_29906);
xnor UO_780 (O_780,N_29850,N_29616);
nor UO_781 (O_781,N_29401,N_29611);
or UO_782 (O_782,N_29962,N_29999);
or UO_783 (O_783,N_29675,N_29475);
and UO_784 (O_784,N_29978,N_29881);
nor UO_785 (O_785,N_29652,N_29996);
nor UO_786 (O_786,N_29482,N_29592);
or UO_787 (O_787,N_29944,N_29419);
or UO_788 (O_788,N_29964,N_29483);
nand UO_789 (O_789,N_29609,N_29913);
and UO_790 (O_790,N_29764,N_29470);
or UO_791 (O_791,N_29770,N_29447);
and UO_792 (O_792,N_29490,N_29505);
or UO_793 (O_793,N_29939,N_29767);
xnor UO_794 (O_794,N_29492,N_29844);
nand UO_795 (O_795,N_29564,N_29921);
and UO_796 (O_796,N_29837,N_29873);
nor UO_797 (O_797,N_29743,N_29954);
nor UO_798 (O_798,N_29951,N_29521);
nand UO_799 (O_799,N_29547,N_29569);
nand UO_800 (O_800,N_29567,N_29634);
or UO_801 (O_801,N_29760,N_29499);
xor UO_802 (O_802,N_29848,N_29426);
xor UO_803 (O_803,N_29595,N_29509);
or UO_804 (O_804,N_29662,N_29845);
nand UO_805 (O_805,N_29866,N_29905);
nand UO_806 (O_806,N_29668,N_29648);
and UO_807 (O_807,N_29530,N_29429);
nor UO_808 (O_808,N_29798,N_29582);
and UO_809 (O_809,N_29800,N_29630);
nor UO_810 (O_810,N_29829,N_29630);
or UO_811 (O_811,N_29914,N_29654);
nor UO_812 (O_812,N_29935,N_29968);
and UO_813 (O_813,N_29611,N_29513);
and UO_814 (O_814,N_29608,N_29966);
and UO_815 (O_815,N_29528,N_29565);
nor UO_816 (O_816,N_29685,N_29852);
or UO_817 (O_817,N_29559,N_29865);
nor UO_818 (O_818,N_29438,N_29927);
nand UO_819 (O_819,N_29561,N_29853);
and UO_820 (O_820,N_29737,N_29992);
nor UO_821 (O_821,N_29973,N_29443);
xnor UO_822 (O_822,N_29957,N_29905);
nand UO_823 (O_823,N_29618,N_29958);
and UO_824 (O_824,N_29825,N_29664);
nor UO_825 (O_825,N_29522,N_29815);
and UO_826 (O_826,N_29781,N_29681);
and UO_827 (O_827,N_29939,N_29478);
nand UO_828 (O_828,N_29817,N_29629);
or UO_829 (O_829,N_29521,N_29998);
or UO_830 (O_830,N_29494,N_29594);
and UO_831 (O_831,N_29703,N_29594);
and UO_832 (O_832,N_29734,N_29992);
nor UO_833 (O_833,N_29542,N_29941);
or UO_834 (O_834,N_29916,N_29803);
xnor UO_835 (O_835,N_29943,N_29691);
or UO_836 (O_836,N_29544,N_29690);
nand UO_837 (O_837,N_29445,N_29462);
nor UO_838 (O_838,N_29903,N_29827);
and UO_839 (O_839,N_29955,N_29745);
nor UO_840 (O_840,N_29915,N_29779);
or UO_841 (O_841,N_29708,N_29956);
and UO_842 (O_842,N_29799,N_29573);
or UO_843 (O_843,N_29739,N_29527);
or UO_844 (O_844,N_29704,N_29898);
or UO_845 (O_845,N_29719,N_29937);
xnor UO_846 (O_846,N_29464,N_29453);
xor UO_847 (O_847,N_29919,N_29944);
or UO_848 (O_848,N_29576,N_29954);
xnor UO_849 (O_849,N_29735,N_29539);
nand UO_850 (O_850,N_29492,N_29643);
or UO_851 (O_851,N_29573,N_29493);
nor UO_852 (O_852,N_29530,N_29783);
nor UO_853 (O_853,N_29871,N_29540);
nand UO_854 (O_854,N_29755,N_29786);
nor UO_855 (O_855,N_29637,N_29565);
and UO_856 (O_856,N_29979,N_29510);
or UO_857 (O_857,N_29632,N_29454);
or UO_858 (O_858,N_29955,N_29866);
and UO_859 (O_859,N_29760,N_29890);
or UO_860 (O_860,N_29488,N_29625);
xor UO_861 (O_861,N_29782,N_29662);
or UO_862 (O_862,N_29501,N_29841);
nor UO_863 (O_863,N_29640,N_29797);
nand UO_864 (O_864,N_29427,N_29884);
nand UO_865 (O_865,N_29908,N_29859);
and UO_866 (O_866,N_29418,N_29839);
and UO_867 (O_867,N_29912,N_29731);
xor UO_868 (O_868,N_29457,N_29750);
nor UO_869 (O_869,N_29851,N_29688);
nand UO_870 (O_870,N_29552,N_29585);
nand UO_871 (O_871,N_29989,N_29569);
xor UO_872 (O_872,N_29958,N_29474);
nor UO_873 (O_873,N_29476,N_29920);
nor UO_874 (O_874,N_29940,N_29504);
or UO_875 (O_875,N_29858,N_29517);
and UO_876 (O_876,N_29603,N_29993);
nand UO_877 (O_877,N_29915,N_29533);
or UO_878 (O_878,N_29498,N_29549);
nor UO_879 (O_879,N_29435,N_29483);
nor UO_880 (O_880,N_29584,N_29508);
xor UO_881 (O_881,N_29686,N_29691);
nor UO_882 (O_882,N_29420,N_29550);
nor UO_883 (O_883,N_29794,N_29846);
and UO_884 (O_884,N_29828,N_29826);
nor UO_885 (O_885,N_29464,N_29501);
nor UO_886 (O_886,N_29799,N_29425);
nand UO_887 (O_887,N_29695,N_29589);
and UO_888 (O_888,N_29658,N_29766);
and UO_889 (O_889,N_29636,N_29757);
nand UO_890 (O_890,N_29578,N_29429);
nand UO_891 (O_891,N_29535,N_29611);
nor UO_892 (O_892,N_29454,N_29816);
nand UO_893 (O_893,N_29569,N_29608);
or UO_894 (O_894,N_29525,N_29539);
nand UO_895 (O_895,N_29738,N_29807);
nor UO_896 (O_896,N_29746,N_29685);
nand UO_897 (O_897,N_29435,N_29816);
nor UO_898 (O_898,N_29428,N_29752);
and UO_899 (O_899,N_29764,N_29886);
xor UO_900 (O_900,N_29850,N_29843);
or UO_901 (O_901,N_29534,N_29717);
nor UO_902 (O_902,N_29532,N_29976);
nor UO_903 (O_903,N_29823,N_29767);
nand UO_904 (O_904,N_29513,N_29481);
nor UO_905 (O_905,N_29829,N_29561);
nand UO_906 (O_906,N_29695,N_29843);
nand UO_907 (O_907,N_29912,N_29900);
xor UO_908 (O_908,N_29788,N_29659);
and UO_909 (O_909,N_29760,N_29671);
nand UO_910 (O_910,N_29901,N_29656);
and UO_911 (O_911,N_29941,N_29834);
xor UO_912 (O_912,N_29739,N_29755);
or UO_913 (O_913,N_29403,N_29504);
nor UO_914 (O_914,N_29487,N_29915);
nand UO_915 (O_915,N_29728,N_29956);
and UO_916 (O_916,N_29481,N_29883);
and UO_917 (O_917,N_29628,N_29895);
and UO_918 (O_918,N_29788,N_29457);
nor UO_919 (O_919,N_29528,N_29502);
and UO_920 (O_920,N_29442,N_29542);
nor UO_921 (O_921,N_29879,N_29832);
or UO_922 (O_922,N_29966,N_29733);
nand UO_923 (O_923,N_29697,N_29823);
nand UO_924 (O_924,N_29835,N_29882);
nand UO_925 (O_925,N_29723,N_29783);
or UO_926 (O_926,N_29666,N_29807);
and UO_927 (O_927,N_29631,N_29574);
and UO_928 (O_928,N_29880,N_29772);
or UO_929 (O_929,N_29525,N_29719);
and UO_930 (O_930,N_29832,N_29843);
nand UO_931 (O_931,N_29842,N_29548);
nand UO_932 (O_932,N_29845,N_29734);
and UO_933 (O_933,N_29697,N_29753);
and UO_934 (O_934,N_29877,N_29487);
nor UO_935 (O_935,N_29523,N_29704);
and UO_936 (O_936,N_29691,N_29603);
or UO_937 (O_937,N_29930,N_29897);
and UO_938 (O_938,N_29493,N_29467);
and UO_939 (O_939,N_29999,N_29431);
nor UO_940 (O_940,N_29683,N_29895);
and UO_941 (O_941,N_29436,N_29472);
nor UO_942 (O_942,N_29504,N_29802);
or UO_943 (O_943,N_29581,N_29957);
nand UO_944 (O_944,N_29911,N_29997);
or UO_945 (O_945,N_29465,N_29841);
and UO_946 (O_946,N_29963,N_29864);
and UO_947 (O_947,N_29465,N_29484);
or UO_948 (O_948,N_29450,N_29445);
nand UO_949 (O_949,N_29540,N_29748);
nor UO_950 (O_950,N_29600,N_29598);
nor UO_951 (O_951,N_29824,N_29972);
nor UO_952 (O_952,N_29627,N_29616);
or UO_953 (O_953,N_29845,N_29933);
nand UO_954 (O_954,N_29549,N_29611);
or UO_955 (O_955,N_29531,N_29792);
xor UO_956 (O_956,N_29438,N_29549);
or UO_957 (O_957,N_29836,N_29830);
and UO_958 (O_958,N_29689,N_29772);
or UO_959 (O_959,N_29681,N_29498);
or UO_960 (O_960,N_29613,N_29916);
or UO_961 (O_961,N_29658,N_29956);
and UO_962 (O_962,N_29956,N_29642);
and UO_963 (O_963,N_29711,N_29650);
nand UO_964 (O_964,N_29409,N_29949);
nand UO_965 (O_965,N_29945,N_29588);
nor UO_966 (O_966,N_29628,N_29601);
and UO_967 (O_967,N_29847,N_29522);
or UO_968 (O_968,N_29629,N_29432);
and UO_969 (O_969,N_29650,N_29618);
or UO_970 (O_970,N_29910,N_29915);
nand UO_971 (O_971,N_29422,N_29822);
or UO_972 (O_972,N_29989,N_29460);
nor UO_973 (O_973,N_29514,N_29814);
and UO_974 (O_974,N_29719,N_29512);
or UO_975 (O_975,N_29966,N_29762);
and UO_976 (O_976,N_29854,N_29971);
and UO_977 (O_977,N_29546,N_29501);
xor UO_978 (O_978,N_29539,N_29823);
nand UO_979 (O_979,N_29955,N_29681);
nand UO_980 (O_980,N_29920,N_29867);
or UO_981 (O_981,N_29508,N_29784);
and UO_982 (O_982,N_29953,N_29422);
and UO_983 (O_983,N_29978,N_29999);
xor UO_984 (O_984,N_29439,N_29768);
or UO_985 (O_985,N_29541,N_29461);
nand UO_986 (O_986,N_29736,N_29901);
or UO_987 (O_987,N_29913,N_29990);
and UO_988 (O_988,N_29779,N_29873);
and UO_989 (O_989,N_29972,N_29435);
and UO_990 (O_990,N_29787,N_29610);
or UO_991 (O_991,N_29958,N_29793);
and UO_992 (O_992,N_29832,N_29547);
nor UO_993 (O_993,N_29920,N_29403);
nor UO_994 (O_994,N_29574,N_29801);
nor UO_995 (O_995,N_29910,N_29411);
or UO_996 (O_996,N_29452,N_29941);
nor UO_997 (O_997,N_29791,N_29741);
or UO_998 (O_998,N_29720,N_29702);
or UO_999 (O_999,N_29983,N_29588);
nand UO_1000 (O_1000,N_29510,N_29646);
or UO_1001 (O_1001,N_29568,N_29516);
and UO_1002 (O_1002,N_29834,N_29897);
and UO_1003 (O_1003,N_29596,N_29841);
nor UO_1004 (O_1004,N_29640,N_29749);
nor UO_1005 (O_1005,N_29796,N_29627);
nor UO_1006 (O_1006,N_29692,N_29993);
and UO_1007 (O_1007,N_29448,N_29635);
nand UO_1008 (O_1008,N_29731,N_29860);
nor UO_1009 (O_1009,N_29497,N_29899);
or UO_1010 (O_1010,N_29975,N_29472);
or UO_1011 (O_1011,N_29965,N_29801);
xor UO_1012 (O_1012,N_29437,N_29648);
and UO_1013 (O_1013,N_29516,N_29461);
nand UO_1014 (O_1014,N_29943,N_29913);
nand UO_1015 (O_1015,N_29985,N_29528);
and UO_1016 (O_1016,N_29588,N_29957);
or UO_1017 (O_1017,N_29562,N_29794);
nor UO_1018 (O_1018,N_29844,N_29636);
or UO_1019 (O_1019,N_29467,N_29542);
nand UO_1020 (O_1020,N_29826,N_29477);
and UO_1021 (O_1021,N_29442,N_29538);
and UO_1022 (O_1022,N_29833,N_29548);
nand UO_1023 (O_1023,N_29730,N_29451);
xnor UO_1024 (O_1024,N_29664,N_29895);
nand UO_1025 (O_1025,N_29704,N_29809);
or UO_1026 (O_1026,N_29411,N_29742);
and UO_1027 (O_1027,N_29954,N_29430);
xor UO_1028 (O_1028,N_29684,N_29828);
nor UO_1029 (O_1029,N_29960,N_29648);
nor UO_1030 (O_1030,N_29513,N_29689);
or UO_1031 (O_1031,N_29871,N_29985);
or UO_1032 (O_1032,N_29957,N_29801);
nor UO_1033 (O_1033,N_29991,N_29938);
and UO_1034 (O_1034,N_29596,N_29970);
nand UO_1035 (O_1035,N_29916,N_29447);
nand UO_1036 (O_1036,N_29699,N_29861);
nor UO_1037 (O_1037,N_29455,N_29493);
nand UO_1038 (O_1038,N_29886,N_29946);
and UO_1039 (O_1039,N_29615,N_29776);
nand UO_1040 (O_1040,N_29430,N_29986);
nand UO_1041 (O_1041,N_29474,N_29809);
nand UO_1042 (O_1042,N_29909,N_29697);
nor UO_1043 (O_1043,N_29584,N_29889);
nand UO_1044 (O_1044,N_29575,N_29645);
or UO_1045 (O_1045,N_29438,N_29972);
and UO_1046 (O_1046,N_29488,N_29616);
and UO_1047 (O_1047,N_29487,N_29594);
or UO_1048 (O_1048,N_29706,N_29400);
nor UO_1049 (O_1049,N_29699,N_29805);
nor UO_1050 (O_1050,N_29530,N_29845);
and UO_1051 (O_1051,N_29646,N_29639);
nor UO_1052 (O_1052,N_29968,N_29685);
or UO_1053 (O_1053,N_29643,N_29943);
or UO_1054 (O_1054,N_29692,N_29793);
or UO_1055 (O_1055,N_29893,N_29946);
nand UO_1056 (O_1056,N_29559,N_29630);
or UO_1057 (O_1057,N_29918,N_29661);
nor UO_1058 (O_1058,N_29853,N_29682);
or UO_1059 (O_1059,N_29912,N_29876);
or UO_1060 (O_1060,N_29455,N_29538);
or UO_1061 (O_1061,N_29879,N_29476);
and UO_1062 (O_1062,N_29553,N_29798);
nand UO_1063 (O_1063,N_29846,N_29556);
and UO_1064 (O_1064,N_29708,N_29835);
xnor UO_1065 (O_1065,N_29501,N_29612);
or UO_1066 (O_1066,N_29527,N_29753);
or UO_1067 (O_1067,N_29805,N_29865);
or UO_1068 (O_1068,N_29933,N_29770);
nand UO_1069 (O_1069,N_29628,N_29757);
nor UO_1070 (O_1070,N_29671,N_29435);
and UO_1071 (O_1071,N_29601,N_29814);
or UO_1072 (O_1072,N_29479,N_29995);
and UO_1073 (O_1073,N_29534,N_29745);
and UO_1074 (O_1074,N_29893,N_29846);
xnor UO_1075 (O_1075,N_29590,N_29485);
nand UO_1076 (O_1076,N_29541,N_29735);
nand UO_1077 (O_1077,N_29968,N_29721);
or UO_1078 (O_1078,N_29442,N_29816);
nand UO_1079 (O_1079,N_29562,N_29637);
nand UO_1080 (O_1080,N_29631,N_29748);
nor UO_1081 (O_1081,N_29901,N_29869);
nor UO_1082 (O_1082,N_29562,N_29546);
nand UO_1083 (O_1083,N_29734,N_29901);
nor UO_1084 (O_1084,N_29782,N_29909);
and UO_1085 (O_1085,N_29864,N_29446);
nand UO_1086 (O_1086,N_29979,N_29622);
nand UO_1087 (O_1087,N_29524,N_29884);
nand UO_1088 (O_1088,N_29543,N_29438);
and UO_1089 (O_1089,N_29810,N_29743);
nor UO_1090 (O_1090,N_29705,N_29935);
xnor UO_1091 (O_1091,N_29459,N_29427);
xnor UO_1092 (O_1092,N_29735,N_29632);
xnor UO_1093 (O_1093,N_29717,N_29634);
xor UO_1094 (O_1094,N_29947,N_29510);
or UO_1095 (O_1095,N_29978,N_29601);
nor UO_1096 (O_1096,N_29425,N_29892);
or UO_1097 (O_1097,N_29779,N_29816);
nor UO_1098 (O_1098,N_29615,N_29910);
nor UO_1099 (O_1099,N_29936,N_29843);
and UO_1100 (O_1100,N_29756,N_29797);
xnor UO_1101 (O_1101,N_29749,N_29921);
nand UO_1102 (O_1102,N_29968,N_29492);
or UO_1103 (O_1103,N_29677,N_29681);
nand UO_1104 (O_1104,N_29492,N_29453);
and UO_1105 (O_1105,N_29739,N_29953);
xnor UO_1106 (O_1106,N_29735,N_29908);
nor UO_1107 (O_1107,N_29688,N_29433);
nor UO_1108 (O_1108,N_29910,N_29627);
and UO_1109 (O_1109,N_29935,N_29863);
nor UO_1110 (O_1110,N_29966,N_29875);
nor UO_1111 (O_1111,N_29446,N_29809);
nand UO_1112 (O_1112,N_29817,N_29400);
or UO_1113 (O_1113,N_29639,N_29626);
and UO_1114 (O_1114,N_29842,N_29973);
nor UO_1115 (O_1115,N_29906,N_29759);
nand UO_1116 (O_1116,N_29820,N_29402);
nor UO_1117 (O_1117,N_29806,N_29592);
and UO_1118 (O_1118,N_29497,N_29912);
nand UO_1119 (O_1119,N_29484,N_29401);
nor UO_1120 (O_1120,N_29479,N_29488);
nand UO_1121 (O_1121,N_29609,N_29786);
nand UO_1122 (O_1122,N_29751,N_29763);
nand UO_1123 (O_1123,N_29857,N_29785);
or UO_1124 (O_1124,N_29558,N_29767);
xnor UO_1125 (O_1125,N_29449,N_29497);
nor UO_1126 (O_1126,N_29564,N_29926);
and UO_1127 (O_1127,N_29480,N_29548);
and UO_1128 (O_1128,N_29739,N_29972);
xnor UO_1129 (O_1129,N_29900,N_29947);
nor UO_1130 (O_1130,N_29535,N_29822);
xor UO_1131 (O_1131,N_29978,N_29896);
and UO_1132 (O_1132,N_29743,N_29926);
and UO_1133 (O_1133,N_29802,N_29519);
nor UO_1134 (O_1134,N_29779,N_29604);
xnor UO_1135 (O_1135,N_29783,N_29941);
and UO_1136 (O_1136,N_29512,N_29470);
or UO_1137 (O_1137,N_29636,N_29400);
nand UO_1138 (O_1138,N_29874,N_29741);
nand UO_1139 (O_1139,N_29577,N_29423);
nand UO_1140 (O_1140,N_29785,N_29899);
nand UO_1141 (O_1141,N_29480,N_29728);
nor UO_1142 (O_1142,N_29612,N_29998);
and UO_1143 (O_1143,N_29577,N_29918);
and UO_1144 (O_1144,N_29669,N_29613);
nand UO_1145 (O_1145,N_29577,N_29473);
xnor UO_1146 (O_1146,N_29449,N_29824);
nor UO_1147 (O_1147,N_29853,N_29490);
nand UO_1148 (O_1148,N_29651,N_29672);
or UO_1149 (O_1149,N_29852,N_29715);
nand UO_1150 (O_1150,N_29778,N_29983);
nand UO_1151 (O_1151,N_29846,N_29929);
nor UO_1152 (O_1152,N_29688,N_29662);
nor UO_1153 (O_1153,N_29850,N_29652);
nor UO_1154 (O_1154,N_29421,N_29780);
or UO_1155 (O_1155,N_29923,N_29671);
nor UO_1156 (O_1156,N_29630,N_29654);
and UO_1157 (O_1157,N_29948,N_29851);
and UO_1158 (O_1158,N_29909,N_29659);
nor UO_1159 (O_1159,N_29980,N_29809);
and UO_1160 (O_1160,N_29673,N_29573);
or UO_1161 (O_1161,N_29648,N_29724);
or UO_1162 (O_1162,N_29996,N_29683);
nand UO_1163 (O_1163,N_29798,N_29863);
nand UO_1164 (O_1164,N_29614,N_29503);
or UO_1165 (O_1165,N_29775,N_29621);
xnor UO_1166 (O_1166,N_29813,N_29989);
xnor UO_1167 (O_1167,N_29545,N_29634);
xor UO_1168 (O_1168,N_29620,N_29551);
nor UO_1169 (O_1169,N_29693,N_29439);
or UO_1170 (O_1170,N_29741,N_29759);
or UO_1171 (O_1171,N_29502,N_29457);
and UO_1172 (O_1172,N_29946,N_29439);
or UO_1173 (O_1173,N_29741,N_29606);
nand UO_1174 (O_1174,N_29658,N_29870);
nand UO_1175 (O_1175,N_29400,N_29696);
or UO_1176 (O_1176,N_29824,N_29730);
xnor UO_1177 (O_1177,N_29456,N_29761);
and UO_1178 (O_1178,N_29965,N_29808);
and UO_1179 (O_1179,N_29524,N_29880);
nand UO_1180 (O_1180,N_29471,N_29991);
or UO_1181 (O_1181,N_29742,N_29543);
nor UO_1182 (O_1182,N_29569,N_29853);
nand UO_1183 (O_1183,N_29430,N_29514);
nor UO_1184 (O_1184,N_29924,N_29418);
nor UO_1185 (O_1185,N_29669,N_29610);
or UO_1186 (O_1186,N_29918,N_29437);
nor UO_1187 (O_1187,N_29534,N_29898);
nor UO_1188 (O_1188,N_29455,N_29762);
xor UO_1189 (O_1189,N_29630,N_29737);
or UO_1190 (O_1190,N_29980,N_29799);
nand UO_1191 (O_1191,N_29485,N_29596);
xnor UO_1192 (O_1192,N_29712,N_29430);
and UO_1193 (O_1193,N_29842,N_29938);
and UO_1194 (O_1194,N_29872,N_29478);
nor UO_1195 (O_1195,N_29797,N_29574);
and UO_1196 (O_1196,N_29704,N_29481);
xor UO_1197 (O_1197,N_29675,N_29869);
xor UO_1198 (O_1198,N_29509,N_29990);
nor UO_1199 (O_1199,N_29860,N_29440);
or UO_1200 (O_1200,N_29906,N_29640);
or UO_1201 (O_1201,N_29532,N_29626);
nor UO_1202 (O_1202,N_29921,N_29908);
nor UO_1203 (O_1203,N_29688,N_29550);
nand UO_1204 (O_1204,N_29615,N_29420);
nand UO_1205 (O_1205,N_29734,N_29965);
xor UO_1206 (O_1206,N_29412,N_29599);
xor UO_1207 (O_1207,N_29877,N_29567);
and UO_1208 (O_1208,N_29588,N_29523);
nand UO_1209 (O_1209,N_29964,N_29624);
or UO_1210 (O_1210,N_29963,N_29853);
nand UO_1211 (O_1211,N_29938,N_29745);
nor UO_1212 (O_1212,N_29416,N_29505);
nor UO_1213 (O_1213,N_29970,N_29585);
and UO_1214 (O_1214,N_29648,N_29786);
nor UO_1215 (O_1215,N_29861,N_29922);
nor UO_1216 (O_1216,N_29591,N_29914);
xnor UO_1217 (O_1217,N_29781,N_29721);
or UO_1218 (O_1218,N_29478,N_29837);
or UO_1219 (O_1219,N_29879,N_29945);
nor UO_1220 (O_1220,N_29599,N_29529);
or UO_1221 (O_1221,N_29693,N_29524);
nand UO_1222 (O_1222,N_29449,N_29640);
and UO_1223 (O_1223,N_29836,N_29987);
nand UO_1224 (O_1224,N_29816,N_29857);
nor UO_1225 (O_1225,N_29600,N_29501);
nor UO_1226 (O_1226,N_29851,N_29968);
or UO_1227 (O_1227,N_29666,N_29710);
and UO_1228 (O_1228,N_29652,N_29521);
or UO_1229 (O_1229,N_29902,N_29568);
xor UO_1230 (O_1230,N_29996,N_29994);
and UO_1231 (O_1231,N_29980,N_29910);
and UO_1232 (O_1232,N_29945,N_29970);
xnor UO_1233 (O_1233,N_29969,N_29479);
or UO_1234 (O_1234,N_29931,N_29772);
xor UO_1235 (O_1235,N_29907,N_29520);
or UO_1236 (O_1236,N_29697,N_29618);
and UO_1237 (O_1237,N_29871,N_29756);
nor UO_1238 (O_1238,N_29499,N_29840);
or UO_1239 (O_1239,N_29896,N_29946);
nor UO_1240 (O_1240,N_29413,N_29963);
and UO_1241 (O_1241,N_29737,N_29776);
or UO_1242 (O_1242,N_29702,N_29617);
or UO_1243 (O_1243,N_29816,N_29594);
nand UO_1244 (O_1244,N_29910,N_29889);
nand UO_1245 (O_1245,N_29974,N_29932);
nand UO_1246 (O_1246,N_29832,N_29513);
nor UO_1247 (O_1247,N_29617,N_29912);
or UO_1248 (O_1248,N_29974,N_29865);
and UO_1249 (O_1249,N_29879,N_29762);
or UO_1250 (O_1250,N_29483,N_29770);
nor UO_1251 (O_1251,N_29735,N_29769);
or UO_1252 (O_1252,N_29820,N_29811);
and UO_1253 (O_1253,N_29813,N_29742);
and UO_1254 (O_1254,N_29735,N_29422);
and UO_1255 (O_1255,N_29523,N_29473);
nor UO_1256 (O_1256,N_29815,N_29710);
and UO_1257 (O_1257,N_29704,N_29741);
or UO_1258 (O_1258,N_29940,N_29607);
nand UO_1259 (O_1259,N_29637,N_29617);
and UO_1260 (O_1260,N_29604,N_29455);
nor UO_1261 (O_1261,N_29452,N_29914);
nand UO_1262 (O_1262,N_29674,N_29494);
and UO_1263 (O_1263,N_29633,N_29761);
nor UO_1264 (O_1264,N_29895,N_29974);
nor UO_1265 (O_1265,N_29424,N_29676);
and UO_1266 (O_1266,N_29901,N_29727);
nand UO_1267 (O_1267,N_29548,N_29694);
xor UO_1268 (O_1268,N_29946,N_29685);
and UO_1269 (O_1269,N_29960,N_29538);
xor UO_1270 (O_1270,N_29512,N_29959);
and UO_1271 (O_1271,N_29588,N_29423);
nor UO_1272 (O_1272,N_29621,N_29840);
nor UO_1273 (O_1273,N_29962,N_29899);
nand UO_1274 (O_1274,N_29535,N_29492);
and UO_1275 (O_1275,N_29653,N_29650);
nand UO_1276 (O_1276,N_29833,N_29877);
nand UO_1277 (O_1277,N_29687,N_29918);
xnor UO_1278 (O_1278,N_29643,N_29731);
or UO_1279 (O_1279,N_29532,N_29619);
or UO_1280 (O_1280,N_29809,N_29613);
nor UO_1281 (O_1281,N_29721,N_29463);
and UO_1282 (O_1282,N_29542,N_29768);
and UO_1283 (O_1283,N_29981,N_29837);
and UO_1284 (O_1284,N_29476,N_29438);
nand UO_1285 (O_1285,N_29564,N_29718);
nor UO_1286 (O_1286,N_29790,N_29837);
nand UO_1287 (O_1287,N_29422,N_29912);
and UO_1288 (O_1288,N_29757,N_29906);
nor UO_1289 (O_1289,N_29843,N_29818);
and UO_1290 (O_1290,N_29620,N_29779);
and UO_1291 (O_1291,N_29910,N_29730);
nand UO_1292 (O_1292,N_29449,N_29695);
nand UO_1293 (O_1293,N_29949,N_29455);
or UO_1294 (O_1294,N_29573,N_29593);
or UO_1295 (O_1295,N_29686,N_29742);
and UO_1296 (O_1296,N_29785,N_29850);
nor UO_1297 (O_1297,N_29475,N_29814);
or UO_1298 (O_1298,N_29978,N_29633);
nor UO_1299 (O_1299,N_29439,N_29939);
nand UO_1300 (O_1300,N_29911,N_29545);
nand UO_1301 (O_1301,N_29754,N_29580);
or UO_1302 (O_1302,N_29743,N_29953);
and UO_1303 (O_1303,N_29641,N_29784);
nor UO_1304 (O_1304,N_29645,N_29424);
and UO_1305 (O_1305,N_29823,N_29477);
or UO_1306 (O_1306,N_29670,N_29914);
or UO_1307 (O_1307,N_29508,N_29561);
or UO_1308 (O_1308,N_29474,N_29954);
or UO_1309 (O_1309,N_29942,N_29900);
xor UO_1310 (O_1310,N_29473,N_29949);
and UO_1311 (O_1311,N_29896,N_29546);
nand UO_1312 (O_1312,N_29489,N_29771);
and UO_1313 (O_1313,N_29431,N_29446);
xnor UO_1314 (O_1314,N_29596,N_29626);
nor UO_1315 (O_1315,N_29772,N_29996);
nand UO_1316 (O_1316,N_29424,N_29870);
or UO_1317 (O_1317,N_29773,N_29767);
nor UO_1318 (O_1318,N_29433,N_29622);
nand UO_1319 (O_1319,N_29626,N_29795);
and UO_1320 (O_1320,N_29607,N_29725);
or UO_1321 (O_1321,N_29720,N_29979);
nand UO_1322 (O_1322,N_29664,N_29993);
nand UO_1323 (O_1323,N_29635,N_29530);
or UO_1324 (O_1324,N_29473,N_29960);
nor UO_1325 (O_1325,N_29513,N_29529);
or UO_1326 (O_1326,N_29476,N_29470);
nor UO_1327 (O_1327,N_29930,N_29531);
or UO_1328 (O_1328,N_29646,N_29643);
and UO_1329 (O_1329,N_29679,N_29771);
nor UO_1330 (O_1330,N_29708,N_29946);
nor UO_1331 (O_1331,N_29525,N_29958);
nor UO_1332 (O_1332,N_29799,N_29446);
nand UO_1333 (O_1333,N_29487,N_29788);
nand UO_1334 (O_1334,N_29957,N_29984);
or UO_1335 (O_1335,N_29788,N_29646);
and UO_1336 (O_1336,N_29735,N_29832);
and UO_1337 (O_1337,N_29696,N_29916);
or UO_1338 (O_1338,N_29610,N_29467);
nand UO_1339 (O_1339,N_29741,N_29979);
and UO_1340 (O_1340,N_29729,N_29774);
nand UO_1341 (O_1341,N_29581,N_29829);
xor UO_1342 (O_1342,N_29592,N_29755);
nor UO_1343 (O_1343,N_29518,N_29433);
or UO_1344 (O_1344,N_29844,N_29779);
or UO_1345 (O_1345,N_29988,N_29538);
nor UO_1346 (O_1346,N_29894,N_29601);
and UO_1347 (O_1347,N_29533,N_29464);
nand UO_1348 (O_1348,N_29829,N_29413);
or UO_1349 (O_1349,N_29812,N_29486);
nor UO_1350 (O_1350,N_29928,N_29624);
xor UO_1351 (O_1351,N_29996,N_29696);
nand UO_1352 (O_1352,N_29821,N_29460);
nand UO_1353 (O_1353,N_29894,N_29872);
nor UO_1354 (O_1354,N_29706,N_29520);
or UO_1355 (O_1355,N_29472,N_29791);
nor UO_1356 (O_1356,N_29898,N_29969);
or UO_1357 (O_1357,N_29921,N_29617);
and UO_1358 (O_1358,N_29501,N_29732);
or UO_1359 (O_1359,N_29713,N_29463);
and UO_1360 (O_1360,N_29560,N_29556);
nand UO_1361 (O_1361,N_29781,N_29752);
and UO_1362 (O_1362,N_29791,N_29958);
nand UO_1363 (O_1363,N_29621,N_29828);
or UO_1364 (O_1364,N_29610,N_29695);
nor UO_1365 (O_1365,N_29555,N_29754);
or UO_1366 (O_1366,N_29891,N_29763);
or UO_1367 (O_1367,N_29440,N_29660);
nor UO_1368 (O_1368,N_29560,N_29986);
nand UO_1369 (O_1369,N_29485,N_29957);
nor UO_1370 (O_1370,N_29412,N_29697);
nand UO_1371 (O_1371,N_29518,N_29995);
and UO_1372 (O_1372,N_29686,N_29925);
nand UO_1373 (O_1373,N_29922,N_29636);
nand UO_1374 (O_1374,N_29409,N_29891);
nor UO_1375 (O_1375,N_29863,N_29669);
nor UO_1376 (O_1376,N_29888,N_29589);
or UO_1377 (O_1377,N_29841,N_29471);
nor UO_1378 (O_1378,N_29566,N_29957);
xnor UO_1379 (O_1379,N_29541,N_29483);
nand UO_1380 (O_1380,N_29610,N_29824);
and UO_1381 (O_1381,N_29815,N_29963);
and UO_1382 (O_1382,N_29555,N_29614);
xnor UO_1383 (O_1383,N_29477,N_29619);
or UO_1384 (O_1384,N_29817,N_29489);
or UO_1385 (O_1385,N_29680,N_29411);
and UO_1386 (O_1386,N_29705,N_29792);
and UO_1387 (O_1387,N_29494,N_29926);
and UO_1388 (O_1388,N_29539,N_29980);
xor UO_1389 (O_1389,N_29824,N_29650);
xor UO_1390 (O_1390,N_29878,N_29856);
or UO_1391 (O_1391,N_29779,N_29976);
and UO_1392 (O_1392,N_29931,N_29921);
or UO_1393 (O_1393,N_29683,N_29402);
nor UO_1394 (O_1394,N_29497,N_29583);
nand UO_1395 (O_1395,N_29532,N_29628);
nand UO_1396 (O_1396,N_29483,N_29911);
nand UO_1397 (O_1397,N_29447,N_29454);
and UO_1398 (O_1398,N_29975,N_29567);
nand UO_1399 (O_1399,N_29708,N_29536);
and UO_1400 (O_1400,N_29932,N_29701);
or UO_1401 (O_1401,N_29615,N_29820);
xor UO_1402 (O_1402,N_29521,N_29640);
and UO_1403 (O_1403,N_29994,N_29792);
and UO_1404 (O_1404,N_29897,N_29805);
and UO_1405 (O_1405,N_29731,N_29734);
and UO_1406 (O_1406,N_29967,N_29581);
nand UO_1407 (O_1407,N_29480,N_29490);
or UO_1408 (O_1408,N_29982,N_29768);
xnor UO_1409 (O_1409,N_29625,N_29596);
nand UO_1410 (O_1410,N_29581,N_29457);
nand UO_1411 (O_1411,N_29853,N_29517);
xor UO_1412 (O_1412,N_29495,N_29537);
and UO_1413 (O_1413,N_29502,N_29722);
xnor UO_1414 (O_1414,N_29893,N_29947);
nand UO_1415 (O_1415,N_29613,N_29792);
nand UO_1416 (O_1416,N_29862,N_29572);
nor UO_1417 (O_1417,N_29900,N_29637);
nand UO_1418 (O_1418,N_29579,N_29954);
nor UO_1419 (O_1419,N_29927,N_29811);
or UO_1420 (O_1420,N_29801,N_29684);
nand UO_1421 (O_1421,N_29877,N_29492);
nand UO_1422 (O_1422,N_29451,N_29876);
nand UO_1423 (O_1423,N_29655,N_29552);
and UO_1424 (O_1424,N_29538,N_29830);
nor UO_1425 (O_1425,N_29960,N_29748);
or UO_1426 (O_1426,N_29605,N_29443);
nor UO_1427 (O_1427,N_29907,N_29496);
or UO_1428 (O_1428,N_29849,N_29941);
and UO_1429 (O_1429,N_29605,N_29951);
or UO_1430 (O_1430,N_29541,N_29584);
and UO_1431 (O_1431,N_29535,N_29485);
or UO_1432 (O_1432,N_29519,N_29719);
and UO_1433 (O_1433,N_29919,N_29996);
xnor UO_1434 (O_1434,N_29888,N_29934);
nor UO_1435 (O_1435,N_29532,N_29499);
and UO_1436 (O_1436,N_29534,N_29434);
xor UO_1437 (O_1437,N_29810,N_29778);
nor UO_1438 (O_1438,N_29905,N_29737);
nor UO_1439 (O_1439,N_29959,N_29815);
nand UO_1440 (O_1440,N_29756,N_29980);
nor UO_1441 (O_1441,N_29739,N_29763);
nor UO_1442 (O_1442,N_29827,N_29474);
nand UO_1443 (O_1443,N_29455,N_29872);
or UO_1444 (O_1444,N_29815,N_29977);
nand UO_1445 (O_1445,N_29535,N_29724);
nand UO_1446 (O_1446,N_29556,N_29729);
or UO_1447 (O_1447,N_29464,N_29784);
nand UO_1448 (O_1448,N_29999,N_29970);
nor UO_1449 (O_1449,N_29632,N_29519);
nand UO_1450 (O_1450,N_29417,N_29519);
nand UO_1451 (O_1451,N_29500,N_29457);
nor UO_1452 (O_1452,N_29900,N_29801);
nand UO_1453 (O_1453,N_29726,N_29509);
and UO_1454 (O_1454,N_29766,N_29863);
or UO_1455 (O_1455,N_29510,N_29799);
xor UO_1456 (O_1456,N_29958,N_29686);
and UO_1457 (O_1457,N_29899,N_29848);
nand UO_1458 (O_1458,N_29481,N_29417);
xnor UO_1459 (O_1459,N_29738,N_29850);
and UO_1460 (O_1460,N_29808,N_29708);
nand UO_1461 (O_1461,N_29913,N_29790);
nand UO_1462 (O_1462,N_29421,N_29763);
nor UO_1463 (O_1463,N_29879,N_29925);
nand UO_1464 (O_1464,N_29778,N_29421);
and UO_1465 (O_1465,N_29537,N_29610);
and UO_1466 (O_1466,N_29453,N_29549);
or UO_1467 (O_1467,N_29865,N_29534);
and UO_1468 (O_1468,N_29906,N_29775);
nor UO_1469 (O_1469,N_29460,N_29714);
or UO_1470 (O_1470,N_29663,N_29790);
nand UO_1471 (O_1471,N_29853,N_29440);
and UO_1472 (O_1472,N_29431,N_29591);
nand UO_1473 (O_1473,N_29767,N_29664);
and UO_1474 (O_1474,N_29845,N_29902);
nand UO_1475 (O_1475,N_29492,N_29974);
nand UO_1476 (O_1476,N_29936,N_29628);
xor UO_1477 (O_1477,N_29499,N_29818);
nand UO_1478 (O_1478,N_29726,N_29675);
and UO_1479 (O_1479,N_29761,N_29765);
nor UO_1480 (O_1480,N_29565,N_29464);
nand UO_1481 (O_1481,N_29833,N_29462);
or UO_1482 (O_1482,N_29790,N_29735);
and UO_1483 (O_1483,N_29419,N_29867);
nor UO_1484 (O_1484,N_29449,N_29486);
and UO_1485 (O_1485,N_29779,N_29505);
or UO_1486 (O_1486,N_29578,N_29738);
xor UO_1487 (O_1487,N_29624,N_29644);
nor UO_1488 (O_1488,N_29931,N_29605);
or UO_1489 (O_1489,N_29723,N_29414);
nor UO_1490 (O_1490,N_29464,N_29539);
nor UO_1491 (O_1491,N_29915,N_29770);
nor UO_1492 (O_1492,N_29699,N_29617);
nand UO_1493 (O_1493,N_29501,N_29453);
xnor UO_1494 (O_1494,N_29676,N_29545);
nand UO_1495 (O_1495,N_29811,N_29685);
nand UO_1496 (O_1496,N_29410,N_29404);
or UO_1497 (O_1497,N_29560,N_29856);
nand UO_1498 (O_1498,N_29483,N_29742);
and UO_1499 (O_1499,N_29879,N_29912);
or UO_1500 (O_1500,N_29435,N_29678);
nor UO_1501 (O_1501,N_29407,N_29854);
nand UO_1502 (O_1502,N_29698,N_29879);
or UO_1503 (O_1503,N_29436,N_29985);
nand UO_1504 (O_1504,N_29786,N_29863);
or UO_1505 (O_1505,N_29822,N_29883);
nor UO_1506 (O_1506,N_29854,N_29793);
xnor UO_1507 (O_1507,N_29525,N_29888);
or UO_1508 (O_1508,N_29891,N_29978);
xor UO_1509 (O_1509,N_29453,N_29965);
and UO_1510 (O_1510,N_29793,N_29446);
and UO_1511 (O_1511,N_29452,N_29711);
nor UO_1512 (O_1512,N_29850,N_29599);
and UO_1513 (O_1513,N_29914,N_29933);
and UO_1514 (O_1514,N_29548,N_29709);
and UO_1515 (O_1515,N_29736,N_29407);
and UO_1516 (O_1516,N_29677,N_29534);
and UO_1517 (O_1517,N_29419,N_29514);
or UO_1518 (O_1518,N_29715,N_29935);
nand UO_1519 (O_1519,N_29974,N_29630);
nand UO_1520 (O_1520,N_29888,N_29538);
nand UO_1521 (O_1521,N_29788,N_29996);
nor UO_1522 (O_1522,N_29577,N_29791);
and UO_1523 (O_1523,N_29809,N_29789);
nand UO_1524 (O_1524,N_29888,N_29565);
or UO_1525 (O_1525,N_29736,N_29965);
and UO_1526 (O_1526,N_29989,N_29750);
nor UO_1527 (O_1527,N_29671,N_29900);
nand UO_1528 (O_1528,N_29761,N_29987);
and UO_1529 (O_1529,N_29434,N_29795);
nor UO_1530 (O_1530,N_29745,N_29625);
nand UO_1531 (O_1531,N_29514,N_29774);
nor UO_1532 (O_1532,N_29590,N_29801);
nor UO_1533 (O_1533,N_29714,N_29706);
nand UO_1534 (O_1534,N_29411,N_29459);
or UO_1535 (O_1535,N_29687,N_29468);
or UO_1536 (O_1536,N_29659,N_29854);
or UO_1537 (O_1537,N_29542,N_29446);
nand UO_1538 (O_1538,N_29566,N_29553);
or UO_1539 (O_1539,N_29917,N_29652);
or UO_1540 (O_1540,N_29414,N_29936);
or UO_1541 (O_1541,N_29612,N_29984);
xnor UO_1542 (O_1542,N_29868,N_29605);
xor UO_1543 (O_1543,N_29701,N_29677);
nor UO_1544 (O_1544,N_29573,N_29678);
nand UO_1545 (O_1545,N_29834,N_29954);
nand UO_1546 (O_1546,N_29919,N_29841);
nand UO_1547 (O_1547,N_29906,N_29915);
nand UO_1548 (O_1548,N_29614,N_29717);
or UO_1549 (O_1549,N_29630,N_29626);
and UO_1550 (O_1550,N_29603,N_29943);
and UO_1551 (O_1551,N_29580,N_29910);
or UO_1552 (O_1552,N_29764,N_29610);
xnor UO_1553 (O_1553,N_29627,N_29655);
nor UO_1554 (O_1554,N_29957,N_29436);
nor UO_1555 (O_1555,N_29985,N_29734);
xor UO_1556 (O_1556,N_29513,N_29969);
nor UO_1557 (O_1557,N_29810,N_29422);
nor UO_1558 (O_1558,N_29964,N_29908);
and UO_1559 (O_1559,N_29486,N_29445);
and UO_1560 (O_1560,N_29417,N_29617);
nand UO_1561 (O_1561,N_29820,N_29756);
nand UO_1562 (O_1562,N_29612,N_29761);
and UO_1563 (O_1563,N_29959,N_29926);
nor UO_1564 (O_1564,N_29470,N_29748);
and UO_1565 (O_1565,N_29679,N_29559);
or UO_1566 (O_1566,N_29650,N_29837);
nand UO_1567 (O_1567,N_29556,N_29479);
nand UO_1568 (O_1568,N_29756,N_29789);
and UO_1569 (O_1569,N_29695,N_29694);
nand UO_1570 (O_1570,N_29401,N_29672);
and UO_1571 (O_1571,N_29872,N_29752);
nand UO_1572 (O_1572,N_29762,N_29899);
nor UO_1573 (O_1573,N_29988,N_29627);
nand UO_1574 (O_1574,N_29619,N_29681);
and UO_1575 (O_1575,N_29551,N_29791);
nor UO_1576 (O_1576,N_29916,N_29530);
xor UO_1577 (O_1577,N_29913,N_29593);
and UO_1578 (O_1578,N_29841,N_29929);
and UO_1579 (O_1579,N_29490,N_29544);
nand UO_1580 (O_1580,N_29945,N_29779);
and UO_1581 (O_1581,N_29593,N_29874);
and UO_1582 (O_1582,N_29620,N_29452);
nand UO_1583 (O_1583,N_29952,N_29663);
or UO_1584 (O_1584,N_29781,N_29427);
nand UO_1585 (O_1585,N_29924,N_29450);
or UO_1586 (O_1586,N_29728,N_29513);
and UO_1587 (O_1587,N_29601,N_29942);
and UO_1588 (O_1588,N_29761,N_29835);
or UO_1589 (O_1589,N_29432,N_29671);
and UO_1590 (O_1590,N_29930,N_29566);
nor UO_1591 (O_1591,N_29918,N_29948);
nor UO_1592 (O_1592,N_29479,N_29539);
or UO_1593 (O_1593,N_29450,N_29827);
and UO_1594 (O_1594,N_29465,N_29495);
nand UO_1595 (O_1595,N_29929,N_29773);
and UO_1596 (O_1596,N_29422,N_29545);
nand UO_1597 (O_1597,N_29699,N_29882);
nor UO_1598 (O_1598,N_29697,N_29628);
or UO_1599 (O_1599,N_29593,N_29403);
xnor UO_1600 (O_1600,N_29706,N_29565);
xor UO_1601 (O_1601,N_29653,N_29770);
nand UO_1602 (O_1602,N_29575,N_29669);
or UO_1603 (O_1603,N_29746,N_29483);
nand UO_1604 (O_1604,N_29658,N_29911);
nor UO_1605 (O_1605,N_29473,N_29794);
nor UO_1606 (O_1606,N_29583,N_29921);
nand UO_1607 (O_1607,N_29705,N_29965);
nand UO_1608 (O_1608,N_29893,N_29737);
nor UO_1609 (O_1609,N_29655,N_29412);
or UO_1610 (O_1610,N_29425,N_29992);
nand UO_1611 (O_1611,N_29645,N_29526);
or UO_1612 (O_1612,N_29971,N_29559);
nand UO_1613 (O_1613,N_29977,N_29451);
and UO_1614 (O_1614,N_29973,N_29847);
xor UO_1615 (O_1615,N_29907,N_29615);
xor UO_1616 (O_1616,N_29634,N_29790);
or UO_1617 (O_1617,N_29564,N_29413);
or UO_1618 (O_1618,N_29548,N_29938);
xnor UO_1619 (O_1619,N_29712,N_29406);
and UO_1620 (O_1620,N_29686,N_29635);
or UO_1621 (O_1621,N_29419,N_29791);
nor UO_1622 (O_1622,N_29795,N_29412);
nand UO_1623 (O_1623,N_29602,N_29847);
xnor UO_1624 (O_1624,N_29667,N_29425);
nand UO_1625 (O_1625,N_29521,N_29878);
nor UO_1626 (O_1626,N_29457,N_29792);
nand UO_1627 (O_1627,N_29558,N_29746);
nor UO_1628 (O_1628,N_29953,N_29960);
and UO_1629 (O_1629,N_29722,N_29560);
nor UO_1630 (O_1630,N_29721,N_29718);
or UO_1631 (O_1631,N_29815,N_29713);
and UO_1632 (O_1632,N_29505,N_29889);
or UO_1633 (O_1633,N_29561,N_29982);
xnor UO_1634 (O_1634,N_29596,N_29713);
nand UO_1635 (O_1635,N_29548,N_29773);
nor UO_1636 (O_1636,N_29458,N_29716);
and UO_1637 (O_1637,N_29866,N_29774);
nand UO_1638 (O_1638,N_29432,N_29638);
nor UO_1639 (O_1639,N_29471,N_29642);
nor UO_1640 (O_1640,N_29803,N_29411);
or UO_1641 (O_1641,N_29639,N_29871);
and UO_1642 (O_1642,N_29858,N_29906);
or UO_1643 (O_1643,N_29745,N_29905);
and UO_1644 (O_1644,N_29747,N_29610);
or UO_1645 (O_1645,N_29605,N_29900);
and UO_1646 (O_1646,N_29511,N_29706);
nand UO_1647 (O_1647,N_29836,N_29774);
nand UO_1648 (O_1648,N_29570,N_29416);
nand UO_1649 (O_1649,N_29891,N_29717);
and UO_1650 (O_1650,N_29611,N_29603);
and UO_1651 (O_1651,N_29490,N_29708);
xnor UO_1652 (O_1652,N_29822,N_29996);
and UO_1653 (O_1653,N_29770,N_29949);
and UO_1654 (O_1654,N_29900,N_29782);
and UO_1655 (O_1655,N_29932,N_29929);
and UO_1656 (O_1656,N_29949,N_29508);
and UO_1657 (O_1657,N_29548,N_29519);
nor UO_1658 (O_1658,N_29904,N_29987);
nor UO_1659 (O_1659,N_29509,N_29807);
and UO_1660 (O_1660,N_29774,N_29946);
nand UO_1661 (O_1661,N_29522,N_29534);
nand UO_1662 (O_1662,N_29856,N_29773);
and UO_1663 (O_1663,N_29415,N_29936);
nor UO_1664 (O_1664,N_29468,N_29940);
xnor UO_1665 (O_1665,N_29619,N_29778);
nand UO_1666 (O_1666,N_29640,N_29756);
xnor UO_1667 (O_1667,N_29926,N_29821);
nand UO_1668 (O_1668,N_29870,N_29523);
nand UO_1669 (O_1669,N_29983,N_29802);
and UO_1670 (O_1670,N_29910,N_29505);
or UO_1671 (O_1671,N_29941,N_29576);
or UO_1672 (O_1672,N_29466,N_29404);
nor UO_1673 (O_1673,N_29871,N_29768);
nor UO_1674 (O_1674,N_29586,N_29796);
nor UO_1675 (O_1675,N_29798,N_29416);
nor UO_1676 (O_1676,N_29750,N_29449);
or UO_1677 (O_1677,N_29440,N_29496);
nor UO_1678 (O_1678,N_29871,N_29609);
nand UO_1679 (O_1679,N_29698,N_29846);
nor UO_1680 (O_1680,N_29486,N_29476);
nand UO_1681 (O_1681,N_29760,N_29616);
and UO_1682 (O_1682,N_29730,N_29430);
nor UO_1683 (O_1683,N_29763,N_29407);
or UO_1684 (O_1684,N_29703,N_29547);
xnor UO_1685 (O_1685,N_29903,N_29851);
and UO_1686 (O_1686,N_29852,N_29742);
and UO_1687 (O_1687,N_29815,N_29472);
nor UO_1688 (O_1688,N_29483,N_29722);
and UO_1689 (O_1689,N_29429,N_29988);
nand UO_1690 (O_1690,N_29865,N_29928);
nor UO_1691 (O_1691,N_29684,N_29820);
xor UO_1692 (O_1692,N_29549,N_29677);
and UO_1693 (O_1693,N_29430,N_29516);
nor UO_1694 (O_1694,N_29667,N_29411);
nor UO_1695 (O_1695,N_29730,N_29464);
and UO_1696 (O_1696,N_29867,N_29645);
or UO_1697 (O_1697,N_29675,N_29819);
nor UO_1698 (O_1698,N_29851,N_29879);
xnor UO_1699 (O_1699,N_29478,N_29410);
and UO_1700 (O_1700,N_29668,N_29833);
and UO_1701 (O_1701,N_29571,N_29718);
nor UO_1702 (O_1702,N_29680,N_29688);
and UO_1703 (O_1703,N_29633,N_29796);
nor UO_1704 (O_1704,N_29495,N_29471);
or UO_1705 (O_1705,N_29863,N_29744);
nand UO_1706 (O_1706,N_29646,N_29417);
xnor UO_1707 (O_1707,N_29521,N_29989);
and UO_1708 (O_1708,N_29547,N_29984);
xor UO_1709 (O_1709,N_29412,N_29659);
nand UO_1710 (O_1710,N_29792,N_29452);
nand UO_1711 (O_1711,N_29586,N_29564);
and UO_1712 (O_1712,N_29991,N_29981);
xnor UO_1713 (O_1713,N_29506,N_29675);
nor UO_1714 (O_1714,N_29525,N_29605);
nor UO_1715 (O_1715,N_29810,N_29729);
or UO_1716 (O_1716,N_29459,N_29960);
nor UO_1717 (O_1717,N_29789,N_29729);
nor UO_1718 (O_1718,N_29415,N_29856);
nor UO_1719 (O_1719,N_29411,N_29854);
and UO_1720 (O_1720,N_29703,N_29836);
or UO_1721 (O_1721,N_29908,N_29747);
and UO_1722 (O_1722,N_29615,N_29869);
xor UO_1723 (O_1723,N_29832,N_29992);
nor UO_1724 (O_1724,N_29796,N_29421);
and UO_1725 (O_1725,N_29867,N_29850);
nand UO_1726 (O_1726,N_29691,N_29795);
nand UO_1727 (O_1727,N_29989,N_29967);
or UO_1728 (O_1728,N_29722,N_29503);
or UO_1729 (O_1729,N_29682,N_29420);
and UO_1730 (O_1730,N_29469,N_29985);
or UO_1731 (O_1731,N_29708,N_29970);
nand UO_1732 (O_1732,N_29617,N_29648);
and UO_1733 (O_1733,N_29440,N_29914);
and UO_1734 (O_1734,N_29997,N_29458);
xnor UO_1735 (O_1735,N_29743,N_29518);
nand UO_1736 (O_1736,N_29428,N_29821);
nor UO_1737 (O_1737,N_29770,N_29434);
and UO_1738 (O_1738,N_29988,N_29921);
nor UO_1739 (O_1739,N_29917,N_29882);
or UO_1740 (O_1740,N_29535,N_29700);
or UO_1741 (O_1741,N_29917,N_29638);
nand UO_1742 (O_1742,N_29623,N_29712);
nor UO_1743 (O_1743,N_29989,N_29783);
nor UO_1744 (O_1744,N_29646,N_29853);
and UO_1745 (O_1745,N_29931,N_29523);
or UO_1746 (O_1746,N_29939,N_29604);
nor UO_1747 (O_1747,N_29416,N_29892);
nand UO_1748 (O_1748,N_29671,N_29546);
and UO_1749 (O_1749,N_29706,N_29923);
xnor UO_1750 (O_1750,N_29498,N_29544);
nand UO_1751 (O_1751,N_29774,N_29701);
xnor UO_1752 (O_1752,N_29724,N_29997);
nand UO_1753 (O_1753,N_29705,N_29656);
xor UO_1754 (O_1754,N_29993,N_29956);
nand UO_1755 (O_1755,N_29798,N_29956);
xnor UO_1756 (O_1756,N_29657,N_29695);
nand UO_1757 (O_1757,N_29910,N_29897);
nand UO_1758 (O_1758,N_29914,N_29680);
nor UO_1759 (O_1759,N_29863,N_29572);
nor UO_1760 (O_1760,N_29739,N_29800);
nand UO_1761 (O_1761,N_29947,N_29413);
nor UO_1762 (O_1762,N_29599,N_29792);
xor UO_1763 (O_1763,N_29884,N_29889);
or UO_1764 (O_1764,N_29739,N_29984);
nand UO_1765 (O_1765,N_29500,N_29909);
nand UO_1766 (O_1766,N_29795,N_29950);
nor UO_1767 (O_1767,N_29901,N_29440);
nor UO_1768 (O_1768,N_29475,N_29792);
nand UO_1769 (O_1769,N_29924,N_29566);
nand UO_1770 (O_1770,N_29758,N_29566);
and UO_1771 (O_1771,N_29445,N_29809);
xor UO_1772 (O_1772,N_29997,N_29993);
nor UO_1773 (O_1773,N_29405,N_29864);
nor UO_1774 (O_1774,N_29713,N_29877);
or UO_1775 (O_1775,N_29854,N_29870);
or UO_1776 (O_1776,N_29612,N_29823);
or UO_1777 (O_1777,N_29466,N_29468);
nand UO_1778 (O_1778,N_29924,N_29637);
or UO_1779 (O_1779,N_29862,N_29978);
and UO_1780 (O_1780,N_29500,N_29420);
nand UO_1781 (O_1781,N_29585,N_29874);
or UO_1782 (O_1782,N_29806,N_29911);
or UO_1783 (O_1783,N_29657,N_29931);
nor UO_1784 (O_1784,N_29485,N_29892);
nor UO_1785 (O_1785,N_29496,N_29800);
and UO_1786 (O_1786,N_29700,N_29954);
xnor UO_1787 (O_1787,N_29500,N_29967);
nand UO_1788 (O_1788,N_29910,N_29843);
xor UO_1789 (O_1789,N_29657,N_29782);
or UO_1790 (O_1790,N_29683,N_29805);
nor UO_1791 (O_1791,N_29724,N_29680);
nor UO_1792 (O_1792,N_29982,N_29916);
and UO_1793 (O_1793,N_29822,N_29913);
nand UO_1794 (O_1794,N_29940,N_29548);
and UO_1795 (O_1795,N_29808,N_29909);
nor UO_1796 (O_1796,N_29812,N_29575);
nor UO_1797 (O_1797,N_29927,N_29489);
nor UO_1798 (O_1798,N_29813,N_29446);
and UO_1799 (O_1799,N_29860,N_29810);
and UO_1800 (O_1800,N_29489,N_29765);
and UO_1801 (O_1801,N_29625,N_29851);
nand UO_1802 (O_1802,N_29458,N_29948);
or UO_1803 (O_1803,N_29737,N_29527);
nand UO_1804 (O_1804,N_29513,N_29945);
and UO_1805 (O_1805,N_29558,N_29910);
and UO_1806 (O_1806,N_29800,N_29596);
xnor UO_1807 (O_1807,N_29887,N_29618);
nand UO_1808 (O_1808,N_29623,N_29855);
xnor UO_1809 (O_1809,N_29846,N_29510);
and UO_1810 (O_1810,N_29955,N_29511);
or UO_1811 (O_1811,N_29866,N_29482);
or UO_1812 (O_1812,N_29543,N_29755);
and UO_1813 (O_1813,N_29558,N_29846);
xnor UO_1814 (O_1814,N_29643,N_29525);
nor UO_1815 (O_1815,N_29983,N_29712);
nand UO_1816 (O_1816,N_29647,N_29627);
nor UO_1817 (O_1817,N_29709,N_29474);
nand UO_1818 (O_1818,N_29964,N_29981);
nand UO_1819 (O_1819,N_29971,N_29487);
and UO_1820 (O_1820,N_29561,N_29846);
nand UO_1821 (O_1821,N_29904,N_29769);
or UO_1822 (O_1822,N_29602,N_29927);
and UO_1823 (O_1823,N_29667,N_29896);
nor UO_1824 (O_1824,N_29950,N_29870);
nor UO_1825 (O_1825,N_29444,N_29740);
nor UO_1826 (O_1826,N_29568,N_29612);
or UO_1827 (O_1827,N_29840,N_29837);
and UO_1828 (O_1828,N_29885,N_29680);
nand UO_1829 (O_1829,N_29623,N_29716);
or UO_1830 (O_1830,N_29696,N_29720);
and UO_1831 (O_1831,N_29827,N_29455);
or UO_1832 (O_1832,N_29665,N_29756);
and UO_1833 (O_1833,N_29530,N_29588);
nor UO_1834 (O_1834,N_29660,N_29681);
and UO_1835 (O_1835,N_29655,N_29740);
nand UO_1836 (O_1836,N_29749,N_29488);
xor UO_1837 (O_1837,N_29993,N_29578);
xor UO_1838 (O_1838,N_29631,N_29767);
nand UO_1839 (O_1839,N_29715,N_29756);
nor UO_1840 (O_1840,N_29660,N_29884);
and UO_1841 (O_1841,N_29447,N_29675);
or UO_1842 (O_1842,N_29879,N_29466);
xnor UO_1843 (O_1843,N_29851,N_29712);
xor UO_1844 (O_1844,N_29958,N_29546);
or UO_1845 (O_1845,N_29585,N_29519);
or UO_1846 (O_1846,N_29438,N_29401);
and UO_1847 (O_1847,N_29667,N_29751);
nor UO_1848 (O_1848,N_29513,N_29801);
nor UO_1849 (O_1849,N_29666,N_29820);
nor UO_1850 (O_1850,N_29435,N_29446);
and UO_1851 (O_1851,N_29553,N_29729);
or UO_1852 (O_1852,N_29757,N_29864);
xnor UO_1853 (O_1853,N_29465,N_29787);
or UO_1854 (O_1854,N_29882,N_29887);
nand UO_1855 (O_1855,N_29873,N_29679);
and UO_1856 (O_1856,N_29942,N_29726);
nand UO_1857 (O_1857,N_29491,N_29861);
or UO_1858 (O_1858,N_29829,N_29972);
nand UO_1859 (O_1859,N_29457,N_29910);
xor UO_1860 (O_1860,N_29561,N_29809);
and UO_1861 (O_1861,N_29583,N_29526);
nor UO_1862 (O_1862,N_29731,N_29847);
nor UO_1863 (O_1863,N_29829,N_29641);
and UO_1864 (O_1864,N_29961,N_29495);
xnor UO_1865 (O_1865,N_29435,N_29445);
nand UO_1866 (O_1866,N_29977,N_29637);
nand UO_1867 (O_1867,N_29690,N_29719);
nand UO_1868 (O_1868,N_29822,N_29946);
xnor UO_1869 (O_1869,N_29863,N_29938);
nand UO_1870 (O_1870,N_29584,N_29795);
or UO_1871 (O_1871,N_29521,N_29802);
nor UO_1872 (O_1872,N_29969,N_29657);
or UO_1873 (O_1873,N_29914,N_29493);
and UO_1874 (O_1874,N_29875,N_29672);
or UO_1875 (O_1875,N_29808,N_29913);
nand UO_1876 (O_1876,N_29535,N_29409);
or UO_1877 (O_1877,N_29616,N_29596);
or UO_1878 (O_1878,N_29489,N_29720);
nor UO_1879 (O_1879,N_29615,N_29890);
or UO_1880 (O_1880,N_29987,N_29591);
and UO_1881 (O_1881,N_29736,N_29552);
nor UO_1882 (O_1882,N_29804,N_29979);
nor UO_1883 (O_1883,N_29415,N_29732);
nand UO_1884 (O_1884,N_29642,N_29703);
or UO_1885 (O_1885,N_29694,N_29732);
nand UO_1886 (O_1886,N_29442,N_29418);
or UO_1887 (O_1887,N_29628,N_29439);
or UO_1888 (O_1888,N_29574,N_29924);
nand UO_1889 (O_1889,N_29640,N_29900);
nand UO_1890 (O_1890,N_29689,N_29956);
nor UO_1891 (O_1891,N_29547,N_29546);
and UO_1892 (O_1892,N_29504,N_29552);
xnor UO_1893 (O_1893,N_29844,N_29968);
nor UO_1894 (O_1894,N_29598,N_29534);
nand UO_1895 (O_1895,N_29567,N_29521);
and UO_1896 (O_1896,N_29511,N_29957);
nand UO_1897 (O_1897,N_29658,N_29581);
nand UO_1898 (O_1898,N_29894,N_29693);
xor UO_1899 (O_1899,N_29955,N_29642);
nand UO_1900 (O_1900,N_29732,N_29741);
and UO_1901 (O_1901,N_29406,N_29716);
nand UO_1902 (O_1902,N_29855,N_29786);
or UO_1903 (O_1903,N_29549,N_29758);
nand UO_1904 (O_1904,N_29508,N_29506);
xnor UO_1905 (O_1905,N_29609,N_29608);
nor UO_1906 (O_1906,N_29907,N_29458);
or UO_1907 (O_1907,N_29710,N_29718);
or UO_1908 (O_1908,N_29485,N_29865);
and UO_1909 (O_1909,N_29848,N_29996);
nand UO_1910 (O_1910,N_29717,N_29528);
nor UO_1911 (O_1911,N_29682,N_29948);
or UO_1912 (O_1912,N_29563,N_29494);
or UO_1913 (O_1913,N_29890,N_29556);
nand UO_1914 (O_1914,N_29454,N_29817);
and UO_1915 (O_1915,N_29658,N_29915);
or UO_1916 (O_1916,N_29452,N_29775);
nand UO_1917 (O_1917,N_29798,N_29457);
and UO_1918 (O_1918,N_29485,N_29913);
and UO_1919 (O_1919,N_29417,N_29444);
nand UO_1920 (O_1920,N_29751,N_29915);
xnor UO_1921 (O_1921,N_29802,N_29768);
and UO_1922 (O_1922,N_29506,N_29912);
nand UO_1923 (O_1923,N_29411,N_29767);
and UO_1924 (O_1924,N_29934,N_29698);
or UO_1925 (O_1925,N_29685,N_29622);
nor UO_1926 (O_1926,N_29574,N_29648);
or UO_1927 (O_1927,N_29515,N_29721);
xnor UO_1928 (O_1928,N_29555,N_29468);
or UO_1929 (O_1929,N_29719,N_29503);
or UO_1930 (O_1930,N_29723,N_29602);
and UO_1931 (O_1931,N_29573,N_29629);
and UO_1932 (O_1932,N_29509,N_29814);
and UO_1933 (O_1933,N_29412,N_29813);
and UO_1934 (O_1934,N_29895,N_29715);
nand UO_1935 (O_1935,N_29896,N_29965);
and UO_1936 (O_1936,N_29980,N_29693);
nand UO_1937 (O_1937,N_29485,N_29757);
nand UO_1938 (O_1938,N_29860,N_29982);
nand UO_1939 (O_1939,N_29765,N_29837);
nor UO_1940 (O_1940,N_29625,N_29516);
and UO_1941 (O_1941,N_29727,N_29579);
or UO_1942 (O_1942,N_29405,N_29565);
nor UO_1943 (O_1943,N_29416,N_29561);
or UO_1944 (O_1944,N_29934,N_29981);
nor UO_1945 (O_1945,N_29594,N_29537);
and UO_1946 (O_1946,N_29554,N_29903);
nor UO_1947 (O_1947,N_29931,N_29795);
and UO_1948 (O_1948,N_29930,N_29886);
nand UO_1949 (O_1949,N_29681,N_29939);
nand UO_1950 (O_1950,N_29971,N_29810);
or UO_1951 (O_1951,N_29452,N_29571);
nand UO_1952 (O_1952,N_29693,N_29941);
nand UO_1953 (O_1953,N_29922,N_29670);
nor UO_1954 (O_1954,N_29722,N_29764);
and UO_1955 (O_1955,N_29589,N_29817);
and UO_1956 (O_1956,N_29601,N_29905);
xnor UO_1957 (O_1957,N_29681,N_29796);
nor UO_1958 (O_1958,N_29492,N_29532);
nor UO_1959 (O_1959,N_29821,N_29575);
or UO_1960 (O_1960,N_29695,N_29707);
or UO_1961 (O_1961,N_29532,N_29790);
nor UO_1962 (O_1962,N_29611,N_29676);
and UO_1963 (O_1963,N_29534,N_29992);
and UO_1964 (O_1964,N_29692,N_29836);
xor UO_1965 (O_1965,N_29487,N_29528);
or UO_1966 (O_1966,N_29983,N_29466);
nand UO_1967 (O_1967,N_29576,N_29596);
nand UO_1968 (O_1968,N_29417,N_29746);
nor UO_1969 (O_1969,N_29715,N_29863);
or UO_1970 (O_1970,N_29946,N_29735);
and UO_1971 (O_1971,N_29696,N_29909);
nand UO_1972 (O_1972,N_29511,N_29935);
xor UO_1973 (O_1973,N_29781,N_29791);
nand UO_1974 (O_1974,N_29937,N_29899);
or UO_1975 (O_1975,N_29819,N_29601);
nand UO_1976 (O_1976,N_29971,N_29754);
and UO_1977 (O_1977,N_29858,N_29419);
nor UO_1978 (O_1978,N_29969,N_29719);
and UO_1979 (O_1979,N_29598,N_29645);
nand UO_1980 (O_1980,N_29728,N_29421);
nand UO_1981 (O_1981,N_29421,N_29612);
or UO_1982 (O_1982,N_29837,N_29523);
nor UO_1983 (O_1983,N_29616,N_29990);
xor UO_1984 (O_1984,N_29583,N_29839);
and UO_1985 (O_1985,N_29676,N_29851);
nand UO_1986 (O_1986,N_29637,N_29878);
or UO_1987 (O_1987,N_29417,N_29620);
nand UO_1988 (O_1988,N_29415,N_29581);
nand UO_1989 (O_1989,N_29926,N_29918);
or UO_1990 (O_1990,N_29889,N_29652);
and UO_1991 (O_1991,N_29937,N_29810);
xor UO_1992 (O_1992,N_29995,N_29726);
or UO_1993 (O_1993,N_29554,N_29709);
and UO_1994 (O_1994,N_29742,N_29937);
nor UO_1995 (O_1995,N_29478,N_29689);
and UO_1996 (O_1996,N_29730,N_29870);
nor UO_1997 (O_1997,N_29650,N_29785);
xnor UO_1998 (O_1998,N_29722,N_29945);
and UO_1999 (O_1999,N_29535,N_29678);
and UO_2000 (O_2000,N_29733,N_29476);
nand UO_2001 (O_2001,N_29595,N_29549);
xor UO_2002 (O_2002,N_29839,N_29522);
nand UO_2003 (O_2003,N_29505,N_29842);
nand UO_2004 (O_2004,N_29907,N_29721);
and UO_2005 (O_2005,N_29496,N_29556);
nor UO_2006 (O_2006,N_29793,N_29967);
and UO_2007 (O_2007,N_29819,N_29854);
or UO_2008 (O_2008,N_29736,N_29687);
and UO_2009 (O_2009,N_29481,N_29961);
nand UO_2010 (O_2010,N_29734,N_29946);
xnor UO_2011 (O_2011,N_29504,N_29989);
nor UO_2012 (O_2012,N_29465,N_29965);
xor UO_2013 (O_2013,N_29992,N_29681);
or UO_2014 (O_2014,N_29590,N_29616);
and UO_2015 (O_2015,N_29582,N_29719);
nand UO_2016 (O_2016,N_29976,N_29526);
nor UO_2017 (O_2017,N_29559,N_29864);
nor UO_2018 (O_2018,N_29594,N_29419);
nor UO_2019 (O_2019,N_29520,N_29469);
nor UO_2020 (O_2020,N_29696,N_29738);
nor UO_2021 (O_2021,N_29580,N_29951);
nand UO_2022 (O_2022,N_29989,N_29672);
or UO_2023 (O_2023,N_29532,N_29408);
and UO_2024 (O_2024,N_29778,N_29866);
nand UO_2025 (O_2025,N_29487,N_29584);
or UO_2026 (O_2026,N_29617,N_29952);
nor UO_2027 (O_2027,N_29864,N_29805);
nor UO_2028 (O_2028,N_29633,N_29597);
and UO_2029 (O_2029,N_29707,N_29551);
nor UO_2030 (O_2030,N_29833,N_29487);
nand UO_2031 (O_2031,N_29644,N_29992);
and UO_2032 (O_2032,N_29570,N_29950);
or UO_2033 (O_2033,N_29720,N_29554);
or UO_2034 (O_2034,N_29656,N_29555);
nor UO_2035 (O_2035,N_29884,N_29488);
or UO_2036 (O_2036,N_29756,N_29713);
or UO_2037 (O_2037,N_29552,N_29827);
nor UO_2038 (O_2038,N_29630,N_29747);
and UO_2039 (O_2039,N_29978,N_29586);
nand UO_2040 (O_2040,N_29690,N_29581);
nand UO_2041 (O_2041,N_29790,N_29987);
or UO_2042 (O_2042,N_29688,N_29751);
and UO_2043 (O_2043,N_29883,N_29601);
xnor UO_2044 (O_2044,N_29433,N_29683);
or UO_2045 (O_2045,N_29816,N_29639);
or UO_2046 (O_2046,N_29508,N_29547);
nor UO_2047 (O_2047,N_29596,N_29440);
or UO_2048 (O_2048,N_29442,N_29618);
and UO_2049 (O_2049,N_29809,N_29902);
nor UO_2050 (O_2050,N_29682,N_29423);
xor UO_2051 (O_2051,N_29810,N_29887);
nor UO_2052 (O_2052,N_29586,N_29524);
nor UO_2053 (O_2053,N_29665,N_29549);
xnor UO_2054 (O_2054,N_29742,N_29706);
and UO_2055 (O_2055,N_29910,N_29765);
or UO_2056 (O_2056,N_29789,N_29697);
nor UO_2057 (O_2057,N_29651,N_29641);
or UO_2058 (O_2058,N_29431,N_29556);
or UO_2059 (O_2059,N_29980,N_29930);
nand UO_2060 (O_2060,N_29417,N_29967);
nor UO_2061 (O_2061,N_29963,N_29617);
and UO_2062 (O_2062,N_29561,N_29446);
or UO_2063 (O_2063,N_29737,N_29458);
and UO_2064 (O_2064,N_29685,N_29743);
and UO_2065 (O_2065,N_29995,N_29626);
nor UO_2066 (O_2066,N_29532,N_29691);
or UO_2067 (O_2067,N_29952,N_29901);
or UO_2068 (O_2068,N_29544,N_29639);
xor UO_2069 (O_2069,N_29762,N_29495);
xor UO_2070 (O_2070,N_29736,N_29824);
nor UO_2071 (O_2071,N_29655,N_29931);
and UO_2072 (O_2072,N_29976,N_29533);
xnor UO_2073 (O_2073,N_29885,N_29950);
xor UO_2074 (O_2074,N_29635,N_29644);
nor UO_2075 (O_2075,N_29521,N_29579);
and UO_2076 (O_2076,N_29511,N_29516);
nand UO_2077 (O_2077,N_29633,N_29706);
and UO_2078 (O_2078,N_29496,N_29614);
nor UO_2079 (O_2079,N_29986,N_29948);
nand UO_2080 (O_2080,N_29460,N_29958);
xnor UO_2081 (O_2081,N_29544,N_29641);
and UO_2082 (O_2082,N_29823,N_29592);
or UO_2083 (O_2083,N_29451,N_29735);
and UO_2084 (O_2084,N_29998,N_29694);
or UO_2085 (O_2085,N_29621,N_29439);
nor UO_2086 (O_2086,N_29538,N_29515);
and UO_2087 (O_2087,N_29675,N_29563);
nand UO_2088 (O_2088,N_29776,N_29840);
or UO_2089 (O_2089,N_29571,N_29855);
xnor UO_2090 (O_2090,N_29694,N_29516);
and UO_2091 (O_2091,N_29809,N_29832);
or UO_2092 (O_2092,N_29428,N_29709);
nor UO_2093 (O_2093,N_29650,N_29657);
nand UO_2094 (O_2094,N_29504,N_29442);
or UO_2095 (O_2095,N_29759,N_29525);
nand UO_2096 (O_2096,N_29613,N_29474);
nand UO_2097 (O_2097,N_29527,N_29540);
and UO_2098 (O_2098,N_29835,N_29528);
nor UO_2099 (O_2099,N_29560,N_29479);
nor UO_2100 (O_2100,N_29519,N_29967);
or UO_2101 (O_2101,N_29402,N_29574);
nand UO_2102 (O_2102,N_29535,N_29645);
nand UO_2103 (O_2103,N_29678,N_29999);
or UO_2104 (O_2104,N_29481,N_29800);
and UO_2105 (O_2105,N_29767,N_29820);
or UO_2106 (O_2106,N_29999,N_29858);
and UO_2107 (O_2107,N_29810,N_29594);
and UO_2108 (O_2108,N_29849,N_29997);
nand UO_2109 (O_2109,N_29846,N_29484);
nor UO_2110 (O_2110,N_29992,N_29916);
nor UO_2111 (O_2111,N_29701,N_29450);
and UO_2112 (O_2112,N_29896,N_29841);
nand UO_2113 (O_2113,N_29538,N_29700);
nand UO_2114 (O_2114,N_29713,N_29409);
and UO_2115 (O_2115,N_29681,N_29831);
nand UO_2116 (O_2116,N_29408,N_29970);
or UO_2117 (O_2117,N_29818,N_29424);
nor UO_2118 (O_2118,N_29408,N_29419);
nor UO_2119 (O_2119,N_29724,N_29467);
nand UO_2120 (O_2120,N_29894,N_29836);
nand UO_2121 (O_2121,N_29743,N_29511);
and UO_2122 (O_2122,N_29456,N_29764);
nor UO_2123 (O_2123,N_29682,N_29666);
nand UO_2124 (O_2124,N_29653,N_29683);
nor UO_2125 (O_2125,N_29733,N_29478);
nand UO_2126 (O_2126,N_29609,N_29589);
nor UO_2127 (O_2127,N_29637,N_29748);
or UO_2128 (O_2128,N_29883,N_29963);
or UO_2129 (O_2129,N_29833,N_29404);
or UO_2130 (O_2130,N_29691,N_29919);
nor UO_2131 (O_2131,N_29993,N_29482);
and UO_2132 (O_2132,N_29552,N_29718);
and UO_2133 (O_2133,N_29475,N_29433);
or UO_2134 (O_2134,N_29570,N_29462);
and UO_2135 (O_2135,N_29837,N_29881);
nor UO_2136 (O_2136,N_29758,N_29440);
nor UO_2137 (O_2137,N_29892,N_29982);
xnor UO_2138 (O_2138,N_29989,N_29699);
or UO_2139 (O_2139,N_29475,N_29786);
and UO_2140 (O_2140,N_29730,N_29553);
nor UO_2141 (O_2141,N_29905,N_29806);
and UO_2142 (O_2142,N_29447,N_29734);
or UO_2143 (O_2143,N_29866,N_29418);
and UO_2144 (O_2144,N_29724,N_29581);
and UO_2145 (O_2145,N_29761,N_29815);
xnor UO_2146 (O_2146,N_29502,N_29734);
and UO_2147 (O_2147,N_29629,N_29657);
nand UO_2148 (O_2148,N_29803,N_29739);
and UO_2149 (O_2149,N_29719,N_29623);
and UO_2150 (O_2150,N_29747,N_29999);
nor UO_2151 (O_2151,N_29964,N_29659);
xor UO_2152 (O_2152,N_29448,N_29653);
nor UO_2153 (O_2153,N_29606,N_29923);
xnor UO_2154 (O_2154,N_29479,N_29565);
nand UO_2155 (O_2155,N_29768,N_29837);
or UO_2156 (O_2156,N_29626,N_29925);
and UO_2157 (O_2157,N_29603,N_29883);
and UO_2158 (O_2158,N_29426,N_29809);
or UO_2159 (O_2159,N_29450,N_29405);
nand UO_2160 (O_2160,N_29507,N_29677);
or UO_2161 (O_2161,N_29580,N_29736);
xnor UO_2162 (O_2162,N_29718,N_29814);
xor UO_2163 (O_2163,N_29840,N_29963);
xnor UO_2164 (O_2164,N_29994,N_29867);
or UO_2165 (O_2165,N_29843,N_29543);
or UO_2166 (O_2166,N_29982,N_29903);
nor UO_2167 (O_2167,N_29470,N_29674);
nor UO_2168 (O_2168,N_29627,N_29996);
or UO_2169 (O_2169,N_29622,N_29546);
nand UO_2170 (O_2170,N_29963,N_29414);
nor UO_2171 (O_2171,N_29684,N_29595);
nand UO_2172 (O_2172,N_29812,N_29647);
nand UO_2173 (O_2173,N_29765,N_29663);
nand UO_2174 (O_2174,N_29579,N_29630);
xnor UO_2175 (O_2175,N_29821,N_29765);
nor UO_2176 (O_2176,N_29979,N_29850);
nor UO_2177 (O_2177,N_29771,N_29720);
and UO_2178 (O_2178,N_29559,N_29534);
xnor UO_2179 (O_2179,N_29732,N_29733);
or UO_2180 (O_2180,N_29633,N_29835);
or UO_2181 (O_2181,N_29545,N_29416);
nand UO_2182 (O_2182,N_29608,N_29858);
nand UO_2183 (O_2183,N_29825,N_29786);
and UO_2184 (O_2184,N_29911,N_29631);
and UO_2185 (O_2185,N_29666,N_29927);
nor UO_2186 (O_2186,N_29479,N_29486);
and UO_2187 (O_2187,N_29453,N_29566);
or UO_2188 (O_2188,N_29600,N_29618);
nor UO_2189 (O_2189,N_29914,N_29771);
nor UO_2190 (O_2190,N_29763,N_29637);
or UO_2191 (O_2191,N_29426,N_29649);
and UO_2192 (O_2192,N_29484,N_29572);
and UO_2193 (O_2193,N_29905,N_29533);
nand UO_2194 (O_2194,N_29762,N_29804);
nor UO_2195 (O_2195,N_29838,N_29859);
nor UO_2196 (O_2196,N_29699,N_29995);
nor UO_2197 (O_2197,N_29838,N_29690);
and UO_2198 (O_2198,N_29765,N_29535);
nand UO_2199 (O_2199,N_29554,N_29493);
or UO_2200 (O_2200,N_29603,N_29753);
nor UO_2201 (O_2201,N_29544,N_29506);
and UO_2202 (O_2202,N_29768,N_29748);
nand UO_2203 (O_2203,N_29927,N_29663);
and UO_2204 (O_2204,N_29648,N_29901);
and UO_2205 (O_2205,N_29962,N_29936);
or UO_2206 (O_2206,N_29748,N_29412);
and UO_2207 (O_2207,N_29579,N_29626);
and UO_2208 (O_2208,N_29915,N_29675);
nand UO_2209 (O_2209,N_29932,N_29654);
nor UO_2210 (O_2210,N_29929,N_29924);
nor UO_2211 (O_2211,N_29433,N_29412);
nor UO_2212 (O_2212,N_29824,N_29900);
xnor UO_2213 (O_2213,N_29842,N_29487);
or UO_2214 (O_2214,N_29900,N_29805);
nor UO_2215 (O_2215,N_29753,N_29971);
nand UO_2216 (O_2216,N_29402,N_29762);
and UO_2217 (O_2217,N_29897,N_29844);
nand UO_2218 (O_2218,N_29699,N_29996);
and UO_2219 (O_2219,N_29814,N_29864);
and UO_2220 (O_2220,N_29836,N_29449);
and UO_2221 (O_2221,N_29820,N_29418);
or UO_2222 (O_2222,N_29879,N_29537);
nor UO_2223 (O_2223,N_29500,N_29569);
or UO_2224 (O_2224,N_29699,N_29871);
and UO_2225 (O_2225,N_29897,N_29813);
nor UO_2226 (O_2226,N_29486,N_29770);
nand UO_2227 (O_2227,N_29578,N_29711);
nand UO_2228 (O_2228,N_29958,N_29468);
nor UO_2229 (O_2229,N_29516,N_29774);
and UO_2230 (O_2230,N_29850,N_29678);
nor UO_2231 (O_2231,N_29526,N_29459);
nand UO_2232 (O_2232,N_29794,N_29626);
and UO_2233 (O_2233,N_29958,N_29735);
and UO_2234 (O_2234,N_29412,N_29521);
or UO_2235 (O_2235,N_29975,N_29634);
nand UO_2236 (O_2236,N_29703,N_29557);
or UO_2237 (O_2237,N_29489,N_29692);
xor UO_2238 (O_2238,N_29449,N_29408);
nand UO_2239 (O_2239,N_29837,N_29858);
nand UO_2240 (O_2240,N_29813,N_29697);
or UO_2241 (O_2241,N_29750,N_29677);
nor UO_2242 (O_2242,N_29904,N_29811);
or UO_2243 (O_2243,N_29863,N_29880);
and UO_2244 (O_2244,N_29855,N_29525);
or UO_2245 (O_2245,N_29480,N_29979);
or UO_2246 (O_2246,N_29602,N_29944);
and UO_2247 (O_2247,N_29860,N_29786);
nand UO_2248 (O_2248,N_29951,N_29581);
and UO_2249 (O_2249,N_29904,N_29938);
or UO_2250 (O_2250,N_29471,N_29846);
nand UO_2251 (O_2251,N_29599,N_29834);
nand UO_2252 (O_2252,N_29412,N_29661);
nand UO_2253 (O_2253,N_29568,N_29785);
nand UO_2254 (O_2254,N_29596,N_29834);
or UO_2255 (O_2255,N_29479,N_29784);
and UO_2256 (O_2256,N_29822,N_29670);
or UO_2257 (O_2257,N_29671,N_29797);
and UO_2258 (O_2258,N_29675,N_29629);
and UO_2259 (O_2259,N_29427,N_29644);
nor UO_2260 (O_2260,N_29474,N_29942);
and UO_2261 (O_2261,N_29840,N_29560);
and UO_2262 (O_2262,N_29693,N_29715);
nand UO_2263 (O_2263,N_29560,N_29933);
or UO_2264 (O_2264,N_29590,N_29948);
xnor UO_2265 (O_2265,N_29794,N_29660);
nor UO_2266 (O_2266,N_29820,N_29791);
nor UO_2267 (O_2267,N_29722,N_29944);
nand UO_2268 (O_2268,N_29696,N_29994);
or UO_2269 (O_2269,N_29792,N_29676);
nor UO_2270 (O_2270,N_29932,N_29830);
nand UO_2271 (O_2271,N_29716,N_29895);
xor UO_2272 (O_2272,N_29785,N_29988);
nor UO_2273 (O_2273,N_29553,N_29425);
or UO_2274 (O_2274,N_29872,N_29699);
nand UO_2275 (O_2275,N_29456,N_29798);
and UO_2276 (O_2276,N_29965,N_29757);
and UO_2277 (O_2277,N_29950,N_29630);
nor UO_2278 (O_2278,N_29647,N_29726);
xor UO_2279 (O_2279,N_29450,N_29960);
nor UO_2280 (O_2280,N_29424,N_29502);
nor UO_2281 (O_2281,N_29579,N_29411);
nor UO_2282 (O_2282,N_29789,N_29519);
and UO_2283 (O_2283,N_29652,N_29820);
nor UO_2284 (O_2284,N_29953,N_29892);
and UO_2285 (O_2285,N_29966,N_29995);
or UO_2286 (O_2286,N_29793,N_29775);
nand UO_2287 (O_2287,N_29423,N_29424);
and UO_2288 (O_2288,N_29862,N_29722);
and UO_2289 (O_2289,N_29506,N_29970);
or UO_2290 (O_2290,N_29526,N_29529);
nand UO_2291 (O_2291,N_29558,N_29597);
nand UO_2292 (O_2292,N_29855,N_29481);
or UO_2293 (O_2293,N_29441,N_29449);
and UO_2294 (O_2294,N_29838,N_29615);
nor UO_2295 (O_2295,N_29891,N_29609);
nand UO_2296 (O_2296,N_29673,N_29472);
or UO_2297 (O_2297,N_29955,N_29779);
and UO_2298 (O_2298,N_29976,N_29885);
or UO_2299 (O_2299,N_29667,N_29855);
nand UO_2300 (O_2300,N_29467,N_29729);
nor UO_2301 (O_2301,N_29401,N_29510);
nor UO_2302 (O_2302,N_29708,N_29715);
and UO_2303 (O_2303,N_29450,N_29640);
nand UO_2304 (O_2304,N_29910,N_29520);
nand UO_2305 (O_2305,N_29602,N_29971);
nor UO_2306 (O_2306,N_29588,N_29669);
xor UO_2307 (O_2307,N_29901,N_29654);
and UO_2308 (O_2308,N_29653,N_29808);
or UO_2309 (O_2309,N_29598,N_29979);
nor UO_2310 (O_2310,N_29472,N_29691);
nor UO_2311 (O_2311,N_29926,N_29892);
nor UO_2312 (O_2312,N_29532,N_29929);
or UO_2313 (O_2313,N_29543,N_29876);
or UO_2314 (O_2314,N_29748,N_29676);
nand UO_2315 (O_2315,N_29616,N_29517);
nand UO_2316 (O_2316,N_29449,N_29737);
nor UO_2317 (O_2317,N_29812,N_29893);
and UO_2318 (O_2318,N_29603,N_29426);
and UO_2319 (O_2319,N_29881,N_29726);
xnor UO_2320 (O_2320,N_29624,N_29726);
xor UO_2321 (O_2321,N_29951,N_29421);
and UO_2322 (O_2322,N_29422,N_29474);
and UO_2323 (O_2323,N_29635,N_29715);
and UO_2324 (O_2324,N_29655,N_29936);
or UO_2325 (O_2325,N_29960,N_29442);
nor UO_2326 (O_2326,N_29410,N_29430);
and UO_2327 (O_2327,N_29824,N_29805);
or UO_2328 (O_2328,N_29420,N_29962);
nand UO_2329 (O_2329,N_29795,N_29790);
xor UO_2330 (O_2330,N_29608,N_29903);
and UO_2331 (O_2331,N_29817,N_29998);
nor UO_2332 (O_2332,N_29626,N_29883);
or UO_2333 (O_2333,N_29503,N_29966);
or UO_2334 (O_2334,N_29905,N_29874);
and UO_2335 (O_2335,N_29508,N_29909);
nor UO_2336 (O_2336,N_29589,N_29558);
nor UO_2337 (O_2337,N_29665,N_29877);
or UO_2338 (O_2338,N_29535,N_29651);
xnor UO_2339 (O_2339,N_29757,N_29830);
nand UO_2340 (O_2340,N_29423,N_29901);
xnor UO_2341 (O_2341,N_29832,N_29853);
nand UO_2342 (O_2342,N_29896,N_29783);
nor UO_2343 (O_2343,N_29450,N_29657);
and UO_2344 (O_2344,N_29616,N_29962);
nand UO_2345 (O_2345,N_29531,N_29887);
or UO_2346 (O_2346,N_29455,N_29922);
xor UO_2347 (O_2347,N_29415,N_29711);
and UO_2348 (O_2348,N_29434,N_29576);
nor UO_2349 (O_2349,N_29538,N_29964);
and UO_2350 (O_2350,N_29727,N_29971);
or UO_2351 (O_2351,N_29541,N_29908);
or UO_2352 (O_2352,N_29879,N_29592);
nand UO_2353 (O_2353,N_29884,N_29708);
nor UO_2354 (O_2354,N_29567,N_29615);
and UO_2355 (O_2355,N_29434,N_29677);
nor UO_2356 (O_2356,N_29648,N_29927);
nor UO_2357 (O_2357,N_29510,N_29794);
and UO_2358 (O_2358,N_29769,N_29418);
nor UO_2359 (O_2359,N_29705,N_29580);
nor UO_2360 (O_2360,N_29729,N_29726);
nor UO_2361 (O_2361,N_29838,N_29700);
or UO_2362 (O_2362,N_29610,N_29416);
nand UO_2363 (O_2363,N_29878,N_29926);
or UO_2364 (O_2364,N_29529,N_29463);
and UO_2365 (O_2365,N_29888,N_29701);
nor UO_2366 (O_2366,N_29669,N_29646);
or UO_2367 (O_2367,N_29689,N_29800);
xor UO_2368 (O_2368,N_29794,N_29590);
nand UO_2369 (O_2369,N_29800,N_29578);
or UO_2370 (O_2370,N_29890,N_29862);
and UO_2371 (O_2371,N_29614,N_29944);
nand UO_2372 (O_2372,N_29692,N_29711);
or UO_2373 (O_2373,N_29668,N_29991);
or UO_2374 (O_2374,N_29582,N_29770);
nand UO_2375 (O_2375,N_29844,N_29827);
nor UO_2376 (O_2376,N_29417,N_29682);
nor UO_2377 (O_2377,N_29603,N_29550);
or UO_2378 (O_2378,N_29487,N_29741);
nand UO_2379 (O_2379,N_29573,N_29663);
nor UO_2380 (O_2380,N_29896,N_29493);
nor UO_2381 (O_2381,N_29722,N_29991);
and UO_2382 (O_2382,N_29902,N_29993);
nand UO_2383 (O_2383,N_29457,N_29489);
nor UO_2384 (O_2384,N_29837,N_29898);
and UO_2385 (O_2385,N_29541,N_29581);
xnor UO_2386 (O_2386,N_29644,N_29614);
nor UO_2387 (O_2387,N_29469,N_29506);
nand UO_2388 (O_2388,N_29411,N_29857);
or UO_2389 (O_2389,N_29586,N_29805);
and UO_2390 (O_2390,N_29582,N_29552);
or UO_2391 (O_2391,N_29946,N_29689);
nand UO_2392 (O_2392,N_29736,N_29604);
nand UO_2393 (O_2393,N_29654,N_29753);
xor UO_2394 (O_2394,N_29566,N_29749);
or UO_2395 (O_2395,N_29662,N_29834);
xor UO_2396 (O_2396,N_29693,N_29773);
nor UO_2397 (O_2397,N_29797,N_29682);
and UO_2398 (O_2398,N_29927,N_29590);
and UO_2399 (O_2399,N_29524,N_29904);
nand UO_2400 (O_2400,N_29582,N_29497);
xnor UO_2401 (O_2401,N_29403,N_29597);
nand UO_2402 (O_2402,N_29991,N_29765);
xnor UO_2403 (O_2403,N_29682,N_29583);
nand UO_2404 (O_2404,N_29554,N_29990);
xnor UO_2405 (O_2405,N_29836,N_29814);
and UO_2406 (O_2406,N_29564,N_29931);
or UO_2407 (O_2407,N_29590,N_29739);
xor UO_2408 (O_2408,N_29696,N_29796);
nor UO_2409 (O_2409,N_29487,N_29510);
and UO_2410 (O_2410,N_29798,N_29945);
or UO_2411 (O_2411,N_29557,N_29635);
nor UO_2412 (O_2412,N_29891,N_29533);
xnor UO_2413 (O_2413,N_29972,N_29436);
and UO_2414 (O_2414,N_29458,N_29856);
nand UO_2415 (O_2415,N_29740,N_29575);
nand UO_2416 (O_2416,N_29455,N_29545);
and UO_2417 (O_2417,N_29602,N_29674);
or UO_2418 (O_2418,N_29651,N_29974);
nor UO_2419 (O_2419,N_29831,N_29522);
and UO_2420 (O_2420,N_29905,N_29418);
nor UO_2421 (O_2421,N_29689,N_29721);
or UO_2422 (O_2422,N_29537,N_29772);
or UO_2423 (O_2423,N_29956,N_29431);
or UO_2424 (O_2424,N_29527,N_29720);
nor UO_2425 (O_2425,N_29411,N_29977);
xnor UO_2426 (O_2426,N_29817,N_29642);
or UO_2427 (O_2427,N_29631,N_29471);
nor UO_2428 (O_2428,N_29613,N_29604);
or UO_2429 (O_2429,N_29888,N_29531);
nor UO_2430 (O_2430,N_29665,N_29674);
nor UO_2431 (O_2431,N_29449,N_29818);
nand UO_2432 (O_2432,N_29617,N_29454);
or UO_2433 (O_2433,N_29413,N_29909);
nand UO_2434 (O_2434,N_29473,N_29593);
nor UO_2435 (O_2435,N_29663,N_29945);
and UO_2436 (O_2436,N_29761,N_29599);
nand UO_2437 (O_2437,N_29995,N_29534);
xor UO_2438 (O_2438,N_29414,N_29820);
and UO_2439 (O_2439,N_29703,N_29752);
nor UO_2440 (O_2440,N_29716,N_29836);
or UO_2441 (O_2441,N_29736,N_29595);
nor UO_2442 (O_2442,N_29801,N_29767);
nand UO_2443 (O_2443,N_29807,N_29906);
nor UO_2444 (O_2444,N_29795,N_29884);
and UO_2445 (O_2445,N_29804,N_29783);
and UO_2446 (O_2446,N_29608,N_29829);
nor UO_2447 (O_2447,N_29740,N_29587);
nor UO_2448 (O_2448,N_29899,N_29513);
nand UO_2449 (O_2449,N_29752,N_29606);
nand UO_2450 (O_2450,N_29646,N_29717);
and UO_2451 (O_2451,N_29926,N_29936);
nor UO_2452 (O_2452,N_29727,N_29966);
xnor UO_2453 (O_2453,N_29460,N_29402);
nor UO_2454 (O_2454,N_29716,N_29944);
and UO_2455 (O_2455,N_29468,N_29782);
nand UO_2456 (O_2456,N_29543,N_29952);
xor UO_2457 (O_2457,N_29616,N_29887);
nor UO_2458 (O_2458,N_29909,N_29775);
nand UO_2459 (O_2459,N_29878,N_29545);
nor UO_2460 (O_2460,N_29532,N_29988);
nor UO_2461 (O_2461,N_29838,N_29561);
nor UO_2462 (O_2462,N_29552,N_29839);
or UO_2463 (O_2463,N_29975,N_29739);
nor UO_2464 (O_2464,N_29552,N_29854);
or UO_2465 (O_2465,N_29448,N_29988);
nor UO_2466 (O_2466,N_29725,N_29945);
or UO_2467 (O_2467,N_29875,N_29640);
nor UO_2468 (O_2468,N_29739,N_29644);
or UO_2469 (O_2469,N_29556,N_29832);
and UO_2470 (O_2470,N_29689,N_29443);
or UO_2471 (O_2471,N_29485,N_29930);
and UO_2472 (O_2472,N_29776,N_29901);
and UO_2473 (O_2473,N_29927,N_29909);
and UO_2474 (O_2474,N_29899,N_29828);
xor UO_2475 (O_2475,N_29459,N_29425);
or UO_2476 (O_2476,N_29695,N_29705);
nor UO_2477 (O_2477,N_29642,N_29828);
and UO_2478 (O_2478,N_29817,N_29827);
or UO_2479 (O_2479,N_29709,N_29973);
nor UO_2480 (O_2480,N_29688,N_29965);
nor UO_2481 (O_2481,N_29763,N_29953);
nor UO_2482 (O_2482,N_29914,N_29732);
and UO_2483 (O_2483,N_29837,N_29885);
nand UO_2484 (O_2484,N_29737,N_29921);
nand UO_2485 (O_2485,N_29414,N_29824);
nor UO_2486 (O_2486,N_29540,N_29489);
nor UO_2487 (O_2487,N_29565,N_29422);
nand UO_2488 (O_2488,N_29682,N_29424);
or UO_2489 (O_2489,N_29430,N_29840);
xor UO_2490 (O_2490,N_29419,N_29557);
and UO_2491 (O_2491,N_29615,N_29481);
nor UO_2492 (O_2492,N_29931,N_29680);
and UO_2493 (O_2493,N_29569,N_29581);
and UO_2494 (O_2494,N_29755,N_29854);
and UO_2495 (O_2495,N_29800,N_29681);
nor UO_2496 (O_2496,N_29732,N_29413);
and UO_2497 (O_2497,N_29996,N_29608);
or UO_2498 (O_2498,N_29932,N_29652);
nor UO_2499 (O_2499,N_29679,N_29605);
nand UO_2500 (O_2500,N_29538,N_29761);
nand UO_2501 (O_2501,N_29761,N_29660);
nand UO_2502 (O_2502,N_29402,N_29622);
nor UO_2503 (O_2503,N_29975,N_29531);
and UO_2504 (O_2504,N_29985,N_29805);
or UO_2505 (O_2505,N_29874,N_29820);
and UO_2506 (O_2506,N_29565,N_29489);
nor UO_2507 (O_2507,N_29509,N_29485);
and UO_2508 (O_2508,N_29969,N_29709);
nand UO_2509 (O_2509,N_29719,N_29571);
xnor UO_2510 (O_2510,N_29720,N_29860);
and UO_2511 (O_2511,N_29964,N_29984);
or UO_2512 (O_2512,N_29687,N_29798);
xor UO_2513 (O_2513,N_29515,N_29645);
nor UO_2514 (O_2514,N_29576,N_29463);
and UO_2515 (O_2515,N_29922,N_29789);
nand UO_2516 (O_2516,N_29501,N_29783);
nand UO_2517 (O_2517,N_29810,N_29510);
or UO_2518 (O_2518,N_29415,N_29819);
nor UO_2519 (O_2519,N_29683,N_29957);
and UO_2520 (O_2520,N_29460,N_29497);
nor UO_2521 (O_2521,N_29793,N_29922);
nor UO_2522 (O_2522,N_29939,N_29447);
xor UO_2523 (O_2523,N_29514,N_29435);
xnor UO_2524 (O_2524,N_29457,N_29485);
nor UO_2525 (O_2525,N_29506,N_29610);
nor UO_2526 (O_2526,N_29612,N_29854);
and UO_2527 (O_2527,N_29824,N_29937);
and UO_2528 (O_2528,N_29556,N_29591);
nor UO_2529 (O_2529,N_29928,N_29592);
xor UO_2530 (O_2530,N_29619,N_29612);
nand UO_2531 (O_2531,N_29784,N_29909);
or UO_2532 (O_2532,N_29511,N_29839);
nor UO_2533 (O_2533,N_29450,N_29505);
and UO_2534 (O_2534,N_29437,N_29887);
or UO_2535 (O_2535,N_29770,N_29472);
nor UO_2536 (O_2536,N_29484,N_29984);
nor UO_2537 (O_2537,N_29658,N_29419);
and UO_2538 (O_2538,N_29485,N_29726);
or UO_2539 (O_2539,N_29891,N_29519);
and UO_2540 (O_2540,N_29732,N_29510);
nand UO_2541 (O_2541,N_29704,N_29472);
nand UO_2542 (O_2542,N_29965,N_29852);
or UO_2543 (O_2543,N_29500,N_29889);
and UO_2544 (O_2544,N_29951,N_29526);
nor UO_2545 (O_2545,N_29724,N_29406);
or UO_2546 (O_2546,N_29403,N_29653);
or UO_2547 (O_2547,N_29997,N_29401);
and UO_2548 (O_2548,N_29954,N_29409);
nor UO_2549 (O_2549,N_29436,N_29824);
nand UO_2550 (O_2550,N_29784,N_29401);
nand UO_2551 (O_2551,N_29420,N_29975);
nand UO_2552 (O_2552,N_29412,N_29487);
and UO_2553 (O_2553,N_29789,N_29515);
nor UO_2554 (O_2554,N_29531,N_29747);
xor UO_2555 (O_2555,N_29741,N_29664);
nand UO_2556 (O_2556,N_29585,N_29904);
xor UO_2557 (O_2557,N_29750,N_29683);
nor UO_2558 (O_2558,N_29905,N_29939);
and UO_2559 (O_2559,N_29790,N_29410);
and UO_2560 (O_2560,N_29756,N_29924);
or UO_2561 (O_2561,N_29581,N_29412);
or UO_2562 (O_2562,N_29564,N_29405);
or UO_2563 (O_2563,N_29660,N_29421);
and UO_2564 (O_2564,N_29495,N_29730);
xor UO_2565 (O_2565,N_29424,N_29515);
or UO_2566 (O_2566,N_29495,N_29560);
nor UO_2567 (O_2567,N_29987,N_29651);
nor UO_2568 (O_2568,N_29463,N_29538);
or UO_2569 (O_2569,N_29504,N_29591);
and UO_2570 (O_2570,N_29875,N_29809);
or UO_2571 (O_2571,N_29870,N_29546);
xor UO_2572 (O_2572,N_29895,N_29972);
nor UO_2573 (O_2573,N_29451,N_29937);
nor UO_2574 (O_2574,N_29428,N_29468);
and UO_2575 (O_2575,N_29424,N_29595);
xnor UO_2576 (O_2576,N_29499,N_29691);
nor UO_2577 (O_2577,N_29525,N_29811);
or UO_2578 (O_2578,N_29750,N_29581);
nand UO_2579 (O_2579,N_29766,N_29799);
nand UO_2580 (O_2580,N_29957,N_29490);
and UO_2581 (O_2581,N_29467,N_29751);
nand UO_2582 (O_2582,N_29977,N_29510);
or UO_2583 (O_2583,N_29893,N_29414);
nand UO_2584 (O_2584,N_29555,N_29465);
and UO_2585 (O_2585,N_29820,N_29471);
or UO_2586 (O_2586,N_29552,N_29432);
nor UO_2587 (O_2587,N_29780,N_29930);
nor UO_2588 (O_2588,N_29590,N_29880);
nor UO_2589 (O_2589,N_29567,N_29954);
and UO_2590 (O_2590,N_29574,N_29660);
or UO_2591 (O_2591,N_29522,N_29914);
nor UO_2592 (O_2592,N_29434,N_29953);
and UO_2593 (O_2593,N_29722,N_29726);
nand UO_2594 (O_2594,N_29417,N_29826);
nand UO_2595 (O_2595,N_29421,N_29859);
xor UO_2596 (O_2596,N_29582,N_29963);
and UO_2597 (O_2597,N_29693,N_29871);
and UO_2598 (O_2598,N_29423,N_29547);
nor UO_2599 (O_2599,N_29826,N_29939);
nand UO_2600 (O_2600,N_29480,N_29557);
nor UO_2601 (O_2601,N_29998,N_29766);
and UO_2602 (O_2602,N_29549,N_29512);
xor UO_2603 (O_2603,N_29564,N_29763);
nor UO_2604 (O_2604,N_29898,N_29751);
nand UO_2605 (O_2605,N_29695,N_29940);
nand UO_2606 (O_2606,N_29731,N_29512);
nor UO_2607 (O_2607,N_29872,N_29481);
and UO_2608 (O_2608,N_29859,N_29491);
and UO_2609 (O_2609,N_29408,N_29629);
and UO_2610 (O_2610,N_29791,N_29722);
nand UO_2611 (O_2611,N_29776,N_29743);
and UO_2612 (O_2612,N_29437,N_29977);
nand UO_2613 (O_2613,N_29590,N_29419);
nor UO_2614 (O_2614,N_29738,N_29970);
nor UO_2615 (O_2615,N_29413,N_29892);
and UO_2616 (O_2616,N_29985,N_29754);
nand UO_2617 (O_2617,N_29490,N_29435);
nor UO_2618 (O_2618,N_29523,N_29674);
nor UO_2619 (O_2619,N_29613,N_29561);
and UO_2620 (O_2620,N_29623,N_29984);
or UO_2621 (O_2621,N_29935,N_29686);
nand UO_2622 (O_2622,N_29886,N_29899);
and UO_2623 (O_2623,N_29621,N_29507);
nand UO_2624 (O_2624,N_29615,N_29642);
or UO_2625 (O_2625,N_29411,N_29533);
or UO_2626 (O_2626,N_29574,N_29618);
nand UO_2627 (O_2627,N_29689,N_29847);
nor UO_2628 (O_2628,N_29737,N_29915);
nor UO_2629 (O_2629,N_29521,N_29458);
and UO_2630 (O_2630,N_29829,N_29860);
or UO_2631 (O_2631,N_29535,N_29959);
and UO_2632 (O_2632,N_29664,N_29473);
and UO_2633 (O_2633,N_29879,N_29560);
nor UO_2634 (O_2634,N_29401,N_29419);
nor UO_2635 (O_2635,N_29502,N_29673);
xor UO_2636 (O_2636,N_29877,N_29423);
or UO_2637 (O_2637,N_29442,N_29526);
nor UO_2638 (O_2638,N_29722,N_29691);
or UO_2639 (O_2639,N_29809,N_29941);
xnor UO_2640 (O_2640,N_29613,N_29422);
nor UO_2641 (O_2641,N_29518,N_29868);
and UO_2642 (O_2642,N_29982,N_29890);
nor UO_2643 (O_2643,N_29737,N_29721);
nand UO_2644 (O_2644,N_29729,N_29541);
and UO_2645 (O_2645,N_29823,N_29589);
or UO_2646 (O_2646,N_29528,N_29635);
xor UO_2647 (O_2647,N_29824,N_29614);
and UO_2648 (O_2648,N_29764,N_29465);
nand UO_2649 (O_2649,N_29724,N_29767);
nor UO_2650 (O_2650,N_29456,N_29978);
nand UO_2651 (O_2651,N_29960,N_29795);
nor UO_2652 (O_2652,N_29833,N_29968);
nand UO_2653 (O_2653,N_29479,N_29541);
nand UO_2654 (O_2654,N_29541,N_29587);
or UO_2655 (O_2655,N_29599,N_29400);
and UO_2656 (O_2656,N_29792,N_29940);
nand UO_2657 (O_2657,N_29951,N_29509);
xor UO_2658 (O_2658,N_29994,N_29468);
nor UO_2659 (O_2659,N_29675,N_29436);
nand UO_2660 (O_2660,N_29895,N_29912);
nand UO_2661 (O_2661,N_29963,N_29729);
or UO_2662 (O_2662,N_29497,N_29868);
and UO_2663 (O_2663,N_29929,N_29611);
or UO_2664 (O_2664,N_29626,N_29587);
and UO_2665 (O_2665,N_29572,N_29773);
xor UO_2666 (O_2666,N_29930,N_29605);
nor UO_2667 (O_2667,N_29510,N_29560);
nor UO_2668 (O_2668,N_29625,N_29751);
nand UO_2669 (O_2669,N_29881,N_29513);
nor UO_2670 (O_2670,N_29488,N_29964);
nand UO_2671 (O_2671,N_29985,N_29942);
nand UO_2672 (O_2672,N_29420,N_29742);
or UO_2673 (O_2673,N_29865,N_29410);
nand UO_2674 (O_2674,N_29684,N_29804);
or UO_2675 (O_2675,N_29401,N_29941);
nor UO_2676 (O_2676,N_29622,N_29879);
xnor UO_2677 (O_2677,N_29713,N_29889);
nand UO_2678 (O_2678,N_29703,N_29895);
xor UO_2679 (O_2679,N_29899,N_29961);
and UO_2680 (O_2680,N_29440,N_29781);
nand UO_2681 (O_2681,N_29541,N_29432);
or UO_2682 (O_2682,N_29874,N_29606);
nand UO_2683 (O_2683,N_29468,N_29653);
nand UO_2684 (O_2684,N_29867,N_29626);
and UO_2685 (O_2685,N_29639,N_29671);
and UO_2686 (O_2686,N_29847,N_29740);
or UO_2687 (O_2687,N_29432,N_29466);
or UO_2688 (O_2688,N_29422,N_29903);
and UO_2689 (O_2689,N_29712,N_29409);
xor UO_2690 (O_2690,N_29415,N_29627);
nor UO_2691 (O_2691,N_29764,N_29425);
and UO_2692 (O_2692,N_29431,N_29685);
nand UO_2693 (O_2693,N_29724,N_29610);
xnor UO_2694 (O_2694,N_29873,N_29454);
nand UO_2695 (O_2695,N_29918,N_29507);
or UO_2696 (O_2696,N_29709,N_29681);
or UO_2697 (O_2697,N_29475,N_29495);
nand UO_2698 (O_2698,N_29853,N_29614);
nand UO_2699 (O_2699,N_29524,N_29956);
xor UO_2700 (O_2700,N_29972,N_29660);
or UO_2701 (O_2701,N_29466,N_29822);
xnor UO_2702 (O_2702,N_29979,N_29910);
nand UO_2703 (O_2703,N_29503,N_29847);
nor UO_2704 (O_2704,N_29912,N_29994);
and UO_2705 (O_2705,N_29473,N_29678);
nand UO_2706 (O_2706,N_29813,N_29781);
and UO_2707 (O_2707,N_29654,N_29736);
nand UO_2708 (O_2708,N_29412,N_29741);
nand UO_2709 (O_2709,N_29909,N_29501);
and UO_2710 (O_2710,N_29785,N_29657);
and UO_2711 (O_2711,N_29682,N_29826);
nand UO_2712 (O_2712,N_29607,N_29693);
nor UO_2713 (O_2713,N_29709,N_29620);
and UO_2714 (O_2714,N_29818,N_29960);
and UO_2715 (O_2715,N_29806,N_29509);
or UO_2716 (O_2716,N_29580,N_29992);
xnor UO_2717 (O_2717,N_29741,N_29528);
and UO_2718 (O_2718,N_29555,N_29420);
nor UO_2719 (O_2719,N_29477,N_29845);
nor UO_2720 (O_2720,N_29966,N_29447);
nand UO_2721 (O_2721,N_29581,N_29797);
and UO_2722 (O_2722,N_29534,N_29734);
nor UO_2723 (O_2723,N_29943,N_29832);
or UO_2724 (O_2724,N_29488,N_29786);
or UO_2725 (O_2725,N_29984,N_29579);
nor UO_2726 (O_2726,N_29489,N_29612);
nor UO_2727 (O_2727,N_29424,N_29863);
nand UO_2728 (O_2728,N_29848,N_29972);
nand UO_2729 (O_2729,N_29806,N_29964);
nor UO_2730 (O_2730,N_29931,N_29555);
nand UO_2731 (O_2731,N_29490,N_29514);
or UO_2732 (O_2732,N_29700,N_29830);
nor UO_2733 (O_2733,N_29717,N_29963);
nor UO_2734 (O_2734,N_29438,N_29809);
xnor UO_2735 (O_2735,N_29570,N_29452);
or UO_2736 (O_2736,N_29581,N_29886);
or UO_2737 (O_2737,N_29523,N_29590);
nand UO_2738 (O_2738,N_29719,N_29622);
nand UO_2739 (O_2739,N_29652,N_29416);
xnor UO_2740 (O_2740,N_29955,N_29407);
nand UO_2741 (O_2741,N_29649,N_29947);
and UO_2742 (O_2742,N_29617,N_29818);
nand UO_2743 (O_2743,N_29984,N_29947);
or UO_2744 (O_2744,N_29692,N_29466);
nand UO_2745 (O_2745,N_29508,N_29891);
nor UO_2746 (O_2746,N_29607,N_29961);
nand UO_2747 (O_2747,N_29865,N_29771);
nand UO_2748 (O_2748,N_29975,N_29876);
or UO_2749 (O_2749,N_29897,N_29859);
and UO_2750 (O_2750,N_29712,N_29546);
nand UO_2751 (O_2751,N_29757,N_29493);
and UO_2752 (O_2752,N_29813,N_29948);
nand UO_2753 (O_2753,N_29788,N_29590);
nor UO_2754 (O_2754,N_29450,N_29920);
nand UO_2755 (O_2755,N_29537,N_29510);
nor UO_2756 (O_2756,N_29844,N_29758);
and UO_2757 (O_2757,N_29492,N_29584);
and UO_2758 (O_2758,N_29858,N_29417);
nand UO_2759 (O_2759,N_29835,N_29870);
or UO_2760 (O_2760,N_29470,N_29858);
or UO_2761 (O_2761,N_29694,N_29484);
and UO_2762 (O_2762,N_29951,N_29644);
or UO_2763 (O_2763,N_29725,N_29421);
or UO_2764 (O_2764,N_29883,N_29801);
and UO_2765 (O_2765,N_29990,N_29730);
nor UO_2766 (O_2766,N_29645,N_29943);
nand UO_2767 (O_2767,N_29952,N_29624);
xnor UO_2768 (O_2768,N_29602,N_29445);
and UO_2769 (O_2769,N_29616,N_29402);
nor UO_2770 (O_2770,N_29581,N_29414);
nor UO_2771 (O_2771,N_29652,N_29618);
nor UO_2772 (O_2772,N_29502,N_29809);
nor UO_2773 (O_2773,N_29464,N_29733);
and UO_2774 (O_2774,N_29784,N_29733);
or UO_2775 (O_2775,N_29817,N_29565);
nand UO_2776 (O_2776,N_29996,N_29454);
or UO_2777 (O_2777,N_29445,N_29742);
nand UO_2778 (O_2778,N_29897,N_29905);
xnor UO_2779 (O_2779,N_29965,N_29926);
nand UO_2780 (O_2780,N_29975,N_29522);
nor UO_2781 (O_2781,N_29769,N_29757);
nand UO_2782 (O_2782,N_29783,N_29757);
nor UO_2783 (O_2783,N_29577,N_29870);
nor UO_2784 (O_2784,N_29534,N_29642);
nand UO_2785 (O_2785,N_29915,N_29990);
and UO_2786 (O_2786,N_29790,N_29803);
nor UO_2787 (O_2787,N_29612,N_29462);
nand UO_2788 (O_2788,N_29889,N_29422);
xnor UO_2789 (O_2789,N_29781,N_29605);
or UO_2790 (O_2790,N_29427,N_29496);
and UO_2791 (O_2791,N_29719,N_29450);
and UO_2792 (O_2792,N_29724,N_29737);
or UO_2793 (O_2793,N_29437,N_29922);
nor UO_2794 (O_2794,N_29876,N_29914);
or UO_2795 (O_2795,N_29671,N_29547);
nor UO_2796 (O_2796,N_29537,N_29863);
or UO_2797 (O_2797,N_29969,N_29666);
and UO_2798 (O_2798,N_29953,N_29543);
xor UO_2799 (O_2799,N_29971,N_29730);
nor UO_2800 (O_2800,N_29816,N_29731);
nand UO_2801 (O_2801,N_29889,N_29907);
nor UO_2802 (O_2802,N_29856,N_29466);
and UO_2803 (O_2803,N_29722,N_29696);
and UO_2804 (O_2804,N_29713,N_29813);
and UO_2805 (O_2805,N_29632,N_29933);
or UO_2806 (O_2806,N_29887,N_29979);
nor UO_2807 (O_2807,N_29803,N_29896);
or UO_2808 (O_2808,N_29729,N_29978);
xor UO_2809 (O_2809,N_29926,N_29596);
xnor UO_2810 (O_2810,N_29698,N_29543);
nand UO_2811 (O_2811,N_29728,N_29570);
nand UO_2812 (O_2812,N_29601,N_29727);
or UO_2813 (O_2813,N_29903,N_29587);
or UO_2814 (O_2814,N_29457,N_29642);
nand UO_2815 (O_2815,N_29829,N_29923);
nand UO_2816 (O_2816,N_29820,N_29729);
nor UO_2817 (O_2817,N_29669,N_29823);
or UO_2818 (O_2818,N_29535,N_29437);
or UO_2819 (O_2819,N_29761,N_29666);
xnor UO_2820 (O_2820,N_29426,N_29652);
or UO_2821 (O_2821,N_29977,N_29568);
or UO_2822 (O_2822,N_29864,N_29634);
and UO_2823 (O_2823,N_29800,N_29573);
and UO_2824 (O_2824,N_29853,N_29427);
and UO_2825 (O_2825,N_29705,N_29826);
nor UO_2826 (O_2826,N_29990,N_29451);
nand UO_2827 (O_2827,N_29514,N_29613);
and UO_2828 (O_2828,N_29887,N_29716);
or UO_2829 (O_2829,N_29855,N_29466);
nand UO_2830 (O_2830,N_29679,N_29658);
and UO_2831 (O_2831,N_29550,N_29771);
nor UO_2832 (O_2832,N_29916,N_29618);
nand UO_2833 (O_2833,N_29810,N_29861);
nand UO_2834 (O_2834,N_29417,N_29683);
or UO_2835 (O_2835,N_29490,N_29644);
or UO_2836 (O_2836,N_29831,N_29915);
nor UO_2837 (O_2837,N_29697,N_29606);
nor UO_2838 (O_2838,N_29510,N_29542);
nand UO_2839 (O_2839,N_29896,N_29857);
nand UO_2840 (O_2840,N_29480,N_29449);
and UO_2841 (O_2841,N_29675,N_29634);
nor UO_2842 (O_2842,N_29996,N_29671);
nand UO_2843 (O_2843,N_29462,N_29556);
or UO_2844 (O_2844,N_29743,N_29852);
nand UO_2845 (O_2845,N_29977,N_29897);
and UO_2846 (O_2846,N_29549,N_29440);
nand UO_2847 (O_2847,N_29779,N_29499);
nor UO_2848 (O_2848,N_29533,N_29934);
and UO_2849 (O_2849,N_29839,N_29521);
and UO_2850 (O_2850,N_29725,N_29751);
and UO_2851 (O_2851,N_29791,N_29511);
or UO_2852 (O_2852,N_29541,N_29612);
or UO_2853 (O_2853,N_29422,N_29435);
nor UO_2854 (O_2854,N_29493,N_29549);
or UO_2855 (O_2855,N_29824,N_29873);
or UO_2856 (O_2856,N_29417,N_29870);
xor UO_2857 (O_2857,N_29459,N_29833);
nand UO_2858 (O_2858,N_29621,N_29921);
xor UO_2859 (O_2859,N_29636,N_29789);
or UO_2860 (O_2860,N_29793,N_29983);
nand UO_2861 (O_2861,N_29782,N_29467);
and UO_2862 (O_2862,N_29840,N_29784);
nor UO_2863 (O_2863,N_29726,N_29672);
nand UO_2864 (O_2864,N_29472,N_29817);
xor UO_2865 (O_2865,N_29778,N_29843);
and UO_2866 (O_2866,N_29487,N_29897);
and UO_2867 (O_2867,N_29840,N_29777);
nand UO_2868 (O_2868,N_29626,N_29848);
or UO_2869 (O_2869,N_29813,N_29487);
or UO_2870 (O_2870,N_29929,N_29772);
nor UO_2871 (O_2871,N_29883,N_29817);
and UO_2872 (O_2872,N_29968,N_29938);
and UO_2873 (O_2873,N_29457,N_29648);
nor UO_2874 (O_2874,N_29421,N_29710);
or UO_2875 (O_2875,N_29791,N_29945);
nor UO_2876 (O_2876,N_29771,N_29432);
nand UO_2877 (O_2877,N_29822,N_29404);
nand UO_2878 (O_2878,N_29651,N_29788);
and UO_2879 (O_2879,N_29958,N_29811);
nor UO_2880 (O_2880,N_29951,N_29666);
and UO_2881 (O_2881,N_29689,N_29585);
nand UO_2882 (O_2882,N_29929,N_29576);
nor UO_2883 (O_2883,N_29922,N_29451);
nand UO_2884 (O_2884,N_29750,N_29972);
or UO_2885 (O_2885,N_29607,N_29830);
and UO_2886 (O_2886,N_29794,N_29637);
or UO_2887 (O_2887,N_29814,N_29625);
xor UO_2888 (O_2888,N_29955,N_29424);
nor UO_2889 (O_2889,N_29836,N_29805);
nor UO_2890 (O_2890,N_29701,N_29695);
nor UO_2891 (O_2891,N_29917,N_29961);
and UO_2892 (O_2892,N_29479,N_29626);
xor UO_2893 (O_2893,N_29615,N_29510);
and UO_2894 (O_2894,N_29612,N_29788);
or UO_2895 (O_2895,N_29476,N_29734);
nor UO_2896 (O_2896,N_29556,N_29906);
nand UO_2897 (O_2897,N_29913,N_29707);
nor UO_2898 (O_2898,N_29916,N_29764);
xor UO_2899 (O_2899,N_29965,N_29698);
xnor UO_2900 (O_2900,N_29565,N_29434);
and UO_2901 (O_2901,N_29865,N_29760);
nor UO_2902 (O_2902,N_29681,N_29712);
and UO_2903 (O_2903,N_29404,N_29733);
xnor UO_2904 (O_2904,N_29690,N_29799);
nor UO_2905 (O_2905,N_29540,N_29597);
or UO_2906 (O_2906,N_29916,N_29874);
nor UO_2907 (O_2907,N_29877,N_29851);
xnor UO_2908 (O_2908,N_29985,N_29798);
nand UO_2909 (O_2909,N_29677,N_29450);
or UO_2910 (O_2910,N_29959,N_29447);
nand UO_2911 (O_2911,N_29438,N_29672);
and UO_2912 (O_2912,N_29438,N_29468);
and UO_2913 (O_2913,N_29477,N_29991);
nor UO_2914 (O_2914,N_29628,N_29771);
nor UO_2915 (O_2915,N_29590,N_29619);
or UO_2916 (O_2916,N_29798,N_29616);
nand UO_2917 (O_2917,N_29969,N_29919);
nand UO_2918 (O_2918,N_29725,N_29978);
nor UO_2919 (O_2919,N_29951,N_29721);
nand UO_2920 (O_2920,N_29523,N_29738);
or UO_2921 (O_2921,N_29519,N_29701);
nor UO_2922 (O_2922,N_29954,N_29610);
xor UO_2923 (O_2923,N_29501,N_29948);
nor UO_2924 (O_2924,N_29482,N_29623);
or UO_2925 (O_2925,N_29899,N_29463);
and UO_2926 (O_2926,N_29938,N_29556);
or UO_2927 (O_2927,N_29930,N_29801);
xnor UO_2928 (O_2928,N_29914,N_29525);
and UO_2929 (O_2929,N_29766,N_29625);
nand UO_2930 (O_2930,N_29448,N_29978);
and UO_2931 (O_2931,N_29520,N_29952);
nor UO_2932 (O_2932,N_29592,N_29777);
and UO_2933 (O_2933,N_29855,N_29856);
or UO_2934 (O_2934,N_29736,N_29730);
xnor UO_2935 (O_2935,N_29649,N_29517);
nor UO_2936 (O_2936,N_29494,N_29843);
nand UO_2937 (O_2937,N_29409,N_29698);
nor UO_2938 (O_2938,N_29923,N_29620);
nand UO_2939 (O_2939,N_29796,N_29478);
or UO_2940 (O_2940,N_29738,N_29534);
xnor UO_2941 (O_2941,N_29446,N_29863);
and UO_2942 (O_2942,N_29643,N_29781);
nand UO_2943 (O_2943,N_29452,N_29947);
or UO_2944 (O_2944,N_29827,N_29921);
nor UO_2945 (O_2945,N_29918,N_29676);
nand UO_2946 (O_2946,N_29770,N_29789);
nor UO_2947 (O_2947,N_29468,N_29761);
nand UO_2948 (O_2948,N_29529,N_29664);
or UO_2949 (O_2949,N_29471,N_29960);
nand UO_2950 (O_2950,N_29611,N_29723);
nor UO_2951 (O_2951,N_29822,N_29767);
nand UO_2952 (O_2952,N_29756,N_29577);
nand UO_2953 (O_2953,N_29685,N_29666);
and UO_2954 (O_2954,N_29523,N_29707);
or UO_2955 (O_2955,N_29573,N_29544);
or UO_2956 (O_2956,N_29961,N_29900);
or UO_2957 (O_2957,N_29603,N_29671);
and UO_2958 (O_2958,N_29922,N_29826);
and UO_2959 (O_2959,N_29850,N_29735);
and UO_2960 (O_2960,N_29581,N_29406);
and UO_2961 (O_2961,N_29527,N_29897);
nand UO_2962 (O_2962,N_29624,N_29854);
and UO_2963 (O_2963,N_29681,N_29515);
xnor UO_2964 (O_2964,N_29552,N_29573);
and UO_2965 (O_2965,N_29955,N_29532);
xor UO_2966 (O_2966,N_29529,N_29616);
xor UO_2967 (O_2967,N_29778,N_29442);
nor UO_2968 (O_2968,N_29967,N_29842);
or UO_2969 (O_2969,N_29555,N_29547);
nor UO_2970 (O_2970,N_29417,N_29832);
xor UO_2971 (O_2971,N_29626,N_29550);
nand UO_2972 (O_2972,N_29990,N_29542);
xnor UO_2973 (O_2973,N_29800,N_29878);
and UO_2974 (O_2974,N_29702,N_29824);
nand UO_2975 (O_2975,N_29906,N_29551);
nand UO_2976 (O_2976,N_29697,N_29695);
xor UO_2977 (O_2977,N_29637,N_29795);
or UO_2978 (O_2978,N_29696,N_29534);
nor UO_2979 (O_2979,N_29439,N_29487);
nor UO_2980 (O_2980,N_29922,N_29805);
nor UO_2981 (O_2981,N_29420,N_29900);
or UO_2982 (O_2982,N_29692,N_29400);
and UO_2983 (O_2983,N_29551,N_29572);
nand UO_2984 (O_2984,N_29509,N_29537);
nor UO_2985 (O_2985,N_29909,N_29953);
nand UO_2986 (O_2986,N_29762,N_29803);
nand UO_2987 (O_2987,N_29839,N_29909);
nor UO_2988 (O_2988,N_29701,N_29822);
nand UO_2989 (O_2989,N_29670,N_29777);
and UO_2990 (O_2990,N_29452,N_29915);
nor UO_2991 (O_2991,N_29714,N_29609);
nor UO_2992 (O_2992,N_29951,N_29782);
nand UO_2993 (O_2993,N_29493,N_29835);
or UO_2994 (O_2994,N_29685,N_29898);
nor UO_2995 (O_2995,N_29719,N_29655);
nor UO_2996 (O_2996,N_29699,N_29459);
xor UO_2997 (O_2997,N_29495,N_29401);
and UO_2998 (O_2998,N_29403,N_29898);
nor UO_2999 (O_2999,N_29862,N_29992);
or UO_3000 (O_3000,N_29806,N_29670);
and UO_3001 (O_3001,N_29743,N_29858);
nand UO_3002 (O_3002,N_29429,N_29745);
nor UO_3003 (O_3003,N_29825,N_29441);
or UO_3004 (O_3004,N_29897,N_29654);
nand UO_3005 (O_3005,N_29653,N_29560);
and UO_3006 (O_3006,N_29853,N_29710);
nor UO_3007 (O_3007,N_29416,N_29993);
nor UO_3008 (O_3008,N_29823,N_29601);
xnor UO_3009 (O_3009,N_29448,N_29590);
and UO_3010 (O_3010,N_29471,N_29909);
nand UO_3011 (O_3011,N_29829,N_29855);
nand UO_3012 (O_3012,N_29772,N_29924);
or UO_3013 (O_3013,N_29929,N_29974);
or UO_3014 (O_3014,N_29859,N_29878);
xnor UO_3015 (O_3015,N_29461,N_29667);
xor UO_3016 (O_3016,N_29641,N_29760);
and UO_3017 (O_3017,N_29527,N_29458);
nor UO_3018 (O_3018,N_29683,N_29673);
nor UO_3019 (O_3019,N_29658,N_29462);
or UO_3020 (O_3020,N_29407,N_29832);
and UO_3021 (O_3021,N_29596,N_29753);
or UO_3022 (O_3022,N_29422,N_29693);
nand UO_3023 (O_3023,N_29575,N_29551);
nor UO_3024 (O_3024,N_29488,N_29482);
nor UO_3025 (O_3025,N_29481,N_29429);
nand UO_3026 (O_3026,N_29957,N_29509);
nand UO_3027 (O_3027,N_29924,N_29708);
and UO_3028 (O_3028,N_29861,N_29524);
or UO_3029 (O_3029,N_29470,N_29649);
nand UO_3030 (O_3030,N_29888,N_29922);
nor UO_3031 (O_3031,N_29643,N_29575);
and UO_3032 (O_3032,N_29774,N_29538);
or UO_3033 (O_3033,N_29855,N_29943);
xnor UO_3034 (O_3034,N_29678,N_29636);
nand UO_3035 (O_3035,N_29732,N_29856);
and UO_3036 (O_3036,N_29425,N_29754);
or UO_3037 (O_3037,N_29583,N_29690);
nand UO_3038 (O_3038,N_29800,N_29735);
nand UO_3039 (O_3039,N_29707,N_29457);
nand UO_3040 (O_3040,N_29601,N_29720);
nand UO_3041 (O_3041,N_29780,N_29617);
and UO_3042 (O_3042,N_29745,N_29701);
and UO_3043 (O_3043,N_29881,N_29631);
nor UO_3044 (O_3044,N_29802,N_29786);
nor UO_3045 (O_3045,N_29834,N_29855);
or UO_3046 (O_3046,N_29868,N_29885);
or UO_3047 (O_3047,N_29534,N_29520);
nand UO_3048 (O_3048,N_29632,N_29544);
nand UO_3049 (O_3049,N_29674,N_29645);
nand UO_3050 (O_3050,N_29738,N_29793);
nand UO_3051 (O_3051,N_29981,N_29543);
nand UO_3052 (O_3052,N_29605,N_29491);
or UO_3053 (O_3053,N_29409,N_29733);
or UO_3054 (O_3054,N_29934,N_29624);
xnor UO_3055 (O_3055,N_29685,N_29810);
and UO_3056 (O_3056,N_29707,N_29922);
xnor UO_3057 (O_3057,N_29816,N_29446);
nand UO_3058 (O_3058,N_29632,N_29676);
and UO_3059 (O_3059,N_29680,N_29822);
xor UO_3060 (O_3060,N_29638,N_29793);
or UO_3061 (O_3061,N_29439,N_29843);
nand UO_3062 (O_3062,N_29532,N_29994);
nor UO_3063 (O_3063,N_29825,N_29560);
nor UO_3064 (O_3064,N_29549,N_29617);
and UO_3065 (O_3065,N_29588,N_29831);
xor UO_3066 (O_3066,N_29831,N_29552);
xnor UO_3067 (O_3067,N_29998,N_29999);
or UO_3068 (O_3068,N_29647,N_29653);
or UO_3069 (O_3069,N_29781,N_29845);
nand UO_3070 (O_3070,N_29881,N_29945);
nand UO_3071 (O_3071,N_29850,N_29676);
nand UO_3072 (O_3072,N_29998,N_29712);
nand UO_3073 (O_3073,N_29455,N_29796);
or UO_3074 (O_3074,N_29564,N_29427);
xor UO_3075 (O_3075,N_29736,N_29572);
and UO_3076 (O_3076,N_29790,N_29915);
or UO_3077 (O_3077,N_29849,N_29909);
or UO_3078 (O_3078,N_29731,N_29609);
and UO_3079 (O_3079,N_29428,N_29808);
nand UO_3080 (O_3080,N_29414,N_29528);
or UO_3081 (O_3081,N_29985,N_29617);
xor UO_3082 (O_3082,N_29948,N_29702);
and UO_3083 (O_3083,N_29552,N_29716);
nand UO_3084 (O_3084,N_29556,N_29916);
nand UO_3085 (O_3085,N_29936,N_29541);
nand UO_3086 (O_3086,N_29951,N_29585);
or UO_3087 (O_3087,N_29878,N_29539);
nor UO_3088 (O_3088,N_29648,N_29886);
or UO_3089 (O_3089,N_29999,N_29797);
nor UO_3090 (O_3090,N_29641,N_29458);
nor UO_3091 (O_3091,N_29569,N_29592);
xor UO_3092 (O_3092,N_29520,N_29501);
nor UO_3093 (O_3093,N_29985,N_29608);
nand UO_3094 (O_3094,N_29914,N_29609);
and UO_3095 (O_3095,N_29612,N_29887);
and UO_3096 (O_3096,N_29701,N_29970);
and UO_3097 (O_3097,N_29861,N_29881);
nand UO_3098 (O_3098,N_29756,N_29533);
or UO_3099 (O_3099,N_29613,N_29491);
or UO_3100 (O_3100,N_29507,N_29791);
or UO_3101 (O_3101,N_29528,N_29670);
nor UO_3102 (O_3102,N_29606,N_29904);
xnor UO_3103 (O_3103,N_29540,N_29470);
nor UO_3104 (O_3104,N_29821,N_29816);
or UO_3105 (O_3105,N_29550,N_29636);
or UO_3106 (O_3106,N_29759,N_29882);
and UO_3107 (O_3107,N_29430,N_29884);
nor UO_3108 (O_3108,N_29687,N_29595);
nand UO_3109 (O_3109,N_29999,N_29631);
or UO_3110 (O_3110,N_29432,N_29709);
nor UO_3111 (O_3111,N_29488,N_29713);
or UO_3112 (O_3112,N_29816,N_29974);
nand UO_3113 (O_3113,N_29409,N_29990);
and UO_3114 (O_3114,N_29849,N_29525);
nor UO_3115 (O_3115,N_29864,N_29503);
nor UO_3116 (O_3116,N_29587,N_29796);
and UO_3117 (O_3117,N_29983,N_29890);
nand UO_3118 (O_3118,N_29820,N_29520);
and UO_3119 (O_3119,N_29923,N_29421);
and UO_3120 (O_3120,N_29424,N_29452);
or UO_3121 (O_3121,N_29881,N_29547);
or UO_3122 (O_3122,N_29931,N_29452);
xnor UO_3123 (O_3123,N_29609,N_29491);
or UO_3124 (O_3124,N_29908,N_29814);
and UO_3125 (O_3125,N_29666,N_29745);
xnor UO_3126 (O_3126,N_29565,N_29572);
and UO_3127 (O_3127,N_29876,N_29872);
nor UO_3128 (O_3128,N_29902,N_29433);
xnor UO_3129 (O_3129,N_29578,N_29610);
nand UO_3130 (O_3130,N_29493,N_29900);
nand UO_3131 (O_3131,N_29706,N_29986);
and UO_3132 (O_3132,N_29893,N_29839);
xnor UO_3133 (O_3133,N_29618,N_29513);
or UO_3134 (O_3134,N_29827,N_29645);
nor UO_3135 (O_3135,N_29927,N_29816);
nand UO_3136 (O_3136,N_29663,N_29978);
nor UO_3137 (O_3137,N_29862,N_29899);
nand UO_3138 (O_3138,N_29433,N_29724);
nor UO_3139 (O_3139,N_29797,N_29517);
nor UO_3140 (O_3140,N_29619,N_29875);
nand UO_3141 (O_3141,N_29581,N_29692);
and UO_3142 (O_3142,N_29755,N_29450);
or UO_3143 (O_3143,N_29954,N_29669);
and UO_3144 (O_3144,N_29579,N_29732);
xor UO_3145 (O_3145,N_29675,N_29770);
xor UO_3146 (O_3146,N_29857,N_29533);
nand UO_3147 (O_3147,N_29877,N_29945);
or UO_3148 (O_3148,N_29646,N_29493);
or UO_3149 (O_3149,N_29693,N_29661);
nor UO_3150 (O_3150,N_29985,N_29996);
nor UO_3151 (O_3151,N_29718,N_29458);
and UO_3152 (O_3152,N_29452,N_29852);
nor UO_3153 (O_3153,N_29490,N_29933);
and UO_3154 (O_3154,N_29532,N_29908);
and UO_3155 (O_3155,N_29694,N_29882);
or UO_3156 (O_3156,N_29457,N_29544);
and UO_3157 (O_3157,N_29804,N_29484);
or UO_3158 (O_3158,N_29761,N_29613);
nand UO_3159 (O_3159,N_29599,N_29415);
nor UO_3160 (O_3160,N_29461,N_29950);
or UO_3161 (O_3161,N_29449,N_29838);
xnor UO_3162 (O_3162,N_29952,N_29869);
or UO_3163 (O_3163,N_29489,N_29558);
nor UO_3164 (O_3164,N_29789,N_29676);
nor UO_3165 (O_3165,N_29441,N_29724);
and UO_3166 (O_3166,N_29888,N_29562);
nand UO_3167 (O_3167,N_29758,N_29435);
nand UO_3168 (O_3168,N_29458,N_29630);
or UO_3169 (O_3169,N_29981,N_29748);
and UO_3170 (O_3170,N_29446,N_29643);
nor UO_3171 (O_3171,N_29965,N_29762);
and UO_3172 (O_3172,N_29955,N_29962);
nor UO_3173 (O_3173,N_29562,N_29400);
nor UO_3174 (O_3174,N_29648,N_29730);
nor UO_3175 (O_3175,N_29629,N_29520);
nor UO_3176 (O_3176,N_29948,N_29503);
nor UO_3177 (O_3177,N_29904,N_29618);
xor UO_3178 (O_3178,N_29826,N_29715);
or UO_3179 (O_3179,N_29773,N_29851);
and UO_3180 (O_3180,N_29937,N_29586);
or UO_3181 (O_3181,N_29590,N_29418);
and UO_3182 (O_3182,N_29518,N_29994);
xor UO_3183 (O_3183,N_29694,N_29684);
nand UO_3184 (O_3184,N_29411,N_29682);
nor UO_3185 (O_3185,N_29623,N_29924);
or UO_3186 (O_3186,N_29943,N_29915);
and UO_3187 (O_3187,N_29931,N_29504);
nand UO_3188 (O_3188,N_29410,N_29516);
and UO_3189 (O_3189,N_29605,N_29583);
nand UO_3190 (O_3190,N_29905,N_29961);
and UO_3191 (O_3191,N_29872,N_29757);
or UO_3192 (O_3192,N_29554,N_29786);
xor UO_3193 (O_3193,N_29762,N_29695);
or UO_3194 (O_3194,N_29860,N_29700);
and UO_3195 (O_3195,N_29997,N_29743);
xor UO_3196 (O_3196,N_29677,N_29901);
nor UO_3197 (O_3197,N_29535,N_29968);
nor UO_3198 (O_3198,N_29997,N_29710);
or UO_3199 (O_3199,N_29941,N_29870);
and UO_3200 (O_3200,N_29497,N_29527);
nor UO_3201 (O_3201,N_29689,N_29591);
or UO_3202 (O_3202,N_29770,N_29806);
nand UO_3203 (O_3203,N_29841,N_29831);
xor UO_3204 (O_3204,N_29666,N_29567);
nand UO_3205 (O_3205,N_29604,N_29456);
or UO_3206 (O_3206,N_29454,N_29599);
and UO_3207 (O_3207,N_29739,N_29832);
nor UO_3208 (O_3208,N_29547,N_29446);
or UO_3209 (O_3209,N_29538,N_29421);
nand UO_3210 (O_3210,N_29903,N_29856);
nor UO_3211 (O_3211,N_29938,N_29455);
or UO_3212 (O_3212,N_29918,N_29967);
nor UO_3213 (O_3213,N_29733,N_29990);
nand UO_3214 (O_3214,N_29733,N_29622);
nand UO_3215 (O_3215,N_29448,N_29793);
and UO_3216 (O_3216,N_29908,N_29681);
nand UO_3217 (O_3217,N_29667,N_29796);
nand UO_3218 (O_3218,N_29425,N_29883);
xor UO_3219 (O_3219,N_29804,N_29462);
or UO_3220 (O_3220,N_29702,N_29774);
nor UO_3221 (O_3221,N_29534,N_29570);
nand UO_3222 (O_3222,N_29723,N_29721);
and UO_3223 (O_3223,N_29637,N_29849);
or UO_3224 (O_3224,N_29903,N_29528);
nor UO_3225 (O_3225,N_29944,N_29646);
or UO_3226 (O_3226,N_29921,N_29715);
or UO_3227 (O_3227,N_29513,N_29449);
or UO_3228 (O_3228,N_29638,N_29854);
and UO_3229 (O_3229,N_29804,N_29517);
or UO_3230 (O_3230,N_29506,N_29496);
or UO_3231 (O_3231,N_29725,N_29444);
nand UO_3232 (O_3232,N_29728,N_29824);
xnor UO_3233 (O_3233,N_29971,N_29895);
xnor UO_3234 (O_3234,N_29932,N_29477);
nand UO_3235 (O_3235,N_29543,N_29785);
xnor UO_3236 (O_3236,N_29815,N_29783);
nor UO_3237 (O_3237,N_29952,N_29425);
or UO_3238 (O_3238,N_29564,N_29524);
nand UO_3239 (O_3239,N_29822,N_29531);
nor UO_3240 (O_3240,N_29571,N_29681);
nor UO_3241 (O_3241,N_29525,N_29918);
nand UO_3242 (O_3242,N_29909,N_29442);
and UO_3243 (O_3243,N_29468,N_29948);
and UO_3244 (O_3244,N_29722,N_29977);
or UO_3245 (O_3245,N_29434,N_29678);
or UO_3246 (O_3246,N_29745,N_29559);
xor UO_3247 (O_3247,N_29592,N_29917);
nand UO_3248 (O_3248,N_29640,N_29768);
xnor UO_3249 (O_3249,N_29958,N_29603);
xor UO_3250 (O_3250,N_29401,N_29590);
nor UO_3251 (O_3251,N_29618,N_29530);
nor UO_3252 (O_3252,N_29819,N_29919);
and UO_3253 (O_3253,N_29476,N_29507);
or UO_3254 (O_3254,N_29730,N_29984);
and UO_3255 (O_3255,N_29816,N_29579);
xor UO_3256 (O_3256,N_29831,N_29574);
nand UO_3257 (O_3257,N_29561,N_29670);
or UO_3258 (O_3258,N_29564,N_29801);
or UO_3259 (O_3259,N_29878,N_29886);
xor UO_3260 (O_3260,N_29939,N_29694);
and UO_3261 (O_3261,N_29754,N_29949);
or UO_3262 (O_3262,N_29542,N_29771);
or UO_3263 (O_3263,N_29516,N_29668);
and UO_3264 (O_3264,N_29819,N_29460);
nor UO_3265 (O_3265,N_29601,N_29422);
or UO_3266 (O_3266,N_29472,N_29851);
or UO_3267 (O_3267,N_29588,N_29845);
nor UO_3268 (O_3268,N_29860,N_29439);
and UO_3269 (O_3269,N_29536,N_29893);
nor UO_3270 (O_3270,N_29964,N_29426);
nand UO_3271 (O_3271,N_29502,N_29407);
nor UO_3272 (O_3272,N_29622,N_29806);
and UO_3273 (O_3273,N_29401,N_29901);
nor UO_3274 (O_3274,N_29822,N_29975);
nor UO_3275 (O_3275,N_29482,N_29680);
and UO_3276 (O_3276,N_29586,N_29932);
nor UO_3277 (O_3277,N_29479,N_29595);
and UO_3278 (O_3278,N_29757,N_29758);
xor UO_3279 (O_3279,N_29979,N_29432);
or UO_3280 (O_3280,N_29451,N_29848);
and UO_3281 (O_3281,N_29641,N_29632);
or UO_3282 (O_3282,N_29800,N_29874);
and UO_3283 (O_3283,N_29792,N_29779);
nand UO_3284 (O_3284,N_29805,N_29637);
or UO_3285 (O_3285,N_29912,N_29986);
or UO_3286 (O_3286,N_29953,N_29797);
xnor UO_3287 (O_3287,N_29841,N_29481);
or UO_3288 (O_3288,N_29661,N_29653);
and UO_3289 (O_3289,N_29497,N_29462);
or UO_3290 (O_3290,N_29665,N_29410);
nand UO_3291 (O_3291,N_29849,N_29843);
and UO_3292 (O_3292,N_29720,N_29508);
and UO_3293 (O_3293,N_29676,N_29589);
and UO_3294 (O_3294,N_29993,N_29497);
and UO_3295 (O_3295,N_29665,N_29409);
nor UO_3296 (O_3296,N_29814,N_29674);
or UO_3297 (O_3297,N_29913,N_29996);
and UO_3298 (O_3298,N_29790,N_29751);
or UO_3299 (O_3299,N_29820,N_29778);
or UO_3300 (O_3300,N_29473,N_29516);
or UO_3301 (O_3301,N_29941,N_29821);
nor UO_3302 (O_3302,N_29858,N_29695);
and UO_3303 (O_3303,N_29703,N_29541);
nor UO_3304 (O_3304,N_29945,N_29898);
nand UO_3305 (O_3305,N_29947,N_29986);
or UO_3306 (O_3306,N_29423,N_29695);
nand UO_3307 (O_3307,N_29589,N_29534);
nand UO_3308 (O_3308,N_29907,N_29745);
and UO_3309 (O_3309,N_29675,N_29636);
xor UO_3310 (O_3310,N_29587,N_29787);
xor UO_3311 (O_3311,N_29924,N_29677);
nand UO_3312 (O_3312,N_29868,N_29554);
and UO_3313 (O_3313,N_29420,N_29773);
nand UO_3314 (O_3314,N_29782,N_29688);
and UO_3315 (O_3315,N_29961,N_29715);
or UO_3316 (O_3316,N_29585,N_29723);
nor UO_3317 (O_3317,N_29488,N_29491);
nand UO_3318 (O_3318,N_29516,N_29737);
nand UO_3319 (O_3319,N_29884,N_29448);
xnor UO_3320 (O_3320,N_29988,N_29743);
nor UO_3321 (O_3321,N_29710,N_29955);
nand UO_3322 (O_3322,N_29489,N_29870);
nor UO_3323 (O_3323,N_29484,N_29741);
xor UO_3324 (O_3324,N_29892,N_29980);
or UO_3325 (O_3325,N_29461,N_29499);
or UO_3326 (O_3326,N_29579,N_29788);
or UO_3327 (O_3327,N_29571,N_29667);
and UO_3328 (O_3328,N_29951,N_29664);
and UO_3329 (O_3329,N_29509,N_29423);
nor UO_3330 (O_3330,N_29564,N_29862);
nand UO_3331 (O_3331,N_29609,N_29465);
and UO_3332 (O_3332,N_29649,N_29625);
nand UO_3333 (O_3333,N_29472,N_29624);
or UO_3334 (O_3334,N_29690,N_29928);
and UO_3335 (O_3335,N_29620,N_29723);
and UO_3336 (O_3336,N_29451,N_29869);
xnor UO_3337 (O_3337,N_29921,N_29561);
nor UO_3338 (O_3338,N_29815,N_29615);
nor UO_3339 (O_3339,N_29852,N_29506);
or UO_3340 (O_3340,N_29903,N_29716);
or UO_3341 (O_3341,N_29924,N_29866);
or UO_3342 (O_3342,N_29807,N_29720);
or UO_3343 (O_3343,N_29911,N_29567);
xor UO_3344 (O_3344,N_29528,N_29863);
nor UO_3345 (O_3345,N_29984,N_29493);
xnor UO_3346 (O_3346,N_29874,N_29681);
xnor UO_3347 (O_3347,N_29505,N_29583);
and UO_3348 (O_3348,N_29431,N_29540);
nand UO_3349 (O_3349,N_29832,N_29505);
nand UO_3350 (O_3350,N_29546,N_29878);
and UO_3351 (O_3351,N_29859,N_29977);
nand UO_3352 (O_3352,N_29794,N_29799);
nand UO_3353 (O_3353,N_29663,N_29727);
and UO_3354 (O_3354,N_29577,N_29579);
nor UO_3355 (O_3355,N_29632,N_29497);
nand UO_3356 (O_3356,N_29946,N_29529);
nand UO_3357 (O_3357,N_29745,N_29522);
or UO_3358 (O_3358,N_29558,N_29502);
nand UO_3359 (O_3359,N_29494,N_29766);
or UO_3360 (O_3360,N_29572,N_29524);
nor UO_3361 (O_3361,N_29735,N_29722);
and UO_3362 (O_3362,N_29681,N_29922);
and UO_3363 (O_3363,N_29799,N_29974);
nor UO_3364 (O_3364,N_29467,N_29653);
and UO_3365 (O_3365,N_29635,N_29987);
and UO_3366 (O_3366,N_29422,N_29547);
and UO_3367 (O_3367,N_29651,N_29516);
nor UO_3368 (O_3368,N_29686,N_29949);
and UO_3369 (O_3369,N_29762,N_29701);
xor UO_3370 (O_3370,N_29549,N_29662);
or UO_3371 (O_3371,N_29849,N_29532);
or UO_3372 (O_3372,N_29679,N_29756);
and UO_3373 (O_3373,N_29969,N_29452);
or UO_3374 (O_3374,N_29521,N_29477);
and UO_3375 (O_3375,N_29841,N_29780);
nand UO_3376 (O_3376,N_29499,N_29552);
and UO_3377 (O_3377,N_29780,N_29543);
or UO_3378 (O_3378,N_29699,N_29472);
and UO_3379 (O_3379,N_29715,N_29524);
nand UO_3380 (O_3380,N_29924,N_29769);
and UO_3381 (O_3381,N_29813,N_29439);
xnor UO_3382 (O_3382,N_29794,N_29577);
and UO_3383 (O_3383,N_29657,N_29697);
nor UO_3384 (O_3384,N_29662,N_29784);
or UO_3385 (O_3385,N_29799,N_29913);
and UO_3386 (O_3386,N_29801,N_29880);
nor UO_3387 (O_3387,N_29773,N_29689);
and UO_3388 (O_3388,N_29436,N_29806);
nor UO_3389 (O_3389,N_29568,N_29825);
nor UO_3390 (O_3390,N_29952,N_29995);
nor UO_3391 (O_3391,N_29774,N_29498);
nand UO_3392 (O_3392,N_29894,N_29733);
nand UO_3393 (O_3393,N_29458,N_29923);
nor UO_3394 (O_3394,N_29998,N_29689);
nor UO_3395 (O_3395,N_29943,N_29969);
nand UO_3396 (O_3396,N_29797,N_29499);
and UO_3397 (O_3397,N_29606,N_29812);
and UO_3398 (O_3398,N_29449,N_29409);
or UO_3399 (O_3399,N_29927,N_29600);
nand UO_3400 (O_3400,N_29954,N_29905);
nand UO_3401 (O_3401,N_29734,N_29516);
nand UO_3402 (O_3402,N_29410,N_29669);
nand UO_3403 (O_3403,N_29863,N_29869);
nor UO_3404 (O_3404,N_29665,N_29923);
or UO_3405 (O_3405,N_29979,N_29858);
xnor UO_3406 (O_3406,N_29465,N_29803);
nor UO_3407 (O_3407,N_29802,N_29494);
nand UO_3408 (O_3408,N_29706,N_29809);
nor UO_3409 (O_3409,N_29792,N_29479);
nor UO_3410 (O_3410,N_29559,N_29861);
or UO_3411 (O_3411,N_29945,N_29912);
nand UO_3412 (O_3412,N_29631,N_29411);
nand UO_3413 (O_3413,N_29479,N_29693);
nor UO_3414 (O_3414,N_29472,N_29986);
nand UO_3415 (O_3415,N_29411,N_29864);
or UO_3416 (O_3416,N_29886,N_29447);
and UO_3417 (O_3417,N_29955,N_29654);
nand UO_3418 (O_3418,N_29679,N_29757);
and UO_3419 (O_3419,N_29590,N_29786);
nand UO_3420 (O_3420,N_29496,N_29992);
nor UO_3421 (O_3421,N_29459,N_29968);
or UO_3422 (O_3422,N_29886,N_29873);
nand UO_3423 (O_3423,N_29612,N_29850);
nand UO_3424 (O_3424,N_29482,N_29835);
or UO_3425 (O_3425,N_29964,N_29676);
nor UO_3426 (O_3426,N_29937,N_29828);
nor UO_3427 (O_3427,N_29527,N_29644);
nand UO_3428 (O_3428,N_29932,N_29850);
xor UO_3429 (O_3429,N_29780,N_29988);
nor UO_3430 (O_3430,N_29634,N_29841);
and UO_3431 (O_3431,N_29763,N_29567);
xor UO_3432 (O_3432,N_29578,N_29700);
nor UO_3433 (O_3433,N_29737,N_29664);
nor UO_3434 (O_3434,N_29842,N_29492);
or UO_3435 (O_3435,N_29701,N_29544);
and UO_3436 (O_3436,N_29934,N_29735);
and UO_3437 (O_3437,N_29413,N_29761);
nor UO_3438 (O_3438,N_29498,N_29753);
or UO_3439 (O_3439,N_29801,N_29887);
nor UO_3440 (O_3440,N_29947,N_29603);
xor UO_3441 (O_3441,N_29506,N_29654);
and UO_3442 (O_3442,N_29828,N_29851);
xnor UO_3443 (O_3443,N_29984,N_29531);
xor UO_3444 (O_3444,N_29805,N_29953);
or UO_3445 (O_3445,N_29473,N_29757);
xnor UO_3446 (O_3446,N_29594,N_29956);
nand UO_3447 (O_3447,N_29745,N_29563);
or UO_3448 (O_3448,N_29866,N_29840);
or UO_3449 (O_3449,N_29462,N_29745);
nor UO_3450 (O_3450,N_29707,N_29486);
or UO_3451 (O_3451,N_29440,N_29558);
or UO_3452 (O_3452,N_29667,N_29490);
nor UO_3453 (O_3453,N_29521,N_29789);
nor UO_3454 (O_3454,N_29412,N_29603);
nand UO_3455 (O_3455,N_29825,N_29945);
nand UO_3456 (O_3456,N_29582,N_29890);
and UO_3457 (O_3457,N_29690,N_29715);
xor UO_3458 (O_3458,N_29803,N_29950);
or UO_3459 (O_3459,N_29889,N_29538);
or UO_3460 (O_3460,N_29434,N_29620);
nand UO_3461 (O_3461,N_29759,N_29949);
nor UO_3462 (O_3462,N_29943,N_29688);
nand UO_3463 (O_3463,N_29742,N_29505);
or UO_3464 (O_3464,N_29722,N_29614);
and UO_3465 (O_3465,N_29483,N_29710);
nor UO_3466 (O_3466,N_29940,N_29530);
or UO_3467 (O_3467,N_29647,N_29495);
or UO_3468 (O_3468,N_29973,N_29498);
and UO_3469 (O_3469,N_29497,N_29772);
and UO_3470 (O_3470,N_29487,N_29847);
nand UO_3471 (O_3471,N_29722,N_29766);
and UO_3472 (O_3472,N_29900,N_29404);
xnor UO_3473 (O_3473,N_29753,N_29884);
or UO_3474 (O_3474,N_29761,N_29663);
nor UO_3475 (O_3475,N_29839,N_29470);
or UO_3476 (O_3476,N_29466,N_29621);
nor UO_3477 (O_3477,N_29594,N_29467);
nor UO_3478 (O_3478,N_29454,N_29438);
or UO_3479 (O_3479,N_29480,N_29541);
and UO_3480 (O_3480,N_29753,N_29984);
xnor UO_3481 (O_3481,N_29411,N_29416);
or UO_3482 (O_3482,N_29745,N_29449);
nand UO_3483 (O_3483,N_29896,N_29619);
or UO_3484 (O_3484,N_29981,N_29719);
nor UO_3485 (O_3485,N_29951,N_29778);
or UO_3486 (O_3486,N_29737,N_29860);
nor UO_3487 (O_3487,N_29974,N_29459);
nand UO_3488 (O_3488,N_29428,N_29809);
and UO_3489 (O_3489,N_29508,N_29654);
or UO_3490 (O_3490,N_29685,N_29487);
or UO_3491 (O_3491,N_29413,N_29651);
nor UO_3492 (O_3492,N_29488,N_29431);
xnor UO_3493 (O_3493,N_29903,N_29444);
nand UO_3494 (O_3494,N_29534,N_29740);
or UO_3495 (O_3495,N_29464,N_29479);
nor UO_3496 (O_3496,N_29450,N_29718);
or UO_3497 (O_3497,N_29937,N_29420);
nand UO_3498 (O_3498,N_29593,N_29511);
or UO_3499 (O_3499,N_29781,N_29483);
endmodule