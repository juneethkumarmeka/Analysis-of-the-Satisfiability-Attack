module basic_500_3000_500_6_levels_1xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
or U0 (N_0,In_79,In_467);
nor U1 (N_1,In_478,In_283);
nand U2 (N_2,In_44,In_108);
nand U3 (N_3,In_37,In_155);
and U4 (N_4,In_219,In_414);
nor U5 (N_5,In_50,In_457);
nor U6 (N_6,In_269,In_111);
or U7 (N_7,In_333,In_241);
xnor U8 (N_8,In_82,In_495);
and U9 (N_9,In_254,In_84);
nor U10 (N_10,In_413,In_116);
xnor U11 (N_11,In_90,In_221);
nand U12 (N_12,In_99,In_22);
nand U13 (N_13,In_139,In_443);
nand U14 (N_14,In_253,In_215);
nor U15 (N_15,In_40,In_263);
xor U16 (N_16,In_257,In_119);
nor U17 (N_17,In_249,In_250);
or U18 (N_18,In_173,In_11);
or U19 (N_19,In_49,In_359);
nor U20 (N_20,In_452,In_420);
nor U21 (N_21,In_491,In_304);
or U22 (N_22,In_18,In_123);
and U23 (N_23,In_232,In_193);
or U24 (N_24,In_165,In_252);
and U25 (N_25,In_438,In_83);
and U26 (N_26,In_197,In_318);
nor U27 (N_27,In_421,In_497);
nor U28 (N_28,In_81,In_66);
nand U29 (N_29,In_266,In_207);
nor U30 (N_30,In_374,In_78);
nand U31 (N_31,In_301,In_361);
xor U32 (N_32,In_170,In_213);
nor U33 (N_33,In_483,In_211);
nand U34 (N_34,In_154,In_303);
nor U35 (N_35,In_416,In_292);
or U36 (N_36,In_143,In_187);
or U37 (N_37,In_0,In_490);
nand U38 (N_38,In_175,In_69);
and U39 (N_39,In_429,In_224);
nor U40 (N_40,In_338,In_89);
or U41 (N_41,In_163,In_473);
nor U42 (N_42,In_95,In_86);
or U43 (N_43,In_401,In_470);
nor U44 (N_44,In_279,In_102);
nor U45 (N_45,In_298,In_329);
nor U46 (N_46,In_396,In_212);
nor U47 (N_47,In_291,In_423);
and U48 (N_48,In_267,In_204);
and U49 (N_49,In_88,In_311);
and U50 (N_50,In_237,In_411);
nor U51 (N_51,In_158,In_394);
nor U52 (N_52,In_314,In_129);
and U53 (N_53,In_75,In_475);
nor U54 (N_54,In_272,In_160);
nor U55 (N_55,In_464,In_330);
nand U56 (N_56,In_228,In_476);
or U57 (N_57,In_239,In_182);
nand U58 (N_58,In_342,In_471);
nor U59 (N_59,In_405,In_402);
or U60 (N_60,In_346,In_152);
and U61 (N_61,In_47,In_387);
and U62 (N_62,In_341,In_4);
and U63 (N_63,In_92,In_52);
nand U64 (N_64,In_440,In_373);
nor U65 (N_65,In_313,In_355);
nand U66 (N_66,In_64,In_281);
or U67 (N_67,In_295,In_425);
nand U68 (N_68,In_391,In_100);
and U69 (N_69,In_230,In_348);
nand U70 (N_70,In_337,In_72);
or U71 (N_71,In_290,In_109);
nor U72 (N_72,In_157,In_384);
and U73 (N_73,In_45,In_141);
nor U74 (N_74,In_14,In_179);
and U75 (N_75,In_258,In_225);
or U76 (N_76,In_434,In_181);
or U77 (N_77,In_369,In_243);
and U78 (N_78,In_328,In_6);
and U79 (N_79,In_151,In_125);
nand U80 (N_80,In_455,In_246);
nor U81 (N_81,In_482,In_71);
nand U82 (N_82,In_397,In_13);
nand U83 (N_83,In_188,In_153);
nand U84 (N_84,In_59,In_55);
nor U85 (N_85,In_41,In_262);
and U86 (N_86,In_363,In_68);
and U87 (N_87,In_233,In_8);
or U88 (N_88,In_159,In_323);
and U89 (N_89,In_134,In_302);
and U90 (N_90,In_271,In_85);
or U91 (N_91,In_441,In_210);
nor U92 (N_92,In_354,In_407);
nor U93 (N_93,In_74,In_468);
nor U94 (N_94,In_162,In_378);
or U95 (N_95,In_392,In_260);
and U96 (N_96,In_465,In_280);
or U97 (N_97,In_28,In_347);
and U98 (N_98,In_178,In_317);
nor U99 (N_99,In_353,In_454);
nand U100 (N_100,In_156,In_492);
nor U101 (N_101,In_198,In_493);
nor U102 (N_102,In_240,In_144);
nor U103 (N_103,In_217,In_166);
and U104 (N_104,In_265,In_73);
and U105 (N_105,In_105,In_284);
nand U106 (N_106,In_404,In_51);
and U107 (N_107,In_176,In_344);
or U108 (N_108,In_16,In_360);
and U109 (N_109,In_7,In_499);
or U110 (N_110,In_403,In_481);
nand U111 (N_111,In_278,In_104);
or U112 (N_112,In_136,In_488);
and U113 (N_113,In_444,In_294);
or U114 (N_114,In_222,In_332);
and U115 (N_115,In_371,In_247);
and U116 (N_116,In_458,In_58);
or U117 (N_117,In_277,In_19);
nand U118 (N_118,In_432,In_148);
and U119 (N_119,In_340,In_406);
nor U120 (N_120,In_386,In_375);
or U121 (N_121,In_24,In_435);
or U122 (N_122,In_410,In_31);
nand U123 (N_123,In_103,In_192);
and U124 (N_124,In_286,In_214);
and U125 (N_125,In_57,In_447);
or U126 (N_126,In_107,In_43);
or U127 (N_127,In_255,In_184);
or U128 (N_128,In_362,In_67);
nand U129 (N_129,In_417,In_370);
nand U130 (N_130,In_110,In_489);
nor U131 (N_131,In_10,In_409);
nand U132 (N_132,In_296,In_183);
and U133 (N_133,In_486,In_358);
nor U134 (N_134,In_376,In_439);
and U135 (N_135,In_462,In_149);
or U136 (N_136,In_453,In_431);
or U137 (N_137,In_293,In_124);
or U138 (N_138,In_305,In_244);
and U139 (N_139,In_130,In_216);
nor U140 (N_140,In_32,In_310);
or U141 (N_141,In_274,In_474);
xor U142 (N_142,In_231,In_398);
nor U143 (N_143,In_29,In_379);
and U144 (N_144,In_350,In_117);
nand U145 (N_145,In_199,In_299);
nor U146 (N_146,In_122,In_113);
nand U147 (N_147,In_168,In_128);
and U148 (N_148,In_1,In_325);
nor U149 (N_149,In_200,In_426);
or U150 (N_150,In_3,In_327);
nor U151 (N_151,In_77,In_368);
or U152 (N_152,In_91,In_48);
or U153 (N_153,In_65,In_393);
or U154 (N_154,In_364,In_164);
and U155 (N_155,In_42,In_494);
nand U156 (N_156,In_203,In_308);
nor U157 (N_157,In_261,In_9);
and U158 (N_158,In_140,In_270);
and U159 (N_159,In_285,In_383);
or U160 (N_160,In_142,In_36);
nand U161 (N_161,In_408,In_322);
or U162 (N_162,In_53,In_357);
nor U163 (N_163,In_62,In_196);
nand U164 (N_164,In_23,In_61);
and U165 (N_165,In_147,In_275);
nand U166 (N_166,In_242,In_93);
nor U167 (N_167,In_451,In_132);
nor U168 (N_168,In_177,In_382);
nor U169 (N_169,In_460,In_372);
nor U170 (N_170,In_98,In_380);
xor U171 (N_171,In_76,In_496);
nand U172 (N_172,In_381,In_201);
nor U173 (N_173,In_226,In_498);
nor U174 (N_174,In_238,In_133);
nor U175 (N_175,In_223,In_60);
and U176 (N_176,In_94,In_208);
nand U177 (N_177,In_56,In_87);
nor U178 (N_178,In_436,In_450);
nand U179 (N_179,In_487,In_106);
nor U180 (N_180,In_412,In_194);
and U181 (N_181,In_343,In_264);
nor U182 (N_182,In_39,In_366);
nand U183 (N_183,In_339,In_97);
nand U184 (N_184,In_190,In_389);
nor U185 (N_185,In_399,In_300);
and U186 (N_186,In_126,In_449);
nor U187 (N_187,In_365,In_167);
nor U188 (N_188,In_218,In_114);
nor U189 (N_189,In_477,In_367);
nand U190 (N_190,In_101,In_169);
or U191 (N_191,In_433,In_326);
or U192 (N_192,In_356,In_206);
xnor U193 (N_193,In_479,In_287);
and U194 (N_194,In_485,In_282);
and U195 (N_195,In_120,In_118);
nor U196 (N_196,In_195,In_463);
or U197 (N_197,In_171,In_312);
and U198 (N_198,In_324,In_309);
or U199 (N_199,In_256,In_273);
nand U200 (N_200,In_334,In_186);
nor U201 (N_201,In_459,In_469);
or U202 (N_202,In_227,In_335);
and U203 (N_203,In_202,In_234);
nand U204 (N_204,In_180,In_352);
nand U205 (N_205,In_480,In_437);
nand U206 (N_206,In_388,In_331);
and U207 (N_207,In_54,In_259);
or U208 (N_208,In_5,In_351);
and U209 (N_209,In_424,In_115);
or U210 (N_210,In_427,In_135);
nand U211 (N_211,In_418,In_131);
and U212 (N_212,In_38,In_422);
nand U213 (N_213,In_428,In_336);
nand U214 (N_214,In_289,In_35);
or U215 (N_215,In_191,In_127);
or U216 (N_216,In_172,In_251);
nor U217 (N_217,In_34,In_121);
nand U218 (N_218,In_400,In_80);
nor U219 (N_219,In_138,In_484);
and U220 (N_220,In_315,In_27);
nand U221 (N_221,In_415,In_319);
nand U222 (N_222,In_189,In_112);
and U223 (N_223,In_461,In_390);
or U224 (N_224,In_316,In_321);
xnor U225 (N_225,In_445,In_12);
nand U226 (N_226,In_46,In_26);
or U227 (N_227,In_209,In_466);
nor U228 (N_228,In_472,In_205);
nand U229 (N_229,In_174,In_150);
or U230 (N_230,In_377,In_268);
and U231 (N_231,In_137,In_146);
and U232 (N_232,In_63,In_21);
nand U233 (N_233,In_15,In_145);
or U234 (N_234,In_448,In_442);
and U235 (N_235,In_419,In_288);
and U236 (N_236,In_185,In_17);
and U237 (N_237,In_235,In_349);
and U238 (N_238,In_430,In_307);
or U239 (N_239,In_245,In_229);
nand U240 (N_240,In_25,In_345);
nand U241 (N_241,In_33,In_220);
nand U242 (N_242,In_20,In_30);
or U243 (N_243,In_395,In_248);
nor U244 (N_244,In_96,In_456);
nand U245 (N_245,In_276,In_2);
or U246 (N_246,In_236,In_306);
or U247 (N_247,In_446,In_385);
and U248 (N_248,In_320,In_297);
and U249 (N_249,In_70,In_161);
nand U250 (N_250,In_143,In_98);
or U251 (N_251,In_34,In_137);
or U252 (N_252,In_293,In_363);
and U253 (N_253,In_415,In_38);
and U254 (N_254,In_256,In_223);
or U255 (N_255,In_52,In_367);
nand U256 (N_256,In_486,In_223);
and U257 (N_257,In_443,In_489);
or U258 (N_258,In_194,In_291);
nand U259 (N_259,In_344,In_318);
or U260 (N_260,In_155,In_344);
nand U261 (N_261,In_425,In_448);
nand U262 (N_262,In_457,In_217);
and U263 (N_263,In_148,In_67);
nand U264 (N_264,In_273,In_473);
or U265 (N_265,In_175,In_355);
and U266 (N_266,In_411,In_270);
nand U267 (N_267,In_72,In_136);
or U268 (N_268,In_367,In_384);
and U269 (N_269,In_423,In_345);
nor U270 (N_270,In_58,In_374);
nand U271 (N_271,In_101,In_114);
nor U272 (N_272,In_257,In_207);
nand U273 (N_273,In_483,In_421);
nor U274 (N_274,In_169,In_0);
nand U275 (N_275,In_119,In_354);
and U276 (N_276,In_71,In_301);
nor U277 (N_277,In_420,In_282);
nand U278 (N_278,In_348,In_396);
nand U279 (N_279,In_241,In_250);
nand U280 (N_280,In_177,In_455);
nand U281 (N_281,In_329,In_263);
or U282 (N_282,In_218,In_61);
nor U283 (N_283,In_158,In_449);
or U284 (N_284,In_295,In_343);
or U285 (N_285,In_312,In_7);
nand U286 (N_286,In_140,In_278);
nor U287 (N_287,In_16,In_445);
nand U288 (N_288,In_73,In_387);
and U289 (N_289,In_132,In_475);
and U290 (N_290,In_258,In_315);
or U291 (N_291,In_34,In_204);
or U292 (N_292,In_376,In_174);
or U293 (N_293,In_260,In_245);
and U294 (N_294,In_197,In_484);
and U295 (N_295,In_327,In_124);
and U296 (N_296,In_450,In_428);
or U297 (N_297,In_29,In_415);
nor U298 (N_298,In_109,In_345);
nand U299 (N_299,In_475,In_382);
or U300 (N_300,In_326,In_51);
or U301 (N_301,In_457,In_254);
or U302 (N_302,In_15,In_303);
nand U303 (N_303,In_415,In_264);
and U304 (N_304,In_10,In_231);
or U305 (N_305,In_401,In_295);
and U306 (N_306,In_105,In_249);
nor U307 (N_307,In_476,In_17);
or U308 (N_308,In_300,In_246);
and U309 (N_309,In_125,In_55);
nor U310 (N_310,In_289,In_44);
or U311 (N_311,In_136,In_252);
or U312 (N_312,In_90,In_35);
nor U313 (N_313,In_278,In_16);
nor U314 (N_314,In_317,In_39);
nand U315 (N_315,In_0,In_417);
and U316 (N_316,In_490,In_213);
nor U317 (N_317,In_240,In_105);
or U318 (N_318,In_87,In_352);
nor U319 (N_319,In_289,In_34);
nor U320 (N_320,In_445,In_488);
or U321 (N_321,In_16,In_210);
and U322 (N_322,In_452,In_150);
nand U323 (N_323,In_479,In_360);
and U324 (N_324,In_440,In_96);
and U325 (N_325,In_363,In_132);
nand U326 (N_326,In_421,In_55);
nor U327 (N_327,In_179,In_340);
nor U328 (N_328,In_486,In_35);
nand U329 (N_329,In_462,In_258);
nor U330 (N_330,In_285,In_403);
or U331 (N_331,In_46,In_164);
and U332 (N_332,In_69,In_79);
xnor U333 (N_333,In_99,In_199);
and U334 (N_334,In_422,In_92);
nor U335 (N_335,In_408,In_313);
nand U336 (N_336,In_119,In_190);
nand U337 (N_337,In_354,In_401);
and U338 (N_338,In_272,In_22);
nand U339 (N_339,In_328,In_472);
nand U340 (N_340,In_158,In_402);
and U341 (N_341,In_457,In_370);
nand U342 (N_342,In_336,In_436);
or U343 (N_343,In_32,In_138);
or U344 (N_344,In_216,In_71);
and U345 (N_345,In_41,In_331);
nor U346 (N_346,In_25,In_224);
and U347 (N_347,In_329,In_8);
or U348 (N_348,In_422,In_363);
or U349 (N_349,In_145,In_237);
and U350 (N_350,In_53,In_447);
or U351 (N_351,In_78,In_482);
and U352 (N_352,In_251,In_52);
or U353 (N_353,In_374,In_412);
nor U354 (N_354,In_476,In_73);
nor U355 (N_355,In_115,In_312);
and U356 (N_356,In_143,In_3);
nand U357 (N_357,In_360,In_298);
nor U358 (N_358,In_339,In_174);
nor U359 (N_359,In_233,In_282);
nor U360 (N_360,In_46,In_109);
or U361 (N_361,In_437,In_303);
and U362 (N_362,In_163,In_130);
nor U363 (N_363,In_50,In_33);
nand U364 (N_364,In_329,In_324);
nor U365 (N_365,In_395,In_371);
and U366 (N_366,In_292,In_85);
and U367 (N_367,In_466,In_349);
or U368 (N_368,In_191,In_488);
or U369 (N_369,In_468,In_163);
xor U370 (N_370,In_129,In_194);
nor U371 (N_371,In_127,In_294);
nand U372 (N_372,In_203,In_476);
nand U373 (N_373,In_4,In_396);
nand U374 (N_374,In_420,In_404);
nor U375 (N_375,In_113,In_196);
nor U376 (N_376,In_355,In_60);
nor U377 (N_377,In_240,In_149);
and U378 (N_378,In_345,In_222);
or U379 (N_379,In_203,In_85);
and U380 (N_380,In_5,In_195);
nor U381 (N_381,In_484,In_495);
and U382 (N_382,In_15,In_199);
nor U383 (N_383,In_12,In_119);
or U384 (N_384,In_292,In_168);
nor U385 (N_385,In_402,In_75);
or U386 (N_386,In_304,In_373);
and U387 (N_387,In_282,In_327);
nand U388 (N_388,In_216,In_464);
nand U389 (N_389,In_352,In_409);
nor U390 (N_390,In_30,In_146);
nor U391 (N_391,In_235,In_73);
nand U392 (N_392,In_8,In_243);
nand U393 (N_393,In_48,In_88);
or U394 (N_394,In_13,In_255);
and U395 (N_395,In_188,In_375);
and U396 (N_396,In_5,In_421);
nor U397 (N_397,In_148,In_159);
nand U398 (N_398,In_328,In_212);
and U399 (N_399,In_62,In_220);
and U400 (N_400,In_238,In_45);
nand U401 (N_401,In_193,In_37);
or U402 (N_402,In_49,In_376);
or U403 (N_403,In_217,In_39);
nor U404 (N_404,In_18,In_299);
nor U405 (N_405,In_99,In_35);
nand U406 (N_406,In_475,In_369);
and U407 (N_407,In_358,In_363);
and U408 (N_408,In_204,In_178);
nor U409 (N_409,In_225,In_63);
nand U410 (N_410,In_84,In_158);
or U411 (N_411,In_438,In_278);
nor U412 (N_412,In_124,In_214);
nand U413 (N_413,In_387,In_266);
nor U414 (N_414,In_90,In_130);
nor U415 (N_415,In_330,In_366);
nor U416 (N_416,In_2,In_153);
nand U417 (N_417,In_278,In_233);
nand U418 (N_418,In_295,In_391);
nor U419 (N_419,In_133,In_209);
nand U420 (N_420,In_373,In_329);
and U421 (N_421,In_20,In_129);
and U422 (N_422,In_22,In_37);
and U423 (N_423,In_286,In_183);
nor U424 (N_424,In_148,In_26);
nand U425 (N_425,In_494,In_454);
and U426 (N_426,In_120,In_214);
nor U427 (N_427,In_249,In_148);
and U428 (N_428,In_423,In_201);
and U429 (N_429,In_271,In_368);
nand U430 (N_430,In_302,In_28);
and U431 (N_431,In_469,In_426);
nand U432 (N_432,In_262,In_156);
nand U433 (N_433,In_175,In_109);
and U434 (N_434,In_50,In_445);
nand U435 (N_435,In_495,In_88);
or U436 (N_436,In_101,In_103);
and U437 (N_437,In_373,In_62);
and U438 (N_438,In_104,In_98);
and U439 (N_439,In_433,In_88);
and U440 (N_440,In_482,In_57);
and U441 (N_441,In_462,In_275);
nand U442 (N_442,In_243,In_189);
or U443 (N_443,In_211,In_323);
nand U444 (N_444,In_147,In_281);
nand U445 (N_445,In_498,In_219);
or U446 (N_446,In_496,In_462);
nand U447 (N_447,In_13,In_413);
nor U448 (N_448,In_282,In_410);
and U449 (N_449,In_326,In_353);
nor U450 (N_450,In_257,In_181);
nor U451 (N_451,In_161,In_288);
nand U452 (N_452,In_364,In_436);
nor U453 (N_453,In_414,In_453);
or U454 (N_454,In_452,In_428);
nand U455 (N_455,In_128,In_174);
and U456 (N_456,In_250,In_407);
nand U457 (N_457,In_28,In_383);
nand U458 (N_458,In_194,In_78);
or U459 (N_459,In_234,In_424);
nand U460 (N_460,In_393,In_167);
nor U461 (N_461,In_12,In_473);
or U462 (N_462,In_242,In_29);
nor U463 (N_463,In_146,In_235);
nand U464 (N_464,In_279,In_197);
nor U465 (N_465,In_257,In_40);
nand U466 (N_466,In_356,In_462);
nor U467 (N_467,In_280,In_95);
nor U468 (N_468,In_302,In_253);
or U469 (N_469,In_62,In_206);
or U470 (N_470,In_374,In_246);
and U471 (N_471,In_153,In_302);
or U472 (N_472,In_192,In_464);
or U473 (N_473,In_347,In_21);
or U474 (N_474,In_265,In_290);
nor U475 (N_475,In_218,In_95);
nor U476 (N_476,In_96,In_306);
and U477 (N_477,In_33,In_271);
and U478 (N_478,In_149,In_407);
and U479 (N_479,In_102,In_129);
or U480 (N_480,In_132,In_323);
or U481 (N_481,In_480,In_230);
nand U482 (N_482,In_10,In_374);
nor U483 (N_483,In_459,In_426);
or U484 (N_484,In_341,In_383);
and U485 (N_485,In_380,In_279);
nor U486 (N_486,In_141,In_498);
nor U487 (N_487,In_94,In_135);
nor U488 (N_488,In_23,In_74);
and U489 (N_489,In_384,In_337);
nor U490 (N_490,In_58,In_304);
nand U491 (N_491,In_93,In_26);
and U492 (N_492,In_108,In_380);
and U493 (N_493,In_432,In_301);
nand U494 (N_494,In_293,In_38);
and U495 (N_495,In_58,In_4);
or U496 (N_496,In_267,In_311);
xnor U497 (N_497,In_344,In_225);
nor U498 (N_498,In_302,In_194);
nor U499 (N_499,In_36,In_442);
or U500 (N_500,N_376,N_85);
and U501 (N_501,N_68,N_143);
nand U502 (N_502,N_386,N_388);
or U503 (N_503,N_201,N_95);
nor U504 (N_504,N_403,N_490);
nand U505 (N_505,N_30,N_495);
and U506 (N_506,N_256,N_378);
nor U507 (N_507,N_300,N_374);
and U508 (N_508,N_104,N_191);
and U509 (N_509,N_450,N_250);
nor U510 (N_510,N_213,N_106);
nand U511 (N_511,N_310,N_188);
or U512 (N_512,N_341,N_52);
or U513 (N_513,N_53,N_94);
nand U514 (N_514,N_55,N_211);
nand U515 (N_515,N_416,N_289);
nand U516 (N_516,N_142,N_330);
nor U517 (N_517,N_417,N_286);
nor U518 (N_518,N_379,N_456);
and U519 (N_519,N_327,N_187);
and U520 (N_520,N_414,N_153);
nand U521 (N_521,N_11,N_146);
or U522 (N_522,N_328,N_200);
nand U523 (N_523,N_319,N_465);
nand U524 (N_524,N_151,N_207);
nand U525 (N_525,N_18,N_144);
and U526 (N_526,N_36,N_324);
or U527 (N_527,N_138,N_226);
nor U528 (N_528,N_112,N_359);
nor U529 (N_529,N_62,N_367);
nand U530 (N_530,N_356,N_267);
nand U531 (N_531,N_306,N_409);
and U532 (N_532,N_212,N_473);
or U533 (N_533,N_59,N_202);
nor U534 (N_534,N_440,N_461);
and U535 (N_535,N_186,N_39);
nand U536 (N_536,N_22,N_318);
nor U537 (N_537,N_321,N_363);
or U538 (N_538,N_349,N_469);
nand U539 (N_539,N_154,N_26);
nand U540 (N_540,N_71,N_25);
nor U541 (N_541,N_314,N_257);
or U542 (N_542,N_431,N_271);
or U543 (N_543,N_255,N_315);
nand U544 (N_544,N_459,N_96);
nand U545 (N_545,N_421,N_114);
nand U546 (N_546,N_159,N_79);
nand U547 (N_547,N_84,N_51);
xnor U548 (N_548,N_65,N_441);
and U549 (N_549,N_33,N_467);
nor U550 (N_550,N_357,N_178);
or U551 (N_551,N_122,N_227);
or U552 (N_552,N_451,N_90);
nand U553 (N_553,N_93,N_464);
nand U554 (N_554,N_81,N_82);
nand U555 (N_555,N_17,N_496);
nor U556 (N_556,N_449,N_392);
nor U557 (N_557,N_381,N_393);
nand U558 (N_558,N_167,N_254);
nor U559 (N_559,N_301,N_273);
nor U560 (N_560,N_58,N_194);
or U561 (N_561,N_460,N_48);
nand U562 (N_562,N_360,N_290);
nand U563 (N_563,N_480,N_72);
and U564 (N_564,N_401,N_425);
nand U565 (N_565,N_323,N_325);
or U566 (N_566,N_132,N_492);
nor U567 (N_567,N_408,N_190);
and U568 (N_568,N_279,N_322);
nand U569 (N_569,N_410,N_383);
and U570 (N_570,N_242,N_295);
and U571 (N_571,N_317,N_5);
nor U572 (N_572,N_365,N_377);
or U573 (N_573,N_195,N_110);
or U574 (N_574,N_415,N_162);
or U575 (N_575,N_427,N_37);
and U576 (N_576,N_64,N_373);
or U577 (N_577,N_134,N_193);
nand U578 (N_578,N_40,N_169);
nand U579 (N_579,N_113,N_475);
nor U580 (N_580,N_228,N_312);
or U581 (N_581,N_78,N_168);
or U582 (N_582,N_482,N_351);
and U583 (N_583,N_304,N_494);
nand U584 (N_584,N_176,N_241);
nor U585 (N_585,N_418,N_45);
nor U586 (N_586,N_196,N_185);
nand U587 (N_587,N_223,N_432);
nand U588 (N_588,N_474,N_430);
or U589 (N_589,N_233,N_177);
nand U590 (N_590,N_358,N_265);
nor U591 (N_591,N_152,N_50);
or U592 (N_592,N_471,N_404);
or U593 (N_593,N_136,N_270);
and U594 (N_594,N_102,N_487);
and U595 (N_595,N_15,N_299);
and U596 (N_596,N_197,N_214);
nor U597 (N_597,N_157,N_337);
or U598 (N_598,N_123,N_145);
nor U599 (N_599,N_163,N_345);
nor U600 (N_600,N_115,N_184);
and U601 (N_601,N_209,N_382);
nor U602 (N_602,N_49,N_1);
nor U603 (N_603,N_262,N_420);
nand U604 (N_604,N_246,N_34);
and U605 (N_605,N_275,N_130);
nor U606 (N_606,N_263,N_32);
or U607 (N_607,N_348,N_175);
or U608 (N_608,N_463,N_232);
nor U609 (N_609,N_338,N_125);
nor U610 (N_610,N_428,N_399);
nor U611 (N_611,N_199,N_332);
nor U612 (N_612,N_261,N_334);
nand U613 (N_613,N_483,N_54);
and U614 (N_614,N_274,N_240);
or U615 (N_615,N_479,N_244);
nand U616 (N_616,N_343,N_9);
or U617 (N_617,N_397,N_181);
and U618 (N_618,N_453,N_192);
and U619 (N_619,N_10,N_498);
nand U620 (N_620,N_131,N_83);
and U621 (N_621,N_141,N_251);
nor U622 (N_622,N_385,N_13);
nand U623 (N_623,N_269,N_443);
and U624 (N_624,N_288,N_390);
or U625 (N_625,N_140,N_225);
and U626 (N_626,N_111,N_63);
nand U627 (N_627,N_287,N_444);
and U628 (N_628,N_476,N_423);
nand U629 (N_629,N_245,N_60);
and U630 (N_630,N_331,N_137);
nand U631 (N_631,N_14,N_47);
or U632 (N_632,N_224,N_272);
nor U633 (N_633,N_297,N_88);
or U634 (N_634,N_41,N_98);
or U635 (N_635,N_433,N_165);
or U636 (N_636,N_277,N_481);
or U637 (N_637,N_260,N_326);
nor U638 (N_638,N_66,N_436);
and U639 (N_639,N_252,N_2);
xnor U640 (N_640,N_303,N_160);
nand U641 (N_641,N_283,N_239);
and U642 (N_642,N_400,N_426);
or U643 (N_643,N_222,N_268);
nor U644 (N_644,N_419,N_284);
or U645 (N_645,N_394,N_350);
or U646 (N_646,N_294,N_120);
and U647 (N_647,N_180,N_292);
and U648 (N_648,N_20,N_216);
or U649 (N_649,N_307,N_116);
nor U650 (N_650,N_210,N_109);
and U651 (N_651,N_6,N_352);
and U652 (N_652,N_3,N_305);
nand U653 (N_653,N_155,N_472);
nand U654 (N_654,N_56,N_171);
nor U655 (N_655,N_179,N_445);
nor U656 (N_656,N_121,N_75);
and U657 (N_657,N_221,N_105);
or U658 (N_658,N_434,N_298);
or U659 (N_659,N_347,N_353);
nand U660 (N_660,N_61,N_366);
nor U661 (N_661,N_97,N_135);
or U662 (N_662,N_364,N_354);
and U663 (N_663,N_119,N_296);
or U664 (N_664,N_127,N_340);
or U665 (N_665,N_38,N_69);
nor U666 (N_666,N_398,N_164);
and U667 (N_667,N_489,N_80);
and U668 (N_668,N_203,N_166);
and U669 (N_669,N_107,N_100);
and U670 (N_670,N_174,N_396);
nor U671 (N_671,N_411,N_402);
or U672 (N_672,N_253,N_491);
nor U673 (N_673,N_391,N_124);
and U674 (N_674,N_249,N_258);
and U675 (N_675,N_355,N_435);
nand U676 (N_676,N_466,N_316);
and U677 (N_677,N_139,N_147);
or U678 (N_678,N_219,N_486);
nand U679 (N_679,N_336,N_237);
nor U680 (N_680,N_447,N_329);
nand U681 (N_681,N_372,N_407);
nor U682 (N_682,N_12,N_67);
nor U683 (N_683,N_31,N_198);
and U684 (N_684,N_235,N_468);
and U685 (N_685,N_339,N_276);
nand U686 (N_686,N_344,N_470);
nor U687 (N_687,N_488,N_266);
and U688 (N_688,N_172,N_19);
nand U689 (N_689,N_183,N_234);
nor U690 (N_690,N_293,N_128);
nand U691 (N_691,N_87,N_7);
and U692 (N_692,N_493,N_206);
nand U693 (N_693,N_218,N_362);
nor U694 (N_694,N_92,N_103);
and U695 (N_695,N_4,N_24);
nand U696 (N_696,N_182,N_148);
and U697 (N_697,N_27,N_264);
or U698 (N_698,N_161,N_458);
xnor U699 (N_699,N_446,N_133);
and U700 (N_700,N_497,N_89);
or U701 (N_701,N_230,N_248);
nor U702 (N_702,N_477,N_43);
nand U703 (N_703,N_424,N_76);
and U704 (N_704,N_156,N_108);
and U705 (N_705,N_86,N_77);
nand U706 (N_706,N_346,N_342);
and U707 (N_707,N_380,N_118);
nor U708 (N_708,N_57,N_35);
and U709 (N_709,N_91,N_99);
and U710 (N_710,N_412,N_413);
nor U711 (N_711,N_220,N_208);
nand U712 (N_712,N_454,N_238);
or U713 (N_713,N_117,N_285);
nand U714 (N_714,N_150,N_371);
and U715 (N_715,N_278,N_370);
or U716 (N_716,N_281,N_405);
and U717 (N_717,N_217,N_455);
and U718 (N_718,N_389,N_229);
and U719 (N_719,N_448,N_457);
nand U720 (N_720,N_437,N_499);
or U721 (N_721,N_439,N_243);
or U722 (N_722,N_302,N_231);
or U723 (N_723,N_282,N_368);
nor U724 (N_724,N_387,N_23);
or U725 (N_725,N_173,N_0);
nand U726 (N_726,N_46,N_215);
nand U727 (N_727,N_247,N_259);
and U728 (N_728,N_73,N_452);
nor U729 (N_729,N_126,N_74);
nor U730 (N_730,N_101,N_369);
or U731 (N_731,N_406,N_44);
nor U732 (N_732,N_311,N_28);
nand U733 (N_733,N_375,N_170);
nor U734 (N_734,N_29,N_484);
nor U735 (N_735,N_462,N_205);
nor U736 (N_736,N_313,N_485);
and U737 (N_737,N_149,N_333);
and U738 (N_738,N_422,N_438);
and U739 (N_739,N_478,N_204);
nand U740 (N_740,N_320,N_42);
or U741 (N_741,N_395,N_309);
and U742 (N_742,N_384,N_442);
or U743 (N_743,N_429,N_308);
nand U744 (N_744,N_291,N_70);
nor U745 (N_745,N_361,N_16);
or U746 (N_746,N_280,N_8);
and U747 (N_747,N_21,N_236);
and U748 (N_748,N_189,N_158);
nor U749 (N_749,N_129,N_335);
or U750 (N_750,N_9,N_303);
and U751 (N_751,N_37,N_60);
nor U752 (N_752,N_165,N_73);
nand U753 (N_753,N_15,N_385);
or U754 (N_754,N_474,N_245);
or U755 (N_755,N_111,N_145);
and U756 (N_756,N_375,N_154);
and U757 (N_757,N_259,N_29);
nand U758 (N_758,N_188,N_161);
and U759 (N_759,N_55,N_334);
or U760 (N_760,N_103,N_308);
or U761 (N_761,N_4,N_138);
nand U762 (N_762,N_169,N_95);
and U763 (N_763,N_210,N_265);
and U764 (N_764,N_308,N_324);
or U765 (N_765,N_47,N_182);
or U766 (N_766,N_113,N_81);
or U767 (N_767,N_400,N_448);
nor U768 (N_768,N_16,N_68);
or U769 (N_769,N_372,N_82);
nand U770 (N_770,N_13,N_124);
nand U771 (N_771,N_374,N_439);
nand U772 (N_772,N_166,N_3);
and U773 (N_773,N_87,N_192);
nor U774 (N_774,N_78,N_382);
and U775 (N_775,N_279,N_178);
or U776 (N_776,N_477,N_201);
nor U777 (N_777,N_370,N_0);
nand U778 (N_778,N_397,N_86);
xor U779 (N_779,N_78,N_251);
nand U780 (N_780,N_169,N_383);
nor U781 (N_781,N_80,N_345);
nor U782 (N_782,N_227,N_394);
or U783 (N_783,N_202,N_14);
nand U784 (N_784,N_176,N_299);
xor U785 (N_785,N_376,N_406);
nor U786 (N_786,N_120,N_352);
and U787 (N_787,N_32,N_255);
nor U788 (N_788,N_207,N_275);
nor U789 (N_789,N_364,N_14);
nand U790 (N_790,N_343,N_154);
xnor U791 (N_791,N_489,N_19);
nor U792 (N_792,N_411,N_349);
or U793 (N_793,N_118,N_458);
nand U794 (N_794,N_421,N_383);
or U795 (N_795,N_297,N_39);
nor U796 (N_796,N_195,N_175);
nand U797 (N_797,N_240,N_396);
nand U798 (N_798,N_487,N_417);
nand U799 (N_799,N_152,N_420);
nor U800 (N_800,N_453,N_293);
and U801 (N_801,N_371,N_179);
and U802 (N_802,N_466,N_325);
nor U803 (N_803,N_499,N_336);
and U804 (N_804,N_85,N_185);
and U805 (N_805,N_423,N_24);
nor U806 (N_806,N_245,N_291);
or U807 (N_807,N_366,N_215);
nor U808 (N_808,N_234,N_87);
nor U809 (N_809,N_373,N_269);
nand U810 (N_810,N_498,N_289);
nand U811 (N_811,N_296,N_68);
xor U812 (N_812,N_55,N_222);
nor U813 (N_813,N_274,N_299);
nor U814 (N_814,N_429,N_200);
or U815 (N_815,N_278,N_45);
and U816 (N_816,N_172,N_415);
and U817 (N_817,N_71,N_426);
nor U818 (N_818,N_149,N_0);
nand U819 (N_819,N_441,N_256);
nand U820 (N_820,N_166,N_141);
nor U821 (N_821,N_418,N_460);
and U822 (N_822,N_169,N_131);
and U823 (N_823,N_36,N_422);
nand U824 (N_824,N_85,N_237);
nand U825 (N_825,N_129,N_152);
nand U826 (N_826,N_394,N_211);
xor U827 (N_827,N_487,N_243);
and U828 (N_828,N_238,N_215);
nor U829 (N_829,N_51,N_137);
or U830 (N_830,N_116,N_304);
or U831 (N_831,N_273,N_206);
xnor U832 (N_832,N_340,N_103);
nand U833 (N_833,N_463,N_322);
and U834 (N_834,N_24,N_247);
nand U835 (N_835,N_363,N_269);
and U836 (N_836,N_326,N_31);
nor U837 (N_837,N_257,N_1);
and U838 (N_838,N_308,N_467);
or U839 (N_839,N_9,N_465);
and U840 (N_840,N_93,N_283);
nor U841 (N_841,N_451,N_15);
nand U842 (N_842,N_103,N_394);
and U843 (N_843,N_38,N_297);
nand U844 (N_844,N_51,N_36);
nor U845 (N_845,N_308,N_397);
nor U846 (N_846,N_330,N_6);
or U847 (N_847,N_174,N_52);
nor U848 (N_848,N_384,N_268);
and U849 (N_849,N_372,N_151);
nor U850 (N_850,N_375,N_29);
nand U851 (N_851,N_412,N_75);
nor U852 (N_852,N_47,N_87);
and U853 (N_853,N_456,N_54);
or U854 (N_854,N_156,N_247);
nand U855 (N_855,N_72,N_196);
nand U856 (N_856,N_59,N_167);
nand U857 (N_857,N_270,N_227);
and U858 (N_858,N_221,N_156);
nor U859 (N_859,N_218,N_280);
nor U860 (N_860,N_182,N_188);
or U861 (N_861,N_151,N_39);
or U862 (N_862,N_3,N_148);
or U863 (N_863,N_72,N_438);
and U864 (N_864,N_46,N_306);
nand U865 (N_865,N_476,N_278);
nor U866 (N_866,N_444,N_289);
or U867 (N_867,N_223,N_33);
or U868 (N_868,N_230,N_185);
nand U869 (N_869,N_465,N_402);
xnor U870 (N_870,N_395,N_262);
and U871 (N_871,N_383,N_441);
nand U872 (N_872,N_32,N_289);
nor U873 (N_873,N_67,N_379);
or U874 (N_874,N_200,N_312);
nor U875 (N_875,N_201,N_168);
nand U876 (N_876,N_341,N_258);
nand U877 (N_877,N_173,N_238);
nor U878 (N_878,N_294,N_273);
nand U879 (N_879,N_291,N_372);
or U880 (N_880,N_291,N_338);
nand U881 (N_881,N_464,N_245);
and U882 (N_882,N_59,N_246);
and U883 (N_883,N_362,N_219);
nor U884 (N_884,N_19,N_98);
or U885 (N_885,N_292,N_246);
and U886 (N_886,N_92,N_247);
nor U887 (N_887,N_5,N_312);
nor U888 (N_888,N_240,N_110);
nand U889 (N_889,N_341,N_304);
nor U890 (N_890,N_206,N_53);
nand U891 (N_891,N_76,N_221);
and U892 (N_892,N_129,N_379);
and U893 (N_893,N_391,N_321);
nor U894 (N_894,N_499,N_60);
nor U895 (N_895,N_120,N_2);
or U896 (N_896,N_177,N_72);
nor U897 (N_897,N_232,N_430);
and U898 (N_898,N_98,N_159);
and U899 (N_899,N_241,N_379);
or U900 (N_900,N_478,N_57);
nand U901 (N_901,N_276,N_283);
and U902 (N_902,N_254,N_272);
and U903 (N_903,N_466,N_212);
nor U904 (N_904,N_33,N_190);
and U905 (N_905,N_411,N_403);
and U906 (N_906,N_380,N_253);
nor U907 (N_907,N_153,N_280);
nor U908 (N_908,N_117,N_437);
or U909 (N_909,N_361,N_61);
or U910 (N_910,N_127,N_435);
or U911 (N_911,N_457,N_12);
and U912 (N_912,N_60,N_417);
nor U913 (N_913,N_421,N_273);
nor U914 (N_914,N_103,N_432);
and U915 (N_915,N_303,N_402);
and U916 (N_916,N_347,N_436);
nand U917 (N_917,N_0,N_196);
nor U918 (N_918,N_66,N_13);
nor U919 (N_919,N_254,N_203);
nand U920 (N_920,N_42,N_432);
nor U921 (N_921,N_173,N_222);
or U922 (N_922,N_429,N_146);
nand U923 (N_923,N_75,N_382);
nor U924 (N_924,N_440,N_175);
and U925 (N_925,N_72,N_234);
and U926 (N_926,N_307,N_40);
nand U927 (N_927,N_223,N_408);
or U928 (N_928,N_405,N_4);
nand U929 (N_929,N_323,N_71);
and U930 (N_930,N_145,N_242);
and U931 (N_931,N_486,N_187);
or U932 (N_932,N_207,N_63);
nor U933 (N_933,N_404,N_3);
or U934 (N_934,N_57,N_470);
or U935 (N_935,N_232,N_297);
nand U936 (N_936,N_460,N_233);
nand U937 (N_937,N_245,N_418);
nor U938 (N_938,N_489,N_8);
nor U939 (N_939,N_237,N_170);
nor U940 (N_940,N_13,N_274);
and U941 (N_941,N_368,N_161);
nand U942 (N_942,N_149,N_398);
nor U943 (N_943,N_38,N_113);
or U944 (N_944,N_403,N_26);
nand U945 (N_945,N_331,N_168);
nor U946 (N_946,N_83,N_372);
and U947 (N_947,N_487,N_245);
nand U948 (N_948,N_6,N_2);
or U949 (N_949,N_319,N_416);
and U950 (N_950,N_390,N_12);
nor U951 (N_951,N_117,N_268);
and U952 (N_952,N_145,N_362);
or U953 (N_953,N_479,N_97);
and U954 (N_954,N_122,N_165);
nand U955 (N_955,N_237,N_293);
xor U956 (N_956,N_11,N_341);
or U957 (N_957,N_458,N_257);
nor U958 (N_958,N_149,N_352);
or U959 (N_959,N_89,N_405);
or U960 (N_960,N_481,N_168);
nand U961 (N_961,N_269,N_205);
nand U962 (N_962,N_44,N_40);
or U963 (N_963,N_495,N_384);
nand U964 (N_964,N_249,N_480);
nor U965 (N_965,N_307,N_12);
nor U966 (N_966,N_60,N_318);
or U967 (N_967,N_7,N_205);
or U968 (N_968,N_97,N_163);
or U969 (N_969,N_8,N_99);
and U970 (N_970,N_497,N_302);
or U971 (N_971,N_416,N_35);
and U972 (N_972,N_339,N_200);
or U973 (N_973,N_74,N_497);
nor U974 (N_974,N_360,N_155);
nor U975 (N_975,N_159,N_86);
nand U976 (N_976,N_489,N_476);
or U977 (N_977,N_459,N_178);
and U978 (N_978,N_417,N_176);
and U979 (N_979,N_298,N_35);
or U980 (N_980,N_30,N_184);
or U981 (N_981,N_267,N_323);
nor U982 (N_982,N_393,N_271);
nand U983 (N_983,N_415,N_37);
nand U984 (N_984,N_457,N_471);
nand U985 (N_985,N_364,N_138);
and U986 (N_986,N_346,N_316);
nor U987 (N_987,N_352,N_35);
nand U988 (N_988,N_480,N_286);
or U989 (N_989,N_440,N_317);
nor U990 (N_990,N_31,N_340);
and U991 (N_991,N_250,N_229);
nand U992 (N_992,N_411,N_260);
nand U993 (N_993,N_114,N_487);
nand U994 (N_994,N_167,N_346);
nand U995 (N_995,N_333,N_343);
and U996 (N_996,N_322,N_268);
nor U997 (N_997,N_392,N_402);
nor U998 (N_998,N_436,N_93);
or U999 (N_999,N_303,N_243);
nand U1000 (N_1000,N_892,N_624);
and U1001 (N_1001,N_837,N_815);
nand U1002 (N_1002,N_974,N_926);
nor U1003 (N_1003,N_557,N_764);
nand U1004 (N_1004,N_893,N_544);
nand U1005 (N_1005,N_676,N_716);
nor U1006 (N_1006,N_987,N_977);
or U1007 (N_1007,N_527,N_959);
nand U1008 (N_1008,N_961,N_573);
or U1009 (N_1009,N_902,N_953);
nor U1010 (N_1010,N_737,N_805);
nor U1011 (N_1011,N_526,N_749);
and U1012 (N_1012,N_535,N_909);
or U1013 (N_1013,N_850,N_963);
nand U1014 (N_1014,N_556,N_598);
nor U1015 (N_1015,N_860,N_966);
and U1016 (N_1016,N_777,N_865);
nor U1017 (N_1017,N_757,N_595);
or U1018 (N_1018,N_947,N_866);
or U1019 (N_1019,N_930,N_710);
and U1020 (N_1020,N_628,N_901);
nor U1021 (N_1021,N_761,N_639);
nor U1022 (N_1022,N_612,N_661);
or U1023 (N_1023,N_677,N_680);
and U1024 (N_1024,N_975,N_611);
nand U1025 (N_1025,N_523,N_877);
nand U1026 (N_1026,N_731,N_811);
or U1027 (N_1027,N_991,N_674);
and U1028 (N_1028,N_871,N_851);
and U1029 (N_1029,N_644,N_888);
and U1030 (N_1030,N_565,N_610);
or U1031 (N_1031,N_776,N_671);
or U1032 (N_1032,N_835,N_620);
nand U1033 (N_1033,N_891,N_516);
nand U1034 (N_1034,N_904,N_906);
xor U1035 (N_1035,N_683,N_684);
nor U1036 (N_1036,N_944,N_838);
or U1037 (N_1037,N_941,N_779);
nand U1038 (N_1038,N_699,N_655);
nand U1039 (N_1039,N_668,N_734);
nor U1040 (N_1040,N_694,N_623);
nand U1041 (N_1041,N_969,N_846);
and U1042 (N_1042,N_994,N_613);
nor U1043 (N_1043,N_663,N_708);
nand U1044 (N_1044,N_736,N_809);
nor U1045 (N_1045,N_758,N_840);
nor U1046 (N_1046,N_604,N_932);
and U1047 (N_1047,N_564,N_895);
nand U1048 (N_1048,N_982,N_649);
or U1049 (N_1049,N_659,N_642);
nand U1050 (N_1050,N_512,N_882);
and U1051 (N_1051,N_621,N_687);
and U1052 (N_1052,N_529,N_563);
and U1053 (N_1053,N_810,N_913);
or U1054 (N_1054,N_946,N_648);
nor U1055 (N_1055,N_894,N_647);
and U1056 (N_1056,N_950,N_999);
nor U1057 (N_1057,N_678,N_675);
nand U1058 (N_1058,N_696,N_897);
nand U1059 (N_1059,N_690,N_606);
or U1060 (N_1060,N_691,N_729);
nor U1061 (N_1061,N_856,N_854);
nand U1062 (N_1062,N_834,N_867);
and U1063 (N_1063,N_603,N_539);
nand U1064 (N_1064,N_706,N_599);
or U1065 (N_1065,N_848,N_520);
nor U1066 (N_1066,N_983,N_839);
nor U1067 (N_1067,N_827,N_664);
or U1068 (N_1068,N_920,N_985);
or U1069 (N_1069,N_938,N_797);
and U1070 (N_1070,N_607,N_861);
and U1071 (N_1071,N_928,N_829);
nand U1072 (N_1072,N_552,N_579);
and U1073 (N_1073,N_568,N_917);
and U1074 (N_1074,N_589,N_770);
or U1075 (N_1075,N_547,N_657);
or U1076 (N_1076,N_862,N_772);
and U1077 (N_1077,N_972,N_955);
or U1078 (N_1078,N_681,N_574);
nor U1079 (N_1079,N_537,N_717);
nor U1080 (N_1080,N_625,N_995);
nand U1081 (N_1081,N_821,N_510);
nor U1082 (N_1082,N_986,N_723);
and U1083 (N_1083,N_722,N_857);
nor U1084 (N_1084,N_788,N_619);
nor U1085 (N_1085,N_633,N_618);
and U1086 (N_1086,N_968,N_883);
nor U1087 (N_1087,N_679,N_908);
nor U1088 (N_1088,N_755,N_685);
or U1089 (N_1089,N_748,N_910);
nor U1090 (N_1090,N_984,N_800);
and U1091 (N_1091,N_713,N_597);
or U1092 (N_1092,N_560,N_582);
and U1093 (N_1093,N_514,N_992);
and U1094 (N_1094,N_616,N_732);
and U1095 (N_1095,N_789,N_584);
or U1096 (N_1096,N_912,N_583);
or U1097 (N_1097,N_585,N_501);
and U1098 (N_1098,N_524,N_981);
and U1099 (N_1099,N_960,N_577);
or U1100 (N_1100,N_773,N_817);
or U1101 (N_1101,N_754,N_769);
nand U1102 (N_1102,N_791,N_872);
and U1103 (N_1103,N_643,N_571);
nand U1104 (N_1104,N_795,N_559);
and U1105 (N_1105,N_843,N_651);
nand U1106 (N_1106,N_958,N_799);
or U1107 (N_1107,N_964,N_592);
nand U1108 (N_1108,N_715,N_640);
nor U1109 (N_1109,N_828,N_790);
nor U1110 (N_1110,N_730,N_899);
and U1111 (N_1111,N_540,N_550);
nand U1112 (N_1112,N_515,N_922);
nand U1113 (N_1113,N_634,N_980);
or U1114 (N_1114,N_554,N_979);
nand U1115 (N_1115,N_575,N_822);
and U1116 (N_1116,N_876,N_753);
nand U1117 (N_1117,N_538,N_553);
or U1118 (N_1118,N_855,N_654);
nor U1119 (N_1119,N_505,N_534);
and U1120 (N_1120,N_508,N_636);
or U1121 (N_1121,N_833,N_667);
or U1122 (N_1122,N_509,N_705);
nor U1123 (N_1123,N_836,N_551);
or U1124 (N_1124,N_884,N_545);
nand U1125 (N_1125,N_590,N_914);
nand U1126 (N_1126,N_825,N_927);
or U1127 (N_1127,N_903,N_741);
nor U1128 (N_1128,N_688,N_507);
nor U1129 (N_1129,N_704,N_924);
nor U1130 (N_1130,N_586,N_763);
nor U1131 (N_1131,N_915,N_660);
nand U1132 (N_1132,N_847,N_572);
nand U1133 (N_1133,N_814,N_631);
nand U1134 (N_1134,N_555,N_881);
or U1135 (N_1135,N_600,N_738);
or U1136 (N_1136,N_739,N_907);
nor U1137 (N_1137,N_558,N_998);
nand U1138 (N_1138,N_541,N_637);
or U1139 (N_1139,N_796,N_638);
nor U1140 (N_1140,N_786,N_531);
and U1141 (N_1141,N_911,N_962);
nand U1142 (N_1142,N_858,N_670);
and U1143 (N_1143,N_601,N_775);
nor U1144 (N_1144,N_561,N_549);
nor U1145 (N_1145,N_948,N_543);
and U1146 (N_1146,N_693,N_521);
and U1147 (N_1147,N_824,N_548);
or U1148 (N_1148,N_780,N_935);
nand U1149 (N_1149,N_996,N_719);
or U1150 (N_1150,N_940,N_650);
or U1151 (N_1151,N_803,N_707);
nor U1152 (N_1152,N_874,N_656);
or U1153 (N_1153,N_673,N_502);
and U1154 (N_1154,N_852,N_669);
nand U1155 (N_1155,N_718,N_886);
nor U1156 (N_1156,N_783,N_952);
nor U1157 (N_1157,N_689,N_967);
or U1158 (N_1158,N_826,N_804);
and U1159 (N_1159,N_890,N_939);
xor U1160 (N_1160,N_711,N_933);
and U1161 (N_1161,N_570,N_845);
nor U1162 (N_1162,N_532,N_614);
nand U1163 (N_1163,N_813,N_744);
nor U1164 (N_1164,N_774,N_931);
and U1165 (N_1165,N_989,N_581);
or U1166 (N_1166,N_949,N_746);
or U1167 (N_1167,N_630,N_576);
or U1168 (N_1168,N_849,N_767);
nor U1169 (N_1169,N_937,N_608);
nor U1170 (N_1170,N_990,N_511);
nand U1171 (N_1171,N_808,N_978);
nor U1172 (N_1172,N_735,N_831);
or U1173 (N_1173,N_816,N_566);
nand U1174 (N_1174,N_880,N_602);
nor U1175 (N_1175,N_806,N_760);
nand U1176 (N_1176,N_528,N_712);
and U1177 (N_1177,N_781,N_609);
and U1178 (N_1178,N_569,N_709);
nand U1179 (N_1179,N_820,N_802);
and U1180 (N_1180,N_943,N_728);
xor U1181 (N_1181,N_759,N_853);
nand U1182 (N_1182,N_580,N_665);
and U1183 (N_1183,N_818,N_518);
and U1184 (N_1184,N_971,N_605);
nor U1185 (N_1185,N_762,N_942);
nand U1186 (N_1186,N_951,N_703);
and U1187 (N_1187,N_792,N_506);
and U1188 (N_1188,N_720,N_727);
nor U1189 (N_1189,N_787,N_921);
and U1190 (N_1190,N_751,N_743);
and U1191 (N_1191,N_626,N_645);
or U1192 (N_1192,N_993,N_658);
nor U1193 (N_1193,N_562,N_503);
nand U1194 (N_1194,N_695,N_887);
nor U1195 (N_1195,N_905,N_819);
or U1196 (N_1196,N_578,N_726);
and U1197 (N_1197,N_798,N_682);
nand U1198 (N_1198,N_697,N_522);
and U1199 (N_1199,N_875,N_698);
and U1200 (N_1200,N_794,N_766);
and U1201 (N_1201,N_747,N_517);
nand U1202 (N_1202,N_666,N_740);
nand U1203 (N_1203,N_929,N_878);
and U1204 (N_1204,N_700,N_635);
or U1205 (N_1205,N_646,N_976);
or U1206 (N_1206,N_869,N_652);
nor U1207 (N_1207,N_627,N_807);
nor U1208 (N_1208,N_784,N_587);
nand U1209 (N_1209,N_889,N_785);
and U1210 (N_1210,N_957,N_970);
nand U1211 (N_1211,N_632,N_988);
nand U1212 (N_1212,N_702,N_801);
nor U1213 (N_1213,N_868,N_859);
or U1214 (N_1214,N_742,N_923);
nand U1215 (N_1215,N_916,N_830);
nor U1216 (N_1216,N_641,N_533);
nand U1217 (N_1217,N_546,N_918);
nand U1218 (N_1218,N_863,N_945);
nand U1219 (N_1219,N_844,N_724);
or U1220 (N_1220,N_782,N_870);
or U1221 (N_1221,N_721,N_997);
or U1222 (N_1222,N_841,N_615);
or U1223 (N_1223,N_965,N_596);
or U1224 (N_1224,N_519,N_530);
and U1225 (N_1225,N_525,N_500);
or U1226 (N_1226,N_653,N_591);
nand U1227 (N_1227,N_536,N_542);
or U1228 (N_1228,N_954,N_745);
nand U1229 (N_1229,N_629,N_714);
and U1230 (N_1230,N_567,N_588);
and U1231 (N_1231,N_832,N_919);
nand U1232 (N_1232,N_973,N_823);
nor U1233 (N_1233,N_622,N_879);
nor U1234 (N_1234,N_617,N_765);
nand U1235 (N_1235,N_686,N_768);
or U1236 (N_1236,N_936,N_771);
nor U1237 (N_1237,N_672,N_593);
nand U1238 (N_1238,N_812,N_885);
and U1239 (N_1239,N_956,N_864);
nand U1240 (N_1240,N_873,N_750);
and U1241 (N_1241,N_594,N_752);
or U1242 (N_1242,N_504,N_662);
or U1243 (N_1243,N_692,N_725);
or U1244 (N_1244,N_793,N_934);
nor U1245 (N_1245,N_898,N_778);
xor U1246 (N_1246,N_842,N_513);
and U1247 (N_1247,N_701,N_733);
nor U1248 (N_1248,N_925,N_900);
nand U1249 (N_1249,N_896,N_756);
or U1250 (N_1250,N_767,N_570);
or U1251 (N_1251,N_848,N_943);
and U1252 (N_1252,N_624,N_750);
nand U1253 (N_1253,N_645,N_975);
nand U1254 (N_1254,N_686,N_763);
and U1255 (N_1255,N_835,N_936);
nor U1256 (N_1256,N_984,N_591);
nand U1257 (N_1257,N_783,N_983);
nor U1258 (N_1258,N_723,N_662);
and U1259 (N_1259,N_591,N_923);
or U1260 (N_1260,N_629,N_578);
nand U1261 (N_1261,N_751,N_944);
nand U1262 (N_1262,N_630,N_963);
xnor U1263 (N_1263,N_568,N_649);
and U1264 (N_1264,N_993,N_613);
nand U1265 (N_1265,N_835,N_547);
nand U1266 (N_1266,N_962,N_604);
nand U1267 (N_1267,N_736,N_600);
and U1268 (N_1268,N_932,N_990);
or U1269 (N_1269,N_813,N_803);
nand U1270 (N_1270,N_945,N_544);
and U1271 (N_1271,N_724,N_748);
nor U1272 (N_1272,N_991,N_882);
and U1273 (N_1273,N_525,N_588);
nand U1274 (N_1274,N_831,N_952);
nor U1275 (N_1275,N_547,N_598);
nand U1276 (N_1276,N_616,N_996);
or U1277 (N_1277,N_897,N_609);
nand U1278 (N_1278,N_857,N_719);
or U1279 (N_1279,N_548,N_862);
or U1280 (N_1280,N_786,N_626);
nand U1281 (N_1281,N_756,N_984);
nor U1282 (N_1282,N_751,N_664);
or U1283 (N_1283,N_508,N_836);
or U1284 (N_1284,N_979,N_721);
or U1285 (N_1285,N_553,N_604);
and U1286 (N_1286,N_881,N_796);
nand U1287 (N_1287,N_871,N_575);
nor U1288 (N_1288,N_835,N_979);
nand U1289 (N_1289,N_710,N_774);
or U1290 (N_1290,N_808,N_940);
nor U1291 (N_1291,N_603,N_587);
nand U1292 (N_1292,N_874,N_732);
nand U1293 (N_1293,N_739,N_546);
nor U1294 (N_1294,N_561,N_864);
nor U1295 (N_1295,N_506,N_710);
nor U1296 (N_1296,N_855,N_718);
nor U1297 (N_1297,N_700,N_925);
nor U1298 (N_1298,N_530,N_566);
nor U1299 (N_1299,N_902,N_641);
or U1300 (N_1300,N_673,N_787);
nor U1301 (N_1301,N_645,N_889);
or U1302 (N_1302,N_624,N_860);
nand U1303 (N_1303,N_787,N_684);
or U1304 (N_1304,N_752,N_617);
or U1305 (N_1305,N_550,N_809);
or U1306 (N_1306,N_988,N_830);
or U1307 (N_1307,N_842,N_729);
nand U1308 (N_1308,N_894,N_906);
and U1309 (N_1309,N_845,N_909);
and U1310 (N_1310,N_650,N_935);
or U1311 (N_1311,N_623,N_870);
nand U1312 (N_1312,N_677,N_838);
nor U1313 (N_1313,N_912,N_642);
and U1314 (N_1314,N_562,N_747);
or U1315 (N_1315,N_882,N_541);
or U1316 (N_1316,N_735,N_926);
or U1317 (N_1317,N_843,N_540);
nand U1318 (N_1318,N_510,N_893);
nand U1319 (N_1319,N_674,N_925);
or U1320 (N_1320,N_737,N_958);
nor U1321 (N_1321,N_840,N_837);
or U1322 (N_1322,N_555,N_891);
nor U1323 (N_1323,N_815,N_868);
or U1324 (N_1324,N_820,N_788);
and U1325 (N_1325,N_583,N_528);
and U1326 (N_1326,N_868,N_938);
nand U1327 (N_1327,N_751,N_641);
nor U1328 (N_1328,N_807,N_753);
or U1329 (N_1329,N_734,N_723);
nand U1330 (N_1330,N_588,N_958);
nand U1331 (N_1331,N_567,N_785);
or U1332 (N_1332,N_743,N_500);
nor U1333 (N_1333,N_519,N_537);
nor U1334 (N_1334,N_632,N_788);
or U1335 (N_1335,N_576,N_961);
nand U1336 (N_1336,N_819,N_686);
nor U1337 (N_1337,N_938,N_818);
and U1338 (N_1338,N_635,N_506);
or U1339 (N_1339,N_602,N_964);
nor U1340 (N_1340,N_878,N_730);
nand U1341 (N_1341,N_853,N_627);
nand U1342 (N_1342,N_863,N_821);
nand U1343 (N_1343,N_678,N_998);
or U1344 (N_1344,N_513,N_679);
nor U1345 (N_1345,N_884,N_983);
and U1346 (N_1346,N_957,N_996);
nor U1347 (N_1347,N_974,N_656);
and U1348 (N_1348,N_557,N_727);
or U1349 (N_1349,N_955,N_907);
or U1350 (N_1350,N_762,N_651);
or U1351 (N_1351,N_705,N_605);
and U1352 (N_1352,N_812,N_754);
or U1353 (N_1353,N_721,N_606);
nand U1354 (N_1354,N_965,N_608);
or U1355 (N_1355,N_747,N_799);
nand U1356 (N_1356,N_995,N_969);
nor U1357 (N_1357,N_549,N_727);
nand U1358 (N_1358,N_852,N_975);
nor U1359 (N_1359,N_851,N_821);
nor U1360 (N_1360,N_521,N_578);
and U1361 (N_1361,N_514,N_889);
nand U1362 (N_1362,N_752,N_976);
nor U1363 (N_1363,N_892,N_802);
and U1364 (N_1364,N_829,N_677);
or U1365 (N_1365,N_967,N_756);
or U1366 (N_1366,N_891,N_577);
nor U1367 (N_1367,N_506,N_933);
or U1368 (N_1368,N_800,N_840);
and U1369 (N_1369,N_868,N_805);
nor U1370 (N_1370,N_981,N_840);
and U1371 (N_1371,N_564,N_752);
nand U1372 (N_1372,N_857,N_838);
and U1373 (N_1373,N_836,N_921);
or U1374 (N_1374,N_772,N_541);
and U1375 (N_1375,N_750,N_786);
nor U1376 (N_1376,N_924,N_756);
and U1377 (N_1377,N_694,N_718);
or U1378 (N_1378,N_749,N_558);
and U1379 (N_1379,N_910,N_684);
xor U1380 (N_1380,N_970,N_578);
nand U1381 (N_1381,N_541,N_949);
nor U1382 (N_1382,N_570,N_717);
or U1383 (N_1383,N_975,N_811);
and U1384 (N_1384,N_964,N_506);
nor U1385 (N_1385,N_991,N_708);
nand U1386 (N_1386,N_662,N_817);
and U1387 (N_1387,N_792,N_820);
nor U1388 (N_1388,N_975,N_710);
and U1389 (N_1389,N_828,N_546);
nor U1390 (N_1390,N_716,N_507);
or U1391 (N_1391,N_699,N_631);
nand U1392 (N_1392,N_648,N_639);
or U1393 (N_1393,N_974,N_612);
nand U1394 (N_1394,N_829,N_681);
nor U1395 (N_1395,N_784,N_942);
nor U1396 (N_1396,N_931,N_624);
and U1397 (N_1397,N_654,N_523);
nand U1398 (N_1398,N_849,N_637);
nand U1399 (N_1399,N_565,N_503);
or U1400 (N_1400,N_669,N_816);
or U1401 (N_1401,N_942,N_979);
or U1402 (N_1402,N_575,N_711);
nand U1403 (N_1403,N_526,N_545);
nor U1404 (N_1404,N_673,N_603);
nor U1405 (N_1405,N_619,N_884);
or U1406 (N_1406,N_946,N_759);
nor U1407 (N_1407,N_505,N_548);
and U1408 (N_1408,N_866,N_998);
nand U1409 (N_1409,N_973,N_811);
nand U1410 (N_1410,N_636,N_773);
and U1411 (N_1411,N_719,N_602);
nand U1412 (N_1412,N_807,N_772);
nor U1413 (N_1413,N_782,N_971);
and U1414 (N_1414,N_849,N_704);
nor U1415 (N_1415,N_626,N_530);
and U1416 (N_1416,N_547,N_689);
and U1417 (N_1417,N_611,N_520);
nand U1418 (N_1418,N_636,N_506);
nor U1419 (N_1419,N_753,N_560);
nor U1420 (N_1420,N_882,N_641);
nor U1421 (N_1421,N_983,N_571);
and U1422 (N_1422,N_800,N_908);
nor U1423 (N_1423,N_873,N_696);
nand U1424 (N_1424,N_627,N_732);
nor U1425 (N_1425,N_608,N_936);
nand U1426 (N_1426,N_921,N_767);
nor U1427 (N_1427,N_985,N_706);
nand U1428 (N_1428,N_834,N_859);
nor U1429 (N_1429,N_891,N_901);
or U1430 (N_1430,N_787,N_719);
nor U1431 (N_1431,N_972,N_740);
or U1432 (N_1432,N_513,N_810);
nand U1433 (N_1433,N_636,N_776);
nand U1434 (N_1434,N_965,N_542);
nor U1435 (N_1435,N_640,N_998);
or U1436 (N_1436,N_870,N_504);
and U1437 (N_1437,N_810,N_743);
or U1438 (N_1438,N_568,N_782);
or U1439 (N_1439,N_593,N_637);
and U1440 (N_1440,N_529,N_984);
nor U1441 (N_1441,N_565,N_669);
nor U1442 (N_1442,N_659,N_829);
and U1443 (N_1443,N_963,N_808);
and U1444 (N_1444,N_969,N_941);
and U1445 (N_1445,N_624,N_728);
nand U1446 (N_1446,N_725,N_738);
nand U1447 (N_1447,N_894,N_951);
nand U1448 (N_1448,N_516,N_609);
and U1449 (N_1449,N_868,N_906);
and U1450 (N_1450,N_647,N_967);
nand U1451 (N_1451,N_898,N_735);
nand U1452 (N_1452,N_789,N_606);
or U1453 (N_1453,N_776,N_895);
and U1454 (N_1454,N_507,N_990);
nor U1455 (N_1455,N_889,N_546);
or U1456 (N_1456,N_937,N_709);
and U1457 (N_1457,N_712,N_947);
nor U1458 (N_1458,N_864,N_632);
or U1459 (N_1459,N_999,N_829);
nand U1460 (N_1460,N_648,N_621);
or U1461 (N_1461,N_939,N_884);
or U1462 (N_1462,N_806,N_769);
or U1463 (N_1463,N_865,N_821);
nor U1464 (N_1464,N_530,N_955);
nor U1465 (N_1465,N_505,N_904);
and U1466 (N_1466,N_870,N_796);
nor U1467 (N_1467,N_668,N_713);
or U1468 (N_1468,N_610,N_975);
nand U1469 (N_1469,N_629,N_786);
and U1470 (N_1470,N_588,N_710);
or U1471 (N_1471,N_772,N_633);
nor U1472 (N_1472,N_564,N_849);
nor U1473 (N_1473,N_962,N_968);
nand U1474 (N_1474,N_968,N_713);
or U1475 (N_1475,N_636,N_672);
nor U1476 (N_1476,N_841,N_984);
nand U1477 (N_1477,N_815,N_866);
or U1478 (N_1478,N_813,N_594);
or U1479 (N_1479,N_611,N_598);
nor U1480 (N_1480,N_524,N_586);
or U1481 (N_1481,N_691,N_895);
and U1482 (N_1482,N_602,N_895);
or U1483 (N_1483,N_708,N_811);
or U1484 (N_1484,N_623,N_602);
nand U1485 (N_1485,N_893,N_775);
nand U1486 (N_1486,N_969,N_624);
or U1487 (N_1487,N_870,N_817);
nor U1488 (N_1488,N_512,N_925);
nor U1489 (N_1489,N_780,N_804);
nor U1490 (N_1490,N_508,N_993);
or U1491 (N_1491,N_534,N_936);
or U1492 (N_1492,N_709,N_676);
nand U1493 (N_1493,N_688,N_745);
and U1494 (N_1494,N_918,N_642);
nand U1495 (N_1495,N_891,N_879);
nor U1496 (N_1496,N_923,N_815);
or U1497 (N_1497,N_992,N_975);
nor U1498 (N_1498,N_694,N_956);
and U1499 (N_1499,N_544,N_999);
or U1500 (N_1500,N_1291,N_1033);
nand U1501 (N_1501,N_1281,N_1353);
or U1502 (N_1502,N_1072,N_1354);
nand U1503 (N_1503,N_1025,N_1468);
nor U1504 (N_1504,N_1492,N_1459);
nor U1505 (N_1505,N_1044,N_1175);
or U1506 (N_1506,N_1446,N_1393);
or U1507 (N_1507,N_1023,N_1293);
and U1508 (N_1508,N_1143,N_1482);
or U1509 (N_1509,N_1242,N_1213);
nor U1510 (N_1510,N_1260,N_1038);
and U1511 (N_1511,N_1100,N_1094);
xor U1512 (N_1512,N_1083,N_1109);
and U1513 (N_1513,N_1326,N_1338);
nor U1514 (N_1514,N_1060,N_1208);
nand U1515 (N_1515,N_1209,N_1379);
or U1516 (N_1516,N_1095,N_1494);
or U1517 (N_1517,N_1120,N_1245);
nand U1518 (N_1518,N_1006,N_1133);
or U1519 (N_1519,N_1188,N_1210);
nor U1520 (N_1520,N_1127,N_1452);
or U1521 (N_1521,N_1128,N_1415);
nand U1522 (N_1522,N_1067,N_1309);
or U1523 (N_1523,N_1007,N_1406);
and U1524 (N_1524,N_1091,N_1102);
nand U1525 (N_1525,N_1434,N_1017);
nand U1526 (N_1526,N_1451,N_1380);
nor U1527 (N_1527,N_1024,N_1126);
nand U1528 (N_1528,N_1179,N_1110);
nand U1529 (N_1529,N_1461,N_1337);
nor U1530 (N_1530,N_1063,N_1262);
and U1531 (N_1531,N_1084,N_1105);
or U1532 (N_1532,N_1243,N_1357);
nand U1533 (N_1533,N_1003,N_1117);
nand U1534 (N_1534,N_1294,N_1162);
and U1535 (N_1535,N_1061,N_1151);
or U1536 (N_1536,N_1051,N_1233);
nor U1537 (N_1537,N_1004,N_1403);
or U1538 (N_1538,N_1153,N_1166);
or U1539 (N_1539,N_1464,N_1029);
nor U1540 (N_1540,N_1185,N_1428);
nor U1541 (N_1541,N_1218,N_1457);
or U1542 (N_1542,N_1320,N_1483);
and U1543 (N_1543,N_1042,N_1054);
nor U1544 (N_1544,N_1323,N_1430);
and U1545 (N_1545,N_1168,N_1057);
nand U1546 (N_1546,N_1077,N_1396);
nor U1547 (N_1547,N_1229,N_1377);
nor U1548 (N_1548,N_1497,N_1289);
nor U1549 (N_1549,N_1138,N_1286);
and U1550 (N_1550,N_1453,N_1288);
and U1551 (N_1551,N_1258,N_1496);
nand U1552 (N_1552,N_1181,N_1404);
nor U1553 (N_1553,N_1370,N_1485);
or U1554 (N_1554,N_1295,N_1488);
nand U1555 (N_1555,N_1019,N_1304);
or U1556 (N_1556,N_1463,N_1340);
nand U1557 (N_1557,N_1270,N_1448);
or U1558 (N_1558,N_1145,N_1424);
nor U1559 (N_1559,N_1387,N_1202);
and U1560 (N_1560,N_1158,N_1071);
nor U1561 (N_1561,N_1196,N_1352);
nor U1562 (N_1562,N_1257,N_1194);
and U1563 (N_1563,N_1252,N_1271);
nor U1564 (N_1564,N_1214,N_1419);
and U1565 (N_1565,N_1455,N_1183);
nor U1566 (N_1566,N_1059,N_1384);
nor U1567 (N_1567,N_1479,N_1174);
nand U1568 (N_1568,N_1278,N_1080);
nand U1569 (N_1569,N_1382,N_1435);
nand U1570 (N_1570,N_1316,N_1325);
nor U1571 (N_1571,N_1097,N_1383);
or U1572 (N_1572,N_1114,N_1355);
xor U1573 (N_1573,N_1324,N_1204);
nand U1574 (N_1574,N_1328,N_1232);
and U1575 (N_1575,N_1108,N_1201);
or U1576 (N_1576,N_1001,N_1123);
nor U1577 (N_1577,N_1119,N_1152);
nand U1578 (N_1578,N_1409,N_1010);
nand U1579 (N_1579,N_1423,N_1172);
nand U1580 (N_1580,N_1200,N_1161);
nor U1581 (N_1581,N_1334,N_1400);
and U1582 (N_1582,N_1312,N_1125);
and U1583 (N_1583,N_1250,N_1111);
nand U1584 (N_1584,N_1347,N_1239);
nand U1585 (N_1585,N_1122,N_1366);
or U1586 (N_1586,N_1171,N_1187);
nand U1587 (N_1587,N_1362,N_1064);
or U1588 (N_1588,N_1360,N_1277);
or U1589 (N_1589,N_1189,N_1197);
nand U1590 (N_1590,N_1165,N_1154);
nand U1591 (N_1591,N_1432,N_1043);
nand U1592 (N_1592,N_1264,N_1163);
or U1593 (N_1593,N_1317,N_1244);
nor U1594 (N_1594,N_1478,N_1235);
nand U1595 (N_1595,N_1037,N_1009);
and U1596 (N_1596,N_1199,N_1306);
nand U1597 (N_1597,N_1206,N_1450);
nand U1598 (N_1598,N_1065,N_1259);
nor U1599 (N_1599,N_1315,N_1443);
or U1600 (N_1600,N_1449,N_1290);
nor U1601 (N_1601,N_1129,N_1481);
nor U1602 (N_1602,N_1429,N_1373);
or U1603 (N_1603,N_1343,N_1364);
or U1604 (N_1604,N_1155,N_1268);
nand U1605 (N_1605,N_1124,N_1253);
nand U1606 (N_1606,N_1300,N_1287);
nor U1607 (N_1607,N_1472,N_1205);
nor U1608 (N_1608,N_1282,N_1191);
nor U1609 (N_1609,N_1134,N_1490);
and U1610 (N_1610,N_1420,N_1305);
nand U1611 (N_1611,N_1195,N_1034);
and U1612 (N_1612,N_1401,N_1027);
and U1613 (N_1613,N_1280,N_1345);
and U1614 (N_1614,N_1180,N_1327);
or U1615 (N_1615,N_1381,N_1351);
nand U1616 (N_1616,N_1186,N_1053);
xor U1617 (N_1617,N_1035,N_1417);
and U1618 (N_1618,N_1056,N_1068);
or U1619 (N_1619,N_1395,N_1426);
and U1620 (N_1620,N_1495,N_1410);
nand U1621 (N_1621,N_1150,N_1149);
nor U1622 (N_1622,N_1005,N_1237);
nor U1623 (N_1623,N_1225,N_1299);
or U1624 (N_1624,N_1474,N_1477);
nor U1625 (N_1625,N_1031,N_1412);
and U1626 (N_1626,N_1444,N_1392);
and U1627 (N_1627,N_1263,N_1062);
and U1628 (N_1628,N_1275,N_1069);
or U1629 (N_1629,N_1096,N_1026);
or U1630 (N_1630,N_1178,N_1020);
nor U1631 (N_1631,N_1389,N_1480);
and U1632 (N_1632,N_1141,N_1462);
or U1633 (N_1633,N_1303,N_1476);
nor U1634 (N_1634,N_1090,N_1422);
nand U1635 (N_1635,N_1081,N_1115);
nand U1636 (N_1636,N_1106,N_1397);
xor U1637 (N_1637,N_1301,N_1248);
nand U1638 (N_1638,N_1283,N_1159);
and U1639 (N_1639,N_1169,N_1398);
nand U1640 (N_1640,N_1346,N_1460);
nand U1641 (N_1641,N_1344,N_1222);
and U1642 (N_1642,N_1269,N_1164);
and U1643 (N_1643,N_1319,N_1399);
and U1644 (N_1644,N_1231,N_1030);
nand U1645 (N_1645,N_1002,N_1086);
and U1646 (N_1646,N_1131,N_1167);
or U1647 (N_1647,N_1285,N_1484);
and U1648 (N_1648,N_1219,N_1296);
or U1649 (N_1649,N_1372,N_1238);
nor U1650 (N_1650,N_1058,N_1411);
nor U1651 (N_1651,N_1032,N_1413);
xor U1652 (N_1652,N_1021,N_1273);
nand U1653 (N_1653,N_1156,N_1491);
nor U1654 (N_1654,N_1227,N_1447);
or U1655 (N_1655,N_1466,N_1331);
nand U1656 (N_1656,N_1028,N_1112);
nand U1657 (N_1657,N_1313,N_1217);
and U1658 (N_1658,N_1458,N_1298);
nand U1659 (N_1659,N_1135,N_1438);
xor U1660 (N_1660,N_1440,N_1335);
nand U1661 (N_1661,N_1104,N_1469);
nor U1662 (N_1662,N_1487,N_1433);
or U1663 (N_1663,N_1241,N_1016);
nor U1664 (N_1664,N_1365,N_1473);
and U1665 (N_1665,N_1101,N_1050);
or U1666 (N_1666,N_1049,N_1394);
nor U1667 (N_1667,N_1246,N_1333);
nand U1668 (N_1668,N_1272,N_1047);
and U1669 (N_1669,N_1216,N_1307);
or U1670 (N_1670,N_1220,N_1203);
and U1671 (N_1671,N_1092,N_1425);
and U1672 (N_1672,N_1274,N_1236);
or U1673 (N_1673,N_1385,N_1022);
nand U1674 (N_1674,N_1427,N_1107);
nand U1675 (N_1675,N_1066,N_1489);
and U1676 (N_1676,N_1160,N_1140);
or U1677 (N_1677,N_1402,N_1329);
or U1678 (N_1678,N_1375,N_1391);
nor U1679 (N_1679,N_1089,N_1261);
nor U1680 (N_1680,N_1118,N_1332);
nor U1681 (N_1681,N_1074,N_1011);
nand U1682 (N_1682,N_1078,N_1190);
or U1683 (N_1683,N_1418,N_1405);
nor U1684 (N_1684,N_1292,N_1040);
or U1685 (N_1685,N_1308,N_1130);
or U1686 (N_1686,N_1465,N_1018);
nor U1687 (N_1687,N_1142,N_1076);
nor U1688 (N_1688,N_1085,N_1079);
or U1689 (N_1689,N_1098,N_1211);
nor U1690 (N_1690,N_1247,N_1358);
nor U1691 (N_1691,N_1265,N_1173);
nor U1692 (N_1692,N_1414,N_1014);
nor U1693 (N_1693,N_1256,N_1249);
nor U1694 (N_1694,N_1371,N_1475);
and U1695 (N_1695,N_1498,N_1055);
nand U1696 (N_1696,N_1039,N_1445);
and U1697 (N_1697,N_1369,N_1048);
nor U1698 (N_1698,N_1228,N_1436);
or U1699 (N_1699,N_1416,N_1349);
nand U1700 (N_1700,N_1284,N_1215);
or U1701 (N_1701,N_1182,N_1013);
nand U1702 (N_1702,N_1439,N_1266);
nand U1703 (N_1703,N_1221,N_1407);
or U1704 (N_1704,N_1431,N_1116);
or U1705 (N_1705,N_1467,N_1255);
nand U1706 (N_1706,N_1052,N_1234);
xnor U1707 (N_1707,N_1192,N_1302);
nand U1708 (N_1708,N_1374,N_1207);
nand U1709 (N_1709,N_1437,N_1359);
and U1710 (N_1710,N_1336,N_1224);
and U1711 (N_1711,N_1486,N_1330);
nor U1712 (N_1712,N_1147,N_1139);
nor U1713 (N_1713,N_1000,N_1240);
nand U1714 (N_1714,N_1388,N_1198);
nand U1715 (N_1715,N_1454,N_1223);
and U1716 (N_1716,N_1442,N_1297);
or U1717 (N_1717,N_1041,N_1251);
or U1718 (N_1718,N_1132,N_1361);
nor U1719 (N_1719,N_1350,N_1144);
or U1720 (N_1720,N_1348,N_1046);
nand U1721 (N_1721,N_1070,N_1441);
nor U1722 (N_1722,N_1367,N_1157);
nor U1723 (N_1723,N_1356,N_1339);
nor U1724 (N_1724,N_1073,N_1036);
nand U1725 (N_1725,N_1082,N_1212);
and U1726 (N_1726,N_1176,N_1177);
nand U1727 (N_1727,N_1408,N_1254);
nor U1728 (N_1728,N_1146,N_1008);
or U1729 (N_1729,N_1421,N_1088);
and U1730 (N_1730,N_1279,N_1015);
or U1731 (N_1731,N_1012,N_1193);
and U1732 (N_1732,N_1321,N_1045);
and U1733 (N_1733,N_1121,N_1311);
or U1734 (N_1734,N_1226,N_1342);
and U1735 (N_1735,N_1170,N_1230);
nand U1736 (N_1736,N_1276,N_1363);
and U1737 (N_1737,N_1137,N_1314);
and U1738 (N_1738,N_1499,N_1113);
and U1739 (N_1739,N_1493,N_1376);
nand U1740 (N_1740,N_1136,N_1368);
nand U1741 (N_1741,N_1093,N_1470);
nor U1742 (N_1742,N_1184,N_1148);
and U1743 (N_1743,N_1318,N_1087);
or U1744 (N_1744,N_1471,N_1341);
or U1745 (N_1745,N_1267,N_1390);
nor U1746 (N_1746,N_1456,N_1103);
and U1747 (N_1747,N_1310,N_1075);
nor U1748 (N_1748,N_1322,N_1386);
nand U1749 (N_1749,N_1378,N_1099);
nor U1750 (N_1750,N_1106,N_1162);
nand U1751 (N_1751,N_1323,N_1355);
nand U1752 (N_1752,N_1373,N_1218);
nor U1753 (N_1753,N_1183,N_1149);
or U1754 (N_1754,N_1454,N_1080);
or U1755 (N_1755,N_1464,N_1459);
nand U1756 (N_1756,N_1178,N_1085);
nand U1757 (N_1757,N_1137,N_1127);
nand U1758 (N_1758,N_1278,N_1455);
or U1759 (N_1759,N_1227,N_1396);
and U1760 (N_1760,N_1196,N_1101);
or U1761 (N_1761,N_1110,N_1116);
nor U1762 (N_1762,N_1127,N_1172);
nand U1763 (N_1763,N_1043,N_1168);
and U1764 (N_1764,N_1056,N_1120);
and U1765 (N_1765,N_1116,N_1445);
and U1766 (N_1766,N_1262,N_1480);
and U1767 (N_1767,N_1040,N_1315);
or U1768 (N_1768,N_1289,N_1376);
and U1769 (N_1769,N_1346,N_1487);
nand U1770 (N_1770,N_1418,N_1078);
nand U1771 (N_1771,N_1132,N_1072);
and U1772 (N_1772,N_1234,N_1226);
nor U1773 (N_1773,N_1474,N_1060);
or U1774 (N_1774,N_1493,N_1490);
or U1775 (N_1775,N_1170,N_1042);
or U1776 (N_1776,N_1371,N_1108);
and U1777 (N_1777,N_1482,N_1122);
or U1778 (N_1778,N_1353,N_1028);
and U1779 (N_1779,N_1244,N_1254);
and U1780 (N_1780,N_1161,N_1244);
or U1781 (N_1781,N_1296,N_1388);
nor U1782 (N_1782,N_1024,N_1415);
and U1783 (N_1783,N_1055,N_1150);
nor U1784 (N_1784,N_1184,N_1337);
and U1785 (N_1785,N_1037,N_1200);
nor U1786 (N_1786,N_1389,N_1418);
nand U1787 (N_1787,N_1054,N_1048);
and U1788 (N_1788,N_1075,N_1497);
nor U1789 (N_1789,N_1009,N_1016);
or U1790 (N_1790,N_1451,N_1155);
nand U1791 (N_1791,N_1444,N_1450);
nand U1792 (N_1792,N_1122,N_1249);
and U1793 (N_1793,N_1411,N_1243);
nand U1794 (N_1794,N_1031,N_1072);
nor U1795 (N_1795,N_1307,N_1380);
and U1796 (N_1796,N_1401,N_1336);
and U1797 (N_1797,N_1040,N_1461);
or U1798 (N_1798,N_1442,N_1429);
or U1799 (N_1799,N_1205,N_1370);
and U1800 (N_1800,N_1102,N_1251);
nand U1801 (N_1801,N_1392,N_1220);
nand U1802 (N_1802,N_1032,N_1109);
or U1803 (N_1803,N_1275,N_1409);
and U1804 (N_1804,N_1126,N_1188);
nand U1805 (N_1805,N_1265,N_1077);
or U1806 (N_1806,N_1182,N_1214);
nand U1807 (N_1807,N_1076,N_1117);
or U1808 (N_1808,N_1235,N_1191);
nand U1809 (N_1809,N_1128,N_1383);
nand U1810 (N_1810,N_1179,N_1408);
nor U1811 (N_1811,N_1124,N_1404);
nor U1812 (N_1812,N_1274,N_1286);
or U1813 (N_1813,N_1369,N_1423);
nor U1814 (N_1814,N_1285,N_1485);
and U1815 (N_1815,N_1447,N_1328);
nand U1816 (N_1816,N_1091,N_1046);
or U1817 (N_1817,N_1435,N_1318);
or U1818 (N_1818,N_1069,N_1225);
or U1819 (N_1819,N_1439,N_1237);
nand U1820 (N_1820,N_1129,N_1190);
or U1821 (N_1821,N_1445,N_1130);
nand U1822 (N_1822,N_1336,N_1118);
nor U1823 (N_1823,N_1009,N_1474);
nor U1824 (N_1824,N_1438,N_1335);
or U1825 (N_1825,N_1251,N_1252);
or U1826 (N_1826,N_1078,N_1479);
and U1827 (N_1827,N_1348,N_1486);
and U1828 (N_1828,N_1161,N_1137);
nor U1829 (N_1829,N_1238,N_1258);
nor U1830 (N_1830,N_1013,N_1259);
or U1831 (N_1831,N_1185,N_1346);
nor U1832 (N_1832,N_1073,N_1242);
nand U1833 (N_1833,N_1101,N_1408);
nand U1834 (N_1834,N_1104,N_1296);
nor U1835 (N_1835,N_1437,N_1236);
nand U1836 (N_1836,N_1295,N_1174);
and U1837 (N_1837,N_1161,N_1012);
and U1838 (N_1838,N_1109,N_1414);
nor U1839 (N_1839,N_1041,N_1094);
and U1840 (N_1840,N_1005,N_1242);
nand U1841 (N_1841,N_1170,N_1246);
and U1842 (N_1842,N_1401,N_1482);
and U1843 (N_1843,N_1097,N_1291);
or U1844 (N_1844,N_1481,N_1336);
nand U1845 (N_1845,N_1431,N_1363);
nand U1846 (N_1846,N_1499,N_1175);
nand U1847 (N_1847,N_1207,N_1462);
and U1848 (N_1848,N_1257,N_1059);
or U1849 (N_1849,N_1149,N_1026);
and U1850 (N_1850,N_1399,N_1465);
and U1851 (N_1851,N_1345,N_1046);
and U1852 (N_1852,N_1016,N_1100);
nand U1853 (N_1853,N_1203,N_1030);
nand U1854 (N_1854,N_1104,N_1459);
nor U1855 (N_1855,N_1100,N_1379);
or U1856 (N_1856,N_1286,N_1300);
nand U1857 (N_1857,N_1427,N_1396);
nand U1858 (N_1858,N_1378,N_1252);
and U1859 (N_1859,N_1415,N_1021);
nor U1860 (N_1860,N_1372,N_1196);
nand U1861 (N_1861,N_1092,N_1048);
and U1862 (N_1862,N_1163,N_1171);
or U1863 (N_1863,N_1408,N_1104);
nor U1864 (N_1864,N_1346,N_1490);
and U1865 (N_1865,N_1416,N_1037);
nor U1866 (N_1866,N_1035,N_1167);
or U1867 (N_1867,N_1295,N_1032);
nor U1868 (N_1868,N_1356,N_1475);
nor U1869 (N_1869,N_1346,N_1228);
and U1870 (N_1870,N_1220,N_1314);
nand U1871 (N_1871,N_1342,N_1275);
nor U1872 (N_1872,N_1221,N_1382);
and U1873 (N_1873,N_1370,N_1484);
and U1874 (N_1874,N_1374,N_1421);
or U1875 (N_1875,N_1168,N_1259);
or U1876 (N_1876,N_1350,N_1197);
nor U1877 (N_1877,N_1080,N_1252);
or U1878 (N_1878,N_1225,N_1046);
nor U1879 (N_1879,N_1030,N_1254);
and U1880 (N_1880,N_1359,N_1136);
or U1881 (N_1881,N_1001,N_1273);
nand U1882 (N_1882,N_1020,N_1123);
or U1883 (N_1883,N_1408,N_1194);
and U1884 (N_1884,N_1386,N_1154);
nor U1885 (N_1885,N_1303,N_1166);
and U1886 (N_1886,N_1209,N_1327);
nand U1887 (N_1887,N_1118,N_1490);
and U1888 (N_1888,N_1189,N_1284);
and U1889 (N_1889,N_1110,N_1321);
nand U1890 (N_1890,N_1016,N_1111);
nand U1891 (N_1891,N_1331,N_1256);
nor U1892 (N_1892,N_1101,N_1372);
nor U1893 (N_1893,N_1054,N_1178);
or U1894 (N_1894,N_1211,N_1256);
nand U1895 (N_1895,N_1003,N_1490);
nor U1896 (N_1896,N_1353,N_1077);
nand U1897 (N_1897,N_1460,N_1258);
xor U1898 (N_1898,N_1014,N_1181);
nand U1899 (N_1899,N_1211,N_1270);
or U1900 (N_1900,N_1027,N_1158);
nand U1901 (N_1901,N_1136,N_1216);
nand U1902 (N_1902,N_1254,N_1057);
or U1903 (N_1903,N_1031,N_1012);
or U1904 (N_1904,N_1138,N_1116);
nor U1905 (N_1905,N_1099,N_1181);
and U1906 (N_1906,N_1156,N_1438);
nor U1907 (N_1907,N_1033,N_1027);
nand U1908 (N_1908,N_1053,N_1326);
nand U1909 (N_1909,N_1461,N_1098);
nand U1910 (N_1910,N_1150,N_1135);
nand U1911 (N_1911,N_1002,N_1362);
or U1912 (N_1912,N_1350,N_1096);
and U1913 (N_1913,N_1096,N_1145);
nor U1914 (N_1914,N_1152,N_1111);
and U1915 (N_1915,N_1007,N_1171);
and U1916 (N_1916,N_1317,N_1210);
and U1917 (N_1917,N_1338,N_1319);
nand U1918 (N_1918,N_1329,N_1303);
or U1919 (N_1919,N_1256,N_1324);
and U1920 (N_1920,N_1463,N_1318);
nand U1921 (N_1921,N_1351,N_1196);
or U1922 (N_1922,N_1196,N_1397);
nand U1923 (N_1923,N_1115,N_1060);
and U1924 (N_1924,N_1471,N_1306);
nor U1925 (N_1925,N_1423,N_1243);
nand U1926 (N_1926,N_1250,N_1124);
xor U1927 (N_1927,N_1375,N_1234);
nand U1928 (N_1928,N_1427,N_1213);
and U1929 (N_1929,N_1066,N_1338);
nor U1930 (N_1930,N_1164,N_1289);
and U1931 (N_1931,N_1095,N_1312);
nor U1932 (N_1932,N_1432,N_1239);
and U1933 (N_1933,N_1403,N_1493);
nor U1934 (N_1934,N_1362,N_1163);
and U1935 (N_1935,N_1174,N_1006);
or U1936 (N_1936,N_1323,N_1043);
nor U1937 (N_1937,N_1097,N_1119);
nand U1938 (N_1938,N_1143,N_1066);
nor U1939 (N_1939,N_1466,N_1164);
and U1940 (N_1940,N_1452,N_1135);
nand U1941 (N_1941,N_1421,N_1063);
nor U1942 (N_1942,N_1230,N_1409);
nor U1943 (N_1943,N_1205,N_1163);
or U1944 (N_1944,N_1417,N_1331);
nand U1945 (N_1945,N_1277,N_1492);
nor U1946 (N_1946,N_1023,N_1252);
nand U1947 (N_1947,N_1295,N_1354);
and U1948 (N_1948,N_1228,N_1432);
and U1949 (N_1949,N_1496,N_1265);
and U1950 (N_1950,N_1095,N_1066);
nand U1951 (N_1951,N_1458,N_1105);
nand U1952 (N_1952,N_1439,N_1389);
nand U1953 (N_1953,N_1398,N_1239);
or U1954 (N_1954,N_1239,N_1134);
or U1955 (N_1955,N_1039,N_1300);
or U1956 (N_1956,N_1188,N_1484);
nand U1957 (N_1957,N_1072,N_1454);
nand U1958 (N_1958,N_1034,N_1099);
nor U1959 (N_1959,N_1486,N_1394);
nand U1960 (N_1960,N_1415,N_1265);
and U1961 (N_1961,N_1480,N_1044);
nor U1962 (N_1962,N_1323,N_1450);
and U1963 (N_1963,N_1404,N_1164);
and U1964 (N_1964,N_1029,N_1207);
or U1965 (N_1965,N_1084,N_1359);
or U1966 (N_1966,N_1463,N_1199);
and U1967 (N_1967,N_1462,N_1220);
nand U1968 (N_1968,N_1460,N_1437);
or U1969 (N_1969,N_1063,N_1328);
nand U1970 (N_1970,N_1380,N_1479);
or U1971 (N_1971,N_1434,N_1197);
nor U1972 (N_1972,N_1300,N_1093);
and U1973 (N_1973,N_1282,N_1262);
nor U1974 (N_1974,N_1212,N_1271);
nand U1975 (N_1975,N_1425,N_1119);
and U1976 (N_1976,N_1041,N_1454);
nand U1977 (N_1977,N_1218,N_1252);
nand U1978 (N_1978,N_1203,N_1135);
and U1979 (N_1979,N_1191,N_1315);
nor U1980 (N_1980,N_1237,N_1354);
and U1981 (N_1981,N_1417,N_1300);
nand U1982 (N_1982,N_1397,N_1034);
and U1983 (N_1983,N_1065,N_1049);
or U1984 (N_1984,N_1284,N_1243);
or U1985 (N_1985,N_1134,N_1095);
and U1986 (N_1986,N_1141,N_1167);
nor U1987 (N_1987,N_1015,N_1370);
and U1988 (N_1988,N_1093,N_1380);
nand U1989 (N_1989,N_1217,N_1141);
nand U1990 (N_1990,N_1306,N_1425);
nand U1991 (N_1991,N_1214,N_1006);
or U1992 (N_1992,N_1410,N_1451);
nor U1993 (N_1993,N_1119,N_1107);
and U1994 (N_1994,N_1155,N_1119);
and U1995 (N_1995,N_1205,N_1317);
or U1996 (N_1996,N_1083,N_1089);
and U1997 (N_1997,N_1141,N_1150);
or U1998 (N_1998,N_1275,N_1416);
nor U1999 (N_1999,N_1468,N_1265);
or U2000 (N_2000,N_1717,N_1895);
nand U2001 (N_2001,N_1552,N_1825);
and U2002 (N_2002,N_1819,N_1760);
nand U2003 (N_2003,N_1912,N_1518);
nor U2004 (N_2004,N_1848,N_1959);
and U2005 (N_2005,N_1777,N_1581);
nand U2006 (N_2006,N_1748,N_1798);
and U2007 (N_2007,N_1619,N_1878);
or U2008 (N_2008,N_1902,N_1697);
nor U2009 (N_2009,N_1663,N_1953);
nor U2010 (N_2010,N_1835,N_1855);
nand U2011 (N_2011,N_1651,N_1683);
nand U2012 (N_2012,N_1719,N_1767);
nor U2013 (N_2013,N_1824,N_1631);
nand U2014 (N_2014,N_1685,N_1979);
and U2015 (N_2015,N_1968,N_1560);
or U2016 (N_2016,N_1638,N_1654);
nand U2017 (N_2017,N_1917,N_1556);
and U2018 (N_2018,N_1984,N_1576);
and U2019 (N_2019,N_1947,N_1675);
or U2020 (N_2020,N_1692,N_1971);
or U2021 (N_2021,N_1589,N_1973);
or U2022 (N_2022,N_1682,N_1528);
or U2023 (N_2023,N_1543,N_1989);
nor U2024 (N_2024,N_1563,N_1826);
nor U2025 (N_2025,N_1665,N_1550);
nand U2026 (N_2026,N_1766,N_1564);
nand U2027 (N_2027,N_1752,N_1694);
and U2028 (N_2028,N_1660,N_1741);
and U2029 (N_2029,N_1929,N_1736);
nor U2030 (N_2030,N_1801,N_1879);
and U2031 (N_2031,N_1785,N_1987);
or U2032 (N_2032,N_1862,N_1504);
nor U2033 (N_2033,N_1779,N_1740);
and U2034 (N_2034,N_1699,N_1964);
nor U2035 (N_2035,N_1679,N_1904);
nand U2036 (N_2036,N_1960,N_1911);
and U2037 (N_2037,N_1820,N_1704);
nand U2038 (N_2038,N_1745,N_1958);
nor U2039 (N_2039,N_1537,N_1611);
and U2040 (N_2040,N_1982,N_1976);
nor U2041 (N_2041,N_1787,N_1930);
nand U2042 (N_2042,N_1540,N_1530);
and U2043 (N_2043,N_1617,N_1937);
nand U2044 (N_2044,N_1952,N_1782);
or U2045 (N_2045,N_1738,N_1807);
and U2046 (N_2046,N_1702,N_1889);
or U2047 (N_2047,N_1843,N_1859);
nand U2048 (N_2048,N_1844,N_1541);
or U2049 (N_2049,N_1673,N_1969);
or U2050 (N_2050,N_1532,N_1938);
or U2051 (N_2051,N_1815,N_1732);
nor U2052 (N_2052,N_1858,N_1579);
nand U2053 (N_2053,N_1840,N_1788);
nand U2054 (N_2054,N_1927,N_1737);
or U2055 (N_2055,N_1972,N_1750);
and U2056 (N_2056,N_1551,N_1547);
and U2057 (N_2057,N_1925,N_1574);
nor U2058 (N_2058,N_1535,N_1950);
and U2059 (N_2059,N_1948,N_1897);
or U2060 (N_2060,N_1691,N_1956);
or U2061 (N_2061,N_1771,N_1890);
or U2062 (N_2062,N_1503,N_1722);
nor U2063 (N_2063,N_1726,N_1507);
nor U2064 (N_2064,N_1666,N_1941);
or U2065 (N_2065,N_1505,N_1981);
nor U2066 (N_2066,N_1733,N_1523);
nand U2067 (N_2067,N_1565,N_1983);
nor U2068 (N_2068,N_1570,N_1659);
nor U2069 (N_2069,N_1729,N_1715);
nand U2070 (N_2070,N_1880,N_1887);
or U2071 (N_2071,N_1914,N_1567);
nand U2072 (N_2072,N_1922,N_1831);
nand U2073 (N_2073,N_1525,N_1545);
nor U2074 (N_2074,N_1793,N_1866);
nand U2075 (N_2075,N_1686,N_1796);
and U2076 (N_2076,N_1841,N_1915);
nand U2077 (N_2077,N_1652,N_1705);
or U2078 (N_2078,N_1778,N_1749);
nand U2079 (N_2079,N_1781,N_1818);
nor U2080 (N_2080,N_1808,N_1830);
nand U2081 (N_2081,N_1951,N_1728);
or U2082 (N_2082,N_1802,N_1690);
and U2083 (N_2083,N_1613,N_1761);
nand U2084 (N_2084,N_1648,N_1508);
nand U2085 (N_2085,N_1626,N_1711);
nand U2086 (N_2086,N_1521,N_1907);
nor U2087 (N_2087,N_1998,N_1513);
nor U2088 (N_2088,N_1562,N_1944);
or U2089 (N_2089,N_1608,N_1763);
and U2090 (N_2090,N_1789,N_1924);
and U2091 (N_2091,N_1901,N_1999);
nor U2092 (N_2092,N_1721,N_1689);
nor U2093 (N_2093,N_1517,N_1881);
nand U2094 (N_2094,N_1587,N_1975);
nand U2095 (N_2095,N_1609,N_1602);
and U2096 (N_2096,N_1616,N_1569);
nor U2097 (N_2097,N_1669,N_1856);
and U2098 (N_2098,N_1643,N_1918);
nor U2099 (N_2099,N_1622,N_1592);
nand U2100 (N_2100,N_1672,N_1603);
and U2101 (N_2101,N_1629,N_1997);
or U2102 (N_2102,N_1853,N_1606);
nand U2103 (N_2103,N_1714,N_1799);
or U2104 (N_2104,N_1939,N_1966);
nor U2105 (N_2105,N_1557,N_1571);
nor U2106 (N_2106,N_1600,N_1764);
and U2107 (N_2107,N_1515,N_1632);
and U2108 (N_2108,N_1842,N_1886);
and U2109 (N_2109,N_1942,N_1935);
nand U2110 (N_2110,N_1809,N_1583);
and U2111 (N_2111,N_1709,N_1712);
nor U2112 (N_2112,N_1865,N_1783);
nand U2113 (N_2113,N_1829,N_1821);
or U2114 (N_2114,N_1575,N_1816);
and U2115 (N_2115,N_1899,N_1586);
nor U2116 (N_2116,N_1769,N_1693);
nand U2117 (N_2117,N_1957,N_1871);
or U2118 (N_2118,N_1710,N_1936);
or U2119 (N_2119,N_1706,N_1870);
nor U2120 (N_2120,N_1839,N_1896);
or U2121 (N_2121,N_1657,N_1772);
nand U2122 (N_2122,N_1684,N_1773);
xor U2123 (N_2123,N_1644,N_1727);
nor U2124 (N_2124,N_1620,N_1755);
nand U2125 (N_2125,N_1633,N_1864);
and U2126 (N_2126,N_1625,N_1618);
nor U2127 (N_2127,N_1582,N_1892);
and U2128 (N_2128,N_1661,N_1790);
nand U2129 (N_2129,N_1640,N_1656);
or U2130 (N_2130,N_1558,N_1992);
nand U2131 (N_2131,N_1877,N_1822);
and U2132 (N_2132,N_1810,N_1642);
or U2133 (N_2133,N_1614,N_1655);
and U2134 (N_2134,N_1650,N_1718);
nand U2135 (N_2135,N_1512,N_1792);
nand U2136 (N_2136,N_1533,N_1529);
and U2137 (N_2137,N_1610,N_1524);
and U2138 (N_2138,N_1599,N_1875);
nor U2139 (N_2139,N_1553,N_1851);
nand U2140 (N_2140,N_1963,N_1544);
nor U2141 (N_2141,N_1874,N_1688);
nand U2142 (N_2142,N_1986,N_1542);
or U2143 (N_2143,N_1676,N_1628);
and U2144 (N_2144,N_1501,N_1817);
nor U2145 (N_2145,N_1857,N_1635);
or U2146 (N_2146,N_1756,N_1703);
nor U2147 (N_2147,N_1903,N_1891);
nor U2148 (N_2148,N_1906,N_1667);
or U2149 (N_2149,N_1630,N_1978);
and U2150 (N_2150,N_1566,N_1647);
and U2151 (N_2151,N_1955,N_1607);
nand U2152 (N_2152,N_1765,N_1724);
or U2153 (N_2153,N_1725,N_1876);
and U2154 (N_2154,N_1716,N_1931);
nand U2155 (N_2155,N_1527,N_1753);
or U2156 (N_2156,N_1572,N_1554);
nor U2157 (N_2157,N_1775,N_1872);
nor U2158 (N_2158,N_1578,N_1649);
nor U2159 (N_2159,N_1923,N_1908);
xor U2160 (N_2160,N_1624,N_1873);
nor U2161 (N_2161,N_1698,N_1921);
nand U2162 (N_2162,N_1744,N_1637);
and U2163 (N_2163,N_1894,N_1510);
nor U2164 (N_2164,N_1597,N_1674);
and U2165 (N_2165,N_1636,N_1701);
and U2166 (N_2166,N_1746,N_1759);
and U2167 (N_2167,N_1993,N_1700);
nand U2168 (N_2168,N_1511,N_1634);
nor U2169 (N_2169,N_1786,N_1627);
or U2170 (N_2170,N_1990,N_1568);
or U2171 (N_2171,N_1834,N_1670);
or U2172 (N_2172,N_1531,N_1730);
nor U2173 (N_2173,N_1645,N_1590);
or U2174 (N_2174,N_1933,N_1754);
or U2175 (N_2175,N_1945,N_1776);
nor U2176 (N_2176,N_1995,N_1814);
nor U2177 (N_2177,N_1584,N_1900);
nor U2178 (N_2178,N_1926,N_1580);
or U2179 (N_2179,N_1967,N_1910);
and U2180 (N_2180,N_1615,N_1561);
and U2181 (N_2181,N_1795,N_1591);
nor U2182 (N_2182,N_1811,N_1852);
and U2183 (N_2183,N_1536,N_1823);
nor U2184 (N_2184,N_1604,N_1598);
or U2185 (N_2185,N_1713,N_1758);
or U2186 (N_2186,N_1885,N_1555);
nor U2187 (N_2187,N_1680,N_1919);
nand U2188 (N_2188,N_1520,N_1803);
and U2189 (N_2189,N_1805,N_1863);
nor U2190 (N_2190,N_1883,N_1977);
nor U2191 (N_2191,N_1707,N_1946);
nand U2192 (N_2192,N_1641,N_1739);
nand U2193 (N_2193,N_1596,N_1743);
nor U2194 (N_2194,N_1949,N_1588);
nand U2195 (N_2195,N_1595,N_1836);
nor U2196 (N_2196,N_1884,N_1671);
nor U2197 (N_2197,N_1846,N_1577);
nor U2198 (N_2198,N_1509,N_1784);
and U2199 (N_2199,N_1849,N_1593);
and U2200 (N_2200,N_1845,N_1800);
nand U2201 (N_2201,N_1548,N_1549);
and U2202 (N_2202,N_1573,N_1687);
or U2203 (N_2203,N_1882,N_1832);
nor U2204 (N_2204,N_1519,N_1988);
nor U2205 (N_2205,N_1954,N_1861);
or U2206 (N_2206,N_1774,N_1888);
nor U2207 (N_2207,N_1623,N_1920);
and U2208 (N_2208,N_1742,N_1898);
and U2209 (N_2209,N_1860,N_1522);
or U2210 (N_2210,N_1678,N_1962);
and U2211 (N_2211,N_1996,N_1500);
nor U2212 (N_2212,N_1601,N_1677);
nand U2213 (N_2213,N_1806,N_1850);
and U2214 (N_2214,N_1664,N_1970);
nand U2215 (N_2215,N_1867,N_1838);
or U2216 (N_2216,N_1893,N_1646);
nand U2217 (N_2217,N_1827,N_1681);
nor U2218 (N_2218,N_1594,N_1934);
nand U2219 (N_2219,N_1723,N_1514);
or U2220 (N_2220,N_1854,N_1980);
nand U2221 (N_2221,N_1943,N_1991);
nor U2222 (N_2222,N_1961,N_1791);
and U2223 (N_2223,N_1668,N_1794);
or U2224 (N_2224,N_1940,N_1869);
or U2225 (N_2225,N_1658,N_1813);
and U2226 (N_2226,N_1502,N_1708);
nor U2227 (N_2227,N_1731,N_1516);
nor U2228 (N_2228,N_1928,N_1735);
or U2229 (N_2229,N_1612,N_1538);
nor U2230 (N_2230,N_1770,N_1762);
nor U2231 (N_2231,N_1605,N_1837);
nand U2232 (N_2232,N_1747,N_1780);
nor U2233 (N_2233,N_1757,N_1812);
nor U2234 (N_2234,N_1828,N_1506);
nor U2235 (N_2235,N_1768,N_1585);
nand U2236 (N_2236,N_1751,N_1994);
or U2237 (N_2237,N_1720,N_1847);
or U2238 (N_2238,N_1833,N_1909);
or U2239 (N_2239,N_1916,N_1534);
or U2240 (N_2240,N_1539,N_1965);
or U2241 (N_2241,N_1734,N_1797);
or U2242 (N_2242,N_1804,N_1559);
nand U2243 (N_2243,N_1913,N_1905);
xnor U2244 (N_2244,N_1653,N_1974);
and U2245 (N_2245,N_1639,N_1695);
or U2246 (N_2246,N_1932,N_1868);
nand U2247 (N_2247,N_1621,N_1985);
and U2248 (N_2248,N_1546,N_1662);
nand U2249 (N_2249,N_1696,N_1526);
nand U2250 (N_2250,N_1727,N_1927);
nor U2251 (N_2251,N_1537,N_1654);
and U2252 (N_2252,N_1847,N_1729);
and U2253 (N_2253,N_1804,N_1682);
nor U2254 (N_2254,N_1923,N_1624);
nand U2255 (N_2255,N_1781,N_1942);
nor U2256 (N_2256,N_1657,N_1619);
nor U2257 (N_2257,N_1656,N_1840);
nand U2258 (N_2258,N_1887,N_1927);
nor U2259 (N_2259,N_1811,N_1613);
nor U2260 (N_2260,N_1812,N_1528);
or U2261 (N_2261,N_1811,N_1597);
or U2262 (N_2262,N_1869,N_1897);
or U2263 (N_2263,N_1688,N_1814);
nor U2264 (N_2264,N_1572,N_1845);
xnor U2265 (N_2265,N_1744,N_1540);
and U2266 (N_2266,N_1772,N_1726);
nor U2267 (N_2267,N_1909,N_1786);
nor U2268 (N_2268,N_1999,N_1688);
nand U2269 (N_2269,N_1500,N_1547);
or U2270 (N_2270,N_1877,N_1835);
nand U2271 (N_2271,N_1611,N_1855);
and U2272 (N_2272,N_1864,N_1887);
and U2273 (N_2273,N_1681,N_1698);
nand U2274 (N_2274,N_1610,N_1553);
or U2275 (N_2275,N_1903,N_1975);
or U2276 (N_2276,N_1673,N_1891);
nand U2277 (N_2277,N_1500,N_1984);
or U2278 (N_2278,N_1792,N_1675);
and U2279 (N_2279,N_1643,N_1748);
and U2280 (N_2280,N_1584,N_1760);
and U2281 (N_2281,N_1660,N_1865);
nor U2282 (N_2282,N_1575,N_1859);
nand U2283 (N_2283,N_1673,N_1524);
nand U2284 (N_2284,N_1936,N_1546);
or U2285 (N_2285,N_1571,N_1788);
nand U2286 (N_2286,N_1786,N_1706);
nand U2287 (N_2287,N_1993,N_1637);
nor U2288 (N_2288,N_1778,N_1723);
and U2289 (N_2289,N_1865,N_1770);
nand U2290 (N_2290,N_1605,N_1629);
nand U2291 (N_2291,N_1882,N_1741);
nand U2292 (N_2292,N_1520,N_1582);
nand U2293 (N_2293,N_1781,N_1767);
nor U2294 (N_2294,N_1857,N_1568);
or U2295 (N_2295,N_1641,N_1534);
nand U2296 (N_2296,N_1850,N_1902);
nand U2297 (N_2297,N_1920,N_1795);
nand U2298 (N_2298,N_1912,N_1955);
and U2299 (N_2299,N_1567,N_1858);
or U2300 (N_2300,N_1600,N_1890);
or U2301 (N_2301,N_1982,N_1569);
and U2302 (N_2302,N_1962,N_1929);
and U2303 (N_2303,N_1670,N_1845);
nor U2304 (N_2304,N_1694,N_1647);
or U2305 (N_2305,N_1750,N_1553);
nand U2306 (N_2306,N_1768,N_1570);
or U2307 (N_2307,N_1854,N_1600);
nor U2308 (N_2308,N_1534,N_1873);
nor U2309 (N_2309,N_1600,N_1621);
or U2310 (N_2310,N_1959,N_1894);
nand U2311 (N_2311,N_1744,N_1960);
nor U2312 (N_2312,N_1901,N_1600);
nand U2313 (N_2313,N_1819,N_1937);
nor U2314 (N_2314,N_1912,N_1570);
nor U2315 (N_2315,N_1820,N_1834);
or U2316 (N_2316,N_1579,N_1991);
nand U2317 (N_2317,N_1779,N_1962);
nand U2318 (N_2318,N_1632,N_1745);
nor U2319 (N_2319,N_1571,N_1629);
nand U2320 (N_2320,N_1816,N_1778);
nand U2321 (N_2321,N_1519,N_1890);
or U2322 (N_2322,N_1847,N_1641);
or U2323 (N_2323,N_1787,N_1580);
nor U2324 (N_2324,N_1547,N_1857);
nor U2325 (N_2325,N_1771,N_1790);
or U2326 (N_2326,N_1658,N_1770);
nand U2327 (N_2327,N_1738,N_1921);
nand U2328 (N_2328,N_1769,N_1973);
and U2329 (N_2329,N_1791,N_1809);
nand U2330 (N_2330,N_1656,N_1518);
or U2331 (N_2331,N_1663,N_1813);
nor U2332 (N_2332,N_1929,N_1607);
or U2333 (N_2333,N_1968,N_1691);
and U2334 (N_2334,N_1903,N_1720);
or U2335 (N_2335,N_1757,N_1539);
nor U2336 (N_2336,N_1687,N_1967);
nand U2337 (N_2337,N_1993,N_1593);
and U2338 (N_2338,N_1733,N_1767);
nand U2339 (N_2339,N_1757,N_1810);
and U2340 (N_2340,N_1961,N_1726);
nand U2341 (N_2341,N_1518,N_1901);
and U2342 (N_2342,N_1558,N_1893);
or U2343 (N_2343,N_1966,N_1548);
and U2344 (N_2344,N_1939,N_1760);
nor U2345 (N_2345,N_1792,N_1694);
or U2346 (N_2346,N_1613,N_1576);
nor U2347 (N_2347,N_1736,N_1544);
nor U2348 (N_2348,N_1530,N_1760);
and U2349 (N_2349,N_1826,N_1600);
or U2350 (N_2350,N_1910,N_1782);
nor U2351 (N_2351,N_1959,N_1803);
nor U2352 (N_2352,N_1522,N_1706);
nor U2353 (N_2353,N_1653,N_1832);
nor U2354 (N_2354,N_1770,N_1941);
nand U2355 (N_2355,N_1970,N_1619);
and U2356 (N_2356,N_1940,N_1704);
nor U2357 (N_2357,N_1877,N_1872);
or U2358 (N_2358,N_1956,N_1569);
nor U2359 (N_2359,N_1917,N_1549);
and U2360 (N_2360,N_1516,N_1980);
and U2361 (N_2361,N_1538,N_1695);
and U2362 (N_2362,N_1695,N_1730);
nand U2363 (N_2363,N_1705,N_1583);
or U2364 (N_2364,N_1866,N_1624);
nand U2365 (N_2365,N_1607,N_1858);
nand U2366 (N_2366,N_1802,N_1524);
nand U2367 (N_2367,N_1510,N_1845);
or U2368 (N_2368,N_1947,N_1727);
nor U2369 (N_2369,N_1838,N_1777);
or U2370 (N_2370,N_1865,N_1998);
nand U2371 (N_2371,N_1723,N_1689);
nor U2372 (N_2372,N_1992,N_1668);
and U2373 (N_2373,N_1533,N_1797);
nand U2374 (N_2374,N_1602,N_1980);
and U2375 (N_2375,N_1847,N_1651);
or U2376 (N_2376,N_1684,N_1658);
nand U2377 (N_2377,N_1690,N_1731);
nand U2378 (N_2378,N_1749,N_1821);
nor U2379 (N_2379,N_1775,N_1906);
and U2380 (N_2380,N_1637,N_1734);
nor U2381 (N_2381,N_1771,N_1936);
or U2382 (N_2382,N_1899,N_1989);
and U2383 (N_2383,N_1599,N_1951);
or U2384 (N_2384,N_1571,N_1607);
nor U2385 (N_2385,N_1788,N_1846);
nor U2386 (N_2386,N_1880,N_1721);
or U2387 (N_2387,N_1697,N_1755);
or U2388 (N_2388,N_1527,N_1945);
or U2389 (N_2389,N_1681,N_1598);
nand U2390 (N_2390,N_1557,N_1945);
nand U2391 (N_2391,N_1579,N_1757);
and U2392 (N_2392,N_1754,N_1514);
nand U2393 (N_2393,N_1983,N_1842);
and U2394 (N_2394,N_1994,N_1699);
nor U2395 (N_2395,N_1874,N_1923);
nor U2396 (N_2396,N_1565,N_1523);
and U2397 (N_2397,N_1935,N_1501);
and U2398 (N_2398,N_1974,N_1884);
or U2399 (N_2399,N_1534,N_1527);
or U2400 (N_2400,N_1621,N_1636);
and U2401 (N_2401,N_1558,N_1989);
nand U2402 (N_2402,N_1506,N_1837);
nor U2403 (N_2403,N_1831,N_1633);
or U2404 (N_2404,N_1611,N_1623);
and U2405 (N_2405,N_1622,N_1590);
nand U2406 (N_2406,N_1738,N_1870);
nand U2407 (N_2407,N_1873,N_1916);
or U2408 (N_2408,N_1734,N_1812);
nor U2409 (N_2409,N_1599,N_1546);
and U2410 (N_2410,N_1590,N_1615);
and U2411 (N_2411,N_1580,N_1829);
or U2412 (N_2412,N_1798,N_1698);
nor U2413 (N_2413,N_1736,N_1696);
or U2414 (N_2414,N_1760,N_1686);
nand U2415 (N_2415,N_1864,N_1522);
nand U2416 (N_2416,N_1652,N_1539);
or U2417 (N_2417,N_1590,N_1505);
nor U2418 (N_2418,N_1889,N_1878);
nand U2419 (N_2419,N_1820,N_1685);
and U2420 (N_2420,N_1815,N_1673);
nor U2421 (N_2421,N_1580,N_1974);
or U2422 (N_2422,N_1725,N_1711);
nor U2423 (N_2423,N_1562,N_1670);
and U2424 (N_2424,N_1723,N_1966);
nor U2425 (N_2425,N_1957,N_1858);
and U2426 (N_2426,N_1834,N_1661);
nor U2427 (N_2427,N_1793,N_1979);
and U2428 (N_2428,N_1963,N_1910);
nor U2429 (N_2429,N_1581,N_1617);
or U2430 (N_2430,N_1975,N_1706);
nand U2431 (N_2431,N_1643,N_1617);
nand U2432 (N_2432,N_1768,N_1538);
nor U2433 (N_2433,N_1588,N_1881);
nand U2434 (N_2434,N_1940,N_1765);
nor U2435 (N_2435,N_1925,N_1753);
or U2436 (N_2436,N_1734,N_1886);
nand U2437 (N_2437,N_1797,N_1690);
and U2438 (N_2438,N_1863,N_1998);
nand U2439 (N_2439,N_1702,N_1593);
nor U2440 (N_2440,N_1695,N_1561);
and U2441 (N_2441,N_1828,N_1762);
nand U2442 (N_2442,N_1873,N_1886);
or U2443 (N_2443,N_1785,N_1705);
nand U2444 (N_2444,N_1766,N_1778);
and U2445 (N_2445,N_1851,N_1747);
nor U2446 (N_2446,N_1817,N_1529);
nand U2447 (N_2447,N_1615,N_1631);
nor U2448 (N_2448,N_1818,N_1827);
and U2449 (N_2449,N_1558,N_1568);
or U2450 (N_2450,N_1792,N_1597);
or U2451 (N_2451,N_1819,N_1578);
nand U2452 (N_2452,N_1902,N_1710);
nor U2453 (N_2453,N_1754,N_1908);
or U2454 (N_2454,N_1703,N_1589);
nand U2455 (N_2455,N_1831,N_1824);
and U2456 (N_2456,N_1959,N_1526);
nor U2457 (N_2457,N_1876,N_1830);
and U2458 (N_2458,N_1853,N_1825);
nor U2459 (N_2459,N_1586,N_1578);
nor U2460 (N_2460,N_1652,N_1994);
nor U2461 (N_2461,N_1553,N_1589);
and U2462 (N_2462,N_1908,N_1885);
nor U2463 (N_2463,N_1694,N_1873);
and U2464 (N_2464,N_1514,N_1984);
nand U2465 (N_2465,N_1536,N_1874);
nor U2466 (N_2466,N_1723,N_1528);
or U2467 (N_2467,N_1793,N_1671);
nand U2468 (N_2468,N_1770,N_1991);
nor U2469 (N_2469,N_1563,N_1643);
nand U2470 (N_2470,N_1662,N_1729);
and U2471 (N_2471,N_1938,N_1564);
nor U2472 (N_2472,N_1501,N_1655);
nand U2473 (N_2473,N_1846,N_1771);
nor U2474 (N_2474,N_1703,N_1888);
and U2475 (N_2475,N_1743,N_1504);
nand U2476 (N_2476,N_1809,N_1782);
and U2477 (N_2477,N_1728,N_1706);
nor U2478 (N_2478,N_1947,N_1978);
and U2479 (N_2479,N_1733,N_1937);
nand U2480 (N_2480,N_1940,N_1819);
nand U2481 (N_2481,N_1868,N_1646);
and U2482 (N_2482,N_1851,N_1923);
and U2483 (N_2483,N_1669,N_1720);
and U2484 (N_2484,N_1565,N_1811);
nand U2485 (N_2485,N_1742,N_1892);
nor U2486 (N_2486,N_1511,N_1616);
and U2487 (N_2487,N_1963,N_1873);
xor U2488 (N_2488,N_1795,N_1857);
or U2489 (N_2489,N_1741,N_1977);
or U2490 (N_2490,N_1693,N_1662);
nor U2491 (N_2491,N_1915,N_1927);
or U2492 (N_2492,N_1969,N_1709);
and U2493 (N_2493,N_1795,N_1533);
nand U2494 (N_2494,N_1763,N_1658);
xnor U2495 (N_2495,N_1941,N_1640);
nor U2496 (N_2496,N_1946,N_1869);
nor U2497 (N_2497,N_1616,N_1725);
nor U2498 (N_2498,N_1578,N_1708);
nor U2499 (N_2499,N_1643,N_1644);
nor U2500 (N_2500,N_2388,N_2408);
nand U2501 (N_2501,N_2372,N_2105);
nand U2502 (N_2502,N_2420,N_2196);
and U2503 (N_2503,N_2450,N_2265);
or U2504 (N_2504,N_2473,N_2235);
nand U2505 (N_2505,N_2064,N_2367);
nor U2506 (N_2506,N_2491,N_2212);
nand U2507 (N_2507,N_2488,N_2287);
or U2508 (N_2508,N_2003,N_2271);
and U2509 (N_2509,N_2415,N_2382);
nor U2510 (N_2510,N_2493,N_2411);
nor U2511 (N_2511,N_2170,N_2446);
or U2512 (N_2512,N_2209,N_2156);
or U2513 (N_2513,N_2466,N_2144);
nor U2514 (N_2514,N_2109,N_2073);
nand U2515 (N_2515,N_2464,N_2190);
and U2516 (N_2516,N_2165,N_2447);
nand U2517 (N_2517,N_2090,N_2045);
nand U2518 (N_2518,N_2387,N_2282);
and U2519 (N_2519,N_2023,N_2286);
nor U2520 (N_2520,N_2344,N_2469);
or U2521 (N_2521,N_2160,N_2189);
nand U2522 (N_2522,N_2242,N_2080);
or U2523 (N_2523,N_2324,N_2036);
or U2524 (N_2524,N_2245,N_2475);
and U2525 (N_2525,N_2322,N_2375);
and U2526 (N_2526,N_2078,N_2187);
or U2527 (N_2527,N_2363,N_2340);
and U2528 (N_2528,N_2397,N_2347);
nand U2529 (N_2529,N_2024,N_2285);
nand U2530 (N_2530,N_2010,N_2383);
nor U2531 (N_2531,N_2412,N_2207);
and U2532 (N_2532,N_2120,N_2208);
nand U2533 (N_2533,N_2311,N_2349);
and U2534 (N_2534,N_2146,N_2027);
or U2535 (N_2535,N_2484,N_2468);
and U2536 (N_2536,N_2039,N_2172);
nor U2537 (N_2537,N_2424,N_2335);
nor U2538 (N_2538,N_2358,N_2401);
and U2539 (N_2539,N_2485,N_2396);
or U2540 (N_2540,N_2257,N_2050);
nor U2541 (N_2541,N_2432,N_2317);
nor U2542 (N_2542,N_2251,N_2046);
or U2543 (N_2543,N_2250,N_2325);
and U2544 (N_2544,N_2370,N_2122);
nor U2545 (N_2545,N_2153,N_2161);
and U2546 (N_2546,N_2244,N_2422);
or U2547 (N_2547,N_2198,N_2402);
nand U2548 (N_2548,N_2148,N_2117);
nand U2549 (N_2549,N_2276,N_2259);
nor U2550 (N_2550,N_2186,N_2226);
and U2551 (N_2551,N_2478,N_2489);
or U2552 (N_2552,N_2483,N_2328);
or U2553 (N_2553,N_2055,N_2427);
nand U2554 (N_2554,N_2037,N_2356);
nor U2555 (N_2555,N_2275,N_2229);
nand U2556 (N_2556,N_2200,N_2185);
nor U2557 (N_2557,N_2127,N_2273);
and U2558 (N_2558,N_2091,N_2075);
and U2559 (N_2559,N_2194,N_2232);
or U2560 (N_2560,N_2240,N_2231);
or U2561 (N_2561,N_2135,N_2426);
nor U2562 (N_2562,N_2291,N_2206);
nand U2563 (N_2563,N_2013,N_2171);
nand U2564 (N_2564,N_2087,N_2454);
xor U2565 (N_2565,N_2445,N_2284);
or U2566 (N_2566,N_2204,N_2494);
nand U2567 (N_2567,N_2292,N_2314);
or U2568 (N_2568,N_2131,N_2044);
nand U2569 (N_2569,N_2352,N_2130);
and U2570 (N_2570,N_2453,N_2268);
and U2571 (N_2571,N_2498,N_2107);
nor U2572 (N_2572,N_2041,N_2100);
nand U2573 (N_2573,N_2093,N_2178);
or U2574 (N_2574,N_2428,N_2294);
nand U2575 (N_2575,N_2318,N_2042);
nand U2576 (N_2576,N_2440,N_2342);
nand U2577 (N_2577,N_2374,N_2476);
nand U2578 (N_2578,N_2048,N_2461);
or U2579 (N_2579,N_2327,N_2174);
nor U2580 (N_2580,N_2067,N_2459);
nand U2581 (N_2581,N_2357,N_2136);
and U2582 (N_2582,N_2029,N_2183);
nand U2583 (N_2583,N_2492,N_2418);
nor U2584 (N_2584,N_2191,N_2398);
nand U2585 (N_2585,N_2243,N_2002);
nor U2586 (N_2586,N_2474,N_2128);
nor U2587 (N_2587,N_2407,N_2481);
nor U2588 (N_2588,N_2393,N_2306);
and U2589 (N_2589,N_2015,N_2147);
or U2590 (N_2590,N_2364,N_2155);
or U2591 (N_2591,N_2004,N_2225);
and U2592 (N_2592,N_2213,N_2081);
nand U2593 (N_2593,N_2009,N_2070);
nand U2594 (N_2594,N_2026,N_2490);
nand U2595 (N_2595,N_2439,N_2366);
and U2596 (N_2596,N_2083,N_2233);
or U2597 (N_2597,N_2216,N_2258);
nor U2598 (N_2598,N_2381,N_2179);
and U2599 (N_2599,N_2436,N_2343);
or U2600 (N_2600,N_2162,N_2479);
nor U2601 (N_2601,N_2017,N_2221);
and U2602 (N_2602,N_2463,N_2077);
nand U2603 (N_2603,N_2047,N_2059);
or U2604 (N_2604,N_2058,N_2220);
or U2605 (N_2605,N_2019,N_2329);
nand U2606 (N_2606,N_2166,N_2458);
nor U2607 (N_2607,N_2201,N_2448);
nand U2608 (N_2608,N_2142,N_2319);
nand U2609 (N_2609,N_2305,N_2111);
nand U2610 (N_2610,N_2112,N_2061);
nor U2611 (N_2611,N_2301,N_2123);
nand U2612 (N_2612,N_2380,N_2316);
and U2613 (N_2613,N_2031,N_2006);
and U2614 (N_2614,N_2132,N_2098);
nor U2615 (N_2615,N_2323,N_2043);
and U2616 (N_2616,N_2433,N_2270);
nand U2617 (N_2617,N_2126,N_2088);
and U2618 (N_2618,N_2145,N_2192);
and U2619 (N_2619,N_2134,N_2496);
and U2620 (N_2620,N_2435,N_2076);
and U2621 (N_2621,N_2255,N_2133);
nand U2622 (N_2622,N_2264,N_2330);
nor U2623 (N_2623,N_2106,N_2038);
and U2624 (N_2624,N_2000,N_2379);
nor U2625 (N_2625,N_2182,N_2210);
nand U2626 (N_2626,N_2066,N_2230);
or U2627 (N_2627,N_2332,N_2497);
nor U2628 (N_2628,N_2272,N_2211);
nor U2629 (N_2629,N_2071,N_2267);
or U2630 (N_2630,N_2274,N_2199);
nor U2631 (N_2631,N_2032,N_2296);
and U2632 (N_2632,N_2337,N_2302);
or U2633 (N_2633,N_2254,N_2069);
and U2634 (N_2634,N_2280,N_2228);
and U2635 (N_2635,N_2290,N_2121);
nand U2636 (N_2636,N_2470,N_2092);
nand U2637 (N_2637,N_2389,N_2108);
or U2638 (N_2638,N_2115,N_2193);
or U2639 (N_2639,N_2089,N_2472);
nor U2640 (N_2640,N_2239,N_2394);
nand U2641 (N_2641,N_2152,N_2443);
and U2642 (N_2642,N_2410,N_2214);
and U2643 (N_2643,N_2406,N_2345);
or U2644 (N_2644,N_2390,N_2241);
nand U2645 (N_2645,N_2279,N_2346);
nor U2646 (N_2646,N_2278,N_2224);
nand U2647 (N_2647,N_2262,N_2405);
or U2648 (N_2648,N_2360,N_2359);
and U2649 (N_2649,N_2139,N_2299);
nand U2650 (N_2650,N_2096,N_2400);
and U2651 (N_2651,N_2320,N_2203);
or U2652 (N_2652,N_2223,N_2289);
or U2653 (N_2653,N_2137,N_2403);
nand U2654 (N_2654,N_2028,N_2072);
or U2655 (N_2655,N_2177,N_2065);
nand U2656 (N_2656,N_2103,N_2168);
or U2657 (N_2657,N_2423,N_2124);
and U2658 (N_2658,N_2295,N_2007);
and U2659 (N_2659,N_2351,N_2012);
nor U2660 (N_2660,N_2238,N_2429);
or U2661 (N_2661,N_2033,N_2062);
nand U2662 (N_2662,N_2247,N_2151);
or U2663 (N_2663,N_2253,N_2414);
nor U2664 (N_2664,N_2163,N_2074);
or U2665 (N_2665,N_2315,N_2308);
nand U2666 (N_2666,N_2277,N_2441);
nor U2667 (N_2667,N_2113,N_2021);
nand U2668 (N_2668,N_2348,N_2499);
and U2669 (N_2669,N_2495,N_2261);
nand U2670 (N_2670,N_2222,N_2056);
nor U2671 (N_2671,N_2362,N_2181);
nor U2672 (N_2672,N_2378,N_2237);
or U2673 (N_2673,N_2263,N_2086);
nor U2674 (N_2674,N_2022,N_2283);
or U2675 (N_2675,N_2060,N_2079);
and U2676 (N_2676,N_2057,N_2350);
nand U2677 (N_2677,N_2312,N_2456);
nor U2678 (N_2678,N_2377,N_2434);
or U2679 (N_2679,N_2460,N_2102);
and U2680 (N_2680,N_2125,N_2154);
or U2681 (N_2681,N_2413,N_2197);
nor U2682 (N_2682,N_2099,N_2008);
or U2683 (N_2683,N_2252,N_2467);
nand U2684 (N_2684,N_2035,N_2040);
nand U2685 (N_2685,N_2425,N_2334);
or U2686 (N_2686,N_2246,N_2150);
nor U2687 (N_2687,N_2471,N_2399);
and U2688 (N_2688,N_2333,N_2063);
or U2689 (N_2689,N_2431,N_2053);
and U2690 (N_2690,N_2480,N_2438);
and U2691 (N_2691,N_2234,N_2068);
and U2692 (N_2692,N_2095,N_2001);
nand U2693 (N_2693,N_2462,N_2114);
and U2694 (N_2694,N_2129,N_2011);
nor U2695 (N_2695,N_2336,N_2376);
nand U2696 (N_2696,N_2217,N_2384);
and U2697 (N_2697,N_2169,N_2385);
or U2698 (N_2698,N_2157,N_2373);
or U2699 (N_2699,N_2417,N_2298);
and U2700 (N_2700,N_2110,N_2149);
and U2701 (N_2701,N_2341,N_2138);
and U2702 (N_2702,N_2020,N_2353);
nand U2703 (N_2703,N_2202,N_2014);
nand U2704 (N_2704,N_2310,N_2248);
and U2705 (N_2705,N_2386,N_2005);
or U2706 (N_2706,N_2085,N_2368);
and U2707 (N_2707,N_2084,N_2309);
nor U2708 (N_2708,N_2404,N_2256);
nand U2709 (N_2709,N_2052,N_2219);
or U2710 (N_2710,N_2140,N_2188);
or U2711 (N_2711,N_2281,N_2249);
and U2712 (N_2712,N_2167,N_2184);
nand U2713 (N_2713,N_2116,N_2051);
and U2714 (N_2714,N_2430,N_2101);
nor U2715 (N_2715,N_2164,N_2195);
nand U2716 (N_2716,N_2371,N_2049);
nor U2717 (N_2717,N_2326,N_2218);
or U2718 (N_2718,N_2354,N_2339);
and U2719 (N_2719,N_2082,N_2444);
or U2720 (N_2720,N_2416,N_2173);
and U2721 (N_2721,N_2391,N_2094);
nor U2722 (N_2722,N_2016,N_2452);
nand U2723 (N_2723,N_2392,N_2260);
and U2724 (N_2724,N_2437,N_2409);
nor U2725 (N_2725,N_2269,N_2457);
nand U2726 (N_2726,N_2421,N_2297);
or U2727 (N_2727,N_2175,N_2355);
or U2728 (N_2728,N_2451,N_2442);
nor U2729 (N_2729,N_2300,N_2487);
nor U2730 (N_2730,N_2180,N_2215);
and U2731 (N_2731,N_2365,N_2034);
or U2732 (N_2732,N_2303,N_2176);
or U2733 (N_2733,N_2455,N_2118);
nor U2734 (N_2734,N_2236,N_2449);
nand U2735 (N_2735,N_2486,N_2338);
and U2736 (N_2736,N_2119,N_2477);
and U2737 (N_2737,N_2025,N_2482);
or U2738 (N_2738,N_2143,N_2266);
nor U2739 (N_2739,N_2395,N_2054);
nand U2740 (N_2740,N_2293,N_2331);
and U2741 (N_2741,N_2159,N_2141);
nor U2742 (N_2742,N_2465,N_2205);
nand U2743 (N_2743,N_2419,N_2361);
or U2744 (N_2744,N_2030,N_2104);
and U2745 (N_2745,N_2307,N_2304);
and U2746 (N_2746,N_2018,N_2313);
or U2747 (N_2747,N_2321,N_2369);
nor U2748 (N_2748,N_2097,N_2227);
nand U2749 (N_2749,N_2158,N_2288);
nand U2750 (N_2750,N_2381,N_2121);
nand U2751 (N_2751,N_2416,N_2085);
nor U2752 (N_2752,N_2331,N_2180);
or U2753 (N_2753,N_2431,N_2171);
and U2754 (N_2754,N_2138,N_2008);
nand U2755 (N_2755,N_2332,N_2406);
nor U2756 (N_2756,N_2332,N_2210);
nor U2757 (N_2757,N_2043,N_2370);
or U2758 (N_2758,N_2235,N_2428);
or U2759 (N_2759,N_2022,N_2154);
or U2760 (N_2760,N_2369,N_2247);
or U2761 (N_2761,N_2301,N_2477);
or U2762 (N_2762,N_2115,N_2295);
nand U2763 (N_2763,N_2348,N_2336);
or U2764 (N_2764,N_2006,N_2066);
or U2765 (N_2765,N_2445,N_2490);
and U2766 (N_2766,N_2467,N_2123);
or U2767 (N_2767,N_2221,N_2035);
nor U2768 (N_2768,N_2292,N_2313);
nand U2769 (N_2769,N_2188,N_2308);
nor U2770 (N_2770,N_2006,N_2336);
nor U2771 (N_2771,N_2342,N_2388);
and U2772 (N_2772,N_2019,N_2193);
or U2773 (N_2773,N_2453,N_2071);
nor U2774 (N_2774,N_2430,N_2431);
nor U2775 (N_2775,N_2256,N_2344);
and U2776 (N_2776,N_2260,N_2153);
or U2777 (N_2777,N_2387,N_2465);
nand U2778 (N_2778,N_2034,N_2234);
or U2779 (N_2779,N_2477,N_2047);
nand U2780 (N_2780,N_2273,N_2051);
and U2781 (N_2781,N_2213,N_2170);
nor U2782 (N_2782,N_2401,N_2144);
nor U2783 (N_2783,N_2380,N_2292);
nand U2784 (N_2784,N_2010,N_2411);
nand U2785 (N_2785,N_2071,N_2401);
and U2786 (N_2786,N_2286,N_2202);
or U2787 (N_2787,N_2241,N_2379);
or U2788 (N_2788,N_2488,N_2373);
or U2789 (N_2789,N_2495,N_2334);
nor U2790 (N_2790,N_2081,N_2390);
nor U2791 (N_2791,N_2398,N_2372);
and U2792 (N_2792,N_2365,N_2147);
nor U2793 (N_2793,N_2195,N_2346);
nor U2794 (N_2794,N_2388,N_2492);
nand U2795 (N_2795,N_2003,N_2481);
or U2796 (N_2796,N_2407,N_2406);
or U2797 (N_2797,N_2198,N_2193);
nor U2798 (N_2798,N_2111,N_2331);
or U2799 (N_2799,N_2216,N_2320);
or U2800 (N_2800,N_2101,N_2389);
or U2801 (N_2801,N_2169,N_2448);
and U2802 (N_2802,N_2166,N_2024);
nand U2803 (N_2803,N_2458,N_2071);
and U2804 (N_2804,N_2007,N_2104);
nand U2805 (N_2805,N_2222,N_2488);
nor U2806 (N_2806,N_2493,N_2110);
and U2807 (N_2807,N_2225,N_2097);
and U2808 (N_2808,N_2239,N_2246);
nand U2809 (N_2809,N_2161,N_2390);
nor U2810 (N_2810,N_2484,N_2217);
or U2811 (N_2811,N_2103,N_2459);
and U2812 (N_2812,N_2465,N_2451);
or U2813 (N_2813,N_2451,N_2135);
nor U2814 (N_2814,N_2185,N_2176);
and U2815 (N_2815,N_2133,N_2264);
and U2816 (N_2816,N_2404,N_2137);
and U2817 (N_2817,N_2394,N_2139);
or U2818 (N_2818,N_2381,N_2224);
nor U2819 (N_2819,N_2165,N_2061);
nand U2820 (N_2820,N_2150,N_2182);
or U2821 (N_2821,N_2254,N_2220);
nand U2822 (N_2822,N_2194,N_2349);
or U2823 (N_2823,N_2301,N_2261);
nor U2824 (N_2824,N_2012,N_2087);
or U2825 (N_2825,N_2110,N_2036);
nand U2826 (N_2826,N_2402,N_2207);
or U2827 (N_2827,N_2478,N_2081);
and U2828 (N_2828,N_2060,N_2419);
nand U2829 (N_2829,N_2340,N_2123);
nor U2830 (N_2830,N_2311,N_2140);
nand U2831 (N_2831,N_2264,N_2418);
nand U2832 (N_2832,N_2185,N_2114);
nand U2833 (N_2833,N_2307,N_2377);
nand U2834 (N_2834,N_2182,N_2163);
and U2835 (N_2835,N_2130,N_2412);
or U2836 (N_2836,N_2210,N_2262);
nand U2837 (N_2837,N_2247,N_2217);
nand U2838 (N_2838,N_2352,N_2357);
nand U2839 (N_2839,N_2126,N_2143);
and U2840 (N_2840,N_2418,N_2167);
or U2841 (N_2841,N_2272,N_2315);
nor U2842 (N_2842,N_2232,N_2420);
and U2843 (N_2843,N_2022,N_2198);
or U2844 (N_2844,N_2117,N_2392);
or U2845 (N_2845,N_2327,N_2370);
nor U2846 (N_2846,N_2445,N_2141);
nor U2847 (N_2847,N_2016,N_2119);
or U2848 (N_2848,N_2416,N_2297);
nand U2849 (N_2849,N_2298,N_2395);
and U2850 (N_2850,N_2252,N_2125);
and U2851 (N_2851,N_2227,N_2243);
and U2852 (N_2852,N_2422,N_2174);
nand U2853 (N_2853,N_2441,N_2282);
or U2854 (N_2854,N_2479,N_2303);
and U2855 (N_2855,N_2298,N_2398);
nor U2856 (N_2856,N_2308,N_2084);
nand U2857 (N_2857,N_2170,N_2376);
nor U2858 (N_2858,N_2194,N_2021);
nand U2859 (N_2859,N_2170,N_2215);
or U2860 (N_2860,N_2250,N_2114);
nand U2861 (N_2861,N_2109,N_2209);
nand U2862 (N_2862,N_2352,N_2113);
nand U2863 (N_2863,N_2178,N_2268);
nand U2864 (N_2864,N_2092,N_2046);
nor U2865 (N_2865,N_2122,N_2440);
or U2866 (N_2866,N_2472,N_2475);
nand U2867 (N_2867,N_2474,N_2473);
and U2868 (N_2868,N_2390,N_2269);
or U2869 (N_2869,N_2383,N_2054);
or U2870 (N_2870,N_2211,N_2310);
and U2871 (N_2871,N_2275,N_2207);
or U2872 (N_2872,N_2168,N_2224);
nor U2873 (N_2873,N_2015,N_2053);
nor U2874 (N_2874,N_2347,N_2089);
nor U2875 (N_2875,N_2023,N_2049);
or U2876 (N_2876,N_2036,N_2469);
nor U2877 (N_2877,N_2188,N_2250);
or U2878 (N_2878,N_2110,N_2164);
nor U2879 (N_2879,N_2322,N_2496);
nor U2880 (N_2880,N_2472,N_2196);
or U2881 (N_2881,N_2382,N_2450);
or U2882 (N_2882,N_2243,N_2079);
and U2883 (N_2883,N_2390,N_2028);
or U2884 (N_2884,N_2078,N_2255);
nor U2885 (N_2885,N_2428,N_2234);
nand U2886 (N_2886,N_2387,N_2274);
nor U2887 (N_2887,N_2474,N_2269);
nand U2888 (N_2888,N_2134,N_2246);
or U2889 (N_2889,N_2343,N_2117);
and U2890 (N_2890,N_2077,N_2449);
nand U2891 (N_2891,N_2372,N_2113);
and U2892 (N_2892,N_2120,N_2280);
or U2893 (N_2893,N_2285,N_2471);
nand U2894 (N_2894,N_2403,N_2295);
nor U2895 (N_2895,N_2066,N_2214);
and U2896 (N_2896,N_2085,N_2177);
nand U2897 (N_2897,N_2388,N_2131);
or U2898 (N_2898,N_2143,N_2084);
or U2899 (N_2899,N_2203,N_2171);
nand U2900 (N_2900,N_2411,N_2247);
and U2901 (N_2901,N_2058,N_2446);
nor U2902 (N_2902,N_2122,N_2102);
nand U2903 (N_2903,N_2383,N_2309);
xnor U2904 (N_2904,N_2425,N_2309);
nand U2905 (N_2905,N_2421,N_2140);
and U2906 (N_2906,N_2259,N_2114);
or U2907 (N_2907,N_2099,N_2479);
and U2908 (N_2908,N_2143,N_2138);
nand U2909 (N_2909,N_2334,N_2157);
and U2910 (N_2910,N_2284,N_2293);
or U2911 (N_2911,N_2104,N_2058);
or U2912 (N_2912,N_2214,N_2495);
or U2913 (N_2913,N_2464,N_2484);
and U2914 (N_2914,N_2251,N_2481);
and U2915 (N_2915,N_2483,N_2265);
nand U2916 (N_2916,N_2467,N_2409);
and U2917 (N_2917,N_2307,N_2029);
and U2918 (N_2918,N_2197,N_2135);
or U2919 (N_2919,N_2017,N_2396);
and U2920 (N_2920,N_2387,N_2084);
or U2921 (N_2921,N_2478,N_2038);
nand U2922 (N_2922,N_2363,N_2221);
nand U2923 (N_2923,N_2143,N_2183);
nor U2924 (N_2924,N_2164,N_2209);
and U2925 (N_2925,N_2233,N_2242);
or U2926 (N_2926,N_2091,N_2439);
nor U2927 (N_2927,N_2235,N_2379);
nor U2928 (N_2928,N_2276,N_2076);
nor U2929 (N_2929,N_2376,N_2082);
or U2930 (N_2930,N_2270,N_2466);
xnor U2931 (N_2931,N_2016,N_2099);
nand U2932 (N_2932,N_2004,N_2253);
nand U2933 (N_2933,N_2258,N_2364);
nor U2934 (N_2934,N_2021,N_2035);
or U2935 (N_2935,N_2054,N_2218);
and U2936 (N_2936,N_2403,N_2124);
or U2937 (N_2937,N_2023,N_2440);
and U2938 (N_2938,N_2375,N_2356);
or U2939 (N_2939,N_2408,N_2406);
nand U2940 (N_2940,N_2301,N_2082);
nor U2941 (N_2941,N_2304,N_2114);
and U2942 (N_2942,N_2258,N_2018);
and U2943 (N_2943,N_2163,N_2304);
nand U2944 (N_2944,N_2391,N_2385);
and U2945 (N_2945,N_2222,N_2092);
or U2946 (N_2946,N_2070,N_2411);
nor U2947 (N_2947,N_2297,N_2310);
nand U2948 (N_2948,N_2171,N_2119);
nor U2949 (N_2949,N_2440,N_2367);
or U2950 (N_2950,N_2215,N_2452);
or U2951 (N_2951,N_2024,N_2064);
nor U2952 (N_2952,N_2114,N_2146);
or U2953 (N_2953,N_2344,N_2380);
and U2954 (N_2954,N_2036,N_2136);
nand U2955 (N_2955,N_2403,N_2063);
nand U2956 (N_2956,N_2253,N_2182);
nor U2957 (N_2957,N_2165,N_2054);
or U2958 (N_2958,N_2165,N_2167);
nand U2959 (N_2959,N_2179,N_2080);
nor U2960 (N_2960,N_2253,N_2317);
and U2961 (N_2961,N_2462,N_2098);
or U2962 (N_2962,N_2035,N_2036);
or U2963 (N_2963,N_2442,N_2492);
or U2964 (N_2964,N_2377,N_2011);
or U2965 (N_2965,N_2218,N_2128);
or U2966 (N_2966,N_2448,N_2340);
or U2967 (N_2967,N_2299,N_2279);
and U2968 (N_2968,N_2038,N_2293);
nor U2969 (N_2969,N_2374,N_2186);
nand U2970 (N_2970,N_2348,N_2490);
nor U2971 (N_2971,N_2049,N_2120);
nor U2972 (N_2972,N_2106,N_2109);
nand U2973 (N_2973,N_2201,N_2267);
or U2974 (N_2974,N_2354,N_2030);
nand U2975 (N_2975,N_2004,N_2090);
nor U2976 (N_2976,N_2413,N_2247);
or U2977 (N_2977,N_2318,N_2062);
nand U2978 (N_2978,N_2006,N_2327);
and U2979 (N_2979,N_2459,N_2034);
and U2980 (N_2980,N_2263,N_2159);
and U2981 (N_2981,N_2022,N_2044);
nand U2982 (N_2982,N_2131,N_2028);
nor U2983 (N_2983,N_2124,N_2324);
nor U2984 (N_2984,N_2054,N_2307);
or U2985 (N_2985,N_2021,N_2139);
and U2986 (N_2986,N_2166,N_2008);
nand U2987 (N_2987,N_2463,N_2045);
nand U2988 (N_2988,N_2061,N_2457);
nor U2989 (N_2989,N_2450,N_2072);
and U2990 (N_2990,N_2356,N_2339);
nor U2991 (N_2991,N_2380,N_2436);
nor U2992 (N_2992,N_2271,N_2153);
and U2993 (N_2993,N_2414,N_2141);
nor U2994 (N_2994,N_2495,N_2381);
nand U2995 (N_2995,N_2061,N_2025);
nor U2996 (N_2996,N_2230,N_2212);
xor U2997 (N_2997,N_2117,N_2195);
and U2998 (N_2998,N_2248,N_2374);
nor U2999 (N_2999,N_2253,N_2461);
or UO_0 (O_0,N_2504,N_2627);
or UO_1 (O_1,N_2834,N_2761);
and UO_2 (O_2,N_2605,N_2900);
nand UO_3 (O_3,N_2954,N_2674);
nand UO_4 (O_4,N_2688,N_2727);
and UO_5 (O_5,N_2712,N_2860);
nor UO_6 (O_6,N_2572,N_2752);
nor UO_7 (O_7,N_2971,N_2799);
and UO_8 (O_8,N_2975,N_2938);
nor UO_9 (O_9,N_2555,N_2581);
nor UO_10 (O_10,N_2503,N_2873);
nor UO_11 (O_11,N_2556,N_2675);
and UO_12 (O_12,N_2726,N_2601);
nand UO_13 (O_13,N_2550,N_2853);
or UO_14 (O_14,N_2604,N_2725);
nand UO_15 (O_15,N_2665,N_2732);
nand UO_16 (O_16,N_2586,N_2989);
or UO_17 (O_17,N_2753,N_2751);
or UO_18 (O_18,N_2817,N_2673);
nor UO_19 (O_19,N_2606,N_2870);
xnor UO_20 (O_20,N_2646,N_2561);
nand UO_21 (O_21,N_2831,N_2632);
or UO_22 (O_22,N_2956,N_2655);
nor UO_23 (O_23,N_2827,N_2592);
nor UO_24 (O_24,N_2825,N_2829);
and UO_25 (O_25,N_2837,N_2843);
nor UO_26 (O_26,N_2519,N_2536);
and UO_27 (O_27,N_2777,N_2734);
nand UO_28 (O_28,N_2925,N_2551);
nand UO_29 (O_29,N_2541,N_2995);
or UO_30 (O_30,N_2931,N_2939);
or UO_31 (O_31,N_2908,N_2877);
nand UO_32 (O_32,N_2540,N_2524);
or UO_33 (O_33,N_2861,N_2537);
or UO_34 (O_34,N_2669,N_2576);
nand UO_35 (O_35,N_2636,N_2695);
nand UO_36 (O_36,N_2641,N_2905);
nor UO_37 (O_37,N_2949,N_2608);
nand UO_38 (O_38,N_2667,N_2657);
nand UO_39 (O_39,N_2659,N_2681);
or UO_40 (O_40,N_2912,N_2992);
nor UO_41 (O_41,N_2934,N_2922);
nor UO_42 (O_42,N_2525,N_2617);
nand UO_43 (O_43,N_2963,N_2784);
nor UO_44 (O_44,N_2693,N_2991);
nor UO_45 (O_45,N_2863,N_2595);
or UO_46 (O_46,N_2663,N_2756);
nor UO_47 (O_47,N_2534,N_2542);
nor UO_48 (O_48,N_2684,N_2848);
nand UO_49 (O_49,N_2505,N_2891);
nor UO_50 (O_50,N_2716,N_2506);
or UO_51 (O_51,N_2921,N_2547);
nand UO_52 (O_52,N_2762,N_2836);
or UO_53 (O_53,N_2806,N_2520);
and UO_54 (O_54,N_2973,N_2988);
nand UO_55 (O_55,N_2630,N_2633);
and UO_56 (O_56,N_2867,N_2924);
nor UO_57 (O_57,N_2927,N_2917);
nor UO_58 (O_58,N_2888,N_2708);
or UO_59 (O_59,N_2598,N_2911);
and UO_60 (O_60,N_2903,N_2749);
nand UO_61 (O_61,N_2782,N_2559);
and UO_62 (O_62,N_2514,N_2558);
or UO_63 (O_63,N_2634,N_2985);
or UO_64 (O_64,N_2745,N_2878);
nand UO_65 (O_65,N_2585,N_2666);
nand UO_66 (O_66,N_2826,N_2578);
or UO_67 (O_67,N_2647,N_2687);
nor UO_68 (O_68,N_2818,N_2807);
nor UO_69 (O_69,N_2517,N_2719);
or UO_70 (O_70,N_2960,N_2770);
nor UO_71 (O_71,N_2968,N_2746);
and UO_72 (O_72,N_2625,N_2933);
nand UO_73 (O_73,N_2685,N_2683);
nor UO_74 (O_74,N_2564,N_2796);
or UO_75 (O_75,N_2652,N_2722);
or UO_76 (O_76,N_2729,N_2629);
nor UO_77 (O_77,N_2760,N_2950);
nor UO_78 (O_78,N_2898,N_2914);
nand UO_79 (O_79,N_2513,N_2713);
or UO_80 (O_80,N_2679,N_2563);
and UO_81 (O_81,N_2830,N_2887);
and UO_82 (O_82,N_2781,N_2590);
nor UO_83 (O_83,N_2615,N_2866);
nand UO_84 (O_84,N_2603,N_2672);
and UO_85 (O_85,N_2723,N_2599);
or UO_86 (O_86,N_2802,N_2509);
nor UO_87 (O_87,N_2821,N_2893);
or UO_88 (O_88,N_2735,N_2668);
nand UO_89 (O_89,N_2923,N_2913);
and UO_90 (O_90,N_2650,N_2835);
nand UO_91 (O_91,N_2699,N_2886);
nor UO_92 (O_92,N_2611,N_2801);
nand UO_93 (O_93,N_2724,N_2850);
nor UO_94 (O_94,N_2677,N_2872);
and UO_95 (O_95,N_2983,N_2895);
nor UO_96 (O_96,N_2842,N_2771);
and UO_97 (O_97,N_2705,N_2910);
or UO_98 (O_98,N_2528,N_2526);
nor UO_99 (O_99,N_2553,N_2757);
nor UO_100 (O_100,N_2822,N_2743);
nor UO_101 (O_101,N_2808,N_2964);
nor UO_102 (O_102,N_2738,N_2736);
nand UO_103 (O_103,N_2941,N_2859);
nor UO_104 (O_104,N_2588,N_2907);
nor UO_105 (O_105,N_2943,N_2763);
nor UO_106 (O_106,N_2994,N_2730);
or UO_107 (O_107,N_2889,N_2621);
and UO_108 (O_108,N_2974,N_2548);
and UO_109 (O_109,N_2814,N_2996);
nand UO_110 (O_110,N_2946,N_2562);
and UO_111 (O_111,N_2501,N_2747);
or UO_112 (O_112,N_2987,N_2717);
and UO_113 (O_113,N_2841,N_2820);
or UO_114 (O_114,N_2686,N_2631);
nor UO_115 (O_115,N_2809,N_2651);
nor UO_116 (O_116,N_2883,N_2890);
and UO_117 (O_117,N_2929,N_2546);
and UO_118 (O_118,N_2765,N_2543);
nor UO_119 (O_119,N_2823,N_2942);
or UO_120 (O_120,N_2754,N_2544);
nor UO_121 (O_121,N_2567,N_2869);
nand UO_122 (O_122,N_2847,N_2703);
or UO_123 (O_123,N_2856,N_2709);
nand UO_124 (O_124,N_2791,N_2694);
nor UO_125 (O_125,N_2602,N_2584);
or UO_126 (O_126,N_2769,N_2803);
nand UO_127 (O_127,N_2515,N_2502);
or UO_128 (O_128,N_2570,N_2928);
and UO_129 (O_129,N_2951,N_2858);
and UO_130 (O_130,N_2653,N_2824);
or UO_131 (O_131,N_2610,N_2804);
nand UO_132 (O_132,N_2772,N_2786);
or UO_133 (O_133,N_2879,N_2533);
nor UO_134 (O_134,N_2612,N_2812);
nor UO_135 (O_135,N_2768,N_2748);
or UO_136 (O_136,N_2697,N_2969);
nor UO_137 (O_137,N_2696,N_2982);
and UO_138 (O_138,N_2737,N_2638);
nor UO_139 (O_139,N_2521,N_2511);
nor UO_140 (O_140,N_2618,N_2930);
nor UO_141 (O_141,N_2776,N_2915);
or UO_142 (O_142,N_2701,N_2876);
and UO_143 (O_143,N_2865,N_2523);
nand UO_144 (O_144,N_2901,N_2654);
and UO_145 (O_145,N_2792,N_2899);
or UO_146 (O_146,N_2571,N_2845);
or UO_147 (O_147,N_2645,N_2678);
or UO_148 (O_148,N_2980,N_2794);
nor UO_149 (O_149,N_2906,N_2958);
nand UO_150 (O_150,N_2984,N_2874);
nor UO_151 (O_151,N_2690,N_2628);
and UO_152 (O_152,N_2692,N_2970);
nor UO_153 (O_153,N_2864,N_2575);
nor UO_154 (O_154,N_2805,N_2711);
and UO_155 (O_155,N_2739,N_2977);
nand UO_156 (O_156,N_2779,N_2593);
nand UO_157 (O_157,N_2600,N_2662);
nand UO_158 (O_158,N_2766,N_2518);
or UO_159 (O_159,N_2787,N_2851);
nand UO_160 (O_160,N_2531,N_2702);
or UO_161 (O_161,N_2670,N_2828);
and UO_162 (O_162,N_2707,N_2948);
and UO_163 (O_163,N_2635,N_2959);
or UO_164 (O_164,N_2759,N_2965);
nand UO_165 (O_165,N_2839,N_2691);
xnor UO_166 (O_166,N_2616,N_2909);
and UO_167 (O_167,N_2740,N_2795);
or UO_168 (O_168,N_2955,N_2833);
or UO_169 (O_169,N_2619,N_2952);
nor UO_170 (O_170,N_2706,N_2516);
and UO_171 (O_171,N_2966,N_2932);
nand UO_172 (O_172,N_2815,N_2643);
nor UO_173 (O_173,N_2591,N_2767);
or UO_174 (O_174,N_2990,N_2811);
or UO_175 (O_175,N_2785,N_2800);
or UO_176 (O_176,N_2671,N_2979);
and UO_177 (O_177,N_2844,N_2728);
and UO_178 (O_178,N_2577,N_2507);
nor UO_179 (O_179,N_2580,N_2937);
or UO_180 (O_180,N_2545,N_2897);
or UO_181 (O_181,N_2918,N_2640);
nand UO_182 (O_182,N_2565,N_2981);
and UO_183 (O_183,N_2510,N_2557);
nor UO_184 (O_184,N_2579,N_2780);
or UO_185 (O_185,N_2552,N_2527);
or UO_186 (O_186,N_2620,N_2904);
and UO_187 (O_187,N_2976,N_2953);
nand UO_188 (O_188,N_2832,N_2649);
nor UO_189 (O_189,N_2962,N_2894);
or UO_190 (O_190,N_2849,N_2744);
or UO_191 (O_191,N_2607,N_2664);
or UO_192 (O_192,N_2945,N_2500);
nand UO_193 (O_193,N_2919,N_2597);
nand UO_194 (O_194,N_2682,N_2700);
and UO_195 (O_195,N_2775,N_2731);
or UO_196 (O_196,N_2582,N_2566);
and UO_197 (O_197,N_2720,N_2885);
or UO_198 (O_198,N_2854,N_2940);
nor UO_199 (O_199,N_2587,N_2742);
nand UO_200 (O_200,N_2522,N_2755);
nand UO_201 (O_201,N_2790,N_2978);
nand UO_202 (O_202,N_2609,N_2594);
or UO_203 (O_203,N_2778,N_2661);
nor UO_204 (O_204,N_2997,N_2758);
nor UO_205 (O_205,N_2733,N_2644);
xor UO_206 (O_206,N_2986,N_2624);
or UO_207 (O_207,N_2596,N_2947);
or UO_208 (O_208,N_2783,N_2680);
nor UO_209 (O_209,N_2656,N_2623);
nand UO_210 (O_210,N_2999,N_2813);
nor UO_211 (O_211,N_2855,N_2935);
or UO_212 (O_212,N_2569,N_2718);
nand UO_213 (O_213,N_2875,N_2613);
and UO_214 (O_214,N_2857,N_2741);
nand UO_215 (O_215,N_2944,N_2838);
nor UO_216 (O_216,N_2816,N_2715);
or UO_217 (O_217,N_2626,N_2936);
nor UO_218 (O_218,N_2589,N_2920);
and UO_219 (O_219,N_2710,N_2573);
and UO_220 (O_220,N_2793,N_2789);
nand UO_221 (O_221,N_2614,N_2862);
and UO_222 (O_222,N_2639,N_2798);
nand UO_223 (O_223,N_2840,N_2574);
and UO_224 (O_224,N_2773,N_2902);
and UO_225 (O_225,N_2512,N_2568);
nand UO_226 (O_226,N_2750,N_2993);
nor UO_227 (O_227,N_2714,N_2689);
nand UO_228 (O_228,N_2797,N_2868);
nand UO_229 (O_229,N_2882,N_2967);
and UO_230 (O_230,N_2622,N_2508);
nand UO_231 (O_231,N_2698,N_2764);
nand UO_232 (O_232,N_2554,N_2819);
nand UO_233 (O_233,N_2810,N_2880);
and UO_234 (O_234,N_2530,N_2539);
and UO_235 (O_235,N_2704,N_2871);
or UO_236 (O_236,N_2972,N_2642);
or UO_237 (O_237,N_2676,N_2535);
or UO_238 (O_238,N_2721,N_2538);
and UO_239 (O_239,N_2658,N_2892);
xor UO_240 (O_240,N_2660,N_2583);
nor UO_241 (O_241,N_2916,N_2852);
nor UO_242 (O_242,N_2884,N_2896);
and UO_243 (O_243,N_2846,N_2529);
nand UO_244 (O_244,N_2532,N_2560);
nor UO_245 (O_245,N_2637,N_2926);
xnor UO_246 (O_246,N_2957,N_2788);
nand UO_247 (O_247,N_2648,N_2549);
and UO_248 (O_248,N_2881,N_2774);
and UO_249 (O_249,N_2961,N_2998);
or UO_250 (O_250,N_2681,N_2975);
nor UO_251 (O_251,N_2941,N_2959);
nand UO_252 (O_252,N_2774,N_2671);
and UO_253 (O_253,N_2641,N_2927);
or UO_254 (O_254,N_2507,N_2911);
nand UO_255 (O_255,N_2695,N_2692);
and UO_256 (O_256,N_2819,N_2537);
or UO_257 (O_257,N_2868,N_2810);
and UO_258 (O_258,N_2585,N_2695);
or UO_259 (O_259,N_2859,N_2608);
nand UO_260 (O_260,N_2659,N_2683);
or UO_261 (O_261,N_2898,N_2795);
and UO_262 (O_262,N_2881,N_2804);
or UO_263 (O_263,N_2905,N_2547);
and UO_264 (O_264,N_2552,N_2630);
nor UO_265 (O_265,N_2895,N_2682);
or UO_266 (O_266,N_2913,N_2788);
nand UO_267 (O_267,N_2616,N_2723);
nand UO_268 (O_268,N_2865,N_2616);
or UO_269 (O_269,N_2955,N_2953);
nor UO_270 (O_270,N_2825,N_2700);
or UO_271 (O_271,N_2599,N_2893);
or UO_272 (O_272,N_2972,N_2527);
or UO_273 (O_273,N_2800,N_2677);
or UO_274 (O_274,N_2513,N_2784);
nand UO_275 (O_275,N_2886,N_2860);
or UO_276 (O_276,N_2515,N_2694);
and UO_277 (O_277,N_2716,N_2944);
or UO_278 (O_278,N_2718,N_2708);
nor UO_279 (O_279,N_2755,N_2649);
nor UO_280 (O_280,N_2821,N_2963);
and UO_281 (O_281,N_2776,N_2544);
xnor UO_282 (O_282,N_2617,N_2662);
nand UO_283 (O_283,N_2948,N_2922);
or UO_284 (O_284,N_2670,N_2555);
and UO_285 (O_285,N_2876,N_2969);
or UO_286 (O_286,N_2509,N_2649);
nand UO_287 (O_287,N_2910,N_2846);
nand UO_288 (O_288,N_2555,N_2565);
nor UO_289 (O_289,N_2928,N_2717);
and UO_290 (O_290,N_2520,N_2538);
nor UO_291 (O_291,N_2933,N_2705);
nor UO_292 (O_292,N_2630,N_2744);
nor UO_293 (O_293,N_2635,N_2533);
nand UO_294 (O_294,N_2987,N_2920);
or UO_295 (O_295,N_2765,N_2703);
nand UO_296 (O_296,N_2949,N_2703);
and UO_297 (O_297,N_2760,N_2986);
nand UO_298 (O_298,N_2734,N_2782);
nor UO_299 (O_299,N_2946,N_2983);
or UO_300 (O_300,N_2530,N_2543);
and UO_301 (O_301,N_2990,N_2558);
or UO_302 (O_302,N_2935,N_2926);
and UO_303 (O_303,N_2865,N_2781);
nor UO_304 (O_304,N_2790,N_2830);
nand UO_305 (O_305,N_2677,N_2972);
or UO_306 (O_306,N_2886,N_2623);
and UO_307 (O_307,N_2965,N_2656);
xor UO_308 (O_308,N_2527,N_2591);
nor UO_309 (O_309,N_2888,N_2700);
or UO_310 (O_310,N_2734,N_2792);
or UO_311 (O_311,N_2513,N_2503);
nor UO_312 (O_312,N_2667,N_2757);
nand UO_313 (O_313,N_2989,N_2959);
nand UO_314 (O_314,N_2782,N_2505);
or UO_315 (O_315,N_2732,N_2887);
nor UO_316 (O_316,N_2791,N_2530);
nor UO_317 (O_317,N_2781,N_2752);
or UO_318 (O_318,N_2745,N_2604);
or UO_319 (O_319,N_2632,N_2630);
nor UO_320 (O_320,N_2711,N_2961);
and UO_321 (O_321,N_2590,N_2785);
or UO_322 (O_322,N_2733,N_2627);
nand UO_323 (O_323,N_2744,N_2569);
nand UO_324 (O_324,N_2516,N_2689);
nand UO_325 (O_325,N_2606,N_2789);
nand UO_326 (O_326,N_2534,N_2607);
xor UO_327 (O_327,N_2664,N_2882);
and UO_328 (O_328,N_2542,N_2777);
nor UO_329 (O_329,N_2921,N_2600);
nand UO_330 (O_330,N_2738,N_2810);
nor UO_331 (O_331,N_2509,N_2992);
or UO_332 (O_332,N_2781,N_2547);
nor UO_333 (O_333,N_2846,N_2746);
or UO_334 (O_334,N_2695,N_2860);
nand UO_335 (O_335,N_2948,N_2822);
xnor UO_336 (O_336,N_2822,N_2533);
and UO_337 (O_337,N_2554,N_2796);
or UO_338 (O_338,N_2520,N_2866);
or UO_339 (O_339,N_2537,N_2648);
nand UO_340 (O_340,N_2763,N_2519);
or UO_341 (O_341,N_2616,N_2545);
and UO_342 (O_342,N_2560,N_2718);
or UO_343 (O_343,N_2728,N_2618);
xor UO_344 (O_344,N_2979,N_2707);
or UO_345 (O_345,N_2994,N_2772);
nor UO_346 (O_346,N_2868,N_2646);
and UO_347 (O_347,N_2594,N_2801);
nor UO_348 (O_348,N_2905,N_2535);
nand UO_349 (O_349,N_2898,N_2963);
nand UO_350 (O_350,N_2644,N_2706);
or UO_351 (O_351,N_2628,N_2905);
and UO_352 (O_352,N_2562,N_2978);
or UO_353 (O_353,N_2911,N_2585);
and UO_354 (O_354,N_2715,N_2741);
xor UO_355 (O_355,N_2728,N_2868);
and UO_356 (O_356,N_2638,N_2550);
nand UO_357 (O_357,N_2820,N_2879);
nor UO_358 (O_358,N_2885,N_2505);
nor UO_359 (O_359,N_2582,N_2579);
or UO_360 (O_360,N_2997,N_2740);
nor UO_361 (O_361,N_2919,N_2736);
nor UO_362 (O_362,N_2563,N_2577);
nor UO_363 (O_363,N_2636,N_2681);
nor UO_364 (O_364,N_2914,N_2658);
nor UO_365 (O_365,N_2638,N_2609);
or UO_366 (O_366,N_2572,N_2932);
nand UO_367 (O_367,N_2794,N_2753);
and UO_368 (O_368,N_2712,N_2694);
nor UO_369 (O_369,N_2622,N_2638);
nand UO_370 (O_370,N_2698,N_2578);
nor UO_371 (O_371,N_2660,N_2504);
or UO_372 (O_372,N_2556,N_2702);
and UO_373 (O_373,N_2732,N_2906);
nand UO_374 (O_374,N_2513,N_2881);
nand UO_375 (O_375,N_2817,N_2795);
nor UO_376 (O_376,N_2578,N_2914);
or UO_377 (O_377,N_2662,N_2914);
and UO_378 (O_378,N_2732,N_2862);
and UO_379 (O_379,N_2878,N_2960);
and UO_380 (O_380,N_2805,N_2513);
or UO_381 (O_381,N_2759,N_2533);
nand UO_382 (O_382,N_2546,N_2692);
nor UO_383 (O_383,N_2717,N_2881);
or UO_384 (O_384,N_2690,N_2751);
and UO_385 (O_385,N_2741,N_2699);
nor UO_386 (O_386,N_2952,N_2720);
or UO_387 (O_387,N_2836,N_2791);
nor UO_388 (O_388,N_2612,N_2947);
nor UO_389 (O_389,N_2941,N_2682);
nor UO_390 (O_390,N_2771,N_2908);
and UO_391 (O_391,N_2753,N_2752);
nand UO_392 (O_392,N_2876,N_2738);
nand UO_393 (O_393,N_2632,N_2811);
nor UO_394 (O_394,N_2501,N_2551);
nor UO_395 (O_395,N_2553,N_2506);
and UO_396 (O_396,N_2907,N_2779);
nor UO_397 (O_397,N_2597,N_2603);
or UO_398 (O_398,N_2800,N_2577);
or UO_399 (O_399,N_2846,N_2853);
and UO_400 (O_400,N_2506,N_2672);
or UO_401 (O_401,N_2926,N_2575);
nor UO_402 (O_402,N_2945,N_2628);
nor UO_403 (O_403,N_2674,N_2640);
or UO_404 (O_404,N_2804,N_2715);
and UO_405 (O_405,N_2949,N_2922);
nand UO_406 (O_406,N_2711,N_2712);
and UO_407 (O_407,N_2644,N_2963);
nand UO_408 (O_408,N_2637,N_2580);
nand UO_409 (O_409,N_2878,N_2584);
and UO_410 (O_410,N_2826,N_2503);
nor UO_411 (O_411,N_2805,N_2610);
nor UO_412 (O_412,N_2697,N_2642);
nor UO_413 (O_413,N_2743,N_2765);
or UO_414 (O_414,N_2799,N_2896);
and UO_415 (O_415,N_2767,N_2995);
or UO_416 (O_416,N_2582,N_2872);
or UO_417 (O_417,N_2718,N_2648);
nand UO_418 (O_418,N_2567,N_2634);
nor UO_419 (O_419,N_2710,N_2933);
or UO_420 (O_420,N_2940,N_2864);
xnor UO_421 (O_421,N_2732,N_2528);
or UO_422 (O_422,N_2985,N_2769);
xor UO_423 (O_423,N_2603,N_2652);
or UO_424 (O_424,N_2585,N_2915);
nor UO_425 (O_425,N_2942,N_2880);
nand UO_426 (O_426,N_2695,N_2989);
nor UO_427 (O_427,N_2680,N_2944);
and UO_428 (O_428,N_2696,N_2587);
nand UO_429 (O_429,N_2868,N_2866);
and UO_430 (O_430,N_2594,N_2836);
and UO_431 (O_431,N_2934,N_2835);
and UO_432 (O_432,N_2955,N_2754);
and UO_433 (O_433,N_2824,N_2573);
nand UO_434 (O_434,N_2725,N_2950);
or UO_435 (O_435,N_2513,N_2674);
or UO_436 (O_436,N_2880,N_2780);
or UO_437 (O_437,N_2820,N_2976);
or UO_438 (O_438,N_2859,N_2843);
and UO_439 (O_439,N_2982,N_2608);
or UO_440 (O_440,N_2954,N_2857);
nor UO_441 (O_441,N_2642,N_2824);
or UO_442 (O_442,N_2689,N_2572);
and UO_443 (O_443,N_2847,N_2648);
and UO_444 (O_444,N_2711,N_2642);
nor UO_445 (O_445,N_2501,N_2939);
or UO_446 (O_446,N_2895,N_2963);
or UO_447 (O_447,N_2612,N_2927);
or UO_448 (O_448,N_2515,N_2689);
nand UO_449 (O_449,N_2696,N_2512);
and UO_450 (O_450,N_2626,N_2592);
or UO_451 (O_451,N_2650,N_2742);
nor UO_452 (O_452,N_2817,N_2762);
and UO_453 (O_453,N_2540,N_2510);
nor UO_454 (O_454,N_2721,N_2595);
nor UO_455 (O_455,N_2638,N_2940);
or UO_456 (O_456,N_2859,N_2805);
and UO_457 (O_457,N_2876,N_2933);
nand UO_458 (O_458,N_2792,N_2775);
or UO_459 (O_459,N_2718,N_2988);
and UO_460 (O_460,N_2833,N_2639);
nand UO_461 (O_461,N_2544,N_2583);
or UO_462 (O_462,N_2779,N_2849);
or UO_463 (O_463,N_2534,N_2603);
nand UO_464 (O_464,N_2513,N_2574);
and UO_465 (O_465,N_2671,N_2536);
or UO_466 (O_466,N_2793,N_2591);
nor UO_467 (O_467,N_2589,N_2793);
nor UO_468 (O_468,N_2623,N_2855);
and UO_469 (O_469,N_2778,N_2502);
and UO_470 (O_470,N_2574,N_2768);
or UO_471 (O_471,N_2922,N_2824);
nor UO_472 (O_472,N_2753,N_2908);
and UO_473 (O_473,N_2617,N_2934);
nor UO_474 (O_474,N_2715,N_2711);
and UO_475 (O_475,N_2806,N_2859);
nand UO_476 (O_476,N_2656,N_2648);
or UO_477 (O_477,N_2883,N_2588);
nand UO_478 (O_478,N_2512,N_2825);
nand UO_479 (O_479,N_2911,N_2874);
or UO_480 (O_480,N_2831,N_2755);
or UO_481 (O_481,N_2878,N_2709);
or UO_482 (O_482,N_2883,N_2524);
nand UO_483 (O_483,N_2606,N_2593);
and UO_484 (O_484,N_2695,N_2740);
nor UO_485 (O_485,N_2758,N_2946);
nor UO_486 (O_486,N_2825,N_2557);
nand UO_487 (O_487,N_2721,N_2711);
nand UO_488 (O_488,N_2767,N_2501);
nand UO_489 (O_489,N_2972,N_2732);
nand UO_490 (O_490,N_2980,N_2677);
nand UO_491 (O_491,N_2698,N_2713);
and UO_492 (O_492,N_2842,N_2749);
and UO_493 (O_493,N_2692,N_2523);
nand UO_494 (O_494,N_2935,N_2520);
nand UO_495 (O_495,N_2523,N_2789);
nor UO_496 (O_496,N_2871,N_2893);
nand UO_497 (O_497,N_2859,N_2711);
nor UO_498 (O_498,N_2607,N_2871);
xnor UO_499 (O_499,N_2944,N_2520);
endmodule