module basic_1500_15000_2000_20_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
and U0 (N_0,In_482,In_699);
or U1 (N_1,In_1222,In_192);
nand U2 (N_2,In_458,In_323);
xor U3 (N_3,In_606,In_655);
and U4 (N_4,In_101,In_940);
nand U5 (N_5,In_1106,In_598);
xnor U6 (N_6,In_1048,In_1346);
xor U7 (N_7,In_1432,In_924);
and U8 (N_8,In_1399,In_232);
nor U9 (N_9,In_1219,In_823);
or U10 (N_10,In_736,In_28);
nor U11 (N_11,In_1333,In_202);
or U12 (N_12,In_1436,In_3);
or U13 (N_13,In_480,In_949);
or U14 (N_14,In_1282,In_463);
or U15 (N_15,In_399,In_1166);
nor U16 (N_16,In_1255,In_631);
xor U17 (N_17,In_1110,In_1138);
nor U18 (N_18,In_14,In_1074);
xnor U19 (N_19,In_967,In_899);
nand U20 (N_20,In_1189,In_607);
nor U21 (N_21,In_617,In_793);
nor U22 (N_22,In_682,In_853);
nand U23 (N_23,In_544,In_389);
or U24 (N_24,In_1190,In_1331);
and U25 (N_25,In_444,In_415);
nor U26 (N_26,In_918,In_1366);
nor U27 (N_27,In_983,In_107);
nor U28 (N_28,In_720,In_417);
xnor U29 (N_29,In_751,In_223);
nand U30 (N_30,In_85,In_669);
nand U31 (N_31,In_622,In_260);
nand U32 (N_32,In_1414,In_222);
and U33 (N_33,In_718,In_1152);
and U34 (N_34,In_987,In_1443);
nand U35 (N_35,In_973,In_1373);
or U36 (N_36,In_1266,In_476);
nand U37 (N_37,In_1109,In_1306);
and U38 (N_38,In_186,In_836);
nor U39 (N_39,In_840,In_339);
or U40 (N_40,In_795,In_1481);
nand U41 (N_41,In_1176,In_1003);
or U42 (N_42,In_1403,In_882);
nand U43 (N_43,In_1288,In_52);
nand U44 (N_44,In_988,In_997);
nor U45 (N_45,In_818,In_861);
or U46 (N_46,In_250,In_198);
nor U47 (N_47,In_1320,In_21);
xnor U48 (N_48,In_262,In_938);
or U49 (N_49,In_128,In_602);
xor U50 (N_50,In_1238,In_568);
or U51 (N_51,In_91,In_756);
nor U52 (N_52,In_98,In_303);
or U53 (N_53,In_584,In_1398);
nor U54 (N_54,In_75,In_1465);
or U55 (N_55,In_204,In_541);
xnor U56 (N_56,In_1305,In_1204);
and U57 (N_57,In_1397,In_182);
nand U58 (N_58,In_764,In_230);
or U59 (N_59,In_167,In_134);
or U60 (N_60,In_800,In_1224);
nor U61 (N_61,In_935,In_299);
and U62 (N_62,In_1000,In_1364);
nand U63 (N_63,In_1310,In_445);
and U64 (N_64,In_760,In_958);
nor U65 (N_65,In_583,In_707);
nor U66 (N_66,In_995,In_290);
and U67 (N_67,In_1066,In_252);
xnor U68 (N_68,In_1335,In_99);
nor U69 (N_69,In_5,In_1326);
nor U70 (N_70,In_833,In_1108);
xor U71 (N_71,In_542,In_1495);
and U72 (N_72,In_1134,In_1304);
and U73 (N_73,In_1265,In_535);
and U74 (N_74,In_670,In_636);
nand U75 (N_75,In_1328,In_275);
or U76 (N_76,In_126,In_742);
and U77 (N_77,In_272,In_708);
nor U78 (N_78,In_559,In_891);
nand U79 (N_79,In_1433,In_928);
or U80 (N_80,In_520,In_100);
and U81 (N_81,In_828,In_672);
and U82 (N_82,In_214,In_454);
xnor U83 (N_83,In_306,In_730);
and U84 (N_84,In_1118,In_1478);
or U85 (N_85,In_1231,In_1389);
nor U86 (N_86,In_845,In_379);
or U87 (N_87,In_336,In_1269);
nand U88 (N_88,In_436,In_337);
and U89 (N_89,In_917,In_439);
xnor U90 (N_90,In_1124,In_1);
or U91 (N_91,In_936,In_1182);
and U92 (N_92,In_572,In_733);
nor U93 (N_93,In_1390,In_452);
or U94 (N_94,In_150,In_1498);
nand U95 (N_95,In_407,In_1327);
nor U96 (N_96,In_660,In_1466);
and U97 (N_97,In_525,In_1216);
xor U98 (N_98,In_16,In_194);
and U99 (N_99,In_221,In_191);
and U100 (N_100,In_470,In_772);
and U101 (N_101,In_780,In_1160);
xnor U102 (N_102,In_560,In_1242);
xor U103 (N_103,In_1289,In_1484);
nand U104 (N_104,In_693,In_355);
or U105 (N_105,In_239,In_685);
and U106 (N_106,In_69,In_59);
xnor U107 (N_107,In_1139,In_634);
and U108 (N_108,In_29,In_295);
and U109 (N_109,In_589,In_748);
nand U110 (N_110,In_1451,In_1161);
nand U111 (N_111,In_26,In_130);
nand U112 (N_112,In_757,In_1114);
or U113 (N_113,In_1345,In_383);
nor U114 (N_114,In_15,In_1344);
nand U115 (N_115,In_618,In_969);
nor U116 (N_116,In_428,In_1301);
nor U117 (N_117,In_719,In_803);
nor U118 (N_118,In_1019,In_785);
nand U119 (N_119,In_856,In_1240);
or U120 (N_120,In_243,In_276);
nand U121 (N_121,In_207,In_1375);
nor U122 (N_122,In_1386,In_1130);
nor U123 (N_123,In_249,In_448);
nor U124 (N_124,In_479,In_145);
nand U125 (N_125,In_673,In_1428);
and U126 (N_126,In_909,In_13);
or U127 (N_127,In_373,In_846);
nor U128 (N_128,In_1449,In_284);
xor U129 (N_129,In_1281,In_1084);
or U130 (N_130,In_1332,In_787);
and U131 (N_131,In_1150,In_1214);
or U132 (N_132,In_1351,In_279);
nor U133 (N_133,In_11,In_906);
or U134 (N_134,In_1181,In_540);
or U135 (N_135,In_644,In_131);
xnor U136 (N_136,In_521,In_885);
xnor U137 (N_137,In_380,In_574);
and U138 (N_138,In_531,In_1058);
nand U139 (N_139,In_226,In_1378);
nand U140 (N_140,In_73,In_97);
nor U141 (N_141,In_1250,In_1025);
xor U142 (N_142,In_61,In_653);
nor U143 (N_143,In_976,In_1232);
and U144 (N_144,In_913,In_791);
nand U145 (N_145,In_1452,In_1081);
nor U146 (N_146,In_985,In_60);
or U147 (N_147,In_512,In_273);
or U148 (N_148,In_1268,In_608);
xor U149 (N_149,In_922,In_1086);
nor U150 (N_150,In_446,In_316);
or U151 (N_151,In_370,In_1413);
nand U152 (N_152,In_1491,In_705);
or U153 (N_153,In_674,In_318);
xor U154 (N_154,In_1132,In_132);
nor U155 (N_155,In_44,In_907);
nand U156 (N_156,In_175,In_650);
nor U157 (N_157,In_286,In_478);
xor U158 (N_158,In_1294,In_633);
xor U159 (N_159,In_713,In_986);
and U160 (N_160,In_263,In_1317);
nand U161 (N_161,In_630,In_1402);
and U162 (N_162,In_1278,In_1051);
nor U163 (N_163,In_364,In_140);
or U164 (N_164,In_962,In_1434);
or U165 (N_165,In_582,In_768);
or U166 (N_166,In_1133,In_1361);
nand U167 (N_167,In_1087,In_806);
or U168 (N_168,In_530,In_504);
nor U169 (N_169,In_663,In_1370);
or U170 (N_170,In_597,In_1191);
nor U171 (N_171,In_819,In_624);
nand U172 (N_172,In_1226,In_36);
xor U173 (N_173,In_409,In_950);
nand U174 (N_174,In_765,In_556);
and U175 (N_175,In_683,In_1239);
or U176 (N_176,In_159,In_83);
nand U177 (N_177,In_895,In_1492);
xor U178 (N_178,In_205,In_702);
or U179 (N_179,In_112,In_1355);
and U180 (N_180,In_942,In_627);
or U181 (N_181,In_166,In_511);
nand U182 (N_182,In_1448,In_543);
or U183 (N_183,In_1485,In_300);
xor U184 (N_184,In_1196,In_999);
nor U185 (N_185,In_93,In_340);
and U186 (N_186,In_488,In_1356);
xor U187 (N_187,In_1046,In_966);
nand U188 (N_188,In_1392,In_1274);
or U189 (N_189,In_536,In_578);
xor U190 (N_190,In_516,In_697);
or U191 (N_191,In_956,In_657);
or U192 (N_192,In_255,In_392);
nor U193 (N_193,In_1153,In_125);
or U194 (N_194,In_643,In_884);
and U195 (N_195,In_947,In_731);
or U196 (N_196,In_430,In_1312);
and U197 (N_197,In_1168,In_1243);
nand U198 (N_198,In_518,In_1263);
and U199 (N_199,In_1457,In_844);
and U200 (N_200,In_527,In_359);
xor U201 (N_201,In_197,In_94);
nor U202 (N_202,In_798,In_157);
xnor U203 (N_203,In_700,In_441);
and U204 (N_204,In_502,In_203);
nor U205 (N_205,In_331,In_473);
xnor U206 (N_206,In_40,In_408);
and U207 (N_207,In_839,In_244);
and U208 (N_208,In_1468,In_1050);
nand U209 (N_209,In_301,In_570);
nand U210 (N_210,In_320,In_1163);
or U211 (N_211,In_309,In_465);
or U212 (N_212,In_442,In_837);
xor U213 (N_213,In_941,In_858);
nor U214 (N_214,In_121,In_782);
xor U215 (N_215,In_1387,In_790);
or U216 (N_216,In_1273,In_304);
and U217 (N_217,In_1447,In_971);
xor U218 (N_218,In_1032,In_1444);
nor U219 (N_219,In_163,In_522);
nand U220 (N_220,In_783,In_176);
xor U221 (N_221,In_1143,In_1127);
nand U222 (N_222,In_857,In_737);
or U223 (N_223,In_208,In_1302);
nor U224 (N_224,In_1353,In_654);
nor U225 (N_225,In_691,In_240);
xor U226 (N_226,In_665,In_57);
nand U227 (N_227,In_330,In_362);
nand U228 (N_228,In_546,In_868);
xnor U229 (N_229,In_1029,In_1494);
nor U230 (N_230,In_398,In_241);
xor U231 (N_231,In_538,In_614);
nor U232 (N_232,In_460,In_1102);
nor U233 (N_233,In_396,In_804);
and U234 (N_234,In_789,In_174);
nor U235 (N_235,In_9,In_348);
nand U236 (N_236,In_964,In_490);
nand U237 (N_237,In_1094,In_802);
or U238 (N_238,In_646,In_84);
and U239 (N_239,In_573,In_1264);
and U240 (N_240,In_886,In_977);
nor U241 (N_241,In_686,In_1195);
xor U242 (N_242,In_338,In_1069);
and U243 (N_243,In_1194,In_509);
and U244 (N_244,In_600,In_280);
or U245 (N_245,In_270,In_1441);
or U246 (N_246,In_1169,In_1272);
and U247 (N_247,In_137,In_327);
nor U248 (N_248,In_1121,In_228);
xor U249 (N_249,In_1296,In_218);
xnor U250 (N_250,In_1128,In_829);
and U251 (N_251,In_952,In_1340);
or U252 (N_252,In_1417,In_55);
or U253 (N_253,In_943,In_1343);
xor U254 (N_254,In_1082,In_1091);
nor U255 (N_255,In_7,In_177);
and U256 (N_256,In_1024,In_1453);
or U257 (N_257,In_4,In_1093);
and U258 (N_258,In_755,In_824);
or U259 (N_259,In_1309,In_659);
nand U260 (N_260,In_1446,In_92);
xor U261 (N_261,In_854,In_1313);
xnor U262 (N_262,In_813,In_210);
and U263 (N_263,In_30,In_1475);
nor U264 (N_264,In_491,In_638);
and U265 (N_265,In_1275,In_1077);
nor U266 (N_266,In_1499,In_1419);
nand U267 (N_267,In_403,In_213);
or U268 (N_268,In_1183,In_763);
or U269 (N_269,In_124,In_767);
and U270 (N_270,In_179,In_1290);
xnor U271 (N_271,In_248,In_1007);
or U272 (N_272,In_413,In_265);
and U273 (N_273,In_576,In_1113);
or U274 (N_274,In_1096,In_1371);
or U275 (N_275,In_732,In_388);
nor U276 (N_276,In_78,In_225);
or U277 (N_277,In_1440,In_571);
nor U278 (N_278,In_443,In_1173);
nor U279 (N_279,In_1103,In_189);
nand U280 (N_280,In_1119,In_314);
or U281 (N_281,In_387,In_497);
nor U282 (N_282,In_1473,In_877);
or U283 (N_283,In_120,In_164);
nor U284 (N_284,In_305,In_524);
and U285 (N_285,In_1365,In_440);
or U286 (N_286,In_48,In_165);
and U287 (N_287,In_489,In_54);
nand U288 (N_288,In_896,In_1225);
and U289 (N_289,In_492,In_661);
nand U290 (N_290,In_462,In_1111);
xor U291 (N_291,In_784,In_1089);
xnor U292 (N_292,In_1394,In_515);
nor U293 (N_293,In_135,In_1013);
nor U294 (N_294,In_1076,In_822);
nor U295 (N_295,In_860,In_507);
nor U296 (N_296,In_25,In_158);
and U297 (N_297,In_1405,In_1396);
nand U298 (N_298,In_1129,In_1197);
nand U299 (N_299,In_1164,In_212);
nand U300 (N_300,In_1229,In_1431);
or U301 (N_301,In_1249,In_1022);
nor U302 (N_302,In_1159,In_549);
nand U303 (N_303,In_1360,In_698);
nand U304 (N_304,In_209,In_1459);
nand U305 (N_305,In_1385,In_266);
and U306 (N_306,In_914,In_1410);
xor U307 (N_307,In_168,In_623);
xnor U308 (N_308,In_1271,In_1324);
nand U309 (N_309,In_769,In_741);
xor U310 (N_310,In_471,In_1174);
and U311 (N_311,In_668,In_1137);
or U312 (N_312,In_236,In_775);
nor U313 (N_313,In_1206,In_781);
nand U314 (N_314,In_122,In_1262);
or U315 (N_315,In_1064,In_905);
nand U316 (N_316,In_561,In_395);
nor U317 (N_317,In_196,In_1252);
nand U318 (N_318,In_103,In_1049);
nor U319 (N_319,In_1101,In_715);
nand U320 (N_320,In_172,In_678);
or U321 (N_321,In_495,In_1020);
xor U322 (N_322,In_153,In_483);
and U323 (N_323,In_838,In_827);
nor U324 (N_324,In_1338,In_1208);
xor U325 (N_325,In_567,In_351);
or U326 (N_326,In_1329,In_24);
xor U327 (N_327,In_1071,In_423);
nor U328 (N_328,In_1053,In_350);
and U329 (N_329,In_1415,In_19);
or U330 (N_330,In_1199,In_506);
xnor U331 (N_331,In_894,In_1001);
or U332 (N_332,In_467,In_345);
xnor U333 (N_333,In_363,In_863);
and U334 (N_334,In_1186,In_960);
or U335 (N_335,In_1156,In_777);
nand U336 (N_336,In_310,In_902);
nand U337 (N_337,In_1455,In_1471);
and U338 (N_338,In_1162,In_1055);
and U339 (N_339,In_1435,In_711);
xnor U340 (N_340,In_325,In_2);
xnor U341 (N_341,In_499,In_927);
or U342 (N_342,In_1154,In_173);
or U343 (N_343,In_1456,In_1472);
nand U344 (N_344,In_1052,In_1057);
and U345 (N_345,In_1292,In_105);
nand U346 (N_346,In_770,In_981);
nand U347 (N_347,In_820,In_369);
and U348 (N_348,In_365,In_215);
or U349 (N_349,In_752,In_1337);
nor U350 (N_350,In_461,In_817);
and U351 (N_351,In_133,In_911);
or U352 (N_352,In_593,In_948);
xnor U353 (N_353,In_539,In_1223);
and U354 (N_354,In_689,In_779);
or U355 (N_355,In_859,In_1234);
xnor U356 (N_356,In_464,In_621);
and U357 (N_357,In_455,In_206);
or U358 (N_358,In_487,In_450);
nor U359 (N_359,In_919,In_493);
and U360 (N_360,In_712,In_356);
or U361 (N_361,In_587,In_88);
or U362 (N_362,In_1438,In_420);
xnor U363 (N_363,In_1044,In_537);
or U364 (N_364,In_302,In_469);
nor U365 (N_365,In_151,In_613);
xnor U366 (N_366,In_1170,In_1388);
nor U367 (N_367,In_1316,In_288);
nor U368 (N_368,In_1145,In_475);
nand U369 (N_369,In_216,In_968);
nor U370 (N_370,In_271,In_1270);
xor U371 (N_371,In_904,In_852);
xor U372 (N_372,In_994,In_1303);
or U373 (N_373,In_1008,In_34);
and U374 (N_374,In_550,In_1033);
nand U375 (N_375,In_1318,In_1072);
and U376 (N_376,In_890,In_727);
nand U377 (N_377,In_372,In_378);
nor U378 (N_378,In_610,In_217);
xor U379 (N_379,In_1464,In_1314);
and U380 (N_380,In_897,In_1136);
xnor U381 (N_381,In_662,In_677);
nand U382 (N_382,In_1251,In_1241);
or U383 (N_383,In_1348,In_869);
and U384 (N_384,In_706,In_1235);
and U385 (N_385,In_998,In_1477);
xnor U386 (N_386,In_447,In_119);
and U387 (N_387,In_1259,In_346);
and U388 (N_388,In_709,In_514);
and U389 (N_389,In_315,In_332);
xor U390 (N_390,In_235,In_1015);
nor U391 (N_391,In_557,In_1401);
and U392 (N_392,In_933,In_234);
nand U393 (N_393,In_811,In_810);
nand U394 (N_394,In_82,In_776);
nor U395 (N_395,In_1165,In_1233);
nand U396 (N_396,In_1247,In_70);
xnor U397 (N_397,In_23,In_426);
and U398 (N_398,In_666,In_1230);
or U399 (N_399,In_552,In_797);
and U400 (N_400,In_20,In_865);
and U401 (N_401,In_1178,In_625);
nor U402 (N_402,In_590,In_558);
nor U403 (N_403,In_116,In_190);
or U404 (N_404,In_429,In_1209);
nand U405 (N_405,In_1404,In_1253);
or U406 (N_406,In_1146,In_594);
nor U407 (N_407,In_843,In_771);
xor U408 (N_408,In_1228,In_1285);
and U409 (N_409,In_1227,In_67);
nor U410 (N_410,In_89,In_519);
nor U411 (N_411,In_642,In_451);
xnor U412 (N_412,In_115,In_626);
or U413 (N_413,In_898,In_1424);
nand U414 (N_414,In_805,In_438);
xor U415 (N_415,In_1104,In_269);
or U416 (N_416,In_1377,In_146);
nand U417 (N_417,In_1418,In_274);
nor U418 (N_418,In_71,In_658);
nor U419 (N_419,In_242,In_1040);
xor U420 (N_420,In_1042,In_915);
or U421 (N_421,In_1379,In_1490);
nor U422 (N_422,In_901,In_548);
xnor U423 (N_423,In_246,In_889);
and U424 (N_424,In_384,In_750);
xor U425 (N_425,In_1372,In_993);
nor U426 (N_426,In_433,In_611);
nand U427 (N_427,In_321,In_1244);
nor U428 (N_428,In_1427,In_1256);
or U429 (N_429,In_377,In_866);
xor U430 (N_430,In_1261,In_291);
and U431 (N_431,In_457,In_932);
nand U432 (N_432,In_199,In_910);
and U433 (N_433,In_601,In_1210);
nand U434 (N_434,In_652,In_569);
nor U435 (N_435,In_1157,In_996);
xor U436 (N_436,In_141,In_357);
or U437 (N_437,In_687,In_864);
xor U438 (N_438,In_870,In_411);
or U439 (N_439,In_888,In_435);
and U440 (N_440,In_788,In_1442);
or U441 (N_441,In_1085,In_334);
nor U442 (N_442,In_22,In_1423);
xnor U443 (N_443,In_466,In_1488);
and U444 (N_444,In_841,In_76);
and U445 (N_445,In_812,In_0);
nor U446 (N_446,In_233,In_1391);
xnor U447 (N_447,In_1167,In_908);
and U448 (N_448,In_312,In_1445);
nor U449 (N_449,In_148,In_679);
or U450 (N_450,In_1339,In_1382);
and U451 (N_451,In_1158,In_595);
or U452 (N_452,In_688,In_343);
or U453 (N_453,In_287,In_1062);
and U454 (N_454,In_1358,In_825);
xnor U455 (N_455,In_1131,In_529);
xnor U456 (N_456,In_1116,In_219);
nand U457 (N_457,In_503,In_1286);
xor U458 (N_458,In_1437,In_1115);
and U459 (N_459,In_1407,In_612);
nor U460 (N_460,In_1347,In_875);
and U461 (N_461,In_1205,In_39);
xor U462 (N_462,In_835,In_201);
xor U463 (N_463,In_188,In_974);
and U464 (N_464,In_1011,In_562);
xnor U465 (N_465,In_628,In_358);
or U466 (N_466,In_1267,In_386);
nor U467 (N_467,In_1034,In_1039);
and U468 (N_468,In_79,In_645);
or U469 (N_469,In_934,In_459);
xor U470 (N_470,In_245,In_496);
nor U471 (N_471,In_110,In_1080);
nand U472 (N_472,In_566,In_6);
nor U473 (N_473,In_294,In_640);
and U474 (N_474,In_526,In_575);
and U475 (N_475,In_1036,In_1248);
nand U476 (N_476,In_296,In_1421);
nor U477 (N_477,In_410,In_424);
nand U478 (N_478,In_1175,In_978);
xnor U479 (N_479,In_390,In_937);
nand U480 (N_480,In_807,In_912);
xnor U481 (N_481,In_1321,In_326);
and U482 (N_482,In_1357,In_1381);
nand U483 (N_483,In_56,In_1097);
xnor U484 (N_484,In_1212,In_1350);
xnor U485 (N_485,In_1349,In_809);
nor U486 (N_486,In_258,In_1454);
nand U487 (N_487,In_1125,In_449);
and U488 (N_488,In_283,In_38);
and U489 (N_489,In_874,In_778);
xor U490 (N_490,In_903,In_726);
nand U491 (N_491,In_1079,In_1211);
or U492 (N_492,In_1151,In_375);
nand U493 (N_493,In_8,In_849);
and U494 (N_494,In_961,In_106);
xor U495 (N_495,In_425,In_847);
or U496 (N_496,In_183,In_1469);
and U497 (N_497,In_412,In_171);
or U498 (N_498,In_231,In_74);
nor U499 (N_499,In_1009,In_1218);
nor U500 (N_500,In_794,In_616);
or U501 (N_501,In_421,In_494);
nor U502 (N_502,In_344,In_629);
nor U503 (N_503,In_238,In_501);
and U504 (N_504,In_746,In_739);
xnor U505 (N_505,In_729,In_563);
nand U506 (N_506,In_1018,In_1461);
xor U507 (N_507,In_1179,In_955);
nor U508 (N_508,In_523,In_1245);
and U509 (N_509,In_588,In_268);
xnor U510 (N_510,In_1412,In_1221);
nand U511 (N_511,In_477,In_152);
nand U512 (N_512,In_17,In_615);
nor U513 (N_513,In_508,In_1439);
nor U514 (N_514,In_254,In_366);
nor U515 (N_515,In_592,In_329);
or U516 (N_516,In_65,In_160);
nor U517 (N_517,In_871,In_872);
nor U518 (N_518,In_80,In_714);
and U519 (N_519,In_35,In_1400);
nand U520 (N_520,In_322,In_484);
and U521 (N_521,In_1458,In_367);
or U522 (N_522,In_1023,In_311);
nor U523 (N_523,In_1254,In_347);
nand U524 (N_524,In_81,In_1016);
and U525 (N_525,In_251,In_123);
nand U526 (N_526,In_277,In_970);
nand U527 (N_527,In_1192,In_391);
and U528 (N_528,In_639,In_51);
or U529 (N_529,In_635,In_814);
or U530 (N_530,In_808,In_127);
nand U531 (N_531,In_1148,In_887);
or U532 (N_532,In_1393,In_418);
and U533 (N_533,In_1482,In_144);
and U534 (N_534,In_1330,In_1470);
nand U535 (N_535,In_1200,In_1140);
or U536 (N_536,In_975,In_278);
nand U537 (N_537,In_1284,In_1429);
and U538 (N_538,In_1369,In_1298);
and U539 (N_539,In_754,In_565);
or U540 (N_540,In_1277,In_1107);
and U541 (N_541,In_930,In_257);
or U542 (N_542,In_187,In_114);
nand U543 (N_543,In_63,In_945);
xnor U544 (N_544,In_647,In_848);
xor U545 (N_545,In_883,In_1342);
and U546 (N_546,In_551,In_282);
and U547 (N_547,In_799,In_842);
nand U548 (N_548,In_341,In_113);
xor U549 (N_549,In_1213,In_354);
nand U550 (N_550,In_66,In_18);
nand U551 (N_551,In_850,In_1246);
and U552 (N_552,In_43,In_786);
or U553 (N_553,In_517,In_432);
and U554 (N_554,In_1004,In_892);
and U555 (N_555,In_500,In_1217);
and U556 (N_556,In_528,In_1406);
or U557 (N_557,In_1100,In_723);
nand U558 (N_558,In_1188,In_87);
or U559 (N_559,In_142,In_876);
or U560 (N_560,In_599,In_1352);
or U561 (N_561,In_603,In_1493);
and U562 (N_562,In_72,In_696);
nand U563 (N_563,In_564,In_1319);
nand U564 (N_564,In_37,In_1430);
or U565 (N_565,In_716,In_1038);
nor U566 (N_566,In_664,In_703);
nand U567 (N_567,In_1293,In_402);
xor U568 (N_568,In_1368,In_86);
xor U569 (N_569,In_481,In_1460);
nor U570 (N_570,In_979,In_1047);
nor U571 (N_571,In_297,In_1300);
and U572 (N_572,In_1483,In_931);
xor U573 (N_573,In_437,In_1476);
nor U574 (N_574,In_1450,In_200);
xnor U575 (N_575,In_900,In_247);
and U576 (N_576,In_32,In_267);
nor U577 (N_577,In_62,In_1341);
or U578 (N_578,In_796,In_831);
nand U579 (N_579,In_1276,In_939);
nor U580 (N_580,In_1287,In_1122);
nand U581 (N_581,In_1060,In_743);
xnor U582 (N_582,In_1180,In_342);
or U583 (N_583,In_138,In_281);
nand U584 (N_584,In_102,In_701);
xor U585 (N_585,In_944,In_879);
or U586 (N_586,In_256,In_609);
and U587 (N_587,In_434,In_361);
and U588 (N_588,In_534,In_1202);
and U589 (N_589,In_761,In_547);
xor U590 (N_590,In_953,In_585);
nand U591 (N_591,In_880,In_989);
or U592 (N_592,In_64,In_376);
or U593 (N_593,In_992,In_619);
nand U594 (N_594,In_472,In_648);
nor U595 (N_595,In_555,In_53);
or U596 (N_596,In_1334,In_10);
nor U597 (N_597,In_946,In_990);
nor U598 (N_598,In_1063,In_1092);
nor U599 (N_599,In_1236,In_724);
nand U600 (N_600,In_710,In_725);
nand U601 (N_601,In_1408,In_1027);
nor U602 (N_602,In_129,In_1463);
or U603 (N_603,In_1384,In_1141);
and U604 (N_604,In_117,In_759);
nand U605 (N_605,In_104,In_397);
xor U606 (N_606,In_1420,In_1041);
nand U607 (N_607,In_1315,In_510);
or U608 (N_608,In_695,In_456);
and U609 (N_609,In_747,In_1257);
or U610 (N_610,In_317,In_728);
nand U611 (N_611,In_313,In_1067);
or U612 (N_612,In_1376,In_1098);
xnor U613 (N_613,In_453,In_773);
or U614 (N_614,In_758,In_984);
nand U615 (N_615,In_649,In_965);
nand U616 (N_616,In_1177,In_1367);
nand U617 (N_617,In_1155,In_972);
nor U618 (N_618,In_1322,In_1123);
and U619 (N_619,In_353,In_684);
and U620 (N_620,In_826,In_957);
or U621 (N_621,In_1487,In_285);
nand U622 (N_622,In_31,In_1083);
or U623 (N_623,In_298,In_1117);
nand U624 (N_624,In_1297,In_498);
and U625 (N_625,In_33,In_414);
xor U626 (N_626,In_744,In_405);
and U627 (N_627,In_1090,In_371);
or U628 (N_628,In_118,In_1035);
xor U629 (N_629,In_431,In_1010);
nor U630 (N_630,In_959,In_360);
nand U631 (N_631,In_505,In_1215);
or U632 (N_632,In_1031,In_416);
nand U633 (N_633,In_193,In_1354);
or U634 (N_634,In_42,In_532);
nand U635 (N_635,In_227,In_259);
xor U636 (N_636,In_333,In_1185);
nor U637 (N_637,In_1184,In_1480);
xor U638 (N_638,In_792,In_963);
xor U639 (N_639,In_162,In_1078);
nand U640 (N_640,In_155,In_139);
and U641 (N_641,In_692,In_632);
and U642 (N_642,In_136,In_154);
nor U643 (N_643,In_738,In_307);
nor U644 (N_644,In_1486,In_328);
xor U645 (N_645,In_980,In_1021);
nand U646 (N_646,In_220,In_1198);
nor U647 (N_647,In_422,In_926);
nand U648 (N_648,In_181,In_178);
and U649 (N_649,In_1005,In_766);
nand U650 (N_650,In_229,In_878);
and U651 (N_651,In_393,In_1425);
xor U652 (N_652,In_1073,In_385);
and U653 (N_653,In_1489,In_1359);
xor U654 (N_654,In_1323,In_671);
or U655 (N_655,In_195,In_382);
and U656 (N_656,In_1307,In_1207);
and U657 (N_657,In_1237,In_717);
nor U658 (N_658,In_921,In_873);
xnor U659 (N_659,In_96,In_581);
nor U660 (N_660,In_1383,In_149);
and U661 (N_661,In_1112,In_694);
or U662 (N_662,In_596,In_1380);
and U663 (N_663,In_1409,In_533);
nor U664 (N_664,In_1126,In_1362);
nand U665 (N_665,In_1054,In_308);
or U666 (N_666,In_855,In_253);
xnor U667 (N_667,In_830,In_184);
nand U668 (N_668,In_954,In_47);
nand U669 (N_669,In_50,In_762);
nor U670 (N_670,In_1014,In_468);
and U671 (N_671,In_1467,In_1193);
xor U672 (N_672,In_916,In_815);
nor U673 (N_673,In_1496,In_1043);
xnor U674 (N_674,In_925,In_293);
xor U675 (N_675,In_591,In_1336);
or U676 (N_676,In_292,In_335);
and U677 (N_677,In_394,In_90);
and U678 (N_678,In_920,In_681);
and U679 (N_679,In_1075,In_400);
or U680 (N_680,In_774,In_641);
nor U681 (N_681,In_1030,In_1006);
and U682 (N_682,In_368,In_991);
nor U683 (N_683,In_1135,In_237);
and U684 (N_684,In_1187,In_41);
xnor U685 (N_685,In_95,In_111);
or U686 (N_686,In_324,In_406);
or U687 (N_687,In_404,In_1280);
xnor U688 (N_688,In_1416,In_816);
or U689 (N_689,In_419,In_1120);
nor U690 (N_690,In_77,In_108);
nand U691 (N_691,In_951,In_734);
nor U692 (N_692,In_1065,In_722);
or U693 (N_693,In_1395,In_264);
nand U694 (N_694,In_224,In_656);
and U695 (N_695,In_1012,In_579);
nand U696 (N_696,In_1056,In_374);
or U697 (N_697,In_1061,In_1325);
nand U698 (N_698,In_801,In_1299);
nand U699 (N_699,In_1147,In_735);
or U700 (N_700,In_161,In_1422);
xor U701 (N_701,In_319,In_1295);
nand U702 (N_702,In_12,In_381);
nand U703 (N_703,In_676,In_893);
nand U704 (N_704,In_675,In_620);
and U705 (N_705,In_45,In_1144);
or U706 (N_706,In_834,In_1172);
and U707 (N_707,In_261,In_862);
or U708 (N_708,In_1149,In_553);
nor U709 (N_709,In_1203,In_1171);
nor U710 (N_710,In_580,In_604);
or U711 (N_711,In_680,In_586);
xor U712 (N_712,In_289,In_1308);
or U713 (N_713,In_821,In_401);
nand U714 (N_714,In_46,In_1479);
nand U715 (N_715,In_1142,In_867);
or U716 (N_716,In_147,In_1426);
and U717 (N_717,In_349,In_753);
xnor U718 (N_718,In_58,In_1095);
nand U719 (N_719,In_577,In_1374);
nand U720 (N_720,In_651,In_1002);
xor U721 (N_721,In_211,In_1363);
and U722 (N_722,In_1311,In_185);
xnor U723 (N_723,In_1291,In_180);
nor U724 (N_724,In_170,In_486);
or U725 (N_725,In_1070,In_169);
nand U726 (N_726,In_690,In_1017);
nand U727 (N_727,In_851,In_1258);
and U728 (N_728,In_1474,In_745);
nor U729 (N_729,In_143,In_49);
xor U730 (N_730,In_740,In_637);
or U731 (N_731,In_1497,In_667);
or U732 (N_732,In_1411,In_1068);
and U733 (N_733,In_1028,In_513);
nor U734 (N_734,In_1220,In_1099);
or U735 (N_735,In_27,In_545);
nand U736 (N_736,In_352,In_554);
and U737 (N_737,In_1462,In_923);
xor U738 (N_738,In_1059,In_485);
and U739 (N_739,In_68,In_156);
nand U740 (N_740,In_427,In_1045);
xor U741 (N_741,In_1037,In_474);
and U742 (N_742,In_929,In_1088);
and U743 (N_743,In_1201,In_605);
nand U744 (N_744,In_881,In_749);
or U745 (N_745,In_109,In_1279);
nor U746 (N_746,In_704,In_1026);
or U747 (N_747,In_1283,In_1105);
xnor U748 (N_748,In_1260,In_721);
xnor U749 (N_749,In_832,In_982);
or U750 (N_750,N_104,N_352);
nor U751 (N_751,N_651,N_165);
or U752 (N_752,N_297,N_551);
nand U753 (N_753,N_122,N_356);
nor U754 (N_754,N_686,N_484);
xor U755 (N_755,N_503,N_205);
nand U756 (N_756,N_4,N_8);
xor U757 (N_757,N_408,N_574);
nand U758 (N_758,N_79,N_101);
xor U759 (N_759,N_94,N_346);
or U760 (N_760,N_507,N_398);
xnor U761 (N_761,N_441,N_570);
or U762 (N_762,N_344,N_690);
xor U763 (N_763,N_583,N_508);
xnor U764 (N_764,N_3,N_68);
or U765 (N_765,N_34,N_232);
xnor U766 (N_766,N_440,N_279);
nand U767 (N_767,N_577,N_543);
xnor U768 (N_768,N_728,N_207);
nand U769 (N_769,N_123,N_477);
nand U770 (N_770,N_269,N_677);
and U771 (N_771,N_271,N_92);
nand U772 (N_772,N_748,N_303);
nand U773 (N_773,N_411,N_376);
nand U774 (N_774,N_709,N_304);
nand U775 (N_775,N_203,N_613);
xnor U776 (N_776,N_697,N_121);
and U777 (N_777,N_609,N_89);
or U778 (N_778,N_417,N_369);
nor U779 (N_779,N_248,N_14);
xor U780 (N_780,N_572,N_740);
xor U781 (N_781,N_505,N_40);
and U782 (N_782,N_323,N_42);
xnor U783 (N_783,N_224,N_465);
and U784 (N_784,N_612,N_11);
or U785 (N_785,N_578,N_495);
or U786 (N_786,N_448,N_559);
nand U787 (N_787,N_67,N_584);
or U788 (N_788,N_134,N_424);
nor U789 (N_789,N_245,N_145);
xnor U790 (N_790,N_679,N_227);
or U791 (N_791,N_148,N_236);
or U792 (N_792,N_235,N_418);
or U793 (N_793,N_293,N_478);
and U794 (N_794,N_514,N_288);
xnor U795 (N_795,N_317,N_394);
xnor U796 (N_796,N_19,N_568);
and U797 (N_797,N_582,N_545);
nand U798 (N_798,N_382,N_307);
or U799 (N_799,N_305,N_160);
xor U800 (N_800,N_125,N_387);
nand U801 (N_801,N_602,N_311);
nand U802 (N_802,N_729,N_180);
nand U803 (N_803,N_513,N_113);
nor U804 (N_804,N_519,N_187);
or U805 (N_805,N_206,N_381);
nor U806 (N_806,N_678,N_73);
xnor U807 (N_807,N_164,N_749);
and U808 (N_808,N_611,N_191);
or U809 (N_809,N_44,N_472);
nand U810 (N_810,N_524,N_209);
or U811 (N_811,N_357,N_5);
and U812 (N_812,N_721,N_447);
and U813 (N_813,N_174,N_727);
or U814 (N_814,N_274,N_22);
and U815 (N_815,N_7,N_47);
nand U816 (N_816,N_676,N_641);
xor U817 (N_817,N_497,N_407);
nor U818 (N_818,N_404,N_623);
xnor U819 (N_819,N_363,N_354);
xnor U820 (N_820,N_646,N_100);
xnor U821 (N_821,N_56,N_217);
nor U822 (N_822,N_747,N_26);
and U823 (N_823,N_512,N_239);
xnor U824 (N_824,N_390,N_720);
nand U825 (N_825,N_333,N_462);
or U826 (N_826,N_419,N_242);
xnor U827 (N_827,N_395,N_310);
nor U828 (N_828,N_548,N_314);
xnor U829 (N_829,N_214,N_605);
xnor U830 (N_830,N_147,N_322);
xor U831 (N_831,N_345,N_416);
and U832 (N_832,N_195,N_177);
or U833 (N_833,N_439,N_673);
xor U834 (N_834,N_320,N_90);
nand U835 (N_835,N_313,N_653);
xnor U836 (N_836,N_576,N_557);
and U837 (N_837,N_309,N_127);
and U838 (N_838,N_528,N_329);
nand U839 (N_839,N_734,N_318);
nand U840 (N_840,N_263,N_39);
xor U841 (N_841,N_536,N_74);
and U842 (N_842,N_336,N_150);
and U843 (N_843,N_443,N_703);
nand U844 (N_844,N_366,N_731);
xor U845 (N_845,N_81,N_379);
and U846 (N_846,N_485,N_181);
or U847 (N_847,N_292,N_325);
and U848 (N_848,N_80,N_139);
nor U849 (N_849,N_467,N_69);
and U850 (N_850,N_254,N_43);
nand U851 (N_851,N_461,N_434);
and U852 (N_852,N_257,N_533);
xnor U853 (N_853,N_737,N_378);
nor U854 (N_854,N_155,N_712);
nor U855 (N_855,N_661,N_640);
or U856 (N_856,N_573,N_597);
nor U857 (N_857,N_511,N_515);
xor U858 (N_858,N_169,N_581);
nand U859 (N_859,N_371,N_539);
and U860 (N_860,N_625,N_107);
and U861 (N_861,N_744,N_580);
and U862 (N_862,N_685,N_645);
xor U863 (N_863,N_109,N_460);
and U864 (N_864,N_124,N_128);
and U865 (N_865,N_716,N_383);
nand U866 (N_866,N_523,N_98);
xnor U867 (N_867,N_342,N_683);
xnor U868 (N_868,N_339,N_593);
nand U869 (N_869,N_130,N_264);
nand U870 (N_870,N_391,N_655);
or U871 (N_871,N_328,N_273);
and U872 (N_872,N_456,N_52);
nand U873 (N_873,N_149,N_225);
xnor U874 (N_874,N_621,N_525);
nand U875 (N_875,N_569,N_386);
xnor U876 (N_876,N_287,N_385);
or U877 (N_877,N_622,N_498);
xnor U878 (N_878,N_541,N_554);
or U879 (N_879,N_220,N_468);
and U880 (N_880,N_36,N_432);
or U881 (N_881,N_482,N_474);
xnor U882 (N_882,N_204,N_176);
xor U883 (N_883,N_261,N_701);
xnor U884 (N_884,N_630,N_237);
and U885 (N_885,N_367,N_278);
and U886 (N_886,N_563,N_722);
and U887 (N_887,N_571,N_189);
nor U888 (N_888,N_601,N_629);
nor U889 (N_889,N_674,N_732);
nor U890 (N_890,N_470,N_742);
nand U891 (N_891,N_230,N_301);
nand U892 (N_892,N_12,N_486);
nor U893 (N_893,N_114,N_564);
or U894 (N_894,N_276,N_10);
xnor U895 (N_895,N_421,N_294);
nor U896 (N_896,N_561,N_665);
and U897 (N_897,N_603,N_221);
xnor U898 (N_898,N_146,N_565);
nand U899 (N_899,N_494,N_450);
nor U900 (N_900,N_216,N_0);
nand U901 (N_901,N_353,N_83);
nor U902 (N_902,N_540,N_556);
and U903 (N_903,N_59,N_9);
xnor U904 (N_904,N_158,N_96);
or U905 (N_905,N_54,N_585);
nor U906 (N_906,N_704,N_412);
and U907 (N_907,N_17,N_526);
nand U908 (N_908,N_644,N_725);
nor U909 (N_909,N_429,N_469);
and U910 (N_910,N_77,N_186);
or U911 (N_911,N_637,N_184);
or U912 (N_912,N_664,N_696);
or U913 (N_913,N_241,N_509);
and U914 (N_914,N_516,N_153);
nand U915 (N_915,N_534,N_161);
nand U916 (N_916,N_527,N_389);
nand U917 (N_917,N_463,N_688);
nor U918 (N_918,N_250,N_666);
or U919 (N_919,N_546,N_327);
nor U920 (N_920,N_251,N_442);
and U921 (N_921,N_718,N_308);
nand U922 (N_922,N_143,N_185);
nand U923 (N_923,N_595,N_506);
and U924 (N_924,N_399,N_97);
xor U925 (N_925,N_178,N_446);
and U926 (N_926,N_544,N_420);
nand U927 (N_927,N_340,N_550);
or U928 (N_928,N_351,N_63);
nand U929 (N_929,N_402,N_364);
xnor U930 (N_930,N_710,N_436);
xnor U931 (N_931,N_156,N_634);
or U932 (N_932,N_218,N_431);
nand U933 (N_933,N_427,N_70);
nor U934 (N_934,N_532,N_607);
and U935 (N_935,N_142,N_682);
and U936 (N_936,N_587,N_739);
xnor U937 (N_937,N_566,N_35);
and U938 (N_938,N_562,N_610);
and U939 (N_939,N_302,N_691);
or U940 (N_940,N_542,N_95);
nand U941 (N_941,N_642,N_670);
xor U942 (N_942,N_370,N_105);
xnor U943 (N_943,N_211,N_93);
or U944 (N_944,N_192,N_244);
and U945 (N_945,N_531,N_708);
and U946 (N_946,N_72,N_730);
xor U947 (N_947,N_16,N_591);
xnor U948 (N_948,N_510,N_380);
and U949 (N_949,N_694,N_137);
nor U950 (N_950,N_598,N_193);
nand U951 (N_951,N_428,N_499);
or U952 (N_952,N_493,N_736);
nor U953 (N_953,N_501,N_616);
nor U954 (N_954,N_31,N_140);
or U955 (N_955,N_112,N_290);
or U956 (N_956,N_648,N_633);
or U957 (N_957,N_312,N_702);
or U958 (N_958,N_680,N_32);
nor U959 (N_959,N_13,N_457);
and U960 (N_960,N_48,N_592);
nor U961 (N_961,N_372,N_451);
or U962 (N_962,N_348,N_455);
xnor U963 (N_963,N_295,N_479);
or U964 (N_964,N_267,N_154);
nor U965 (N_965,N_152,N_58);
xnor U966 (N_966,N_619,N_259);
and U967 (N_967,N_330,N_663);
nand U968 (N_968,N_368,N_215);
xor U969 (N_969,N_1,N_504);
nand U970 (N_970,N_473,N_131);
xnor U971 (N_971,N_392,N_714);
or U972 (N_972,N_413,N_537);
and U973 (N_973,N_453,N_713);
nand U974 (N_974,N_198,N_409);
nand U975 (N_975,N_624,N_200);
and U976 (N_976,N_699,N_30);
xor U977 (N_977,N_384,N_549);
nor U978 (N_978,N_449,N_600);
and U979 (N_979,N_700,N_615);
xor U980 (N_980,N_291,N_268);
xnor U981 (N_981,N_102,N_163);
or U982 (N_982,N_628,N_84);
and U983 (N_983,N_21,N_425);
nand U984 (N_984,N_452,N_481);
xor U985 (N_985,N_282,N_272);
nand U986 (N_986,N_338,N_111);
nand U987 (N_987,N_639,N_162);
nand U988 (N_988,N_491,N_256);
or U989 (N_989,N_350,N_606);
xnor U990 (N_990,N_689,N_657);
xor U991 (N_991,N_671,N_698);
nor U992 (N_992,N_316,N_135);
nor U993 (N_993,N_166,N_41);
nor U994 (N_994,N_49,N_253);
or U995 (N_995,N_575,N_590);
and U996 (N_996,N_226,N_299);
nor U997 (N_997,N_589,N_334);
or U998 (N_998,N_660,N_435);
or U999 (N_999,N_471,N_315);
nor U1000 (N_1000,N_500,N_129);
nand U1001 (N_1001,N_182,N_324);
and U1002 (N_1002,N_197,N_620);
nand U1003 (N_1003,N_170,N_306);
and U1004 (N_1004,N_717,N_62);
nor U1005 (N_1005,N_119,N_480);
or U1006 (N_1006,N_24,N_144);
or U1007 (N_1007,N_520,N_496);
or U1008 (N_1008,N_711,N_535);
and U1009 (N_1009,N_281,N_103);
nor U1010 (N_1010,N_374,N_458);
nor U1011 (N_1011,N_745,N_654);
or U1012 (N_1012,N_159,N_579);
and U1013 (N_1013,N_631,N_355);
or U1014 (N_1014,N_265,N_201);
nor U1015 (N_1015,N_706,N_401);
nand U1016 (N_1016,N_614,N_558);
nor U1017 (N_1017,N_502,N_560);
nor U1018 (N_1018,N_229,N_567);
xor U1019 (N_1019,N_538,N_393);
xor U1020 (N_1020,N_332,N_466);
and U1021 (N_1021,N_406,N_596);
xor U1022 (N_1022,N_57,N_289);
nor U1023 (N_1023,N_475,N_132);
and U1024 (N_1024,N_360,N_247);
xor U1025 (N_1025,N_275,N_51);
nand U1026 (N_1026,N_110,N_437);
nor U1027 (N_1027,N_280,N_108);
nand U1028 (N_1028,N_555,N_599);
xor U1029 (N_1029,N_675,N_78);
and U1030 (N_1030,N_202,N_423);
or U1031 (N_1031,N_547,N_87);
or U1032 (N_1032,N_37,N_38);
nand U1033 (N_1033,N_341,N_672);
or U1034 (N_1034,N_695,N_438);
xnor U1035 (N_1035,N_213,N_662);
nand U1036 (N_1036,N_359,N_426);
nor U1037 (N_1037,N_743,N_444);
or U1038 (N_1038,N_219,N_183);
nand U1039 (N_1039,N_64,N_405);
or U1040 (N_1040,N_377,N_488);
xor U1041 (N_1041,N_246,N_483);
nor U1042 (N_1042,N_117,N_82);
or U1043 (N_1043,N_430,N_414);
nand U1044 (N_1044,N_415,N_319);
or U1045 (N_1045,N_2,N_298);
and U1046 (N_1046,N_724,N_553);
xor U1047 (N_1047,N_733,N_618);
and U1048 (N_1048,N_656,N_681);
and U1049 (N_1049,N_85,N_445);
xor U1050 (N_1050,N_530,N_643);
nand U1051 (N_1051,N_266,N_529);
xor U1052 (N_1052,N_326,N_588);
nand U1053 (N_1053,N_25,N_106);
or U1054 (N_1054,N_157,N_422);
or U1055 (N_1055,N_626,N_632);
xnor U1056 (N_1056,N_228,N_321);
or U1057 (N_1057,N_331,N_636);
xor U1058 (N_1058,N_116,N_586);
xnor U1059 (N_1059,N_151,N_88);
or U1060 (N_1060,N_126,N_735);
nand U1061 (N_1061,N_120,N_46);
nor U1062 (N_1062,N_53,N_617);
or U1063 (N_1063,N_15,N_238);
nand U1064 (N_1064,N_521,N_362);
nor U1065 (N_1065,N_270,N_190);
nand U1066 (N_1066,N_692,N_517);
xnor U1067 (N_1067,N_365,N_349);
or U1068 (N_1068,N_723,N_23);
or U1069 (N_1069,N_172,N_173);
or U1070 (N_1070,N_454,N_693);
or U1071 (N_1071,N_50,N_489);
or U1072 (N_1072,N_86,N_61);
nand U1073 (N_1073,N_658,N_196);
nor U1074 (N_1074,N_296,N_55);
and U1075 (N_1075,N_285,N_388);
or U1076 (N_1076,N_179,N_726);
and U1077 (N_1077,N_136,N_627);
xor U1078 (N_1078,N_258,N_233);
or U1079 (N_1079,N_222,N_28);
xor U1080 (N_1080,N_171,N_33);
nor U1081 (N_1081,N_403,N_719);
nor U1082 (N_1082,N_487,N_212);
and U1083 (N_1083,N_231,N_659);
nor U1084 (N_1084,N_284,N_223);
and U1085 (N_1085,N_175,N_60);
nand U1086 (N_1086,N_260,N_115);
xnor U1087 (N_1087,N_707,N_335);
nor U1088 (N_1088,N_194,N_652);
or U1089 (N_1089,N_76,N_65);
or U1090 (N_1090,N_343,N_373);
or U1091 (N_1091,N_684,N_188);
nor U1092 (N_1092,N_262,N_300);
and U1093 (N_1093,N_492,N_649);
or U1094 (N_1094,N_141,N_518);
nor U1095 (N_1095,N_27,N_667);
or U1096 (N_1096,N_208,N_277);
and U1097 (N_1097,N_29,N_252);
or U1098 (N_1098,N_650,N_669);
nand U1099 (N_1099,N_167,N_400);
or U1100 (N_1100,N_635,N_375);
nand U1101 (N_1101,N_240,N_210);
nor U1102 (N_1102,N_337,N_234);
or U1103 (N_1103,N_522,N_286);
or U1104 (N_1104,N_118,N_255);
nand U1105 (N_1105,N_199,N_715);
or U1106 (N_1106,N_249,N_459);
or U1107 (N_1107,N_66,N_138);
nand U1108 (N_1108,N_608,N_687);
or U1109 (N_1109,N_91,N_741);
nor U1110 (N_1110,N_99,N_133);
xnor U1111 (N_1111,N_738,N_604);
or U1112 (N_1112,N_18,N_638);
and U1113 (N_1113,N_410,N_283);
nand U1114 (N_1114,N_396,N_45);
xnor U1115 (N_1115,N_361,N_490);
nand U1116 (N_1116,N_6,N_746);
nand U1117 (N_1117,N_647,N_168);
and U1118 (N_1118,N_433,N_464);
nor U1119 (N_1119,N_20,N_476);
or U1120 (N_1120,N_358,N_397);
and U1121 (N_1121,N_668,N_243);
nand U1122 (N_1122,N_705,N_71);
xor U1123 (N_1123,N_594,N_552);
and U1124 (N_1124,N_75,N_347);
or U1125 (N_1125,N_196,N_461);
nor U1126 (N_1126,N_33,N_689);
nor U1127 (N_1127,N_383,N_428);
xor U1128 (N_1128,N_431,N_41);
and U1129 (N_1129,N_338,N_242);
nor U1130 (N_1130,N_269,N_607);
nor U1131 (N_1131,N_735,N_349);
and U1132 (N_1132,N_174,N_700);
xnor U1133 (N_1133,N_229,N_697);
or U1134 (N_1134,N_557,N_60);
xnor U1135 (N_1135,N_591,N_427);
xor U1136 (N_1136,N_592,N_248);
and U1137 (N_1137,N_364,N_75);
xnor U1138 (N_1138,N_695,N_341);
xnor U1139 (N_1139,N_142,N_394);
nor U1140 (N_1140,N_360,N_601);
or U1141 (N_1141,N_37,N_14);
xor U1142 (N_1142,N_149,N_49);
nor U1143 (N_1143,N_73,N_362);
nand U1144 (N_1144,N_211,N_510);
nand U1145 (N_1145,N_70,N_250);
nand U1146 (N_1146,N_559,N_257);
nor U1147 (N_1147,N_195,N_217);
nor U1148 (N_1148,N_634,N_668);
and U1149 (N_1149,N_78,N_326);
xor U1150 (N_1150,N_617,N_394);
xor U1151 (N_1151,N_627,N_340);
nor U1152 (N_1152,N_578,N_651);
nand U1153 (N_1153,N_678,N_349);
nor U1154 (N_1154,N_521,N_252);
nor U1155 (N_1155,N_327,N_300);
or U1156 (N_1156,N_743,N_572);
nor U1157 (N_1157,N_202,N_536);
xor U1158 (N_1158,N_506,N_304);
nor U1159 (N_1159,N_71,N_567);
or U1160 (N_1160,N_429,N_244);
nor U1161 (N_1161,N_736,N_421);
nand U1162 (N_1162,N_477,N_618);
nand U1163 (N_1163,N_239,N_256);
xnor U1164 (N_1164,N_648,N_367);
xnor U1165 (N_1165,N_108,N_734);
xnor U1166 (N_1166,N_54,N_175);
xnor U1167 (N_1167,N_426,N_61);
nor U1168 (N_1168,N_11,N_136);
xnor U1169 (N_1169,N_328,N_265);
nor U1170 (N_1170,N_273,N_512);
or U1171 (N_1171,N_444,N_620);
nor U1172 (N_1172,N_499,N_124);
nand U1173 (N_1173,N_295,N_434);
and U1174 (N_1174,N_178,N_211);
nand U1175 (N_1175,N_167,N_557);
and U1176 (N_1176,N_272,N_346);
or U1177 (N_1177,N_736,N_673);
and U1178 (N_1178,N_350,N_509);
or U1179 (N_1179,N_567,N_603);
nor U1180 (N_1180,N_365,N_570);
or U1181 (N_1181,N_731,N_368);
nand U1182 (N_1182,N_394,N_613);
xor U1183 (N_1183,N_467,N_710);
nand U1184 (N_1184,N_213,N_132);
and U1185 (N_1185,N_458,N_577);
or U1186 (N_1186,N_44,N_452);
nor U1187 (N_1187,N_532,N_241);
xor U1188 (N_1188,N_280,N_225);
nand U1189 (N_1189,N_603,N_258);
and U1190 (N_1190,N_740,N_662);
xor U1191 (N_1191,N_455,N_432);
xnor U1192 (N_1192,N_434,N_94);
nor U1193 (N_1193,N_270,N_389);
xnor U1194 (N_1194,N_471,N_116);
or U1195 (N_1195,N_722,N_465);
or U1196 (N_1196,N_417,N_557);
and U1197 (N_1197,N_99,N_422);
or U1198 (N_1198,N_669,N_95);
or U1199 (N_1199,N_251,N_426);
nand U1200 (N_1200,N_629,N_294);
and U1201 (N_1201,N_645,N_23);
or U1202 (N_1202,N_85,N_712);
nor U1203 (N_1203,N_725,N_170);
and U1204 (N_1204,N_709,N_566);
nor U1205 (N_1205,N_8,N_740);
nor U1206 (N_1206,N_576,N_192);
nand U1207 (N_1207,N_558,N_199);
or U1208 (N_1208,N_577,N_471);
and U1209 (N_1209,N_211,N_738);
nor U1210 (N_1210,N_441,N_470);
and U1211 (N_1211,N_343,N_495);
xnor U1212 (N_1212,N_629,N_87);
and U1213 (N_1213,N_255,N_682);
xor U1214 (N_1214,N_619,N_32);
and U1215 (N_1215,N_671,N_494);
xor U1216 (N_1216,N_200,N_27);
xnor U1217 (N_1217,N_533,N_511);
nor U1218 (N_1218,N_95,N_295);
xnor U1219 (N_1219,N_274,N_464);
xor U1220 (N_1220,N_660,N_140);
and U1221 (N_1221,N_13,N_102);
nand U1222 (N_1222,N_534,N_521);
or U1223 (N_1223,N_584,N_369);
xnor U1224 (N_1224,N_113,N_611);
and U1225 (N_1225,N_274,N_117);
nor U1226 (N_1226,N_648,N_327);
nand U1227 (N_1227,N_289,N_244);
xnor U1228 (N_1228,N_521,N_131);
nor U1229 (N_1229,N_324,N_416);
nand U1230 (N_1230,N_517,N_651);
xnor U1231 (N_1231,N_373,N_748);
or U1232 (N_1232,N_121,N_618);
and U1233 (N_1233,N_462,N_127);
nand U1234 (N_1234,N_60,N_85);
or U1235 (N_1235,N_167,N_330);
nor U1236 (N_1236,N_617,N_536);
or U1237 (N_1237,N_239,N_557);
nand U1238 (N_1238,N_442,N_172);
nand U1239 (N_1239,N_738,N_601);
or U1240 (N_1240,N_684,N_682);
nor U1241 (N_1241,N_167,N_60);
nor U1242 (N_1242,N_734,N_439);
xor U1243 (N_1243,N_345,N_152);
nor U1244 (N_1244,N_128,N_143);
nor U1245 (N_1245,N_328,N_16);
and U1246 (N_1246,N_416,N_613);
or U1247 (N_1247,N_263,N_557);
nor U1248 (N_1248,N_640,N_345);
nand U1249 (N_1249,N_14,N_483);
and U1250 (N_1250,N_597,N_161);
nor U1251 (N_1251,N_253,N_72);
and U1252 (N_1252,N_630,N_142);
or U1253 (N_1253,N_121,N_57);
xnor U1254 (N_1254,N_345,N_287);
or U1255 (N_1255,N_228,N_25);
nand U1256 (N_1256,N_666,N_127);
or U1257 (N_1257,N_281,N_404);
xor U1258 (N_1258,N_709,N_264);
or U1259 (N_1259,N_219,N_644);
nor U1260 (N_1260,N_300,N_310);
or U1261 (N_1261,N_357,N_343);
xnor U1262 (N_1262,N_376,N_577);
nor U1263 (N_1263,N_614,N_189);
and U1264 (N_1264,N_229,N_413);
nand U1265 (N_1265,N_546,N_383);
nor U1266 (N_1266,N_320,N_198);
and U1267 (N_1267,N_573,N_105);
or U1268 (N_1268,N_670,N_369);
nor U1269 (N_1269,N_225,N_99);
nand U1270 (N_1270,N_648,N_335);
xor U1271 (N_1271,N_599,N_258);
xnor U1272 (N_1272,N_624,N_126);
nand U1273 (N_1273,N_665,N_523);
and U1274 (N_1274,N_62,N_136);
nor U1275 (N_1275,N_144,N_434);
and U1276 (N_1276,N_597,N_156);
nor U1277 (N_1277,N_716,N_279);
or U1278 (N_1278,N_741,N_496);
xor U1279 (N_1279,N_468,N_253);
nor U1280 (N_1280,N_467,N_129);
xor U1281 (N_1281,N_299,N_305);
and U1282 (N_1282,N_610,N_497);
and U1283 (N_1283,N_314,N_732);
xor U1284 (N_1284,N_572,N_538);
and U1285 (N_1285,N_75,N_79);
nor U1286 (N_1286,N_6,N_308);
nor U1287 (N_1287,N_91,N_102);
and U1288 (N_1288,N_162,N_290);
or U1289 (N_1289,N_653,N_133);
xnor U1290 (N_1290,N_660,N_226);
or U1291 (N_1291,N_666,N_133);
nand U1292 (N_1292,N_132,N_402);
nor U1293 (N_1293,N_92,N_714);
nand U1294 (N_1294,N_252,N_170);
or U1295 (N_1295,N_738,N_482);
nand U1296 (N_1296,N_235,N_482);
and U1297 (N_1297,N_195,N_568);
and U1298 (N_1298,N_662,N_523);
nor U1299 (N_1299,N_317,N_226);
nand U1300 (N_1300,N_685,N_678);
or U1301 (N_1301,N_520,N_12);
nor U1302 (N_1302,N_440,N_153);
or U1303 (N_1303,N_86,N_395);
nand U1304 (N_1304,N_584,N_568);
and U1305 (N_1305,N_49,N_182);
and U1306 (N_1306,N_119,N_549);
and U1307 (N_1307,N_608,N_605);
xor U1308 (N_1308,N_504,N_69);
xnor U1309 (N_1309,N_470,N_317);
xor U1310 (N_1310,N_592,N_391);
xor U1311 (N_1311,N_368,N_720);
nor U1312 (N_1312,N_494,N_8);
xnor U1313 (N_1313,N_31,N_329);
nor U1314 (N_1314,N_43,N_706);
or U1315 (N_1315,N_175,N_652);
nor U1316 (N_1316,N_336,N_679);
nand U1317 (N_1317,N_310,N_482);
nand U1318 (N_1318,N_378,N_456);
xnor U1319 (N_1319,N_290,N_46);
and U1320 (N_1320,N_719,N_112);
nand U1321 (N_1321,N_368,N_116);
xnor U1322 (N_1322,N_37,N_388);
xnor U1323 (N_1323,N_602,N_94);
and U1324 (N_1324,N_534,N_399);
nand U1325 (N_1325,N_715,N_131);
or U1326 (N_1326,N_562,N_103);
or U1327 (N_1327,N_611,N_369);
or U1328 (N_1328,N_361,N_256);
and U1329 (N_1329,N_574,N_326);
nand U1330 (N_1330,N_371,N_382);
nor U1331 (N_1331,N_444,N_327);
nand U1332 (N_1332,N_190,N_105);
xnor U1333 (N_1333,N_569,N_495);
and U1334 (N_1334,N_393,N_295);
xor U1335 (N_1335,N_169,N_702);
xor U1336 (N_1336,N_462,N_201);
or U1337 (N_1337,N_38,N_508);
nor U1338 (N_1338,N_638,N_603);
nor U1339 (N_1339,N_115,N_111);
or U1340 (N_1340,N_328,N_613);
nor U1341 (N_1341,N_108,N_374);
or U1342 (N_1342,N_12,N_10);
nand U1343 (N_1343,N_648,N_135);
nor U1344 (N_1344,N_54,N_482);
nor U1345 (N_1345,N_501,N_59);
and U1346 (N_1346,N_69,N_554);
and U1347 (N_1347,N_141,N_569);
nand U1348 (N_1348,N_658,N_205);
nor U1349 (N_1349,N_744,N_468);
and U1350 (N_1350,N_645,N_732);
xnor U1351 (N_1351,N_613,N_400);
nand U1352 (N_1352,N_210,N_454);
or U1353 (N_1353,N_209,N_319);
nor U1354 (N_1354,N_162,N_620);
or U1355 (N_1355,N_680,N_327);
nor U1356 (N_1356,N_686,N_350);
and U1357 (N_1357,N_385,N_339);
and U1358 (N_1358,N_68,N_467);
or U1359 (N_1359,N_327,N_748);
nand U1360 (N_1360,N_484,N_644);
xnor U1361 (N_1361,N_746,N_421);
nand U1362 (N_1362,N_684,N_350);
xnor U1363 (N_1363,N_555,N_634);
xor U1364 (N_1364,N_37,N_325);
nor U1365 (N_1365,N_610,N_28);
nor U1366 (N_1366,N_26,N_10);
nor U1367 (N_1367,N_76,N_162);
nand U1368 (N_1368,N_576,N_473);
nor U1369 (N_1369,N_202,N_88);
or U1370 (N_1370,N_488,N_496);
or U1371 (N_1371,N_159,N_198);
and U1372 (N_1372,N_149,N_688);
nor U1373 (N_1373,N_130,N_400);
nor U1374 (N_1374,N_471,N_681);
nor U1375 (N_1375,N_654,N_143);
nand U1376 (N_1376,N_48,N_653);
xnor U1377 (N_1377,N_525,N_675);
nor U1378 (N_1378,N_703,N_420);
xor U1379 (N_1379,N_703,N_631);
nand U1380 (N_1380,N_527,N_485);
xnor U1381 (N_1381,N_653,N_177);
and U1382 (N_1382,N_217,N_184);
nor U1383 (N_1383,N_427,N_173);
nor U1384 (N_1384,N_255,N_157);
nand U1385 (N_1385,N_360,N_313);
and U1386 (N_1386,N_190,N_397);
xnor U1387 (N_1387,N_452,N_713);
nor U1388 (N_1388,N_465,N_47);
or U1389 (N_1389,N_577,N_80);
xnor U1390 (N_1390,N_713,N_302);
or U1391 (N_1391,N_37,N_159);
or U1392 (N_1392,N_326,N_6);
nand U1393 (N_1393,N_652,N_727);
nand U1394 (N_1394,N_646,N_560);
nor U1395 (N_1395,N_593,N_114);
xor U1396 (N_1396,N_506,N_300);
and U1397 (N_1397,N_637,N_54);
nand U1398 (N_1398,N_560,N_37);
or U1399 (N_1399,N_308,N_9);
or U1400 (N_1400,N_453,N_643);
or U1401 (N_1401,N_63,N_455);
xor U1402 (N_1402,N_372,N_29);
or U1403 (N_1403,N_736,N_663);
xnor U1404 (N_1404,N_675,N_272);
xor U1405 (N_1405,N_276,N_200);
xor U1406 (N_1406,N_218,N_466);
nand U1407 (N_1407,N_256,N_652);
nor U1408 (N_1408,N_498,N_343);
or U1409 (N_1409,N_747,N_464);
nor U1410 (N_1410,N_246,N_148);
nand U1411 (N_1411,N_688,N_74);
nand U1412 (N_1412,N_23,N_407);
and U1413 (N_1413,N_2,N_482);
and U1414 (N_1414,N_688,N_298);
and U1415 (N_1415,N_174,N_169);
nor U1416 (N_1416,N_310,N_737);
xor U1417 (N_1417,N_620,N_297);
xor U1418 (N_1418,N_162,N_415);
and U1419 (N_1419,N_629,N_95);
xnor U1420 (N_1420,N_581,N_438);
xor U1421 (N_1421,N_578,N_105);
nor U1422 (N_1422,N_179,N_311);
or U1423 (N_1423,N_91,N_748);
nor U1424 (N_1424,N_484,N_204);
xnor U1425 (N_1425,N_276,N_512);
nand U1426 (N_1426,N_743,N_73);
nand U1427 (N_1427,N_662,N_60);
nor U1428 (N_1428,N_40,N_441);
nand U1429 (N_1429,N_641,N_661);
nor U1430 (N_1430,N_736,N_143);
or U1431 (N_1431,N_739,N_428);
xor U1432 (N_1432,N_551,N_565);
nor U1433 (N_1433,N_335,N_305);
and U1434 (N_1434,N_445,N_395);
or U1435 (N_1435,N_119,N_72);
nand U1436 (N_1436,N_95,N_505);
nor U1437 (N_1437,N_401,N_348);
or U1438 (N_1438,N_363,N_275);
xor U1439 (N_1439,N_622,N_403);
and U1440 (N_1440,N_437,N_417);
and U1441 (N_1441,N_217,N_624);
xnor U1442 (N_1442,N_654,N_656);
or U1443 (N_1443,N_519,N_31);
nor U1444 (N_1444,N_455,N_163);
nor U1445 (N_1445,N_179,N_745);
and U1446 (N_1446,N_146,N_140);
nor U1447 (N_1447,N_335,N_98);
and U1448 (N_1448,N_129,N_517);
and U1449 (N_1449,N_89,N_506);
nor U1450 (N_1450,N_411,N_457);
or U1451 (N_1451,N_40,N_65);
xor U1452 (N_1452,N_470,N_725);
nand U1453 (N_1453,N_351,N_100);
nor U1454 (N_1454,N_7,N_744);
or U1455 (N_1455,N_610,N_147);
xor U1456 (N_1456,N_319,N_336);
nor U1457 (N_1457,N_146,N_382);
nor U1458 (N_1458,N_712,N_277);
xor U1459 (N_1459,N_534,N_52);
and U1460 (N_1460,N_214,N_446);
or U1461 (N_1461,N_370,N_688);
xnor U1462 (N_1462,N_253,N_88);
xor U1463 (N_1463,N_246,N_41);
nand U1464 (N_1464,N_541,N_349);
nor U1465 (N_1465,N_451,N_443);
nand U1466 (N_1466,N_469,N_468);
nand U1467 (N_1467,N_74,N_698);
and U1468 (N_1468,N_74,N_178);
nand U1469 (N_1469,N_510,N_188);
xor U1470 (N_1470,N_537,N_72);
nor U1471 (N_1471,N_265,N_695);
and U1472 (N_1472,N_106,N_239);
nor U1473 (N_1473,N_294,N_498);
nand U1474 (N_1474,N_561,N_483);
xnor U1475 (N_1475,N_705,N_252);
or U1476 (N_1476,N_201,N_340);
and U1477 (N_1477,N_249,N_223);
or U1478 (N_1478,N_33,N_511);
and U1479 (N_1479,N_645,N_253);
and U1480 (N_1480,N_263,N_679);
nor U1481 (N_1481,N_284,N_26);
and U1482 (N_1482,N_674,N_509);
and U1483 (N_1483,N_429,N_494);
nor U1484 (N_1484,N_551,N_427);
and U1485 (N_1485,N_440,N_131);
and U1486 (N_1486,N_30,N_138);
or U1487 (N_1487,N_131,N_663);
nand U1488 (N_1488,N_653,N_483);
xor U1489 (N_1489,N_27,N_461);
nand U1490 (N_1490,N_401,N_731);
or U1491 (N_1491,N_103,N_193);
xnor U1492 (N_1492,N_411,N_571);
xor U1493 (N_1493,N_3,N_184);
and U1494 (N_1494,N_682,N_220);
and U1495 (N_1495,N_698,N_433);
nand U1496 (N_1496,N_550,N_691);
xnor U1497 (N_1497,N_410,N_45);
or U1498 (N_1498,N_538,N_559);
xnor U1499 (N_1499,N_78,N_194);
xnor U1500 (N_1500,N_1057,N_1413);
and U1501 (N_1501,N_855,N_866);
nand U1502 (N_1502,N_1375,N_1472);
or U1503 (N_1503,N_1348,N_1447);
and U1504 (N_1504,N_905,N_1175);
or U1505 (N_1505,N_1405,N_812);
nand U1506 (N_1506,N_1191,N_1371);
nor U1507 (N_1507,N_1242,N_1250);
nand U1508 (N_1508,N_1215,N_1489);
or U1509 (N_1509,N_822,N_1309);
and U1510 (N_1510,N_1243,N_1248);
nand U1511 (N_1511,N_1380,N_987);
nor U1512 (N_1512,N_1293,N_1184);
nand U1513 (N_1513,N_1171,N_1263);
or U1514 (N_1514,N_1276,N_862);
and U1515 (N_1515,N_1000,N_1435);
nand U1516 (N_1516,N_1361,N_770);
and U1517 (N_1517,N_1335,N_1238);
and U1518 (N_1518,N_1189,N_1245);
xor U1519 (N_1519,N_841,N_1100);
and U1520 (N_1520,N_1305,N_773);
nor U1521 (N_1521,N_858,N_985);
nand U1522 (N_1522,N_1469,N_1442);
or U1523 (N_1523,N_1239,N_818);
nor U1524 (N_1524,N_1164,N_942);
xor U1525 (N_1525,N_1384,N_1343);
nor U1526 (N_1526,N_1203,N_1251);
or U1527 (N_1527,N_1271,N_1226);
or U1528 (N_1528,N_922,N_1446);
and U1529 (N_1529,N_783,N_850);
or U1530 (N_1530,N_1381,N_786);
xor U1531 (N_1531,N_823,N_1112);
and U1532 (N_1532,N_1399,N_1428);
nor U1533 (N_1533,N_1369,N_1159);
nand U1534 (N_1534,N_1105,N_1430);
nand U1535 (N_1535,N_1227,N_1037);
nand U1536 (N_1536,N_1198,N_1476);
xor U1537 (N_1537,N_1456,N_986);
and U1538 (N_1538,N_901,N_1039);
nor U1539 (N_1539,N_1196,N_1424);
or U1540 (N_1540,N_873,N_930);
and U1541 (N_1541,N_1033,N_996);
xor U1542 (N_1542,N_1177,N_1449);
xor U1543 (N_1543,N_1154,N_1475);
and U1544 (N_1544,N_1054,N_1099);
nor U1545 (N_1545,N_1032,N_1160);
xnor U1546 (N_1546,N_1264,N_1342);
nor U1547 (N_1547,N_766,N_1417);
or U1548 (N_1548,N_1454,N_1019);
nor U1549 (N_1549,N_1185,N_1444);
nand U1550 (N_1550,N_848,N_1117);
or U1551 (N_1551,N_1025,N_1055);
and U1552 (N_1552,N_924,N_1073);
or U1553 (N_1553,N_958,N_1300);
or U1554 (N_1554,N_1115,N_1045);
and U1555 (N_1555,N_1436,N_1034);
nand U1556 (N_1556,N_1443,N_1323);
or U1557 (N_1557,N_1230,N_1273);
or U1558 (N_1558,N_1471,N_1272);
nor U1559 (N_1559,N_1079,N_871);
nor U1560 (N_1560,N_1004,N_1278);
and U1561 (N_1561,N_897,N_1458);
nand U1562 (N_1562,N_831,N_751);
nand U1563 (N_1563,N_923,N_874);
nor U1564 (N_1564,N_767,N_1247);
xnor U1565 (N_1565,N_1216,N_938);
and U1566 (N_1566,N_1410,N_1485);
xor U1567 (N_1567,N_1061,N_808);
xnor U1568 (N_1568,N_1134,N_1155);
or U1569 (N_1569,N_1144,N_1122);
and U1570 (N_1570,N_1492,N_828);
or U1571 (N_1571,N_1167,N_1332);
nand U1572 (N_1572,N_950,N_1150);
or U1573 (N_1573,N_1451,N_877);
nor U1574 (N_1574,N_991,N_1081);
xor U1575 (N_1575,N_1253,N_1224);
nor U1576 (N_1576,N_1408,N_943);
or U1577 (N_1577,N_1268,N_1313);
nand U1578 (N_1578,N_1360,N_1455);
xnor U1579 (N_1579,N_830,N_1161);
xor U1580 (N_1580,N_929,N_1119);
or U1581 (N_1581,N_976,N_1098);
nor U1582 (N_1582,N_1209,N_1064);
nand U1583 (N_1583,N_953,N_968);
nand U1584 (N_1584,N_1016,N_1307);
xnor U1585 (N_1585,N_1212,N_913);
nand U1586 (N_1586,N_1074,N_1445);
nor U1587 (N_1587,N_1474,N_1072);
nand U1588 (N_1588,N_944,N_1101);
nand U1589 (N_1589,N_945,N_1292);
xnor U1590 (N_1590,N_979,N_967);
or U1591 (N_1591,N_1056,N_834);
nand U1592 (N_1592,N_1063,N_1046);
nor U1593 (N_1593,N_1133,N_1314);
and U1594 (N_1594,N_1481,N_1421);
nor U1595 (N_1595,N_1350,N_1179);
nand U1596 (N_1596,N_1165,N_964);
or U1597 (N_1597,N_925,N_1131);
nand U1598 (N_1598,N_1206,N_965);
xor U1599 (N_1599,N_1174,N_1409);
and U1600 (N_1600,N_875,N_1254);
or U1601 (N_1601,N_1108,N_1194);
nand U1602 (N_1602,N_1013,N_960);
and U1603 (N_1603,N_817,N_1319);
nand U1604 (N_1604,N_1383,N_1301);
nor U1605 (N_1605,N_956,N_1386);
nand U1606 (N_1606,N_1240,N_1279);
or U1607 (N_1607,N_1130,N_792);
and U1608 (N_1608,N_1494,N_813);
nor U1609 (N_1609,N_1364,N_1008);
and U1610 (N_1610,N_762,N_961);
nor U1611 (N_1611,N_1420,N_889);
xor U1612 (N_1612,N_1357,N_1393);
nand U1613 (N_1613,N_833,N_849);
nor U1614 (N_1614,N_1087,N_883);
xor U1615 (N_1615,N_843,N_1295);
nand U1616 (N_1616,N_752,N_1459);
or U1617 (N_1617,N_769,N_832);
nand U1618 (N_1618,N_993,N_1345);
or U1619 (N_1619,N_963,N_1488);
and U1620 (N_1620,N_1389,N_1135);
xnor U1621 (N_1621,N_1036,N_1014);
and U1622 (N_1622,N_1022,N_1329);
xnor U1623 (N_1623,N_1235,N_840);
nor U1624 (N_1624,N_1395,N_1390);
and U1625 (N_1625,N_1152,N_1321);
xnor U1626 (N_1626,N_1249,N_1180);
or U1627 (N_1627,N_915,N_1480);
or U1628 (N_1628,N_797,N_1285);
or U1629 (N_1629,N_937,N_1170);
or U1630 (N_1630,N_1225,N_1116);
nand U1631 (N_1631,N_1317,N_1414);
nand U1632 (N_1632,N_1286,N_1487);
nand U1633 (N_1633,N_894,N_1477);
xor U1634 (N_1634,N_1190,N_1288);
and U1635 (N_1635,N_750,N_983);
nand U1636 (N_1636,N_1402,N_1188);
nand U1637 (N_1637,N_779,N_1450);
xnor U1638 (N_1638,N_997,N_1388);
nor U1639 (N_1639,N_860,N_815);
or U1640 (N_1640,N_1151,N_857);
nand U1641 (N_1641,N_878,N_899);
nor U1642 (N_1642,N_887,N_1229);
or U1643 (N_1643,N_911,N_1473);
nand U1644 (N_1644,N_1166,N_959);
and U1645 (N_1645,N_816,N_934);
nand U1646 (N_1646,N_1440,N_1035);
xor U1647 (N_1647,N_1128,N_1283);
and U1648 (N_1648,N_1241,N_876);
nand U1649 (N_1649,N_1124,N_1193);
and U1650 (N_1650,N_785,N_1096);
nor U1651 (N_1651,N_1065,N_916);
nor U1652 (N_1652,N_1137,N_829);
and U1653 (N_1653,N_1041,N_1269);
nand U1654 (N_1654,N_1322,N_1419);
nand U1655 (N_1655,N_806,N_1136);
and U1656 (N_1656,N_1094,N_1259);
nor U1657 (N_1657,N_1303,N_879);
xnor U1658 (N_1658,N_1059,N_775);
xor U1659 (N_1659,N_814,N_1341);
nand U1660 (N_1660,N_1316,N_1090);
nand U1661 (N_1661,N_1298,N_776);
xor U1662 (N_1662,N_870,N_1483);
nand U1663 (N_1663,N_1182,N_1205);
nor U1664 (N_1664,N_1132,N_1318);
or U1665 (N_1665,N_978,N_892);
nor U1666 (N_1666,N_1261,N_1222);
and U1667 (N_1667,N_1213,N_1416);
xor U1668 (N_1668,N_1289,N_970);
or U1669 (N_1669,N_1429,N_1018);
nand U1670 (N_1670,N_1311,N_1398);
xor U1671 (N_1671,N_795,N_758);
and U1672 (N_1672,N_1491,N_1060);
xnor U1673 (N_1673,N_1049,N_1040);
nor U1674 (N_1674,N_1392,N_914);
nor U1675 (N_1675,N_1376,N_1200);
nor U1676 (N_1676,N_819,N_1156);
xnor U1677 (N_1677,N_1221,N_1172);
or U1678 (N_1678,N_1084,N_1365);
or U1679 (N_1679,N_984,N_1207);
nor U1680 (N_1680,N_1490,N_1328);
xor U1681 (N_1681,N_888,N_1223);
xnor U1682 (N_1682,N_824,N_895);
xor U1683 (N_1683,N_1220,N_1062);
and U1684 (N_1684,N_1274,N_1373);
or U1685 (N_1685,N_992,N_952);
nand U1686 (N_1686,N_1479,N_847);
nand U1687 (N_1687,N_1423,N_759);
nor U1688 (N_1688,N_898,N_1187);
or U1689 (N_1689,N_1176,N_1030);
xor U1690 (N_1690,N_761,N_1181);
nand U1691 (N_1691,N_1277,N_1403);
or U1692 (N_1692,N_1326,N_900);
or U1693 (N_1693,N_1106,N_908);
xnor U1694 (N_1694,N_1366,N_753);
xnor U1695 (N_1695,N_1299,N_1431);
nand U1696 (N_1696,N_1109,N_1005);
and U1697 (N_1697,N_1140,N_846);
nor U1698 (N_1698,N_1453,N_890);
or U1699 (N_1699,N_1282,N_1486);
or U1700 (N_1700,N_1201,N_1434);
nand U1701 (N_1701,N_1262,N_1021);
and U1702 (N_1702,N_1338,N_801);
xor U1703 (N_1703,N_755,N_1493);
xor U1704 (N_1704,N_864,N_1382);
nand U1705 (N_1705,N_1192,N_1400);
and U1706 (N_1706,N_868,N_1051);
xor U1707 (N_1707,N_826,N_1157);
or U1708 (N_1708,N_856,N_1337);
nand U1709 (N_1709,N_1378,N_1080);
and U1710 (N_1710,N_1359,N_804);
nor U1711 (N_1711,N_1024,N_951);
nand U1712 (N_1712,N_1147,N_1267);
xor U1713 (N_1713,N_1071,N_1053);
nor U1714 (N_1714,N_1448,N_1415);
nand U1715 (N_1715,N_1139,N_771);
and U1716 (N_1716,N_949,N_981);
xor U1717 (N_1717,N_1391,N_884);
xnor U1718 (N_1718,N_1102,N_1197);
or U1719 (N_1719,N_948,N_1125);
and U1720 (N_1720,N_798,N_893);
nor U1721 (N_1721,N_763,N_1009);
and U1722 (N_1722,N_861,N_1347);
xnor U1723 (N_1723,N_1266,N_1284);
nand U1724 (N_1724,N_772,N_1237);
nor U1725 (N_1725,N_1233,N_1302);
and U1726 (N_1726,N_1070,N_1126);
or U1727 (N_1727,N_907,N_971);
nor U1728 (N_1728,N_1252,N_863);
xnor U1729 (N_1729,N_1367,N_1394);
nand U1730 (N_1730,N_844,N_1387);
or U1731 (N_1731,N_955,N_1002);
xor U1732 (N_1732,N_975,N_757);
nor U1733 (N_1733,N_1129,N_1256);
nor U1734 (N_1734,N_1017,N_1228);
nor U1735 (N_1735,N_935,N_1412);
xor U1736 (N_1736,N_1330,N_789);
nor U1737 (N_1737,N_1068,N_1260);
nand U1738 (N_1738,N_1495,N_1110);
nor U1739 (N_1739,N_1346,N_768);
nor U1740 (N_1740,N_1461,N_1003);
xor U1741 (N_1741,N_1370,N_778);
xor U1742 (N_1742,N_1173,N_932);
nand U1743 (N_1743,N_1291,N_793);
nor U1744 (N_1744,N_1236,N_1287);
and U1745 (N_1745,N_854,N_1437);
or U1746 (N_1746,N_1464,N_1385);
xor U1747 (N_1747,N_836,N_919);
or U1748 (N_1748,N_1031,N_946);
nand U1749 (N_1749,N_1093,N_982);
nor U1750 (N_1750,N_1324,N_1149);
nand U1751 (N_1751,N_1496,N_1012);
and U1752 (N_1752,N_1028,N_1499);
and U1753 (N_1753,N_774,N_859);
nand U1754 (N_1754,N_784,N_1452);
or U1755 (N_1755,N_1426,N_1107);
and U1756 (N_1756,N_1463,N_1076);
or U1757 (N_1757,N_802,N_1083);
nand U1758 (N_1758,N_1441,N_1211);
or U1759 (N_1759,N_1497,N_1265);
nor U1760 (N_1760,N_809,N_962);
or U1761 (N_1761,N_1086,N_1075);
nand U1762 (N_1762,N_882,N_782);
nand U1763 (N_1763,N_853,N_931);
nor U1764 (N_1764,N_1010,N_1162);
xnor U1765 (N_1765,N_906,N_839);
xnor U1766 (N_1766,N_1304,N_1433);
xnor U1767 (N_1767,N_1484,N_842);
nand U1768 (N_1768,N_1275,N_1320);
nand U1769 (N_1769,N_995,N_1043);
and U1770 (N_1770,N_794,N_1315);
nand U1771 (N_1771,N_1186,N_1308);
or U1772 (N_1772,N_1042,N_936);
xor U1773 (N_1773,N_998,N_1118);
and U1774 (N_1774,N_1310,N_1358);
or U1775 (N_1775,N_1354,N_1097);
nor U1776 (N_1776,N_1396,N_1246);
or U1777 (N_1777,N_1406,N_954);
xnor U1778 (N_1778,N_1336,N_1457);
or U1779 (N_1779,N_803,N_760);
xnor U1780 (N_1780,N_1427,N_1082);
xnor U1781 (N_1781,N_1141,N_1026);
nor U1782 (N_1782,N_1178,N_1123);
or U1783 (N_1783,N_1334,N_1407);
or U1784 (N_1784,N_1029,N_1217);
nand U1785 (N_1785,N_1163,N_902);
or U1786 (N_1786,N_957,N_1044);
nand U1787 (N_1787,N_1023,N_1498);
or U1788 (N_1788,N_990,N_1127);
and U1789 (N_1789,N_810,N_781);
nor U1790 (N_1790,N_1258,N_1052);
nand U1791 (N_1791,N_1377,N_1462);
xnor U1792 (N_1792,N_921,N_1296);
or U1793 (N_1793,N_845,N_791);
xor U1794 (N_1794,N_787,N_1356);
nor U1795 (N_1795,N_1006,N_764);
and U1796 (N_1796,N_827,N_1183);
nand U1797 (N_1797,N_1363,N_1210);
and U1798 (N_1798,N_928,N_800);
xnor U1799 (N_1799,N_1111,N_1244);
nand U1800 (N_1800,N_969,N_989);
xor U1801 (N_1801,N_1050,N_1425);
or U1802 (N_1802,N_1143,N_1048);
or U1803 (N_1803,N_807,N_1104);
xnor U1804 (N_1804,N_1482,N_1372);
nand U1805 (N_1805,N_1066,N_1114);
nand U1806 (N_1806,N_1418,N_973);
nor U1807 (N_1807,N_1219,N_999);
or U1808 (N_1808,N_1011,N_1439);
nand U1809 (N_1809,N_1208,N_903);
nand U1810 (N_1810,N_1362,N_1047);
nand U1811 (N_1811,N_1411,N_851);
nor U1812 (N_1812,N_1020,N_1379);
xnor U1813 (N_1813,N_1460,N_1333);
nand U1814 (N_1814,N_788,N_927);
nand U1815 (N_1815,N_918,N_1325);
or U1816 (N_1816,N_1120,N_1113);
nand U1817 (N_1817,N_780,N_939);
or U1818 (N_1818,N_891,N_1397);
nand U1819 (N_1819,N_1467,N_972);
nor U1820 (N_1820,N_1015,N_1281);
nand U1821 (N_1821,N_1312,N_1327);
or U1822 (N_1822,N_1199,N_777);
nor U1823 (N_1823,N_1195,N_1438);
or U1824 (N_1824,N_1145,N_920);
nand U1825 (N_1825,N_1255,N_756);
and U1826 (N_1826,N_1085,N_1422);
nand U1827 (N_1827,N_974,N_1148);
and U1828 (N_1828,N_926,N_1306);
xnor U1829 (N_1829,N_933,N_1294);
and U1830 (N_1830,N_1058,N_941);
or U1831 (N_1831,N_796,N_904);
nor U1832 (N_1832,N_865,N_988);
nor U1833 (N_1833,N_1218,N_977);
and U1834 (N_1834,N_1103,N_917);
or U1835 (N_1835,N_980,N_881);
or U1836 (N_1836,N_1432,N_838);
or U1837 (N_1837,N_1091,N_1466);
nand U1838 (N_1838,N_1121,N_1404);
xor U1839 (N_1839,N_1297,N_1089);
xnor U1840 (N_1840,N_1355,N_820);
xor U1841 (N_1841,N_1478,N_1067);
and U1842 (N_1842,N_790,N_754);
nand U1843 (N_1843,N_1078,N_1232);
nand U1844 (N_1844,N_994,N_910);
and U1845 (N_1845,N_765,N_1401);
nor U1846 (N_1846,N_1465,N_1468);
nand U1847 (N_1847,N_1027,N_940);
nor U1848 (N_1848,N_835,N_825);
and U1849 (N_1849,N_1038,N_1290);
nand U1850 (N_1850,N_1280,N_896);
nand U1851 (N_1851,N_869,N_1158);
or U1852 (N_1852,N_805,N_799);
or U1853 (N_1853,N_837,N_1257);
nor U1854 (N_1854,N_811,N_1368);
xnor U1855 (N_1855,N_1234,N_909);
nand U1856 (N_1856,N_1088,N_912);
nor U1857 (N_1857,N_1153,N_947);
xor U1858 (N_1858,N_885,N_1231);
nor U1859 (N_1859,N_867,N_1270);
and U1860 (N_1860,N_1092,N_1001);
or U1861 (N_1861,N_1344,N_1069);
xnor U1862 (N_1862,N_1142,N_1138);
nor U1863 (N_1863,N_966,N_1340);
xor U1864 (N_1864,N_1353,N_872);
and U1865 (N_1865,N_1331,N_821);
or U1866 (N_1866,N_1339,N_1204);
xor U1867 (N_1867,N_1146,N_1351);
nand U1868 (N_1868,N_886,N_1349);
nor U1869 (N_1869,N_1007,N_1352);
and U1870 (N_1870,N_1374,N_880);
and U1871 (N_1871,N_852,N_1169);
nand U1872 (N_1872,N_1214,N_1077);
or U1873 (N_1873,N_1470,N_1168);
xor U1874 (N_1874,N_1202,N_1095);
or U1875 (N_1875,N_750,N_1279);
and U1876 (N_1876,N_942,N_1460);
nand U1877 (N_1877,N_891,N_1207);
and U1878 (N_1878,N_1347,N_1406);
and U1879 (N_1879,N_1443,N_857);
xor U1880 (N_1880,N_1185,N_1448);
or U1881 (N_1881,N_953,N_1000);
and U1882 (N_1882,N_1011,N_1106);
xnor U1883 (N_1883,N_1273,N_1015);
and U1884 (N_1884,N_1331,N_1029);
nand U1885 (N_1885,N_1080,N_1162);
or U1886 (N_1886,N_1096,N_1351);
xor U1887 (N_1887,N_996,N_830);
nor U1888 (N_1888,N_1179,N_1112);
xnor U1889 (N_1889,N_1252,N_1320);
and U1890 (N_1890,N_1395,N_1103);
nor U1891 (N_1891,N_819,N_1244);
nand U1892 (N_1892,N_1058,N_1444);
and U1893 (N_1893,N_1245,N_1062);
and U1894 (N_1894,N_1435,N_847);
xor U1895 (N_1895,N_1163,N_925);
xor U1896 (N_1896,N_1132,N_1224);
xnor U1897 (N_1897,N_903,N_864);
nor U1898 (N_1898,N_1150,N_1484);
or U1899 (N_1899,N_1449,N_1239);
nor U1900 (N_1900,N_948,N_763);
nor U1901 (N_1901,N_1486,N_1304);
nand U1902 (N_1902,N_1035,N_1413);
and U1903 (N_1903,N_993,N_1373);
xnor U1904 (N_1904,N_1155,N_784);
nor U1905 (N_1905,N_1394,N_1334);
xor U1906 (N_1906,N_1217,N_878);
nand U1907 (N_1907,N_1250,N_952);
xnor U1908 (N_1908,N_874,N_1340);
nor U1909 (N_1909,N_975,N_1121);
nand U1910 (N_1910,N_848,N_1268);
nor U1911 (N_1911,N_1246,N_1042);
nor U1912 (N_1912,N_1247,N_1406);
and U1913 (N_1913,N_1203,N_1239);
xor U1914 (N_1914,N_794,N_1432);
xnor U1915 (N_1915,N_806,N_844);
or U1916 (N_1916,N_901,N_1192);
xor U1917 (N_1917,N_1439,N_1302);
nor U1918 (N_1918,N_869,N_1409);
or U1919 (N_1919,N_1333,N_1187);
nor U1920 (N_1920,N_1165,N_1496);
and U1921 (N_1921,N_1072,N_1379);
or U1922 (N_1922,N_1114,N_910);
xnor U1923 (N_1923,N_866,N_1274);
nor U1924 (N_1924,N_918,N_1048);
or U1925 (N_1925,N_864,N_1141);
or U1926 (N_1926,N_965,N_1076);
nand U1927 (N_1927,N_1108,N_1150);
nor U1928 (N_1928,N_1087,N_1323);
xnor U1929 (N_1929,N_950,N_1215);
nand U1930 (N_1930,N_1008,N_1265);
xnor U1931 (N_1931,N_777,N_880);
xor U1932 (N_1932,N_867,N_1277);
xnor U1933 (N_1933,N_1251,N_1417);
or U1934 (N_1934,N_1309,N_1390);
or U1935 (N_1935,N_1347,N_1166);
or U1936 (N_1936,N_1248,N_1082);
nand U1937 (N_1937,N_912,N_857);
and U1938 (N_1938,N_855,N_1268);
and U1939 (N_1939,N_1379,N_1196);
and U1940 (N_1940,N_1164,N_808);
or U1941 (N_1941,N_878,N_1064);
and U1942 (N_1942,N_1448,N_1005);
nor U1943 (N_1943,N_816,N_1208);
or U1944 (N_1944,N_858,N_1361);
nand U1945 (N_1945,N_945,N_1256);
xnor U1946 (N_1946,N_1378,N_785);
or U1947 (N_1947,N_1305,N_1115);
or U1948 (N_1948,N_1337,N_813);
xnor U1949 (N_1949,N_1290,N_913);
nor U1950 (N_1950,N_799,N_1007);
xor U1951 (N_1951,N_762,N_1174);
xnor U1952 (N_1952,N_1160,N_970);
and U1953 (N_1953,N_1482,N_1304);
or U1954 (N_1954,N_1057,N_1213);
nand U1955 (N_1955,N_1405,N_1390);
or U1956 (N_1956,N_1050,N_886);
or U1957 (N_1957,N_1187,N_1305);
and U1958 (N_1958,N_1033,N_1414);
nand U1959 (N_1959,N_1115,N_1133);
and U1960 (N_1960,N_1184,N_990);
and U1961 (N_1961,N_1489,N_1081);
xnor U1962 (N_1962,N_1198,N_793);
and U1963 (N_1963,N_1034,N_1014);
nand U1964 (N_1964,N_1047,N_1265);
and U1965 (N_1965,N_770,N_843);
or U1966 (N_1966,N_1218,N_1006);
or U1967 (N_1967,N_1313,N_825);
xnor U1968 (N_1968,N_784,N_1154);
and U1969 (N_1969,N_1237,N_867);
or U1970 (N_1970,N_850,N_1454);
and U1971 (N_1971,N_989,N_1282);
and U1972 (N_1972,N_1492,N_1288);
and U1973 (N_1973,N_806,N_950);
nor U1974 (N_1974,N_1434,N_1388);
nand U1975 (N_1975,N_882,N_1079);
xnor U1976 (N_1976,N_921,N_765);
and U1977 (N_1977,N_1094,N_774);
nand U1978 (N_1978,N_1365,N_1080);
or U1979 (N_1979,N_1404,N_1166);
and U1980 (N_1980,N_1397,N_811);
xnor U1981 (N_1981,N_1366,N_1320);
nor U1982 (N_1982,N_1318,N_1344);
nand U1983 (N_1983,N_798,N_1417);
or U1984 (N_1984,N_859,N_950);
xnor U1985 (N_1985,N_912,N_1256);
nand U1986 (N_1986,N_1460,N_1424);
and U1987 (N_1987,N_1181,N_973);
nand U1988 (N_1988,N_792,N_1033);
xnor U1989 (N_1989,N_1394,N_1391);
nand U1990 (N_1990,N_1174,N_813);
nand U1991 (N_1991,N_1009,N_1056);
or U1992 (N_1992,N_1412,N_918);
xnor U1993 (N_1993,N_1024,N_1066);
and U1994 (N_1994,N_831,N_1128);
nand U1995 (N_1995,N_792,N_966);
nand U1996 (N_1996,N_1336,N_1029);
nand U1997 (N_1997,N_1230,N_1222);
nor U1998 (N_1998,N_1205,N_755);
nor U1999 (N_1999,N_1461,N_776);
nand U2000 (N_2000,N_1354,N_1400);
nand U2001 (N_2001,N_796,N_1480);
and U2002 (N_2002,N_784,N_774);
nand U2003 (N_2003,N_1107,N_1009);
xor U2004 (N_2004,N_879,N_1267);
nor U2005 (N_2005,N_914,N_1343);
xor U2006 (N_2006,N_752,N_1460);
nor U2007 (N_2007,N_928,N_821);
nand U2008 (N_2008,N_929,N_786);
and U2009 (N_2009,N_934,N_1023);
nor U2010 (N_2010,N_980,N_1291);
xnor U2011 (N_2011,N_1476,N_1352);
nand U2012 (N_2012,N_859,N_981);
or U2013 (N_2013,N_1478,N_871);
and U2014 (N_2014,N_868,N_1106);
xnor U2015 (N_2015,N_1070,N_1178);
xor U2016 (N_2016,N_1273,N_1223);
nor U2017 (N_2017,N_756,N_968);
xor U2018 (N_2018,N_937,N_1415);
nor U2019 (N_2019,N_818,N_1167);
or U2020 (N_2020,N_1227,N_1011);
and U2021 (N_2021,N_1396,N_1025);
xor U2022 (N_2022,N_1034,N_1359);
nand U2023 (N_2023,N_1003,N_1023);
xor U2024 (N_2024,N_1244,N_1233);
nor U2025 (N_2025,N_1135,N_962);
or U2026 (N_2026,N_1039,N_1126);
nand U2027 (N_2027,N_1427,N_767);
xnor U2028 (N_2028,N_833,N_1318);
or U2029 (N_2029,N_818,N_1265);
xnor U2030 (N_2030,N_1022,N_1229);
xnor U2031 (N_2031,N_1429,N_1347);
or U2032 (N_2032,N_1433,N_1372);
nand U2033 (N_2033,N_960,N_1477);
or U2034 (N_2034,N_1214,N_1308);
xor U2035 (N_2035,N_1373,N_959);
and U2036 (N_2036,N_1121,N_993);
xnor U2037 (N_2037,N_1297,N_840);
nor U2038 (N_2038,N_1213,N_1438);
and U2039 (N_2039,N_1229,N_775);
or U2040 (N_2040,N_1402,N_1305);
or U2041 (N_2041,N_906,N_976);
xnor U2042 (N_2042,N_934,N_1195);
or U2043 (N_2043,N_1102,N_1431);
xnor U2044 (N_2044,N_1035,N_1288);
or U2045 (N_2045,N_1041,N_1012);
and U2046 (N_2046,N_974,N_1089);
nor U2047 (N_2047,N_1061,N_780);
or U2048 (N_2048,N_964,N_954);
or U2049 (N_2049,N_1042,N_1329);
nand U2050 (N_2050,N_1059,N_1413);
xor U2051 (N_2051,N_1084,N_1478);
and U2052 (N_2052,N_1071,N_1442);
nor U2053 (N_2053,N_806,N_1428);
or U2054 (N_2054,N_837,N_1019);
nor U2055 (N_2055,N_1222,N_801);
xor U2056 (N_2056,N_870,N_1140);
nand U2057 (N_2057,N_1114,N_1337);
nor U2058 (N_2058,N_957,N_839);
and U2059 (N_2059,N_1283,N_1203);
or U2060 (N_2060,N_1404,N_910);
nor U2061 (N_2061,N_755,N_872);
nor U2062 (N_2062,N_1396,N_847);
xor U2063 (N_2063,N_921,N_1140);
and U2064 (N_2064,N_1422,N_908);
and U2065 (N_2065,N_1464,N_831);
nand U2066 (N_2066,N_1261,N_828);
or U2067 (N_2067,N_993,N_1300);
xnor U2068 (N_2068,N_1265,N_763);
xor U2069 (N_2069,N_1004,N_942);
or U2070 (N_2070,N_1219,N_1426);
and U2071 (N_2071,N_893,N_1338);
nand U2072 (N_2072,N_1460,N_1216);
xnor U2073 (N_2073,N_1415,N_823);
nand U2074 (N_2074,N_1481,N_971);
xnor U2075 (N_2075,N_1498,N_1239);
nor U2076 (N_2076,N_836,N_858);
nor U2077 (N_2077,N_783,N_1294);
nor U2078 (N_2078,N_1036,N_854);
nor U2079 (N_2079,N_1211,N_1454);
xor U2080 (N_2080,N_840,N_1216);
and U2081 (N_2081,N_862,N_987);
or U2082 (N_2082,N_1043,N_1437);
nand U2083 (N_2083,N_791,N_873);
or U2084 (N_2084,N_1266,N_886);
xnor U2085 (N_2085,N_779,N_1138);
nor U2086 (N_2086,N_923,N_776);
nor U2087 (N_2087,N_1136,N_933);
nand U2088 (N_2088,N_860,N_861);
xor U2089 (N_2089,N_1288,N_1135);
nor U2090 (N_2090,N_1047,N_948);
nor U2091 (N_2091,N_1188,N_1004);
nand U2092 (N_2092,N_973,N_795);
nor U2093 (N_2093,N_1034,N_1128);
or U2094 (N_2094,N_962,N_1067);
nor U2095 (N_2095,N_1467,N_876);
xor U2096 (N_2096,N_1021,N_897);
xnor U2097 (N_2097,N_1217,N_780);
xnor U2098 (N_2098,N_1154,N_956);
nor U2099 (N_2099,N_1135,N_1153);
xor U2100 (N_2100,N_1309,N_850);
or U2101 (N_2101,N_1440,N_950);
or U2102 (N_2102,N_922,N_821);
or U2103 (N_2103,N_925,N_946);
or U2104 (N_2104,N_1445,N_1010);
nand U2105 (N_2105,N_1121,N_1087);
nand U2106 (N_2106,N_998,N_1195);
and U2107 (N_2107,N_807,N_1313);
nor U2108 (N_2108,N_1253,N_1164);
nand U2109 (N_2109,N_1292,N_1211);
and U2110 (N_2110,N_1081,N_1311);
nand U2111 (N_2111,N_1111,N_1031);
nor U2112 (N_2112,N_798,N_1282);
and U2113 (N_2113,N_756,N_1397);
or U2114 (N_2114,N_1239,N_1009);
xnor U2115 (N_2115,N_949,N_1376);
xor U2116 (N_2116,N_1321,N_1072);
or U2117 (N_2117,N_1340,N_1286);
or U2118 (N_2118,N_989,N_861);
nor U2119 (N_2119,N_947,N_1038);
xnor U2120 (N_2120,N_762,N_826);
or U2121 (N_2121,N_1390,N_868);
xnor U2122 (N_2122,N_795,N_1437);
or U2123 (N_2123,N_1466,N_867);
xor U2124 (N_2124,N_1002,N_1228);
nor U2125 (N_2125,N_1098,N_1176);
nor U2126 (N_2126,N_1087,N_1064);
or U2127 (N_2127,N_1015,N_1156);
nor U2128 (N_2128,N_1313,N_1447);
and U2129 (N_2129,N_778,N_1001);
xnor U2130 (N_2130,N_978,N_941);
xnor U2131 (N_2131,N_1160,N_1263);
or U2132 (N_2132,N_1278,N_777);
nand U2133 (N_2133,N_972,N_1447);
and U2134 (N_2134,N_1375,N_788);
nand U2135 (N_2135,N_1003,N_850);
and U2136 (N_2136,N_871,N_1227);
or U2137 (N_2137,N_1280,N_1444);
and U2138 (N_2138,N_1207,N_1154);
nor U2139 (N_2139,N_802,N_1350);
nor U2140 (N_2140,N_1254,N_843);
or U2141 (N_2141,N_796,N_1073);
or U2142 (N_2142,N_1203,N_888);
nor U2143 (N_2143,N_996,N_1043);
nand U2144 (N_2144,N_1150,N_1337);
and U2145 (N_2145,N_1197,N_1445);
xnor U2146 (N_2146,N_927,N_837);
nand U2147 (N_2147,N_871,N_1248);
or U2148 (N_2148,N_953,N_1490);
nand U2149 (N_2149,N_1085,N_1047);
or U2150 (N_2150,N_1403,N_934);
nand U2151 (N_2151,N_1288,N_802);
nor U2152 (N_2152,N_1234,N_1008);
and U2153 (N_2153,N_1189,N_975);
nand U2154 (N_2154,N_1076,N_1047);
xor U2155 (N_2155,N_1239,N_758);
and U2156 (N_2156,N_1261,N_852);
and U2157 (N_2157,N_1019,N_1274);
nor U2158 (N_2158,N_842,N_959);
nand U2159 (N_2159,N_1477,N_1156);
xor U2160 (N_2160,N_1397,N_1353);
nor U2161 (N_2161,N_1197,N_971);
nor U2162 (N_2162,N_1364,N_1147);
nor U2163 (N_2163,N_1160,N_1142);
xor U2164 (N_2164,N_1474,N_1075);
nor U2165 (N_2165,N_1294,N_1428);
nor U2166 (N_2166,N_929,N_791);
or U2167 (N_2167,N_784,N_1249);
nand U2168 (N_2168,N_1262,N_815);
xnor U2169 (N_2169,N_1210,N_1403);
and U2170 (N_2170,N_884,N_1472);
and U2171 (N_2171,N_1226,N_946);
or U2172 (N_2172,N_1442,N_1091);
nand U2173 (N_2173,N_1379,N_846);
or U2174 (N_2174,N_1231,N_1221);
nand U2175 (N_2175,N_1362,N_978);
nor U2176 (N_2176,N_1433,N_893);
and U2177 (N_2177,N_1210,N_970);
xnor U2178 (N_2178,N_949,N_756);
xor U2179 (N_2179,N_1240,N_893);
or U2180 (N_2180,N_1385,N_1029);
or U2181 (N_2181,N_1382,N_1142);
nor U2182 (N_2182,N_912,N_939);
and U2183 (N_2183,N_981,N_1155);
and U2184 (N_2184,N_937,N_1492);
xor U2185 (N_2185,N_1450,N_1200);
nand U2186 (N_2186,N_1120,N_825);
nand U2187 (N_2187,N_1418,N_1349);
or U2188 (N_2188,N_975,N_1396);
and U2189 (N_2189,N_775,N_1248);
nand U2190 (N_2190,N_1212,N_1354);
xor U2191 (N_2191,N_1311,N_930);
nand U2192 (N_2192,N_1320,N_1352);
xnor U2193 (N_2193,N_886,N_1404);
or U2194 (N_2194,N_1175,N_961);
xnor U2195 (N_2195,N_784,N_957);
nor U2196 (N_2196,N_1355,N_1224);
nand U2197 (N_2197,N_1431,N_1002);
or U2198 (N_2198,N_1176,N_846);
or U2199 (N_2199,N_1380,N_823);
nand U2200 (N_2200,N_1099,N_791);
nand U2201 (N_2201,N_1360,N_883);
nor U2202 (N_2202,N_912,N_1326);
nand U2203 (N_2203,N_792,N_1000);
nand U2204 (N_2204,N_1424,N_1073);
and U2205 (N_2205,N_993,N_1271);
nor U2206 (N_2206,N_767,N_987);
or U2207 (N_2207,N_1281,N_1039);
nand U2208 (N_2208,N_1426,N_1143);
nor U2209 (N_2209,N_887,N_1076);
or U2210 (N_2210,N_867,N_843);
and U2211 (N_2211,N_921,N_941);
nor U2212 (N_2212,N_875,N_1120);
and U2213 (N_2213,N_1363,N_1030);
xnor U2214 (N_2214,N_1401,N_855);
xnor U2215 (N_2215,N_1080,N_832);
xnor U2216 (N_2216,N_1175,N_1094);
nand U2217 (N_2217,N_917,N_1326);
and U2218 (N_2218,N_1149,N_1024);
nor U2219 (N_2219,N_1062,N_923);
nand U2220 (N_2220,N_1029,N_1051);
xor U2221 (N_2221,N_1418,N_1270);
and U2222 (N_2222,N_1310,N_1247);
or U2223 (N_2223,N_1083,N_1082);
or U2224 (N_2224,N_1079,N_1194);
xor U2225 (N_2225,N_1243,N_1474);
and U2226 (N_2226,N_1440,N_1304);
nor U2227 (N_2227,N_1209,N_787);
and U2228 (N_2228,N_849,N_1360);
nand U2229 (N_2229,N_771,N_772);
and U2230 (N_2230,N_1211,N_1093);
or U2231 (N_2231,N_1456,N_1282);
and U2232 (N_2232,N_879,N_1254);
xnor U2233 (N_2233,N_1240,N_1170);
or U2234 (N_2234,N_1307,N_882);
xnor U2235 (N_2235,N_1369,N_1276);
nand U2236 (N_2236,N_1144,N_946);
or U2237 (N_2237,N_911,N_933);
nand U2238 (N_2238,N_751,N_1116);
and U2239 (N_2239,N_1201,N_1321);
nand U2240 (N_2240,N_1159,N_1387);
nor U2241 (N_2241,N_1143,N_1275);
nor U2242 (N_2242,N_1040,N_1227);
and U2243 (N_2243,N_965,N_1089);
xor U2244 (N_2244,N_1243,N_1405);
and U2245 (N_2245,N_1231,N_773);
or U2246 (N_2246,N_839,N_1137);
xor U2247 (N_2247,N_878,N_1189);
or U2248 (N_2248,N_1362,N_1398);
xnor U2249 (N_2249,N_1386,N_895);
and U2250 (N_2250,N_1763,N_1650);
or U2251 (N_2251,N_1896,N_1515);
nand U2252 (N_2252,N_1785,N_1816);
nor U2253 (N_2253,N_1807,N_1502);
nor U2254 (N_2254,N_1843,N_1659);
nand U2255 (N_2255,N_2104,N_1969);
xor U2256 (N_2256,N_1806,N_1715);
or U2257 (N_2257,N_2053,N_2051);
nand U2258 (N_2258,N_1780,N_2159);
nor U2259 (N_2259,N_1908,N_2010);
xor U2260 (N_2260,N_2094,N_1689);
and U2261 (N_2261,N_1724,N_2204);
nor U2262 (N_2262,N_1797,N_1964);
xor U2263 (N_2263,N_1722,N_1586);
xnor U2264 (N_2264,N_1915,N_2167);
and U2265 (N_2265,N_1905,N_1680);
and U2266 (N_2266,N_1948,N_1830);
and U2267 (N_2267,N_1765,N_1539);
or U2268 (N_2268,N_1654,N_1818);
xor U2269 (N_2269,N_1717,N_2004);
and U2270 (N_2270,N_2067,N_2138);
and U2271 (N_2271,N_1546,N_1850);
and U2272 (N_2272,N_1718,N_2030);
or U2273 (N_2273,N_1930,N_1821);
nor U2274 (N_2274,N_1679,N_2171);
xnor U2275 (N_2275,N_1708,N_1662);
xor U2276 (N_2276,N_1879,N_1921);
and U2277 (N_2277,N_2020,N_1699);
and U2278 (N_2278,N_1723,N_1836);
xor U2279 (N_2279,N_1865,N_1660);
and U2280 (N_2280,N_1883,N_1601);
nor U2281 (N_2281,N_1748,N_1968);
nor U2282 (N_2282,N_2113,N_2063);
xnor U2283 (N_2283,N_1619,N_1542);
nand U2284 (N_2284,N_2182,N_1511);
nand U2285 (N_2285,N_2196,N_2207);
or U2286 (N_2286,N_1885,N_2213);
nor U2287 (N_2287,N_2183,N_1953);
nor U2288 (N_2288,N_1752,N_2043);
nand U2289 (N_2289,N_1976,N_2189);
xnor U2290 (N_2290,N_1649,N_2119);
xnor U2291 (N_2291,N_1570,N_1922);
nand U2292 (N_2292,N_1794,N_1656);
and U2293 (N_2293,N_1954,N_2146);
and U2294 (N_2294,N_2118,N_1674);
and U2295 (N_2295,N_1851,N_1558);
nand U2296 (N_2296,N_1683,N_1886);
nand U2297 (N_2297,N_1581,N_1670);
and U2298 (N_2298,N_1913,N_1735);
nand U2299 (N_2299,N_2084,N_1653);
and U2300 (N_2300,N_1661,N_1827);
and U2301 (N_2301,N_1703,N_1860);
xnor U2302 (N_2302,N_1527,N_1629);
nand U2303 (N_2303,N_1852,N_1758);
nor U2304 (N_2304,N_2122,N_1749);
nor U2305 (N_2305,N_1576,N_2247);
nor U2306 (N_2306,N_1872,N_1988);
xor U2307 (N_2307,N_1590,N_1598);
xor U2308 (N_2308,N_1993,N_1516);
nand U2309 (N_2309,N_1589,N_2163);
or U2310 (N_2310,N_2034,N_1652);
nor U2311 (N_2311,N_1769,N_1623);
and U2312 (N_2312,N_1826,N_1991);
xnor U2313 (N_2313,N_1919,N_1588);
nor U2314 (N_2314,N_1644,N_2139);
or U2315 (N_2315,N_1714,N_1880);
or U2316 (N_2316,N_1537,N_2227);
or U2317 (N_2317,N_2150,N_1973);
xor U2318 (N_2318,N_1551,N_1825);
nor U2319 (N_2319,N_1543,N_2086);
and U2320 (N_2320,N_1738,N_1732);
and U2321 (N_2321,N_2080,N_1895);
or U2322 (N_2322,N_1697,N_1974);
nor U2323 (N_2323,N_1664,N_1638);
or U2324 (N_2324,N_1631,N_1521);
or U2325 (N_2325,N_2050,N_2068);
nand U2326 (N_2326,N_1898,N_1873);
or U2327 (N_2327,N_2040,N_2166);
nand U2328 (N_2328,N_1877,N_1848);
nor U2329 (N_2329,N_1986,N_1677);
and U2330 (N_2330,N_1550,N_2237);
and U2331 (N_2331,N_1512,N_1666);
nand U2332 (N_2332,N_1995,N_2110);
nand U2333 (N_2333,N_2126,N_2142);
nor U2334 (N_2334,N_1795,N_2085);
xnor U2335 (N_2335,N_1870,N_2195);
xnor U2336 (N_2336,N_2021,N_1894);
nand U2337 (N_2337,N_2046,N_1610);
nand U2338 (N_2338,N_1582,N_2002);
nand U2339 (N_2339,N_1944,N_1892);
and U2340 (N_2340,N_2107,N_1834);
nand U2341 (N_2341,N_2136,N_1636);
and U2342 (N_2342,N_2135,N_1630);
xnor U2343 (N_2343,N_1632,N_2091);
and U2344 (N_2344,N_2095,N_2064);
or U2345 (N_2345,N_1591,N_1524);
nand U2346 (N_2346,N_1575,N_1997);
nor U2347 (N_2347,N_1801,N_1923);
nor U2348 (N_2348,N_1691,N_1726);
and U2349 (N_2349,N_2203,N_1853);
xnor U2350 (N_2350,N_1561,N_2016);
nand U2351 (N_2351,N_1890,N_1688);
or U2352 (N_2352,N_1784,N_1901);
and U2353 (N_2353,N_1713,N_1909);
or U2354 (N_2354,N_1854,N_1846);
nor U2355 (N_2355,N_1721,N_1531);
or U2356 (N_2356,N_1685,N_2089);
and U2357 (N_2357,N_1538,N_2047);
and U2358 (N_2358,N_2137,N_1599);
and U2359 (N_2359,N_1560,N_2200);
nor U2360 (N_2360,N_1771,N_1557);
or U2361 (N_2361,N_1869,N_1505);
nand U2362 (N_2362,N_1960,N_1866);
xnor U2363 (N_2363,N_2023,N_1907);
xnor U2364 (N_2364,N_2233,N_1779);
xor U2365 (N_2365,N_1967,N_1868);
nand U2366 (N_2366,N_2031,N_2129);
xnor U2367 (N_2367,N_2014,N_1978);
and U2368 (N_2368,N_1965,N_2108);
nand U2369 (N_2369,N_2155,N_1528);
and U2370 (N_2370,N_1642,N_1882);
nor U2371 (N_2371,N_1935,N_2032);
or U2372 (N_2372,N_1768,N_1867);
and U2373 (N_2373,N_1809,N_1700);
and U2374 (N_2374,N_2199,N_2071);
and U2375 (N_2375,N_2222,N_2097);
nand U2376 (N_2376,N_2215,N_2123);
nor U2377 (N_2377,N_1747,N_2157);
and U2378 (N_2378,N_2147,N_2012);
nand U2379 (N_2379,N_2039,N_1663);
xnor U2380 (N_2380,N_1501,N_2077);
xnor U2381 (N_2381,N_1676,N_1789);
xor U2382 (N_2382,N_2038,N_1634);
and U2383 (N_2383,N_1686,N_2160);
and U2384 (N_2384,N_1962,N_1972);
and U2385 (N_2385,N_1567,N_2178);
nor U2386 (N_2386,N_2078,N_2114);
nand U2387 (N_2387,N_1932,N_1790);
xor U2388 (N_2388,N_1861,N_1568);
nand U2389 (N_2389,N_2045,N_1817);
xor U2390 (N_2390,N_2090,N_1504);
xor U2391 (N_2391,N_1767,N_1753);
nand U2392 (N_2392,N_1966,N_2061);
and U2393 (N_2393,N_1849,N_1645);
nor U2394 (N_2394,N_1600,N_1984);
nand U2395 (N_2395,N_2223,N_1982);
nand U2396 (N_2396,N_1667,N_1971);
and U2397 (N_2397,N_2056,N_2141);
or U2398 (N_2398,N_2060,N_2205);
or U2399 (N_2399,N_1938,N_1555);
nor U2400 (N_2400,N_1863,N_2172);
and U2401 (N_2401,N_1940,N_1937);
and U2402 (N_2402,N_2239,N_1736);
nor U2403 (N_2403,N_1627,N_1594);
or U2404 (N_2404,N_1742,N_2101);
or U2405 (N_2405,N_1727,N_2028);
nor U2406 (N_2406,N_1888,N_1673);
and U2407 (N_2407,N_2217,N_1605);
nor U2408 (N_2408,N_2076,N_2226);
and U2409 (N_2409,N_1757,N_1719);
nor U2410 (N_2410,N_1616,N_1773);
and U2411 (N_2411,N_1633,N_1712);
and U2412 (N_2412,N_1815,N_2069);
and U2413 (N_2413,N_1730,N_2022);
xnor U2414 (N_2414,N_2165,N_1945);
or U2415 (N_2415,N_1977,N_1927);
nor U2416 (N_2416,N_1777,N_2121);
xnor U2417 (N_2417,N_1658,N_1517);
nor U2418 (N_2418,N_2229,N_2162);
nor U2419 (N_2419,N_1548,N_1609);
and U2420 (N_2420,N_2209,N_1637);
or U2421 (N_2421,N_2065,N_1625);
or U2422 (N_2422,N_1696,N_1597);
xor U2423 (N_2423,N_1547,N_2170);
nor U2424 (N_2424,N_2211,N_1914);
xor U2425 (N_2425,N_1731,N_1793);
nor U2426 (N_2426,N_2099,N_1740);
xnor U2427 (N_2427,N_2049,N_2009);
nand U2428 (N_2428,N_1733,N_2241);
and U2429 (N_2429,N_1655,N_1545);
and U2430 (N_2430,N_2216,N_1618);
xor U2431 (N_2431,N_1862,N_1620);
xnor U2432 (N_2432,N_1856,N_1711);
xor U2433 (N_2433,N_2242,N_1871);
nand U2434 (N_2434,N_1897,N_1509);
or U2435 (N_2435,N_2100,N_1554);
or U2436 (N_2436,N_1626,N_1621);
xor U2437 (N_2437,N_2088,N_2194);
xnor U2438 (N_2438,N_1580,N_1955);
and U2439 (N_2439,N_1884,N_1902);
or U2440 (N_2440,N_1690,N_1893);
xnor U2441 (N_2441,N_2231,N_1952);
nand U2442 (N_2442,N_1613,N_1530);
xnor U2443 (N_2443,N_2026,N_2057);
nor U2444 (N_2444,N_1604,N_1762);
xor U2445 (N_2445,N_1682,N_2234);
or U2446 (N_2446,N_1774,N_2249);
nor U2447 (N_2447,N_1936,N_2192);
xnor U2448 (N_2448,N_2072,N_1958);
nand U2449 (N_2449,N_1819,N_1624);
or U2450 (N_2450,N_2131,N_2149);
and U2451 (N_2451,N_1508,N_2143);
and U2452 (N_2452,N_1611,N_1615);
nand U2453 (N_2453,N_2188,N_1864);
nand U2454 (N_2454,N_2001,N_2158);
xor U2455 (N_2455,N_2175,N_1549);
and U2456 (N_2456,N_1787,N_1529);
or U2457 (N_2457,N_1845,N_1559);
or U2458 (N_2458,N_1603,N_2082);
nor U2459 (N_2459,N_1791,N_1985);
or U2460 (N_2460,N_1887,N_1566);
or U2461 (N_2461,N_1800,N_1841);
and U2462 (N_2462,N_2134,N_1904);
or U2463 (N_2463,N_1743,N_2116);
or U2464 (N_2464,N_2236,N_2228);
and U2465 (N_2465,N_1999,N_1987);
nand U2466 (N_2466,N_1577,N_1705);
nand U2467 (N_2467,N_1755,N_1823);
nand U2468 (N_2468,N_2066,N_1716);
nand U2469 (N_2469,N_1992,N_1593);
nor U2470 (N_2470,N_1961,N_1617);
xor U2471 (N_2471,N_2218,N_2235);
xnor U2472 (N_2472,N_1831,N_1776);
nand U2473 (N_2473,N_1729,N_2240);
and U2474 (N_2474,N_1553,N_2024);
nor U2475 (N_2475,N_1595,N_2059);
nor U2476 (N_2476,N_1500,N_2062);
and U2477 (N_2477,N_2036,N_1647);
xnor U2478 (N_2478,N_1878,N_1983);
xor U2479 (N_2479,N_1641,N_2106);
nand U2480 (N_2480,N_1507,N_1701);
nand U2481 (N_2481,N_1926,N_1764);
nand U2482 (N_2482,N_1788,N_1684);
xnor U2483 (N_2483,N_1704,N_2103);
nand U2484 (N_2484,N_2187,N_1710);
nor U2485 (N_2485,N_1906,N_1772);
or U2486 (N_2486,N_1796,N_2245);
xor U2487 (N_2487,N_1759,N_2221);
nand U2488 (N_2488,N_1891,N_2007);
xor U2489 (N_2489,N_2055,N_1635);
and U2490 (N_2490,N_1881,N_2130);
or U2491 (N_2491,N_2093,N_1828);
nand U2492 (N_2492,N_1824,N_1996);
xor U2493 (N_2493,N_1859,N_1844);
and U2494 (N_2494,N_2058,N_1837);
nor U2495 (N_2495,N_1858,N_1675);
xor U2496 (N_2496,N_2140,N_1963);
and U2497 (N_2497,N_1565,N_1707);
xor U2498 (N_2498,N_1681,N_1916);
nand U2499 (N_2499,N_2161,N_2180);
or U2500 (N_2500,N_2185,N_2193);
xor U2501 (N_2501,N_1933,N_1770);
nor U2502 (N_2502,N_2246,N_1744);
or U2503 (N_2503,N_1563,N_2115);
nor U2504 (N_2504,N_2079,N_2151);
nor U2505 (N_2505,N_1783,N_1875);
nor U2506 (N_2506,N_1781,N_2224);
nand U2507 (N_2507,N_1737,N_2073);
nand U2508 (N_2508,N_1510,N_1669);
nand U2509 (N_2509,N_1556,N_2176);
xnor U2510 (N_2510,N_2190,N_1693);
nand U2511 (N_2511,N_2052,N_1812);
nand U2512 (N_2512,N_2128,N_2003);
nor U2513 (N_2513,N_2173,N_2181);
and U2514 (N_2514,N_2238,N_2035);
or U2515 (N_2515,N_1678,N_2109);
nand U2516 (N_2516,N_1842,N_1799);
and U2517 (N_2517,N_2054,N_1741);
and U2518 (N_2518,N_2210,N_1622);
nor U2519 (N_2519,N_1728,N_1998);
xor U2520 (N_2520,N_1506,N_1518);
nand U2521 (N_2521,N_1924,N_1946);
nand U2522 (N_2522,N_1803,N_2015);
xnor U2523 (N_2523,N_1949,N_1750);
xnor U2524 (N_2524,N_1651,N_2202);
nor U2525 (N_2525,N_1928,N_2042);
nor U2526 (N_2526,N_1592,N_1668);
and U2527 (N_2527,N_1950,N_1792);
nand U2528 (N_2528,N_1646,N_2144);
nor U2529 (N_2529,N_1573,N_1709);
and U2530 (N_2530,N_1602,N_1943);
nor U2531 (N_2531,N_1813,N_2017);
nor U2532 (N_2532,N_1571,N_1990);
xnor U2533 (N_2533,N_2197,N_2184);
and U2534 (N_2534,N_1811,N_1534);
nand U2535 (N_2535,N_1912,N_1725);
and U2536 (N_2536,N_1694,N_1734);
and U2537 (N_2537,N_1931,N_2156);
xnor U2538 (N_2538,N_1766,N_1775);
or U2539 (N_2539,N_1840,N_2008);
nor U2540 (N_2540,N_2125,N_1918);
or U2541 (N_2541,N_1939,N_2244);
nor U2542 (N_2542,N_1564,N_2033);
and U2543 (N_2543,N_2225,N_2198);
or U2544 (N_2544,N_1910,N_2111);
and U2545 (N_2545,N_1628,N_1925);
and U2546 (N_2546,N_1804,N_2092);
or U2547 (N_2547,N_1941,N_1739);
or U2548 (N_2548,N_1643,N_1980);
or U2549 (N_2549,N_2041,N_1596);
or U2550 (N_2550,N_1706,N_1900);
nand U2551 (N_2551,N_1981,N_2191);
nor U2552 (N_2552,N_2152,N_2081);
nor U2553 (N_2553,N_1698,N_1513);
nor U2554 (N_2554,N_1526,N_1665);
nand U2555 (N_2555,N_2018,N_1520);
nor U2556 (N_2556,N_1754,N_1874);
nor U2557 (N_2557,N_1857,N_2248);
nand U2558 (N_2558,N_1720,N_2075);
xor U2559 (N_2559,N_1970,N_2120);
nand U2560 (N_2560,N_2153,N_1745);
or U2561 (N_2561,N_1947,N_1798);
nor U2562 (N_2562,N_1687,N_2005);
and U2563 (N_2563,N_2117,N_1522);
nor U2564 (N_2564,N_1917,N_2025);
nand U2565 (N_2565,N_2102,N_1756);
or U2566 (N_2566,N_1929,N_2029);
nand U2567 (N_2567,N_1503,N_1514);
xor U2568 (N_2568,N_1778,N_1648);
xor U2569 (N_2569,N_1523,N_1786);
nor U2570 (N_2570,N_2169,N_2208);
xor U2571 (N_2571,N_2174,N_1585);
or U2572 (N_2572,N_2164,N_2044);
nor U2573 (N_2573,N_1607,N_1671);
nor U2574 (N_2574,N_1672,N_2124);
nor U2575 (N_2575,N_2127,N_1572);
nand U2576 (N_2576,N_2214,N_1805);
and U2577 (N_2577,N_2132,N_1535);
and U2578 (N_2578,N_1994,N_1899);
nor U2579 (N_2579,N_1934,N_1957);
nor U2580 (N_2580,N_1839,N_2168);
xor U2581 (N_2581,N_1889,N_2027);
nand U2582 (N_2582,N_1657,N_1536);
and U2583 (N_2583,N_1583,N_2006);
xor U2584 (N_2584,N_2011,N_1562);
nor U2585 (N_2585,N_1835,N_2186);
or U2586 (N_2586,N_1606,N_1832);
nor U2587 (N_2587,N_1847,N_2048);
nor U2588 (N_2588,N_1608,N_1833);
and U2589 (N_2589,N_2070,N_2206);
nand U2590 (N_2590,N_1519,N_1920);
or U2591 (N_2591,N_1951,N_1574);
or U2592 (N_2592,N_2243,N_1702);
or U2593 (N_2593,N_1956,N_2133);
or U2594 (N_2594,N_1584,N_1829);
nor U2595 (N_2595,N_1525,N_2013);
nand U2596 (N_2596,N_1810,N_2148);
nand U2597 (N_2597,N_1541,N_1578);
nor U2598 (N_2598,N_1569,N_1820);
or U2599 (N_2599,N_1692,N_1838);
xor U2600 (N_2600,N_2037,N_2083);
nor U2601 (N_2601,N_1975,N_2230);
and U2602 (N_2602,N_1761,N_2000);
nor U2603 (N_2603,N_1760,N_1822);
and U2604 (N_2604,N_1959,N_2177);
nand U2605 (N_2605,N_1552,N_1911);
xor U2606 (N_2606,N_2105,N_1782);
nand U2607 (N_2607,N_1855,N_1808);
or U2608 (N_2608,N_2212,N_2087);
nor U2609 (N_2609,N_2232,N_1942);
and U2610 (N_2610,N_2019,N_2074);
or U2611 (N_2611,N_1814,N_1540);
xnor U2612 (N_2612,N_1587,N_2220);
or U2613 (N_2613,N_1640,N_1639);
nor U2614 (N_2614,N_2219,N_1544);
and U2615 (N_2615,N_1612,N_1876);
nand U2616 (N_2616,N_1903,N_2154);
nor U2617 (N_2617,N_2096,N_1533);
and U2618 (N_2618,N_1532,N_2179);
nor U2619 (N_2619,N_1979,N_1579);
xor U2620 (N_2620,N_1695,N_1614);
and U2621 (N_2621,N_2201,N_1802);
or U2622 (N_2622,N_2145,N_2098);
and U2623 (N_2623,N_1746,N_1989);
and U2624 (N_2624,N_1751,N_2112);
and U2625 (N_2625,N_1910,N_1861);
xor U2626 (N_2626,N_2177,N_2104);
and U2627 (N_2627,N_1648,N_2157);
nand U2628 (N_2628,N_1686,N_1746);
and U2629 (N_2629,N_2142,N_1832);
xor U2630 (N_2630,N_2036,N_1910);
or U2631 (N_2631,N_2024,N_1609);
xor U2632 (N_2632,N_2047,N_2063);
or U2633 (N_2633,N_1607,N_1602);
nand U2634 (N_2634,N_1706,N_2093);
xnor U2635 (N_2635,N_2162,N_1650);
and U2636 (N_2636,N_1992,N_1658);
xor U2637 (N_2637,N_1571,N_1831);
or U2638 (N_2638,N_2078,N_1883);
nor U2639 (N_2639,N_2124,N_1891);
nand U2640 (N_2640,N_2184,N_1800);
nor U2641 (N_2641,N_2228,N_1879);
or U2642 (N_2642,N_2234,N_1721);
nand U2643 (N_2643,N_1724,N_1679);
nand U2644 (N_2644,N_1965,N_2117);
or U2645 (N_2645,N_2101,N_1842);
xnor U2646 (N_2646,N_1596,N_1713);
and U2647 (N_2647,N_1999,N_1644);
nor U2648 (N_2648,N_1826,N_1714);
xnor U2649 (N_2649,N_2231,N_1855);
xnor U2650 (N_2650,N_1887,N_1763);
xor U2651 (N_2651,N_1753,N_2117);
nand U2652 (N_2652,N_1769,N_2015);
nor U2653 (N_2653,N_1856,N_1517);
or U2654 (N_2654,N_1505,N_1911);
xnor U2655 (N_2655,N_1512,N_1926);
or U2656 (N_2656,N_2235,N_1772);
nand U2657 (N_2657,N_1745,N_2115);
or U2658 (N_2658,N_1969,N_1877);
xnor U2659 (N_2659,N_2044,N_1918);
nand U2660 (N_2660,N_2066,N_2223);
nor U2661 (N_2661,N_1722,N_1780);
or U2662 (N_2662,N_1812,N_2243);
or U2663 (N_2663,N_2094,N_2197);
nand U2664 (N_2664,N_1953,N_2249);
nor U2665 (N_2665,N_1502,N_1680);
nor U2666 (N_2666,N_2041,N_2138);
nand U2667 (N_2667,N_1626,N_1671);
xor U2668 (N_2668,N_2169,N_2069);
nor U2669 (N_2669,N_1874,N_1768);
and U2670 (N_2670,N_1602,N_1637);
nand U2671 (N_2671,N_2005,N_1976);
and U2672 (N_2672,N_2203,N_1804);
and U2673 (N_2673,N_2116,N_1614);
nand U2674 (N_2674,N_1829,N_2047);
or U2675 (N_2675,N_1759,N_1719);
nand U2676 (N_2676,N_1809,N_1510);
nand U2677 (N_2677,N_1969,N_2245);
nand U2678 (N_2678,N_1653,N_1989);
xnor U2679 (N_2679,N_1798,N_1754);
xnor U2680 (N_2680,N_1619,N_2018);
and U2681 (N_2681,N_2209,N_1717);
or U2682 (N_2682,N_1942,N_1864);
nor U2683 (N_2683,N_1700,N_1578);
nand U2684 (N_2684,N_1911,N_2223);
or U2685 (N_2685,N_1935,N_2159);
nand U2686 (N_2686,N_1834,N_2184);
or U2687 (N_2687,N_2065,N_1554);
nor U2688 (N_2688,N_1611,N_2233);
or U2689 (N_2689,N_2184,N_1564);
nand U2690 (N_2690,N_1641,N_2196);
nor U2691 (N_2691,N_1512,N_1656);
or U2692 (N_2692,N_1805,N_1770);
nor U2693 (N_2693,N_1989,N_1529);
nand U2694 (N_2694,N_1727,N_2009);
or U2695 (N_2695,N_2127,N_2214);
and U2696 (N_2696,N_1623,N_1519);
nand U2697 (N_2697,N_1690,N_1779);
nor U2698 (N_2698,N_1900,N_2028);
and U2699 (N_2699,N_2110,N_1914);
and U2700 (N_2700,N_1687,N_1881);
nand U2701 (N_2701,N_2235,N_1921);
and U2702 (N_2702,N_1915,N_1727);
or U2703 (N_2703,N_1956,N_1780);
xnor U2704 (N_2704,N_1532,N_1985);
nand U2705 (N_2705,N_1782,N_2119);
nor U2706 (N_2706,N_1571,N_1737);
xnor U2707 (N_2707,N_1913,N_1505);
nand U2708 (N_2708,N_2205,N_2240);
nand U2709 (N_2709,N_1782,N_2162);
nand U2710 (N_2710,N_1853,N_2037);
nor U2711 (N_2711,N_2113,N_2071);
nand U2712 (N_2712,N_2234,N_1618);
or U2713 (N_2713,N_1611,N_2014);
nor U2714 (N_2714,N_1800,N_2145);
nor U2715 (N_2715,N_1673,N_1989);
or U2716 (N_2716,N_1639,N_1775);
or U2717 (N_2717,N_1952,N_1883);
or U2718 (N_2718,N_2067,N_1789);
nand U2719 (N_2719,N_1640,N_1506);
nand U2720 (N_2720,N_1871,N_2012);
and U2721 (N_2721,N_2100,N_1933);
and U2722 (N_2722,N_1976,N_1912);
nand U2723 (N_2723,N_2064,N_1881);
or U2724 (N_2724,N_2115,N_1800);
or U2725 (N_2725,N_2091,N_1582);
nand U2726 (N_2726,N_1532,N_1627);
and U2727 (N_2727,N_1760,N_2039);
nor U2728 (N_2728,N_2165,N_1910);
or U2729 (N_2729,N_1656,N_1537);
xor U2730 (N_2730,N_2206,N_2239);
or U2731 (N_2731,N_2149,N_1602);
nand U2732 (N_2732,N_2062,N_1742);
or U2733 (N_2733,N_2166,N_1986);
nand U2734 (N_2734,N_1854,N_2163);
or U2735 (N_2735,N_1957,N_1602);
or U2736 (N_2736,N_1857,N_2084);
xnor U2737 (N_2737,N_2073,N_1773);
nand U2738 (N_2738,N_2089,N_1532);
or U2739 (N_2739,N_2015,N_1888);
nand U2740 (N_2740,N_2156,N_1781);
and U2741 (N_2741,N_1621,N_1557);
nand U2742 (N_2742,N_2117,N_1782);
or U2743 (N_2743,N_1552,N_2054);
nor U2744 (N_2744,N_1782,N_1861);
xor U2745 (N_2745,N_2032,N_1899);
nor U2746 (N_2746,N_1883,N_1787);
xnor U2747 (N_2747,N_2229,N_2037);
nand U2748 (N_2748,N_1511,N_1627);
xnor U2749 (N_2749,N_1568,N_1775);
xor U2750 (N_2750,N_2006,N_2015);
nor U2751 (N_2751,N_1504,N_1852);
nand U2752 (N_2752,N_2165,N_1907);
or U2753 (N_2753,N_1932,N_1822);
and U2754 (N_2754,N_2079,N_1967);
and U2755 (N_2755,N_1985,N_2236);
nor U2756 (N_2756,N_2063,N_1687);
nand U2757 (N_2757,N_2137,N_1778);
nor U2758 (N_2758,N_1754,N_1888);
or U2759 (N_2759,N_1881,N_1878);
xnor U2760 (N_2760,N_1710,N_1518);
xnor U2761 (N_2761,N_2182,N_2003);
xnor U2762 (N_2762,N_2023,N_1689);
and U2763 (N_2763,N_1702,N_1642);
and U2764 (N_2764,N_2041,N_1595);
nor U2765 (N_2765,N_1685,N_1989);
nor U2766 (N_2766,N_2092,N_2010);
xor U2767 (N_2767,N_1930,N_1844);
nand U2768 (N_2768,N_1827,N_1972);
or U2769 (N_2769,N_1615,N_1724);
or U2770 (N_2770,N_1560,N_2009);
nor U2771 (N_2771,N_2169,N_1968);
nand U2772 (N_2772,N_2059,N_1666);
nor U2773 (N_2773,N_2159,N_2033);
and U2774 (N_2774,N_1807,N_1513);
nand U2775 (N_2775,N_2113,N_1695);
and U2776 (N_2776,N_1803,N_2221);
and U2777 (N_2777,N_1612,N_1995);
xor U2778 (N_2778,N_2218,N_1736);
and U2779 (N_2779,N_1945,N_2191);
nand U2780 (N_2780,N_2028,N_2006);
nand U2781 (N_2781,N_1637,N_1646);
and U2782 (N_2782,N_1824,N_1965);
and U2783 (N_2783,N_1741,N_1819);
and U2784 (N_2784,N_2032,N_1849);
and U2785 (N_2785,N_1516,N_1505);
and U2786 (N_2786,N_1643,N_1877);
or U2787 (N_2787,N_1718,N_1819);
xor U2788 (N_2788,N_1919,N_1545);
or U2789 (N_2789,N_2056,N_1956);
xor U2790 (N_2790,N_2076,N_1684);
and U2791 (N_2791,N_1884,N_1988);
xnor U2792 (N_2792,N_1620,N_2008);
xor U2793 (N_2793,N_1747,N_1865);
nor U2794 (N_2794,N_1557,N_2076);
nand U2795 (N_2795,N_1918,N_1829);
xnor U2796 (N_2796,N_2057,N_1852);
and U2797 (N_2797,N_2074,N_2107);
and U2798 (N_2798,N_2067,N_2032);
and U2799 (N_2799,N_2171,N_1771);
or U2800 (N_2800,N_1746,N_1755);
and U2801 (N_2801,N_1749,N_1710);
and U2802 (N_2802,N_1793,N_1711);
nor U2803 (N_2803,N_1778,N_1659);
and U2804 (N_2804,N_1882,N_1580);
xor U2805 (N_2805,N_1847,N_2193);
or U2806 (N_2806,N_2197,N_1525);
nor U2807 (N_2807,N_1879,N_2103);
xnor U2808 (N_2808,N_2197,N_2025);
and U2809 (N_2809,N_1912,N_2238);
nand U2810 (N_2810,N_1540,N_1703);
or U2811 (N_2811,N_1879,N_2235);
nand U2812 (N_2812,N_2012,N_2071);
nand U2813 (N_2813,N_1825,N_1978);
and U2814 (N_2814,N_1755,N_1867);
xnor U2815 (N_2815,N_1745,N_1668);
and U2816 (N_2816,N_2155,N_1723);
or U2817 (N_2817,N_1886,N_2000);
xor U2818 (N_2818,N_1750,N_2105);
nand U2819 (N_2819,N_2110,N_1830);
nor U2820 (N_2820,N_2116,N_2171);
xor U2821 (N_2821,N_1938,N_2130);
nor U2822 (N_2822,N_2091,N_1505);
or U2823 (N_2823,N_1684,N_1671);
and U2824 (N_2824,N_1518,N_2056);
nand U2825 (N_2825,N_1694,N_1547);
nand U2826 (N_2826,N_1532,N_1785);
and U2827 (N_2827,N_2029,N_1636);
nor U2828 (N_2828,N_1731,N_1785);
xor U2829 (N_2829,N_1593,N_1876);
nand U2830 (N_2830,N_1672,N_2225);
nand U2831 (N_2831,N_2115,N_2149);
nor U2832 (N_2832,N_1778,N_1643);
nor U2833 (N_2833,N_2226,N_1945);
or U2834 (N_2834,N_1967,N_1579);
nand U2835 (N_2835,N_1504,N_1729);
nor U2836 (N_2836,N_1731,N_1887);
nand U2837 (N_2837,N_1879,N_1571);
and U2838 (N_2838,N_1742,N_1679);
or U2839 (N_2839,N_1778,N_2150);
or U2840 (N_2840,N_1824,N_1679);
xnor U2841 (N_2841,N_1988,N_2059);
and U2842 (N_2842,N_1760,N_1685);
and U2843 (N_2843,N_1935,N_2246);
nor U2844 (N_2844,N_1938,N_2025);
and U2845 (N_2845,N_1843,N_1884);
nand U2846 (N_2846,N_1659,N_2201);
or U2847 (N_2847,N_1551,N_1926);
xor U2848 (N_2848,N_1612,N_2225);
nor U2849 (N_2849,N_1820,N_1759);
nand U2850 (N_2850,N_1505,N_2132);
nor U2851 (N_2851,N_1536,N_2120);
xnor U2852 (N_2852,N_1961,N_1927);
xor U2853 (N_2853,N_2186,N_1542);
or U2854 (N_2854,N_2144,N_1707);
nor U2855 (N_2855,N_1696,N_1831);
xnor U2856 (N_2856,N_2190,N_2127);
nor U2857 (N_2857,N_1717,N_1829);
and U2858 (N_2858,N_1763,N_2049);
or U2859 (N_2859,N_1992,N_1833);
xnor U2860 (N_2860,N_2006,N_1622);
nor U2861 (N_2861,N_2075,N_1976);
nand U2862 (N_2862,N_1847,N_1546);
nor U2863 (N_2863,N_1849,N_2088);
and U2864 (N_2864,N_2071,N_1745);
nor U2865 (N_2865,N_1810,N_1742);
nand U2866 (N_2866,N_2010,N_1800);
and U2867 (N_2867,N_1741,N_1840);
and U2868 (N_2868,N_1874,N_2058);
xor U2869 (N_2869,N_1669,N_1555);
nor U2870 (N_2870,N_1997,N_1926);
or U2871 (N_2871,N_2171,N_1956);
and U2872 (N_2872,N_2245,N_1868);
nor U2873 (N_2873,N_1535,N_1866);
nor U2874 (N_2874,N_1763,N_1709);
or U2875 (N_2875,N_1709,N_1684);
nand U2876 (N_2876,N_1672,N_2203);
nor U2877 (N_2877,N_2181,N_1886);
xnor U2878 (N_2878,N_1635,N_1977);
nand U2879 (N_2879,N_1972,N_1887);
nand U2880 (N_2880,N_1697,N_1783);
or U2881 (N_2881,N_2193,N_1887);
and U2882 (N_2882,N_1963,N_1967);
xor U2883 (N_2883,N_1637,N_2040);
or U2884 (N_2884,N_2085,N_1833);
nand U2885 (N_2885,N_2193,N_1926);
nor U2886 (N_2886,N_2009,N_1592);
nand U2887 (N_2887,N_1642,N_1617);
xor U2888 (N_2888,N_2110,N_2028);
nor U2889 (N_2889,N_2025,N_1637);
nand U2890 (N_2890,N_2021,N_1814);
nor U2891 (N_2891,N_1929,N_1873);
and U2892 (N_2892,N_2056,N_2020);
and U2893 (N_2893,N_1518,N_1508);
nor U2894 (N_2894,N_2125,N_1800);
nor U2895 (N_2895,N_1737,N_1654);
and U2896 (N_2896,N_1717,N_1727);
and U2897 (N_2897,N_1953,N_1942);
or U2898 (N_2898,N_1969,N_1833);
and U2899 (N_2899,N_2003,N_2176);
xor U2900 (N_2900,N_1854,N_2164);
and U2901 (N_2901,N_2232,N_2201);
xor U2902 (N_2902,N_1724,N_1544);
nor U2903 (N_2903,N_1588,N_1818);
xor U2904 (N_2904,N_1958,N_1565);
or U2905 (N_2905,N_2190,N_1533);
and U2906 (N_2906,N_2198,N_1643);
or U2907 (N_2907,N_1627,N_1990);
and U2908 (N_2908,N_1755,N_1545);
nand U2909 (N_2909,N_1578,N_1664);
or U2910 (N_2910,N_1842,N_2099);
and U2911 (N_2911,N_1881,N_1913);
nor U2912 (N_2912,N_1721,N_1527);
nor U2913 (N_2913,N_1842,N_2038);
nor U2914 (N_2914,N_2046,N_1522);
xnor U2915 (N_2915,N_1797,N_2095);
nand U2916 (N_2916,N_1867,N_1662);
or U2917 (N_2917,N_2098,N_1640);
or U2918 (N_2918,N_1571,N_2041);
nor U2919 (N_2919,N_1651,N_1907);
and U2920 (N_2920,N_2148,N_2015);
nor U2921 (N_2921,N_1546,N_1548);
or U2922 (N_2922,N_1922,N_1941);
or U2923 (N_2923,N_1944,N_1714);
nor U2924 (N_2924,N_1594,N_1847);
nor U2925 (N_2925,N_1680,N_2103);
nand U2926 (N_2926,N_1522,N_1700);
nor U2927 (N_2927,N_2086,N_1525);
and U2928 (N_2928,N_2193,N_1671);
nor U2929 (N_2929,N_1696,N_1744);
xnor U2930 (N_2930,N_1770,N_2067);
xor U2931 (N_2931,N_1977,N_1570);
nor U2932 (N_2932,N_1973,N_1653);
nand U2933 (N_2933,N_2085,N_2038);
and U2934 (N_2934,N_1941,N_2070);
nor U2935 (N_2935,N_2047,N_1565);
and U2936 (N_2936,N_2057,N_1839);
xnor U2937 (N_2937,N_2110,N_1500);
nor U2938 (N_2938,N_2094,N_1836);
nand U2939 (N_2939,N_2085,N_1719);
nor U2940 (N_2940,N_1730,N_2194);
nand U2941 (N_2941,N_1981,N_1520);
nor U2942 (N_2942,N_2077,N_2078);
nand U2943 (N_2943,N_2241,N_1862);
xnor U2944 (N_2944,N_1556,N_2130);
xor U2945 (N_2945,N_2198,N_1859);
or U2946 (N_2946,N_1564,N_2120);
and U2947 (N_2947,N_1673,N_1804);
or U2948 (N_2948,N_1767,N_1911);
nor U2949 (N_2949,N_1748,N_2050);
xnor U2950 (N_2950,N_1797,N_2023);
or U2951 (N_2951,N_1837,N_1969);
nor U2952 (N_2952,N_1985,N_1663);
or U2953 (N_2953,N_1933,N_1789);
or U2954 (N_2954,N_1780,N_1591);
and U2955 (N_2955,N_1552,N_1744);
and U2956 (N_2956,N_1610,N_1605);
nand U2957 (N_2957,N_1664,N_1807);
nand U2958 (N_2958,N_2242,N_1601);
nand U2959 (N_2959,N_1772,N_1781);
nand U2960 (N_2960,N_1611,N_1741);
nor U2961 (N_2961,N_2056,N_1791);
nand U2962 (N_2962,N_1640,N_2175);
nor U2963 (N_2963,N_1697,N_2110);
or U2964 (N_2964,N_1547,N_1726);
or U2965 (N_2965,N_2126,N_2067);
nand U2966 (N_2966,N_1784,N_1532);
nor U2967 (N_2967,N_1674,N_1886);
nor U2968 (N_2968,N_1594,N_1518);
and U2969 (N_2969,N_1822,N_2119);
nand U2970 (N_2970,N_1857,N_2141);
and U2971 (N_2971,N_2177,N_1821);
or U2972 (N_2972,N_1887,N_1546);
xnor U2973 (N_2973,N_1840,N_2127);
or U2974 (N_2974,N_1614,N_2128);
nor U2975 (N_2975,N_1656,N_2047);
nor U2976 (N_2976,N_1909,N_1536);
xor U2977 (N_2977,N_1745,N_1764);
or U2978 (N_2978,N_1928,N_1555);
xor U2979 (N_2979,N_1634,N_1533);
nor U2980 (N_2980,N_1587,N_1581);
and U2981 (N_2981,N_1559,N_2220);
and U2982 (N_2982,N_1552,N_1922);
xor U2983 (N_2983,N_1502,N_2171);
xor U2984 (N_2984,N_2185,N_2236);
and U2985 (N_2985,N_1561,N_2117);
or U2986 (N_2986,N_1926,N_2196);
or U2987 (N_2987,N_2127,N_1667);
xnor U2988 (N_2988,N_1873,N_2119);
xnor U2989 (N_2989,N_1871,N_1907);
xnor U2990 (N_2990,N_1589,N_1922);
or U2991 (N_2991,N_2173,N_1899);
nor U2992 (N_2992,N_1985,N_1584);
or U2993 (N_2993,N_1601,N_1802);
xor U2994 (N_2994,N_2243,N_2043);
xnor U2995 (N_2995,N_2168,N_1620);
and U2996 (N_2996,N_2223,N_1530);
and U2997 (N_2997,N_2047,N_1591);
xor U2998 (N_2998,N_1821,N_2046);
and U2999 (N_2999,N_2249,N_2158);
nand U3000 (N_3000,N_2825,N_2656);
nand U3001 (N_3001,N_2351,N_2484);
nand U3002 (N_3002,N_2695,N_2383);
or U3003 (N_3003,N_2456,N_2890);
nand U3004 (N_3004,N_2437,N_2726);
nor U3005 (N_3005,N_2862,N_2812);
nand U3006 (N_3006,N_2655,N_2733);
xnor U3007 (N_3007,N_2700,N_2849);
and U3008 (N_3008,N_2837,N_2449);
xnor U3009 (N_3009,N_2791,N_2478);
nor U3010 (N_3010,N_2601,N_2672);
and U3011 (N_3011,N_2707,N_2839);
nand U3012 (N_3012,N_2856,N_2471);
nand U3013 (N_3013,N_2539,N_2399);
xor U3014 (N_3014,N_2586,N_2336);
or U3015 (N_3015,N_2271,N_2516);
and U3016 (N_3016,N_2703,N_2795);
and U3017 (N_3017,N_2773,N_2623);
and U3018 (N_3018,N_2536,N_2507);
nand U3019 (N_3019,N_2296,N_2658);
nand U3020 (N_3020,N_2528,N_2662);
and U3021 (N_3021,N_2250,N_2879);
nor U3022 (N_3022,N_2769,N_2923);
nor U3023 (N_3023,N_2360,N_2522);
xor U3024 (N_3024,N_2397,N_2706);
nor U3025 (N_3025,N_2266,N_2572);
nor U3026 (N_3026,N_2465,N_2431);
nand U3027 (N_3027,N_2318,N_2817);
and U3028 (N_3028,N_2993,N_2282);
and U3029 (N_3029,N_2682,N_2367);
xor U3030 (N_3030,N_2571,N_2736);
nor U3031 (N_3031,N_2622,N_2480);
nand U3032 (N_3032,N_2959,N_2541);
xnor U3033 (N_3033,N_2713,N_2928);
nor U3034 (N_3034,N_2676,N_2389);
nor U3035 (N_3035,N_2366,N_2967);
or U3036 (N_3036,N_2816,N_2467);
xnor U3037 (N_3037,N_2438,N_2691);
xnor U3038 (N_3038,N_2504,N_2954);
xor U3039 (N_3039,N_2882,N_2529);
nor U3040 (N_3040,N_2569,N_2908);
and U3041 (N_3041,N_2960,N_2759);
xnor U3042 (N_3042,N_2711,N_2457);
or U3043 (N_3043,N_2341,N_2941);
nor U3044 (N_3044,N_2517,N_2490);
nor U3045 (N_3045,N_2940,N_2981);
and U3046 (N_3046,N_2998,N_2428);
xnor U3047 (N_3047,N_2270,N_2258);
or U3048 (N_3048,N_2446,N_2283);
nor U3049 (N_3049,N_2485,N_2920);
nor U3050 (N_3050,N_2558,N_2990);
xor U3051 (N_3051,N_2398,N_2820);
xor U3052 (N_3052,N_2393,N_2810);
and U3053 (N_3053,N_2892,N_2802);
nor U3054 (N_3054,N_2272,N_2740);
nor U3055 (N_3055,N_2780,N_2945);
and U3056 (N_3056,N_2306,N_2727);
nor U3057 (N_3057,N_2347,N_2563);
nor U3058 (N_3058,N_2801,N_2657);
nand U3059 (N_3059,N_2404,N_2771);
nor U3060 (N_3060,N_2909,N_2374);
and U3061 (N_3061,N_2854,N_2865);
nand U3062 (N_3062,N_2997,N_2363);
and U3063 (N_3063,N_2721,N_2723);
or U3064 (N_3064,N_2503,N_2352);
nand U3065 (N_3065,N_2524,N_2551);
nand U3066 (N_3066,N_2262,N_2679);
nor U3067 (N_3067,N_2819,N_2957);
or U3068 (N_3068,N_2387,N_2379);
nand U3069 (N_3069,N_2894,N_2337);
xor U3070 (N_3070,N_2953,N_2520);
nor U3071 (N_3071,N_2423,N_2553);
and U3072 (N_3072,N_2312,N_2823);
nor U3073 (N_3073,N_2858,N_2965);
nand U3074 (N_3074,N_2895,N_2749);
or U3075 (N_3075,N_2978,N_2492);
nor U3076 (N_3076,N_2372,N_2401);
or U3077 (N_3077,N_2932,N_2639);
xnor U3078 (N_3078,N_2955,N_2434);
nand U3079 (N_3079,N_2712,N_2716);
nand U3080 (N_3080,N_2991,N_2265);
or U3081 (N_3081,N_2883,N_2783);
or U3082 (N_3082,N_2540,N_2976);
nor U3083 (N_3083,N_2566,N_2380);
nor U3084 (N_3084,N_2725,N_2884);
nand U3085 (N_3085,N_2453,N_2979);
or U3086 (N_3086,N_2370,N_2581);
or U3087 (N_3087,N_2415,N_2869);
nand U3088 (N_3088,N_2530,N_2995);
xor U3089 (N_3089,N_2373,N_2785);
xor U3090 (N_3090,N_2589,N_2252);
or U3091 (N_3091,N_2324,N_2685);
and U3092 (N_3092,N_2844,N_2444);
nor U3093 (N_3093,N_2325,N_2512);
and U3094 (N_3094,N_2307,N_2973);
nor U3095 (N_3095,N_2760,N_2546);
nand U3096 (N_3096,N_2793,N_2537);
nand U3097 (N_3097,N_2510,N_2410);
nor U3098 (N_3098,N_2321,N_2877);
or U3099 (N_3099,N_2855,N_2396);
xnor U3100 (N_3100,N_2643,N_2582);
or U3101 (N_3101,N_2259,N_2843);
nand U3102 (N_3102,N_2511,N_2746);
nor U3103 (N_3103,N_2634,N_2915);
nand U3104 (N_3104,N_2278,N_2319);
nor U3105 (N_3105,N_2591,N_2413);
xnor U3106 (N_3106,N_2481,N_2277);
nand U3107 (N_3107,N_2600,N_2982);
or U3108 (N_3108,N_2489,N_2905);
xor U3109 (N_3109,N_2356,N_2803);
and U3110 (N_3110,N_2742,N_2487);
xor U3111 (N_3111,N_2650,N_2758);
nor U3112 (N_3112,N_2432,N_2964);
and U3113 (N_3113,N_2901,N_2867);
nand U3114 (N_3114,N_2702,N_2663);
nand U3115 (N_3115,N_2382,N_2753);
nor U3116 (N_3116,N_2464,N_2888);
nor U3117 (N_3117,N_2354,N_2564);
and U3118 (N_3118,N_2988,N_2458);
or U3119 (N_3119,N_2309,N_2267);
or U3120 (N_3120,N_2784,N_2754);
nor U3121 (N_3121,N_2942,N_2521);
and U3122 (N_3122,N_2949,N_2455);
nand U3123 (N_3123,N_2255,N_2575);
xor U3124 (N_3124,N_2527,N_2597);
or U3125 (N_3125,N_2669,N_2590);
nor U3126 (N_3126,N_2872,N_2547);
nand U3127 (N_3127,N_2303,N_2871);
nand U3128 (N_3128,N_2776,N_2963);
nor U3129 (N_3129,N_2514,N_2598);
and U3130 (N_3130,N_2983,N_2419);
or U3131 (N_3131,N_2705,N_2509);
and U3132 (N_3132,N_2305,N_2254);
and U3133 (N_3133,N_2608,N_2615);
or U3134 (N_3134,N_2889,N_2280);
xor U3135 (N_3135,N_2893,N_2744);
nor U3136 (N_3136,N_2294,N_2787);
or U3137 (N_3137,N_2253,N_2745);
xnor U3138 (N_3138,N_2421,N_2824);
nor U3139 (N_3139,N_2934,N_2675);
or U3140 (N_3140,N_2317,N_2999);
nor U3141 (N_3141,N_2606,N_2962);
or U3142 (N_3142,N_2427,N_2343);
or U3143 (N_3143,N_2483,N_2304);
and U3144 (N_3144,N_2922,N_2442);
xor U3145 (N_3145,N_2469,N_2627);
nor U3146 (N_3146,N_2491,N_2969);
xnor U3147 (N_3147,N_2666,N_2903);
nor U3148 (N_3148,N_2985,N_2972);
or U3149 (N_3149,N_2439,N_2472);
nand U3150 (N_3150,N_2835,N_2475);
nand U3151 (N_3151,N_2261,N_2523);
xnor U3152 (N_3152,N_2554,N_2690);
and U3153 (N_3153,N_2878,N_2273);
nand U3154 (N_3154,N_2394,N_2930);
or U3155 (N_3155,N_2532,N_2741);
or U3156 (N_3156,N_2381,N_2284);
or U3157 (N_3157,N_2989,N_2755);
or U3158 (N_3158,N_2290,N_2699);
nor U3159 (N_3159,N_2479,N_2897);
or U3160 (N_3160,N_2376,N_2593);
or U3161 (N_3161,N_2619,N_2287);
xor U3162 (N_3162,N_2804,N_2943);
or U3163 (N_3163,N_2834,N_2543);
and U3164 (N_3164,N_2344,N_2454);
and U3165 (N_3165,N_2762,N_2687);
or U3166 (N_3166,N_2299,N_2334);
or U3167 (N_3167,N_2734,N_2561);
or U3168 (N_3168,N_2829,N_2335);
nor U3169 (N_3169,N_2917,N_2946);
nor U3170 (N_3170,N_2671,N_2632);
xor U3171 (N_3171,N_2345,N_2339);
and U3172 (N_3172,N_2377,N_2718);
nor U3173 (N_3173,N_2417,N_2407);
nor U3174 (N_3174,N_2493,N_2704);
xor U3175 (N_3175,N_2866,N_2297);
nor U3176 (N_3176,N_2412,N_2416);
and U3177 (N_3177,N_2364,N_2692);
xnor U3178 (N_3178,N_2580,N_2559);
xnor U3179 (N_3179,N_2501,N_2560);
or U3180 (N_3180,N_2293,N_2617);
nand U3181 (N_3181,N_2519,N_2956);
nor U3182 (N_3182,N_2260,N_2912);
and U3183 (N_3183,N_2395,N_2518);
xor U3184 (N_3184,N_2570,N_2616);
nand U3185 (N_3185,N_2833,N_2567);
nor U3186 (N_3186,N_2426,N_2974);
or U3187 (N_3187,N_2391,N_2463);
and U3188 (N_3188,N_2595,N_2587);
nand U3189 (N_3189,N_2907,N_2680);
or U3190 (N_3190,N_2630,N_2330);
and U3191 (N_3191,N_2276,N_2980);
or U3192 (N_3192,N_2275,N_2288);
and U3193 (N_3193,N_2654,N_2422);
and U3194 (N_3194,N_2896,N_2286);
xor U3195 (N_3195,N_2975,N_2406);
nand U3196 (N_3196,N_2788,N_2933);
xnor U3197 (N_3197,N_2592,N_2482);
and U3198 (N_3198,N_2314,N_2384);
nand U3199 (N_3199,N_2846,N_2459);
nor U3200 (N_3200,N_2938,N_2611);
nand U3201 (N_3201,N_2329,N_2388);
or U3202 (N_3202,N_2424,N_2362);
nor U3203 (N_3203,N_2534,N_2440);
and U3204 (N_3204,N_2496,N_2774);
xor U3205 (N_3205,N_2697,N_2451);
or U3206 (N_3206,N_2289,N_2499);
nand U3207 (N_3207,N_2301,N_2961);
xnor U3208 (N_3208,N_2651,N_2328);
nand U3209 (N_3209,N_2316,N_2996);
nor U3210 (N_3210,N_2526,N_2686);
or U3211 (N_3211,N_2710,N_2333);
and U3212 (N_3212,N_2902,N_2931);
or U3213 (N_3213,N_2694,N_2548);
and U3214 (N_3214,N_2640,N_2256);
and U3215 (N_3215,N_2637,N_2462);
xnor U3216 (N_3216,N_2612,N_2660);
xnor U3217 (N_3217,N_2533,N_2635);
or U3218 (N_3218,N_2557,N_2750);
nand U3219 (N_3219,N_2891,N_2913);
nand U3220 (N_3220,N_2914,N_2850);
xnor U3221 (N_3221,N_2859,N_2925);
nand U3222 (N_3222,N_2770,N_2778);
and U3223 (N_3223,N_2450,N_2798);
and U3224 (N_3224,N_2822,N_2556);
nand U3225 (N_3225,N_2429,N_2729);
nor U3226 (N_3226,N_2781,N_2782);
xnor U3227 (N_3227,N_2452,N_2719);
and U3228 (N_3228,N_2748,N_2468);
and U3229 (N_3229,N_2645,N_2506);
or U3230 (N_3230,N_2573,N_2677);
and U3231 (N_3231,N_2358,N_2665);
nor U3232 (N_3232,N_2851,N_2311);
and U3233 (N_3233,N_2433,N_2313);
and U3234 (N_3234,N_2772,N_2994);
and U3235 (N_3235,N_2880,N_2411);
nor U3236 (N_3236,N_2498,N_2470);
nand U3237 (N_3237,N_2904,N_2420);
nor U3238 (N_3238,N_2565,N_2838);
xnor U3239 (N_3239,N_2495,N_2323);
nor U3240 (N_3240,N_2709,N_2535);
or U3241 (N_3241,N_2935,N_2629);
or U3242 (N_3242,N_2873,N_2831);
nand U3243 (N_3243,N_2870,N_2257);
xor U3244 (N_3244,N_2269,N_2731);
xor U3245 (N_3245,N_2579,N_2308);
and U3246 (N_3246,N_2594,N_2898);
or U3247 (N_3247,N_2326,N_2390);
xnor U3248 (N_3248,N_2385,N_2614);
or U3249 (N_3249,N_2921,N_2797);
nor U3250 (N_3250,N_2408,N_2845);
nor U3251 (N_3251,N_2724,N_2631);
and U3252 (N_3252,N_2368,N_2950);
nor U3253 (N_3253,N_2435,N_2545);
nor U3254 (N_3254,N_2610,N_2585);
xor U3255 (N_3255,N_2924,N_2720);
nand U3256 (N_3256,N_2853,N_2550);
nand U3257 (N_3257,N_2661,N_2796);
xnor U3258 (N_3258,N_2863,N_2375);
xnor U3259 (N_3259,N_2642,N_2678);
xnor U3260 (N_3260,N_2386,N_2701);
nand U3261 (N_3261,N_2937,N_2715);
and U3262 (N_3262,N_2332,N_2602);
nand U3263 (N_3263,N_2653,N_2728);
or U3264 (N_3264,N_2830,N_2327);
nand U3265 (N_3265,N_2681,N_2357);
xor U3266 (N_3266,N_2737,N_2477);
xor U3267 (N_3267,N_2418,N_2378);
xnor U3268 (N_3268,N_2881,N_2730);
nand U3269 (N_3269,N_2636,N_2840);
xor U3270 (N_3270,N_2876,N_2751);
nor U3271 (N_3271,N_2900,N_2578);
and U3272 (N_3272,N_2779,N_2315);
nand U3273 (N_3273,N_2806,N_2861);
nand U3274 (N_3274,N_2574,N_2576);
nand U3275 (N_3275,N_2497,N_2402);
or U3276 (N_3276,N_2609,N_2599);
nand U3277 (N_3277,N_2683,N_2624);
xnor U3278 (N_3278,N_2777,N_2353);
or U3279 (N_3279,N_2841,N_2966);
and U3280 (N_3280,N_2805,N_2350);
nand U3281 (N_3281,N_2268,N_2562);
nor U3282 (N_3282,N_2811,N_2868);
nor U3283 (N_3283,N_2508,N_2371);
or U3284 (N_3284,N_2929,N_2414);
nand U3285 (N_3285,N_2899,N_2515);
and U3286 (N_3286,N_2461,N_2583);
nand U3287 (N_3287,N_2939,N_2466);
and U3288 (N_3288,N_2918,N_2500);
nor U3289 (N_3289,N_2927,N_2906);
nand U3290 (N_3290,N_2664,N_2628);
and U3291 (N_3291,N_2425,N_2310);
or U3292 (N_3292,N_2970,N_2405);
nand U3293 (N_3293,N_2355,N_2349);
and U3294 (N_3294,N_2476,N_2836);
or U3295 (N_3295,N_2673,N_2342);
and U3296 (N_3296,N_2298,N_2369);
xnor U3297 (N_3297,N_2292,N_2847);
nand U3298 (N_3298,N_2944,N_2502);
or U3299 (N_3299,N_2505,N_2910);
and U3300 (N_3300,N_2513,N_2735);
or U3301 (N_3301,N_2605,N_2264);
nor U3302 (N_3302,N_2460,N_2821);
nor U3303 (N_3303,N_2951,N_2768);
nand U3304 (N_3304,N_2948,N_2625);
xnor U3305 (N_3305,N_2430,N_2874);
nand U3306 (N_3306,N_2714,N_2864);
nand U3307 (N_3307,N_2747,N_2732);
and U3308 (N_3308,N_2621,N_2474);
nor U3309 (N_3309,N_2765,N_2764);
nand U3310 (N_3310,N_2852,N_2633);
or U3311 (N_3311,N_2799,N_2911);
and U3312 (N_3312,N_2525,N_2626);
nor U3313 (N_3313,N_2977,N_2544);
nor U3314 (N_3314,N_2322,N_2947);
and U3315 (N_3315,N_2409,N_2738);
nor U3316 (N_3316,N_2403,N_2443);
or U3317 (N_3317,N_2887,N_2584);
xnor U3318 (N_3318,N_2618,N_2644);
nand U3319 (N_3319,N_2486,N_2767);
xnor U3320 (N_3320,N_2641,N_2684);
nand U3321 (N_3321,N_2531,N_2549);
nand U3322 (N_3322,N_2320,N_2281);
and U3323 (N_3323,N_2604,N_2722);
nand U3324 (N_3324,N_2987,N_2365);
or U3325 (N_3325,N_2886,N_2648);
and U3326 (N_3326,N_2302,N_2436);
nor U3327 (N_3327,N_2448,N_2668);
nand U3328 (N_3328,N_2992,N_2274);
or U3329 (N_3329,N_2984,N_2445);
and U3330 (N_3330,N_2542,N_2986);
or U3331 (N_3331,N_2743,N_2649);
xnor U3332 (N_3332,N_2473,N_2818);
or U3333 (N_3333,N_2832,N_2971);
xor U3334 (N_3334,N_2291,N_2752);
nor U3335 (N_3335,N_2647,N_2958);
or U3336 (N_3336,N_2757,N_2577);
nand U3337 (N_3337,N_2809,N_2646);
nand U3338 (N_3338,N_2674,N_2689);
xnor U3339 (N_3339,N_2775,N_2800);
nor U3340 (N_3340,N_2359,N_2620);
and U3341 (N_3341,N_2652,N_2552);
nor U3342 (N_3342,N_2696,N_2613);
nand U3343 (N_3343,N_2708,N_2607);
nand U3344 (N_3344,N_2828,N_2936);
nor U3345 (N_3345,N_2968,N_2588);
and U3346 (N_3346,N_2790,N_2763);
nor U3347 (N_3347,N_2285,N_2340);
nand U3348 (N_3348,N_2670,N_2348);
and U3349 (N_3349,N_2447,N_2698);
nand U3350 (N_3350,N_2952,N_2826);
nand U3351 (N_3351,N_2361,N_2392);
and U3352 (N_3352,N_2693,N_2596);
xnor U3353 (N_3353,N_2300,N_2717);
xnor U3354 (N_3354,N_2814,N_2813);
and U3355 (N_3355,N_2346,N_2786);
or U3356 (N_3356,N_2794,N_2761);
nor U3357 (N_3357,N_2756,N_2568);
xor U3358 (N_3358,N_2659,N_2441);
nand U3359 (N_3359,N_2857,N_2808);
or U3360 (N_3360,N_2815,N_2827);
nor U3361 (N_3361,N_2916,N_2638);
xnor U3362 (N_3362,N_2842,N_2789);
or U3363 (N_3363,N_2331,N_2885);
nor U3364 (N_3364,N_2766,N_2603);
or U3365 (N_3365,N_2488,N_2848);
or U3366 (N_3366,N_2263,N_2688);
and U3367 (N_3367,N_2792,N_2860);
nor U3368 (N_3368,N_2919,N_2338);
or U3369 (N_3369,N_2538,N_2555);
and U3370 (N_3370,N_2400,N_2807);
nor U3371 (N_3371,N_2875,N_2295);
nand U3372 (N_3372,N_2926,N_2251);
and U3373 (N_3373,N_2279,N_2494);
and U3374 (N_3374,N_2667,N_2739);
xnor U3375 (N_3375,N_2908,N_2474);
nor U3376 (N_3376,N_2950,N_2885);
and U3377 (N_3377,N_2816,N_2478);
nor U3378 (N_3378,N_2605,N_2646);
xor U3379 (N_3379,N_2589,N_2262);
xnor U3380 (N_3380,N_2482,N_2896);
nor U3381 (N_3381,N_2560,N_2336);
and U3382 (N_3382,N_2582,N_2874);
and U3383 (N_3383,N_2909,N_2958);
nor U3384 (N_3384,N_2330,N_2876);
and U3385 (N_3385,N_2422,N_2667);
nor U3386 (N_3386,N_2837,N_2884);
nor U3387 (N_3387,N_2343,N_2402);
and U3388 (N_3388,N_2310,N_2470);
nor U3389 (N_3389,N_2906,N_2984);
or U3390 (N_3390,N_2688,N_2646);
or U3391 (N_3391,N_2950,N_2578);
or U3392 (N_3392,N_2306,N_2453);
xnor U3393 (N_3393,N_2659,N_2969);
nor U3394 (N_3394,N_2532,N_2261);
nand U3395 (N_3395,N_2922,N_2380);
nand U3396 (N_3396,N_2422,N_2912);
xnor U3397 (N_3397,N_2424,N_2974);
and U3398 (N_3398,N_2785,N_2358);
xnor U3399 (N_3399,N_2992,N_2426);
xnor U3400 (N_3400,N_2251,N_2908);
and U3401 (N_3401,N_2671,N_2910);
xor U3402 (N_3402,N_2251,N_2353);
nor U3403 (N_3403,N_2716,N_2310);
nand U3404 (N_3404,N_2457,N_2906);
nand U3405 (N_3405,N_2778,N_2437);
nand U3406 (N_3406,N_2840,N_2622);
xnor U3407 (N_3407,N_2911,N_2832);
or U3408 (N_3408,N_2978,N_2330);
and U3409 (N_3409,N_2817,N_2861);
nand U3410 (N_3410,N_2450,N_2456);
nand U3411 (N_3411,N_2723,N_2949);
nand U3412 (N_3412,N_2748,N_2689);
or U3413 (N_3413,N_2562,N_2690);
nand U3414 (N_3414,N_2844,N_2546);
nand U3415 (N_3415,N_2754,N_2939);
and U3416 (N_3416,N_2314,N_2621);
and U3417 (N_3417,N_2508,N_2740);
nor U3418 (N_3418,N_2886,N_2650);
nand U3419 (N_3419,N_2802,N_2363);
xnor U3420 (N_3420,N_2615,N_2308);
nor U3421 (N_3421,N_2429,N_2889);
nor U3422 (N_3422,N_2615,N_2911);
or U3423 (N_3423,N_2717,N_2543);
nor U3424 (N_3424,N_2438,N_2330);
nand U3425 (N_3425,N_2567,N_2922);
and U3426 (N_3426,N_2464,N_2313);
and U3427 (N_3427,N_2893,N_2658);
and U3428 (N_3428,N_2646,N_2524);
or U3429 (N_3429,N_2280,N_2432);
nor U3430 (N_3430,N_2893,N_2680);
nor U3431 (N_3431,N_2810,N_2278);
or U3432 (N_3432,N_2661,N_2603);
or U3433 (N_3433,N_2862,N_2726);
or U3434 (N_3434,N_2349,N_2268);
xnor U3435 (N_3435,N_2574,N_2992);
xor U3436 (N_3436,N_2914,N_2544);
xnor U3437 (N_3437,N_2274,N_2881);
nand U3438 (N_3438,N_2824,N_2521);
nor U3439 (N_3439,N_2272,N_2842);
nand U3440 (N_3440,N_2296,N_2684);
nand U3441 (N_3441,N_2690,N_2755);
or U3442 (N_3442,N_2538,N_2307);
nand U3443 (N_3443,N_2600,N_2275);
xor U3444 (N_3444,N_2340,N_2514);
nor U3445 (N_3445,N_2965,N_2379);
nor U3446 (N_3446,N_2314,N_2397);
nor U3447 (N_3447,N_2954,N_2870);
xnor U3448 (N_3448,N_2447,N_2565);
nor U3449 (N_3449,N_2456,N_2517);
nand U3450 (N_3450,N_2445,N_2535);
nand U3451 (N_3451,N_2899,N_2272);
nor U3452 (N_3452,N_2994,N_2633);
and U3453 (N_3453,N_2728,N_2842);
xnor U3454 (N_3454,N_2592,N_2624);
nor U3455 (N_3455,N_2414,N_2659);
nand U3456 (N_3456,N_2706,N_2838);
xnor U3457 (N_3457,N_2551,N_2717);
and U3458 (N_3458,N_2606,N_2681);
nand U3459 (N_3459,N_2604,N_2743);
nor U3460 (N_3460,N_2932,N_2620);
or U3461 (N_3461,N_2914,N_2829);
and U3462 (N_3462,N_2389,N_2551);
or U3463 (N_3463,N_2584,N_2617);
nand U3464 (N_3464,N_2844,N_2386);
xor U3465 (N_3465,N_2946,N_2810);
and U3466 (N_3466,N_2865,N_2800);
nand U3467 (N_3467,N_2286,N_2897);
or U3468 (N_3468,N_2403,N_2374);
or U3469 (N_3469,N_2488,N_2520);
nor U3470 (N_3470,N_2827,N_2718);
and U3471 (N_3471,N_2399,N_2559);
nor U3472 (N_3472,N_2483,N_2840);
or U3473 (N_3473,N_2547,N_2949);
xor U3474 (N_3474,N_2530,N_2526);
nand U3475 (N_3475,N_2342,N_2850);
nor U3476 (N_3476,N_2752,N_2676);
nor U3477 (N_3477,N_2262,N_2393);
and U3478 (N_3478,N_2518,N_2574);
or U3479 (N_3479,N_2885,N_2639);
or U3480 (N_3480,N_2772,N_2860);
xor U3481 (N_3481,N_2690,N_2858);
and U3482 (N_3482,N_2869,N_2391);
and U3483 (N_3483,N_2318,N_2420);
or U3484 (N_3484,N_2481,N_2657);
and U3485 (N_3485,N_2404,N_2678);
and U3486 (N_3486,N_2890,N_2568);
or U3487 (N_3487,N_2952,N_2964);
xnor U3488 (N_3488,N_2629,N_2726);
nor U3489 (N_3489,N_2455,N_2666);
nor U3490 (N_3490,N_2836,N_2634);
or U3491 (N_3491,N_2288,N_2903);
or U3492 (N_3492,N_2623,N_2984);
and U3493 (N_3493,N_2621,N_2920);
and U3494 (N_3494,N_2259,N_2436);
nor U3495 (N_3495,N_2501,N_2929);
or U3496 (N_3496,N_2895,N_2615);
xor U3497 (N_3497,N_2401,N_2308);
and U3498 (N_3498,N_2282,N_2373);
nand U3499 (N_3499,N_2808,N_2329);
or U3500 (N_3500,N_2957,N_2424);
or U3501 (N_3501,N_2541,N_2379);
or U3502 (N_3502,N_2451,N_2867);
xnor U3503 (N_3503,N_2265,N_2995);
nand U3504 (N_3504,N_2460,N_2842);
and U3505 (N_3505,N_2624,N_2897);
and U3506 (N_3506,N_2259,N_2669);
nor U3507 (N_3507,N_2897,N_2539);
and U3508 (N_3508,N_2785,N_2963);
and U3509 (N_3509,N_2261,N_2495);
and U3510 (N_3510,N_2538,N_2562);
xnor U3511 (N_3511,N_2780,N_2423);
and U3512 (N_3512,N_2327,N_2530);
and U3513 (N_3513,N_2350,N_2645);
nor U3514 (N_3514,N_2722,N_2297);
or U3515 (N_3515,N_2401,N_2472);
or U3516 (N_3516,N_2707,N_2271);
and U3517 (N_3517,N_2627,N_2454);
nand U3518 (N_3518,N_2538,N_2999);
nor U3519 (N_3519,N_2356,N_2381);
or U3520 (N_3520,N_2518,N_2431);
nor U3521 (N_3521,N_2564,N_2378);
and U3522 (N_3522,N_2954,N_2953);
nor U3523 (N_3523,N_2677,N_2482);
and U3524 (N_3524,N_2784,N_2790);
and U3525 (N_3525,N_2517,N_2682);
xnor U3526 (N_3526,N_2886,N_2713);
or U3527 (N_3527,N_2872,N_2551);
xnor U3528 (N_3528,N_2704,N_2310);
or U3529 (N_3529,N_2471,N_2561);
nor U3530 (N_3530,N_2290,N_2545);
nor U3531 (N_3531,N_2607,N_2804);
nor U3532 (N_3532,N_2311,N_2679);
nand U3533 (N_3533,N_2293,N_2678);
xor U3534 (N_3534,N_2640,N_2734);
nand U3535 (N_3535,N_2554,N_2337);
nand U3536 (N_3536,N_2588,N_2786);
nor U3537 (N_3537,N_2709,N_2754);
xor U3538 (N_3538,N_2420,N_2667);
and U3539 (N_3539,N_2908,N_2699);
or U3540 (N_3540,N_2352,N_2401);
xor U3541 (N_3541,N_2484,N_2520);
nor U3542 (N_3542,N_2956,N_2891);
and U3543 (N_3543,N_2758,N_2900);
and U3544 (N_3544,N_2989,N_2507);
and U3545 (N_3545,N_2458,N_2538);
nand U3546 (N_3546,N_2406,N_2927);
nand U3547 (N_3547,N_2677,N_2598);
nand U3548 (N_3548,N_2432,N_2892);
nor U3549 (N_3549,N_2341,N_2623);
or U3550 (N_3550,N_2382,N_2713);
or U3551 (N_3551,N_2868,N_2388);
xnor U3552 (N_3552,N_2384,N_2379);
nor U3553 (N_3553,N_2954,N_2261);
xor U3554 (N_3554,N_2512,N_2376);
nand U3555 (N_3555,N_2853,N_2844);
or U3556 (N_3556,N_2283,N_2707);
nand U3557 (N_3557,N_2469,N_2455);
nand U3558 (N_3558,N_2696,N_2965);
nand U3559 (N_3559,N_2304,N_2370);
and U3560 (N_3560,N_2426,N_2479);
nor U3561 (N_3561,N_2330,N_2975);
xnor U3562 (N_3562,N_2695,N_2301);
nor U3563 (N_3563,N_2414,N_2405);
or U3564 (N_3564,N_2663,N_2689);
or U3565 (N_3565,N_2285,N_2934);
and U3566 (N_3566,N_2905,N_2591);
and U3567 (N_3567,N_2959,N_2924);
and U3568 (N_3568,N_2274,N_2848);
nand U3569 (N_3569,N_2955,N_2468);
or U3570 (N_3570,N_2634,N_2447);
xor U3571 (N_3571,N_2445,N_2873);
nor U3572 (N_3572,N_2583,N_2610);
xnor U3573 (N_3573,N_2856,N_2943);
nor U3574 (N_3574,N_2380,N_2894);
and U3575 (N_3575,N_2779,N_2924);
nor U3576 (N_3576,N_2498,N_2963);
or U3577 (N_3577,N_2466,N_2722);
and U3578 (N_3578,N_2961,N_2923);
and U3579 (N_3579,N_2456,N_2426);
or U3580 (N_3580,N_2963,N_2401);
xnor U3581 (N_3581,N_2622,N_2645);
nand U3582 (N_3582,N_2494,N_2524);
nor U3583 (N_3583,N_2747,N_2964);
nor U3584 (N_3584,N_2993,N_2354);
xnor U3585 (N_3585,N_2534,N_2263);
xnor U3586 (N_3586,N_2291,N_2971);
or U3587 (N_3587,N_2741,N_2941);
xor U3588 (N_3588,N_2635,N_2320);
xor U3589 (N_3589,N_2614,N_2559);
or U3590 (N_3590,N_2610,N_2619);
nand U3591 (N_3591,N_2776,N_2636);
or U3592 (N_3592,N_2563,N_2301);
nor U3593 (N_3593,N_2953,N_2538);
nand U3594 (N_3594,N_2583,N_2941);
nor U3595 (N_3595,N_2863,N_2653);
or U3596 (N_3596,N_2841,N_2322);
and U3597 (N_3597,N_2421,N_2990);
nor U3598 (N_3598,N_2961,N_2295);
and U3599 (N_3599,N_2784,N_2761);
xor U3600 (N_3600,N_2975,N_2543);
or U3601 (N_3601,N_2469,N_2890);
or U3602 (N_3602,N_2331,N_2509);
or U3603 (N_3603,N_2713,N_2806);
nor U3604 (N_3604,N_2971,N_2967);
xnor U3605 (N_3605,N_2531,N_2545);
nor U3606 (N_3606,N_2628,N_2700);
or U3607 (N_3607,N_2421,N_2777);
xor U3608 (N_3608,N_2989,N_2667);
and U3609 (N_3609,N_2990,N_2368);
and U3610 (N_3610,N_2316,N_2509);
nor U3611 (N_3611,N_2931,N_2818);
or U3612 (N_3612,N_2879,N_2323);
nor U3613 (N_3613,N_2879,N_2702);
or U3614 (N_3614,N_2557,N_2522);
nor U3615 (N_3615,N_2452,N_2435);
or U3616 (N_3616,N_2743,N_2315);
or U3617 (N_3617,N_2274,N_2730);
xnor U3618 (N_3618,N_2950,N_2341);
nor U3619 (N_3619,N_2343,N_2714);
or U3620 (N_3620,N_2460,N_2671);
nor U3621 (N_3621,N_2656,N_2914);
nor U3622 (N_3622,N_2396,N_2280);
xnor U3623 (N_3623,N_2360,N_2434);
or U3624 (N_3624,N_2883,N_2542);
and U3625 (N_3625,N_2538,N_2398);
xnor U3626 (N_3626,N_2475,N_2862);
nor U3627 (N_3627,N_2501,N_2747);
nor U3628 (N_3628,N_2679,N_2680);
nor U3629 (N_3629,N_2433,N_2829);
xnor U3630 (N_3630,N_2314,N_2948);
or U3631 (N_3631,N_2490,N_2401);
and U3632 (N_3632,N_2648,N_2733);
or U3633 (N_3633,N_2836,N_2616);
and U3634 (N_3634,N_2383,N_2287);
xnor U3635 (N_3635,N_2497,N_2769);
nor U3636 (N_3636,N_2664,N_2393);
nor U3637 (N_3637,N_2409,N_2699);
nand U3638 (N_3638,N_2332,N_2280);
or U3639 (N_3639,N_2284,N_2398);
and U3640 (N_3640,N_2294,N_2279);
xor U3641 (N_3641,N_2500,N_2584);
nand U3642 (N_3642,N_2644,N_2468);
nand U3643 (N_3643,N_2987,N_2834);
and U3644 (N_3644,N_2914,N_2314);
and U3645 (N_3645,N_2313,N_2396);
xor U3646 (N_3646,N_2904,N_2874);
nor U3647 (N_3647,N_2534,N_2881);
nand U3648 (N_3648,N_2386,N_2804);
xor U3649 (N_3649,N_2375,N_2775);
nand U3650 (N_3650,N_2809,N_2705);
or U3651 (N_3651,N_2310,N_2777);
xnor U3652 (N_3652,N_2993,N_2760);
xor U3653 (N_3653,N_2556,N_2475);
nor U3654 (N_3654,N_2866,N_2499);
and U3655 (N_3655,N_2689,N_2380);
xor U3656 (N_3656,N_2317,N_2486);
or U3657 (N_3657,N_2918,N_2267);
and U3658 (N_3658,N_2665,N_2987);
and U3659 (N_3659,N_2903,N_2590);
nor U3660 (N_3660,N_2921,N_2591);
and U3661 (N_3661,N_2297,N_2792);
nor U3662 (N_3662,N_2357,N_2330);
or U3663 (N_3663,N_2717,N_2351);
xor U3664 (N_3664,N_2455,N_2860);
xor U3665 (N_3665,N_2820,N_2254);
nor U3666 (N_3666,N_2403,N_2468);
and U3667 (N_3667,N_2747,N_2560);
and U3668 (N_3668,N_2615,N_2485);
or U3669 (N_3669,N_2274,N_2325);
nor U3670 (N_3670,N_2813,N_2889);
xor U3671 (N_3671,N_2713,N_2590);
or U3672 (N_3672,N_2924,N_2595);
nand U3673 (N_3673,N_2287,N_2995);
nand U3674 (N_3674,N_2586,N_2864);
and U3675 (N_3675,N_2888,N_2920);
nand U3676 (N_3676,N_2991,N_2732);
nor U3677 (N_3677,N_2943,N_2526);
or U3678 (N_3678,N_2806,N_2955);
or U3679 (N_3679,N_2810,N_2274);
and U3680 (N_3680,N_2720,N_2714);
nand U3681 (N_3681,N_2267,N_2647);
xnor U3682 (N_3682,N_2737,N_2910);
and U3683 (N_3683,N_2959,N_2324);
xnor U3684 (N_3684,N_2775,N_2665);
and U3685 (N_3685,N_2924,N_2668);
and U3686 (N_3686,N_2406,N_2492);
nor U3687 (N_3687,N_2392,N_2944);
and U3688 (N_3688,N_2845,N_2594);
or U3689 (N_3689,N_2459,N_2422);
nor U3690 (N_3690,N_2991,N_2874);
nand U3691 (N_3691,N_2503,N_2635);
xnor U3692 (N_3692,N_2867,N_2803);
nor U3693 (N_3693,N_2411,N_2672);
nand U3694 (N_3694,N_2694,N_2262);
or U3695 (N_3695,N_2401,N_2619);
or U3696 (N_3696,N_2732,N_2424);
xnor U3697 (N_3697,N_2940,N_2992);
or U3698 (N_3698,N_2303,N_2607);
or U3699 (N_3699,N_2932,N_2319);
nand U3700 (N_3700,N_2339,N_2741);
or U3701 (N_3701,N_2677,N_2445);
or U3702 (N_3702,N_2393,N_2996);
and U3703 (N_3703,N_2430,N_2533);
xnor U3704 (N_3704,N_2894,N_2832);
or U3705 (N_3705,N_2565,N_2294);
or U3706 (N_3706,N_2894,N_2273);
nor U3707 (N_3707,N_2748,N_2709);
nand U3708 (N_3708,N_2730,N_2705);
and U3709 (N_3709,N_2459,N_2797);
or U3710 (N_3710,N_2502,N_2797);
nor U3711 (N_3711,N_2436,N_2458);
and U3712 (N_3712,N_2379,N_2552);
or U3713 (N_3713,N_2408,N_2290);
nand U3714 (N_3714,N_2995,N_2510);
xor U3715 (N_3715,N_2560,N_2603);
nor U3716 (N_3716,N_2376,N_2397);
or U3717 (N_3717,N_2823,N_2854);
nand U3718 (N_3718,N_2958,N_2660);
or U3719 (N_3719,N_2772,N_2819);
or U3720 (N_3720,N_2566,N_2716);
or U3721 (N_3721,N_2433,N_2547);
and U3722 (N_3722,N_2332,N_2895);
and U3723 (N_3723,N_2794,N_2618);
nand U3724 (N_3724,N_2797,N_2619);
nor U3725 (N_3725,N_2977,N_2949);
nand U3726 (N_3726,N_2583,N_2483);
nor U3727 (N_3727,N_2353,N_2792);
or U3728 (N_3728,N_2715,N_2975);
nand U3729 (N_3729,N_2399,N_2891);
or U3730 (N_3730,N_2618,N_2927);
xor U3731 (N_3731,N_2526,N_2772);
nand U3732 (N_3732,N_2751,N_2834);
or U3733 (N_3733,N_2840,N_2545);
nor U3734 (N_3734,N_2455,N_2496);
or U3735 (N_3735,N_2504,N_2682);
or U3736 (N_3736,N_2699,N_2695);
nor U3737 (N_3737,N_2571,N_2755);
and U3738 (N_3738,N_2568,N_2969);
nand U3739 (N_3739,N_2775,N_2653);
nand U3740 (N_3740,N_2713,N_2982);
or U3741 (N_3741,N_2573,N_2623);
and U3742 (N_3742,N_2373,N_2903);
xor U3743 (N_3743,N_2532,N_2698);
or U3744 (N_3744,N_2386,N_2715);
nor U3745 (N_3745,N_2974,N_2382);
nand U3746 (N_3746,N_2426,N_2418);
nor U3747 (N_3747,N_2814,N_2312);
xor U3748 (N_3748,N_2432,N_2603);
xor U3749 (N_3749,N_2844,N_2515);
xnor U3750 (N_3750,N_3206,N_3497);
nand U3751 (N_3751,N_3371,N_3722);
and U3752 (N_3752,N_3131,N_3681);
or U3753 (N_3753,N_3664,N_3199);
nand U3754 (N_3754,N_3038,N_3093);
and U3755 (N_3755,N_3384,N_3082);
or U3756 (N_3756,N_3215,N_3053);
nand U3757 (N_3757,N_3685,N_3579);
and U3758 (N_3758,N_3250,N_3203);
or U3759 (N_3759,N_3401,N_3555);
or U3760 (N_3760,N_3455,N_3020);
nor U3761 (N_3761,N_3421,N_3018);
nand U3762 (N_3762,N_3631,N_3533);
nand U3763 (N_3763,N_3575,N_3657);
nand U3764 (N_3764,N_3314,N_3336);
or U3765 (N_3765,N_3247,N_3243);
nand U3766 (N_3766,N_3283,N_3282);
and U3767 (N_3767,N_3504,N_3196);
nor U3768 (N_3768,N_3150,N_3456);
xnor U3769 (N_3769,N_3597,N_3677);
xnor U3770 (N_3770,N_3094,N_3168);
xnor U3771 (N_3771,N_3568,N_3034);
and U3772 (N_3772,N_3558,N_3029);
or U3773 (N_3773,N_3182,N_3599);
nor U3774 (N_3774,N_3682,N_3185);
xor U3775 (N_3775,N_3554,N_3274);
nor U3776 (N_3776,N_3586,N_3704);
nor U3777 (N_3777,N_3736,N_3201);
xnor U3778 (N_3778,N_3382,N_3633);
nand U3779 (N_3779,N_3543,N_3662);
and U3780 (N_3780,N_3214,N_3403);
or U3781 (N_3781,N_3112,N_3672);
nor U3782 (N_3782,N_3589,N_3535);
xnor U3783 (N_3783,N_3080,N_3102);
nor U3784 (N_3784,N_3576,N_3103);
nor U3785 (N_3785,N_3278,N_3075);
xor U3786 (N_3786,N_3588,N_3227);
or U3787 (N_3787,N_3390,N_3095);
and U3788 (N_3788,N_3607,N_3132);
xor U3789 (N_3789,N_3123,N_3129);
and U3790 (N_3790,N_3530,N_3621);
nand U3791 (N_3791,N_3559,N_3479);
and U3792 (N_3792,N_3210,N_3313);
nor U3793 (N_3793,N_3581,N_3602);
nor U3794 (N_3794,N_3548,N_3748);
and U3795 (N_3795,N_3295,N_3276);
and U3796 (N_3796,N_3078,N_3051);
nand U3797 (N_3797,N_3083,N_3057);
nand U3798 (N_3798,N_3126,N_3560);
nand U3799 (N_3799,N_3244,N_3228);
nor U3800 (N_3800,N_3337,N_3236);
or U3801 (N_3801,N_3515,N_3204);
xor U3802 (N_3802,N_3149,N_3041);
nand U3803 (N_3803,N_3605,N_3121);
xor U3804 (N_3804,N_3398,N_3361);
nor U3805 (N_3805,N_3011,N_3137);
nor U3806 (N_3806,N_3623,N_3175);
and U3807 (N_3807,N_3578,N_3342);
or U3808 (N_3808,N_3715,N_3143);
xnor U3809 (N_3809,N_3574,N_3180);
nand U3810 (N_3810,N_3408,N_3417);
xnor U3811 (N_3811,N_3307,N_3510);
and U3812 (N_3812,N_3135,N_3644);
nand U3813 (N_3813,N_3404,N_3161);
or U3814 (N_3814,N_3419,N_3154);
or U3815 (N_3815,N_3289,N_3267);
and U3816 (N_3816,N_3077,N_3364);
nand U3817 (N_3817,N_3489,N_3517);
and U3818 (N_3818,N_3625,N_3117);
and U3819 (N_3819,N_3136,N_3360);
xnor U3820 (N_3820,N_3606,N_3348);
xor U3821 (N_3821,N_3202,N_3380);
and U3822 (N_3822,N_3663,N_3655);
and U3823 (N_3823,N_3690,N_3622);
or U3824 (N_3824,N_3349,N_3618);
xor U3825 (N_3825,N_3749,N_3465);
or U3826 (N_3826,N_3138,N_3067);
nand U3827 (N_3827,N_3509,N_3039);
xnor U3828 (N_3828,N_3650,N_3340);
xnor U3829 (N_3829,N_3587,N_3482);
xor U3830 (N_3830,N_3061,N_3629);
and U3831 (N_3831,N_3259,N_3166);
and U3832 (N_3832,N_3221,N_3661);
xor U3833 (N_3833,N_3414,N_3462);
and U3834 (N_3834,N_3298,N_3415);
or U3835 (N_3835,N_3590,N_3518);
nand U3836 (N_3836,N_3321,N_3411);
nor U3837 (N_3837,N_3301,N_3226);
nor U3838 (N_3838,N_3596,N_3467);
or U3839 (N_3839,N_3127,N_3604);
and U3840 (N_3840,N_3104,N_3015);
nor U3841 (N_3841,N_3213,N_3146);
nand U3842 (N_3842,N_3688,N_3721);
nand U3843 (N_3843,N_3211,N_3252);
nor U3844 (N_3844,N_3447,N_3148);
nor U3845 (N_3845,N_3217,N_3553);
and U3846 (N_3846,N_3372,N_3028);
xnor U3847 (N_3847,N_3643,N_3675);
nand U3848 (N_3848,N_3732,N_3220);
nor U3849 (N_3849,N_3583,N_3229);
and U3850 (N_3850,N_3058,N_3035);
and U3851 (N_3851,N_3043,N_3004);
xor U3852 (N_3852,N_3648,N_3144);
xnor U3853 (N_3853,N_3552,N_3435);
nand U3854 (N_3854,N_3355,N_3641);
nand U3855 (N_3855,N_3725,N_3717);
and U3856 (N_3856,N_3177,N_3413);
or U3857 (N_3857,N_3585,N_3487);
xor U3858 (N_3858,N_3345,N_3294);
or U3859 (N_3859,N_3626,N_3022);
nand U3860 (N_3860,N_3503,N_3007);
or U3861 (N_3861,N_3079,N_3716);
and U3862 (N_3862,N_3176,N_3318);
and U3863 (N_3863,N_3042,N_3676);
nand U3864 (N_3864,N_3446,N_3532);
nand U3865 (N_3865,N_3156,N_3316);
and U3866 (N_3866,N_3021,N_3733);
xnor U3867 (N_3867,N_3331,N_3139);
and U3868 (N_3868,N_3737,N_3678);
and U3869 (N_3869,N_3433,N_3466);
nand U3870 (N_3870,N_3001,N_3153);
nor U3871 (N_3871,N_3550,N_3346);
and U3872 (N_3872,N_3191,N_3065);
or U3873 (N_3873,N_3481,N_3164);
nor U3874 (N_3874,N_3740,N_3549);
nor U3875 (N_3875,N_3375,N_3174);
and U3876 (N_3876,N_3580,N_3335);
nor U3877 (N_3877,N_3428,N_3223);
xnor U3878 (N_3878,N_3113,N_3698);
nor U3879 (N_3879,N_3306,N_3598);
nand U3880 (N_3880,N_3271,N_3438);
and U3881 (N_3881,N_3285,N_3312);
or U3882 (N_3882,N_3024,N_3697);
and U3883 (N_3883,N_3458,N_3656);
nor U3884 (N_3884,N_3570,N_3195);
and U3885 (N_3885,N_3234,N_3556);
and U3886 (N_3886,N_3383,N_3488);
nor U3887 (N_3887,N_3516,N_3388);
xnor U3888 (N_3888,N_3064,N_3734);
and U3889 (N_3889,N_3396,N_3612);
nor U3890 (N_3890,N_3457,N_3299);
nor U3891 (N_3891,N_3665,N_3014);
nand U3892 (N_3892,N_3054,N_3424);
and U3893 (N_3893,N_3531,N_3241);
nor U3894 (N_3894,N_3119,N_3702);
nand U3895 (N_3895,N_3357,N_3448);
nor U3896 (N_3896,N_3513,N_3235);
xnor U3897 (N_3897,N_3128,N_3432);
or U3898 (N_3898,N_3184,N_3072);
nor U3899 (N_3899,N_3052,N_3615);
xor U3900 (N_3900,N_3060,N_3367);
and U3901 (N_3901,N_3744,N_3567);
and U3902 (N_3902,N_3461,N_3670);
or U3903 (N_3903,N_3339,N_3275);
nand U3904 (N_3904,N_3394,N_3356);
nand U3905 (N_3905,N_3699,N_3397);
or U3906 (N_3906,N_3070,N_3671);
nand U3907 (N_3907,N_3037,N_3059);
and U3908 (N_3908,N_3290,N_3085);
or U3909 (N_3909,N_3653,N_3245);
xor U3910 (N_3910,N_3157,N_3608);
nand U3911 (N_3911,N_3141,N_3105);
nor U3912 (N_3912,N_3118,N_3689);
or U3913 (N_3913,N_3536,N_3257);
xor U3914 (N_3914,N_3440,N_3714);
xor U3915 (N_3915,N_3557,N_3476);
xnor U3916 (N_3916,N_3473,N_3529);
nor U3917 (N_3917,N_3495,N_3659);
nand U3918 (N_3918,N_3286,N_3571);
or U3919 (N_3919,N_3296,N_3452);
nor U3920 (N_3920,N_3418,N_3023);
xnor U3921 (N_3921,N_3179,N_3183);
and U3922 (N_3922,N_3212,N_3122);
xnor U3923 (N_3923,N_3524,N_3399);
or U3924 (N_3924,N_3333,N_3280);
nor U3925 (N_3925,N_3522,N_3101);
and U3926 (N_3926,N_3377,N_3044);
and U3927 (N_3927,N_3100,N_3310);
nor U3928 (N_3928,N_3000,N_3572);
nor U3929 (N_3929,N_3158,N_3695);
and U3930 (N_3930,N_3469,N_3266);
nand U3931 (N_3931,N_3025,N_3088);
and U3932 (N_3932,N_3630,N_3406);
and U3933 (N_3933,N_3528,N_3613);
nor U3934 (N_3934,N_3620,N_3674);
nor U3935 (N_3935,N_3254,N_3315);
or U3936 (N_3936,N_3525,N_3405);
nor U3937 (N_3937,N_3638,N_3099);
xnor U3938 (N_3938,N_3288,N_3222);
nand U3939 (N_3939,N_3480,N_3096);
and U3940 (N_3940,N_3645,N_3486);
nand U3941 (N_3941,N_3281,N_3628);
nand U3942 (N_3942,N_3305,N_3500);
nand U3943 (N_3943,N_3352,N_3443);
nand U3944 (N_3944,N_3727,N_3186);
xnor U3945 (N_3945,N_3592,N_3474);
nor U3946 (N_3946,N_3232,N_3219);
nor U3947 (N_3947,N_3603,N_3498);
or U3948 (N_3948,N_3036,N_3068);
nand U3949 (N_3949,N_3169,N_3718);
xnor U3950 (N_3950,N_3673,N_3263);
and U3951 (N_3951,N_3111,N_3430);
nand U3952 (N_3952,N_3649,N_3086);
nand U3953 (N_3953,N_3048,N_3198);
and U3954 (N_3954,N_3279,N_3125);
xor U3955 (N_3955,N_3055,N_3172);
nor U3956 (N_3956,N_3326,N_3651);
nand U3957 (N_3957,N_3292,N_3304);
xnor U3958 (N_3958,N_3499,N_3087);
xor U3959 (N_3959,N_3565,N_3165);
nor U3960 (N_3960,N_3680,N_3062);
xnor U3961 (N_3961,N_3066,N_3287);
xnor U3962 (N_3962,N_3691,N_3505);
nor U3963 (N_3963,N_3492,N_3426);
or U3964 (N_3964,N_3140,N_3109);
xnor U3965 (N_3965,N_3442,N_3047);
nor U3966 (N_3966,N_3658,N_3425);
xnor U3967 (N_3967,N_3713,N_3610);
nand U3968 (N_3968,N_3297,N_3233);
xor U3969 (N_3969,N_3684,N_3441);
and U3970 (N_3970,N_3003,N_3728);
and U3971 (N_3971,N_3193,N_3483);
nand U3972 (N_3972,N_3563,N_3319);
and U3973 (N_3973,N_3601,N_3016);
nor U3974 (N_3974,N_3347,N_3092);
nand U3975 (N_3975,N_3723,N_3694);
and U3976 (N_3976,N_3258,N_3343);
nor U3977 (N_3977,N_3365,N_3485);
nor U3978 (N_3978,N_3617,N_3218);
or U3979 (N_3979,N_3107,N_3017);
or U3980 (N_3980,N_3063,N_3423);
and U3981 (N_3981,N_3667,N_3409);
or U3982 (N_3982,N_3071,N_3260);
nor U3983 (N_3983,N_3152,N_3027);
nand U3984 (N_3984,N_3046,N_3090);
nand U3985 (N_3985,N_3073,N_3130);
and U3986 (N_3986,N_3159,N_3208);
or U3987 (N_3987,N_3050,N_3692);
nand U3988 (N_3988,N_3545,N_3106);
xnor U3989 (N_3989,N_3407,N_3256);
or U3990 (N_3990,N_3323,N_3354);
nor U3991 (N_3991,N_3619,N_3431);
xnor U3992 (N_3992,N_3526,N_3115);
or U3993 (N_3993,N_3049,N_3708);
nor U3994 (N_3994,N_3197,N_3255);
and U3995 (N_3995,N_3300,N_3178);
xor U3996 (N_3996,N_3520,N_3155);
and U3997 (N_3997,N_3593,N_3006);
nor U3998 (N_3998,N_3710,N_3436);
nor U3999 (N_3999,N_3389,N_3262);
and U4000 (N_4000,N_3703,N_3696);
and U4001 (N_4001,N_3668,N_3546);
or U4002 (N_4002,N_3634,N_3540);
nand U4003 (N_4003,N_3216,N_3493);
and U4004 (N_4004,N_3616,N_3181);
nor U4005 (N_4005,N_3705,N_3133);
xor U4006 (N_4006,N_3368,N_3472);
and U4007 (N_4007,N_3496,N_3344);
or U4008 (N_4008,N_3439,N_3163);
and U4009 (N_4009,N_3277,N_3484);
or U4010 (N_4010,N_3449,N_3272);
and U4011 (N_4011,N_3074,N_3012);
nor U4012 (N_4012,N_3366,N_3194);
xor U4013 (N_4013,N_3248,N_3200);
xor U4014 (N_4014,N_3464,N_3293);
nor U4015 (N_4015,N_3393,N_3056);
nand U4016 (N_4016,N_3162,N_3238);
or U4017 (N_4017,N_3745,N_3110);
and U4018 (N_4018,N_3450,N_3720);
or U4019 (N_4019,N_3097,N_3730);
xnor U4020 (N_4020,N_3437,N_3330);
or U4021 (N_4021,N_3249,N_3521);
nand U4022 (N_4022,N_3420,N_3683);
xnor U4023 (N_4023,N_3679,N_3666);
xor U4024 (N_4024,N_3009,N_3541);
or U4025 (N_4025,N_3328,N_3635);
and U4026 (N_4026,N_3322,N_3539);
nor U4027 (N_4027,N_3600,N_3040);
xnor U4028 (N_4028,N_3624,N_3729);
or U4029 (N_4029,N_3142,N_3444);
or U4030 (N_4030,N_3669,N_3076);
and U4031 (N_4031,N_3577,N_3329);
nor U4032 (N_4032,N_3542,N_3654);
nand U4033 (N_4033,N_3463,N_3231);
nor U4034 (N_4034,N_3741,N_3005);
xor U4035 (N_4035,N_3726,N_3353);
and U4036 (N_4036,N_3719,N_3108);
nor U4037 (N_4037,N_3124,N_3120);
nor U4038 (N_4038,N_3362,N_3030);
nor U4039 (N_4039,N_3145,N_3477);
nor U4040 (N_4040,N_3660,N_3370);
nand U4041 (N_4041,N_3646,N_3026);
xor U4042 (N_4042,N_3743,N_3114);
and U4043 (N_4043,N_3427,N_3460);
nand U4044 (N_4044,N_3591,N_3302);
or U4045 (N_4045,N_3475,N_3359);
xnor U4046 (N_4046,N_3738,N_3724);
xnor U4047 (N_4047,N_3230,N_3400);
xnor U4048 (N_4048,N_3392,N_3511);
or U4049 (N_4049,N_3735,N_3687);
nand U4050 (N_4050,N_3471,N_3647);
xor U4051 (N_4051,N_3116,N_3091);
or U4052 (N_4052,N_3265,N_3273);
xor U4053 (N_4053,N_3746,N_3742);
xnor U4054 (N_4054,N_3391,N_3381);
and U4055 (N_4055,N_3527,N_3454);
xnor U4056 (N_4056,N_3317,N_3642);
and U4057 (N_4057,N_3269,N_3595);
nand U4058 (N_4058,N_3551,N_3636);
and U4059 (N_4059,N_3611,N_3261);
xor U4060 (N_4060,N_3594,N_3445);
or U4061 (N_4061,N_3686,N_3325);
or U4062 (N_4062,N_3709,N_3700);
xor U4063 (N_4063,N_3013,N_3309);
xnor U4064 (N_4064,N_3303,N_3209);
nor U4065 (N_4065,N_3350,N_3308);
and U4066 (N_4066,N_3490,N_3147);
and U4067 (N_4067,N_3523,N_3379);
nand U4068 (N_4068,N_3731,N_3045);
and U4069 (N_4069,N_3502,N_3134);
or U4070 (N_4070,N_3151,N_3453);
xnor U4071 (N_4071,N_3501,N_3098);
and U4072 (N_4072,N_3268,N_3341);
xnor U4073 (N_4073,N_3569,N_3002);
xor U4074 (N_4074,N_3459,N_3224);
xnor U4075 (N_4075,N_3084,N_3416);
nor U4076 (N_4076,N_3514,N_3701);
and U4077 (N_4077,N_3205,N_3468);
or U4078 (N_4078,N_3332,N_3562);
xnor U4079 (N_4079,N_3639,N_3019);
or U4080 (N_4080,N_3190,N_3519);
nand U4081 (N_4081,N_3627,N_3253);
nand U4082 (N_4082,N_3320,N_3351);
xnor U4083 (N_4083,N_3363,N_3652);
nand U4084 (N_4084,N_3395,N_3251);
nor U4085 (N_4085,N_3010,N_3207);
nand U4086 (N_4086,N_3173,N_3582);
or U4087 (N_4087,N_3707,N_3566);
nor U4088 (N_4088,N_3189,N_3291);
and U4089 (N_4089,N_3422,N_3544);
xor U4090 (N_4090,N_3170,N_3561);
nor U4091 (N_4091,N_3327,N_3270);
or U4092 (N_4092,N_3160,N_3237);
or U4093 (N_4093,N_3494,N_3069);
xor U4094 (N_4094,N_3188,N_3008);
or U4095 (N_4095,N_3374,N_3376);
nor U4096 (N_4096,N_3081,N_3031);
or U4097 (N_4097,N_3507,N_3338);
nor U4098 (N_4098,N_3451,N_3609);
nor U4099 (N_4099,N_3614,N_3225);
nand U4100 (N_4100,N_3412,N_3706);
xnor U4101 (N_4101,N_3311,N_3640);
xnor U4102 (N_4102,N_3369,N_3711);
nand U4103 (N_4103,N_3089,N_3693);
xnor U4104 (N_4104,N_3508,N_3512);
nand U4105 (N_4105,N_3239,N_3564);
or U4106 (N_4106,N_3584,N_3470);
nand U4107 (N_4107,N_3739,N_3242);
and U4108 (N_4108,N_3402,N_3324);
xnor U4109 (N_4109,N_3385,N_3334);
xnor U4110 (N_4110,N_3032,N_3284);
nand U4111 (N_4111,N_3378,N_3547);
nor U4112 (N_4112,N_3573,N_3538);
xnor U4113 (N_4113,N_3171,N_3491);
nor U4114 (N_4114,N_3478,N_3386);
nand U4115 (N_4115,N_3264,N_3373);
and U4116 (N_4116,N_3358,N_3187);
nor U4117 (N_4117,N_3167,N_3506);
xnor U4118 (N_4118,N_3632,N_3537);
xor U4119 (N_4119,N_3637,N_3534);
and U4120 (N_4120,N_3033,N_3246);
xor U4121 (N_4121,N_3429,N_3240);
or U4122 (N_4122,N_3387,N_3747);
nand U4123 (N_4123,N_3410,N_3712);
nand U4124 (N_4124,N_3434,N_3192);
and U4125 (N_4125,N_3162,N_3284);
xor U4126 (N_4126,N_3060,N_3225);
xor U4127 (N_4127,N_3283,N_3049);
nor U4128 (N_4128,N_3517,N_3481);
nor U4129 (N_4129,N_3456,N_3103);
xnor U4130 (N_4130,N_3163,N_3595);
xnor U4131 (N_4131,N_3023,N_3633);
xnor U4132 (N_4132,N_3389,N_3605);
or U4133 (N_4133,N_3379,N_3485);
or U4134 (N_4134,N_3012,N_3535);
and U4135 (N_4135,N_3316,N_3551);
or U4136 (N_4136,N_3463,N_3513);
nor U4137 (N_4137,N_3065,N_3699);
nand U4138 (N_4138,N_3202,N_3036);
nor U4139 (N_4139,N_3265,N_3529);
and U4140 (N_4140,N_3155,N_3458);
and U4141 (N_4141,N_3595,N_3526);
or U4142 (N_4142,N_3407,N_3408);
and U4143 (N_4143,N_3598,N_3372);
and U4144 (N_4144,N_3086,N_3105);
nor U4145 (N_4145,N_3719,N_3121);
or U4146 (N_4146,N_3246,N_3455);
nand U4147 (N_4147,N_3519,N_3334);
or U4148 (N_4148,N_3326,N_3515);
xor U4149 (N_4149,N_3434,N_3671);
or U4150 (N_4150,N_3273,N_3291);
xnor U4151 (N_4151,N_3670,N_3201);
and U4152 (N_4152,N_3191,N_3657);
xnor U4153 (N_4153,N_3387,N_3401);
and U4154 (N_4154,N_3087,N_3496);
or U4155 (N_4155,N_3209,N_3092);
xor U4156 (N_4156,N_3015,N_3216);
nand U4157 (N_4157,N_3266,N_3394);
nand U4158 (N_4158,N_3075,N_3521);
nand U4159 (N_4159,N_3621,N_3431);
or U4160 (N_4160,N_3199,N_3584);
nand U4161 (N_4161,N_3566,N_3218);
and U4162 (N_4162,N_3054,N_3650);
and U4163 (N_4163,N_3662,N_3518);
nand U4164 (N_4164,N_3491,N_3595);
and U4165 (N_4165,N_3667,N_3565);
and U4166 (N_4166,N_3227,N_3125);
or U4167 (N_4167,N_3382,N_3550);
or U4168 (N_4168,N_3069,N_3612);
or U4169 (N_4169,N_3204,N_3474);
or U4170 (N_4170,N_3593,N_3317);
or U4171 (N_4171,N_3734,N_3641);
xnor U4172 (N_4172,N_3313,N_3260);
xnor U4173 (N_4173,N_3529,N_3371);
nor U4174 (N_4174,N_3072,N_3466);
and U4175 (N_4175,N_3517,N_3713);
or U4176 (N_4176,N_3568,N_3128);
xor U4177 (N_4177,N_3299,N_3111);
and U4178 (N_4178,N_3023,N_3067);
xor U4179 (N_4179,N_3495,N_3052);
or U4180 (N_4180,N_3148,N_3036);
or U4181 (N_4181,N_3515,N_3396);
and U4182 (N_4182,N_3728,N_3192);
nand U4183 (N_4183,N_3274,N_3711);
xnor U4184 (N_4184,N_3345,N_3136);
nor U4185 (N_4185,N_3342,N_3631);
or U4186 (N_4186,N_3387,N_3408);
nor U4187 (N_4187,N_3659,N_3090);
nand U4188 (N_4188,N_3561,N_3557);
nor U4189 (N_4189,N_3039,N_3431);
xnor U4190 (N_4190,N_3419,N_3052);
or U4191 (N_4191,N_3669,N_3374);
or U4192 (N_4192,N_3562,N_3283);
and U4193 (N_4193,N_3699,N_3716);
nand U4194 (N_4194,N_3415,N_3567);
nor U4195 (N_4195,N_3730,N_3339);
xor U4196 (N_4196,N_3105,N_3178);
and U4197 (N_4197,N_3061,N_3459);
nand U4198 (N_4198,N_3155,N_3328);
xnor U4199 (N_4199,N_3466,N_3167);
xnor U4200 (N_4200,N_3366,N_3487);
nand U4201 (N_4201,N_3575,N_3369);
xnor U4202 (N_4202,N_3656,N_3205);
nand U4203 (N_4203,N_3377,N_3129);
nor U4204 (N_4204,N_3207,N_3017);
xor U4205 (N_4205,N_3090,N_3655);
xnor U4206 (N_4206,N_3455,N_3091);
xnor U4207 (N_4207,N_3243,N_3287);
and U4208 (N_4208,N_3415,N_3401);
and U4209 (N_4209,N_3169,N_3721);
or U4210 (N_4210,N_3358,N_3099);
or U4211 (N_4211,N_3319,N_3248);
or U4212 (N_4212,N_3518,N_3211);
or U4213 (N_4213,N_3190,N_3344);
xor U4214 (N_4214,N_3164,N_3244);
nand U4215 (N_4215,N_3682,N_3595);
or U4216 (N_4216,N_3504,N_3015);
nand U4217 (N_4217,N_3201,N_3726);
nand U4218 (N_4218,N_3019,N_3347);
and U4219 (N_4219,N_3711,N_3674);
nand U4220 (N_4220,N_3024,N_3346);
or U4221 (N_4221,N_3385,N_3481);
nand U4222 (N_4222,N_3169,N_3206);
nand U4223 (N_4223,N_3619,N_3621);
or U4224 (N_4224,N_3584,N_3001);
and U4225 (N_4225,N_3601,N_3302);
and U4226 (N_4226,N_3390,N_3458);
nor U4227 (N_4227,N_3679,N_3688);
nand U4228 (N_4228,N_3690,N_3610);
and U4229 (N_4229,N_3536,N_3439);
nor U4230 (N_4230,N_3261,N_3305);
nand U4231 (N_4231,N_3415,N_3265);
and U4232 (N_4232,N_3283,N_3515);
nand U4233 (N_4233,N_3030,N_3643);
and U4234 (N_4234,N_3567,N_3524);
and U4235 (N_4235,N_3443,N_3262);
or U4236 (N_4236,N_3457,N_3312);
xor U4237 (N_4237,N_3641,N_3441);
nand U4238 (N_4238,N_3724,N_3100);
nor U4239 (N_4239,N_3630,N_3333);
nor U4240 (N_4240,N_3041,N_3021);
or U4241 (N_4241,N_3067,N_3103);
xor U4242 (N_4242,N_3651,N_3462);
xor U4243 (N_4243,N_3143,N_3678);
nor U4244 (N_4244,N_3501,N_3055);
nand U4245 (N_4245,N_3321,N_3695);
nor U4246 (N_4246,N_3703,N_3579);
nand U4247 (N_4247,N_3507,N_3705);
nand U4248 (N_4248,N_3477,N_3484);
and U4249 (N_4249,N_3475,N_3704);
xor U4250 (N_4250,N_3615,N_3744);
nand U4251 (N_4251,N_3102,N_3082);
nor U4252 (N_4252,N_3155,N_3287);
nand U4253 (N_4253,N_3375,N_3490);
nor U4254 (N_4254,N_3140,N_3170);
or U4255 (N_4255,N_3652,N_3514);
nand U4256 (N_4256,N_3411,N_3701);
or U4257 (N_4257,N_3218,N_3707);
or U4258 (N_4258,N_3007,N_3637);
xor U4259 (N_4259,N_3159,N_3624);
xor U4260 (N_4260,N_3142,N_3091);
or U4261 (N_4261,N_3477,N_3736);
xor U4262 (N_4262,N_3532,N_3742);
or U4263 (N_4263,N_3368,N_3041);
xnor U4264 (N_4264,N_3327,N_3631);
nor U4265 (N_4265,N_3610,N_3395);
or U4266 (N_4266,N_3256,N_3735);
nor U4267 (N_4267,N_3194,N_3126);
nand U4268 (N_4268,N_3359,N_3189);
and U4269 (N_4269,N_3571,N_3001);
nor U4270 (N_4270,N_3075,N_3373);
and U4271 (N_4271,N_3664,N_3651);
xnor U4272 (N_4272,N_3632,N_3284);
xnor U4273 (N_4273,N_3395,N_3048);
and U4274 (N_4274,N_3063,N_3360);
and U4275 (N_4275,N_3077,N_3173);
and U4276 (N_4276,N_3034,N_3330);
or U4277 (N_4277,N_3095,N_3655);
or U4278 (N_4278,N_3159,N_3359);
and U4279 (N_4279,N_3542,N_3283);
or U4280 (N_4280,N_3681,N_3619);
nor U4281 (N_4281,N_3267,N_3331);
or U4282 (N_4282,N_3424,N_3231);
nor U4283 (N_4283,N_3346,N_3418);
xnor U4284 (N_4284,N_3274,N_3514);
and U4285 (N_4285,N_3261,N_3313);
nand U4286 (N_4286,N_3102,N_3479);
or U4287 (N_4287,N_3539,N_3737);
nand U4288 (N_4288,N_3582,N_3698);
xor U4289 (N_4289,N_3589,N_3428);
xor U4290 (N_4290,N_3695,N_3550);
or U4291 (N_4291,N_3349,N_3218);
nor U4292 (N_4292,N_3184,N_3198);
nor U4293 (N_4293,N_3176,N_3685);
xor U4294 (N_4294,N_3588,N_3011);
nor U4295 (N_4295,N_3123,N_3598);
xnor U4296 (N_4296,N_3550,N_3211);
nor U4297 (N_4297,N_3191,N_3117);
xnor U4298 (N_4298,N_3476,N_3024);
and U4299 (N_4299,N_3237,N_3636);
nor U4300 (N_4300,N_3389,N_3459);
nor U4301 (N_4301,N_3502,N_3226);
nand U4302 (N_4302,N_3261,N_3724);
or U4303 (N_4303,N_3004,N_3531);
and U4304 (N_4304,N_3206,N_3027);
xnor U4305 (N_4305,N_3571,N_3134);
nor U4306 (N_4306,N_3268,N_3469);
or U4307 (N_4307,N_3059,N_3724);
xor U4308 (N_4308,N_3603,N_3376);
nand U4309 (N_4309,N_3388,N_3048);
nor U4310 (N_4310,N_3286,N_3007);
and U4311 (N_4311,N_3401,N_3571);
and U4312 (N_4312,N_3689,N_3051);
nor U4313 (N_4313,N_3136,N_3125);
or U4314 (N_4314,N_3045,N_3202);
xor U4315 (N_4315,N_3519,N_3551);
nand U4316 (N_4316,N_3030,N_3430);
or U4317 (N_4317,N_3530,N_3424);
nor U4318 (N_4318,N_3613,N_3724);
xor U4319 (N_4319,N_3220,N_3020);
or U4320 (N_4320,N_3500,N_3524);
nand U4321 (N_4321,N_3485,N_3486);
nand U4322 (N_4322,N_3510,N_3363);
and U4323 (N_4323,N_3728,N_3107);
and U4324 (N_4324,N_3122,N_3291);
and U4325 (N_4325,N_3267,N_3597);
and U4326 (N_4326,N_3148,N_3479);
or U4327 (N_4327,N_3400,N_3725);
and U4328 (N_4328,N_3619,N_3073);
and U4329 (N_4329,N_3041,N_3319);
or U4330 (N_4330,N_3395,N_3068);
nand U4331 (N_4331,N_3464,N_3690);
or U4332 (N_4332,N_3317,N_3411);
nand U4333 (N_4333,N_3380,N_3370);
or U4334 (N_4334,N_3731,N_3258);
and U4335 (N_4335,N_3690,N_3175);
and U4336 (N_4336,N_3126,N_3444);
nand U4337 (N_4337,N_3173,N_3344);
or U4338 (N_4338,N_3503,N_3000);
and U4339 (N_4339,N_3231,N_3095);
nand U4340 (N_4340,N_3097,N_3366);
and U4341 (N_4341,N_3006,N_3044);
nand U4342 (N_4342,N_3294,N_3550);
nor U4343 (N_4343,N_3317,N_3600);
xor U4344 (N_4344,N_3077,N_3285);
nor U4345 (N_4345,N_3023,N_3392);
and U4346 (N_4346,N_3230,N_3014);
and U4347 (N_4347,N_3200,N_3316);
nor U4348 (N_4348,N_3628,N_3111);
or U4349 (N_4349,N_3447,N_3101);
nand U4350 (N_4350,N_3230,N_3387);
or U4351 (N_4351,N_3178,N_3465);
xnor U4352 (N_4352,N_3538,N_3641);
or U4353 (N_4353,N_3707,N_3426);
or U4354 (N_4354,N_3588,N_3343);
nor U4355 (N_4355,N_3477,N_3334);
xor U4356 (N_4356,N_3687,N_3741);
or U4357 (N_4357,N_3090,N_3451);
xor U4358 (N_4358,N_3237,N_3425);
nor U4359 (N_4359,N_3204,N_3465);
nor U4360 (N_4360,N_3646,N_3032);
nor U4361 (N_4361,N_3271,N_3731);
or U4362 (N_4362,N_3222,N_3375);
nand U4363 (N_4363,N_3025,N_3506);
nand U4364 (N_4364,N_3155,N_3680);
nor U4365 (N_4365,N_3718,N_3422);
xor U4366 (N_4366,N_3581,N_3415);
nor U4367 (N_4367,N_3604,N_3320);
nand U4368 (N_4368,N_3084,N_3593);
and U4369 (N_4369,N_3426,N_3474);
xor U4370 (N_4370,N_3140,N_3313);
xor U4371 (N_4371,N_3200,N_3550);
and U4372 (N_4372,N_3363,N_3619);
nor U4373 (N_4373,N_3359,N_3512);
nand U4374 (N_4374,N_3577,N_3330);
or U4375 (N_4375,N_3287,N_3333);
and U4376 (N_4376,N_3465,N_3274);
or U4377 (N_4377,N_3513,N_3460);
and U4378 (N_4378,N_3149,N_3393);
nor U4379 (N_4379,N_3642,N_3436);
nor U4380 (N_4380,N_3702,N_3125);
nand U4381 (N_4381,N_3180,N_3094);
and U4382 (N_4382,N_3001,N_3017);
and U4383 (N_4383,N_3345,N_3296);
or U4384 (N_4384,N_3732,N_3191);
or U4385 (N_4385,N_3566,N_3079);
and U4386 (N_4386,N_3313,N_3089);
nand U4387 (N_4387,N_3465,N_3307);
xor U4388 (N_4388,N_3468,N_3600);
and U4389 (N_4389,N_3631,N_3744);
or U4390 (N_4390,N_3578,N_3453);
and U4391 (N_4391,N_3432,N_3172);
xor U4392 (N_4392,N_3447,N_3669);
nor U4393 (N_4393,N_3114,N_3486);
xnor U4394 (N_4394,N_3342,N_3375);
nand U4395 (N_4395,N_3303,N_3063);
nand U4396 (N_4396,N_3181,N_3631);
or U4397 (N_4397,N_3644,N_3558);
nand U4398 (N_4398,N_3502,N_3515);
nor U4399 (N_4399,N_3699,N_3118);
or U4400 (N_4400,N_3264,N_3404);
nand U4401 (N_4401,N_3547,N_3054);
or U4402 (N_4402,N_3393,N_3748);
xnor U4403 (N_4403,N_3178,N_3017);
nand U4404 (N_4404,N_3146,N_3423);
xor U4405 (N_4405,N_3481,N_3173);
and U4406 (N_4406,N_3423,N_3135);
xnor U4407 (N_4407,N_3353,N_3480);
or U4408 (N_4408,N_3596,N_3466);
xor U4409 (N_4409,N_3430,N_3672);
or U4410 (N_4410,N_3486,N_3233);
nor U4411 (N_4411,N_3191,N_3238);
xnor U4412 (N_4412,N_3510,N_3589);
nor U4413 (N_4413,N_3272,N_3695);
or U4414 (N_4414,N_3119,N_3674);
xor U4415 (N_4415,N_3636,N_3717);
nor U4416 (N_4416,N_3284,N_3639);
and U4417 (N_4417,N_3223,N_3670);
and U4418 (N_4418,N_3641,N_3173);
nor U4419 (N_4419,N_3616,N_3208);
xnor U4420 (N_4420,N_3084,N_3318);
xor U4421 (N_4421,N_3153,N_3355);
or U4422 (N_4422,N_3235,N_3585);
xor U4423 (N_4423,N_3355,N_3489);
and U4424 (N_4424,N_3106,N_3602);
nor U4425 (N_4425,N_3312,N_3205);
and U4426 (N_4426,N_3155,N_3118);
xor U4427 (N_4427,N_3047,N_3492);
nand U4428 (N_4428,N_3677,N_3340);
nand U4429 (N_4429,N_3237,N_3484);
or U4430 (N_4430,N_3106,N_3422);
or U4431 (N_4431,N_3701,N_3595);
xor U4432 (N_4432,N_3422,N_3268);
nor U4433 (N_4433,N_3307,N_3002);
or U4434 (N_4434,N_3113,N_3148);
and U4435 (N_4435,N_3134,N_3023);
and U4436 (N_4436,N_3026,N_3324);
xor U4437 (N_4437,N_3246,N_3504);
nand U4438 (N_4438,N_3244,N_3189);
or U4439 (N_4439,N_3662,N_3066);
or U4440 (N_4440,N_3185,N_3708);
or U4441 (N_4441,N_3449,N_3414);
or U4442 (N_4442,N_3568,N_3567);
nand U4443 (N_4443,N_3448,N_3555);
or U4444 (N_4444,N_3004,N_3069);
xnor U4445 (N_4445,N_3739,N_3221);
nand U4446 (N_4446,N_3673,N_3445);
and U4447 (N_4447,N_3287,N_3343);
and U4448 (N_4448,N_3426,N_3161);
and U4449 (N_4449,N_3539,N_3332);
and U4450 (N_4450,N_3337,N_3389);
xor U4451 (N_4451,N_3471,N_3005);
xnor U4452 (N_4452,N_3317,N_3277);
and U4453 (N_4453,N_3473,N_3231);
xnor U4454 (N_4454,N_3054,N_3719);
nor U4455 (N_4455,N_3661,N_3399);
nor U4456 (N_4456,N_3563,N_3573);
xnor U4457 (N_4457,N_3147,N_3201);
nand U4458 (N_4458,N_3208,N_3408);
nor U4459 (N_4459,N_3662,N_3475);
xnor U4460 (N_4460,N_3522,N_3285);
nor U4461 (N_4461,N_3099,N_3402);
or U4462 (N_4462,N_3341,N_3083);
nor U4463 (N_4463,N_3276,N_3538);
nand U4464 (N_4464,N_3015,N_3716);
or U4465 (N_4465,N_3211,N_3392);
and U4466 (N_4466,N_3140,N_3615);
nand U4467 (N_4467,N_3261,N_3237);
or U4468 (N_4468,N_3294,N_3224);
nand U4469 (N_4469,N_3078,N_3065);
nand U4470 (N_4470,N_3571,N_3347);
or U4471 (N_4471,N_3058,N_3571);
nand U4472 (N_4472,N_3736,N_3622);
or U4473 (N_4473,N_3287,N_3615);
or U4474 (N_4474,N_3098,N_3223);
or U4475 (N_4475,N_3005,N_3273);
nand U4476 (N_4476,N_3381,N_3695);
or U4477 (N_4477,N_3089,N_3369);
or U4478 (N_4478,N_3412,N_3230);
xnor U4479 (N_4479,N_3611,N_3683);
nor U4480 (N_4480,N_3301,N_3449);
nand U4481 (N_4481,N_3609,N_3039);
xor U4482 (N_4482,N_3261,N_3641);
nand U4483 (N_4483,N_3151,N_3047);
nand U4484 (N_4484,N_3742,N_3724);
nand U4485 (N_4485,N_3695,N_3391);
nand U4486 (N_4486,N_3555,N_3526);
or U4487 (N_4487,N_3277,N_3062);
and U4488 (N_4488,N_3576,N_3169);
xnor U4489 (N_4489,N_3586,N_3598);
or U4490 (N_4490,N_3728,N_3746);
or U4491 (N_4491,N_3261,N_3233);
xor U4492 (N_4492,N_3511,N_3240);
nand U4493 (N_4493,N_3237,N_3453);
and U4494 (N_4494,N_3669,N_3177);
and U4495 (N_4495,N_3124,N_3549);
or U4496 (N_4496,N_3327,N_3478);
nand U4497 (N_4497,N_3060,N_3226);
and U4498 (N_4498,N_3449,N_3307);
nand U4499 (N_4499,N_3115,N_3144);
nand U4500 (N_4500,N_4319,N_3842);
xor U4501 (N_4501,N_3957,N_4333);
or U4502 (N_4502,N_3774,N_4050);
nand U4503 (N_4503,N_4488,N_3947);
xnor U4504 (N_4504,N_3963,N_4002);
or U4505 (N_4505,N_4350,N_4043);
and U4506 (N_4506,N_4389,N_4300);
or U4507 (N_4507,N_4192,N_4038);
or U4508 (N_4508,N_4453,N_3802);
or U4509 (N_4509,N_4281,N_4267);
xnor U4510 (N_4510,N_4285,N_3845);
xnor U4511 (N_4511,N_4308,N_4134);
or U4512 (N_4512,N_4107,N_4046);
and U4513 (N_4513,N_3884,N_3970);
nor U4514 (N_4514,N_4339,N_3992);
and U4515 (N_4515,N_4039,N_4233);
nand U4516 (N_4516,N_4313,N_4380);
xor U4517 (N_4517,N_4329,N_4222);
or U4518 (N_4518,N_4030,N_4179);
or U4519 (N_4519,N_3852,N_4425);
and U4520 (N_4520,N_4460,N_3848);
or U4521 (N_4521,N_4141,N_4013);
nand U4522 (N_4522,N_4060,N_4074);
nand U4523 (N_4523,N_4177,N_4098);
and U4524 (N_4524,N_3795,N_3889);
or U4525 (N_4525,N_3960,N_4197);
nand U4526 (N_4526,N_3891,N_4398);
or U4527 (N_4527,N_4131,N_3765);
xnor U4528 (N_4528,N_4409,N_3792);
nand U4529 (N_4529,N_4076,N_3926);
nand U4530 (N_4530,N_4492,N_4372);
xor U4531 (N_4531,N_3937,N_4396);
nor U4532 (N_4532,N_4408,N_4143);
xnor U4533 (N_4533,N_4364,N_4070);
nand U4534 (N_4534,N_4496,N_3978);
nor U4535 (N_4535,N_4108,N_4101);
nor U4536 (N_4536,N_4142,N_3850);
or U4537 (N_4537,N_3953,N_4088);
nand U4538 (N_4538,N_3951,N_4041);
nand U4539 (N_4539,N_4036,N_4348);
xor U4540 (N_4540,N_4057,N_4152);
and U4541 (N_4541,N_4354,N_4176);
and U4542 (N_4542,N_3982,N_4357);
nor U4543 (N_4543,N_4309,N_3836);
xor U4544 (N_4544,N_4145,N_4017);
or U4545 (N_4545,N_3780,N_3824);
nor U4546 (N_4546,N_4273,N_4183);
or U4547 (N_4547,N_3858,N_4307);
or U4548 (N_4548,N_4336,N_4465);
nand U4549 (N_4549,N_3775,N_3837);
and U4550 (N_4550,N_4114,N_4356);
and U4551 (N_4551,N_4399,N_3994);
or U4552 (N_4552,N_4201,N_4000);
nor U4553 (N_4553,N_3799,N_3929);
nor U4554 (N_4554,N_3855,N_3877);
nand U4555 (N_4555,N_3965,N_3844);
and U4556 (N_4556,N_3777,N_3804);
and U4557 (N_4557,N_3898,N_4462);
nand U4558 (N_4558,N_4213,N_4484);
nor U4559 (N_4559,N_4432,N_4424);
xor U4560 (N_4560,N_3909,N_3961);
xor U4561 (N_4561,N_4353,N_3991);
and U4562 (N_4562,N_3779,N_3820);
nor U4563 (N_4563,N_3969,N_4054);
nand U4564 (N_4564,N_3871,N_4387);
xor U4565 (N_4565,N_4044,N_4137);
nor U4566 (N_4566,N_4006,N_4414);
nand U4567 (N_4567,N_4156,N_4181);
xor U4568 (N_4568,N_3921,N_3757);
nand U4569 (N_4569,N_4199,N_4022);
and U4570 (N_4570,N_3800,N_4327);
nor U4571 (N_4571,N_4328,N_4477);
xnor U4572 (N_4572,N_4311,N_4234);
or U4573 (N_4573,N_4175,N_4272);
or U4574 (N_4574,N_4191,N_4338);
and U4575 (N_4575,N_4132,N_3834);
nand U4576 (N_4576,N_4130,N_4047);
xor U4577 (N_4577,N_4069,N_3812);
nand U4578 (N_4578,N_3752,N_4445);
nand U4579 (N_4579,N_4485,N_4472);
xnor U4580 (N_4580,N_4037,N_4276);
nor U4581 (N_4581,N_4349,N_4494);
and U4582 (N_4582,N_4253,N_3958);
nand U4583 (N_4583,N_4119,N_3797);
nor U4584 (N_4584,N_4094,N_3764);
nand U4585 (N_4585,N_4158,N_3928);
and U4586 (N_4586,N_4301,N_3756);
nor U4587 (N_4587,N_3810,N_4490);
or U4588 (N_4588,N_4383,N_3959);
and U4589 (N_4589,N_3856,N_3945);
xor U4590 (N_4590,N_3995,N_4246);
and U4591 (N_4591,N_4099,N_4478);
and U4592 (N_4592,N_3843,N_4026);
nand U4593 (N_4593,N_3751,N_4025);
nand U4594 (N_4594,N_3789,N_4100);
nor U4595 (N_4595,N_4255,N_4284);
or U4596 (N_4596,N_3750,N_4450);
nor U4597 (N_4597,N_4148,N_3767);
or U4598 (N_4598,N_4056,N_3754);
xnor U4599 (N_4599,N_4404,N_3830);
or U4600 (N_4600,N_4227,N_4342);
or U4601 (N_4601,N_4378,N_4420);
and U4602 (N_4602,N_4335,N_3999);
nand U4603 (N_4603,N_4391,N_4105);
and U4604 (N_4604,N_4304,N_4456);
xnor U4605 (N_4605,N_3861,N_4080);
and U4606 (N_4606,N_4412,N_4431);
xnor U4607 (N_4607,N_3972,N_4280);
nand U4608 (N_4608,N_4402,N_3930);
or U4609 (N_4609,N_3847,N_4097);
nor U4610 (N_4610,N_4318,N_3949);
xor U4611 (N_4611,N_4242,N_3897);
and U4612 (N_4612,N_4049,N_4212);
and U4613 (N_4613,N_4205,N_4452);
nand U4614 (N_4614,N_4157,N_4249);
nand U4615 (N_4615,N_4454,N_4189);
xnor U4616 (N_4616,N_3827,N_4180);
nand U4617 (N_4617,N_4194,N_3760);
and U4618 (N_4618,N_4208,N_3910);
or U4619 (N_4619,N_4048,N_4239);
nor U4620 (N_4620,N_4103,N_3817);
and U4621 (N_4621,N_4340,N_4209);
and U4622 (N_4622,N_3872,N_4407);
xor U4623 (N_4623,N_4173,N_3942);
xnor U4624 (N_4624,N_4294,N_4457);
or U4625 (N_4625,N_4190,N_4287);
nand U4626 (N_4626,N_4331,N_4323);
nand U4627 (N_4627,N_4009,N_4362);
or U4628 (N_4628,N_4256,N_4116);
xor U4629 (N_4629,N_4240,N_4369);
and U4630 (N_4630,N_4363,N_4202);
nand U4631 (N_4631,N_4018,N_4257);
xor U4632 (N_4632,N_4437,N_4266);
or U4633 (N_4633,N_4358,N_4123);
and U4634 (N_4634,N_3905,N_4035);
nor U4635 (N_4635,N_4376,N_4317);
nor U4636 (N_4636,N_4290,N_4250);
and U4637 (N_4637,N_3798,N_3809);
xor U4638 (N_4638,N_4258,N_3900);
and U4639 (N_4639,N_3860,N_3796);
and U4640 (N_4640,N_3785,N_4118);
nor U4641 (N_4641,N_4235,N_3946);
and U4642 (N_4642,N_3769,N_3966);
xnor U4643 (N_4643,N_3955,N_3968);
and U4644 (N_4644,N_4373,N_4019);
xnor U4645 (N_4645,N_3857,N_3893);
nand U4646 (N_4646,N_4368,N_4226);
nor U4647 (N_4647,N_4138,N_3977);
nor U4648 (N_4648,N_4384,N_4436);
and U4649 (N_4649,N_3826,N_4014);
nor U4650 (N_4650,N_4071,N_3781);
nand U4651 (N_4651,N_4341,N_3924);
xor U4652 (N_4652,N_3931,N_3918);
xnor U4653 (N_4653,N_3934,N_3914);
or U4654 (N_4654,N_3818,N_4073);
nor U4655 (N_4655,N_4236,N_4172);
xnor U4656 (N_4656,N_4162,N_4068);
xnor U4657 (N_4657,N_4230,N_3899);
xor U4658 (N_4658,N_4493,N_4149);
nor U4659 (N_4659,N_4064,N_4449);
or U4660 (N_4660,N_4343,N_4476);
or U4661 (N_4661,N_3993,N_4229);
xnor U4662 (N_4662,N_4031,N_4413);
and U4663 (N_4663,N_4169,N_3788);
and U4664 (N_4664,N_3948,N_4161);
xor U4665 (N_4665,N_4248,N_3906);
nor U4666 (N_4666,N_3973,N_4252);
or U4667 (N_4667,N_4232,N_3922);
or U4668 (N_4668,N_3892,N_4090);
and U4669 (N_4669,N_3763,N_4001);
or U4670 (N_4670,N_4458,N_3941);
nand U4671 (N_4671,N_4224,N_3815);
nor U4672 (N_4672,N_4059,N_4225);
nand U4673 (N_4673,N_3886,N_3793);
nor U4674 (N_4674,N_4111,N_4447);
nor U4675 (N_4675,N_4461,N_4207);
nor U4676 (N_4676,N_3944,N_3878);
and U4677 (N_4677,N_4159,N_4125);
nand U4678 (N_4678,N_4223,N_3894);
and U4679 (N_4679,N_3819,N_3870);
and U4680 (N_4680,N_3933,N_4174);
or U4681 (N_4681,N_4321,N_3987);
nand U4682 (N_4682,N_4245,N_3831);
nand U4683 (N_4683,N_3825,N_4204);
nor U4684 (N_4684,N_4216,N_3854);
nor U4685 (N_4685,N_4238,N_4467);
or U4686 (N_4686,N_3998,N_4433);
nor U4687 (N_4687,N_4347,N_4489);
and U4688 (N_4688,N_4371,N_4063);
nand U4689 (N_4689,N_3916,N_4320);
or U4690 (N_4690,N_3985,N_3983);
and U4691 (N_4691,N_4382,N_4422);
nor U4692 (N_4692,N_3940,N_4167);
or U4693 (N_4693,N_3919,N_3823);
xor U4694 (N_4694,N_4040,N_4163);
nor U4695 (N_4695,N_3901,N_4196);
nand U4696 (N_4696,N_4473,N_3841);
nand U4697 (N_4697,N_4471,N_4155);
xnor U4698 (N_4698,N_4463,N_4055);
or U4699 (N_4699,N_4361,N_4482);
or U4700 (N_4700,N_4077,N_3816);
nor U4701 (N_4701,N_4128,N_3996);
or U4702 (N_4702,N_3876,N_4359);
or U4703 (N_4703,N_3853,N_3768);
or U4704 (N_4704,N_4394,N_4299);
or U4705 (N_4705,N_4459,N_3927);
and U4706 (N_4706,N_3821,N_4440);
xor U4707 (N_4707,N_3862,N_3962);
nand U4708 (N_4708,N_4279,N_4122);
and U4709 (N_4709,N_4254,N_4165);
and U4710 (N_4710,N_4296,N_4016);
nor U4711 (N_4711,N_4314,N_3975);
and U4712 (N_4712,N_4110,N_3976);
nand U4713 (N_4713,N_3932,N_4075);
and U4714 (N_4714,N_4292,N_3829);
nand U4715 (N_4715,N_4102,N_3908);
nor U4716 (N_4716,N_3935,N_3791);
nor U4717 (N_4717,N_4298,N_4390);
nor U4718 (N_4718,N_4305,N_4346);
nor U4719 (N_4719,N_3806,N_3846);
nor U4720 (N_4720,N_3794,N_4497);
or U4721 (N_4721,N_4464,N_3887);
xor U4722 (N_4722,N_4186,N_4092);
nand U4723 (N_4723,N_3849,N_3863);
xor U4724 (N_4724,N_3867,N_3784);
nand U4725 (N_4725,N_4042,N_4171);
xor U4726 (N_4726,N_4259,N_4062);
nor U4727 (N_4727,N_4081,N_3864);
xor U4728 (N_4728,N_4291,N_4244);
nand U4729 (N_4729,N_4469,N_4451);
xnor U4730 (N_4730,N_4220,N_4481);
xor U4731 (N_4731,N_3790,N_4061);
nor U4732 (N_4732,N_3895,N_3776);
and U4733 (N_4733,N_3954,N_4405);
nand U4734 (N_4734,N_4164,N_4410);
and U4735 (N_4735,N_4427,N_4474);
or U4736 (N_4736,N_3911,N_4153);
and U4737 (N_4737,N_4243,N_3939);
nand U4738 (N_4738,N_4441,N_3913);
nand U4739 (N_4739,N_4136,N_4140);
nor U4740 (N_4740,N_4417,N_3786);
and U4741 (N_4741,N_4444,N_4486);
xnor U4742 (N_4742,N_4182,N_4218);
nand U4743 (N_4743,N_4005,N_3880);
nor U4744 (N_4744,N_4475,N_3805);
nand U4745 (N_4745,N_4032,N_3936);
or U4746 (N_4746,N_3950,N_3762);
or U4747 (N_4747,N_3925,N_4127);
xor U4748 (N_4748,N_4195,N_4126);
nor U4749 (N_4749,N_4271,N_4282);
nor U4750 (N_4750,N_4479,N_3866);
nor U4751 (N_4751,N_4446,N_4367);
nor U4752 (N_4752,N_4206,N_4360);
xnor U4753 (N_4753,N_4406,N_4093);
or U4754 (N_4754,N_4228,N_4231);
nand U4755 (N_4755,N_3920,N_3865);
or U4756 (N_4756,N_3778,N_4147);
xor U4757 (N_4757,N_3967,N_4265);
nand U4758 (N_4758,N_4428,N_4277);
nand U4759 (N_4759,N_3938,N_4072);
xnor U4760 (N_4760,N_3868,N_4135);
or U4761 (N_4761,N_4418,N_4388);
nor U4762 (N_4762,N_4113,N_4095);
nor U4763 (N_4763,N_3988,N_4144);
and U4764 (N_4764,N_4434,N_4468);
nand U4765 (N_4765,N_4416,N_3885);
or U4766 (N_4766,N_4400,N_3952);
xor U4767 (N_4767,N_4010,N_4210);
nand U4768 (N_4768,N_3882,N_3755);
xor U4769 (N_4769,N_4193,N_4045);
xnor U4770 (N_4770,N_4442,N_4324);
and U4771 (N_4771,N_3770,N_4084);
xor U4772 (N_4772,N_4310,N_3851);
or U4773 (N_4773,N_4215,N_4067);
nand U4774 (N_4774,N_4011,N_4133);
or U4775 (N_4775,N_4237,N_3981);
or U4776 (N_4776,N_3801,N_3903);
or U4777 (N_4777,N_4426,N_4033);
nor U4778 (N_4778,N_4200,N_3771);
xor U4779 (N_4779,N_4377,N_4397);
nand U4780 (N_4780,N_4295,N_4121);
xor U4781 (N_4781,N_3964,N_3971);
or U4782 (N_4782,N_4015,N_4470);
or U4783 (N_4783,N_4268,N_4029);
or U4784 (N_4784,N_4495,N_4124);
and U4785 (N_4785,N_3807,N_3917);
xnor U4786 (N_4786,N_4109,N_3803);
nand U4787 (N_4787,N_4352,N_4374);
xor U4788 (N_4788,N_4221,N_4269);
nand U4789 (N_4789,N_3956,N_4178);
nand U4790 (N_4790,N_4115,N_4379);
or U4791 (N_4791,N_3890,N_4286);
nand U4792 (N_4792,N_3896,N_3813);
nor U4793 (N_4793,N_4219,N_3874);
nor U4794 (N_4794,N_4293,N_4430);
nor U4795 (N_4795,N_4435,N_4448);
nor U4796 (N_4796,N_4117,N_3943);
nor U4797 (N_4797,N_4315,N_4283);
xnor U4798 (N_4798,N_4421,N_4278);
or U4799 (N_4799,N_4012,N_4326);
xnor U4800 (N_4800,N_4483,N_4274);
xor U4801 (N_4801,N_4386,N_4403);
and U4802 (N_4802,N_4185,N_4270);
and U4803 (N_4803,N_3984,N_4297);
nor U4804 (N_4804,N_4198,N_4241);
nand U4805 (N_4805,N_4251,N_3873);
nor U4806 (N_4806,N_4146,N_4170);
and U4807 (N_4807,N_4112,N_4129);
or U4808 (N_4808,N_3989,N_4027);
nor U4809 (N_4809,N_4086,N_4082);
nor U4810 (N_4810,N_3881,N_4154);
and U4811 (N_4811,N_3811,N_4499);
xor U4812 (N_4812,N_4303,N_4085);
nand U4813 (N_4813,N_3990,N_3753);
nor U4814 (N_4814,N_4139,N_4260);
or U4815 (N_4815,N_4187,N_3838);
xor U4816 (N_4816,N_4151,N_3758);
and U4817 (N_4817,N_4007,N_3822);
or U4818 (N_4818,N_4375,N_3907);
nor U4819 (N_4819,N_4289,N_3904);
nor U4820 (N_4820,N_4487,N_4275);
nor U4821 (N_4821,N_4079,N_3814);
or U4822 (N_4822,N_4381,N_3915);
nor U4823 (N_4823,N_4439,N_3839);
or U4824 (N_4824,N_4312,N_3787);
nor U4825 (N_4825,N_3997,N_3974);
and U4826 (N_4826,N_4491,N_4203);
xor U4827 (N_4827,N_4217,N_3912);
nand U4828 (N_4828,N_4150,N_4288);
and U4829 (N_4829,N_4423,N_4322);
and U4830 (N_4830,N_4438,N_3902);
xnor U4831 (N_4831,N_4392,N_3783);
xnor U4832 (N_4832,N_4316,N_4332);
nand U4833 (N_4833,N_4366,N_4020);
xor U4834 (N_4834,N_3828,N_3869);
nand U4835 (N_4835,N_4091,N_4023);
nor U4836 (N_4836,N_4106,N_4003);
nand U4837 (N_4837,N_3782,N_4053);
xor U4838 (N_4838,N_4443,N_4188);
or U4839 (N_4839,N_3759,N_4058);
or U4840 (N_4840,N_3766,N_4355);
nor U4841 (N_4841,N_4051,N_4345);
and U4842 (N_4842,N_4104,N_4034);
or U4843 (N_4843,N_4415,N_3835);
nand U4844 (N_4844,N_3923,N_4344);
nand U4845 (N_4845,N_4306,N_3979);
xor U4846 (N_4846,N_3833,N_3875);
nand U4847 (N_4847,N_4184,N_4004);
xnor U4848 (N_4848,N_4089,N_3832);
nor U4849 (N_4849,N_4466,N_4393);
xor U4850 (N_4850,N_4498,N_4401);
and U4851 (N_4851,N_4411,N_4096);
xor U4852 (N_4852,N_4083,N_4365);
nand U4853 (N_4853,N_4211,N_4078);
xor U4854 (N_4854,N_4264,N_4052);
nand U4855 (N_4855,N_4087,N_4160);
nor U4856 (N_4856,N_3808,N_3772);
nand U4857 (N_4857,N_3883,N_3840);
nor U4858 (N_4858,N_4395,N_4455);
xnor U4859 (N_4859,N_4370,N_3761);
and U4860 (N_4860,N_3859,N_4261);
nand U4861 (N_4861,N_4480,N_3986);
nor U4862 (N_4862,N_4021,N_4024);
nand U4863 (N_4863,N_4263,N_4028);
or U4864 (N_4864,N_4008,N_3980);
and U4865 (N_4865,N_4337,N_4302);
xor U4866 (N_4866,N_4351,N_4330);
nand U4867 (N_4867,N_4419,N_4262);
or U4868 (N_4868,N_4120,N_4385);
or U4869 (N_4869,N_4429,N_4066);
nor U4870 (N_4870,N_3879,N_4065);
and U4871 (N_4871,N_4214,N_3888);
or U4872 (N_4872,N_4166,N_4168);
and U4873 (N_4873,N_4247,N_4325);
xnor U4874 (N_4874,N_4334,N_3773);
or U4875 (N_4875,N_4320,N_4376);
or U4876 (N_4876,N_3799,N_4223);
or U4877 (N_4877,N_4306,N_3786);
xnor U4878 (N_4878,N_4259,N_4448);
or U4879 (N_4879,N_4177,N_4037);
or U4880 (N_4880,N_4450,N_4356);
and U4881 (N_4881,N_3947,N_4238);
xnor U4882 (N_4882,N_3763,N_4018);
or U4883 (N_4883,N_4497,N_4488);
and U4884 (N_4884,N_4232,N_4280);
or U4885 (N_4885,N_3767,N_4362);
or U4886 (N_4886,N_4193,N_3802);
and U4887 (N_4887,N_3903,N_4392);
or U4888 (N_4888,N_3914,N_4466);
xor U4889 (N_4889,N_4460,N_4022);
or U4890 (N_4890,N_4303,N_3808);
nand U4891 (N_4891,N_4162,N_3781);
nor U4892 (N_4892,N_3971,N_4193);
or U4893 (N_4893,N_4065,N_3778);
and U4894 (N_4894,N_3939,N_3763);
and U4895 (N_4895,N_4393,N_4107);
nand U4896 (N_4896,N_4254,N_3914);
or U4897 (N_4897,N_4305,N_4303);
and U4898 (N_4898,N_4462,N_4353);
or U4899 (N_4899,N_4114,N_4165);
or U4900 (N_4900,N_4430,N_4083);
or U4901 (N_4901,N_4398,N_3930);
nand U4902 (N_4902,N_4400,N_4058);
or U4903 (N_4903,N_3970,N_4400);
or U4904 (N_4904,N_4004,N_3824);
or U4905 (N_4905,N_4211,N_3836);
nand U4906 (N_4906,N_4211,N_3945);
nand U4907 (N_4907,N_3972,N_4166);
or U4908 (N_4908,N_3923,N_4165);
or U4909 (N_4909,N_3833,N_4182);
and U4910 (N_4910,N_4274,N_4459);
nor U4911 (N_4911,N_4235,N_4417);
nand U4912 (N_4912,N_4314,N_3755);
xnor U4913 (N_4913,N_3889,N_4150);
nand U4914 (N_4914,N_4290,N_3923);
and U4915 (N_4915,N_4361,N_4457);
nor U4916 (N_4916,N_3883,N_4127);
or U4917 (N_4917,N_3810,N_4025);
nand U4918 (N_4918,N_4143,N_3828);
and U4919 (N_4919,N_4471,N_4291);
nand U4920 (N_4920,N_4171,N_4364);
or U4921 (N_4921,N_3876,N_3778);
or U4922 (N_4922,N_4411,N_4297);
nand U4923 (N_4923,N_4133,N_4450);
and U4924 (N_4924,N_4417,N_4418);
nor U4925 (N_4925,N_3898,N_3843);
or U4926 (N_4926,N_4067,N_3776);
nor U4927 (N_4927,N_4386,N_4191);
or U4928 (N_4928,N_3932,N_3942);
xor U4929 (N_4929,N_4308,N_4235);
nand U4930 (N_4930,N_4477,N_3829);
nor U4931 (N_4931,N_3897,N_4033);
nand U4932 (N_4932,N_4329,N_4236);
or U4933 (N_4933,N_3944,N_3806);
nor U4934 (N_4934,N_4001,N_4235);
or U4935 (N_4935,N_4381,N_3794);
or U4936 (N_4936,N_3857,N_4356);
or U4937 (N_4937,N_4302,N_4229);
xnor U4938 (N_4938,N_4226,N_4165);
xnor U4939 (N_4939,N_4015,N_4317);
xnor U4940 (N_4940,N_3895,N_4008);
nand U4941 (N_4941,N_4211,N_4063);
nor U4942 (N_4942,N_4340,N_3762);
nor U4943 (N_4943,N_4030,N_4161);
xnor U4944 (N_4944,N_4008,N_4435);
and U4945 (N_4945,N_4217,N_3856);
nor U4946 (N_4946,N_3770,N_3848);
and U4947 (N_4947,N_3878,N_4336);
nor U4948 (N_4948,N_4378,N_4083);
nor U4949 (N_4949,N_4096,N_4189);
xnor U4950 (N_4950,N_4240,N_3943);
nor U4951 (N_4951,N_4325,N_3812);
or U4952 (N_4952,N_3908,N_3798);
xnor U4953 (N_4953,N_4174,N_4447);
nand U4954 (N_4954,N_4257,N_4125);
and U4955 (N_4955,N_4127,N_4480);
nand U4956 (N_4956,N_3759,N_4280);
xor U4957 (N_4957,N_4193,N_4385);
and U4958 (N_4958,N_3848,N_4307);
nand U4959 (N_4959,N_4485,N_3853);
or U4960 (N_4960,N_3870,N_4329);
or U4961 (N_4961,N_4303,N_3836);
nand U4962 (N_4962,N_4043,N_4295);
xnor U4963 (N_4963,N_4083,N_3948);
nor U4964 (N_4964,N_4455,N_3949);
nor U4965 (N_4965,N_4277,N_3956);
and U4966 (N_4966,N_4430,N_3855);
nor U4967 (N_4967,N_3901,N_4306);
nor U4968 (N_4968,N_3762,N_4125);
and U4969 (N_4969,N_3821,N_3898);
nor U4970 (N_4970,N_3798,N_4242);
xnor U4971 (N_4971,N_3872,N_4199);
nor U4972 (N_4972,N_3930,N_4430);
nand U4973 (N_4973,N_3828,N_3842);
nand U4974 (N_4974,N_4200,N_3880);
and U4975 (N_4975,N_4166,N_4099);
or U4976 (N_4976,N_4441,N_4341);
xnor U4977 (N_4977,N_4457,N_4173);
or U4978 (N_4978,N_4332,N_4462);
nand U4979 (N_4979,N_4396,N_4005);
xor U4980 (N_4980,N_3768,N_4040);
xor U4981 (N_4981,N_3896,N_4015);
nand U4982 (N_4982,N_4113,N_4094);
nor U4983 (N_4983,N_4202,N_4335);
or U4984 (N_4984,N_3926,N_4172);
nor U4985 (N_4985,N_3866,N_4231);
xor U4986 (N_4986,N_4301,N_4150);
nor U4987 (N_4987,N_3755,N_4498);
and U4988 (N_4988,N_4426,N_3964);
nand U4989 (N_4989,N_3864,N_3816);
nor U4990 (N_4990,N_3946,N_4226);
nor U4991 (N_4991,N_4244,N_4241);
nand U4992 (N_4992,N_4244,N_3754);
nor U4993 (N_4993,N_3760,N_4007);
nor U4994 (N_4994,N_4106,N_3943);
nor U4995 (N_4995,N_4467,N_4086);
xnor U4996 (N_4996,N_3875,N_4164);
nor U4997 (N_4997,N_4460,N_4254);
or U4998 (N_4998,N_3930,N_4326);
or U4999 (N_4999,N_4029,N_4414);
or U5000 (N_5000,N_3902,N_3968);
and U5001 (N_5001,N_4054,N_4326);
nand U5002 (N_5002,N_4473,N_4421);
or U5003 (N_5003,N_4336,N_3918);
or U5004 (N_5004,N_3975,N_3807);
nor U5005 (N_5005,N_4133,N_4187);
or U5006 (N_5006,N_4209,N_3771);
nand U5007 (N_5007,N_4029,N_4039);
xor U5008 (N_5008,N_4408,N_4475);
nand U5009 (N_5009,N_3932,N_4479);
nand U5010 (N_5010,N_4083,N_4370);
and U5011 (N_5011,N_3807,N_3752);
and U5012 (N_5012,N_4262,N_4019);
nand U5013 (N_5013,N_3905,N_4175);
nor U5014 (N_5014,N_4122,N_4277);
nand U5015 (N_5015,N_4399,N_4345);
nor U5016 (N_5016,N_4465,N_4400);
or U5017 (N_5017,N_4274,N_3973);
nor U5018 (N_5018,N_4195,N_4409);
and U5019 (N_5019,N_3865,N_3986);
nand U5020 (N_5020,N_4368,N_4032);
xnor U5021 (N_5021,N_4429,N_4198);
xor U5022 (N_5022,N_3802,N_4112);
or U5023 (N_5023,N_4190,N_4192);
nor U5024 (N_5024,N_4334,N_4465);
nand U5025 (N_5025,N_4071,N_4007);
xor U5026 (N_5026,N_3908,N_4342);
nor U5027 (N_5027,N_3776,N_4043);
nor U5028 (N_5028,N_3867,N_3751);
nor U5029 (N_5029,N_4094,N_4133);
nand U5030 (N_5030,N_3808,N_4418);
nand U5031 (N_5031,N_3806,N_3945);
nor U5032 (N_5032,N_4094,N_4119);
nor U5033 (N_5033,N_4369,N_3838);
xor U5034 (N_5034,N_4304,N_3936);
and U5035 (N_5035,N_3769,N_4394);
or U5036 (N_5036,N_3873,N_3761);
and U5037 (N_5037,N_4400,N_3954);
nor U5038 (N_5038,N_3903,N_4353);
and U5039 (N_5039,N_4077,N_4302);
and U5040 (N_5040,N_3795,N_3789);
nor U5041 (N_5041,N_3772,N_4132);
xnor U5042 (N_5042,N_4231,N_4293);
nand U5043 (N_5043,N_3863,N_3935);
xor U5044 (N_5044,N_4080,N_4100);
and U5045 (N_5045,N_4446,N_4293);
or U5046 (N_5046,N_4124,N_4028);
and U5047 (N_5047,N_4132,N_4015);
and U5048 (N_5048,N_3905,N_4486);
or U5049 (N_5049,N_4221,N_3961);
or U5050 (N_5050,N_4052,N_4407);
nor U5051 (N_5051,N_4262,N_4439);
or U5052 (N_5052,N_4085,N_3977);
and U5053 (N_5053,N_4177,N_4305);
xnor U5054 (N_5054,N_4219,N_4118);
or U5055 (N_5055,N_4039,N_3752);
and U5056 (N_5056,N_4490,N_3965);
and U5057 (N_5057,N_4212,N_3804);
xnor U5058 (N_5058,N_4153,N_4365);
nor U5059 (N_5059,N_4332,N_4127);
and U5060 (N_5060,N_4132,N_4364);
or U5061 (N_5061,N_4223,N_4257);
xnor U5062 (N_5062,N_4245,N_4430);
xnor U5063 (N_5063,N_3838,N_4258);
or U5064 (N_5064,N_3972,N_4076);
xor U5065 (N_5065,N_4158,N_4132);
and U5066 (N_5066,N_4143,N_4064);
nor U5067 (N_5067,N_4228,N_3928);
xnor U5068 (N_5068,N_3761,N_4129);
or U5069 (N_5069,N_3944,N_4336);
nand U5070 (N_5070,N_4351,N_4004);
nand U5071 (N_5071,N_4497,N_4016);
or U5072 (N_5072,N_4175,N_4251);
xnor U5073 (N_5073,N_3818,N_3880);
or U5074 (N_5074,N_4084,N_4129);
nand U5075 (N_5075,N_4227,N_3793);
xor U5076 (N_5076,N_3950,N_4174);
nor U5077 (N_5077,N_4264,N_3867);
nor U5078 (N_5078,N_4365,N_4360);
or U5079 (N_5079,N_4159,N_3778);
or U5080 (N_5080,N_3976,N_4337);
and U5081 (N_5081,N_4289,N_3846);
nand U5082 (N_5082,N_3835,N_4268);
nand U5083 (N_5083,N_4001,N_4393);
or U5084 (N_5084,N_4240,N_4467);
or U5085 (N_5085,N_4453,N_3892);
xor U5086 (N_5086,N_3961,N_4008);
nor U5087 (N_5087,N_4391,N_4448);
xnor U5088 (N_5088,N_4303,N_3753);
nand U5089 (N_5089,N_4440,N_4386);
or U5090 (N_5090,N_3861,N_3885);
xor U5091 (N_5091,N_3981,N_4401);
xnor U5092 (N_5092,N_4306,N_4028);
nor U5093 (N_5093,N_4185,N_4308);
or U5094 (N_5094,N_3892,N_4475);
nand U5095 (N_5095,N_3932,N_4152);
xor U5096 (N_5096,N_3842,N_4391);
xor U5097 (N_5097,N_3901,N_4413);
xor U5098 (N_5098,N_4000,N_3856);
xnor U5099 (N_5099,N_3932,N_4410);
nand U5100 (N_5100,N_3800,N_4381);
xnor U5101 (N_5101,N_4048,N_4297);
or U5102 (N_5102,N_4072,N_4233);
and U5103 (N_5103,N_4181,N_4127);
nor U5104 (N_5104,N_3854,N_4325);
xnor U5105 (N_5105,N_4368,N_4110);
nand U5106 (N_5106,N_4122,N_3978);
and U5107 (N_5107,N_3909,N_4492);
nand U5108 (N_5108,N_3831,N_4102);
nand U5109 (N_5109,N_3890,N_3912);
or U5110 (N_5110,N_3764,N_4348);
xnor U5111 (N_5111,N_3782,N_4366);
and U5112 (N_5112,N_3916,N_4169);
xor U5113 (N_5113,N_4456,N_4467);
and U5114 (N_5114,N_4017,N_3941);
and U5115 (N_5115,N_3759,N_4412);
or U5116 (N_5116,N_3917,N_4098);
nand U5117 (N_5117,N_3977,N_4429);
and U5118 (N_5118,N_3768,N_4222);
xnor U5119 (N_5119,N_4159,N_3837);
and U5120 (N_5120,N_4340,N_3752);
and U5121 (N_5121,N_3923,N_4275);
xnor U5122 (N_5122,N_3753,N_3760);
nor U5123 (N_5123,N_4147,N_4071);
nor U5124 (N_5124,N_4259,N_3936);
nor U5125 (N_5125,N_4281,N_3960);
xor U5126 (N_5126,N_4416,N_4443);
or U5127 (N_5127,N_4249,N_4282);
nor U5128 (N_5128,N_4085,N_3865);
xor U5129 (N_5129,N_4077,N_4347);
xor U5130 (N_5130,N_4238,N_4384);
nand U5131 (N_5131,N_3847,N_4339);
and U5132 (N_5132,N_4309,N_4338);
xor U5133 (N_5133,N_4440,N_4377);
and U5134 (N_5134,N_4284,N_3935);
or U5135 (N_5135,N_4018,N_3943);
xor U5136 (N_5136,N_4074,N_4195);
and U5137 (N_5137,N_4484,N_4384);
and U5138 (N_5138,N_4268,N_4213);
or U5139 (N_5139,N_3837,N_4478);
and U5140 (N_5140,N_3898,N_4365);
xor U5141 (N_5141,N_4016,N_4231);
or U5142 (N_5142,N_3761,N_3959);
nand U5143 (N_5143,N_4186,N_4194);
xor U5144 (N_5144,N_3774,N_4213);
and U5145 (N_5145,N_4484,N_4118);
nand U5146 (N_5146,N_4011,N_4023);
nand U5147 (N_5147,N_4346,N_4216);
or U5148 (N_5148,N_4043,N_3997);
and U5149 (N_5149,N_3819,N_4061);
nor U5150 (N_5150,N_4477,N_4009);
nor U5151 (N_5151,N_3872,N_4157);
nand U5152 (N_5152,N_4426,N_4091);
or U5153 (N_5153,N_4420,N_4183);
or U5154 (N_5154,N_4167,N_4077);
and U5155 (N_5155,N_3858,N_4426);
or U5156 (N_5156,N_4293,N_4468);
nand U5157 (N_5157,N_3907,N_4087);
and U5158 (N_5158,N_3923,N_3751);
nor U5159 (N_5159,N_4123,N_3908);
and U5160 (N_5160,N_4208,N_4248);
and U5161 (N_5161,N_4317,N_4439);
nand U5162 (N_5162,N_3894,N_4415);
xor U5163 (N_5163,N_4296,N_4123);
or U5164 (N_5164,N_4302,N_4218);
and U5165 (N_5165,N_3903,N_4426);
or U5166 (N_5166,N_3962,N_4404);
or U5167 (N_5167,N_3774,N_4175);
nor U5168 (N_5168,N_3751,N_4288);
xor U5169 (N_5169,N_4083,N_4031);
nand U5170 (N_5170,N_4049,N_4373);
or U5171 (N_5171,N_4372,N_3964);
nor U5172 (N_5172,N_3866,N_4010);
xor U5173 (N_5173,N_4347,N_3807);
xor U5174 (N_5174,N_4308,N_4224);
or U5175 (N_5175,N_3874,N_4269);
nor U5176 (N_5176,N_4010,N_3927);
or U5177 (N_5177,N_4073,N_4027);
nand U5178 (N_5178,N_4056,N_3834);
or U5179 (N_5179,N_4124,N_3998);
nand U5180 (N_5180,N_4251,N_3854);
nor U5181 (N_5181,N_4281,N_4211);
and U5182 (N_5182,N_3818,N_4058);
xor U5183 (N_5183,N_3829,N_3894);
nor U5184 (N_5184,N_3869,N_4027);
and U5185 (N_5185,N_4306,N_3848);
nand U5186 (N_5186,N_4243,N_3856);
nand U5187 (N_5187,N_4410,N_4253);
nand U5188 (N_5188,N_3922,N_4215);
nor U5189 (N_5189,N_4454,N_4403);
xor U5190 (N_5190,N_4325,N_4017);
nand U5191 (N_5191,N_4065,N_4074);
and U5192 (N_5192,N_3957,N_3862);
xnor U5193 (N_5193,N_3974,N_3816);
or U5194 (N_5194,N_4286,N_4093);
nand U5195 (N_5195,N_4031,N_3974);
nor U5196 (N_5196,N_4042,N_4355);
xor U5197 (N_5197,N_4059,N_4438);
and U5198 (N_5198,N_3931,N_4070);
and U5199 (N_5199,N_4380,N_3805);
and U5200 (N_5200,N_3787,N_3968);
and U5201 (N_5201,N_4401,N_4165);
nand U5202 (N_5202,N_3873,N_3770);
xor U5203 (N_5203,N_4433,N_3863);
xor U5204 (N_5204,N_4379,N_4421);
or U5205 (N_5205,N_3757,N_4385);
nand U5206 (N_5206,N_4477,N_4164);
and U5207 (N_5207,N_4083,N_4159);
and U5208 (N_5208,N_3847,N_3961);
nand U5209 (N_5209,N_3946,N_4176);
xor U5210 (N_5210,N_3786,N_3867);
xnor U5211 (N_5211,N_3953,N_4129);
or U5212 (N_5212,N_4131,N_4211);
or U5213 (N_5213,N_4325,N_4284);
xnor U5214 (N_5214,N_3936,N_3765);
nor U5215 (N_5215,N_4020,N_3813);
xnor U5216 (N_5216,N_4446,N_3910);
xnor U5217 (N_5217,N_4095,N_4439);
and U5218 (N_5218,N_3946,N_4141);
nor U5219 (N_5219,N_4044,N_3854);
xnor U5220 (N_5220,N_3938,N_4423);
or U5221 (N_5221,N_4109,N_4344);
nand U5222 (N_5222,N_4087,N_3835);
xor U5223 (N_5223,N_4451,N_4238);
xor U5224 (N_5224,N_3786,N_3938);
nor U5225 (N_5225,N_4368,N_4275);
or U5226 (N_5226,N_4167,N_4360);
xnor U5227 (N_5227,N_4004,N_4179);
xor U5228 (N_5228,N_3937,N_4474);
and U5229 (N_5229,N_4422,N_3834);
nand U5230 (N_5230,N_4168,N_4352);
nor U5231 (N_5231,N_4257,N_4044);
xnor U5232 (N_5232,N_4492,N_4357);
and U5233 (N_5233,N_3850,N_4294);
nor U5234 (N_5234,N_3760,N_4056);
or U5235 (N_5235,N_3916,N_4450);
xor U5236 (N_5236,N_4358,N_4345);
or U5237 (N_5237,N_4410,N_4190);
and U5238 (N_5238,N_4291,N_4499);
nand U5239 (N_5239,N_3831,N_4029);
nor U5240 (N_5240,N_4041,N_4476);
or U5241 (N_5241,N_4453,N_3973);
or U5242 (N_5242,N_3896,N_4487);
nand U5243 (N_5243,N_4053,N_3858);
xnor U5244 (N_5244,N_4106,N_4217);
or U5245 (N_5245,N_4112,N_3855);
xnor U5246 (N_5246,N_3778,N_4223);
nand U5247 (N_5247,N_3816,N_4266);
xnor U5248 (N_5248,N_3795,N_4427);
or U5249 (N_5249,N_4226,N_3973);
nor U5250 (N_5250,N_4964,N_4884);
and U5251 (N_5251,N_4643,N_4892);
nand U5252 (N_5252,N_4834,N_4963);
nand U5253 (N_5253,N_4636,N_4865);
xnor U5254 (N_5254,N_5199,N_5109);
xor U5255 (N_5255,N_4811,N_5085);
xnor U5256 (N_5256,N_4995,N_4640);
nor U5257 (N_5257,N_5039,N_5058);
or U5258 (N_5258,N_5002,N_4912);
and U5259 (N_5259,N_5108,N_5219);
or U5260 (N_5260,N_4977,N_5176);
nor U5261 (N_5261,N_5225,N_5053);
or U5262 (N_5262,N_4530,N_4953);
nor U5263 (N_5263,N_4587,N_5060);
and U5264 (N_5264,N_5040,N_5131);
nor U5265 (N_5265,N_4999,N_4829);
xnor U5266 (N_5266,N_5232,N_5181);
nand U5267 (N_5267,N_5212,N_4684);
xor U5268 (N_5268,N_5047,N_4942);
or U5269 (N_5269,N_5187,N_4806);
and U5270 (N_5270,N_4694,N_4590);
xor U5271 (N_5271,N_4853,N_5037);
and U5272 (N_5272,N_4544,N_4948);
and U5273 (N_5273,N_4648,N_4864);
xnor U5274 (N_5274,N_5208,N_5149);
nand U5275 (N_5275,N_5209,N_4619);
nand U5276 (N_5276,N_4786,N_4564);
and U5277 (N_5277,N_4875,N_5028);
nand U5278 (N_5278,N_4848,N_5115);
or U5279 (N_5279,N_5159,N_4622);
nor U5280 (N_5280,N_4722,N_4777);
nand U5281 (N_5281,N_4713,N_5175);
nor U5282 (N_5282,N_4667,N_5155);
and U5283 (N_5283,N_5200,N_5196);
nor U5284 (N_5284,N_5154,N_4647);
nand U5285 (N_5285,N_4968,N_5026);
nand U5286 (N_5286,N_4687,N_4551);
nand U5287 (N_5287,N_4927,N_5103);
and U5288 (N_5288,N_5099,N_4507);
nor U5289 (N_5289,N_4816,N_4693);
xor U5290 (N_5290,N_5239,N_4882);
or U5291 (N_5291,N_4833,N_4651);
xnor U5292 (N_5292,N_5158,N_5083);
nand U5293 (N_5293,N_4594,N_4610);
or U5294 (N_5294,N_4889,N_4653);
and U5295 (N_5295,N_5038,N_4872);
or U5296 (N_5296,N_5162,N_4918);
xor U5297 (N_5297,N_4985,N_4814);
nand U5298 (N_5298,N_5195,N_4979);
xnor U5299 (N_5299,N_5086,N_4876);
and U5300 (N_5300,N_4855,N_5122);
and U5301 (N_5301,N_4705,N_5100);
and U5302 (N_5302,N_5130,N_5226);
nand U5303 (N_5303,N_4515,N_5142);
or U5304 (N_5304,N_4677,N_4781);
nand U5305 (N_5305,N_4826,N_4524);
and U5306 (N_5306,N_4700,N_4762);
and U5307 (N_5307,N_4825,N_4642);
or U5308 (N_5308,N_4748,N_4623);
nor U5309 (N_5309,N_4930,N_4792);
and U5310 (N_5310,N_5121,N_5170);
and U5311 (N_5311,N_4947,N_4899);
and U5312 (N_5312,N_4612,N_4845);
or U5313 (N_5313,N_4661,N_4746);
or U5314 (N_5314,N_5182,N_4593);
and U5315 (N_5315,N_5198,N_4574);
nand U5316 (N_5316,N_4832,N_4863);
nor U5317 (N_5317,N_4624,N_4670);
or U5318 (N_5318,N_4949,N_5206);
nor U5319 (N_5319,N_5042,N_4718);
and U5320 (N_5320,N_4727,N_4675);
nor U5321 (N_5321,N_4567,N_4691);
nand U5322 (N_5322,N_4514,N_4758);
nor U5323 (N_5323,N_5202,N_5024);
nor U5324 (N_5324,N_5217,N_5106);
xnor U5325 (N_5325,N_4537,N_4943);
and U5326 (N_5326,N_4645,N_4969);
and U5327 (N_5327,N_5203,N_5236);
nor U5328 (N_5328,N_5059,N_4965);
nand U5329 (N_5329,N_4575,N_4534);
nor U5330 (N_5330,N_4794,N_5055);
and U5331 (N_5331,N_4751,N_5129);
nor U5332 (N_5332,N_4565,N_4808);
or U5333 (N_5333,N_4989,N_5051);
xor U5334 (N_5334,N_5163,N_4732);
nor U5335 (N_5335,N_5010,N_5091);
nand U5336 (N_5336,N_4598,N_4662);
and U5337 (N_5337,N_4789,N_4917);
xnor U5338 (N_5338,N_4996,N_4827);
nand U5339 (N_5339,N_4915,N_5152);
xor U5340 (N_5340,N_4576,N_4568);
or U5341 (N_5341,N_5032,N_5140);
nor U5342 (N_5342,N_4980,N_4778);
or U5343 (N_5343,N_4922,N_4756);
and U5344 (N_5344,N_4743,N_4885);
nor U5345 (N_5345,N_5007,N_4951);
or U5346 (N_5346,N_4771,N_4752);
and U5347 (N_5347,N_4591,N_5240);
or U5348 (N_5348,N_5213,N_5043);
nor U5349 (N_5349,N_5146,N_4729);
and U5350 (N_5350,N_4831,N_5123);
and U5351 (N_5351,N_5183,N_5223);
xor U5352 (N_5352,N_4874,N_5077);
nand U5353 (N_5353,N_4563,N_4525);
or U5354 (N_5354,N_4749,N_4997);
nand U5355 (N_5355,N_4570,N_4500);
and U5356 (N_5356,N_4739,N_4747);
and U5357 (N_5357,N_5171,N_4618);
nor U5358 (N_5358,N_4984,N_5005);
xnor U5359 (N_5359,N_4824,N_4844);
nand U5360 (N_5360,N_5070,N_5227);
nor U5361 (N_5361,N_4501,N_4956);
nand U5362 (N_5362,N_5220,N_5003);
nand U5363 (N_5363,N_4615,N_4579);
and U5364 (N_5364,N_4644,N_4923);
nor U5365 (N_5365,N_5090,N_4913);
xor U5366 (N_5366,N_4711,N_4611);
or U5367 (N_5367,N_4641,N_5161);
or U5368 (N_5368,N_4503,N_5111);
or U5369 (N_5369,N_5190,N_4728);
or U5370 (N_5370,N_4552,N_5120);
xnor U5371 (N_5371,N_5218,N_5101);
and U5372 (N_5372,N_5082,N_4585);
nor U5373 (N_5373,N_5192,N_4907);
and U5374 (N_5374,N_4933,N_4650);
or U5375 (N_5375,N_4818,N_5138);
nand U5376 (N_5376,N_4835,N_5094);
or U5377 (N_5377,N_4609,N_4955);
or U5378 (N_5378,N_4723,N_4788);
nor U5379 (N_5379,N_4992,N_4580);
or U5380 (N_5380,N_5157,N_5097);
and U5381 (N_5381,N_4937,N_4562);
nand U5382 (N_5382,N_5143,N_4897);
nor U5383 (N_5383,N_5098,N_4740);
and U5384 (N_5384,N_5233,N_5249);
or U5385 (N_5385,N_4720,N_5001);
and U5386 (N_5386,N_4873,N_4970);
or U5387 (N_5387,N_4940,N_4664);
xnor U5388 (N_5388,N_4902,N_4685);
xor U5389 (N_5389,N_4961,N_4819);
xnor U5390 (N_5390,N_4856,N_4802);
and U5391 (N_5391,N_5193,N_5179);
or U5392 (N_5392,N_5046,N_4896);
nand U5393 (N_5393,N_4517,N_4633);
nor U5394 (N_5394,N_4854,N_4506);
or U5395 (N_5395,N_4924,N_4546);
nor U5396 (N_5396,N_4582,N_5160);
nand U5397 (N_5397,N_4656,N_4674);
or U5398 (N_5398,N_4688,N_4566);
and U5399 (N_5399,N_4807,N_4671);
or U5400 (N_5400,N_5063,N_4836);
xnor U5401 (N_5401,N_4878,N_4695);
nor U5402 (N_5402,N_4932,N_4978);
nand U5403 (N_5403,N_4604,N_4815);
nor U5404 (N_5404,N_4862,N_4505);
and U5405 (N_5405,N_4668,N_5229);
nand U5406 (N_5406,N_4513,N_4663);
nand U5407 (N_5407,N_5128,N_4511);
nand U5408 (N_5408,N_4911,N_5102);
nand U5409 (N_5409,N_5132,N_4657);
nor U5410 (N_5410,N_4621,N_4957);
and U5411 (N_5411,N_4542,N_5107);
or U5412 (N_5412,N_4608,N_4529);
nand U5413 (N_5413,N_4921,N_5216);
nor U5414 (N_5414,N_4712,N_4860);
or U5415 (N_5415,N_5167,N_4635);
xor U5416 (N_5416,N_4793,N_4795);
xor U5417 (N_5417,N_5177,N_5237);
and U5418 (N_5418,N_4724,N_5114);
xor U5419 (N_5419,N_5073,N_4810);
or U5420 (N_5420,N_4981,N_5041);
xor U5421 (N_5421,N_4689,N_4665);
nand U5422 (N_5422,N_4573,N_4772);
nand U5423 (N_5423,N_4502,N_4553);
nand U5424 (N_5424,N_4757,N_4540);
nor U5425 (N_5425,N_4851,N_5168);
nor U5426 (N_5426,N_4904,N_4822);
nor U5427 (N_5427,N_5210,N_4843);
nor U5428 (N_5428,N_5222,N_4523);
xnor U5429 (N_5429,N_4522,N_4555);
nand U5430 (N_5430,N_5069,N_4559);
nor U5431 (N_5431,N_5119,N_4881);
or U5432 (N_5432,N_4737,N_4914);
nor U5433 (N_5433,N_4767,N_5049);
xor U5434 (N_5434,N_4931,N_4982);
xor U5435 (N_5435,N_4731,N_5105);
nor U5436 (N_5436,N_4649,N_5000);
or U5437 (N_5437,N_5078,N_4859);
nor U5438 (N_5438,N_4742,N_5201);
xnor U5439 (N_5439,N_5173,N_5188);
xor U5440 (N_5440,N_5015,N_4697);
nor U5441 (N_5441,N_4538,N_4683);
nor U5442 (N_5442,N_4784,N_4646);
and U5443 (N_5443,N_4894,N_4541);
or U5444 (N_5444,N_5124,N_4583);
nor U5445 (N_5445,N_4597,N_4941);
xor U5446 (N_5446,N_4763,N_5189);
xor U5447 (N_5447,N_4858,N_4797);
and U5448 (N_5448,N_4625,N_5095);
or U5449 (N_5449,N_4837,N_4715);
and U5450 (N_5450,N_5075,N_5224);
nor U5451 (N_5451,N_4741,N_4905);
nand U5452 (N_5452,N_4765,N_4993);
nand U5453 (N_5453,N_5062,N_5084);
or U5454 (N_5454,N_4954,N_4764);
or U5455 (N_5455,N_4850,N_4880);
xnor U5456 (N_5456,N_4959,N_4785);
or U5457 (N_5457,N_5054,N_4888);
nand U5458 (N_5458,N_4659,N_4990);
nor U5459 (N_5459,N_4950,N_5166);
or U5460 (N_5460,N_4547,N_4536);
xor U5461 (N_5461,N_5074,N_4886);
xnor U5462 (N_5462,N_4589,N_4561);
xnor U5463 (N_5463,N_4987,N_5065);
nand U5464 (N_5464,N_5031,N_5066);
xnor U5465 (N_5465,N_5126,N_5081);
nand U5466 (N_5466,N_4637,N_5165);
and U5467 (N_5467,N_4813,N_4577);
nor U5468 (N_5468,N_4706,N_4988);
or U5469 (N_5469,N_4588,N_5139);
or U5470 (N_5470,N_5241,N_4535);
and U5471 (N_5471,N_5141,N_5221);
nor U5472 (N_5472,N_5185,N_4703);
xnor U5473 (N_5473,N_5174,N_4782);
nor U5474 (N_5474,N_4779,N_4869);
and U5475 (N_5475,N_4678,N_5080);
or U5476 (N_5476,N_4744,N_4972);
or U5477 (N_5477,N_4632,N_5104);
and U5478 (N_5478,N_4708,N_5035);
nand U5479 (N_5479,N_4898,N_4745);
or U5480 (N_5480,N_4849,N_5019);
or U5481 (N_5481,N_4631,N_5044);
or U5482 (N_5482,N_5033,N_5089);
and U5483 (N_5483,N_4692,N_5172);
or U5484 (N_5484,N_4916,N_4944);
and U5485 (N_5485,N_4600,N_5145);
and U5486 (N_5486,N_5048,N_4614);
nor U5487 (N_5487,N_4601,N_5092);
nand U5488 (N_5488,N_4550,N_5071);
xnor U5489 (N_5489,N_4710,N_5178);
nand U5490 (N_5490,N_4870,N_4738);
and U5491 (N_5491,N_5093,N_4929);
xor U5492 (N_5492,N_4669,N_4630);
xor U5493 (N_5493,N_4962,N_5025);
nand U5494 (N_5494,N_5235,N_4966);
or U5495 (N_5495,N_4787,N_5087);
and U5496 (N_5496,N_4868,N_5197);
and U5497 (N_5497,N_5151,N_5234);
xnor U5498 (N_5498,N_4660,N_5045);
nor U5499 (N_5499,N_4769,N_5133);
nor U5500 (N_5500,N_5022,N_5238);
and U5501 (N_5501,N_4726,N_4548);
xnor U5502 (N_5502,N_5214,N_4891);
and U5503 (N_5503,N_5050,N_4557);
nand U5504 (N_5504,N_5052,N_4909);
nor U5505 (N_5505,N_4560,N_4804);
and U5506 (N_5506,N_5036,N_4699);
or U5507 (N_5507,N_4531,N_4596);
nor U5508 (N_5508,N_4799,N_5164);
xor U5509 (N_5509,N_5156,N_4759);
xnor U5510 (N_5510,N_4971,N_4903);
xnor U5511 (N_5511,N_4846,N_4516);
or U5512 (N_5512,N_4952,N_4701);
or U5513 (N_5513,N_4673,N_5191);
xnor U5514 (N_5514,N_5112,N_4817);
nor U5515 (N_5515,N_4602,N_4543);
xnor U5516 (N_5516,N_4519,N_5246);
or U5517 (N_5517,N_4986,N_5244);
or U5518 (N_5518,N_5029,N_4805);
nor U5519 (N_5519,N_4617,N_4508);
nor U5520 (N_5520,N_5245,N_4877);
xnor U5521 (N_5521,N_5008,N_4681);
xnor U5522 (N_5522,N_4975,N_5067);
and U5523 (N_5523,N_5110,N_4571);
and U5524 (N_5524,N_4934,N_4628);
nand U5525 (N_5525,N_4796,N_4714);
nor U5526 (N_5526,N_4823,N_5180);
nand U5527 (N_5527,N_4928,N_4716);
or U5528 (N_5528,N_4919,N_4960);
or U5529 (N_5529,N_4702,N_5230);
nor U5530 (N_5530,N_5207,N_4783);
and U5531 (N_5531,N_4842,N_4812);
nand U5532 (N_5532,N_5057,N_4866);
and U5533 (N_5533,N_4549,N_4613);
nor U5534 (N_5534,N_4974,N_4533);
nand U5535 (N_5535,N_4606,N_5134);
or U5536 (N_5536,N_4890,N_4935);
nand U5537 (N_5537,N_4761,N_5061);
xnor U5538 (N_5538,N_4775,N_4821);
or U5539 (N_5539,N_4696,N_5018);
and U5540 (N_5540,N_5248,N_4605);
nor U5541 (N_5541,N_4750,N_4838);
nand U5542 (N_5542,N_5215,N_4730);
nor U5543 (N_5543,N_4840,N_4906);
and U5544 (N_5544,N_4753,N_4509);
or U5545 (N_5545,N_4798,N_4766);
nor U5546 (N_5546,N_4627,N_5006);
xor U5547 (N_5547,N_4801,N_5009);
or U5548 (N_5548,N_4857,N_4910);
and U5549 (N_5549,N_5064,N_4773);
nor U5550 (N_5550,N_4901,N_4735);
or U5551 (N_5551,N_5135,N_4569);
xor U5552 (N_5552,N_4768,N_4629);
or U5553 (N_5553,N_5136,N_4676);
nand U5554 (N_5554,N_4666,N_5211);
and U5555 (N_5555,N_4945,N_4558);
xnor U5556 (N_5556,N_4780,N_5034);
nand U5557 (N_5557,N_4755,N_4704);
nor U5558 (N_5558,N_4652,N_5186);
xor U5559 (N_5559,N_4698,N_4686);
or U5560 (N_5560,N_4908,N_4672);
nor U5561 (N_5561,N_4938,N_4626);
nor U5562 (N_5562,N_4800,N_4867);
and U5563 (N_5563,N_5169,N_4839);
nand U5564 (N_5564,N_4682,N_4770);
and U5565 (N_5565,N_4871,N_4690);
xor U5566 (N_5566,N_4599,N_4991);
or U5567 (N_5567,N_4754,N_4595);
and U5568 (N_5568,N_4946,N_5088);
or U5569 (N_5569,N_4920,N_4654);
nor U5570 (N_5570,N_5056,N_4539);
or U5571 (N_5571,N_4581,N_5228);
xnor U5572 (N_5572,N_5023,N_5243);
nand U5573 (N_5573,N_5012,N_4900);
xnor U5574 (N_5574,N_4994,N_4658);
or U5575 (N_5575,N_5072,N_4717);
xnor U5576 (N_5576,N_4586,N_4887);
nor U5577 (N_5577,N_5011,N_5004);
xnor U5578 (N_5578,N_4830,N_5014);
or U5579 (N_5579,N_4725,N_5231);
and U5580 (N_5580,N_4734,N_4847);
xor U5581 (N_5581,N_4526,N_4879);
and U5582 (N_5582,N_5016,N_4592);
or U5583 (N_5583,N_4841,N_5117);
or U5584 (N_5584,N_4584,N_4510);
and U5585 (N_5585,N_4709,N_5021);
nor U5586 (N_5586,N_5127,N_4820);
nor U5587 (N_5587,N_4936,N_5148);
xor U5588 (N_5588,N_5118,N_5079);
and U5589 (N_5589,N_5030,N_5125);
or U5590 (N_5590,N_5153,N_4973);
or U5591 (N_5591,N_4926,N_5013);
nor U5592 (N_5592,N_4861,N_4776);
nor U5593 (N_5593,N_4828,N_5205);
or U5594 (N_5594,N_4578,N_4556);
nor U5595 (N_5595,N_4736,N_4532);
or U5596 (N_5596,N_4518,N_4554);
and U5597 (N_5597,N_5204,N_4719);
or U5598 (N_5598,N_4883,N_4572);
xor U5599 (N_5599,N_4958,N_5113);
xor U5600 (N_5600,N_5150,N_5027);
and U5601 (N_5601,N_4620,N_4809);
or U5602 (N_5602,N_4545,N_4504);
and U5603 (N_5603,N_4607,N_5020);
nor U5604 (N_5604,N_5137,N_4707);
nand U5605 (N_5605,N_5147,N_4512);
or U5606 (N_5606,N_5068,N_5017);
and U5607 (N_5607,N_4967,N_5184);
nand U5608 (N_5608,N_4679,N_4852);
xor U5609 (N_5609,N_4803,N_4760);
xnor U5610 (N_5610,N_4528,N_5144);
nor U5611 (N_5611,N_4634,N_5194);
xnor U5612 (N_5612,N_4998,N_4790);
and U5613 (N_5613,N_4521,N_4639);
or U5614 (N_5614,N_5116,N_4791);
nor U5615 (N_5615,N_5076,N_4527);
and U5616 (N_5616,N_4774,N_4733);
xor U5617 (N_5617,N_4638,N_4616);
nand U5618 (N_5618,N_4983,N_4603);
nor U5619 (N_5619,N_5247,N_4976);
nor U5620 (N_5620,N_4939,N_4655);
xnor U5621 (N_5621,N_4895,N_4680);
nand U5622 (N_5622,N_5242,N_4520);
nor U5623 (N_5623,N_5096,N_4925);
nor U5624 (N_5624,N_4893,N_4721);
and U5625 (N_5625,N_4973,N_5009);
nand U5626 (N_5626,N_4658,N_4694);
xor U5627 (N_5627,N_4522,N_4741);
or U5628 (N_5628,N_4589,N_5122);
xnor U5629 (N_5629,N_4547,N_4777);
nand U5630 (N_5630,N_4847,N_5004);
xor U5631 (N_5631,N_4777,N_4689);
nand U5632 (N_5632,N_5093,N_4964);
nand U5633 (N_5633,N_4878,N_4703);
nor U5634 (N_5634,N_5093,N_4858);
xor U5635 (N_5635,N_4652,N_4551);
xor U5636 (N_5636,N_4554,N_5203);
and U5637 (N_5637,N_4782,N_4717);
nand U5638 (N_5638,N_5042,N_4891);
nor U5639 (N_5639,N_4985,N_5156);
or U5640 (N_5640,N_5234,N_4777);
nand U5641 (N_5641,N_4552,N_5207);
nand U5642 (N_5642,N_4544,N_4864);
or U5643 (N_5643,N_4758,N_4756);
and U5644 (N_5644,N_4515,N_4974);
and U5645 (N_5645,N_5099,N_5157);
nor U5646 (N_5646,N_4920,N_5099);
xnor U5647 (N_5647,N_4896,N_4952);
nand U5648 (N_5648,N_5110,N_5069);
nand U5649 (N_5649,N_4765,N_5249);
nand U5650 (N_5650,N_4808,N_4872);
and U5651 (N_5651,N_4727,N_4778);
and U5652 (N_5652,N_4620,N_5104);
xor U5653 (N_5653,N_5219,N_4747);
and U5654 (N_5654,N_4904,N_4814);
and U5655 (N_5655,N_4514,N_4573);
or U5656 (N_5656,N_4957,N_5190);
xnor U5657 (N_5657,N_4602,N_5169);
and U5658 (N_5658,N_4746,N_4624);
or U5659 (N_5659,N_4822,N_4653);
nand U5660 (N_5660,N_5150,N_4909);
or U5661 (N_5661,N_4867,N_4786);
and U5662 (N_5662,N_4652,N_4618);
nand U5663 (N_5663,N_4771,N_5218);
nor U5664 (N_5664,N_4512,N_4925);
xnor U5665 (N_5665,N_4984,N_4752);
nor U5666 (N_5666,N_4961,N_4853);
nand U5667 (N_5667,N_5118,N_4636);
xnor U5668 (N_5668,N_5185,N_4742);
and U5669 (N_5669,N_4536,N_4736);
nand U5670 (N_5670,N_4643,N_4970);
nand U5671 (N_5671,N_4627,N_4997);
and U5672 (N_5672,N_5148,N_5140);
nor U5673 (N_5673,N_4827,N_4988);
xnor U5674 (N_5674,N_4508,N_5082);
or U5675 (N_5675,N_4843,N_4522);
nor U5676 (N_5676,N_5080,N_4590);
and U5677 (N_5677,N_4961,N_4804);
nand U5678 (N_5678,N_5148,N_4783);
and U5679 (N_5679,N_4579,N_4715);
xnor U5680 (N_5680,N_5091,N_4532);
xor U5681 (N_5681,N_5201,N_5072);
and U5682 (N_5682,N_5026,N_5051);
or U5683 (N_5683,N_4890,N_5009);
nand U5684 (N_5684,N_5080,N_5243);
and U5685 (N_5685,N_4736,N_5027);
nand U5686 (N_5686,N_4754,N_4789);
nor U5687 (N_5687,N_4836,N_4769);
xor U5688 (N_5688,N_5130,N_4599);
and U5689 (N_5689,N_4838,N_5006);
nor U5690 (N_5690,N_4864,N_4724);
xor U5691 (N_5691,N_4690,N_4547);
nor U5692 (N_5692,N_4865,N_4931);
nor U5693 (N_5693,N_4634,N_5000);
xnor U5694 (N_5694,N_4799,N_4693);
xnor U5695 (N_5695,N_4516,N_4805);
and U5696 (N_5696,N_4942,N_4604);
and U5697 (N_5697,N_5073,N_4606);
xnor U5698 (N_5698,N_4873,N_4646);
nor U5699 (N_5699,N_4777,N_5025);
nor U5700 (N_5700,N_5132,N_5065);
nand U5701 (N_5701,N_5073,N_5188);
or U5702 (N_5702,N_5026,N_4749);
nand U5703 (N_5703,N_5008,N_5001);
and U5704 (N_5704,N_5236,N_5031);
and U5705 (N_5705,N_4972,N_5064);
xor U5706 (N_5706,N_4839,N_5138);
or U5707 (N_5707,N_4595,N_4809);
and U5708 (N_5708,N_4770,N_5056);
and U5709 (N_5709,N_5038,N_5208);
or U5710 (N_5710,N_4759,N_4767);
and U5711 (N_5711,N_4852,N_4524);
nand U5712 (N_5712,N_4760,N_4816);
nor U5713 (N_5713,N_4675,N_4506);
xnor U5714 (N_5714,N_4806,N_4748);
and U5715 (N_5715,N_4908,N_5115);
xor U5716 (N_5716,N_4537,N_5041);
and U5717 (N_5717,N_4731,N_4969);
nor U5718 (N_5718,N_4631,N_4855);
and U5719 (N_5719,N_5246,N_4617);
nand U5720 (N_5720,N_5116,N_4738);
and U5721 (N_5721,N_4587,N_5249);
nand U5722 (N_5722,N_4932,N_4707);
nand U5723 (N_5723,N_4816,N_4978);
and U5724 (N_5724,N_4915,N_4722);
nor U5725 (N_5725,N_4992,N_4801);
or U5726 (N_5726,N_4601,N_4511);
nand U5727 (N_5727,N_4979,N_5249);
nor U5728 (N_5728,N_5217,N_4825);
nand U5729 (N_5729,N_4853,N_4802);
nand U5730 (N_5730,N_5168,N_5069);
nand U5731 (N_5731,N_4523,N_5240);
xnor U5732 (N_5732,N_4758,N_4924);
nand U5733 (N_5733,N_4916,N_5107);
and U5734 (N_5734,N_5040,N_5027);
or U5735 (N_5735,N_4719,N_5170);
and U5736 (N_5736,N_4512,N_4665);
or U5737 (N_5737,N_5249,N_5016);
or U5738 (N_5738,N_5000,N_4615);
nand U5739 (N_5739,N_4634,N_5244);
and U5740 (N_5740,N_4970,N_4590);
or U5741 (N_5741,N_5202,N_5026);
nor U5742 (N_5742,N_4972,N_5169);
nand U5743 (N_5743,N_4883,N_5239);
and U5744 (N_5744,N_4598,N_5172);
nor U5745 (N_5745,N_4832,N_4976);
nor U5746 (N_5746,N_5058,N_4713);
nor U5747 (N_5747,N_4952,N_5074);
nand U5748 (N_5748,N_4756,N_5171);
nand U5749 (N_5749,N_5011,N_4927);
and U5750 (N_5750,N_5072,N_4565);
xnor U5751 (N_5751,N_4757,N_4775);
nand U5752 (N_5752,N_4716,N_4509);
nor U5753 (N_5753,N_5035,N_4698);
nor U5754 (N_5754,N_5047,N_4747);
or U5755 (N_5755,N_5018,N_5042);
nand U5756 (N_5756,N_5045,N_5245);
xor U5757 (N_5757,N_4770,N_5079);
nor U5758 (N_5758,N_4963,N_5024);
xor U5759 (N_5759,N_5088,N_4896);
nor U5760 (N_5760,N_4660,N_4670);
nor U5761 (N_5761,N_4782,N_5058);
nand U5762 (N_5762,N_4837,N_4835);
xnor U5763 (N_5763,N_5056,N_5044);
and U5764 (N_5764,N_4812,N_4555);
or U5765 (N_5765,N_4514,N_5138);
or U5766 (N_5766,N_4681,N_4659);
or U5767 (N_5767,N_4690,N_4511);
xnor U5768 (N_5768,N_5188,N_4943);
nand U5769 (N_5769,N_4856,N_5028);
or U5770 (N_5770,N_4514,N_4977);
and U5771 (N_5771,N_4501,N_5193);
xor U5772 (N_5772,N_5027,N_4704);
or U5773 (N_5773,N_5115,N_5155);
xor U5774 (N_5774,N_4526,N_4613);
xor U5775 (N_5775,N_5017,N_4931);
and U5776 (N_5776,N_5159,N_5017);
or U5777 (N_5777,N_4794,N_5067);
or U5778 (N_5778,N_5212,N_4874);
or U5779 (N_5779,N_4899,N_4822);
nand U5780 (N_5780,N_4626,N_5091);
nor U5781 (N_5781,N_5002,N_4995);
nand U5782 (N_5782,N_5117,N_5236);
and U5783 (N_5783,N_4849,N_4784);
nand U5784 (N_5784,N_4901,N_4701);
nand U5785 (N_5785,N_4813,N_4684);
or U5786 (N_5786,N_4539,N_5083);
nor U5787 (N_5787,N_5159,N_5139);
and U5788 (N_5788,N_5158,N_4550);
nor U5789 (N_5789,N_4726,N_5206);
xnor U5790 (N_5790,N_4633,N_4813);
and U5791 (N_5791,N_5203,N_4571);
xor U5792 (N_5792,N_5119,N_4596);
nand U5793 (N_5793,N_5166,N_4537);
nand U5794 (N_5794,N_4770,N_4941);
nand U5795 (N_5795,N_4882,N_5051);
or U5796 (N_5796,N_4660,N_4900);
nor U5797 (N_5797,N_4883,N_4560);
or U5798 (N_5798,N_4750,N_4526);
or U5799 (N_5799,N_5239,N_5095);
nand U5800 (N_5800,N_4785,N_5096);
xnor U5801 (N_5801,N_5125,N_4956);
xor U5802 (N_5802,N_5214,N_4590);
or U5803 (N_5803,N_4538,N_4944);
nand U5804 (N_5804,N_5129,N_4986);
and U5805 (N_5805,N_5206,N_4999);
xor U5806 (N_5806,N_4680,N_4559);
and U5807 (N_5807,N_4873,N_5051);
nand U5808 (N_5808,N_5179,N_5089);
nor U5809 (N_5809,N_5179,N_5068);
nor U5810 (N_5810,N_4989,N_4815);
and U5811 (N_5811,N_4944,N_4572);
or U5812 (N_5812,N_4772,N_4636);
and U5813 (N_5813,N_5198,N_4704);
or U5814 (N_5814,N_5245,N_4897);
or U5815 (N_5815,N_4884,N_5086);
nand U5816 (N_5816,N_5116,N_4548);
xnor U5817 (N_5817,N_4635,N_4647);
nand U5818 (N_5818,N_5027,N_4956);
nand U5819 (N_5819,N_4721,N_5103);
xnor U5820 (N_5820,N_5229,N_4539);
nor U5821 (N_5821,N_4606,N_4897);
xor U5822 (N_5822,N_4887,N_4800);
nor U5823 (N_5823,N_4510,N_5125);
and U5824 (N_5824,N_5123,N_4648);
nand U5825 (N_5825,N_5094,N_4818);
and U5826 (N_5826,N_4991,N_4520);
or U5827 (N_5827,N_5010,N_4662);
nor U5828 (N_5828,N_5160,N_4511);
and U5829 (N_5829,N_5107,N_4958);
and U5830 (N_5830,N_4675,N_4898);
or U5831 (N_5831,N_5243,N_5019);
and U5832 (N_5832,N_4649,N_5038);
or U5833 (N_5833,N_4571,N_4637);
or U5834 (N_5834,N_4519,N_5186);
or U5835 (N_5835,N_5150,N_5163);
nor U5836 (N_5836,N_4931,N_4733);
nor U5837 (N_5837,N_5091,N_5023);
nor U5838 (N_5838,N_5147,N_4992);
nor U5839 (N_5839,N_4644,N_4835);
and U5840 (N_5840,N_5042,N_4797);
or U5841 (N_5841,N_5228,N_5211);
xnor U5842 (N_5842,N_4760,N_4882);
xor U5843 (N_5843,N_5012,N_4739);
nor U5844 (N_5844,N_5038,N_4759);
and U5845 (N_5845,N_4794,N_5047);
nor U5846 (N_5846,N_4635,N_4778);
or U5847 (N_5847,N_4679,N_4980);
nand U5848 (N_5848,N_5067,N_4664);
and U5849 (N_5849,N_4834,N_5111);
or U5850 (N_5850,N_4785,N_5032);
and U5851 (N_5851,N_5061,N_4849);
and U5852 (N_5852,N_5106,N_5022);
nand U5853 (N_5853,N_4552,N_5087);
xor U5854 (N_5854,N_4981,N_4577);
xnor U5855 (N_5855,N_5178,N_4946);
xor U5856 (N_5856,N_5189,N_4828);
or U5857 (N_5857,N_5065,N_5064);
and U5858 (N_5858,N_4636,N_4922);
and U5859 (N_5859,N_5086,N_4532);
nor U5860 (N_5860,N_4990,N_5111);
nor U5861 (N_5861,N_4725,N_4947);
xor U5862 (N_5862,N_5101,N_4666);
xnor U5863 (N_5863,N_4896,N_5027);
or U5864 (N_5864,N_5127,N_4909);
nor U5865 (N_5865,N_4814,N_4936);
and U5866 (N_5866,N_4574,N_4549);
xnor U5867 (N_5867,N_4690,N_4512);
nand U5868 (N_5868,N_4961,N_5137);
nor U5869 (N_5869,N_4679,N_4813);
xor U5870 (N_5870,N_4634,N_4933);
or U5871 (N_5871,N_4626,N_5076);
nor U5872 (N_5872,N_5109,N_4540);
nand U5873 (N_5873,N_5067,N_5175);
or U5874 (N_5874,N_5191,N_4730);
xor U5875 (N_5875,N_4568,N_5225);
and U5876 (N_5876,N_5163,N_4718);
or U5877 (N_5877,N_4905,N_4632);
xor U5878 (N_5878,N_5026,N_4992);
nand U5879 (N_5879,N_4721,N_4758);
and U5880 (N_5880,N_4804,N_5143);
nand U5881 (N_5881,N_4592,N_4855);
or U5882 (N_5882,N_4503,N_4542);
or U5883 (N_5883,N_4761,N_5032);
and U5884 (N_5884,N_4585,N_5126);
xor U5885 (N_5885,N_4560,N_4532);
xor U5886 (N_5886,N_4793,N_4987);
xnor U5887 (N_5887,N_4934,N_4640);
nand U5888 (N_5888,N_4558,N_4609);
xnor U5889 (N_5889,N_4716,N_4505);
xor U5890 (N_5890,N_4557,N_4587);
nand U5891 (N_5891,N_5060,N_4671);
xnor U5892 (N_5892,N_4627,N_5111);
nor U5893 (N_5893,N_4525,N_4561);
and U5894 (N_5894,N_4778,N_5084);
nor U5895 (N_5895,N_4843,N_5017);
nand U5896 (N_5896,N_4918,N_5170);
nand U5897 (N_5897,N_5152,N_4905);
nor U5898 (N_5898,N_4975,N_4722);
and U5899 (N_5899,N_5045,N_4762);
xor U5900 (N_5900,N_4875,N_5178);
and U5901 (N_5901,N_5091,N_5201);
nand U5902 (N_5902,N_4635,N_4539);
or U5903 (N_5903,N_5033,N_4730);
or U5904 (N_5904,N_4799,N_5247);
or U5905 (N_5905,N_5031,N_4652);
or U5906 (N_5906,N_4953,N_5173);
or U5907 (N_5907,N_4778,N_5231);
nand U5908 (N_5908,N_4786,N_4616);
nor U5909 (N_5909,N_5226,N_4856);
or U5910 (N_5910,N_4791,N_5036);
or U5911 (N_5911,N_4757,N_4851);
nor U5912 (N_5912,N_5100,N_4577);
nand U5913 (N_5913,N_5202,N_4609);
or U5914 (N_5914,N_5120,N_5116);
nor U5915 (N_5915,N_5182,N_5104);
nand U5916 (N_5916,N_4829,N_4549);
and U5917 (N_5917,N_5242,N_4781);
or U5918 (N_5918,N_4592,N_4946);
or U5919 (N_5919,N_4961,N_4812);
nand U5920 (N_5920,N_4826,N_5075);
nand U5921 (N_5921,N_4899,N_4579);
or U5922 (N_5922,N_4827,N_4820);
xor U5923 (N_5923,N_4845,N_4989);
or U5924 (N_5924,N_4739,N_5103);
nand U5925 (N_5925,N_5029,N_4909);
xnor U5926 (N_5926,N_4527,N_4938);
nor U5927 (N_5927,N_4649,N_4607);
and U5928 (N_5928,N_5022,N_5143);
xor U5929 (N_5929,N_4870,N_5223);
and U5930 (N_5930,N_5044,N_4529);
or U5931 (N_5931,N_5210,N_4544);
nor U5932 (N_5932,N_4906,N_4521);
xnor U5933 (N_5933,N_4862,N_4709);
or U5934 (N_5934,N_4688,N_4548);
and U5935 (N_5935,N_5101,N_5114);
or U5936 (N_5936,N_5030,N_4936);
nand U5937 (N_5937,N_4956,N_4635);
xnor U5938 (N_5938,N_5104,N_4712);
and U5939 (N_5939,N_4788,N_4876);
or U5940 (N_5940,N_5077,N_4541);
and U5941 (N_5941,N_5091,N_4777);
or U5942 (N_5942,N_5175,N_5205);
nand U5943 (N_5943,N_5152,N_4660);
nor U5944 (N_5944,N_4930,N_5236);
or U5945 (N_5945,N_5054,N_5126);
or U5946 (N_5946,N_5135,N_5211);
and U5947 (N_5947,N_4541,N_5168);
nand U5948 (N_5948,N_4983,N_4631);
nor U5949 (N_5949,N_4883,N_5057);
xor U5950 (N_5950,N_5038,N_4978);
or U5951 (N_5951,N_4504,N_5076);
and U5952 (N_5952,N_4773,N_4799);
xor U5953 (N_5953,N_4709,N_4540);
xnor U5954 (N_5954,N_4635,N_4918);
nor U5955 (N_5955,N_4951,N_4666);
nand U5956 (N_5956,N_4517,N_5204);
nand U5957 (N_5957,N_4800,N_4972);
nand U5958 (N_5958,N_5220,N_5163);
nor U5959 (N_5959,N_4566,N_4992);
or U5960 (N_5960,N_4981,N_4771);
xor U5961 (N_5961,N_4748,N_5078);
and U5962 (N_5962,N_4641,N_4567);
xnor U5963 (N_5963,N_5227,N_4521);
nand U5964 (N_5964,N_5249,N_5076);
xnor U5965 (N_5965,N_4615,N_5198);
nor U5966 (N_5966,N_5210,N_4909);
nand U5967 (N_5967,N_4762,N_4537);
xnor U5968 (N_5968,N_4671,N_5066);
xnor U5969 (N_5969,N_4719,N_4811);
xor U5970 (N_5970,N_5179,N_4893);
nor U5971 (N_5971,N_4560,N_4756);
and U5972 (N_5972,N_4711,N_4714);
or U5973 (N_5973,N_5150,N_4640);
nor U5974 (N_5974,N_5129,N_5163);
or U5975 (N_5975,N_4625,N_4580);
xor U5976 (N_5976,N_5012,N_5058);
and U5977 (N_5977,N_4870,N_4641);
xnor U5978 (N_5978,N_4538,N_4911);
and U5979 (N_5979,N_4616,N_4811);
nor U5980 (N_5980,N_4937,N_5171);
xnor U5981 (N_5981,N_5212,N_4895);
xor U5982 (N_5982,N_5195,N_4763);
and U5983 (N_5983,N_5036,N_4606);
or U5984 (N_5984,N_4999,N_4967);
nand U5985 (N_5985,N_5182,N_4811);
nand U5986 (N_5986,N_4914,N_4709);
nand U5987 (N_5987,N_4584,N_4566);
xor U5988 (N_5988,N_4539,N_4744);
or U5989 (N_5989,N_4552,N_4582);
nor U5990 (N_5990,N_4909,N_4829);
or U5991 (N_5991,N_5141,N_4682);
nand U5992 (N_5992,N_4500,N_5213);
nand U5993 (N_5993,N_4501,N_4839);
xnor U5994 (N_5994,N_5124,N_5022);
and U5995 (N_5995,N_4908,N_4834);
nand U5996 (N_5996,N_4941,N_4877);
nand U5997 (N_5997,N_4904,N_4753);
nor U5998 (N_5998,N_4541,N_4657);
nor U5999 (N_5999,N_4814,N_5106);
and U6000 (N_6000,N_5350,N_5573);
nand U6001 (N_6001,N_5799,N_5561);
and U6002 (N_6002,N_5272,N_5914);
and U6003 (N_6003,N_5655,N_5433);
or U6004 (N_6004,N_5834,N_5641);
nor U6005 (N_6005,N_5690,N_5780);
xor U6006 (N_6006,N_5625,N_5736);
nor U6007 (N_6007,N_5367,N_5552);
nand U6008 (N_6008,N_5339,N_5730);
or U6009 (N_6009,N_5623,N_5802);
or U6010 (N_6010,N_5444,N_5527);
xor U6011 (N_6011,N_5772,N_5855);
nand U6012 (N_6012,N_5825,N_5266);
nor U6013 (N_6013,N_5335,N_5828);
or U6014 (N_6014,N_5943,N_5845);
nor U6015 (N_6015,N_5995,N_5742);
nor U6016 (N_6016,N_5747,N_5530);
or U6017 (N_6017,N_5949,N_5313);
or U6018 (N_6018,N_5725,N_5422);
nor U6019 (N_6019,N_5559,N_5776);
or U6020 (N_6020,N_5554,N_5865);
nand U6021 (N_6021,N_5654,N_5715);
nor U6022 (N_6022,N_5340,N_5890);
nand U6023 (N_6023,N_5366,N_5569);
or U6024 (N_6024,N_5806,N_5465);
and U6025 (N_6025,N_5735,N_5851);
nor U6026 (N_6026,N_5476,N_5485);
nand U6027 (N_6027,N_5797,N_5817);
nand U6028 (N_6028,N_5646,N_5885);
nor U6029 (N_6029,N_5666,N_5628);
and U6030 (N_6030,N_5721,N_5436);
nor U6031 (N_6031,N_5457,N_5892);
and U6032 (N_6032,N_5270,N_5349);
or U6033 (N_6033,N_5674,N_5374);
and U6034 (N_6034,N_5363,N_5344);
nand U6035 (N_6035,N_5526,N_5603);
and U6036 (N_6036,N_5588,N_5846);
or U6037 (N_6037,N_5460,N_5399);
nor U6038 (N_6038,N_5508,N_5777);
and U6039 (N_6039,N_5307,N_5861);
nand U6040 (N_6040,N_5522,N_5440);
nand U6041 (N_6041,N_5420,N_5556);
or U6042 (N_6042,N_5380,N_5788);
and U6043 (N_6043,N_5587,N_5970);
and U6044 (N_6044,N_5958,N_5517);
xnor U6045 (N_6045,N_5262,N_5540);
nor U6046 (N_6046,N_5271,N_5868);
nor U6047 (N_6047,N_5787,N_5841);
xor U6048 (N_6048,N_5394,N_5647);
nor U6049 (N_6049,N_5487,N_5660);
or U6050 (N_6050,N_5659,N_5296);
and U6051 (N_6051,N_5823,N_5796);
xnor U6052 (N_6052,N_5734,N_5827);
nand U6053 (N_6053,N_5922,N_5585);
nand U6054 (N_6054,N_5303,N_5677);
nor U6055 (N_6055,N_5935,N_5594);
xor U6056 (N_6056,N_5698,N_5626);
nand U6057 (N_6057,N_5605,N_5467);
nor U6058 (N_6058,N_5604,N_5591);
or U6059 (N_6059,N_5979,N_5863);
xnor U6060 (N_6060,N_5878,N_5864);
xor U6061 (N_6061,N_5386,N_5783);
or U6062 (N_6062,N_5687,N_5983);
or U6063 (N_6063,N_5830,N_5443);
or U6064 (N_6064,N_5456,N_5739);
nand U6065 (N_6065,N_5453,N_5720);
xor U6066 (N_6066,N_5620,N_5390);
and U6067 (N_6067,N_5314,N_5793);
xnor U6068 (N_6068,N_5547,N_5657);
and U6069 (N_6069,N_5592,N_5835);
xnor U6070 (N_6070,N_5961,N_5437);
xor U6071 (N_6071,N_5458,N_5997);
and U6072 (N_6072,N_5651,N_5500);
nand U6073 (N_6073,N_5297,N_5718);
nand U6074 (N_6074,N_5558,N_5385);
nand U6075 (N_6075,N_5857,N_5901);
xor U6076 (N_6076,N_5482,N_5921);
xnor U6077 (N_6077,N_5820,N_5534);
xor U6078 (N_6078,N_5541,N_5496);
nand U6079 (N_6079,N_5630,N_5839);
xor U6080 (N_6080,N_5814,N_5521);
nand U6081 (N_6081,N_5880,N_5583);
nor U6082 (N_6082,N_5732,N_5275);
nor U6083 (N_6083,N_5932,N_5359);
nor U6084 (N_6084,N_5737,N_5751);
xnor U6085 (N_6085,N_5905,N_5408);
xnor U6086 (N_6086,N_5993,N_5778);
and U6087 (N_6087,N_5765,N_5904);
nand U6088 (N_6088,N_5469,N_5356);
nor U6089 (N_6089,N_5947,N_5792);
nor U6090 (N_6090,N_5325,N_5273);
or U6091 (N_6091,N_5658,N_5774);
or U6092 (N_6092,N_5329,N_5381);
or U6093 (N_6093,N_5609,N_5782);
xor U6094 (N_6094,N_5639,N_5608);
nor U6095 (N_6095,N_5531,N_5462);
nor U6096 (N_6096,N_5371,N_5746);
nor U6097 (N_6097,N_5909,N_5405);
nand U6098 (N_6098,N_5689,N_5286);
nor U6099 (N_6099,N_5752,N_5749);
or U6100 (N_6100,N_5757,N_5634);
and U6101 (N_6101,N_5631,N_5343);
nor U6102 (N_6102,N_5299,N_5582);
or U6103 (N_6103,N_5840,N_5451);
nand U6104 (N_6104,N_5669,N_5254);
nor U6105 (N_6105,N_5251,N_5406);
xnor U6106 (N_6106,N_5728,N_5692);
nor U6107 (N_6107,N_5294,N_5425);
nand U6108 (N_6108,N_5267,N_5786);
xor U6109 (N_6109,N_5738,N_5570);
and U6110 (N_6110,N_5445,N_5320);
and U6111 (N_6111,N_5744,N_5317);
nor U6112 (N_6112,N_5599,N_5686);
or U6113 (N_6113,N_5847,N_5719);
and U6114 (N_6114,N_5529,N_5638);
nor U6115 (N_6115,N_5395,N_5428);
nand U6116 (N_6116,N_5672,N_5581);
nand U6117 (N_6117,N_5763,N_5859);
or U6118 (N_6118,N_5986,N_5941);
nor U6119 (N_6119,N_5563,N_5895);
nand U6120 (N_6120,N_5870,N_5546);
or U6121 (N_6121,N_5423,N_5471);
nand U6122 (N_6122,N_5695,N_5759);
nand U6123 (N_6123,N_5333,N_5956);
nand U6124 (N_6124,N_5337,N_5649);
and U6125 (N_6125,N_5486,N_5795);
nor U6126 (N_6126,N_5279,N_5894);
nor U6127 (N_6127,N_5982,N_5421);
nor U6128 (N_6128,N_5580,N_5758);
xor U6129 (N_6129,N_5850,N_5480);
or U6130 (N_6130,N_5537,N_5601);
or U6131 (N_6131,N_5938,N_5283);
or U6132 (N_6132,N_5448,N_5256);
nor U6133 (N_6133,N_5934,N_5391);
xnor U6134 (N_6134,N_5353,N_5998);
or U6135 (N_6135,N_5811,N_5700);
xnor U6136 (N_6136,N_5483,N_5969);
xor U6137 (N_6137,N_5665,N_5576);
or U6138 (N_6138,N_5409,N_5586);
or U6139 (N_6139,N_5532,N_5617);
xor U6140 (N_6140,N_5866,N_5498);
or U6141 (N_6141,N_5449,N_5516);
nor U6142 (N_6142,N_5510,N_5877);
xnor U6143 (N_6143,N_5533,N_5931);
or U6144 (N_6144,N_5775,N_5791);
nand U6145 (N_6145,N_5853,N_5673);
nand U6146 (N_6146,N_5618,N_5964);
or U6147 (N_6147,N_5790,N_5629);
and U6148 (N_6148,N_5745,N_5753);
nand U6149 (N_6149,N_5284,N_5614);
xor U6150 (N_6150,N_5560,N_5447);
and U6151 (N_6151,N_5287,N_5568);
nor U6152 (N_6152,N_5397,N_5567);
nor U6153 (N_6153,N_5536,N_5475);
xor U6154 (N_6154,N_5808,N_5724);
xnor U6155 (N_6155,N_5278,N_5450);
xnor U6156 (N_6156,N_5341,N_5761);
nor U6157 (N_6157,N_5375,N_5731);
or U6158 (N_6158,N_5762,N_5872);
or U6159 (N_6159,N_5807,N_5729);
and U6160 (N_6160,N_5939,N_5966);
nor U6161 (N_6161,N_5685,N_5973);
xnor U6162 (N_6162,N_5255,N_5972);
or U6163 (N_6163,N_5613,N_5891);
xor U6164 (N_6164,N_5810,N_5675);
xor U6165 (N_6165,N_5318,N_5676);
and U6166 (N_6166,N_5948,N_5703);
or U6167 (N_6167,N_5883,N_5670);
or U6168 (N_6168,N_5253,N_5978);
and U6169 (N_6169,N_5364,N_5985);
and U6170 (N_6170,N_5771,N_5477);
or U6171 (N_6171,N_5412,N_5327);
nand U6172 (N_6172,N_5926,N_5881);
and U6173 (N_6173,N_5463,N_5388);
or U6174 (N_6174,N_5597,N_5726);
and U6175 (N_6175,N_5338,N_5438);
xnor U6176 (N_6176,N_5813,N_5678);
or U6177 (N_6177,N_5991,N_5499);
nor U6178 (N_6178,N_5937,N_5306);
xor U6179 (N_6179,N_5512,N_5252);
or U6180 (N_6180,N_5488,N_5379);
nor U6181 (N_6181,N_5497,N_5418);
or U6182 (N_6182,N_5971,N_5697);
and U6183 (N_6183,N_5474,N_5930);
xnor U6184 (N_6184,N_5856,N_5953);
nand U6185 (N_6185,N_5369,N_5387);
or U6186 (N_6186,N_5622,N_5691);
xor U6187 (N_6187,N_5308,N_5923);
nand U6188 (N_6188,N_5976,N_5351);
or U6189 (N_6189,N_5945,N_5555);
or U6190 (N_6190,N_5289,N_5528);
and U6191 (N_6191,N_5564,N_5781);
nor U6192 (N_6192,N_5815,N_5574);
or U6193 (N_6193,N_5332,N_5992);
nor U6194 (N_6194,N_5304,N_5345);
and U6195 (N_6195,N_5519,N_5265);
or U6196 (N_6196,N_5511,N_5382);
nand U6197 (N_6197,N_5714,N_5459);
xor U6198 (N_6198,N_5924,N_5598);
xnor U6199 (N_6199,N_5716,N_5713);
nor U6200 (N_6200,N_5331,N_5292);
and U6201 (N_6201,N_5538,N_5902);
nand U6202 (N_6202,N_5316,N_5352);
or U6203 (N_6203,N_5898,N_5838);
nor U6204 (N_6204,N_5309,N_5627);
or U6205 (N_6205,N_5800,N_5288);
or U6206 (N_6206,N_5565,N_5683);
xnor U6207 (N_6207,N_5431,N_5415);
xnor U6208 (N_6208,N_5944,N_5354);
nor U6209 (N_6209,N_5548,N_5768);
or U6210 (N_6210,N_5504,N_5404);
nand U6211 (N_6211,N_5291,N_5750);
or U6212 (N_6212,N_5518,N_5928);
nor U6213 (N_6213,N_5789,N_5884);
and U6214 (N_6214,N_5442,N_5298);
nor U6215 (N_6215,N_5392,N_5767);
nor U6216 (N_6216,N_5584,N_5430);
or U6217 (N_6217,N_5616,N_5466);
nand U6218 (N_6218,N_5826,N_5876);
nand U6219 (N_6219,N_5461,N_5645);
nand U6220 (N_6220,N_5606,N_5407);
and U6221 (N_6221,N_5416,N_5489);
xor U6222 (N_6222,N_5543,N_5503);
nor U6223 (N_6223,N_5701,N_5957);
and U6224 (N_6224,N_5667,N_5454);
nand U6225 (N_6225,N_5523,N_5871);
xnor U6226 (N_6226,N_5867,N_5577);
nand U6227 (N_6227,N_5899,N_5996);
nor U6228 (N_6228,N_5414,N_5372);
or U6229 (N_6229,N_5711,N_5727);
or U6230 (N_6230,N_5550,N_5401);
or U6231 (N_6231,N_5495,N_5968);
nand U6232 (N_6232,N_5336,N_5611);
or U6233 (N_6233,N_5684,N_5723);
or U6234 (N_6234,N_5837,N_5801);
nor U6235 (N_6235,N_5990,N_5819);
or U6236 (N_6236,N_5671,N_5439);
or U6237 (N_6237,N_5798,N_5912);
xor U6238 (N_6238,N_5854,N_5411);
xnor U6239 (N_6239,N_5693,N_5636);
nand U6240 (N_6240,N_5933,N_5346);
xnor U6241 (N_6241,N_5323,N_5927);
nor U6242 (N_6242,N_5862,N_5621);
nand U6243 (N_6243,N_5707,N_5429);
or U6244 (N_6244,N_5368,N_5410);
or U6245 (N_6245,N_5274,N_5803);
or U6246 (N_6246,N_5302,N_5756);
or U6247 (N_6247,N_5596,N_5648);
nand U6248 (N_6248,N_5980,N_5712);
and U6249 (N_6249,N_5766,N_5696);
nor U6250 (N_6250,N_5310,N_5889);
nand U6251 (N_6251,N_5984,N_5326);
xnor U6252 (N_6252,N_5590,N_5607);
and U6253 (N_6253,N_5858,N_5741);
nand U6254 (N_6254,N_5575,N_5989);
nand U6255 (N_6255,N_5920,N_5962);
or U6256 (N_6256,N_5705,N_5886);
or U6257 (N_6257,N_5571,N_5812);
or U6258 (N_6258,N_5963,N_5681);
nand U6259 (N_6259,N_5427,N_5268);
and U6260 (N_6260,N_5347,N_5328);
and U6261 (N_6261,N_5615,N_5818);
or U6262 (N_6262,N_5915,N_5929);
nor U6263 (N_6263,N_5441,N_5694);
nand U6264 (N_6264,N_5551,N_5999);
or U6265 (N_6265,N_5264,N_5276);
and U6266 (N_6266,N_5794,N_5805);
nand U6267 (N_6267,N_5258,N_5804);
or U6268 (N_6268,N_5882,N_5760);
xnor U6269 (N_6269,N_5589,N_5873);
nor U6270 (N_6270,N_5330,N_5852);
nor U6271 (N_6271,N_5769,N_5373);
and U6272 (N_6272,N_5652,N_5269);
nor U6273 (N_6273,N_5709,N_5295);
and U6274 (N_6274,N_5653,N_5663);
nor U6275 (N_6275,N_5955,N_5773);
nor U6276 (N_6276,N_5965,N_5942);
and U6277 (N_6277,N_5578,N_5925);
nand U6278 (N_6278,N_5779,N_5419);
and U6279 (N_6279,N_5950,N_5688);
and U6280 (N_6280,N_5539,N_5509);
nand U6281 (N_6281,N_5740,N_5770);
nand U6282 (N_6282,N_5301,N_5470);
xnor U6283 (N_6283,N_5897,N_5668);
nand U6284 (N_6284,N_5708,N_5893);
or U6285 (N_6285,N_5610,N_5319);
xor U6286 (N_6286,N_5321,N_5967);
nand U6287 (N_6287,N_5640,N_5393);
nand U6288 (N_6288,N_5849,N_5632);
and U6289 (N_6289,N_5887,N_5472);
xnor U6290 (N_6290,N_5661,N_5911);
nor U6291 (N_6291,N_5282,N_5468);
nor U6292 (N_6292,N_5875,N_5913);
and U6293 (N_6293,N_5959,N_5357);
or U6294 (N_6294,N_5722,N_5277);
or U6295 (N_6295,N_5975,N_5361);
xnor U6296 (N_6296,N_5507,N_5358);
nor U6297 (N_6297,N_5250,N_5842);
nor U6298 (N_6298,N_5637,N_5524);
nor U6299 (N_6299,N_5280,N_5579);
nand U6300 (N_6300,N_5383,N_5664);
nor U6301 (N_6301,N_5384,N_5908);
xnor U6302 (N_6302,N_5733,N_5916);
nor U6303 (N_6303,N_5829,N_5502);
or U6304 (N_6304,N_5822,N_5481);
nand U6305 (N_6305,N_5389,N_5505);
or U6306 (N_6306,N_5981,N_5572);
nor U6307 (N_6307,N_5553,N_5940);
xor U6308 (N_6308,N_5682,N_5900);
nor U6309 (N_6309,N_5377,N_5300);
nor U6310 (N_6310,N_5535,N_5644);
xor U6311 (N_6311,N_5951,N_5513);
and U6312 (N_6312,N_5491,N_5954);
xnor U6313 (N_6313,N_5821,N_5315);
nor U6314 (N_6314,N_5362,N_5493);
and U6315 (N_6315,N_5784,N_5748);
or U6316 (N_6316,N_5642,N_5557);
xor U6317 (N_6317,N_5525,N_5479);
or U6318 (N_6318,N_5816,N_5860);
and U6319 (N_6319,N_5305,N_5595);
and U6320 (N_6320,N_5290,N_5844);
nand U6321 (N_6321,N_5506,N_5478);
and U6322 (N_6322,N_5764,N_5324);
nand U6323 (N_6323,N_5896,N_5717);
or U6324 (N_6324,N_5635,N_5566);
nand U6325 (N_6325,N_5650,N_5473);
and U6326 (N_6326,N_5490,N_5869);
xnor U6327 (N_6327,N_5602,N_5743);
xor U6328 (N_6328,N_5365,N_5633);
and U6329 (N_6329,N_5542,N_5257);
or U6330 (N_6330,N_5600,N_5874);
or U6331 (N_6331,N_5515,N_5879);
nand U6332 (N_6332,N_5403,N_5612);
or U6333 (N_6333,N_5464,N_5263);
and U6334 (N_6334,N_5435,N_5960);
nor U6335 (N_6335,N_5987,N_5400);
nand U6336 (N_6336,N_5396,N_5848);
nor U6337 (N_6337,N_5424,N_5679);
or U6338 (N_6338,N_5699,N_5643);
xor U6339 (N_6339,N_5520,N_5376);
xor U6340 (N_6340,N_5312,N_5662);
or U6341 (N_6341,N_5903,N_5355);
nand U6342 (N_6342,N_5549,N_5494);
nand U6343 (N_6343,N_5936,N_5910);
or U6344 (N_6344,N_5917,N_5706);
nor U6345 (N_6345,N_5452,N_5260);
nor U6346 (N_6346,N_5974,N_5836);
and U6347 (N_6347,N_5833,N_5311);
nand U6348 (N_6348,N_5261,N_5432);
or U6349 (N_6349,N_5514,N_5402);
nor U6350 (N_6350,N_5370,N_5809);
xor U6351 (N_6351,N_5281,N_5624);
nand U6352 (N_6352,N_5755,N_5843);
nand U6353 (N_6353,N_5619,N_5484);
and U6354 (N_6354,N_5426,N_5710);
nand U6355 (N_6355,N_5704,N_5434);
or U6356 (N_6356,N_5501,N_5259);
nor U6357 (N_6357,N_5918,N_5446);
nand U6358 (N_6358,N_5824,N_5702);
and U6359 (N_6359,N_5946,N_5544);
or U6360 (N_6360,N_5455,N_5398);
and U6361 (N_6361,N_5988,N_5831);
and U6362 (N_6362,N_5334,N_5785);
or U6363 (N_6363,N_5952,N_5656);
or U6364 (N_6364,N_5919,N_5994);
nand U6365 (N_6365,N_5417,N_5888);
nand U6366 (N_6366,N_5906,N_5680);
nand U6367 (N_6367,N_5360,N_5593);
and U6368 (N_6368,N_5378,N_5907);
nor U6369 (N_6369,N_5754,N_5545);
or U6370 (N_6370,N_5348,N_5342);
or U6371 (N_6371,N_5285,N_5832);
xnor U6372 (N_6372,N_5413,N_5977);
xor U6373 (N_6373,N_5492,N_5293);
or U6374 (N_6374,N_5562,N_5322);
nand U6375 (N_6375,N_5281,N_5654);
xor U6376 (N_6376,N_5885,N_5998);
or U6377 (N_6377,N_5764,N_5540);
and U6378 (N_6378,N_5842,N_5426);
or U6379 (N_6379,N_5991,N_5905);
and U6380 (N_6380,N_5498,N_5547);
or U6381 (N_6381,N_5958,N_5471);
and U6382 (N_6382,N_5822,N_5642);
and U6383 (N_6383,N_5614,N_5840);
or U6384 (N_6384,N_5301,N_5493);
nor U6385 (N_6385,N_5392,N_5522);
xor U6386 (N_6386,N_5797,N_5410);
nor U6387 (N_6387,N_5857,N_5937);
and U6388 (N_6388,N_5821,N_5914);
xor U6389 (N_6389,N_5742,N_5444);
or U6390 (N_6390,N_5882,N_5641);
xor U6391 (N_6391,N_5791,N_5502);
and U6392 (N_6392,N_5740,N_5522);
and U6393 (N_6393,N_5523,N_5869);
nand U6394 (N_6394,N_5826,N_5397);
and U6395 (N_6395,N_5764,N_5717);
xnor U6396 (N_6396,N_5860,N_5298);
and U6397 (N_6397,N_5766,N_5776);
or U6398 (N_6398,N_5810,N_5263);
or U6399 (N_6399,N_5639,N_5531);
and U6400 (N_6400,N_5930,N_5968);
nand U6401 (N_6401,N_5423,N_5949);
nand U6402 (N_6402,N_5648,N_5921);
xor U6403 (N_6403,N_5324,N_5397);
nor U6404 (N_6404,N_5538,N_5370);
xor U6405 (N_6405,N_5920,N_5301);
xor U6406 (N_6406,N_5639,N_5831);
xnor U6407 (N_6407,N_5663,N_5531);
nand U6408 (N_6408,N_5477,N_5331);
and U6409 (N_6409,N_5643,N_5449);
nand U6410 (N_6410,N_5786,N_5504);
xor U6411 (N_6411,N_5906,N_5619);
nor U6412 (N_6412,N_5726,N_5651);
and U6413 (N_6413,N_5680,N_5789);
and U6414 (N_6414,N_5335,N_5839);
xnor U6415 (N_6415,N_5305,N_5447);
or U6416 (N_6416,N_5634,N_5415);
and U6417 (N_6417,N_5924,N_5468);
nand U6418 (N_6418,N_5670,N_5941);
xnor U6419 (N_6419,N_5316,N_5599);
nand U6420 (N_6420,N_5629,N_5737);
or U6421 (N_6421,N_5764,N_5794);
xnor U6422 (N_6422,N_5579,N_5731);
nand U6423 (N_6423,N_5992,N_5971);
nand U6424 (N_6424,N_5778,N_5329);
nand U6425 (N_6425,N_5946,N_5931);
nor U6426 (N_6426,N_5463,N_5629);
or U6427 (N_6427,N_5940,N_5580);
and U6428 (N_6428,N_5809,N_5374);
and U6429 (N_6429,N_5826,N_5433);
and U6430 (N_6430,N_5952,N_5433);
nor U6431 (N_6431,N_5582,N_5540);
and U6432 (N_6432,N_5975,N_5703);
and U6433 (N_6433,N_5558,N_5418);
or U6434 (N_6434,N_5932,N_5569);
nor U6435 (N_6435,N_5912,N_5476);
nand U6436 (N_6436,N_5288,N_5702);
nand U6437 (N_6437,N_5864,N_5396);
and U6438 (N_6438,N_5259,N_5323);
or U6439 (N_6439,N_5351,N_5873);
or U6440 (N_6440,N_5973,N_5406);
xor U6441 (N_6441,N_5504,N_5887);
nand U6442 (N_6442,N_5559,N_5529);
nand U6443 (N_6443,N_5343,N_5737);
and U6444 (N_6444,N_5931,N_5868);
nand U6445 (N_6445,N_5270,N_5612);
or U6446 (N_6446,N_5476,N_5467);
or U6447 (N_6447,N_5543,N_5955);
and U6448 (N_6448,N_5562,N_5747);
and U6449 (N_6449,N_5459,N_5350);
or U6450 (N_6450,N_5322,N_5872);
or U6451 (N_6451,N_5277,N_5780);
nand U6452 (N_6452,N_5900,N_5417);
or U6453 (N_6453,N_5812,N_5512);
xnor U6454 (N_6454,N_5258,N_5475);
or U6455 (N_6455,N_5648,N_5831);
nand U6456 (N_6456,N_5745,N_5689);
and U6457 (N_6457,N_5756,N_5682);
nor U6458 (N_6458,N_5273,N_5677);
nand U6459 (N_6459,N_5781,N_5447);
or U6460 (N_6460,N_5592,N_5927);
and U6461 (N_6461,N_5900,N_5528);
nand U6462 (N_6462,N_5545,N_5316);
or U6463 (N_6463,N_5303,N_5784);
nand U6464 (N_6464,N_5273,N_5664);
or U6465 (N_6465,N_5488,N_5881);
or U6466 (N_6466,N_5476,N_5738);
nor U6467 (N_6467,N_5450,N_5326);
nand U6468 (N_6468,N_5266,N_5696);
or U6469 (N_6469,N_5579,N_5970);
and U6470 (N_6470,N_5290,N_5475);
and U6471 (N_6471,N_5688,N_5787);
xor U6472 (N_6472,N_5309,N_5436);
and U6473 (N_6473,N_5732,N_5879);
and U6474 (N_6474,N_5904,N_5261);
nand U6475 (N_6475,N_5943,N_5664);
nor U6476 (N_6476,N_5916,N_5479);
xor U6477 (N_6477,N_5250,N_5551);
or U6478 (N_6478,N_5969,N_5847);
and U6479 (N_6479,N_5294,N_5908);
or U6480 (N_6480,N_5493,N_5866);
or U6481 (N_6481,N_5336,N_5346);
nand U6482 (N_6482,N_5804,N_5838);
or U6483 (N_6483,N_5592,N_5909);
nand U6484 (N_6484,N_5719,N_5854);
or U6485 (N_6485,N_5752,N_5287);
xnor U6486 (N_6486,N_5875,N_5342);
and U6487 (N_6487,N_5861,N_5680);
xor U6488 (N_6488,N_5390,N_5626);
nor U6489 (N_6489,N_5508,N_5422);
or U6490 (N_6490,N_5342,N_5675);
xor U6491 (N_6491,N_5830,N_5663);
nor U6492 (N_6492,N_5947,N_5763);
or U6493 (N_6493,N_5673,N_5847);
or U6494 (N_6494,N_5359,N_5855);
or U6495 (N_6495,N_5366,N_5422);
xnor U6496 (N_6496,N_5798,N_5871);
and U6497 (N_6497,N_5960,N_5292);
nand U6498 (N_6498,N_5694,N_5477);
nor U6499 (N_6499,N_5953,N_5464);
or U6500 (N_6500,N_5283,N_5714);
xnor U6501 (N_6501,N_5404,N_5845);
or U6502 (N_6502,N_5283,N_5835);
and U6503 (N_6503,N_5886,N_5883);
or U6504 (N_6504,N_5504,N_5574);
xnor U6505 (N_6505,N_5427,N_5604);
nand U6506 (N_6506,N_5351,N_5774);
and U6507 (N_6507,N_5972,N_5793);
xnor U6508 (N_6508,N_5487,N_5503);
nand U6509 (N_6509,N_5396,N_5516);
xnor U6510 (N_6510,N_5907,N_5290);
nor U6511 (N_6511,N_5277,N_5599);
nand U6512 (N_6512,N_5450,N_5750);
nor U6513 (N_6513,N_5822,N_5394);
nor U6514 (N_6514,N_5742,N_5271);
nand U6515 (N_6515,N_5940,N_5491);
or U6516 (N_6516,N_5420,N_5435);
and U6517 (N_6517,N_5734,N_5283);
nand U6518 (N_6518,N_5973,N_5892);
xor U6519 (N_6519,N_5620,N_5433);
nand U6520 (N_6520,N_5876,N_5948);
xor U6521 (N_6521,N_5571,N_5898);
xor U6522 (N_6522,N_5459,N_5854);
or U6523 (N_6523,N_5839,N_5657);
xor U6524 (N_6524,N_5714,N_5518);
nor U6525 (N_6525,N_5343,N_5728);
or U6526 (N_6526,N_5955,N_5905);
and U6527 (N_6527,N_5908,N_5675);
xor U6528 (N_6528,N_5287,N_5510);
nand U6529 (N_6529,N_5670,N_5352);
or U6530 (N_6530,N_5753,N_5448);
or U6531 (N_6531,N_5793,N_5718);
xor U6532 (N_6532,N_5936,N_5460);
xnor U6533 (N_6533,N_5949,N_5976);
nor U6534 (N_6534,N_5999,N_5798);
xnor U6535 (N_6535,N_5870,N_5617);
or U6536 (N_6536,N_5990,N_5569);
and U6537 (N_6537,N_5572,N_5844);
nor U6538 (N_6538,N_5485,N_5251);
nand U6539 (N_6539,N_5906,N_5769);
xor U6540 (N_6540,N_5478,N_5647);
nand U6541 (N_6541,N_5318,N_5870);
nor U6542 (N_6542,N_5475,N_5321);
nor U6543 (N_6543,N_5709,N_5925);
nand U6544 (N_6544,N_5761,N_5316);
nor U6545 (N_6545,N_5848,N_5613);
nand U6546 (N_6546,N_5572,N_5837);
and U6547 (N_6547,N_5861,N_5487);
or U6548 (N_6548,N_5288,N_5488);
xor U6549 (N_6549,N_5795,N_5641);
and U6550 (N_6550,N_5587,N_5338);
or U6551 (N_6551,N_5558,N_5390);
or U6552 (N_6552,N_5347,N_5593);
or U6553 (N_6553,N_5897,N_5585);
or U6554 (N_6554,N_5414,N_5518);
and U6555 (N_6555,N_5254,N_5986);
nand U6556 (N_6556,N_5884,N_5888);
or U6557 (N_6557,N_5852,N_5523);
or U6558 (N_6558,N_5623,N_5842);
and U6559 (N_6559,N_5276,N_5746);
nand U6560 (N_6560,N_5803,N_5759);
or U6561 (N_6561,N_5564,N_5733);
nand U6562 (N_6562,N_5375,N_5804);
nor U6563 (N_6563,N_5290,N_5723);
or U6564 (N_6564,N_5587,N_5901);
nand U6565 (N_6565,N_5542,N_5379);
nor U6566 (N_6566,N_5876,N_5843);
nand U6567 (N_6567,N_5701,N_5506);
and U6568 (N_6568,N_5626,N_5635);
xnor U6569 (N_6569,N_5794,N_5717);
nor U6570 (N_6570,N_5629,N_5337);
and U6571 (N_6571,N_5371,N_5677);
or U6572 (N_6572,N_5695,N_5501);
nor U6573 (N_6573,N_5511,N_5266);
nor U6574 (N_6574,N_5501,N_5858);
nand U6575 (N_6575,N_5942,N_5992);
nor U6576 (N_6576,N_5315,N_5290);
and U6577 (N_6577,N_5474,N_5905);
nor U6578 (N_6578,N_5539,N_5492);
nor U6579 (N_6579,N_5416,N_5340);
xnor U6580 (N_6580,N_5513,N_5465);
nor U6581 (N_6581,N_5675,N_5365);
or U6582 (N_6582,N_5303,N_5879);
and U6583 (N_6583,N_5385,N_5999);
xnor U6584 (N_6584,N_5290,N_5357);
nand U6585 (N_6585,N_5925,N_5748);
or U6586 (N_6586,N_5799,N_5685);
nand U6587 (N_6587,N_5488,N_5378);
nand U6588 (N_6588,N_5631,N_5721);
xnor U6589 (N_6589,N_5915,N_5279);
xnor U6590 (N_6590,N_5934,N_5518);
nor U6591 (N_6591,N_5317,N_5971);
nor U6592 (N_6592,N_5395,N_5252);
nor U6593 (N_6593,N_5505,N_5842);
xor U6594 (N_6594,N_5286,N_5463);
or U6595 (N_6595,N_5442,N_5925);
and U6596 (N_6596,N_5601,N_5477);
nand U6597 (N_6597,N_5828,N_5977);
and U6598 (N_6598,N_5915,N_5621);
nand U6599 (N_6599,N_5651,N_5404);
nand U6600 (N_6600,N_5342,N_5296);
nor U6601 (N_6601,N_5833,N_5981);
xor U6602 (N_6602,N_5265,N_5979);
nor U6603 (N_6603,N_5656,N_5814);
and U6604 (N_6604,N_5811,N_5871);
nor U6605 (N_6605,N_5667,N_5518);
xor U6606 (N_6606,N_5659,N_5915);
and U6607 (N_6607,N_5897,N_5445);
xnor U6608 (N_6608,N_5329,N_5695);
nand U6609 (N_6609,N_5940,N_5319);
and U6610 (N_6610,N_5269,N_5908);
or U6611 (N_6611,N_5942,N_5481);
nor U6612 (N_6612,N_5595,N_5457);
and U6613 (N_6613,N_5748,N_5629);
or U6614 (N_6614,N_5585,N_5450);
nand U6615 (N_6615,N_5442,N_5786);
nand U6616 (N_6616,N_5697,N_5273);
nand U6617 (N_6617,N_5690,N_5673);
nor U6618 (N_6618,N_5693,N_5894);
xnor U6619 (N_6619,N_5856,N_5305);
nor U6620 (N_6620,N_5408,N_5374);
and U6621 (N_6621,N_5723,N_5742);
nand U6622 (N_6622,N_5254,N_5628);
nor U6623 (N_6623,N_5335,N_5576);
and U6624 (N_6624,N_5657,N_5815);
and U6625 (N_6625,N_5608,N_5795);
and U6626 (N_6626,N_5397,N_5892);
nor U6627 (N_6627,N_5965,N_5439);
nor U6628 (N_6628,N_5911,N_5927);
xnor U6629 (N_6629,N_5813,N_5524);
xor U6630 (N_6630,N_5853,N_5605);
nor U6631 (N_6631,N_5305,N_5410);
and U6632 (N_6632,N_5990,N_5885);
nand U6633 (N_6633,N_5997,N_5840);
nand U6634 (N_6634,N_5533,N_5702);
and U6635 (N_6635,N_5529,N_5979);
and U6636 (N_6636,N_5800,N_5646);
xor U6637 (N_6637,N_5766,N_5292);
nand U6638 (N_6638,N_5997,N_5969);
nor U6639 (N_6639,N_5547,N_5497);
nand U6640 (N_6640,N_5252,N_5277);
or U6641 (N_6641,N_5304,N_5941);
nor U6642 (N_6642,N_5712,N_5527);
nand U6643 (N_6643,N_5607,N_5600);
xnor U6644 (N_6644,N_5268,N_5520);
or U6645 (N_6645,N_5918,N_5520);
xnor U6646 (N_6646,N_5404,N_5438);
nand U6647 (N_6647,N_5303,N_5884);
nor U6648 (N_6648,N_5940,N_5386);
or U6649 (N_6649,N_5967,N_5567);
or U6650 (N_6650,N_5949,N_5887);
and U6651 (N_6651,N_5472,N_5946);
nand U6652 (N_6652,N_5949,N_5893);
or U6653 (N_6653,N_5413,N_5374);
and U6654 (N_6654,N_5543,N_5962);
nand U6655 (N_6655,N_5505,N_5408);
and U6656 (N_6656,N_5520,N_5463);
and U6657 (N_6657,N_5571,N_5498);
or U6658 (N_6658,N_5531,N_5481);
nand U6659 (N_6659,N_5585,N_5497);
xor U6660 (N_6660,N_5676,N_5584);
nand U6661 (N_6661,N_5476,N_5776);
and U6662 (N_6662,N_5538,N_5629);
nand U6663 (N_6663,N_5517,N_5408);
xnor U6664 (N_6664,N_5860,N_5438);
or U6665 (N_6665,N_5941,N_5344);
or U6666 (N_6666,N_5750,N_5534);
nor U6667 (N_6667,N_5263,N_5628);
nor U6668 (N_6668,N_5491,N_5646);
and U6669 (N_6669,N_5811,N_5790);
and U6670 (N_6670,N_5480,N_5251);
and U6671 (N_6671,N_5318,N_5577);
nand U6672 (N_6672,N_5876,N_5643);
nor U6673 (N_6673,N_5406,N_5652);
nor U6674 (N_6674,N_5735,N_5897);
xnor U6675 (N_6675,N_5915,N_5261);
nor U6676 (N_6676,N_5512,N_5736);
nor U6677 (N_6677,N_5289,N_5285);
nand U6678 (N_6678,N_5864,N_5552);
xnor U6679 (N_6679,N_5513,N_5361);
nor U6680 (N_6680,N_5299,N_5518);
xor U6681 (N_6681,N_5879,N_5661);
nand U6682 (N_6682,N_5846,N_5384);
xor U6683 (N_6683,N_5355,N_5958);
and U6684 (N_6684,N_5935,N_5291);
nand U6685 (N_6685,N_5780,N_5598);
or U6686 (N_6686,N_5739,N_5876);
nor U6687 (N_6687,N_5574,N_5472);
nor U6688 (N_6688,N_5629,N_5553);
nand U6689 (N_6689,N_5875,N_5602);
nor U6690 (N_6690,N_5937,N_5961);
xor U6691 (N_6691,N_5278,N_5833);
and U6692 (N_6692,N_5759,N_5918);
nand U6693 (N_6693,N_5938,N_5320);
or U6694 (N_6694,N_5891,N_5818);
nand U6695 (N_6695,N_5761,N_5474);
nand U6696 (N_6696,N_5508,N_5527);
nor U6697 (N_6697,N_5434,N_5898);
or U6698 (N_6698,N_5473,N_5604);
or U6699 (N_6699,N_5347,N_5571);
or U6700 (N_6700,N_5329,N_5831);
nand U6701 (N_6701,N_5756,N_5726);
or U6702 (N_6702,N_5290,N_5744);
or U6703 (N_6703,N_5666,N_5459);
and U6704 (N_6704,N_5774,N_5773);
or U6705 (N_6705,N_5537,N_5270);
nor U6706 (N_6706,N_5702,N_5647);
or U6707 (N_6707,N_5369,N_5314);
or U6708 (N_6708,N_5813,N_5944);
nor U6709 (N_6709,N_5591,N_5780);
and U6710 (N_6710,N_5657,N_5387);
and U6711 (N_6711,N_5424,N_5525);
or U6712 (N_6712,N_5906,N_5440);
nor U6713 (N_6713,N_5839,N_5488);
or U6714 (N_6714,N_5808,N_5435);
and U6715 (N_6715,N_5814,N_5599);
xnor U6716 (N_6716,N_5358,N_5628);
and U6717 (N_6717,N_5747,N_5259);
nor U6718 (N_6718,N_5893,N_5855);
xnor U6719 (N_6719,N_5278,N_5395);
nand U6720 (N_6720,N_5788,N_5473);
nor U6721 (N_6721,N_5547,N_5528);
nor U6722 (N_6722,N_5867,N_5660);
or U6723 (N_6723,N_5932,N_5814);
and U6724 (N_6724,N_5592,N_5794);
or U6725 (N_6725,N_5430,N_5434);
or U6726 (N_6726,N_5506,N_5877);
nand U6727 (N_6727,N_5469,N_5911);
or U6728 (N_6728,N_5790,N_5613);
nand U6729 (N_6729,N_5545,N_5738);
nand U6730 (N_6730,N_5619,N_5857);
or U6731 (N_6731,N_5250,N_5596);
xnor U6732 (N_6732,N_5674,N_5843);
nor U6733 (N_6733,N_5980,N_5737);
nor U6734 (N_6734,N_5526,N_5718);
or U6735 (N_6735,N_5670,N_5739);
nor U6736 (N_6736,N_5856,N_5267);
nor U6737 (N_6737,N_5516,N_5844);
or U6738 (N_6738,N_5482,N_5543);
xor U6739 (N_6739,N_5736,N_5540);
nand U6740 (N_6740,N_5615,N_5871);
nor U6741 (N_6741,N_5254,N_5948);
and U6742 (N_6742,N_5795,N_5986);
or U6743 (N_6743,N_5990,N_5871);
and U6744 (N_6744,N_5287,N_5428);
nand U6745 (N_6745,N_5593,N_5530);
xor U6746 (N_6746,N_5760,N_5544);
nand U6747 (N_6747,N_5923,N_5490);
and U6748 (N_6748,N_5600,N_5596);
and U6749 (N_6749,N_5415,N_5744);
nand U6750 (N_6750,N_6051,N_6707);
nor U6751 (N_6751,N_6115,N_6147);
and U6752 (N_6752,N_6031,N_6064);
nand U6753 (N_6753,N_6069,N_6614);
nor U6754 (N_6754,N_6627,N_6387);
nand U6755 (N_6755,N_6153,N_6388);
or U6756 (N_6756,N_6083,N_6542);
and U6757 (N_6757,N_6246,N_6541);
or U6758 (N_6758,N_6181,N_6450);
or U6759 (N_6759,N_6239,N_6312);
nor U6760 (N_6760,N_6092,N_6468);
nor U6761 (N_6761,N_6566,N_6404);
or U6762 (N_6762,N_6457,N_6607);
xor U6763 (N_6763,N_6482,N_6677);
xnor U6764 (N_6764,N_6276,N_6635);
and U6765 (N_6765,N_6448,N_6271);
or U6766 (N_6766,N_6453,N_6411);
or U6767 (N_6767,N_6503,N_6304);
xnor U6768 (N_6768,N_6099,N_6412);
or U6769 (N_6769,N_6547,N_6416);
nor U6770 (N_6770,N_6152,N_6444);
and U6771 (N_6771,N_6461,N_6192);
nand U6772 (N_6772,N_6221,N_6585);
nor U6773 (N_6773,N_6403,N_6636);
nor U6774 (N_6774,N_6539,N_6743);
xnor U6775 (N_6775,N_6021,N_6420);
or U6776 (N_6776,N_6436,N_6378);
nand U6777 (N_6777,N_6218,N_6699);
nand U6778 (N_6778,N_6311,N_6748);
nor U6779 (N_6779,N_6228,N_6254);
and U6780 (N_6780,N_6201,N_6197);
xor U6781 (N_6781,N_6616,N_6645);
nor U6782 (N_6782,N_6275,N_6247);
xor U6783 (N_6783,N_6065,N_6089);
nand U6784 (N_6784,N_6537,N_6018);
xnor U6785 (N_6785,N_6252,N_6729);
nor U6786 (N_6786,N_6036,N_6113);
xor U6787 (N_6787,N_6694,N_6288);
and U6788 (N_6788,N_6718,N_6193);
nor U6789 (N_6789,N_6467,N_6269);
nor U6790 (N_6790,N_6577,N_6749);
nand U6791 (N_6791,N_6406,N_6075);
xnor U6792 (N_6792,N_6674,N_6141);
xor U6793 (N_6793,N_6574,N_6534);
nor U6794 (N_6794,N_6569,N_6356);
nor U6795 (N_6795,N_6510,N_6701);
nor U6796 (N_6796,N_6671,N_6742);
xor U6797 (N_6797,N_6415,N_6705);
xor U6798 (N_6798,N_6062,N_6626);
and U6799 (N_6799,N_6441,N_6506);
nand U6800 (N_6800,N_6291,N_6085);
and U6801 (N_6801,N_6417,N_6123);
nand U6802 (N_6802,N_6161,N_6522);
and U6803 (N_6803,N_6034,N_6205);
nor U6804 (N_6804,N_6287,N_6678);
or U6805 (N_6805,N_6187,N_6279);
xnor U6806 (N_6806,N_6560,N_6731);
nand U6807 (N_6807,N_6267,N_6054);
and U6808 (N_6808,N_6315,N_6003);
and U6809 (N_6809,N_6140,N_6172);
nor U6810 (N_6810,N_6090,N_6371);
nand U6811 (N_6811,N_6074,N_6298);
xnor U6812 (N_6812,N_6106,N_6086);
and U6813 (N_6813,N_6622,N_6556);
nand U6814 (N_6814,N_6199,N_6377);
nand U6815 (N_6815,N_6326,N_6512);
and U6816 (N_6816,N_6332,N_6084);
xor U6817 (N_6817,N_6219,N_6230);
or U6818 (N_6818,N_6102,N_6588);
and U6819 (N_6819,N_6644,N_6198);
and U6820 (N_6820,N_6047,N_6068);
nand U6821 (N_6821,N_6225,N_6394);
xor U6822 (N_6822,N_6495,N_6268);
nand U6823 (N_6823,N_6568,N_6005);
and U6824 (N_6824,N_6365,N_6306);
nand U6825 (N_6825,N_6144,N_6500);
and U6826 (N_6826,N_6263,N_6392);
and U6827 (N_6827,N_6063,N_6615);
nand U6828 (N_6828,N_6242,N_6032);
xnor U6829 (N_6829,N_6533,N_6060);
or U6830 (N_6830,N_6673,N_6628);
or U6831 (N_6831,N_6231,N_6319);
xnor U6832 (N_6832,N_6698,N_6586);
and U6833 (N_6833,N_6178,N_6447);
xnor U6834 (N_6834,N_6601,N_6372);
and U6835 (N_6835,N_6660,N_6483);
or U6836 (N_6836,N_6346,N_6672);
xnor U6837 (N_6837,N_6619,N_6196);
nor U6838 (N_6838,N_6428,N_6168);
and U6839 (N_6839,N_6736,N_6238);
xnor U6840 (N_6840,N_6719,N_6355);
and U6841 (N_6841,N_6121,N_6166);
or U6842 (N_6842,N_6374,N_6160);
and U6843 (N_6843,N_6425,N_6362);
nand U6844 (N_6844,N_6333,N_6734);
nand U6845 (N_6845,N_6427,N_6264);
xor U6846 (N_6846,N_6173,N_6592);
or U6847 (N_6847,N_6726,N_6024);
xnor U6848 (N_6848,N_6049,N_6532);
and U6849 (N_6849,N_6042,N_6020);
or U6850 (N_6850,N_6286,N_6250);
xor U6851 (N_6851,N_6019,N_6216);
nand U6852 (N_6852,N_6107,N_6243);
and U6853 (N_6853,N_6498,N_6433);
or U6854 (N_6854,N_6108,N_6570);
and U6855 (N_6855,N_6511,N_6361);
xor U6856 (N_6856,N_6475,N_6233);
and U6857 (N_6857,N_6704,N_6697);
and U6858 (N_6858,N_6662,N_6557);
nor U6859 (N_6859,N_6576,N_6001);
or U6860 (N_6860,N_6657,N_6030);
and U6861 (N_6861,N_6353,N_6605);
and U6862 (N_6862,N_6012,N_6105);
nand U6863 (N_6863,N_6190,N_6561);
or U6864 (N_6864,N_6142,N_6617);
xnor U6865 (N_6865,N_6737,N_6307);
nand U6866 (N_6866,N_6469,N_6558);
or U6867 (N_6867,N_6308,N_6708);
xnor U6868 (N_6868,N_6546,N_6352);
and U6869 (N_6869,N_6602,N_6551);
xnor U6870 (N_6870,N_6313,N_6011);
nand U6871 (N_6871,N_6421,N_6621);
xnor U6872 (N_6872,N_6184,N_6473);
nor U6873 (N_6873,N_6257,N_6497);
or U6874 (N_6874,N_6292,N_6229);
or U6875 (N_6875,N_6582,N_6329);
nand U6876 (N_6876,N_6116,N_6414);
and U6877 (N_6877,N_6408,N_6189);
nand U6878 (N_6878,N_6641,N_6055);
and U6879 (N_6879,N_6145,N_6564);
nor U6880 (N_6880,N_6139,N_6659);
xor U6881 (N_6881,N_6266,N_6251);
or U6882 (N_6882,N_6658,N_6452);
and U6883 (N_6883,N_6256,N_6203);
or U6884 (N_6884,N_6097,N_6653);
nand U6885 (N_6885,N_6432,N_6342);
or U6886 (N_6886,N_6481,N_6309);
nand U6887 (N_6887,N_6262,N_6155);
and U6888 (N_6888,N_6126,N_6014);
xor U6889 (N_6889,N_6531,N_6027);
or U6890 (N_6890,N_6245,N_6202);
nor U6891 (N_6891,N_6052,N_6563);
nand U6892 (N_6892,N_6305,N_6594);
xnor U6893 (N_6893,N_6398,N_6259);
or U6894 (N_6894,N_6290,N_6261);
nor U6895 (N_6895,N_6188,N_6150);
nand U6896 (N_6896,N_6265,N_6158);
or U6897 (N_6897,N_6302,N_6136);
or U6898 (N_6898,N_6642,N_6223);
nor U6899 (N_6899,N_6523,N_6367);
nand U6900 (N_6900,N_6480,N_6215);
and U6901 (N_6901,N_6455,N_6395);
or U6902 (N_6902,N_6217,N_6258);
nand U6903 (N_6903,N_6046,N_6285);
or U6904 (N_6904,N_6389,N_6571);
nor U6905 (N_6905,N_6488,N_6204);
nor U6906 (N_6906,N_6000,N_6670);
xnor U6907 (N_6907,N_6578,N_6747);
xor U6908 (N_6908,N_6050,N_6186);
xor U6909 (N_6909,N_6318,N_6565);
nor U6910 (N_6910,N_6584,N_6209);
xnor U6911 (N_6911,N_6338,N_6407);
and U6912 (N_6912,N_6207,N_6723);
nand U6913 (N_6913,N_6526,N_6717);
or U6914 (N_6914,N_6691,N_6351);
xnor U6915 (N_6915,N_6148,N_6667);
nand U6916 (N_6916,N_6727,N_6349);
nand U6917 (N_6917,N_6689,N_6499);
nand U6918 (N_6918,N_6345,N_6104);
xnor U6919 (N_6919,N_6714,N_6735);
nor U6920 (N_6920,N_6026,N_6151);
nor U6921 (N_6921,N_6323,N_6732);
xnor U6922 (N_6922,N_6373,N_6396);
or U6923 (N_6923,N_6112,N_6134);
nand U6924 (N_6924,N_6384,N_6098);
nor U6925 (N_6925,N_6625,N_6170);
nand U6926 (N_6926,N_6103,N_6022);
nand U6927 (N_6927,N_6476,N_6096);
xor U6928 (N_6928,N_6517,N_6439);
nand U6929 (N_6929,N_6359,N_6710);
nor U6930 (N_6930,N_6632,N_6094);
nor U6931 (N_6931,N_6039,N_6399);
nand U6932 (N_6932,N_6273,N_6516);
nand U6933 (N_6933,N_6117,N_6391);
xor U6934 (N_6934,N_6424,N_6715);
or U6935 (N_6935,N_6449,N_6331);
and U6936 (N_6936,N_6240,N_6494);
xnor U6937 (N_6937,N_6082,N_6643);
xor U6938 (N_6938,N_6536,N_6638);
nor U6939 (N_6939,N_6035,N_6131);
and U6940 (N_6940,N_6695,N_6270);
and U6941 (N_6941,N_6222,N_6344);
or U6942 (N_6942,N_6746,N_6593);
nor U6943 (N_6943,N_6525,N_6157);
or U6944 (N_6944,N_6095,N_6640);
or U6945 (N_6945,N_6070,N_6081);
xnor U6946 (N_6946,N_6502,N_6630);
or U6947 (N_6947,N_6277,N_6133);
nor U6948 (N_6948,N_6611,N_6580);
nor U6949 (N_6949,N_6528,N_6652);
or U6950 (N_6950,N_6651,N_6700);
or U6951 (N_6951,N_6281,N_6077);
xnor U6952 (N_6952,N_6490,N_6504);
xnor U6953 (N_6953,N_6101,N_6017);
xnor U6954 (N_6954,N_6744,N_6429);
nand U6955 (N_6955,N_6458,N_6325);
nor U6956 (N_6956,N_6740,N_6129);
nand U6957 (N_6957,N_6016,N_6472);
nor U6958 (N_6958,N_6232,N_6293);
or U6959 (N_6959,N_6381,N_6194);
nor U6960 (N_6960,N_6538,N_6380);
nor U6961 (N_6961,N_6210,N_6501);
or U6962 (N_6962,N_6162,N_6682);
xnor U6963 (N_6963,N_6033,N_6278);
and U6964 (N_6964,N_6587,N_6044);
nor U6965 (N_6965,N_6618,N_6071);
nand U6966 (N_6966,N_6709,N_6169);
xnor U6967 (N_6967,N_6334,N_6581);
nor U6968 (N_6968,N_6175,N_6182);
xnor U6969 (N_6969,N_6513,N_6664);
nand U6970 (N_6970,N_6200,N_6543);
nand U6971 (N_6971,N_6368,N_6048);
nor U6972 (N_6972,N_6343,N_6294);
nor U6973 (N_6973,N_6119,N_6080);
or U6974 (N_6974,N_6623,N_6088);
xor U6975 (N_6975,N_6303,N_6029);
nor U6976 (N_6976,N_6109,N_6478);
xor U6977 (N_6977,N_6053,N_6040);
xor U6978 (N_6978,N_6600,N_6023);
nor U6979 (N_6979,N_6183,N_6057);
and U6980 (N_6980,N_6317,N_6474);
nand U6981 (N_6981,N_6445,N_6419);
nand U6982 (N_6982,N_6702,N_6629);
and U6983 (N_6983,N_6548,N_6728);
nand U6984 (N_6984,N_6604,N_6341);
and U6985 (N_6985,N_6087,N_6227);
or U6986 (N_6986,N_6382,N_6529);
xor U6987 (N_6987,N_6661,N_6454);
nor U6988 (N_6988,N_6350,N_6466);
nor U6989 (N_6989,N_6540,N_6688);
nand U6990 (N_6990,N_6686,N_6634);
nor U6991 (N_6991,N_6248,N_6386);
and U6992 (N_6992,N_6214,N_6195);
xnor U6993 (N_6993,N_6375,N_6310);
nand U6994 (N_6994,N_6559,N_6426);
xor U6995 (N_6995,N_6741,N_6213);
nand U6996 (N_6996,N_6505,N_6675);
xnor U6997 (N_6997,N_6383,N_6613);
and U6998 (N_6998,N_6237,N_6493);
xor U6999 (N_6999,N_6314,N_6212);
and U7000 (N_7000,N_6519,N_6322);
nor U7001 (N_7001,N_6244,N_6620);
xnor U7002 (N_7002,N_6646,N_6509);
nand U7003 (N_7003,N_6685,N_6486);
nor U7004 (N_7004,N_6598,N_6579);
nor U7005 (N_7005,N_6738,N_6220);
or U7006 (N_7006,N_6357,N_6135);
and U7007 (N_7007,N_6535,N_6530);
nand U7008 (N_7008,N_6545,N_6612);
or U7009 (N_7009,N_6006,N_6722);
nand U7010 (N_7010,N_6280,N_6596);
nand U7011 (N_7011,N_6059,N_6226);
or U7012 (N_7012,N_6485,N_6496);
nor U7013 (N_7013,N_6120,N_6008);
and U7014 (N_7014,N_6552,N_6038);
or U7015 (N_7015,N_6324,N_6554);
nand U7016 (N_7016,N_6211,N_6339);
and U7017 (N_7017,N_6358,N_6443);
nor U7018 (N_7018,N_6236,N_6518);
nor U7019 (N_7019,N_6146,N_6297);
and U7020 (N_7020,N_6316,N_6274);
and U7021 (N_7021,N_6440,N_6484);
or U7022 (N_7022,N_6122,N_6492);
and U7023 (N_7023,N_6124,N_6597);
nor U7024 (N_7024,N_6606,N_6056);
nand U7025 (N_7025,N_6460,N_6013);
and U7026 (N_7026,N_6608,N_6347);
or U7027 (N_7027,N_6206,N_6589);
nor U7028 (N_7028,N_6028,N_6521);
or U7029 (N_7029,N_6572,N_6078);
nand U7030 (N_7030,N_6573,N_6591);
xnor U7031 (N_7031,N_6423,N_6363);
or U7032 (N_7032,N_6045,N_6009);
nor U7033 (N_7033,N_6138,N_6149);
or U7034 (N_7034,N_6418,N_6176);
xor U7035 (N_7035,N_6163,N_6300);
nand U7036 (N_7036,N_6154,N_6553);
nor U7037 (N_7037,N_6180,N_6679);
xor U7038 (N_7038,N_6002,N_6650);
and U7039 (N_7039,N_6721,N_6015);
nand U7040 (N_7040,N_6669,N_6434);
nor U7041 (N_7041,N_6520,N_6348);
nand U7042 (N_7042,N_6301,N_6224);
and U7043 (N_7043,N_6711,N_6706);
nand U7044 (N_7044,N_6402,N_6712);
or U7045 (N_7045,N_6463,N_6668);
and U7046 (N_7046,N_6666,N_6143);
nand U7047 (N_7047,N_6165,N_6253);
or U7048 (N_7048,N_6687,N_6507);
and U7049 (N_7049,N_6655,N_6110);
nor U7050 (N_7050,N_6442,N_6007);
and U7051 (N_7051,N_6745,N_6255);
nand U7052 (N_7052,N_6633,N_6451);
xnor U7053 (N_7053,N_6739,N_6730);
nand U7054 (N_7054,N_6562,N_6471);
and U7055 (N_7055,N_6130,N_6465);
and U7056 (N_7056,N_6713,N_6680);
nand U7057 (N_7057,N_6470,N_6693);
nand U7058 (N_7058,N_6164,N_6076);
xnor U7059 (N_7059,N_6438,N_6555);
nor U7060 (N_7060,N_6401,N_6295);
nor U7061 (N_7061,N_6185,N_6079);
nand U7062 (N_7062,N_6128,N_6514);
nor U7063 (N_7063,N_6366,N_6132);
nand U7064 (N_7064,N_6073,N_6456);
nand U7065 (N_7065,N_6590,N_6241);
xor U7066 (N_7066,N_6446,N_6296);
nand U7067 (N_7067,N_6393,N_6696);
and U7068 (N_7068,N_6487,N_6637);
nor U7069 (N_7069,N_6459,N_6327);
nand U7070 (N_7070,N_6025,N_6235);
or U7071 (N_7071,N_6114,N_6369);
or U7072 (N_7072,N_6336,N_6508);
nand U7073 (N_7073,N_6111,N_6370);
and U7074 (N_7074,N_6550,N_6464);
or U7075 (N_7075,N_6272,N_6058);
nand U7076 (N_7076,N_6690,N_6631);
or U7077 (N_7077,N_6527,N_6328);
or U7078 (N_7078,N_6067,N_6665);
nand U7079 (N_7079,N_6249,N_6100);
xor U7080 (N_7080,N_6400,N_6656);
and U7081 (N_7081,N_6093,N_6524);
and U7082 (N_7082,N_6639,N_6654);
nor U7083 (N_7083,N_6376,N_6390);
nand U7084 (N_7084,N_6647,N_6720);
nor U7085 (N_7085,N_6405,N_6649);
and U7086 (N_7086,N_6010,N_6191);
nand U7087 (N_7087,N_6703,N_6208);
nor U7088 (N_7088,N_6360,N_6692);
nor U7089 (N_7089,N_6610,N_6435);
xor U7090 (N_7090,N_6477,N_6066);
and U7091 (N_7091,N_6681,N_6684);
and U7092 (N_7092,N_6379,N_6489);
nor U7093 (N_7093,N_6725,N_6167);
xor U7094 (N_7094,N_6004,N_6284);
and U7095 (N_7095,N_6260,N_6125);
nand U7096 (N_7096,N_6061,N_6159);
or U7097 (N_7097,N_6676,N_6321);
or U7098 (N_7098,N_6544,N_6091);
and U7099 (N_7099,N_6072,N_6364);
or U7100 (N_7100,N_6663,N_6479);
xnor U7101 (N_7101,N_6127,N_6330);
and U7102 (N_7102,N_6724,N_6118);
nor U7103 (N_7103,N_6575,N_6289);
or U7104 (N_7104,N_6171,N_6410);
and U7105 (N_7105,N_6567,N_6549);
or U7106 (N_7106,N_6716,N_6583);
and U7107 (N_7107,N_6422,N_6599);
nand U7108 (N_7108,N_6043,N_6609);
and U7109 (N_7109,N_6179,N_6234);
nand U7110 (N_7110,N_6733,N_6431);
nor U7111 (N_7111,N_6354,N_6337);
or U7112 (N_7112,N_6603,N_6137);
nand U7113 (N_7113,N_6595,N_6156);
nand U7114 (N_7114,N_6177,N_6282);
or U7115 (N_7115,N_6683,N_6283);
or U7116 (N_7116,N_6397,N_6413);
xnor U7117 (N_7117,N_6320,N_6335);
and U7118 (N_7118,N_6299,N_6462);
nor U7119 (N_7119,N_6174,N_6437);
nor U7120 (N_7120,N_6515,N_6340);
xnor U7121 (N_7121,N_6648,N_6385);
xor U7122 (N_7122,N_6409,N_6430);
xor U7123 (N_7123,N_6624,N_6037);
and U7124 (N_7124,N_6041,N_6491);
nand U7125 (N_7125,N_6636,N_6476);
nor U7126 (N_7126,N_6567,N_6385);
or U7127 (N_7127,N_6609,N_6579);
nor U7128 (N_7128,N_6647,N_6590);
or U7129 (N_7129,N_6576,N_6375);
xnor U7130 (N_7130,N_6420,N_6351);
nand U7131 (N_7131,N_6614,N_6682);
xnor U7132 (N_7132,N_6638,N_6033);
xnor U7133 (N_7133,N_6625,N_6503);
nor U7134 (N_7134,N_6644,N_6250);
or U7135 (N_7135,N_6319,N_6738);
nand U7136 (N_7136,N_6385,N_6562);
and U7137 (N_7137,N_6703,N_6638);
or U7138 (N_7138,N_6397,N_6258);
xor U7139 (N_7139,N_6177,N_6104);
nor U7140 (N_7140,N_6216,N_6146);
nor U7141 (N_7141,N_6192,N_6421);
xor U7142 (N_7142,N_6060,N_6053);
and U7143 (N_7143,N_6481,N_6490);
or U7144 (N_7144,N_6224,N_6495);
or U7145 (N_7145,N_6404,N_6005);
xnor U7146 (N_7146,N_6130,N_6290);
or U7147 (N_7147,N_6022,N_6542);
or U7148 (N_7148,N_6177,N_6470);
xnor U7149 (N_7149,N_6520,N_6154);
and U7150 (N_7150,N_6013,N_6539);
or U7151 (N_7151,N_6384,N_6080);
and U7152 (N_7152,N_6142,N_6601);
or U7153 (N_7153,N_6194,N_6682);
nand U7154 (N_7154,N_6121,N_6397);
xnor U7155 (N_7155,N_6247,N_6729);
nor U7156 (N_7156,N_6530,N_6285);
nor U7157 (N_7157,N_6058,N_6151);
or U7158 (N_7158,N_6607,N_6203);
nand U7159 (N_7159,N_6609,N_6334);
nand U7160 (N_7160,N_6621,N_6586);
nor U7161 (N_7161,N_6602,N_6126);
nor U7162 (N_7162,N_6201,N_6614);
xor U7163 (N_7163,N_6632,N_6374);
nand U7164 (N_7164,N_6478,N_6647);
and U7165 (N_7165,N_6078,N_6161);
or U7166 (N_7166,N_6456,N_6466);
and U7167 (N_7167,N_6615,N_6716);
xor U7168 (N_7168,N_6374,N_6544);
or U7169 (N_7169,N_6494,N_6119);
and U7170 (N_7170,N_6443,N_6089);
xnor U7171 (N_7171,N_6436,N_6402);
nand U7172 (N_7172,N_6368,N_6469);
nand U7173 (N_7173,N_6357,N_6175);
nor U7174 (N_7174,N_6505,N_6027);
nor U7175 (N_7175,N_6691,N_6150);
and U7176 (N_7176,N_6205,N_6219);
xor U7177 (N_7177,N_6035,N_6409);
and U7178 (N_7178,N_6122,N_6218);
nor U7179 (N_7179,N_6212,N_6609);
xnor U7180 (N_7180,N_6622,N_6233);
and U7181 (N_7181,N_6715,N_6493);
and U7182 (N_7182,N_6529,N_6254);
xor U7183 (N_7183,N_6343,N_6267);
or U7184 (N_7184,N_6413,N_6628);
or U7185 (N_7185,N_6565,N_6600);
and U7186 (N_7186,N_6242,N_6310);
nand U7187 (N_7187,N_6704,N_6069);
nand U7188 (N_7188,N_6058,N_6285);
nor U7189 (N_7189,N_6456,N_6318);
nor U7190 (N_7190,N_6414,N_6068);
and U7191 (N_7191,N_6448,N_6346);
nand U7192 (N_7192,N_6618,N_6249);
xnor U7193 (N_7193,N_6740,N_6001);
or U7194 (N_7194,N_6337,N_6029);
xnor U7195 (N_7195,N_6025,N_6635);
xor U7196 (N_7196,N_6748,N_6160);
and U7197 (N_7197,N_6444,N_6702);
or U7198 (N_7198,N_6282,N_6446);
or U7199 (N_7199,N_6623,N_6046);
nor U7200 (N_7200,N_6381,N_6207);
nand U7201 (N_7201,N_6661,N_6335);
and U7202 (N_7202,N_6357,N_6071);
nand U7203 (N_7203,N_6110,N_6582);
and U7204 (N_7204,N_6123,N_6698);
nand U7205 (N_7205,N_6054,N_6130);
or U7206 (N_7206,N_6216,N_6600);
nor U7207 (N_7207,N_6221,N_6303);
nand U7208 (N_7208,N_6311,N_6143);
or U7209 (N_7209,N_6149,N_6290);
and U7210 (N_7210,N_6433,N_6190);
nor U7211 (N_7211,N_6102,N_6300);
or U7212 (N_7212,N_6324,N_6168);
or U7213 (N_7213,N_6033,N_6591);
and U7214 (N_7214,N_6612,N_6733);
nand U7215 (N_7215,N_6217,N_6532);
xnor U7216 (N_7216,N_6747,N_6011);
or U7217 (N_7217,N_6179,N_6542);
or U7218 (N_7218,N_6304,N_6699);
xor U7219 (N_7219,N_6715,N_6024);
nor U7220 (N_7220,N_6178,N_6464);
nand U7221 (N_7221,N_6404,N_6121);
or U7222 (N_7222,N_6111,N_6379);
nor U7223 (N_7223,N_6622,N_6673);
nand U7224 (N_7224,N_6593,N_6250);
nor U7225 (N_7225,N_6567,N_6103);
nand U7226 (N_7226,N_6163,N_6369);
nand U7227 (N_7227,N_6237,N_6265);
xnor U7228 (N_7228,N_6240,N_6233);
nor U7229 (N_7229,N_6631,N_6234);
or U7230 (N_7230,N_6281,N_6047);
xnor U7231 (N_7231,N_6295,N_6032);
and U7232 (N_7232,N_6375,N_6192);
and U7233 (N_7233,N_6064,N_6573);
xor U7234 (N_7234,N_6653,N_6276);
nor U7235 (N_7235,N_6641,N_6679);
nand U7236 (N_7236,N_6670,N_6659);
or U7237 (N_7237,N_6003,N_6316);
and U7238 (N_7238,N_6223,N_6616);
nand U7239 (N_7239,N_6310,N_6678);
or U7240 (N_7240,N_6634,N_6610);
xnor U7241 (N_7241,N_6040,N_6218);
xor U7242 (N_7242,N_6596,N_6333);
nand U7243 (N_7243,N_6098,N_6052);
nand U7244 (N_7244,N_6016,N_6720);
nand U7245 (N_7245,N_6495,N_6307);
or U7246 (N_7246,N_6735,N_6455);
or U7247 (N_7247,N_6748,N_6527);
xor U7248 (N_7248,N_6511,N_6538);
and U7249 (N_7249,N_6227,N_6335);
and U7250 (N_7250,N_6211,N_6297);
and U7251 (N_7251,N_6275,N_6613);
xnor U7252 (N_7252,N_6424,N_6262);
nand U7253 (N_7253,N_6602,N_6272);
nor U7254 (N_7254,N_6316,N_6327);
or U7255 (N_7255,N_6161,N_6441);
nand U7256 (N_7256,N_6062,N_6746);
nand U7257 (N_7257,N_6224,N_6392);
or U7258 (N_7258,N_6246,N_6010);
and U7259 (N_7259,N_6001,N_6182);
nor U7260 (N_7260,N_6303,N_6005);
and U7261 (N_7261,N_6685,N_6188);
or U7262 (N_7262,N_6203,N_6258);
and U7263 (N_7263,N_6128,N_6021);
nor U7264 (N_7264,N_6517,N_6138);
xor U7265 (N_7265,N_6184,N_6039);
xor U7266 (N_7266,N_6065,N_6389);
and U7267 (N_7267,N_6100,N_6325);
and U7268 (N_7268,N_6124,N_6184);
and U7269 (N_7269,N_6594,N_6378);
xor U7270 (N_7270,N_6229,N_6433);
xor U7271 (N_7271,N_6125,N_6695);
or U7272 (N_7272,N_6178,N_6348);
or U7273 (N_7273,N_6724,N_6644);
xnor U7274 (N_7274,N_6061,N_6200);
or U7275 (N_7275,N_6563,N_6456);
nor U7276 (N_7276,N_6609,N_6021);
xnor U7277 (N_7277,N_6572,N_6689);
nand U7278 (N_7278,N_6406,N_6399);
or U7279 (N_7279,N_6119,N_6627);
xnor U7280 (N_7280,N_6389,N_6675);
nand U7281 (N_7281,N_6339,N_6549);
or U7282 (N_7282,N_6365,N_6139);
or U7283 (N_7283,N_6608,N_6530);
or U7284 (N_7284,N_6304,N_6442);
nand U7285 (N_7285,N_6164,N_6691);
or U7286 (N_7286,N_6576,N_6687);
or U7287 (N_7287,N_6271,N_6610);
or U7288 (N_7288,N_6003,N_6354);
nor U7289 (N_7289,N_6410,N_6583);
nor U7290 (N_7290,N_6332,N_6644);
or U7291 (N_7291,N_6253,N_6520);
nor U7292 (N_7292,N_6655,N_6661);
nand U7293 (N_7293,N_6458,N_6404);
or U7294 (N_7294,N_6078,N_6132);
nor U7295 (N_7295,N_6392,N_6571);
and U7296 (N_7296,N_6046,N_6303);
nor U7297 (N_7297,N_6115,N_6248);
nand U7298 (N_7298,N_6329,N_6668);
nand U7299 (N_7299,N_6394,N_6220);
nor U7300 (N_7300,N_6245,N_6253);
and U7301 (N_7301,N_6749,N_6381);
and U7302 (N_7302,N_6351,N_6099);
nor U7303 (N_7303,N_6706,N_6635);
nand U7304 (N_7304,N_6305,N_6542);
and U7305 (N_7305,N_6567,N_6677);
nand U7306 (N_7306,N_6451,N_6736);
or U7307 (N_7307,N_6503,N_6076);
or U7308 (N_7308,N_6169,N_6437);
nor U7309 (N_7309,N_6025,N_6444);
and U7310 (N_7310,N_6161,N_6382);
and U7311 (N_7311,N_6519,N_6371);
or U7312 (N_7312,N_6011,N_6303);
and U7313 (N_7313,N_6193,N_6268);
nor U7314 (N_7314,N_6666,N_6194);
xnor U7315 (N_7315,N_6489,N_6481);
xor U7316 (N_7316,N_6711,N_6130);
xor U7317 (N_7317,N_6045,N_6328);
nand U7318 (N_7318,N_6359,N_6398);
xor U7319 (N_7319,N_6143,N_6226);
nand U7320 (N_7320,N_6354,N_6216);
nand U7321 (N_7321,N_6137,N_6706);
nor U7322 (N_7322,N_6578,N_6722);
nand U7323 (N_7323,N_6308,N_6369);
nor U7324 (N_7324,N_6738,N_6182);
nor U7325 (N_7325,N_6046,N_6453);
nand U7326 (N_7326,N_6638,N_6546);
nor U7327 (N_7327,N_6605,N_6361);
nor U7328 (N_7328,N_6485,N_6314);
or U7329 (N_7329,N_6149,N_6029);
xnor U7330 (N_7330,N_6588,N_6375);
nor U7331 (N_7331,N_6661,N_6555);
xor U7332 (N_7332,N_6345,N_6038);
xnor U7333 (N_7333,N_6269,N_6519);
nand U7334 (N_7334,N_6631,N_6657);
nand U7335 (N_7335,N_6664,N_6255);
nor U7336 (N_7336,N_6650,N_6041);
xor U7337 (N_7337,N_6020,N_6601);
nor U7338 (N_7338,N_6470,N_6372);
nor U7339 (N_7339,N_6202,N_6497);
or U7340 (N_7340,N_6585,N_6646);
or U7341 (N_7341,N_6052,N_6048);
nand U7342 (N_7342,N_6420,N_6698);
xor U7343 (N_7343,N_6551,N_6078);
or U7344 (N_7344,N_6268,N_6364);
nor U7345 (N_7345,N_6641,N_6167);
or U7346 (N_7346,N_6312,N_6049);
xnor U7347 (N_7347,N_6677,N_6681);
nand U7348 (N_7348,N_6633,N_6534);
or U7349 (N_7349,N_6507,N_6699);
xnor U7350 (N_7350,N_6298,N_6100);
nor U7351 (N_7351,N_6299,N_6150);
and U7352 (N_7352,N_6500,N_6276);
xnor U7353 (N_7353,N_6252,N_6217);
nor U7354 (N_7354,N_6038,N_6451);
nor U7355 (N_7355,N_6211,N_6675);
or U7356 (N_7356,N_6505,N_6312);
or U7357 (N_7357,N_6415,N_6429);
nor U7358 (N_7358,N_6403,N_6549);
or U7359 (N_7359,N_6619,N_6582);
nor U7360 (N_7360,N_6075,N_6236);
and U7361 (N_7361,N_6420,N_6247);
nand U7362 (N_7362,N_6049,N_6641);
xor U7363 (N_7363,N_6201,N_6207);
and U7364 (N_7364,N_6461,N_6500);
or U7365 (N_7365,N_6694,N_6170);
or U7366 (N_7366,N_6507,N_6084);
nor U7367 (N_7367,N_6370,N_6238);
or U7368 (N_7368,N_6115,N_6456);
nand U7369 (N_7369,N_6667,N_6592);
xnor U7370 (N_7370,N_6112,N_6602);
and U7371 (N_7371,N_6556,N_6277);
and U7372 (N_7372,N_6608,N_6320);
nor U7373 (N_7373,N_6406,N_6335);
xor U7374 (N_7374,N_6722,N_6400);
or U7375 (N_7375,N_6353,N_6059);
nand U7376 (N_7376,N_6665,N_6075);
nand U7377 (N_7377,N_6613,N_6600);
nor U7378 (N_7378,N_6354,N_6547);
or U7379 (N_7379,N_6336,N_6607);
nor U7380 (N_7380,N_6443,N_6457);
or U7381 (N_7381,N_6710,N_6222);
nor U7382 (N_7382,N_6448,N_6406);
nor U7383 (N_7383,N_6356,N_6359);
and U7384 (N_7384,N_6710,N_6625);
and U7385 (N_7385,N_6369,N_6538);
or U7386 (N_7386,N_6382,N_6402);
nor U7387 (N_7387,N_6555,N_6626);
xnor U7388 (N_7388,N_6408,N_6749);
or U7389 (N_7389,N_6043,N_6450);
and U7390 (N_7390,N_6173,N_6237);
nor U7391 (N_7391,N_6513,N_6024);
nand U7392 (N_7392,N_6158,N_6615);
and U7393 (N_7393,N_6607,N_6252);
nor U7394 (N_7394,N_6746,N_6657);
xnor U7395 (N_7395,N_6495,N_6181);
xnor U7396 (N_7396,N_6348,N_6717);
nand U7397 (N_7397,N_6350,N_6747);
nor U7398 (N_7398,N_6412,N_6161);
and U7399 (N_7399,N_6418,N_6143);
xor U7400 (N_7400,N_6569,N_6144);
xnor U7401 (N_7401,N_6012,N_6217);
and U7402 (N_7402,N_6316,N_6662);
nand U7403 (N_7403,N_6201,N_6665);
and U7404 (N_7404,N_6082,N_6702);
or U7405 (N_7405,N_6304,N_6471);
nand U7406 (N_7406,N_6030,N_6154);
nand U7407 (N_7407,N_6239,N_6127);
and U7408 (N_7408,N_6275,N_6013);
and U7409 (N_7409,N_6209,N_6148);
or U7410 (N_7410,N_6710,N_6262);
xor U7411 (N_7411,N_6002,N_6216);
or U7412 (N_7412,N_6130,N_6611);
or U7413 (N_7413,N_6412,N_6657);
and U7414 (N_7414,N_6264,N_6333);
and U7415 (N_7415,N_6216,N_6411);
or U7416 (N_7416,N_6258,N_6328);
xnor U7417 (N_7417,N_6196,N_6416);
nor U7418 (N_7418,N_6245,N_6179);
nand U7419 (N_7419,N_6535,N_6664);
nand U7420 (N_7420,N_6134,N_6409);
xnor U7421 (N_7421,N_6099,N_6620);
nand U7422 (N_7422,N_6085,N_6004);
nor U7423 (N_7423,N_6272,N_6525);
xnor U7424 (N_7424,N_6736,N_6293);
and U7425 (N_7425,N_6417,N_6344);
xor U7426 (N_7426,N_6627,N_6744);
xor U7427 (N_7427,N_6153,N_6315);
or U7428 (N_7428,N_6646,N_6449);
xor U7429 (N_7429,N_6564,N_6706);
and U7430 (N_7430,N_6683,N_6206);
xor U7431 (N_7431,N_6082,N_6679);
or U7432 (N_7432,N_6639,N_6056);
nand U7433 (N_7433,N_6290,N_6195);
or U7434 (N_7434,N_6386,N_6280);
nand U7435 (N_7435,N_6682,N_6698);
xnor U7436 (N_7436,N_6456,N_6622);
nand U7437 (N_7437,N_6711,N_6517);
nor U7438 (N_7438,N_6357,N_6556);
nor U7439 (N_7439,N_6231,N_6065);
xor U7440 (N_7440,N_6696,N_6636);
xnor U7441 (N_7441,N_6500,N_6641);
nand U7442 (N_7442,N_6229,N_6436);
and U7443 (N_7443,N_6355,N_6683);
nor U7444 (N_7444,N_6723,N_6390);
xor U7445 (N_7445,N_6647,N_6028);
or U7446 (N_7446,N_6215,N_6524);
nor U7447 (N_7447,N_6736,N_6067);
nor U7448 (N_7448,N_6347,N_6373);
and U7449 (N_7449,N_6081,N_6706);
and U7450 (N_7450,N_6523,N_6706);
or U7451 (N_7451,N_6606,N_6356);
nor U7452 (N_7452,N_6309,N_6405);
nand U7453 (N_7453,N_6472,N_6614);
or U7454 (N_7454,N_6255,N_6675);
nor U7455 (N_7455,N_6705,N_6294);
and U7456 (N_7456,N_6713,N_6419);
xnor U7457 (N_7457,N_6672,N_6245);
nand U7458 (N_7458,N_6234,N_6317);
or U7459 (N_7459,N_6650,N_6141);
nand U7460 (N_7460,N_6738,N_6562);
nand U7461 (N_7461,N_6529,N_6449);
xor U7462 (N_7462,N_6252,N_6696);
xor U7463 (N_7463,N_6095,N_6255);
and U7464 (N_7464,N_6268,N_6529);
nor U7465 (N_7465,N_6260,N_6681);
xor U7466 (N_7466,N_6170,N_6709);
nor U7467 (N_7467,N_6496,N_6122);
nand U7468 (N_7468,N_6066,N_6190);
or U7469 (N_7469,N_6175,N_6431);
and U7470 (N_7470,N_6246,N_6718);
nor U7471 (N_7471,N_6587,N_6067);
and U7472 (N_7472,N_6558,N_6484);
nand U7473 (N_7473,N_6323,N_6270);
or U7474 (N_7474,N_6385,N_6195);
xor U7475 (N_7475,N_6138,N_6632);
nor U7476 (N_7476,N_6003,N_6094);
nor U7477 (N_7477,N_6665,N_6349);
or U7478 (N_7478,N_6446,N_6205);
and U7479 (N_7479,N_6325,N_6725);
xor U7480 (N_7480,N_6687,N_6580);
nor U7481 (N_7481,N_6613,N_6650);
nand U7482 (N_7482,N_6686,N_6090);
or U7483 (N_7483,N_6118,N_6337);
or U7484 (N_7484,N_6456,N_6529);
nor U7485 (N_7485,N_6585,N_6203);
xor U7486 (N_7486,N_6247,N_6707);
xnor U7487 (N_7487,N_6510,N_6205);
or U7488 (N_7488,N_6571,N_6292);
nor U7489 (N_7489,N_6746,N_6712);
xnor U7490 (N_7490,N_6126,N_6031);
nor U7491 (N_7491,N_6729,N_6447);
xnor U7492 (N_7492,N_6547,N_6194);
or U7493 (N_7493,N_6112,N_6572);
xnor U7494 (N_7494,N_6634,N_6670);
and U7495 (N_7495,N_6642,N_6287);
nand U7496 (N_7496,N_6569,N_6236);
or U7497 (N_7497,N_6621,N_6092);
xor U7498 (N_7498,N_6612,N_6195);
and U7499 (N_7499,N_6283,N_6601);
xnor U7500 (N_7500,N_6845,N_7190);
or U7501 (N_7501,N_7451,N_7339);
nor U7502 (N_7502,N_6868,N_7289);
xor U7503 (N_7503,N_6809,N_6782);
xnor U7504 (N_7504,N_7295,N_6985);
or U7505 (N_7505,N_7262,N_7292);
or U7506 (N_7506,N_6988,N_6944);
nand U7507 (N_7507,N_7017,N_7398);
xor U7508 (N_7508,N_7444,N_6853);
nor U7509 (N_7509,N_7090,N_7142);
and U7510 (N_7510,N_7184,N_6768);
or U7511 (N_7511,N_7153,N_7027);
nor U7512 (N_7512,N_6956,N_7401);
nand U7513 (N_7513,N_7436,N_7166);
or U7514 (N_7514,N_7333,N_6967);
and U7515 (N_7515,N_7112,N_7192);
xnor U7516 (N_7516,N_7254,N_7094);
xor U7517 (N_7517,N_7197,N_7001);
or U7518 (N_7518,N_7404,N_7353);
or U7519 (N_7519,N_7224,N_7259);
nor U7520 (N_7520,N_7117,N_7187);
nand U7521 (N_7521,N_7091,N_7124);
or U7522 (N_7522,N_6839,N_7271);
and U7523 (N_7523,N_7114,N_7273);
nor U7524 (N_7524,N_6923,N_7180);
xor U7525 (N_7525,N_7176,N_7223);
or U7526 (N_7526,N_7391,N_7018);
xor U7527 (N_7527,N_7100,N_7138);
xor U7528 (N_7528,N_7051,N_7127);
xor U7529 (N_7529,N_7032,N_7321);
or U7530 (N_7530,N_7487,N_7287);
nor U7531 (N_7531,N_6996,N_7499);
or U7532 (N_7532,N_7128,N_7496);
or U7533 (N_7533,N_7354,N_7351);
nand U7534 (N_7534,N_6995,N_7244);
nand U7535 (N_7535,N_6767,N_7085);
and U7536 (N_7536,N_7123,N_7039);
or U7537 (N_7537,N_7250,N_6869);
xnor U7538 (N_7538,N_6787,N_7399);
xnor U7539 (N_7539,N_7409,N_6934);
and U7540 (N_7540,N_7479,N_6973);
and U7541 (N_7541,N_7159,N_7408);
nor U7542 (N_7542,N_6805,N_7358);
and U7543 (N_7543,N_6836,N_7331);
nand U7544 (N_7544,N_7055,N_6851);
and U7545 (N_7545,N_7490,N_7300);
nor U7546 (N_7546,N_6966,N_7340);
xor U7547 (N_7547,N_7312,N_7316);
nor U7548 (N_7548,N_7266,N_7483);
nand U7549 (N_7549,N_7420,N_7293);
and U7550 (N_7550,N_7392,N_7275);
nand U7551 (N_7551,N_7462,N_7104);
or U7552 (N_7552,N_6975,N_7194);
nor U7553 (N_7553,N_6825,N_6942);
or U7554 (N_7554,N_7381,N_7103);
xor U7555 (N_7555,N_7133,N_7163);
and U7556 (N_7556,N_6761,N_7208);
xnor U7557 (N_7557,N_7165,N_6838);
xor U7558 (N_7558,N_7081,N_7002);
nor U7559 (N_7559,N_6776,N_7044);
xor U7560 (N_7560,N_7365,N_7364);
nor U7561 (N_7561,N_6846,N_6897);
and U7562 (N_7562,N_7068,N_6870);
and U7563 (N_7563,N_6876,N_6806);
nor U7564 (N_7564,N_7116,N_6951);
and U7565 (N_7565,N_7062,N_7359);
or U7566 (N_7566,N_6879,N_7368);
or U7567 (N_7567,N_7431,N_7129);
or U7568 (N_7568,N_7013,N_7349);
or U7569 (N_7569,N_6913,N_6818);
or U7570 (N_7570,N_6878,N_7132);
xnor U7571 (N_7571,N_7181,N_6779);
or U7572 (N_7572,N_6802,N_7210);
nand U7573 (N_7573,N_6792,N_7171);
xnor U7574 (N_7574,N_7376,N_7414);
and U7575 (N_7575,N_7231,N_7086);
xor U7576 (N_7576,N_6887,N_6997);
nor U7577 (N_7577,N_7216,N_6992);
xnor U7578 (N_7578,N_6953,N_6907);
and U7579 (N_7579,N_6883,N_7387);
nand U7580 (N_7580,N_6841,N_7249);
xor U7581 (N_7581,N_7467,N_7394);
and U7582 (N_7582,N_6824,N_7237);
nand U7583 (N_7583,N_7229,N_7291);
and U7584 (N_7584,N_7480,N_7335);
and U7585 (N_7585,N_6752,N_7155);
or U7586 (N_7586,N_6819,N_7476);
or U7587 (N_7587,N_6989,N_7267);
and U7588 (N_7588,N_7345,N_6990);
nor U7589 (N_7589,N_7481,N_7228);
xor U7590 (N_7590,N_7378,N_7269);
or U7591 (N_7591,N_6908,N_7448);
nand U7592 (N_7592,N_6920,N_7182);
xnor U7593 (N_7593,N_7145,N_6909);
xnor U7594 (N_7594,N_7294,N_7141);
or U7595 (N_7595,N_7168,N_7384);
and U7596 (N_7596,N_7099,N_7074);
nand U7597 (N_7597,N_6837,N_7239);
nand U7598 (N_7598,N_7220,N_7227);
and U7599 (N_7599,N_6919,N_6892);
nor U7600 (N_7600,N_7232,N_6832);
xnor U7601 (N_7601,N_7063,N_6979);
nand U7602 (N_7602,N_7028,N_7463);
and U7603 (N_7603,N_7179,N_7149);
nand U7604 (N_7604,N_7200,N_7111);
xor U7605 (N_7605,N_7242,N_7206);
nand U7606 (N_7606,N_7373,N_6906);
or U7607 (N_7607,N_7494,N_7469);
or U7608 (N_7608,N_7457,N_7336);
xor U7609 (N_7609,N_7139,N_6843);
nor U7610 (N_7610,N_7024,N_6921);
nand U7611 (N_7611,N_7258,N_7067);
xor U7612 (N_7612,N_7105,N_6901);
or U7613 (N_7613,N_7076,N_7298);
xnor U7614 (N_7614,N_7183,N_7393);
nand U7615 (N_7615,N_7043,N_7233);
and U7616 (N_7616,N_7069,N_6866);
xor U7617 (N_7617,N_7033,N_7285);
nor U7618 (N_7618,N_7484,N_7029);
nor U7619 (N_7619,N_7140,N_7157);
xnor U7620 (N_7620,N_7264,N_6881);
or U7621 (N_7621,N_6938,N_7425);
or U7622 (N_7622,N_6964,N_6855);
or U7623 (N_7623,N_6981,N_7022);
xor U7624 (N_7624,N_7198,N_7252);
or U7625 (N_7625,N_7097,N_7428);
nor U7626 (N_7626,N_7397,N_7201);
or U7627 (N_7627,N_7413,N_6960);
nand U7628 (N_7628,N_7489,N_7379);
nand U7629 (N_7629,N_6800,N_7424);
nor U7630 (N_7630,N_7209,N_7311);
nand U7631 (N_7631,N_7486,N_7355);
nor U7632 (N_7632,N_7066,N_7026);
xnor U7633 (N_7633,N_7073,N_6918);
nor U7634 (N_7634,N_7309,N_7301);
xnor U7635 (N_7635,N_6904,N_7202);
or U7636 (N_7636,N_7452,N_7281);
or U7637 (N_7637,N_7418,N_6753);
or U7638 (N_7638,N_7042,N_7341);
and U7639 (N_7639,N_6797,N_7008);
or U7640 (N_7640,N_6929,N_7240);
nand U7641 (N_7641,N_7025,N_6820);
and U7642 (N_7642,N_6927,N_7234);
and U7643 (N_7643,N_6780,N_6860);
nand U7644 (N_7644,N_7477,N_7260);
and U7645 (N_7645,N_7071,N_7326);
and U7646 (N_7646,N_6771,N_7386);
nor U7647 (N_7647,N_7478,N_7310);
or U7648 (N_7648,N_6946,N_7423);
xor U7649 (N_7649,N_7474,N_7348);
nand U7650 (N_7650,N_7322,N_7430);
xor U7651 (N_7651,N_7265,N_7372);
nor U7652 (N_7652,N_7306,N_7460);
and U7653 (N_7653,N_6833,N_6835);
xnor U7654 (N_7654,N_6757,N_6793);
nand U7655 (N_7655,N_7215,N_7064);
nand U7656 (N_7656,N_6970,N_6847);
nand U7657 (N_7657,N_7156,N_6939);
or U7658 (N_7658,N_7172,N_7412);
and U7659 (N_7659,N_6961,N_6755);
or U7660 (N_7660,N_7174,N_6903);
or U7661 (N_7661,N_6854,N_7113);
or U7662 (N_7662,N_6807,N_6922);
nor U7663 (N_7663,N_7052,N_6828);
xnor U7664 (N_7664,N_7261,N_7175);
nor U7665 (N_7665,N_7130,N_7049);
and U7666 (N_7666,N_7263,N_7432);
nor U7667 (N_7667,N_6882,N_6926);
or U7668 (N_7668,N_7251,N_7473);
xor U7669 (N_7669,N_7374,N_7169);
or U7670 (N_7670,N_6982,N_7098);
nor U7671 (N_7671,N_7422,N_7492);
and U7672 (N_7672,N_6827,N_6999);
nand U7673 (N_7673,N_7126,N_6993);
xor U7674 (N_7674,N_6965,N_7065);
or U7675 (N_7675,N_7204,N_7147);
nand U7676 (N_7676,N_6830,N_7257);
or U7677 (N_7677,N_7015,N_7107);
nor U7678 (N_7678,N_7390,N_7010);
nor U7679 (N_7679,N_7199,N_7170);
or U7680 (N_7680,N_7407,N_6900);
or U7681 (N_7681,N_7191,N_7058);
xor U7682 (N_7682,N_7019,N_6814);
nand U7683 (N_7683,N_7054,N_7075);
and U7684 (N_7684,N_7110,N_7135);
or U7685 (N_7685,N_7070,N_7415);
or U7686 (N_7686,N_6987,N_7256);
nor U7687 (N_7687,N_7437,N_7217);
and U7688 (N_7688,N_7461,N_6821);
or U7689 (N_7689,N_7031,N_6874);
nor U7690 (N_7690,N_6849,N_7352);
and U7691 (N_7691,N_7270,N_6758);
or U7692 (N_7692,N_7102,N_6763);
nand U7693 (N_7693,N_7297,N_7343);
nand U7694 (N_7694,N_7303,N_7442);
nor U7695 (N_7695,N_6784,N_7317);
and U7696 (N_7696,N_7230,N_6986);
or U7697 (N_7697,N_7411,N_7361);
xnor U7698 (N_7698,N_6925,N_6816);
nor U7699 (N_7699,N_7417,N_6844);
and U7700 (N_7700,N_6850,N_7421);
and U7701 (N_7701,N_7319,N_7445);
nor U7702 (N_7702,N_7497,N_6813);
xor U7703 (N_7703,N_6886,N_7446);
nor U7704 (N_7704,N_7334,N_6871);
or U7705 (N_7705,N_7009,N_6983);
or U7706 (N_7706,N_6902,N_7125);
and U7707 (N_7707,N_7109,N_6932);
or U7708 (N_7708,N_7093,N_7283);
or U7709 (N_7709,N_7482,N_7402);
nand U7710 (N_7710,N_7385,N_7456);
xnor U7711 (N_7711,N_7164,N_7041);
and U7712 (N_7712,N_7318,N_7214);
nand U7713 (N_7713,N_7106,N_6950);
and U7714 (N_7714,N_7219,N_7225);
nand U7715 (N_7715,N_7324,N_7416);
nand U7716 (N_7716,N_7357,N_6957);
nor U7717 (N_7717,N_7395,N_7455);
nand U7718 (N_7718,N_6875,N_6930);
nand U7719 (N_7719,N_7186,N_7185);
nor U7720 (N_7720,N_7441,N_7344);
xnor U7721 (N_7721,N_7406,N_7320);
and U7722 (N_7722,N_7000,N_6756);
nor U7723 (N_7723,N_6774,N_6941);
nand U7724 (N_7724,N_7274,N_7282);
xnor U7725 (N_7725,N_7003,N_7205);
and U7726 (N_7726,N_7082,N_6783);
or U7727 (N_7727,N_7360,N_7327);
and U7728 (N_7728,N_7447,N_7092);
nand U7729 (N_7729,N_7095,N_7014);
or U7730 (N_7730,N_6865,N_6772);
nor U7731 (N_7731,N_7380,N_7434);
xnor U7732 (N_7732,N_7362,N_7276);
nor U7733 (N_7733,N_7466,N_7196);
and U7734 (N_7734,N_6978,N_7458);
or U7735 (N_7735,N_6750,N_6896);
xnor U7736 (N_7736,N_6893,N_7268);
nor U7737 (N_7737,N_6826,N_7299);
and U7738 (N_7738,N_7011,N_6791);
or U7739 (N_7739,N_7059,N_7167);
nand U7740 (N_7740,N_7211,N_7144);
nand U7741 (N_7741,N_7388,N_7382);
nand U7742 (N_7742,N_6994,N_6895);
xor U7743 (N_7743,N_7405,N_7410);
nor U7744 (N_7744,N_6974,N_7089);
nor U7745 (N_7745,N_6785,N_7366);
and U7746 (N_7746,N_6799,N_7241);
xnor U7747 (N_7747,N_7272,N_7302);
or U7748 (N_7748,N_6773,N_7329);
nor U7749 (N_7749,N_6856,N_7246);
or U7750 (N_7750,N_7435,N_7150);
xor U7751 (N_7751,N_6928,N_7471);
or U7752 (N_7752,N_6891,N_6872);
and U7753 (N_7753,N_6910,N_6977);
or U7754 (N_7754,N_7193,N_7307);
nand U7755 (N_7755,N_7493,N_7060);
or U7756 (N_7756,N_7488,N_7440);
xor U7757 (N_7757,N_6789,N_7450);
nor U7758 (N_7758,N_7396,N_6831);
nor U7759 (N_7759,N_6778,N_7120);
and U7760 (N_7760,N_6889,N_7347);
or U7761 (N_7761,N_7213,N_7243);
nor U7762 (N_7762,N_7449,N_7235);
nand U7763 (N_7763,N_7383,N_7038);
and U7764 (N_7764,N_6984,N_7305);
nand U7765 (N_7765,N_7439,N_6955);
nor U7766 (N_7766,N_6834,N_7346);
and U7767 (N_7767,N_7464,N_7119);
nand U7768 (N_7768,N_6808,N_6890);
nor U7769 (N_7769,N_6848,N_7077);
or U7770 (N_7770,N_6829,N_6781);
nor U7771 (N_7771,N_6940,N_7438);
nor U7772 (N_7772,N_6790,N_7178);
nand U7773 (N_7773,N_7021,N_6823);
and U7774 (N_7774,N_7400,N_7443);
and U7775 (N_7775,N_7048,N_7203);
and U7776 (N_7776,N_7152,N_6911);
nand U7777 (N_7777,N_7255,N_6976);
or U7778 (N_7778,N_7491,N_6867);
nand U7779 (N_7779,N_6817,N_7350);
and U7780 (N_7780,N_6863,N_7296);
nor U7781 (N_7781,N_7007,N_6765);
or U7782 (N_7782,N_7313,N_7495);
nand U7783 (N_7783,N_6760,N_7371);
or U7784 (N_7784,N_7328,N_7108);
nand U7785 (N_7785,N_6840,N_7162);
nor U7786 (N_7786,N_6945,N_6852);
nor U7787 (N_7787,N_7323,N_7173);
xor U7788 (N_7788,N_7101,N_7084);
or U7789 (N_7789,N_7088,N_7047);
xor U7790 (N_7790,N_6899,N_7148);
nor U7791 (N_7791,N_7056,N_7284);
xnor U7792 (N_7792,N_6764,N_7134);
nand U7793 (N_7793,N_7160,N_7330);
and U7794 (N_7794,N_7136,N_7072);
nand U7795 (N_7795,N_6762,N_7034);
or U7796 (N_7796,N_7061,N_7012);
xor U7797 (N_7797,N_7470,N_7121);
or U7798 (N_7798,N_7403,N_6810);
and U7799 (N_7799,N_7226,N_7337);
and U7800 (N_7800,N_6980,N_7485);
nand U7801 (N_7801,N_6858,N_6914);
nor U7802 (N_7802,N_7286,N_7375);
or U7803 (N_7803,N_6759,N_7057);
xnor U7804 (N_7804,N_6898,N_6917);
nor U7805 (N_7805,N_7079,N_7290);
nand U7806 (N_7806,N_6933,N_7037);
and U7807 (N_7807,N_6916,N_6864);
xnor U7808 (N_7808,N_6954,N_7468);
xnor U7809 (N_7809,N_6971,N_6795);
nand U7810 (N_7810,N_7046,N_7221);
xor U7811 (N_7811,N_6754,N_7080);
or U7812 (N_7812,N_6972,N_7115);
nand U7813 (N_7813,N_6794,N_7177);
xor U7814 (N_7814,N_7035,N_7247);
and U7815 (N_7815,N_6777,N_6859);
nand U7816 (N_7816,N_6959,N_6894);
nor U7817 (N_7817,N_6786,N_7369);
xor U7818 (N_7818,N_6842,N_7377);
nand U7819 (N_7819,N_6991,N_6862);
nand U7820 (N_7820,N_7006,N_7189);
and U7821 (N_7821,N_7030,N_7004);
nor U7822 (N_7822,N_6796,N_6766);
and U7823 (N_7823,N_7475,N_6801);
xnor U7824 (N_7824,N_6948,N_6812);
and U7825 (N_7825,N_6751,N_7083);
and U7826 (N_7826,N_7288,N_7137);
xnor U7827 (N_7827,N_7426,N_6798);
and U7828 (N_7828,N_7277,N_7465);
nand U7829 (N_7829,N_7304,N_6885);
or U7830 (N_7830,N_7363,N_7053);
nor U7831 (N_7831,N_6815,N_7161);
or U7832 (N_7832,N_6969,N_7122);
nand U7833 (N_7833,N_7143,N_6861);
and U7834 (N_7834,N_7023,N_7472);
nand U7835 (N_7835,N_6924,N_7096);
nand U7836 (N_7836,N_7338,N_6877);
xnor U7837 (N_7837,N_7154,N_7238);
nor U7838 (N_7838,N_6962,N_6880);
nand U7839 (N_7839,N_6937,N_6943);
nand U7840 (N_7840,N_6963,N_6949);
and U7841 (N_7841,N_7245,N_7195);
xnor U7842 (N_7842,N_6873,N_6905);
nand U7843 (N_7843,N_7040,N_6770);
or U7844 (N_7844,N_6952,N_7087);
nand U7845 (N_7845,N_7280,N_7429);
nand U7846 (N_7846,N_7005,N_7045);
nand U7847 (N_7847,N_7325,N_7236);
and U7848 (N_7848,N_7131,N_6857);
and U7849 (N_7849,N_7253,N_7279);
or U7850 (N_7850,N_7498,N_7433);
and U7851 (N_7851,N_7356,N_7036);
xnor U7852 (N_7852,N_7332,N_7454);
nor U7853 (N_7853,N_7248,N_7078);
nand U7854 (N_7854,N_6936,N_7050);
nor U7855 (N_7855,N_7308,N_6958);
xnor U7856 (N_7856,N_7118,N_6912);
or U7857 (N_7857,N_7151,N_7419);
or U7858 (N_7858,N_7146,N_6931);
nor U7859 (N_7859,N_7342,N_7278);
and U7860 (N_7860,N_7367,N_6811);
nor U7861 (N_7861,N_7315,N_6788);
nor U7862 (N_7862,N_6803,N_6915);
and U7863 (N_7863,N_6947,N_6968);
and U7864 (N_7864,N_7188,N_6804);
nand U7865 (N_7865,N_6884,N_7222);
and U7866 (N_7866,N_6998,N_6775);
and U7867 (N_7867,N_7453,N_6935);
nand U7868 (N_7868,N_6888,N_6822);
or U7869 (N_7869,N_7370,N_7020);
xnor U7870 (N_7870,N_7389,N_7459);
xor U7871 (N_7871,N_7427,N_7158);
and U7872 (N_7872,N_7212,N_7314);
nor U7873 (N_7873,N_6769,N_7016);
nor U7874 (N_7874,N_7218,N_7207);
nor U7875 (N_7875,N_6795,N_7181);
or U7876 (N_7876,N_7343,N_6961);
nor U7877 (N_7877,N_7408,N_6901);
xnor U7878 (N_7878,N_6817,N_7409);
xnor U7879 (N_7879,N_6894,N_7209);
and U7880 (N_7880,N_7084,N_6866);
xnor U7881 (N_7881,N_7289,N_6791);
and U7882 (N_7882,N_7384,N_7175);
nor U7883 (N_7883,N_7343,N_7449);
nor U7884 (N_7884,N_6820,N_6900);
nand U7885 (N_7885,N_7215,N_7461);
xnor U7886 (N_7886,N_7182,N_7330);
and U7887 (N_7887,N_6917,N_7115);
nor U7888 (N_7888,N_7278,N_7271);
xor U7889 (N_7889,N_7254,N_6961);
xnor U7890 (N_7890,N_7384,N_7484);
nor U7891 (N_7891,N_7196,N_6869);
nor U7892 (N_7892,N_6878,N_7213);
nor U7893 (N_7893,N_6979,N_7419);
xnor U7894 (N_7894,N_7080,N_7169);
nor U7895 (N_7895,N_7266,N_7037);
nand U7896 (N_7896,N_6750,N_7039);
nand U7897 (N_7897,N_7412,N_6754);
nand U7898 (N_7898,N_7050,N_7280);
and U7899 (N_7899,N_7276,N_6993);
or U7900 (N_7900,N_6820,N_7313);
and U7901 (N_7901,N_7438,N_7453);
or U7902 (N_7902,N_7177,N_7166);
nand U7903 (N_7903,N_6904,N_7278);
xnor U7904 (N_7904,N_6969,N_7329);
xnor U7905 (N_7905,N_7107,N_6845);
nand U7906 (N_7906,N_6778,N_7425);
nor U7907 (N_7907,N_7492,N_6823);
nand U7908 (N_7908,N_7172,N_6800);
and U7909 (N_7909,N_6797,N_6767);
nand U7910 (N_7910,N_7441,N_6754);
nor U7911 (N_7911,N_7330,N_7334);
and U7912 (N_7912,N_7346,N_6917);
nor U7913 (N_7913,N_6866,N_7110);
nor U7914 (N_7914,N_6810,N_7232);
and U7915 (N_7915,N_7028,N_7056);
nand U7916 (N_7916,N_7064,N_6877);
or U7917 (N_7917,N_6916,N_7385);
and U7918 (N_7918,N_6838,N_7328);
nor U7919 (N_7919,N_7244,N_7480);
and U7920 (N_7920,N_7421,N_7140);
nor U7921 (N_7921,N_6835,N_7124);
xor U7922 (N_7922,N_6764,N_7049);
xor U7923 (N_7923,N_7163,N_6797);
nor U7924 (N_7924,N_6917,N_7025);
or U7925 (N_7925,N_7125,N_6813);
nor U7926 (N_7926,N_7073,N_7120);
or U7927 (N_7927,N_7162,N_7396);
or U7928 (N_7928,N_7119,N_7188);
or U7929 (N_7929,N_7069,N_6868);
or U7930 (N_7930,N_7125,N_6978);
xor U7931 (N_7931,N_6919,N_7201);
nand U7932 (N_7932,N_6946,N_7253);
or U7933 (N_7933,N_6850,N_7298);
or U7934 (N_7934,N_7248,N_7070);
or U7935 (N_7935,N_7214,N_7039);
nor U7936 (N_7936,N_7166,N_6758);
and U7937 (N_7937,N_7460,N_7062);
xor U7938 (N_7938,N_7034,N_6755);
and U7939 (N_7939,N_7431,N_7031);
nor U7940 (N_7940,N_7445,N_6825);
nor U7941 (N_7941,N_7489,N_7371);
nor U7942 (N_7942,N_7213,N_6964);
nor U7943 (N_7943,N_7308,N_7164);
and U7944 (N_7944,N_7085,N_6982);
or U7945 (N_7945,N_7067,N_7415);
or U7946 (N_7946,N_6887,N_7337);
and U7947 (N_7947,N_7191,N_7222);
and U7948 (N_7948,N_7135,N_7112);
nand U7949 (N_7949,N_7281,N_6925);
xor U7950 (N_7950,N_7067,N_7042);
nor U7951 (N_7951,N_7209,N_7382);
nor U7952 (N_7952,N_6848,N_7414);
nor U7953 (N_7953,N_7039,N_7192);
and U7954 (N_7954,N_6761,N_7143);
or U7955 (N_7955,N_7481,N_7032);
nand U7956 (N_7956,N_7222,N_7148);
nand U7957 (N_7957,N_7420,N_6811);
or U7958 (N_7958,N_7140,N_7323);
xor U7959 (N_7959,N_6885,N_7419);
or U7960 (N_7960,N_6751,N_6750);
xor U7961 (N_7961,N_6760,N_7150);
or U7962 (N_7962,N_6754,N_7487);
and U7963 (N_7963,N_7374,N_7184);
nand U7964 (N_7964,N_6778,N_6816);
nor U7965 (N_7965,N_6879,N_7439);
or U7966 (N_7966,N_7460,N_7169);
nor U7967 (N_7967,N_6938,N_7006);
xor U7968 (N_7968,N_7463,N_7489);
or U7969 (N_7969,N_6844,N_7113);
xnor U7970 (N_7970,N_7449,N_7084);
xnor U7971 (N_7971,N_7269,N_7478);
or U7972 (N_7972,N_7114,N_7053);
or U7973 (N_7973,N_7136,N_7260);
nor U7974 (N_7974,N_7447,N_7244);
nor U7975 (N_7975,N_7413,N_6805);
nor U7976 (N_7976,N_6859,N_7053);
xnor U7977 (N_7977,N_7142,N_7247);
and U7978 (N_7978,N_6785,N_7250);
nor U7979 (N_7979,N_7087,N_7254);
and U7980 (N_7980,N_6987,N_7364);
nor U7981 (N_7981,N_7289,N_7186);
nand U7982 (N_7982,N_7136,N_7023);
or U7983 (N_7983,N_7127,N_6952);
and U7984 (N_7984,N_7267,N_7222);
xor U7985 (N_7985,N_6883,N_7245);
nor U7986 (N_7986,N_7210,N_7090);
nand U7987 (N_7987,N_7008,N_7324);
nor U7988 (N_7988,N_7026,N_6848);
or U7989 (N_7989,N_7388,N_6790);
nor U7990 (N_7990,N_7160,N_7122);
nor U7991 (N_7991,N_7163,N_7274);
or U7992 (N_7992,N_7246,N_7408);
or U7993 (N_7993,N_7422,N_7150);
and U7994 (N_7994,N_7163,N_7118);
and U7995 (N_7995,N_7025,N_6991);
xor U7996 (N_7996,N_7277,N_6808);
nand U7997 (N_7997,N_7431,N_6755);
nor U7998 (N_7998,N_6988,N_6833);
xor U7999 (N_7999,N_6919,N_7089);
or U8000 (N_8000,N_6960,N_7486);
nand U8001 (N_8001,N_7023,N_7268);
nand U8002 (N_8002,N_7366,N_6873);
nand U8003 (N_8003,N_6813,N_7085);
nor U8004 (N_8004,N_7144,N_7292);
nor U8005 (N_8005,N_6848,N_7263);
xnor U8006 (N_8006,N_6988,N_6879);
and U8007 (N_8007,N_7090,N_7056);
or U8008 (N_8008,N_6891,N_6827);
and U8009 (N_8009,N_7291,N_6924);
nand U8010 (N_8010,N_7223,N_7355);
nor U8011 (N_8011,N_7038,N_7353);
or U8012 (N_8012,N_7333,N_7258);
nor U8013 (N_8013,N_6791,N_6852);
xnor U8014 (N_8014,N_6861,N_7474);
nand U8015 (N_8015,N_7409,N_7251);
nor U8016 (N_8016,N_7139,N_7368);
nor U8017 (N_8017,N_7287,N_7195);
or U8018 (N_8018,N_6998,N_6831);
or U8019 (N_8019,N_7206,N_6900);
xnor U8020 (N_8020,N_7106,N_7098);
nor U8021 (N_8021,N_7453,N_7195);
nand U8022 (N_8022,N_7086,N_7036);
nand U8023 (N_8023,N_7212,N_6960);
or U8024 (N_8024,N_6807,N_7102);
and U8025 (N_8025,N_7300,N_7370);
or U8026 (N_8026,N_6984,N_6987);
and U8027 (N_8027,N_7447,N_6909);
nand U8028 (N_8028,N_6825,N_7154);
nand U8029 (N_8029,N_7409,N_7056);
and U8030 (N_8030,N_7437,N_7499);
xor U8031 (N_8031,N_7382,N_7454);
and U8032 (N_8032,N_7037,N_6834);
xnor U8033 (N_8033,N_6875,N_6801);
xnor U8034 (N_8034,N_7125,N_7152);
nand U8035 (N_8035,N_6843,N_6865);
and U8036 (N_8036,N_7135,N_7055);
nor U8037 (N_8037,N_7348,N_6890);
or U8038 (N_8038,N_7106,N_6845);
xnor U8039 (N_8039,N_7467,N_7015);
and U8040 (N_8040,N_7376,N_7147);
xor U8041 (N_8041,N_7032,N_7104);
xor U8042 (N_8042,N_7257,N_7031);
nor U8043 (N_8043,N_7203,N_7376);
or U8044 (N_8044,N_7173,N_6777);
xnor U8045 (N_8045,N_7323,N_7312);
and U8046 (N_8046,N_7488,N_7143);
nand U8047 (N_8047,N_6956,N_7259);
nor U8048 (N_8048,N_7298,N_6935);
nand U8049 (N_8049,N_7347,N_7053);
nor U8050 (N_8050,N_6905,N_7322);
nor U8051 (N_8051,N_6973,N_6806);
or U8052 (N_8052,N_7203,N_6922);
and U8053 (N_8053,N_7100,N_7257);
xnor U8054 (N_8054,N_7073,N_6927);
xor U8055 (N_8055,N_6813,N_7157);
and U8056 (N_8056,N_6994,N_7098);
or U8057 (N_8057,N_6873,N_7100);
nor U8058 (N_8058,N_7072,N_6803);
nand U8059 (N_8059,N_7327,N_6807);
nand U8060 (N_8060,N_6885,N_6796);
and U8061 (N_8061,N_7107,N_6957);
nor U8062 (N_8062,N_7203,N_7012);
nand U8063 (N_8063,N_7015,N_7319);
nor U8064 (N_8064,N_7283,N_7188);
nor U8065 (N_8065,N_6846,N_7105);
or U8066 (N_8066,N_7275,N_7343);
and U8067 (N_8067,N_6823,N_6864);
and U8068 (N_8068,N_6818,N_6810);
or U8069 (N_8069,N_7434,N_7489);
xnor U8070 (N_8070,N_7044,N_7483);
or U8071 (N_8071,N_7393,N_6768);
nand U8072 (N_8072,N_7006,N_6780);
nand U8073 (N_8073,N_7150,N_7372);
nand U8074 (N_8074,N_7464,N_6877);
and U8075 (N_8075,N_7401,N_7388);
or U8076 (N_8076,N_7225,N_7441);
nor U8077 (N_8077,N_7413,N_7434);
nand U8078 (N_8078,N_7261,N_7465);
and U8079 (N_8079,N_6942,N_6939);
xnor U8080 (N_8080,N_6947,N_7106);
nand U8081 (N_8081,N_6993,N_6799);
xor U8082 (N_8082,N_7251,N_7355);
nor U8083 (N_8083,N_7363,N_6948);
xnor U8084 (N_8084,N_7060,N_7111);
and U8085 (N_8085,N_6898,N_6809);
xor U8086 (N_8086,N_6920,N_6771);
or U8087 (N_8087,N_7452,N_7295);
or U8088 (N_8088,N_7199,N_6772);
nand U8089 (N_8089,N_6990,N_7189);
xnor U8090 (N_8090,N_6890,N_7223);
and U8091 (N_8091,N_6809,N_6910);
nand U8092 (N_8092,N_6910,N_7465);
or U8093 (N_8093,N_7102,N_6889);
xnor U8094 (N_8094,N_7113,N_7187);
and U8095 (N_8095,N_6816,N_7329);
and U8096 (N_8096,N_7091,N_7231);
xnor U8097 (N_8097,N_7329,N_7099);
nand U8098 (N_8098,N_6818,N_7087);
or U8099 (N_8099,N_6897,N_7371);
nor U8100 (N_8100,N_7491,N_7485);
nand U8101 (N_8101,N_6980,N_7097);
nand U8102 (N_8102,N_7216,N_7023);
xnor U8103 (N_8103,N_6794,N_6875);
xnor U8104 (N_8104,N_7316,N_6924);
nor U8105 (N_8105,N_7379,N_7451);
xnor U8106 (N_8106,N_7086,N_7128);
xnor U8107 (N_8107,N_7130,N_6997);
or U8108 (N_8108,N_7162,N_7118);
or U8109 (N_8109,N_6861,N_7120);
nand U8110 (N_8110,N_6862,N_7248);
xor U8111 (N_8111,N_6901,N_7086);
or U8112 (N_8112,N_7316,N_7266);
nand U8113 (N_8113,N_7470,N_7314);
and U8114 (N_8114,N_7354,N_6949);
or U8115 (N_8115,N_7281,N_7204);
nand U8116 (N_8116,N_7065,N_6891);
and U8117 (N_8117,N_6989,N_6819);
and U8118 (N_8118,N_7150,N_6804);
nor U8119 (N_8119,N_7060,N_7301);
nand U8120 (N_8120,N_7168,N_6837);
xor U8121 (N_8121,N_7222,N_7028);
xnor U8122 (N_8122,N_6816,N_7066);
nand U8123 (N_8123,N_6798,N_7039);
nand U8124 (N_8124,N_7289,N_6804);
or U8125 (N_8125,N_6833,N_7436);
nand U8126 (N_8126,N_7038,N_7237);
nor U8127 (N_8127,N_7494,N_7468);
or U8128 (N_8128,N_6763,N_6895);
and U8129 (N_8129,N_7236,N_7496);
xor U8130 (N_8130,N_7251,N_7415);
xnor U8131 (N_8131,N_7033,N_7214);
nor U8132 (N_8132,N_7325,N_7418);
and U8133 (N_8133,N_6823,N_7193);
or U8134 (N_8134,N_7214,N_7157);
or U8135 (N_8135,N_6964,N_7414);
nand U8136 (N_8136,N_7462,N_7283);
and U8137 (N_8137,N_7487,N_7161);
or U8138 (N_8138,N_7242,N_7131);
xnor U8139 (N_8139,N_7336,N_7190);
nor U8140 (N_8140,N_7125,N_7475);
or U8141 (N_8141,N_7148,N_7040);
nand U8142 (N_8142,N_7104,N_7285);
nor U8143 (N_8143,N_7472,N_7069);
nor U8144 (N_8144,N_7003,N_7387);
or U8145 (N_8145,N_7405,N_6811);
and U8146 (N_8146,N_6807,N_6875);
nor U8147 (N_8147,N_6846,N_6944);
nor U8148 (N_8148,N_7464,N_7120);
nor U8149 (N_8149,N_7110,N_6778);
and U8150 (N_8150,N_7301,N_6776);
or U8151 (N_8151,N_6954,N_7395);
nand U8152 (N_8152,N_7446,N_7042);
and U8153 (N_8153,N_7033,N_7240);
xnor U8154 (N_8154,N_7026,N_7484);
xnor U8155 (N_8155,N_6898,N_7191);
xnor U8156 (N_8156,N_6960,N_7125);
xnor U8157 (N_8157,N_7056,N_7367);
nor U8158 (N_8158,N_7349,N_7015);
and U8159 (N_8159,N_7191,N_7277);
xnor U8160 (N_8160,N_7107,N_6765);
xnor U8161 (N_8161,N_6763,N_7182);
nor U8162 (N_8162,N_7262,N_7434);
nor U8163 (N_8163,N_7351,N_6928);
nand U8164 (N_8164,N_7338,N_7481);
xor U8165 (N_8165,N_6838,N_6808);
xnor U8166 (N_8166,N_6943,N_6782);
nand U8167 (N_8167,N_7268,N_6798);
and U8168 (N_8168,N_7074,N_7403);
or U8169 (N_8169,N_7463,N_6773);
xor U8170 (N_8170,N_6772,N_6961);
and U8171 (N_8171,N_7343,N_7315);
nand U8172 (N_8172,N_7188,N_6814);
xor U8173 (N_8173,N_7109,N_7169);
nor U8174 (N_8174,N_7074,N_6918);
or U8175 (N_8175,N_7270,N_7065);
nor U8176 (N_8176,N_6794,N_7113);
xor U8177 (N_8177,N_7241,N_7177);
and U8178 (N_8178,N_6807,N_7212);
and U8179 (N_8179,N_7078,N_7437);
nor U8180 (N_8180,N_7457,N_7170);
and U8181 (N_8181,N_7128,N_7105);
or U8182 (N_8182,N_7374,N_6807);
xnor U8183 (N_8183,N_6981,N_7023);
nand U8184 (N_8184,N_6780,N_7306);
nor U8185 (N_8185,N_7212,N_6822);
and U8186 (N_8186,N_7372,N_7269);
and U8187 (N_8187,N_7193,N_6816);
and U8188 (N_8188,N_7413,N_7453);
nand U8189 (N_8189,N_7199,N_7460);
xor U8190 (N_8190,N_7242,N_7477);
nand U8191 (N_8191,N_7232,N_6898);
nor U8192 (N_8192,N_6796,N_7492);
nor U8193 (N_8193,N_6839,N_7483);
nor U8194 (N_8194,N_7147,N_7106);
nor U8195 (N_8195,N_7189,N_7457);
or U8196 (N_8196,N_7122,N_7212);
xor U8197 (N_8197,N_7260,N_6962);
nor U8198 (N_8198,N_7168,N_7237);
xnor U8199 (N_8199,N_7059,N_6802);
nor U8200 (N_8200,N_7047,N_6849);
and U8201 (N_8201,N_7305,N_7106);
or U8202 (N_8202,N_6995,N_7304);
and U8203 (N_8203,N_6827,N_7062);
or U8204 (N_8204,N_7212,N_6878);
and U8205 (N_8205,N_7292,N_7410);
and U8206 (N_8206,N_6961,N_6819);
nor U8207 (N_8207,N_7387,N_7490);
or U8208 (N_8208,N_7475,N_7352);
and U8209 (N_8209,N_6846,N_7140);
and U8210 (N_8210,N_6946,N_7232);
xnor U8211 (N_8211,N_7349,N_6850);
nor U8212 (N_8212,N_7004,N_7308);
and U8213 (N_8213,N_7029,N_6786);
nor U8214 (N_8214,N_7096,N_7455);
and U8215 (N_8215,N_7287,N_6905);
or U8216 (N_8216,N_7156,N_6933);
nor U8217 (N_8217,N_7204,N_7242);
or U8218 (N_8218,N_7496,N_7437);
or U8219 (N_8219,N_7172,N_7342);
nor U8220 (N_8220,N_6854,N_7001);
or U8221 (N_8221,N_6796,N_7158);
or U8222 (N_8222,N_7304,N_7039);
nor U8223 (N_8223,N_7359,N_6991);
nor U8224 (N_8224,N_6950,N_7157);
nor U8225 (N_8225,N_6850,N_7392);
or U8226 (N_8226,N_7066,N_6940);
nor U8227 (N_8227,N_6901,N_6911);
xor U8228 (N_8228,N_7127,N_6782);
and U8229 (N_8229,N_7345,N_7136);
and U8230 (N_8230,N_7266,N_6803);
or U8231 (N_8231,N_7402,N_6994);
and U8232 (N_8232,N_6772,N_6760);
nand U8233 (N_8233,N_7234,N_7188);
or U8234 (N_8234,N_7013,N_7205);
and U8235 (N_8235,N_6849,N_7122);
and U8236 (N_8236,N_7028,N_7054);
xnor U8237 (N_8237,N_7283,N_7250);
and U8238 (N_8238,N_7181,N_7216);
and U8239 (N_8239,N_6938,N_6859);
nor U8240 (N_8240,N_7286,N_7099);
xor U8241 (N_8241,N_7457,N_7389);
and U8242 (N_8242,N_6765,N_7085);
nor U8243 (N_8243,N_7058,N_7024);
nor U8244 (N_8244,N_7463,N_7048);
xnor U8245 (N_8245,N_6842,N_6907);
nand U8246 (N_8246,N_6933,N_6862);
or U8247 (N_8247,N_6852,N_7444);
nor U8248 (N_8248,N_7498,N_7280);
and U8249 (N_8249,N_7142,N_7085);
and U8250 (N_8250,N_7978,N_7968);
and U8251 (N_8251,N_7597,N_7504);
nor U8252 (N_8252,N_7598,N_8132);
and U8253 (N_8253,N_7595,N_8004);
nor U8254 (N_8254,N_7743,N_8179);
nor U8255 (N_8255,N_7508,N_8120);
and U8256 (N_8256,N_7678,N_7509);
and U8257 (N_8257,N_7822,N_7856);
and U8258 (N_8258,N_7719,N_8152);
xnor U8259 (N_8259,N_8029,N_7658);
xnor U8260 (N_8260,N_8162,N_7692);
or U8261 (N_8261,N_8195,N_7531);
and U8262 (N_8262,N_7993,N_7904);
xor U8263 (N_8263,N_7611,N_7606);
and U8264 (N_8264,N_7906,N_8196);
nor U8265 (N_8265,N_7757,N_7529);
nor U8266 (N_8266,N_7868,N_7707);
and U8267 (N_8267,N_7849,N_8108);
xor U8268 (N_8268,N_7729,N_8115);
or U8269 (N_8269,N_7960,N_7772);
nand U8270 (N_8270,N_7622,N_7789);
or U8271 (N_8271,N_7565,N_7992);
or U8272 (N_8272,N_7961,N_7862);
xor U8273 (N_8273,N_8185,N_8220);
nand U8274 (N_8274,N_7874,N_7963);
nor U8275 (N_8275,N_7558,N_8032);
nand U8276 (N_8276,N_7875,N_7712);
xnor U8277 (N_8277,N_8138,N_7843);
nor U8278 (N_8278,N_7831,N_7742);
xor U8279 (N_8279,N_7947,N_7932);
nand U8280 (N_8280,N_8170,N_7768);
or U8281 (N_8281,N_7636,N_7846);
and U8282 (N_8282,N_7819,N_8001);
nor U8283 (N_8283,N_8155,N_7762);
and U8284 (N_8284,N_7740,N_7863);
or U8285 (N_8285,N_8190,N_8058);
nor U8286 (N_8286,N_7527,N_7841);
and U8287 (N_8287,N_8079,N_7809);
or U8288 (N_8288,N_7589,N_8098);
nor U8289 (N_8289,N_7745,N_7642);
nor U8290 (N_8290,N_7550,N_8036);
xnor U8291 (N_8291,N_7786,N_7782);
nor U8292 (N_8292,N_8116,N_7832);
nor U8293 (N_8293,N_7921,N_7705);
or U8294 (N_8294,N_7853,N_7990);
nand U8295 (N_8295,N_7821,N_7510);
nand U8296 (N_8296,N_7860,N_8021);
nor U8297 (N_8297,N_8105,N_8171);
nand U8298 (N_8298,N_7922,N_7661);
or U8299 (N_8299,N_7549,N_7895);
xor U8300 (N_8300,N_7674,N_8110);
xnor U8301 (N_8301,N_7938,N_7695);
nor U8302 (N_8302,N_7951,N_7788);
nand U8303 (N_8303,N_7948,N_7744);
nand U8304 (N_8304,N_7865,N_7774);
or U8305 (N_8305,N_8234,N_7842);
and U8306 (N_8306,N_7721,N_8051);
xnor U8307 (N_8307,N_7741,N_8071);
xnor U8308 (N_8308,N_7656,N_7987);
nand U8309 (N_8309,N_7905,N_8164);
nor U8310 (N_8310,N_8072,N_8173);
nand U8311 (N_8311,N_7667,N_7501);
or U8312 (N_8312,N_8163,N_8213);
xor U8313 (N_8313,N_8249,N_8206);
or U8314 (N_8314,N_8134,N_8232);
nor U8315 (N_8315,N_7848,N_7599);
xor U8316 (N_8316,N_7808,N_7626);
or U8317 (N_8317,N_8174,N_8111);
xnor U8318 (N_8318,N_8066,N_7748);
xnor U8319 (N_8319,N_7804,N_8060);
nand U8320 (N_8320,N_7699,N_7720);
nand U8321 (N_8321,N_7864,N_7574);
and U8322 (N_8322,N_8224,N_7533);
xor U8323 (N_8323,N_7725,N_7600);
nor U8324 (N_8324,N_7986,N_7588);
and U8325 (N_8325,N_8052,N_8245);
nand U8326 (N_8326,N_7798,N_7632);
or U8327 (N_8327,N_7939,N_7563);
or U8328 (N_8328,N_7861,N_7970);
or U8329 (N_8329,N_8199,N_7913);
xor U8330 (N_8330,N_7735,N_7594);
and U8331 (N_8331,N_7733,N_8119);
nor U8332 (N_8332,N_7634,N_7572);
or U8333 (N_8333,N_8063,N_8074);
and U8334 (N_8334,N_7648,N_7751);
nand U8335 (N_8335,N_7686,N_8186);
or U8336 (N_8336,N_7871,N_7955);
and U8337 (N_8337,N_7985,N_8028);
xnor U8338 (N_8338,N_7924,N_7994);
nor U8339 (N_8339,N_7631,N_7571);
nand U8340 (N_8340,N_7583,N_7952);
or U8341 (N_8341,N_7564,N_8038);
nand U8342 (N_8342,N_7920,N_7585);
nand U8343 (N_8343,N_8065,N_7666);
nand U8344 (N_8344,N_7612,N_7535);
xor U8345 (N_8345,N_8219,N_8160);
xnor U8346 (N_8346,N_7873,N_7511);
and U8347 (N_8347,N_7543,N_8142);
nor U8348 (N_8348,N_7579,N_7567);
xor U8349 (N_8349,N_8020,N_7542);
xnor U8350 (N_8350,N_7693,N_7797);
and U8351 (N_8351,N_7603,N_7615);
nand U8352 (N_8352,N_8197,N_7655);
nor U8353 (N_8353,N_8240,N_8183);
nand U8354 (N_8354,N_8013,N_8033);
nand U8355 (N_8355,N_7541,N_7709);
or U8356 (N_8356,N_7687,N_8144);
or U8357 (N_8357,N_7890,N_8169);
nor U8358 (N_8358,N_7738,N_7618);
xnor U8359 (N_8359,N_7814,N_8089);
nand U8360 (N_8360,N_8040,N_8178);
and U8361 (N_8361,N_7730,N_7556);
and U8362 (N_8362,N_7880,N_7944);
and U8363 (N_8363,N_7624,N_7749);
xor U8364 (N_8364,N_8137,N_8205);
xor U8365 (N_8365,N_7795,N_7805);
and U8366 (N_8366,N_7647,N_8154);
or U8367 (N_8367,N_7881,N_7607);
nand U8368 (N_8368,N_8136,N_7587);
nand U8369 (N_8369,N_8123,N_8050);
xnor U8370 (N_8370,N_8182,N_7816);
or U8371 (N_8371,N_7654,N_7557);
or U8372 (N_8372,N_7975,N_8076);
nor U8373 (N_8373,N_7806,N_8068);
nand U8374 (N_8374,N_8218,N_8228);
or U8375 (N_8375,N_8189,N_7840);
and U8376 (N_8376,N_7900,N_7803);
nor U8377 (N_8377,N_7991,N_7815);
nor U8378 (N_8378,N_8188,N_8106);
nor U8379 (N_8379,N_8193,N_8044);
nand U8380 (N_8380,N_8203,N_7979);
xnor U8381 (N_8381,N_7857,N_7560);
nand U8382 (N_8382,N_7653,N_7649);
and U8383 (N_8383,N_8034,N_7545);
nand U8384 (N_8384,N_7812,N_8048);
xor U8385 (N_8385,N_8156,N_7909);
or U8386 (N_8386,N_7663,N_7945);
and U8387 (N_8387,N_7982,N_7573);
or U8388 (N_8388,N_7824,N_8147);
and U8389 (N_8389,N_7810,N_8177);
or U8390 (N_8390,N_7536,N_8025);
or U8391 (N_8391,N_7903,N_8039);
nand U8392 (N_8392,N_7767,N_8128);
nand U8393 (N_8393,N_7616,N_8130);
or U8394 (N_8394,N_7604,N_7937);
nand U8395 (N_8395,N_7553,N_7623);
nor U8396 (N_8396,N_7775,N_7879);
or U8397 (N_8397,N_8056,N_8126);
or U8398 (N_8398,N_7681,N_7526);
or U8399 (N_8399,N_8057,N_7581);
and U8400 (N_8400,N_8018,N_7690);
nor U8401 (N_8401,N_7736,N_7839);
and U8402 (N_8402,N_7800,N_8236);
xnor U8403 (N_8403,N_7969,N_7592);
and U8404 (N_8404,N_7908,N_7852);
or U8405 (N_8405,N_8198,N_8204);
nor U8406 (N_8406,N_8209,N_7811);
nand U8407 (N_8407,N_7792,N_7988);
or U8408 (N_8408,N_8062,N_7717);
and U8409 (N_8409,N_8008,N_7566);
xor U8410 (N_8410,N_7701,N_8227);
nor U8411 (N_8411,N_7974,N_7697);
nor U8412 (N_8412,N_7562,N_8093);
nor U8413 (N_8413,N_7910,N_7700);
or U8414 (N_8414,N_7746,N_8006);
nand U8415 (N_8415,N_7949,N_8027);
and U8416 (N_8416,N_8102,N_8166);
or U8417 (N_8417,N_7959,N_7659);
nor U8418 (N_8418,N_7796,N_7635);
or U8419 (N_8419,N_7941,N_7515);
nand U8420 (N_8420,N_7818,N_7828);
xor U8421 (N_8421,N_7911,N_7546);
or U8422 (N_8422,N_7621,N_8181);
and U8423 (N_8423,N_7523,N_7928);
and U8424 (N_8424,N_7966,N_8015);
nor U8425 (N_8425,N_8041,N_8022);
xnor U8426 (N_8426,N_8101,N_8082);
nand U8427 (N_8427,N_7645,N_8139);
nor U8428 (N_8428,N_7844,N_8127);
nand U8429 (N_8429,N_7633,N_7714);
nand U8430 (N_8430,N_7896,N_7544);
xor U8431 (N_8431,N_8109,N_8148);
or U8432 (N_8432,N_7559,N_7826);
nand U8433 (N_8433,N_8248,N_7643);
nand U8434 (N_8434,N_8014,N_7539);
or U8435 (N_8435,N_7813,N_7727);
nand U8436 (N_8436,N_7694,N_7930);
and U8437 (N_8437,N_7750,N_7902);
and U8438 (N_8438,N_7505,N_8229);
and U8439 (N_8439,N_8094,N_7677);
xnor U8440 (N_8440,N_8241,N_8042);
xor U8441 (N_8441,N_8059,N_8045);
xnor U8442 (N_8442,N_8084,N_7779);
nor U8443 (N_8443,N_7981,N_7682);
and U8444 (N_8444,N_8221,N_7520);
nor U8445 (N_8445,N_8216,N_8046);
xnor U8446 (N_8446,N_8244,N_7547);
and U8447 (N_8447,N_8149,N_7680);
xor U8448 (N_8448,N_7799,N_7646);
nand U8449 (N_8449,N_7943,N_8131);
nor U8450 (N_8450,N_7718,N_7827);
or U8451 (N_8451,N_8067,N_7829);
nand U8452 (N_8452,N_7715,N_7926);
or U8453 (N_8453,N_7503,N_7888);
and U8454 (N_8454,N_7538,N_7561);
and U8455 (N_8455,N_8187,N_7785);
or U8456 (N_8456,N_7691,N_8212);
or U8457 (N_8457,N_7847,N_7833);
nand U8458 (N_8458,N_8230,N_8030);
xor U8459 (N_8459,N_7897,N_8200);
and U8460 (N_8460,N_7942,N_8007);
nor U8461 (N_8461,N_7917,N_7953);
xor U8462 (N_8462,N_8242,N_7894);
and U8463 (N_8463,N_8246,N_8153);
or U8464 (N_8464,N_7783,N_7664);
nand U8465 (N_8465,N_7899,N_7790);
or U8466 (N_8466,N_8035,N_8165);
nor U8467 (N_8467,N_7884,N_7644);
or U8468 (N_8468,N_7639,N_7999);
nand U8469 (N_8469,N_8024,N_7867);
or U8470 (N_8470,N_7919,N_7898);
or U8471 (N_8471,N_7688,N_7605);
xnor U8472 (N_8472,N_8210,N_8112);
xnor U8473 (N_8473,N_7802,N_8003);
nand U8474 (N_8474,N_7660,N_8092);
nor U8475 (N_8475,N_7791,N_7784);
nand U8476 (N_8476,N_7555,N_7957);
nand U8477 (N_8477,N_7956,N_7935);
nand U8478 (N_8478,N_7753,N_7914);
xnor U8479 (N_8479,N_8180,N_7502);
and U8480 (N_8480,N_7836,N_7512);
or U8481 (N_8481,N_7958,N_7755);
nor U8482 (N_8482,N_7763,N_8087);
nand U8483 (N_8483,N_8053,N_7596);
nand U8484 (N_8484,N_7859,N_7777);
or U8485 (N_8485,N_7617,N_7886);
nand U8486 (N_8486,N_8151,N_8049);
and U8487 (N_8487,N_7540,N_7773);
or U8488 (N_8488,N_7641,N_7521);
xnor U8489 (N_8489,N_8167,N_8202);
nor U8490 (N_8490,N_7613,N_7670);
nor U8491 (N_8491,N_7837,N_7807);
xor U8492 (N_8492,N_8070,N_8088);
nand U8493 (N_8493,N_7877,N_7996);
nor U8494 (N_8494,N_7619,N_7787);
and U8495 (N_8495,N_8222,N_8168);
nor U8496 (N_8496,N_8031,N_7876);
or U8497 (N_8497,N_8208,N_8114);
xnor U8498 (N_8498,N_7923,N_7780);
xor U8499 (N_8499,N_7927,N_7739);
xor U8500 (N_8500,N_7734,N_8125);
and U8501 (N_8501,N_7967,N_8129);
xnor U8502 (N_8502,N_7609,N_7866);
or U8503 (N_8503,N_7954,N_7834);
and U8504 (N_8504,N_7793,N_7554);
nand U8505 (N_8505,N_7983,N_8017);
and U8506 (N_8506,N_7673,N_7723);
nand U8507 (N_8507,N_8002,N_7569);
nor U8508 (N_8508,N_7964,N_8009);
nand U8509 (N_8509,N_7870,N_7855);
xnor U8510 (N_8510,N_7965,N_7610);
and U8511 (N_8511,N_7912,N_8201);
or U8512 (N_8512,N_8217,N_7684);
and U8513 (N_8513,N_8037,N_7929);
xor U8514 (N_8514,N_8124,N_8226);
nor U8515 (N_8515,N_8077,N_8215);
nor U8516 (N_8516,N_7838,N_7568);
nand U8517 (N_8517,N_7671,N_7851);
xor U8518 (N_8518,N_7758,N_8081);
and U8519 (N_8519,N_7668,N_8150);
nor U8520 (N_8520,N_7931,N_7713);
nand U8521 (N_8521,N_7901,N_8073);
nand U8522 (N_8522,N_7933,N_7591);
and U8523 (N_8523,N_7683,N_7704);
xor U8524 (N_8524,N_7747,N_8104);
xnor U8525 (N_8525,N_8161,N_7845);
nand U8526 (N_8526,N_7760,N_8005);
or U8527 (N_8527,N_7524,N_8145);
nor U8528 (N_8528,N_8157,N_7891);
xnor U8529 (N_8529,N_8107,N_7752);
or U8530 (N_8530,N_7629,N_7578);
nand U8531 (N_8531,N_8141,N_8090);
nand U8532 (N_8532,N_8085,N_7706);
and U8533 (N_8533,N_7710,N_7830);
xor U8534 (N_8534,N_7854,N_8140);
nor U8535 (N_8535,N_8026,N_8103);
nor U8536 (N_8536,N_8225,N_7885);
nand U8537 (N_8537,N_8184,N_7728);
nor U8538 (N_8538,N_7657,N_8192);
nand U8539 (N_8539,N_7577,N_7962);
and U8540 (N_8540,N_7582,N_8023);
nor U8541 (N_8541,N_8135,N_8121);
nand U8542 (N_8542,N_7817,N_7507);
nand U8543 (N_8543,N_7625,N_7835);
nor U8544 (N_8544,N_7925,N_7669);
nor U8545 (N_8545,N_7640,N_8095);
nand U8546 (N_8546,N_8099,N_7513);
xnor U8547 (N_8547,N_8191,N_7602);
nor U8548 (N_8548,N_7548,N_7608);
nor U8549 (N_8549,N_7702,N_8247);
nor U8550 (N_8550,N_7689,N_7576);
or U8551 (N_8551,N_8235,N_7820);
or U8552 (N_8552,N_8237,N_7665);
xor U8553 (N_8553,N_8113,N_7650);
nor U8554 (N_8554,N_7525,N_7940);
xor U8555 (N_8555,N_7638,N_7771);
and U8556 (N_8556,N_7627,N_7892);
nor U8557 (N_8557,N_8012,N_7794);
nand U8558 (N_8558,N_7737,N_7825);
xnor U8559 (N_8559,N_7823,N_7950);
nand U8560 (N_8560,N_8054,N_8097);
and U8561 (N_8561,N_7584,N_7765);
or U8562 (N_8562,N_7869,N_7522);
or U8563 (N_8563,N_8122,N_7882);
and U8564 (N_8564,N_7530,N_7696);
nand U8565 (N_8565,N_7756,N_7801);
and U8566 (N_8566,N_8231,N_7732);
xor U8567 (N_8567,N_8047,N_7685);
or U8568 (N_8568,N_7651,N_7972);
xnor U8569 (N_8569,N_8061,N_8100);
xor U8570 (N_8570,N_7989,N_8233);
nand U8571 (N_8571,N_8158,N_7570);
nand U8572 (N_8572,N_8011,N_8016);
xor U8573 (N_8573,N_7754,N_7893);
xnor U8574 (N_8574,N_7506,N_7973);
nor U8575 (N_8575,N_8143,N_8010);
or U8576 (N_8576,N_8172,N_7628);
nor U8577 (N_8577,N_7593,N_7601);
xnor U8578 (N_8578,N_8019,N_8243);
nand U8579 (N_8579,N_8118,N_8159);
and U8580 (N_8580,N_8091,N_7726);
nor U8581 (N_8581,N_7679,N_7662);
nand U8582 (N_8582,N_7630,N_8207);
or U8583 (N_8583,N_7698,N_7872);
and U8584 (N_8584,N_7676,N_7887);
or U8585 (N_8585,N_7976,N_7769);
and U8586 (N_8586,N_7946,N_7997);
nor U8587 (N_8587,N_7850,N_8146);
nand U8588 (N_8588,N_7761,N_7984);
xor U8589 (N_8589,N_7575,N_7977);
nand U8590 (N_8590,N_8211,N_7980);
nor U8591 (N_8591,N_7934,N_7703);
nand U8592 (N_8592,N_7889,N_7672);
nor U8593 (N_8593,N_8176,N_7532);
or U8594 (N_8594,N_7781,N_7766);
nor U8595 (N_8595,N_7528,N_8223);
xor U8596 (N_8596,N_8080,N_7776);
xnor U8597 (N_8597,N_7534,N_7936);
or U8598 (N_8598,N_7858,N_8086);
xor U8599 (N_8599,N_7759,N_8064);
nand U8600 (N_8600,N_8214,N_8043);
xnor U8601 (N_8601,N_8083,N_8239);
xor U8602 (N_8602,N_7590,N_7652);
or U8603 (N_8603,N_8069,N_7724);
nand U8604 (N_8604,N_7586,N_7770);
nor U8605 (N_8605,N_7998,N_7731);
and U8606 (N_8606,N_8055,N_8238);
and U8607 (N_8607,N_8078,N_7778);
or U8608 (N_8608,N_7883,N_8117);
or U8609 (N_8609,N_7516,N_7552);
xor U8610 (N_8610,N_7878,N_7637);
xor U8611 (N_8611,N_7614,N_7716);
nor U8612 (N_8612,N_7995,N_8194);
and U8613 (N_8613,N_7551,N_7711);
nor U8614 (N_8614,N_7518,N_8000);
or U8615 (N_8615,N_7514,N_7764);
nand U8616 (N_8616,N_7519,N_7971);
xor U8617 (N_8617,N_7620,N_7675);
and U8618 (N_8618,N_7500,N_7907);
nor U8619 (N_8619,N_8075,N_7918);
nor U8620 (N_8620,N_8175,N_8133);
nand U8621 (N_8621,N_7580,N_7915);
or U8622 (N_8622,N_7517,N_7708);
or U8623 (N_8623,N_7722,N_8096);
xnor U8624 (N_8624,N_7916,N_7537);
nor U8625 (N_8625,N_7723,N_7996);
and U8626 (N_8626,N_7646,N_8047);
xor U8627 (N_8627,N_7763,N_7560);
nor U8628 (N_8628,N_7584,N_7994);
xor U8629 (N_8629,N_8068,N_7815);
nand U8630 (N_8630,N_8244,N_8161);
and U8631 (N_8631,N_8110,N_8171);
nor U8632 (N_8632,N_8102,N_7832);
xor U8633 (N_8633,N_8146,N_7505);
and U8634 (N_8634,N_7906,N_7563);
nor U8635 (N_8635,N_8058,N_7573);
and U8636 (N_8636,N_7668,N_7575);
nand U8637 (N_8637,N_7922,N_7572);
nand U8638 (N_8638,N_8165,N_7919);
nor U8639 (N_8639,N_7855,N_8209);
nor U8640 (N_8640,N_7915,N_7663);
xnor U8641 (N_8641,N_7555,N_7630);
and U8642 (N_8642,N_8188,N_7878);
or U8643 (N_8643,N_7617,N_7772);
and U8644 (N_8644,N_7650,N_8060);
xor U8645 (N_8645,N_7864,N_7653);
xnor U8646 (N_8646,N_8137,N_7616);
nand U8647 (N_8647,N_7860,N_7621);
and U8648 (N_8648,N_8205,N_8215);
and U8649 (N_8649,N_8106,N_8011);
nor U8650 (N_8650,N_7513,N_7520);
or U8651 (N_8651,N_8150,N_7537);
and U8652 (N_8652,N_8046,N_7715);
nand U8653 (N_8653,N_8219,N_8005);
or U8654 (N_8654,N_7984,N_7833);
nor U8655 (N_8655,N_7842,N_8084);
or U8656 (N_8656,N_7959,N_7605);
nor U8657 (N_8657,N_8007,N_7967);
xnor U8658 (N_8658,N_8136,N_7800);
xor U8659 (N_8659,N_7765,N_7712);
and U8660 (N_8660,N_7758,N_7938);
and U8661 (N_8661,N_7549,N_7694);
xnor U8662 (N_8662,N_8108,N_8175);
and U8663 (N_8663,N_8180,N_8046);
xnor U8664 (N_8664,N_7996,N_7670);
xnor U8665 (N_8665,N_8234,N_8010);
xor U8666 (N_8666,N_8036,N_7961);
xor U8667 (N_8667,N_8166,N_7934);
xnor U8668 (N_8668,N_7788,N_7990);
and U8669 (N_8669,N_8013,N_7524);
nor U8670 (N_8670,N_7732,N_7855);
and U8671 (N_8671,N_7566,N_7887);
xnor U8672 (N_8672,N_8123,N_7917);
nor U8673 (N_8673,N_8082,N_8031);
xor U8674 (N_8674,N_8109,N_8067);
and U8675 (N_8675,N_7576,N_7641);
xor U8676 (N_8676,N_8102,N_8089);
and U8677 (N_8677,N_7981,N_7582);
xnor U8678 (N_8678,N_7731,N_8118);
and U8679 (N_8679,N_7695,N_7697);
and U8680 (N_8680,N_7751,N_8014);
nand U8681 (N_8681,N_8116,N_8118);
nor U8682 (N_8682,N_7658,N_7877);
xor U8683 (N_8683,N_7665,N_7807);
xnor U8684 (N_8684,N_7704,N_8209);
and U8685 (N_8685,N_7726,N_7803);
nand U8686 (N_8686,N_7848,N_7782);
or U8687 (N_8687,N_8112,N_7502);
nor U8688 (N_8688,N_7928,N_7637);
xor U8689 (N_8689,N_7977,N_8112);
and U8690 (N_8690,N_7560,N_7511);
or U8691 (N_8691,N_7502,N_7553);
nand U8692 (N_8692,N_8083,N_8093);
xor U8693 (N_8693,N_7730,N_7518);
and U8694 (N_8694,N_7824,N_8208);
xor U8695 (N_8695,N_8178,N_7625);
nand U8696 (N_8696,N_7697,N_8200);
nand U8697 (N_8697,N_7786,N_7838);
nand U8698 (N_8698,N_8223,N_8067);
and U8699 (N_8699,N_7576,N_7812);
or U8700 (N_8700,N_8235,N_7844);
nand U8701 (N_8701,N_7670,N_7852);
xor U8702 (N_8702,N_7949,N_8065);
xnor U8703 (N_8703,N_7509,N_8248);
nor U8704 (N_8704,N_7652,N_7819);
or U8705 (N_8705,N_7760,N_8161);
and U8706 (N_8706,N_7905,N_7765);
and U8707 (N_8707,N_7866,N_7723);
xnor U8708 (N_8708,N_8228,N_7794);
and U8709 (N_8709,N_8103,N_7652);
xnor U8710 (N_8710,N_8011,N_7813);
or U8711 (N_8711,N_7812,N_8013);
and U8712 (N_8712,N_7891,N_7998);
or U8713 (N_8713,N_7774,N_7630);
or U8714 (N_8714,N_7650,N_7542);
and U8715 (N_8715,N_7853,N_7905);
nor U8716 (N_8716,N_7939,N_8187);
xor U8717 (N_8717,N_8126,N_7867);
and U8718 (N_8718,N_7760,N_7953);
or U8719 (N_8719,N_7531,N_8057);
nand U8720 (N_8720,N_8167,N_7608);
and U8721 (N_8721,N_8047,N_8193);
nand U8722 (N_8722,N_7699,N_7965);
or U8723 (N_8723,N_8037,N_8010);
nor U8724 (N_8724,N_7697,N_7854);
or U8725 (N_8725,N_7851,N_7922);
nand U8726 (N_8726,N_8091,N_7966);
nand U8727 (N_8727,N_8004,N_7730);
or U8728 (N_8728,N_7742,N_7997);
or U8729 (N_8729,N_8214,N_8031);
xnor U8730 (N_8730,N_7919,N_8181);
or U8731 (N_8731,N_7832,N_8045);
nor U8732 (N_8732,N_7746,N_7798);
nand U8733 (N_8733,N_7569,N_7930);
nor U8734 (N_8734,N_8243,N_7764);
nor U8735 (N_8735,N_7873,N_7640);
and U8736 (N_8736,N_7698,N_7757);
or U8737 (N_8737,N_7863,N_7702);
and U8738 (N_8738,N_7679,N_8117);
nor U8739 (N_8739,N_7626,N_8106);
and U8740 (N_8740,N_7839,N_8005);
and U8741 (N_8741,N_7541,N_7506);
xor U8742 (N_8742,N_7609,N_7627);
nor U8743 (N_8743,N_7853,N_7678);
xnor U8744 (N_8744,N_8206,N_7566);
nor U8745 (N_8745,N_7735,N_7649);
or U8746 (N_8746,N_8064,N_8045);
or U8747 (N_8747,N_7810,N_7919);
nor U8748 (N_8748,N_8173,N_8042);
and U8749 (N_8749,N_7685,N_7537);
nand U8750 (N_8750,N_8167,N_7616);
nor U8751 (N_8751,N_7657,N_7879);
or U8752 (N_8752,N_7961,N_7662);
and U8753 (N_8753,N_7790,N_7931);
nor U8754 (N_8754,N_7544,N_8088);
or U8755 (N_8755,N_7686,N_7543);
xnor U8756 (N_8756,N_8232,N_7999);
xnor U8757 (N_8757,N_7995,N_7958);
and U8758 (N_8758,N_8197,N_7795);
or U8759 (N_8759,N_7942,N_7595);
or U8760 (N_8760,N_8112,N_7916);
and U8761 (N_8761,N_8218,N_8068);
nand U8762 (N_8762,N_7687,N_7866);
nand U8763 (N_8763,N_7852,N_7944);
nor U8764 (N_8764,N_8004,N_7717);
nand U8765 (N_8765,N_8200,N_7961);
and U8766 (N_8766,N_7526,N_7925);
xnor U8767 (N_8767,N_7729,N_8238);
and U8768 (N_8768,N_7908,N_7812);
and U8769 (N_8769,N_7904,N_7625);
nor U8770 (N_8770,N_7756,N_8154);
xnor U8771 (N_8771,N_7966,N_8210);
nor U8772 (N_8772,N_7930,N_8149);
xor U8773 (N_8773,N_8002,N_7817);
or U8774 (N_8774,N_7931,N_7580);
nor U8775 (N_8775,N_7945,N_7643);
nand U8776 (N_8776,N_8128,N_7575);
nor U8777 (N_8777,N_7780,N_8087);
or U8778 (N_8778,N_7815,N_7819);
nand U8779 (N_8779,N_8076,N_8007);
nand U8780 (N_8780,N_7542,N_7800);
or U8781 (N_8781,N_7620,N_8058);
nand U8782 (N_8782,N_8047,N_7931);
nand U8783 (N_8783,N_7744,N_8039);
nand U8784 (N_8784,N_7628,N_7897);
nand U8785 (N_8785,N_8183,N_7599);
or U8786 (N_8786,N_7546,N_8145);
nor U8787 (N_8787,N_8221,N_8001);
and U8788 (N_8788,N_7723,N_7949);
nor U8789 (N_8789,N_7535,N_7905);
xor U8790 (N_8790,N_8129,N_7980);
or U8791 (N_8791,N_8205,N_8122);
or U8792 (N_8792,N_7510,N_7875);
xor U8793 (N_8793,N_7657,N_7842);
xnor U8794 (N_8794,N_7944,N_7732);
nor U8795 (N_8795,N_7953,N_7719);
nand U8796 (N_8796,N_7655,N_8026);
nand U8797 (N_8797,N_8146,N_8077);
or U8798 (N_8798,N_7645,N_7924);
xor U8799 (N_8799,N_8148,N_7969);
nand U8800 (N_8800,N_7614,N_8188);
nor U8801 (N_8801,N_7979,N_7531);
nand U8802 (N_8802,N_7869,N_7880);
or U8803 (N_8803,N_7900,N_8198);
or U8804 (N_8804,N_8126,N_8059);
xor U8805 (N_8805,N_7554,N_8069);
xnor U8806 (N_8806,N_7502,N_8086);
nor U8807 (N_8807,N_7732,N_7878);
and U8808 (N_8808,N_7891,N_7731);
nand U8809 (N_8809,N_7965,N_7738);
xor U8810 (N_8810,N_7644,N_7769);
and U8811 (N_8811,N_7529,N_7564);
nand U8812 (N_8812,N_7724,N_8228);
and U8813 (N_8813,N_7767,N_8024);
and U8814 (N_8814,N_7827,N_7828);
xor U8815 (N_8815,N_8039,N_7559);
nor U8816 (N_8816,N_8226,N_7769);
nand U8817 (N_8817,N_8101,N_7652);
and U8818 (N_8818,N_7865,N_7848);
or U8819 (N_8819,N_7686,N_7847);
or U8820 (N_8820,N_7649,N_8194);
and U8821 (N_8821,N_7854,N_8000);
xnor U8822 (N_8822,N_8246,N_7798);
nor U8823 (N_8823,N_7963,N_8032);
nor U8824 (N_8824,N_7932,N_7904);
nor U8825 (N_8825,N_7586,N_8185);
or U8826 (N_8826,N_8144,N_7637);
xor U8827 (N_8827,N_8112,N_7701);
nor U8828 (N_8828,N_7610,N_8120);
and U8829 (N_8829,N_8127,N_7752);
or U8830 (N_8830,N_7880,N_7567);
and U8831 (N_8831,N_8117,N_8064);
or U8832 (N_8832,N_7526,N_7781);
nor U8833 (N_8833,N_7749,N_8140);
and U8834 (N_8834,N_7773,N_8207);
nor U8835 (N_8835,N_8126,N_7508);
or U8836 (N_8836,N_8104,N_7688);
xnor U8837 (N_8837,N_7957,N_8229);
nor U8838 (N_8838,N_7958,N_7726);
nor U8839 (N_8839,N_7905,N_7759);
xor U8840 (N_8840,N_7506,N_7570);
xnor U8841 (N_8841,N_7632,N_8240);
or U8842 (N_8842,N_8156,N_8007);
or U8843 (N_8843,N_7799,N_8031);
and U8844 (N_8844,N_8233,N_8182);
or U8845 (N_8845,N_8119,N_8146);
xnor U8846 (N_8846,N_7517,N_7997);
nand U8847 (N_8847,N_7851,N_7609);
or U8848 (N_8848,N_7862,N_7939);
xnor U8849 (N_8849,N_7569,N_7863);
xnor U8850 (N_8850,N_7535,N_7730);
xnor U8851 (N_8851,N_8205,N_7690);
nand U8852 (N_8852,N_7523,N_7734);
nand U8853 (N_8853,N_8183,N_8035);
nor U8854 (N_8854,N_7643,N_8068);
nor U8855 (N_8855,N_7664,N_7960);
or U8856 (N_8856,N_7735,N_8170);
nor U8857 (N_8857,N_8180,N_7764);
nand U8858 (N_8858,N_8214,N_8065);
and U8859 (N_8859,N_7878,N_8094);
nand U8860 (N_8860,N_8023,N_8107);
nor U8861 (N_8861,N_8059,N_7855);
or U8862 (N_8862,N_7957,N_7656);
nor U8863 (N_8863,N_7814,N_7957);
nand U8864 (N_8864,N_7973,N_7597);
nor U8865 (N_8865,N_7877,N_7872);
nand U8866 (N_8866,N_8016,N_8079);
and U8867 (N_8867,N_7959,N_7670);
nand U8868 (N_8868,N_7705,N_8117);
or U8869 (N_8869,N_7914,N_7653);
or U8870 (N_8870,N_7592,N_8026);
and U8871 (N_8871,N_7514,N_7843);
or U8872 (N_8872,N_7594,N_8092);
xor U8873 (N_8873,N_7822,N_7553);
nand U8874 (N_8874,N_7725,N_7724);
and U8875 (N_8875,N_7829,N_7963);
xnor U8876 (N_8876,N_8167,N_7614);
nor U8877 (N_8877,N_7901,N_8060);
or U8878 (N_8878,N_7992,N_7808);
nor U8879 (N_8879,N_7518,N_7771);
nand U8880 (N_8880,N_7639,N_8100);
xnor U8881 (N_8881,N_7697,N_7841);
nand U8882 (N_8882,N_7869,N_8089);
or U8883 (N_8883,N_7523,N_7525);
nor U8884 (N_8884,N_8085,N_7624);
xor U8885 (N_8885,N_7978,N_8108);
nor U8886 (N_8886,N_7737,N_7635);
and U8887 (N_8887,N_7849,N_7757);
and U8888 (N_8888,N_7900,N_7819);
nand U8889 (N_8889,N_7892,N_7980);
nand U8890 (N_8890,N_7747,N_7534);
or U8891 (N_8891,N_7748,N_8140);
nand U8892 (N_8892,N_8161,N_7875);
nor U8893 (N_8893,N_8174,N_7630);
xor U8894 (N_8894,N_7566,N_8014);
xor U8895 (N_8895,N_7740,N_7779);
nand U8896 (N_8896,N_7588,N_7940);
or U8897 (N_8897,N_7922,N_8158);
and U8898 (N_8898,N_7552,N_7536);
or U8899 (N_8899,N_8083,N_7530);
or U8900 (N_8900,N_7647,N_7755);
nand U8901 (N_8901,N_7660,N_7537);
or U8902 (N_8902,N_7955,N_8120);
or U8903 (N_8903,N_7792,N_8064);
xnor U8904 (N_8904,N_7548,N_7946);
nor U8905 (N_8905,N_8006,N_8076);
xor U8906 (N_8906,N_7891,N_7651);
nor U8907 (N_8907,N_7919,N_8051);
nand U8908 (N_8908,N_7888,N_7723);
xor U8909 (N_8909,N_7721,N_7837);
nor U8910 (N_8910,N_7886,N_8019);
nand U8911 (N_8911,N_8085,N_7560);
xnor U8912 (N_8912,N_8147,N_7552);
nor U8913 (N_8913,N_7752,N_7854);
or U8914 (N_8914,N_8237,N_7654);
nor U8915 (N_8915,N_7632,N_7920);
xor U8916 (N_8916,N_8145,N_8067);
and U8917 (N_8917,N_7859,N_8192);
or U8918 (N_8918,N_7626,N_8245);
and U8919 (N_8919,N_8099,N_7607);
nor U8920 (N_8920,N_8008,N_7954);
and U8921 (N_8921,N_8112,N_7929);
xor U8922 (N_8922,N_7880,N_7810);
xor U8923 (N_8923,N_7584,N_7728);
nor U8924 (N_8924,N_8196,N_7680);
nor U8925 (N_8925,N_7566,N_7540);
xnor U8926 (N_8926,N_8068,N_7571);
xor U8927 (N_8927,N_8053,N_8000);
nand U8928 (N_8928,N_7842,N_7663);
or U8929 (N_8929,N_7691,N_8023);
and U8930 (N_8930,N_7774,N_7582);
or U8931 (N_8931,N_7511,N_7846);
xor U8932 (N_8932,N_8179,N_8039);
nand U8933 (N_8933,N_8092,N_7683);
xnor U8934 (N_8934,N_8234,N_8033);
and U8935 (N_8935,N_7539,N_8060);
xnor U8936 (N_8936,N_7553,N_7639);
nor U8937 (N_8937,N_7561,N_7954);
nor U8938 (N_8938,N_8019,N_7826);
nand U8939 (N_8939,N_7578,N_7890);
or U8940 (N_8940,N_8106,N_7510);
nand U8941 (N_8941,N_7829,N_7593);
xor U8942 (N_8942,N_7655,N_7819);
xor U8943 (N_8943,N_7739,N_7628);
nand U8944 (N_8944,N_7725,N_7980);
nor U8945 (N_8945,N_8163,N_8170);
xor U8946 (N_8946,N_8021,N_8226);
and U8947 (N_8947,N_8019,N_7783);
xor U8948 (N_8948,N_8188,N_8097);
xor U8949 (N_8949,N_7847,N_7992);
or U8950 (N_8950,N_8105,N_8088);
xor U8951 (N_8951,N_8132,N_7985);
nor U8952 (N_8952,N_7823,N_8165);
and U8953 (N_8953,N_7978,N_7623);
nand U8954 (N_8954,N_8091,N_7548);
nand U8955 (N_8955,N_7737,N_7888);
nand U8956 (N_8956,N_8226,N_7718);
nand U8957 (N_8957,N_7509,N_8070);
and U8958 (N_8958,N_7584,N_7911);
nor U8959 (N_8959,N_7662,N_7858);
nand U8960 (N_8960,N_7994,N_7788);
or U8961 (N_8961,N_8054,N_7730);
nor U8962 (N_8962,N_8213,N_7705);
and U8963 (N_8963,N_8106,N_7985);
nand U8964 (N_8964,N_7540,N_8042);
or U8965 (N_8965,N_7981,N_7508);
nor U8966 (N_8966,N_7597,N_8174);
and U8967 (N_8967,N_7512,N_8018);
or U8968 (N_8968,N_7697,N_7931);
nand U8969 (N_8969,N_7500,N_7710);
nand U8970 (N_8970,N_7985,N_7833);
and U8971 (N_8971,N_7755,N_7776);
nor U8972 (N_8972,N_8140,N_7979);
or U8973 (N_8973,N_8223,N_7899);
and U8974 (N_8974,N_8229,N_7851);
and U8975 (N_8975,N_8121,N_7940);
nor U8976 (N_8976,N_7895,N_8232);
nand U8977 (N_8977,N_7560,N_7970);
xor U8978 (N_8978,N_7804,N_7704);
and U8979 (N_8979,N_7984,N_8159);
and U8980 (N_8980,N_8013,N_7963);
nand U8981 (N_8981,N_7938,N_7747);
nand U8982 (N_8982,N_8111,N_8034);
nor U8983 (N_8983,N_7853,N_7751);
nand U8984 (N_8984,N_8147,N_8026);
and U8985 (N_8985,N_8226,N_7764);
and U8986 (N_8986,N_8211,N_8142);
xor U8987 (N_8987,N_8063,N_8104);
nor U8988 (N_8988,N_7535,N_7944);
nor U8989 (N_8989,N_8007,N_7551);
or U8990 (N_8990,N_7545,N_7739);
and U8991 (N_8991,N_7839,N_8104);
nor U8992 (N_8992,N_8170,N_7808);
nand U8993 (N_8993,N_7531,N_7549);
nand U8994 (N_8994,N_7908,N_8068);
nor U8995 (N_8995,N_8141,N_8205);
nor U8996 (N_8996,N_8035,N_8185);
nand U8997 (N_8997,N_8049,N_7972);
or U8998 (N_8998,N_7508,N_7928);
nor U8999 (N_8999,N_7686,N_7774);
nor U9000 (N_9000,N_8366,N_8945);
and U9001 (N_9001,N_8956,N_8560);
or U9002 (N_9002,N_8903,N_8740);
or U9003 (N_9003,N_8969,N_8389);
nand U9004 (N_9004,N_8306,N_8805);
and U9005 (N_9005,N_8877,N_8581);
or U9006 (N_9006,N_8619,N_8975);
or U9007 (N_9007,N_8984,N_8898);
nor U9008 (N_9008,N_8441,N_8386);
or U9009 (N_9009,N_8497,N_8551);
or U9010 (N_9010,N_8342,N_8841);
nor U9011 (N_9011,N_8762,N_8326);
or U9012 (N_9012,N_8630,N_8746);
nand U9013 (N_9013,N_8256,N_8666);
and U9014 (N_9014,N_8530,N_8252);
or U9015 (N_9015,N_8862,N_8612);
and U9016 (N_9016,N_8960,N_8568);
nand U9017 (N_9017,N_8345,N_8873);
and U9018 (N_9018,N_8452,N_8548);
xnor U9019 (N_9019,N_8533,N_8623);
or U9020 (N_9020,N_8745,N_8406);
xor U9021 (N_9021,N_8624,N_8902);
xor U9022 (N_9022,N_8869,N_8867);
nand U9023 (N_9023,N_8685,N_8737);
or U9024 (N_9024,N_8319,N_8645);
xnor U9025 (N_9025,N_8827,N_8299);
or U9026 (N_9026,N_8423,N_8894);
nor U9027 (N_9027,N_8261,N_8353);
nor U9028 (N_9028,N_8412,N_8838);
nor U9029 (N_9029,N_8783,N_8736);
xor U9030 (N_9030,N_8682,N_8892);
and U9031 (N_9031,N_8443,N_8312);
or U9032 (N_9032,N_8268,N_8959);
and U9033 (N_9033,N_8669,N_8436);
nand U9034 (N_9034,N_8858,N_8393);
nand U9035 (N_9035,N_8333,N_8971);
or U9036 (N_9036,N_8392,N_8912);
xnor U9037 (N_9037,N_8519,N_8621);
nand U9038 (N_9038,N_8395,N_8524);
xor U9039 (N_9039,N_8535,N_8865);
nand U9040 (N_9040,N_8944,N_8507);
nand U9041 (N_9041,N_8954,N_8918);
nor U9042 (N_9042,N_8481,N_8697);
and U9043 (N_9043,N_8778,N_8391);
nor U9044 (N_9044,N_8269,N_8916);
and U9045 (N_9045,N_8492,N_8633);
nand U9046 (N_9046,N_8769,N_8933);
or U9047 (N_9047,N_8584,N_8594);
nor U9048 (N_9048,N_8935,N_8260);
xor U9049 (N_9049,N_8486,N_8801);
nor U9050 (N_9050,N_8262,N_8377);
or U9051 (N_9051,N_8732,N_8637);
or U9052 (N_9052,N_8466,N_8511);
or U9053 (N_9053,N_8907,N_8561);
and U9054 (N_9054,N_8837,N_8836);
or U9055 (N_9055,N_8327,N_8354);
xor U9056 (N_9056,N_8559,N_8698);
or U9057 (N_9057,N_8870,N_8693);
or U9058 (N_9058,N_8920,N_8344);
and U9059 (N_9059,N_8814,N_8609);
nor U9060 (N_9060,N_8845,N_8390);
nor U9061 (N_9061,N_8277,N_8539);
xnor U9062 (N_9062,N_8427,N_8718);
nand U9063 (N_9063,N_8648,N_8315);
and U9064 (N_9064,N_8983,N_8704);
and U9065 (N_9065,N_8947,N_8540);
or U9066 (N_9066,N_8529,N_8781);
xor U9067 (N_9067,N_8639,N_8430);
nand U9068 (N_9068,N_8348,N_8893);
xnor U9069 (N_9069,N_8385,N_8469);
xnor U9070 (N_9070,N_8628,N_8338);
or U9071 (N_9071,N_8713,N_8405);
nand U9072 (N_9072,N_8644,N_8283);
xor U9073 (N_9073,N_8989,N_8946);
and U9074 (N_9074,N_8985,N_8566);
nor U9075 (N_9075,N_8311,N_8929);
or U9076 (N_9076,N_8780,N_8330);
or U9077 (N_9077,N_8349,N_8803);
and U9078 (N_9078,N_8374,N_8942);
nand U9079 (N_9079,N_8501,N_8706);
nor U9080 (N_9080,N_8909,N_8728);
and U9081 (N_9081,N_8683,N_8415);
or U9082 (N_9082,N_8674,N_8589);
nand U9083 (N_9083,N_8958,N_8977);
nand U9084 (N_9084,N_8911,N_8785);
nor U9085 (N_9085,N_8699,N_8284);
and U9086 (N_9086,N_8489,N_8352);
nor U9087 (N_9087,N_8343,N_8538);
nor U9088 (N_9088,N_8308,N_8571);
xnor U9089 (N_9089,N_8477,N_8642);
or U9090 (N_9090,N_8372,N_8378);
nand U9091 (N_9091,N_8886,N_8313);
nand U9092 (N_9092,N_8653,N_8282);
or U9093 (N_9093,N_8362,N_8402);
nor U9094 (N_9094,N_8513,N_8480);
and U9095 (N_9095,N_8413,N_8582);
nor U9096 (N_9096,N_8906,N_8611);
nor U9097 (N_9097,N_8474,N_8657);
and U9098 (N_9098,N_8922,N_8991);
or U9099 (N_9099,N_8305,N_8808);
and U9100 (N_9100,N_8578,N_8748);
and U9101 (N_9101,N_8579,N_8440);
and U9102 (N_9102,N_8339,N_8273);
nand U9103 (N_9103,N_8766,N_8288);
and U9104 (N_9104,N_8455,N_8588);
xnor U9105 (N_9105,N_8450,N_8301);
and U9106 (N_9106,N_8270,N_8847);
nand U9107 (N_9107,N_8461,N_8964);
nand U9108 (N_9108,N_8924,N_8323);
or U9109 (N_9109,N_8563,N_8754);
and U9110 (N_9110,N_8613,N_8722);
xor U9111 (N_9111,N_8379,N_8855);
xor U9112 (N_9112,N_8555,N_8309);
nor U9113 (N_9113,N_8723,N_8788);
nand U9114 (N_9114,N_8360,N_8537);
nor U9115 (N_9115,N_8750,N_8771);
or U9116 (N_9116,N_8546,N_8716);
nor U9117 (N_9117,N_8428,N_8521);
or U9118 (N_9118,N_8665,N_8735);
and U9119 (N_9119,N_8341,N_8979);
nor U9120 (N_9120,N_8557,N_8744);
and U9121 (N_9121,N_8951,N_8266);
xnor U9122 (N_9122,N_8671,N_8363);
nor U9123 (N_9123,N_8523,N_8941);
xor U9124 (N_9124,N_8351,N_8749);
or U9125 (N_9125,N_8967,N_8792);
or U9126 (N_9126,N_8553,N_8705);
nand U9127 (N_9127,N_8518,N_8531);
xnor U9128 (N_9128,N_8791,N_8673);
xor U9129 (N_9129,N_8357,N_8835);
and U9130 (N_9130,N_8765,N_8863);
or U9131 (N_9131,N_8514,N_8310);
and U9132 (N_9132,N_8543,N_8291);
xor U9133 (N_9133,N_8799,N_8418);
nor U9134 (N_9134,N_8250,N_8652);
or U9135 (N_9135,N_8687,N_8451);
or U9136 (N_9136,N_8380,N_8646);
nand U9137 (N_9137,N_8640,N_8331);
and U9138 (N_9138,N_8509,N_8986);
nand U9139 (N_9139,N_8517,N_8585);
and U9140 (N_9140,N_8369,N_8478);
or U9141 (N_9141,N_8251,N_8690);
and U9142 (N_9142,N_8446,N_8729);
nor U9143 (N_9143,N_8700,N_8844);
nand U9144 (N_9144,N_8743,N_8595);
or U9145 (N_9145,N_8404,N_8714);
xor U9146 (N_9146,N_8528,N_8494);
xor U9147 (N_9147,N_8678,N_8365);
and U9148 (N_9148,N_8897,N_8410);
and U9149 (N_9149,N_8321,N_8618);
nor U9150 (N_9150,N_8696,N_8914);
or U9151 (N_9151,N_8820,N_8281);
or U9152 (N_9152,N_8583,N_8275);
and U9153 (N_9153,N_8414,N_8527);
and U9154 (N_9154,N_8794,N_8864);
nand U9155 (N_9155,N_8576,N_8952);
or U9156 (N_9156,N_8751,N_8565);
or U9157 (N_9157,N_8987,N_8634);
or U9158 (N_9158,N_8472,N_8600);
nor U9159 (N_9159,N_8641,N_8426);
nor U9160 (N_9160,N_8775,N_8479);
xnor U9161 (N_9161,N_8998,N_8580);
or U9162 (N_9162,N_8992,N_8325);
nor U9163 (N_9163,N_8361,N_8849);
and U9164 (N_9164,N_8741,N_8953);
or U9165 (N_9165,N_8833,N_8364);
nor U9166 (N_9166,N_8787,N_8295);
xor U9167 (N_9167,N_8937,N_8843);
xor U9168 (N_9168,N_8710,N_8570);
or U9169 (N_9169,N_8448,N_8949);
nand U9170 (N_9170,N_8738,N_8759);
nor U9171 (N_9171,N_8821,N_8485);
xnor U9172 (N_9172,N_8254,N_8468);
or U9173 (N_9173,N_8724,N_8431);
nand U9174 (N_9174,N_8829,N_8770);
and U9175 (N_9175,N_8558,N_8996);
nor U9176 (N_9176,N_8488,N_8635);
nor U9177 (N_9177,N_8381,N_8850);
and U9178 (N_9178,N_8358,N_8972);
nand U9179 (N_9179,N_8449,N_8731);
or U9180 (N_9180,N_8453,N_8715);
or U9181 (N_9181,N_8638,N_8661);
or U9182 (N_9182,N_8675,N_8278);
xor U9183 (N_9183,N_8419,N_8802);
and U9184 (N_9184,N_8471,N_8923);
xnor U9185 (N_9185,N_8672,N_8854);
or U9186 (N_9186,N_8755,N_8296);
and U9187 (N_9187,N_8890,N_8701);
and U9188 (N_9188,N_8320,N_8928);
and U9189 (N_9189,N_8265,N_8515);
xor U9190 (N_9190,N_8614,N_8491);
nand U9191 (N_9191,N_8435,N_8608);
and U9192 (N_9192,N_8655,N_8931);
xnor U9193 (N_9193,N_8574,N_8293);
nor U9194 (N_9194,N_8596,N_8908);
nor U9195 (N_9195,N_8556,N_8948);
nor U9196 (N_9196,N_8981,N_8968);
nor U9197 (N_9197,N_8355,N_8602);
nand U9198 (N_9198,N_8544,N_8569);
and U9199 (N_9199,N_8915,N_8940);
nor U9200 (N_9200,N_8978,N_8962);
and U9201 (N_9201,N_8264,N_8830);
xor U9202 (N_9202,N_8943,N_8495);
and U9203 (N_9203,N_8593,N_8782);
nor U9204 (N_9204,N_8454,N_8840);
nor U9205 (N_9205,N_8885,N_8403);
and U9206 (N_9206,N_8617,N_8417);
xor U9207 (N_9207,N_8689,N_8562);
or U9208 (N_9208,N_8542,N_8373);
and U9209 (N_9209,N_8314,N_8810);
xor U9210 (N_9210,N_8447,N_8707);
and U9211 (N_9211,N_8550,N_8811);
xnor U9212 (N_9212,N_8610,N_8532);
or U9213 (N_9213,N_8879,N_8703);
and U9214 (N_9214,N_8259,N_8368);
xor U9215 (N_9215,N_8966,N_8702);
nor U9216 (N_9216,N_8605,N_8512);
or U9217 (N_9217,N_8625,N_8825);
and U9218 (N_9218,N_8287,N_8334);
nor U9219 (N_9219,N_8302,N_8476);
or U9220 (N_9220,N_8670,N_8656);
or U9221 (N_9221,N_8592,N_8598);
nand U9222 (N_9222,N_8899,N_8408);
and U9223 (N_9223,N_8632,N_8950);
nor U9224 (N_9224,N_8647,N_8257);
nand U9225 (N_9225,N_8806,N_8725);
or U9226 (N_9226,N_8888,N_8988);
or U9227 (N_9227,N_8607,N_8622);
nor U9228 (N_9228,N_8797,N_8397);
or U9229 (N_9229,N_8322,N_8874);
and U9230 (N_9230,N_8603,N_8547);
or U9231 (N_9231,N_8868,N_8575);
nor U9232 (N_9232,N_8332,N_8597);
or U9233 (N_9233,N_8434,N_8601);
xnor U9234 (N_9234,N_8317,N_8955);
nand U9235 (N_9235,N_8846,N_8460);
and U9236 (N_9236,N_8636,N_8359);
nand U9237 (N_9237,N_8875,N_8438);
nor U9238 (N_9238,N_8615,N_8997);
or U9239 (N_9239,N_8534,N_8761);
nor U9240 (N_9240,N_8721,N_8437);
and U9241 (N_9241,N_8668,N_8346);
or U9242 (N_9242,N_8587,N_8429);
or U9243 (N_9243,N_8629,N_8303);
nor U9244 (N_9244,N_8336,N_8384);
or U9245 (N_9245,N_8848,N_8851);
nor U9246 (N_9246,N_8649,N_8289);
nor U9247 (N_9247,N_8932,N_8773);
nor U9248 (N_9248,N_8292,N_8409);
xor U9249 (N_9249,N_8999,N_8457);
and U9250 (N_9250,N_8913,N_8730);
nand U9251 (N_9251,N_8462,N_8300);
nor U9252 (N_9252,N_8679,N_8927);
xnor U9253 (N_9253,N_8880,N_8753);
nor U9254 (N_9254,N_8980,N_8826);
nor U9255 (N_9255,N_8993,N_8733);
nand U9256 (N_9256,N_8482,N_8823);
and U9257 (N_9257,N_8473,N_8508);
xor U9258 (N_9258,N_8526,N_8659);
nand U9259 (N_9259,N_8963,N_8643);
nor U9260 (N_9260,N_8856,N_8859);
nor U9261 (N_9261,N_8459,N_8387);
nand U9262 (N_9262,N_8926,N_8347);
or U9263 (N_9263,N_8763,N_8626);
or U9264 (N_9264,N_8442,N_8272);
and U9265 (N_9265,N_8465,N_8467);
and U9266 (N_9266,N_8554,N_8490);
or U9267 (N_9267,N_8936,N_8662);
or U9268 (N_9268,N_8483,N_8774);
nand U9269 (N_9269,N_8411,N_8620);
nand U9270 (N_9270,N_8340,N_8982);
nor U9271 (N_9271,N_8790,N_8764);
nand U9272 (N_9272,N_8925,N_8376);
or U9273 (N_9273,N_8901,N_8938);
nand U9274 (N_9274,N_8889,N_8917);
xor U9275 (N_9275,N_8274,N_8590);
and U9276 (N_9276,N_8388,N_8734);
xnor U9277 (N_9277,N_8258,N_8502);
xor U9278 (N_9278,N_8536,N_8458);
xnor U9279 (N_9279,N_8255,N_8383);
and U9280 (N_9280,N_8420,N_8712);
nor U9281 (N_9281,N_8768,N_8757);
xor U9282 (N_9282,N_8541,N_8815);
nand U9283 (N_9283,N_8522,N_8416);
nor U9284 (N_9284,N_8930,N_8793);
xor U9285 (N_9285,N_8298,N_8329);
and U9286 (N_9286,N_8719,N_8324);
and U9287 (N_9287,N_8900,N_8573);
nand U9288 (N_9288,N_8800,N_8433);
and U9289 (N_9289,N_8505,N_8817);
or U9290 (N_9290,N_8525,N_8726);
or U9291 (N_9291,N_8267,N_8767);
and U9292 (N_9292,N_8279,N_8905);
or U9293 (N_9293,N_8904,N_8976);
nor U9294 (N_9294,N_8939,N_8887);
and U9295 (N_9295,N_8970,N_8432);
and U9296 (N_9296,N_8684,N_8752);
and U9297 (N_9297,N_8328,N_8842);
or U9298 (N_9298,N_8286,N_8294);
xor U9299 (N_9299,N_8965,N_8396);
xnor U9300 (N_9300,N_8456,N_8382);
and U9301 (N_9301,N_8681,N_8552);
xor U9302 (N_9302,N_8921,N_8470);
xnor U9303 (N_9303,N_8627,N_8853);
and U9304 (N_9304,N_8884,N_8709);
or U9305 (N_9305,N_8496,N_8995);
xnor U9306 (N_9306,N_8816,N_8425);
nand U9307 (N_9307,N_8660,N_8498);
nand U9308 (N_9308,N_8882,N_8439);
or U9309 (N_9309,N_8307,N_8484);
nand U9310 (N_9310,N_8503,N_8394);
and U9311 (N_9311,N_8606,N_8919);
and U9312 (N_9312,N_8756,N_8831);
and U9313 (N_9313,N_8499,N_8974);
xor U9314 (N_9314,N_8798,N_8676);
or U9315 (N_9315,N_8421,N_8688);
or U9316 (N_9316,N_8878,N_8493);
and U9317 (N_9317,N_8549,N_8839);
nor U9318 (N_9318,N_8871,N_8401);
xnor U9319 (N_9319,N_8692,N_8796);
nand U9320 (N_9320,N_8784,N_8777);
nand U9321 (N_9321,N_8818,N_8463);
nand U9322 (N_9322,N_8475,N_8786);
xor U9323 (N_9323,N_8857,N_8304);
or U9324 (N_9324,N_8739,N_8819);
nor U9325 (N_9325,N_8834,N_8895);
nor U9326 (N_9326,N_8370,N_8910);
nor U9327 (N_9327,N_8422,N_8861);
nand U9328 (N_9328,N_8444,N_8650);
nand U9329 (N_9329,N_8487,N_8445);
nand U9330 (N_9330,N_8760,N_8813);
xnor U9331 (N_9331,N_8280,N_8506);
and U9332 (N_9332,N_8654,N_8708);
xnor U9333 (N_9333,N_8658,N_8375);
and U9334 (N_9334,N_8398,N_8290);
nand U9335 (N_9335,N_8318,N_8367);
nor U9336 (N_9336,N_8994,N_8572);
or U9337 (N_9337,N_8567,N_8852);
xnor U9338 (N_9338,N_8500,N_8812);
nand U9339 (N_9339,N_8663,N_8297);
xnor U9340 (N_9340,N_8577,N_8828);
or U9341 (N_9341,N_8711,N_8717);
or U9342 (N_9342,N_8742,N_8695);
and U9343 (N_9343,N_8776,N_8727);
xor U9344 (N_9344,N_8896,N_8961);
nand U9345 (N_9345,N_8832,N_8604);
nor U9346 (N_9346,N_8779,N_8883);
nand U9347 (N_9347,N_8677,N_8680);
nor U9348 (N_9348,N_8337,N_8795);
and U9349 (N_9349,N_8651,N_8520);
nor U9350 (N_9350,N_8424,N_8350);
xnor U9351 (N_9351,N_8957,N_8263);
and U9352 (N_9352,N_8464,N_8371);
nor U9353 (N_9353,N_8510,N_8586);
and U9354 (N_9354,N_8809,N_8758);
nand U9355 (N_9355,N_8591,N_8824);
nand U9356 (N_9356,N_8860,N_8616);
xor U9357 (N_9357,N_8973,N_8545);
xor U9358 (N_9358,N_8876,N_8720);
nand U9359 (N_9359,N_8990,N_8631);
nor U9360 (N_9360,N_8504,N_8399);
nor U9361 (N_9361,N_8807,N_8694);
xor U9362 (N_9362,N_8564,N_8356);
nand U9363 (N_9363,N_8934,N_8772);
xnor U9364 (N_9364,N_8667,N_8804);
nand U9365 (N_9365,N_8335,N_8285);
or U9366 (N_9366,N_8276,N_8866);
nand U9367 (N_9367,N_8686,N_8881);
or U9368 (N_9368,N_8407,N_8253);
or U9369 (N_9369,N_8664,N_8271);
xnor U9370 (N_9370,N_8789,N_8316);
nor U9371 (N_9371,N_8400,N_8891);
and U9372 (N_9372,N_8599,N_8691);
xor U9373 (N_9373,N_8516,N_8747);
or U9374 (N_9374,N_8822,N_8872);
nand U9375 (N_9375,N_8906,N_8968);
and U9376 (N_9376,N_8811,N_8402);
nor U9377 (N_9377,N_8299,N_8641);
xnor U9378 (N_9378,N_8827,N_8346);
or U9379 (N_9379,N_8406,N_8658);
xnor U9380 (N_9380,N_8711,N_8922);
and U9381 (N_9381,N_8272,N_8947);
nand U9382 (N_9382,N_8845,N_8511);
or U9383 (N_9383,N_8481,N_8918);
and U9384 (N_9384,N_8816,N_8526);
nand U9385 (N_9385,N_8312,N_8737);
nand U9386 (N_9386,N_8852,N_8587);
or U9387 (N_9387,N_8819,N_8623);
nor U9388 (N_9388,N_8551,N_8930);
xor U9389 (N_9389,N_8897,N_8704);
and U9390 (N_9390,N_8492,N_8521);
nor U9391 (N_9391,N_8678,N_8807);
xnor U9392 (N_9392,N_8989,N_8360);
nor U9393 (N_9393,N_8341,N_8812);
nand U9394 (N_9394,N_8546,N_8736);
nor U9395 (N_9395,N_8565,N_8870);
and U9396 (N_9396,N_8771,N_8931);
nor U9397 (N_9397,N_8813,N_8927);
or U9398 (N_9398,N_8655,N_8824);
nor U9399 (N_9399,N_8515,N_8559);
or U9400 (N_9400,N_8823,N_8270);
xnor U9401 (N_9401,N_8305,N_8788);
and U9402 (N_9402,N_8810,N_8267);
or U9403 (N_9403,N_8387,N_8371);
and U9404 (N_9404,N_8268,N_8427);
nor U9405 (N_9405,N_8515,N_8414);
or U9406 (N_9406,N_8784,N_8619);
and U9407 (N_9407,N_8977,N_8401);
or U9408 (N_9408,N_8786,N_8677);
and U9409 (N_9409,N_8323,N_8546);
and U9410 (N_9410,N_8583,N_8820);
and U9411 (N_9411,N_8648,N_8853);
and U9412 (N_9412,N_8821,N_8483);
nand U9413 (N_9413,N_8571,N_8548);
and U9414 (N_9414,N_8557,N_8775);
and U9415 (N_9415,N_8560,N_8584);
nand U9416 (N_9416,N_8941,N_8945);
or U9417 (N_9417,N_8760,N_8748);
nor U9418 (N_9418,N_8804,N_8857);
and U9419 (N_9419,N_8251,N_8399);
and U9420 (N_9420,N_8585,N_8740);
or U9421 (N_9421,N_8891,N_8516);
nor U9422 (N_9422,N_8467,N_8857);
nor U9423 (N_9423,N_8289,N_8412);
nand U9424 (N_9424,N_8311,N_8924);
nand U9425 (N_9425,N_8447,N_8994);
xnor U9426 (N_9426,N_8595,N_8683);
nand U9427 (N_9427,N_8831,N_8407);
nor U9428 (N_9428,N_8677,N_8933);
xnor U9429 (N_9429,N_8871,N_8983);
nand U9430 (N_9430,N_8456,N_8794);
or U9431 (N_9431,N_8894,N_8271);
nor U9432 (N_9432,N_8914,N_8831);
nand U9433 (N_9433,N_8613,N_8378);
and U9434 (N_9434,N_8409,N_8565);
xor U9435 (N_9435,N_8519,N_8835);
or U9436 (N_9436,N_8422,N_8935);
or U9437 (N_9437,N_8281,N_8886);
nor U9438 (N_9438,N_8314,N_8610);
nand U9439 (N_9439,N_8671,N_8397);
nor U9440 (N_9440,N_8730,N_8884);
or U9441 (N_9441,N_8349,N_8586);
nand U9442 (N_9442,N_8822,N_8566);
or U9443 (N_9443,N_8854,N_8269);
xnor U9444 (N_9444,N_8914,N_8338);
nor U9445 (N_9445,N_8404,N_8736);
or U9446 (N_9446,N_8917,N_8742);
and U9447 (N_9447,N_8738,N_8291);
nand U9448 (N_9448,N_8702,N_8607);
nand U9449 (N_9449,N_8941,N_8271);
nor U9450 (N_9450,N_8848,N_8901);
xnor U9451 (N_9451,N_8799,N_8713);
and U9452 (N_9452,N_8844,N_8453);
nand U9453 (N_9453,N_8709,N_8596);
and U9454 (N_9454,N_8749,N_8810);
or U9455 (N_9455,N_8839,N_8795);
xor U9456 (N_9456,N_8623,N_8371);
or U9457 (N_9457,N_8825,N_8912);
xnor U9458 (N_9458,N_8780,N_8870);
xor U9459 (N_9459,N_8869,N_8979);
and U9460 (N_9460,N_8755,N_8588);
nor U9461 (N_9461,N_8388,N_8873);
or U9462 (N_9462,N_8468,N_8627);
nand U9463 (N_9463,N_8768,N_8772);
nand U9464 (N_9464,N_8566,N_8771);
xor U9465 (N_9465,N_8657,N_8955);
nor U9466 (N_9466,N_8918,N_8504);
or U9467 (N_9467,N_8734,N_8375);
and U9468 (N_9468,N_8760,N_8438);
or U9469 (N_9469,N_8684,N_8389);
and U9470 (N_9470,N_8810,N_8875);
or U9471 (N_9471,N_8746,N_8987);
and U9472 (N_9472,N_8303,N_8581);
and U9473 (N_9473,N_8366,N_8942);
or U9474 (N_9474,N_8830,N_8579);
nand U9475 (N_9475,N_8964,N_8500);
nand U9476 (N_9476,N_8963,N_8376);
and U9477 (N_9477,N_8656,N_8350);
or U9478 (N_9478,N_8301,N_8490);
or U9479 (N_9479,N_8812,N_8740);
nor U9480 (N_9480,N_8477,N_8400);
nor U9481 (N_9481,N_8622,N_8741);
nand U9482 (N_9482,N_8282,N_8587);
nand U9483 (N_9483,N_8932,N_8731);
and U9484 (N_9484,N_8585,N_8602);
nor U9485 (N_9485,N_8649,N_8915);
nor U9486 (N_9486,N_8804,N_8532);
xor U9487 (N_9487,N_8694,N_8559);
or U9488 (N_9488,N_8738,N_8783);
or U9489 (N_9489,N_8524,N_8879);
xnor U9490 (N_9490,N_8828,N_8552);
and U9491 (N_9491,N_8618,N_8492);
nor U9492 (N_9492,N_8556,N_8690);
and U9493 (N_9493,N_8901,N_8312);
nand U9494 (N_9494,N_8530,N_8646);
nor U9495 (N_9495,N_8928,N_8285);
nand U9496 (N_9496,N_8962,N_8558);
nor U9497 (N_9497,N_8342,N_8600);
xnor U9498 (N_9498,N_8409,N_8748);
or U9499 (N_9499,N_8306,N_8532);
nand U9500 (N_9500,N_8760,N_8910);
xnor U9501 (N_9501,N_8345,N_8936);
or U9502 (N_9502,N_8965,N_8305);
or U9503 (N_9503,N_8864,N_8288);
and U9504 (N_9504,N_8896,N_8713);
and U9505 (N_9505,N_8289,N_8525);
nand U9506 (N_9506,N_8635,N_8811);
xnor U9507 (N_9507,N_8373,N_8941);
xor U9508 (N_9508,N_8737,N_8798);
and U9509 (N_9509,N_8812,N_8270);
and U9510 (N_9510,N_8683,N_8744);
and U9511 (N_9511,N_8373,N_8802);
nor U9512 (N_9512,N_8271,N_8583);
nand U9513 (N_9513,N_8269,N_8888);
and U9514 (N_9514,N_8356,N_8443);
or U9515 (N_9515,N_8565,N_8488);
nor U9516 (N_9516,N_8829,N_8693);
nor U9517 (N_9517,N_8739,N_8590);
nand U9518 (N_9518,N_8635,N_8994);
nand U9519 (N_9519,N_8408,N_8694);
nand U9520 (N_9520,N_8901,N_8561);
or U9521 (N_9521,N_8938,N_8568);
and U9522 (N_9522,N_8433,N_8721);
and U9523 (N_9523,N_8395,N_8668);
nor U9524 (N_9524,N_8292,N_8555);
nor U9525 (N_9525,N_8416,N_8422);
nor U9526 (N_9526,N_8680,N_8383);
nor U9527 (N_9527,N_8623,N_8924);
or U9528 (N_9528,N_8619,N_8424);
or U9529 (N_9529,N_8296,N_8556);
nor U9530 (N_9530,N_8775,N_8546);
nand U9531 (N_9531,N_8524,N_8921);
and U9532 (N_9532,N_8378,N_8376);
xnor U9533 (N_9533,N_8505,N_8867);
nand U9534 (N_9534,N_8551,N_8359);
xor U9535 (N_9535,N_8432,N_8303);
or U9536 (N_9536,N_8800,N_8872);
or U9537 (N_9537,N_8866,N_8831);
nand U9538 (N_9538,N_8463,N_8288);
xnor U9539 (N_9539,N_8479,N_8500);
and U9540 (N_9540,N_8672,N_8621);
and U9541 (N_9541,N_8858,N_8371);
nor U9542 (N_9542,N_8614,N_8803);
xor U9543 (N_9543,N_8436,N_8935);
and U9544 (N_9544,N_8561,N_8369);
xor U9545 (N_9545,N_8666,N_8535);
or U9546 (N_9546,N_8418,N_8687);
xor U9547 (N_9547,N_8446,N_8908);
and U9548 (N_9548,N_8410,N_8652);
nor U9549 (N_9549,N_8909,N_8784);
nand U9550 (N_9550,N_8982,N_8973);
xor U9551 (N_9551,N_8484,N_8664);
nand U9552 (N_9552,N_8439,N_8846);
nand U9553 (N_9553,N_8970,N_8466);
nand U9554 (N_9554,N_8474,N_8877);
nor U9555 (N_9555,N_8599,N_8430);
nor U9556 (N_9556,N_8365,N_8796);
and U9557 (N_9557,N_8650,N_8409);
nor U9558 (N_9558,N_8910,N_8374);
xnor U9559 (N_9559,N_8992,N_8925);
nand U9560 (N_9560,N_8752,N_8573);
nand U9561 (N_9561,N_8560,N_8522);
nand U9562 (N_9562,N_8323,N_8958);
nor U9563 (N_9563,N_8817,N_8457);
or U9564 (N_9564,N_8314,N_8957);
nand U9565 (N_9565,N_8811,N_8421);
xor U9566 (N_9566,N_8968,N_8443);
nor U9567 (N_9567,N_8395,N_8821);
nand U9568 (N_9568,N_8680,N_8805);
nand U9569 (N_9569,N_8476,N_8385);
nand U9570 (N_9570,N_8929,N_8520);
nor U9571 (N_9571,N_8945,N_8482);
or U9572 (N_9572,N_8263,N_8694);
or U9573 (N_9573,N_8590,N_8950);
nand U9574 (N_9574,N_8531,N_8991);
nand U9575 (N_9575,N_8834,N_8297);
nand U9576 (N_9576,N_8375,N_8571);
and U9577 (N_9577,N_8285,N_8585);
nor U9578 (N_9578,N_8584,N_8841);
or U9579 (N_9579,N_8737,N_8511);
or U9580 (N_9580,N_8479,N_8697);
xnor U9581 (N_9581,N_8469,N_8969);
and U9582 (N_9582,N_8356,N_8908);
and U9583 (N_9583,N_8975,N_8672);
nand U9584 (N_9584,N_8292,N_8696);
nor U9585 (N_9585,N_8284,N_8612);
or U9586 (N_9586,N_8250,N_8863);
and U9587 (N_9587,N_8935,N_8639);
nand U9588 (N_9588,N_8511,N_8582);
nand U9589 (N_9589,N_8588,N_8884);
nand U9590 (N_9590,N_8844,N_8646);
or U9591 (N_9591,N_8343,N_8746);
nor U9592 (N_9592,N_8812,N_8641);
nand U9593 (N_9593,N_8808,N_8874);
nand U9594 (N_9594,N_8761,N_8871);
and U9595 (N_9595,N_8898,N_8838);
and U9596 (N_9596,N_8737,N_8928);
and U9597 (N_9597,N_8635,N_8523);
xor U9598 (N_9598,N_8852,N_8658);
xor U9599 (N_9599,N_8320,N_8308);
nand U9600 (N_9600,N_8816,N_8722);
and U9601 (N_9601,N_8605,N_8439);
nand U9602 (N_9602,N_8994,N_8768);
nor U9603 (N_9603,N_8424,N_8918);
xnor U9604 (N_9604,N_8760,N_8592);
xnor U9605 (N_9605,N_8661,N_8420);
nor U9606 (N_9606,N_8494,N_8250);
xnor U9607 (N_9607,N_8895,N_8258);
nor U9608 (N_9608,N_8705,N_8844);
nand U9609 (N_9609,N_8564,N_8997);
or U9610 (N_9610,N_8696,N_8307);
or U9611 (N_9611,N_8484,N_8915);
xor U9612 (N_9612,N_8521,N_8647);
nand U9613 (N_9613,N_8823,N_8634);
xnor U9614 (N_9614,N_8614,N_8535);
xnor U9615 (N_9615,N_8707,N_8349);
and U9616 (N_9616,N_8462,N_8360);
nand U9617 (N_9617,N_8767,N_8408);
xor U9618 (N_9618,N_8347,N_8265);
and U9619 (N_9619,N_8293,N_8468);
nand U9620 (N_9620,N_8260,N_8584);
xor U9621 (N_9621,N_8442,N_8930);
xor U9622 (N_9622,N_8674,N_8784);
nand U9623 (N_9623,N_8987,N_8333);
xor U9624 (N_9624,N_8310,N_8761);
nor U9625 (N_9625,N_8834,N_8273);
nand U9626 (N_9626,N_8333,N_8565);
nor U9627 (N_9627,N_8661,N_8410);
or U9628 (N_9628,N_8286,N_8502);
nor U9629 (N_9629,N_8303,N_8341);
and U9630 (N_9630,N_8551,N_8281);
nand U9631 (N_9631,N_8542,N_8291);
nand U9632 (N_9632,N_8781,N_8695);
nor U9633 (N_9633,N_8944,N_8692);
nand U9634 (N_9634,N_8946,N_8957);
nand U9635 (N_9635,N_8648,N_8295);
nor U9636 (N_9636,N_8600,N_8758);
nor U9637 (N_9637,N_8632,N_8271);
and U9638 (N_9638,N_8890,N_8675);
nor U9639 (N_9639,N_8919,N_8699);
nand U9640 (N_9640,N_8953,N_8543);
xor U9641 (N_9641,N_8690,N_8695);
and U9642 (N_9642,N_8303,N_8579);
xor U9643 (N_9643,N_8483,N_8904);
nor U9644 (N_9644,N_8616,N_8515);
and U9645 (N_9645,N_8594,N_8865);
or U9646 (N_9646,N_8964,N_8412);
and U9647 (N_9647,N_8957,N_8780);
nor U9648 (N_9648,N_8686,N_8690);
and U9649 (N_9649,N_8811,N_8800);
nand U9650 (N_9650,N_8660,N_8603);
xor U9651 (N_9651,N_8807,N_8605);
or U9652 (N_9652,N_8868,N_8614);
or U9653 (N_9653,N_8373,N_8370);
and U9654 (N_9654,N_8901,N_8775);
and U9655 (N_9655,N_8507,N_8680);
or U9656 (N_9656,N_8305,N_8393);
or U9657 (N_9657,N_8302,N_8633);
xnor U9658 (N_9658,N_8375,N_8744);
or U9659 (N_9659,N_8826,N_8790);
nand U9660 (N_9660,N_8813,N_8562);
xnor U9661 (N_9661,N_8651,N_8362);
nor U9662 (N_9662,N_8682,N_8603);
and U9663 (N_9663,N_8871,N_8382);
nor U9664 (N_9664,N_8911,N_8505);
or U9665 (N_9665,N_8659,N_8986);
and U9666 (N_9666,N_8552,N_8262);
nor U9667 (N_9667,N_8628,N_8955);
or U9668 (N_9668,N_8609,N_8330);
nor U9669 (N_9669,N_8732,N_8682);
and U9670 (N_9670,N_8936,N_8631);
or U9671 (N_9671,N_8274,N_8475);
and U9672 (N_9672,N_8836,N_8396);
nand U9673 (N_9673,N_8746,N_8425);
and U9674 (N_9674,N_8939,N_8595);
or U9675 (N_9675,N_8852,N_8765);
nand U9676 (N_9676,N_8823,N_8407);
nand U9677 (N_9677,N_8415,N_8595);
nor U9678 (N_9678,N_8562,N_8543);
nand U9679 (N_9679,N_8901,N_8421);
xnor U9680 (N_9680,N_8727,N_8531);
xor U9681 (N_9681,N_8459,N_8785);
xor U9682 (N_9682,N_8896,N_8860);
nand U9683 (N_9683,N_8992,N_8711);
nor U9684 (N_9684,N_8354,N_8321);
xor U9685 (N_9685,N_8943,N_8859);
xor U9686 (N_9686,N_8554,N_8558);
nor U9687 (N_9687,N_8681,N_8501);
nand U9688 (N_9688,N_8334,N_8344);
and U9689 (N_9689,N_8935,N_8435);
or U9690 (N_9690,N_8447,N_8543);
or U9691 (N_9691,N_8662,N_8445);
or U9692 (N_9692,N_8939,N_8360);
nor U9693 (N_9693,N_8561,N_8791);
nand U9694 (N_9694,N_8963,N_8722);
nand U9695 (N_9695,N_8609,N_8726);
and U9696 (N_9696,N_8427,N_8666);
nor U9697 (N_9697,N_8840,N_8458);
or U9698 (N_9698,N_8364,N_8265);
or U9699 (N_9699,N_8460,N_8568);
nand U9700 (N_9700,N_8368,N_8805);
nand U9701 (N_9701,N_8602,N_8939);
or U9702 (N_9702,N_8637,N_8893);
and U9703 (N_9703,N_8739,N_8263);
or U9704 (N_9704,N_8635,N_8718);
nor U9705 (N_9705,N_8290,N_8943);
and U9706 (N_9706,N_8843,N_8498);
nor U9707 (N_9707,N_8461,N_8364);
or U9708 (N_9708,N_8315,N_8594);
and U9709 (N_9709,N_8296,N_8486);
nand U9710 (N_9710,N_8945,N_8409);
and U9711 (N_9711,N_8252,N_8724);
and U9712 (N_9712,N_8902,N_8596);
and U9713 (N_9713,N_8918,N_8921);
and U9714 (N_9714,N_8545,N_8441);
and U9715 (N_9715,N_8408,N_8252);
and U9716 (N_9716,N_8480,N_8859);
xor U9717 (N_9717,N_8740,N_8757);
xnor U9718 (N_9718,N_8603,N_8279);
and U9719 (N_9719,N_8552,N_8862);
nor U9720 (N_9720,N_8882,N_8555);
or U9721 (N_9721,N_8400,N_8671);
and U9722 (N_9722,N_8827,N_8900);
nor U9723 (N_9723,N_8925,N_8413);
and U9724 (N_9724,N_8284,N_8494);
nor U9725 (N_9725,N_8357,N_8706);
and U9726 (N_9726,N_8329,N_8847);
xor U9727 (N_9727,N_8352,N_8885);
nor U9728 (N_9728,N_8793,N_8383);
nor U9729 (N_9729,N_8301,N_8582);
or U9730 (N_9730,N_8467,N_8653);
nor U9731 (N_9731,N_8474,N_8840);
xnor U9732 (N_9732,N_8366,N_8986);
nor U9733 (N_9733,N_8314,N_8524);
xor U9734 (N_9734,N_8415,N_8378);
or U9735 (N_9735,N_8661,N_8590);
and U9736 (N_9736,N_8936,N_8414);
xnor U9737 (N_9737,N_8276,N_8650);
xor U9738 (N_9738,N_8290,N_8306);
and U9739 (N_9739,N_8947,N_8616);
nand U9740 (N_9740,N_8555,N_8580);
or U9741 (N_9741,N_8475,N_8721);
or U9742 (N_9742,N_8706,N_8823);
and U9743 (N_9743,N_8894,N_8624);
nor U9744 (N_9744,N_8947,N_8919);
and U9745 (N_9745,N_8751,N_8442);
and U9746 (N_9746,N_8445,N_8657);
and U9747 (N_9747,N_8824,N_8279);
xor U9748 (N_9748,N_8333,N_8278);
nor U9749 (N_9749,N_8528,N_8383);
xor U9750 (N_9750,N_9038,N_9188);
nor U9751 (N_9751,N_9171,N_9444);
nand U9752 (N_9752,N_9680,N_9478);
xnor U9753 (N_9753,N_9199,N_9546);
nand U9754 (N_9754,N_9559,N_9715);
xor U9755 (N_9755,N_9636,N_9605);
nand U9756 (N_9756,N_9541,N_9134);
and U9757 (N_9757,N_9613,N_9539);
or U9758 (N_9758,N_9317,N_9273);
or U9759 (N_9759,N_9013,N_9452);
xor U9760 (N_9760,N_9101,N_9544);
or U9761 (N_9761,N_9565,N_9018);
or U9762 (N_9762,N_9529,N_9278);
or U9763 (N_9763,N_9649,N_9638);
xnor U9764 (N_9764,N_9545,N_9575);
or U9765 (N_9765,N_9563,N_9702);
nor U9766 (N_9766,N_9265,N_9472);
or U9767 (N_9767,N_9170,N_9527);
xnor U9768 (N_9768,N_9663,N_9289);
xor U9769 (N_9769,N_9586,N_9524);
xor U9770 (N_9770,N_9651,N_9360);
xor U9771 (N_9771,N_9451,N_9588);
and U9772 (N_9772,N_9479,N_9437);
xnor U9773 (N_9773,N_9198,N_9402);
or U9774 (N_9774,N_9032,N_9507);
or U9775 (N_9775,N_9123,N_9017);
nor U9776 (N_9776,N_9313,N_9733);
and U9777 (N_9777,N_9468,N_9597);
xnor U9778 (N_9778,N_9469,N_9495);
xnor U9779 (N_9779,N_9279,N_9266);
or U9780 (N_9780,N_9028,N_9403);
nand U9781 (N_9781,N_9066,N_9552);
and U9782 (N_9782,N_9150,N_9082);
nand U9783 (N_9783,N_9035,N_9489);
xor U9784 (N_9784,N_9136,N_9111);
nand U9785 (N_9785,N_9294,N_9029);
nand U9786 (N_9786,N_9375,N_9416);
or U9787 (N_9787,N_9555,N_9604);
nor U9788 (N_9788,N_9008,N_9502);
and U9789 (N_9789,N_9582,N_9072);
nor U9790 (N_9790,N_9690,N_9735);
nand U9791 (N_9791,N_9387,N_9205);
nor U9792 (N_9792,N_9526,N_9671);
or U9793 (N_9793,N_9430,N_9664);
xnor U9794 (N_9794,N_9543,N_9599);
nor U9795 (N_9795,N_9094,N_9460);
nor U9796 (N_9796,N_9340,N_9408);
and U9797 (N_9797,N_9076,N_9291);
xor U9798 (N_9798,N_9330,N_9019);
nor U9799 (N_9799,N_9210,N_9711);
and U9800 (N_9800,N_9244,N_9394);
or U9801 (N_9801,N_9481,N_9229);
nand U9802 (N_9802,N_9177,N_9295);
nor U9803 (N_9803,N_9354,N_9088);
xnor U9804 (N_9804,N_9738,N_9127);
xnor U9805 (N_9805,N_9499,N_9104);
xor U9806 (N_9806,N_9496,N_9165);
and U9807 (N_9807,N_9730,N_9531);
or U9808 (N_9808,N_9654,N_9637);
nand U9809 (N_9809,N_9522,N_9155);
or U9810 (N_9810,N_9675,N_9246);
and U9811 (N_9811,N_9158,N_9197);
or U9812 (N_9812,N_9620,N_9748);
nand U9813 (N_9813,N_9454,N_9612);
nor U9814 (N_9814,N_9697,N_9348);
xnor U9815 (N_9815,N_9193,N_9359);
nor U9816 (N_9816,N_9269,N_9583);
and U9817 (N_9817,N_9053,N_9463);
nor U9818 (N_9818,N_9204,N_9364);
nand U9819 (N_9819,N_9371,N_9096);
xnor U9820 (N_9820,N_9144,N_9139);
or U9821 (N_9821,N_9536,N_9594);
nand U9822 (N_9822,N_9011,N_9379);
or U9823 (N_9823,N_9323,N_9712);
and U9824 (N_9824,N_9467,N_9607);
and U9825 (N_9825,N_9519,N_9533);
and U9826 (N_9826,N_9576,N_9180);
xnor U9827 (N_9827,N_9643,N_9322);
nor U9828 (N_9828,N_9215,N_9069);
xnor U9829 (N_9829,N_9551,N_9207);
xnor U9830 (N_9830,N_9698,N_9523);
nor U9831 (N_9831,N_9042,N_9513);
or U9832 (N_9832,N_9587,N_9062);
xnor U9833 (N_9833,N_9296,N_9464);
nand U9834 (N_9834,N_9719,N_9457);
nor U9835 (N_9835,N_9435,N_9001);
nand U9836 (N_9836,N_9486,N_9137);
xor U9837 (N_9837,N_9129,N_9578);
and U9838 (N_9838,N_9271,N_9064);
xor U9839 (N_9839,N_9141,N_9329);
nand U9840 (N_9840,N_9259,N_9181);
nand U9841 (N_9841,N_9439,N_9319);
nand U9842 (N_9842,N_9203,N_9135);
and U9843 (N_9843,N_9316,N_9281);
nand U9844 (N_9844,N_9670,N_9126);
and U9845 (N_9845,N_9216,N_9621);
and U9846 (N_9846,N_9355,N_9174);
nand U9847 (N_9847,N_9110,N_9561);
or U9848 (N_9848,N_9668,N_9485);
or U9849 (N_9849,N_9630,N_9234);
nor U9850 (N_9850,N_9247,N_9374);
xnor U9851 (N_9851,N_9743,N_9061);
nand U9852 (N_9852,N_9221,N_9242);
and U9853 (N_9853,N_9645,N_9039);
or U9854 (N_9854,N_9219,N_9238);
nand U9855 (N_9855,N_9441,N_9253);
xor U9856 (N_9856,N_9570,N_9741);
xnor U9857 (N_9857,N_9386,N_9257);
xor U9858 (N_9858,N_9314,N_9632);
nand U9859 (N_9859,N_9365,N_9609);
and U9860 (N_9860,N_9338,N_9746);
or U9861 (N_9861,N_9227,N_9012);
nor U9862 (N_9862,N_9335,N_9046);
or U9863 (N_9863,N_9413,N_9184);
xor U9864 (N_9864,N_9538,N_9625);
and U9865 (N_9865,N_9107,N_9532);
and U9866 (N_9866,N_9392,N_9410);
nor U9867 (N_9867,N_9717,N_9200);
nand U9868 (N_9868,N_9256,N_9015);
xnor U9869 (N_9869,N_9376,N_9431);
and U9870 (N_9870,N_9488,N_9473);
and U9871 (N_9871,N_9677,N_9385);
nand U9872 (N_9872,N_9665,N_9267);
and U9873 (N_9873,N_9579,N_9742);
and U9874 (N_9874,N_9681,N_9143);
or U9875 (N_9875,N_9725,N_9090);
nand U9876 (N_9876,N_9631,N_9689);
nor U9877 (N_9877,N_9706,N_9600);
and U9878 (N_9878,N_9191,N_9307);
nand U9879 (N_9879,N_9049,N_9142);
xnor U9880 (N_9880,N_9087,N_9352);
nand U9881 (N_9881,N_9065,N_9009);
nor U9882 (N_9882,N_9233,N_9713);
and U9883 (N_9883,N_9145,N_9276);
nand U9884 (N_9884,N_9153,N_9208);
or U9885 (N_9885,N_9151,N_9023);
or U9886 (N_9886,N_9390,N_9258);
and U9887 (N_9887,N_9404,N_9747);
nand U9888 (N_9888,N_9428,N_9367);
or U9889 (N_9889,N_9108,N_9280);
and U9890 (N_9890,N_9550,N_9696);
nor U9891 (N_9891,N_9644,N_9080);
or U9892 (N_9892,N_9617,N_9071);
nor U9893 (N_9893,N_9159,N_9293);
and U9894 (N_9894,N_9138,N_9744);
or U9895 (N_9895,N_9156,N_9119);
and U9896 (N_9896,N_9262,N_9068);
xor U9897 (N_9897,N_9571,N_9333);
or U9898 (N_9898,N_9530,N_9459);
nand U9899 (N_9899,N_9749,N_9427);
and U9900 (N_9900,N_9443,N_9679);
nor U9901 (N_9901,N_9089,N_9225);
xnor U9902 (N_9902,N_9109,N_9121);
xor U9903 (N_9903,N_9056,N_9695);
xor U9904 (N_9904,N_9099,N_9103);
nand U9905 (N_9905,N_9226,N_9206);
xnor U9906 (N_9906,N_9498,N_9036);
nor U9907 (N_9907,N_9569,N_9732);
nand U9908 (N_9908,N_9412,N_9251);
and U9909 (N_9909,N_9243,N_9168);
nand U9910 (N_9910,N_9268,N_9629);
xor U9911 (N_9911,N_9492,N_9615);
nand U9912 (N_9912,N_9384,N_9067);
xor U9913 (N_9913,N_9118,N_9154);
or U9914 (N_9914,N_9389,N_9140);
xnor U9915 (N_9915,N_9051,N_9209);
nand U9916 (N_9916,N_9006,N_9231);
or U9917 (N_9917,N_9000,N_9125);
or U9918 (N_9918,N_9590,N_9426);
xnor U9919 (N_9919,N_9573,N_9098);
xnor U9920 (N_9920,N_9623,N_9641);
nand U9921 (N_9921,N_9595,N_9298);
nor U9922 (N_9922,N_9122,N_9382);
and U9923 (N_9923,N_9239,N_9282);
nor U9924 (N_9924,N_9420,N_9554);
and U9925 (N_9925,N_9511,N_9714);
nand U9926 (N_9926,N_9411,N_9102);
nor U9927 (N_9927,N_9491,N_9556);
nor U9928 (N_9928,N_9718,N_9686);
or U9929 (N_9929,N_9650,N_9339);
nor U9930 (N_9930,N_9020,N_9601);
nand U9931 (N_9931,N_9182,N_9611);
nor U9932 (N_9932,N_9037,N_9584);
and U9933 (N_9933,N_9152,N_9602);
nand U9934 (N_9934,N_9453,N_9351);
nand U9935 (N_9935,N_9106,N_9506);
or U9936 (N_9936,N_9297,N_9358);
and U9937 (N_9937,N_9494,N_9054);
xnor U9938 (N_9938,N_9189,N_9508);
or U9939 (N_9939,N_9349,N_9378);
xnor U9940 (N_9940,N_9445,N_9078);
nor U9941 (N_9941,N_9063,N_9327);
and U9942 (N_9942,N_9025,N_9073);
nor U9943 (N_9943,N_9432,N_9624);
xnor U9944 (N_9944,N_9212,N_9377);
nand U9945 (N_9945,N_9501,N_9470);
and U9946 (N_9946,N_9250,N_9477);
or U9947 (N_9947,N_9283,N_9060);
and U9948 (N_9948,N_9547,N_9716);
nand U9949 (N_9949,N_9031,N_9315);
xnor U9950 (N_9950,N_9085,N_9558);
and U9951 (N_9951,N_9639,N_9326);
xnor U9952 (N_9952,N_9424,N_9731);
or U9953 (N_9953,N_9564,N_9606);
and U9954 (N_9954,N_9074,N_9095);
or U9955 (N_9955,N_9081,N_9528);
nor U9956 (N_9956,N_9535,N_9667);
xor U9957 (N_9957,N_9700,N_9537);
nand U9958 (N_9958,N_9252,N_9172);
nor U9959 (N_9959,N_9516,N_9369);
or U9960 (N_9960,N_9456,N_9007);
xor U9961 (N_9961,N_9448,N_9399);
or U9962 (N_9962,N_9237,N_9033);
and U9963 (N_9963,N_9398,N_9673);
nor U9964 (N_9964,N_9346,N_9483);
and U9965 (N_9965,N_9674,N_9490);
and U9966 (N_9966,N_9397,N_9048);
or U9967 (N_9967,N_9091,N_9447);
and U9968 (N_9968,N_9589,N_9691);
xor U9969 (N_9969,N_9070,N_9699);
nand U9970 (N_9970,N_9693,N_9720);
xnor U9971 (N_9971,N_9423,N_9052);
nand U9972 (N_9972,N_9653,N_9634);
or U9973 (N_9973,N_9647,N_9306);
nor U9974 (N_9974,N_9465,N_9192);
nor U9975 (N_9975,N_9505,N_9041);
xor U9976 (N_9976,N_9503,N_9572);
and U9977 (N_9977,N_9190,N_9474);
or U9978 (N_9978,N_9026,N_9476);
nand U9979 (N_9979,N_9059,N_9414);
xnor U9980 (N_9980,N_9662,N_9254);
nor U9981 (N_9981,N_9740,N_9175);
and U9982 (N_9982,N_9311,N_9131);
nand U9983 (N_9983,N_9727,N_9300);
or U9984 (N_9984,N_9368,N_9415);
or U9985 (N_9985,N_9179,N_9147);
and U9986 (N_9986,N_9284,N_9418);
nor U9987 (N_9987,N_9591,N_9117);
nand U9988 (N_9988,N_9652,N_9353);
xnor U9989 (N_9989,N_9320,N_9497);
xor U9990 (N_9990,N_9553,N_9057);
and U9991 (N_9991,N_9462,N_9304);
xnor U9992 (N_9992,N_9610,N_9666);
or U9993 (N_9993,N_9173,N_9396);
xor U9994 (N_9994,N_9093,N_9211);
xnor U9995 (N_9995,N_9024,N_9482);
and U9996 (N_9996,N_9685,N_9201);
nor U9997 (N_9997,N_9292,N_9092);
and U9998 (N_9998,N_9241,N_9512);
or U9999 (N_9999,N_9707,N_9705);
and U10000 (N_10000,N_9356,N_9183);
nor U10001 (N_10001,N_9022,N_9678);
nor U10002 (N_10002,N_9724,N_9703);
nor U10003 (N_10003,N_9433,N_9466);
nand U10004 (N_10004,N_9186,N_9596);
xnor U10005 (N_10005,N_9161,N_9487);
and U10006 (N_10006,N_9164,N_9240);
nand U10007 (N_10007,N_9342,N_9366);
xor U10008 (N_10008,N_9683,N_9704);
nand U10009 (N_10009,N_9034,N_9562);
or U10010 (N_10010,N_9043,N_9248);
nor U10011 (N_10011,N_9343,N_9658);
nor U10012 (N_10012,N_9633,N_9362);
nor U10013 (N_10013,N_9169,N_9676);
and U10014 (N_10014,N_9272,N_9004);
nor U10015 (N_10015,N_9455,N_9593);
nand U10016 (N_10016,N_9005,N_9220);
and U10017 (N_10017,N_9083,N_9515);
and U10018 (N_10018,N_9185,N_9194);
xor U10019 (N_10019,N_9128,N_9520);
nand U10020 (N_10020,N_9534,N_9657);
and U10021 (N_10021,N_9548,N_9525);
nand U10022 (N_10022,N_9373,N_9400);
xnor U10023 (N_10023,N_9619,N_9660);
or U10024 (N_10024,N_9040,N_9518);
nand U10025 (N_10025,N_9391,N_9228);
and U10026 (N_10026,N_9337,N_9120);
xor U10027 (N_10027,N_9357,N_9687);
nor U10028 (N_10028,N_9328,N_9381);
and U10029 (N_10029,N_9614,N_9149);
or U10030 (N_10030,N_9684,N_9646);
or U10031 (N_10031,N_9648,N_9471);
nor U10032 (N_10032,N_9222,N_9627);
nor U10033 (N_10033,N_9401,N_9440);
nand U10034 (N_10034,N_9510,N_9245);
xor U10035 (N_10035,N_9264,N_9438);
nor U10036 (N_10036,N_9160,N_9585);
nand U10037 (N_10037,N_9318,N_9363);
nand U10038 (N_10038,N_9370,N_9334);
xnor U10039 (N_10039,N_9097,N_9310);
nand U10040 (N_10040,N_9303,N_9050);
or U10041 (N_10041,N_9659,N_9077);
or U10042 (N_10042,N_9736,N_9560);
nor U10043 (N_10043,N_9100,N_9112);
or U10044 (N_10044,N_9235,N_9458);
nand U10045 (N_10045,N_9270,N_9124);
or U10046 (N_10046,N_9500,N_9047);
nand U10047 (N_10047,N_9417,N_9223);
nand U10048 (N_10048,N_9217,N_9285);
nor U10049 (N_10049,N_9726,N_9045);
nand U10050 (N_10050,N_9130,N_9549);
xnor U10051 (N_10051,N_9542,N_9286);
nand U10052 (N_10052,N_9341,N_9301);
and U10053 (N_10053,N_9592,N_9163);
nand U10054 (N_10054,N_9580,N_9419);
nor U10055 (N_10055,N_9655,N_9436);
and U10056 (N_10056,N_9321,N_9232);
and U10057 (N_10057,N_9166,N_9566);
nand U10058 (N_10058,N_9261,N_9079);
or U10059 (N_10059,N_9721,N_9708);
and U10060 (N_10060,N_9148,N_9157);
nor U10061 (N_10061,N_9325,N_9540);
xnor U10062 (N_10062,N_9167,N_9484);
nand U10063 (N_10063,N_9132,N_9475);
nand U10064 (N_10064,N_9196,N_9557);
xor U10065 (N_10065,N_9461,N_9290);
nand U10066 (N_10066,N_9692,N_9701);
nand U10067 (N_10067,N_9324,N_9616);
nor U10068 (N_10068,N_9626,N_9214);
and U10069 (N_10069,N_9003,N_9739);
nor U10070 (N_10070,N_9114,N_9288);
and U10071 (N_10071,N_9187,N_9710);
nand U10072 (N_10072,N_9635,N_9336);
nand U10073 (N_10073,N_9493,N_9661);
nor U10074 (N_10074,N_9302,N_9230);
or U10075 (N_10075,N_9504,N_9380);
or U10076 (N_10076,N_9347,N_9263);
nor U10077 (N_10077,N_9405,N_9332);
nand U10078 (N_10078,N_9305,N_9146);
nand U10079 (N_10079,N_9517,N_9509);
xor U10080 (N_10080,N_9388,N_9021);
nand U10081 (N_10081,N_9656,N_9425);
nand U10082 (N_10082,N_9383,N_9567);
xor U10083 (N_10083,N_9598,N_9084);
and U10084 (N_10084,N_9331,N_9044);
xnor U10085 (N_10085,N_9116,N_9628);
or U10086 (N_10086,N_9027,N_9218);
and U10087 (N_10087,N_9058,N_9195);
nand U10088 (N_10088,N_9075,N_9236);
nand U10089 (N_10089,N_9309,N_9344);
and U10090 (N_10090,N_9734,N_9274);
nor U10091 (N_10091,N_9275,N_9345);
nor U10092 (N_10092,N_9249,N_9113);
xor U10093 (N_10093,N_9133,N_9002);
or U10094 (N_10094,N_9202,N_9224);
and U10095 (N_10095,N_9729,N_9521);
or U10096 (N_10096,N_9213,N_9603);
nand U10097 (N_10097,N_9514,N_9640);
xor U10098 (N_10098,N_9308,N_9010);
nand U10099 (N_10099,N_9723,N_9450);
nand U10100 (N_10100,N_9669,N_9260);
nand U10101 (N_10101,N_9429,N_9372);
nand U10102 (N_10102,N_9030,N_9446);
nand U10103 (N_10103,N_9287,N_9255);
nor U10104 (N_10104,N_9672,N_9722);
xor U10105 (N_10105,N_9480,N_9409);
or U10106 (N_10106,N_9105,N_9682);
and U10107 (N_10107,N_9086,N_9395);
or U10108 (N_10108,N_9178,N_9442);
xor U10109 (N_10109,N_9737,N_9016);
or U10110 (N_10110,N_9449,N_9014);
xnor U10111 (N_10111,N_9622,N_9361);
nor U10112 (N_10112,N_9162,N_9350);
nand U10113 (N_10113,N_9709,N_9642);
nor U10114 (N_10114,N_9277,N_9581);
nor U10115 (N_10115,N_9688,N_9568);
xor U10116 (N_10116,N_9406,N_9728);
xnor U10117 (N_10117,N_9618,N_9421);
nor U10118 (N_10118,N_9407,N_9176);
or U10119 (N_10119,N_9434,N_9393);
xnor U10120 (N_10120,N_9115,N_9608);
nand U10121 (N_10121,N_9055,N_9299);
nand U10122 (N_10122,N_9745,N_9312);
and U10123 (N_10123,N_9422,N_9694);
xnor U10124 (N_10124,N_9574,N_9577);
nor U10125 (N_10125,N_9149,N_9209);
xnor U10126 (N_10126,N_9251,N_9371);
xor U10127 (N_10127,N_9449,N_9676);
nor U10128 (N_10128,N_9543,N_9490);
and U10129 (N_10129,N_9277,N_9200);
or U10130 (N_10130,N_9276,N_9712);
or U10131 (N_10131,N_9319,N_9537);
xnor U10132 (N_10132,N_9389,N_9659);
xnor U10133 (N_10133,N_9391,N_9562);
xnor U10134 (N_10134,N_9524,N_9258);
xor U10135 (N_10135,N_9490,N_9148);
or U10136 (N_10136,N_9528,N_9196);
or U10137 (N_10137,N_9537,N_9361);
and U10138 (N_10138,N_9297,N_9466);
or U10139 (N_10139,N_9061,N_9448);
xnor U10140 (N_10140,N_9210,N_9725);
xnor U10141 (N_10141,N_9248,N_9632);
xnor U10142 (N_10142,N_9624,N_9551);
xnor U10143 (N_10143,N_9231,N_9628);
nand U10144 (N_10144,N_9287,N_9170);
nor U10145 (N_10145,N_9712,N_9602);
xnor U10146 (N_10146,N_9055,N_9075);
nor U10147 (N_10147,N_9729,N_9448);
nand U10148 (N_10148,N_9626,N_9091);
or U10149 (N_10149,N_9605,N_9550);
xnor U10150 (N_10150,N_9611,N_9590);
and U10151 (N_10151,N_9306,N_9349);
or U10152 (N_10152,N_9154,N_9506);
nor U10153 (N_10153,N_9144,N_9711);
and U10154 (N_10154,N_9664,N_9471);
or U10155 (N_10155,N_9471,N_9226);
or U10156 (N_10156,N_9353,N_9569);
and U10157 (N_10157,N_9192,N_9237);
xnor U10158 (N_10158,N_9481,N_9378);
xnor U10159 (N_10159,N_9434,N_9539);
or U10160 (N_10160,N_9503,N_9062);
and U10161 (N_10161,N_9014,N_9027);
nor U10162 (N_10162,N_9600,N_9417);
nor U10163 (N_10163,N_9345,N_9277);
xnor U10164 (N_10164,N_9009,N_9635);
xor U10165 (N_10165,N_9416,N_9012);
and U10166 (N_10166,N_9197,N_9522);
nor U10167 (N_10167,N_9349,N_9168);
or U10168 (N_10168,N_9374,N_9325);
and U10169 (N_10169,N_9391,N_9385);
nor U10170 (N_10170,N_9209,N_9321);
or U10171 (N_10171,N_9319,N_9267);
or U10172 (N_10172,N_9545,N_9028);
nand U10173 (N_10173,N_9671,N_9490);
and U10174 (N_10174,N_9148,N_9249);
nor U10175 (N_10175,N_9352,N_9623);
nor U10176 (N_10176,N_9493,N_9116);
or U10177 (N_10177,N_9122,N_9400);
nand U10178 (N_10178,N_9158,N_9549);
or U10179 (N_10179,N_9721,N_9406);
and U10180 (N_10180,N_9320,N_9361);
nand U10181 (N_10181,N_9622,N_9201);
nand U10182 (N_10182,N_9600,N_9685);
xor U10183 (N_10183,N_9406,N_9660);
and U10184 (N_10184,N_9389,N_9148);
nor U10185 (N_10185,N_9538,N_9748);
or U10186 (N_10186,N_9087,N_9251);
or U10187 (N_10187,N_9292,N_9596);
and U10188 (N_10188,N_9593,N_9211);
or U10189 (N_10189,N_9683,N_9616);
or U10190 (N_10190,N_9232,N_9565);
nand U10191 (N_10191,N_9646,N_9525);
xor U10192 (N_10192,N_9519,N_9254);
nor U10193 (N_10193,N_9281,N_9530);
nor U10194 (N_10194,N_9683,N_9249);
nor U10195 (N_10195,N_9608,N_9577);
and U10196 (N_10196,N_9194,N_9737);
nand U10197 (N_10197,N_9360,N_9354);
or U10198 (N_10198,N_9428,N_9182);
xnor U10199 (N_10199,N_9144,N_9220);
nor U10200 (N_10200,N_9452,N_9514);
nand U10201 (N_10201,N_9448,N_9674);
or U10202 (N_10202,N_9227,N_9344);
or U10203 (N_10203,N_9057,N_9253);
or U10204 (N_10204,N_9020,N_9014);
nand U10205 (N_10205,N_9556,N_9437);
and U10206 (N_10206,N_9158,N_9528);
or U10207 (N_10207,N_9184,N_9093);
nand U10208 (N_10208,N_9167,N_9647);
nor U10209 (N_10209,N_9583,N_9478);
xnor U10210 (N_10210,N_9663,N_9065);
or U10211 (N_10211,N_9281,N_9417);
and U10212 (N_10212,N_9307,N_9374);
nor U10213 (N_10213,N_9430,N_9235);
nand U10214 (N_10214,N_9278,N_9499);
nand U10215 (N_10215,N_9393,N_9048);
xor U10216 (N_10216,N_9271,N_9533);
and U10217 (N_10217,N_9350,N_9237);
and U10218 (N_10218,N_9315,N_9275);
nand U10219 (N_10219,N_9370,N_9236);
xnor U10220 (N_10220,N_9714,N_9612);
xnor U10221 (N_10221,N_9242,N_9552);
nor U10222 (N_10222,N_9198,N_9505);
nand U10223 (N_10223,N_9583,N_9167);
or U10224 (N_10224,N_9297,N_9102);
or U10225 (N_10225,N_9388,N_9547);
nand U10226 (N_10226,N_9553,N_9658);
xor U10227 (N_10227,N_9451,N_9459);
and U10228 (N_10228,N_9238,N_9098);
nor U10229 (N_10229,N_9540,N_9106);
or U10230 (N_10230,N_9466,N_9584);
nor U10231 (N_10231,N_9445,N_9720);
xor U10232 (N_10232,N_9364,N_9481);
xnor U10233 (N_10233,N_9687,N_9277);
or U10234 (N_10234,N_9634,N_9003);
nor U10235 (N_10235,N_9056,N_9300);
or U10236 (N_10236,N_9329,N_9702);
or U10237 (N_10237,N_9677,N_9295);
xor U10238 (N_10238,N_9508,N_9278);
nand U10239 (N_10239,N_9101,N_9699);
nor U10240 (N_10240,N_9062,N_9704);
nor U10241 (N_10241,N_9444,N_9343);
and U10242 (N_10242,N_9206,N_9385);
nand U10243 (N_10243,N_9685,N_9099);
xor U10244 (N_10244,N_9265,N_9609);
nand U10245 (N_10245,N_9380,N_9329);
nor U10246 (N_10246,N_9234,N_9025);
and U10247 (N_10247,N_9017,N_9627);
xor U10248 (N_10248,N_9289,N_9129);
or U10249 (N_10249,N_9099,N_9439);
and U10250 (N_10250,N_9508,N_9258);
and U10251 (N_10251,N_9569,N_9280);
and U10252 (N_10252,N_9104,N_9490);
and U10253 (N_10253,N_9000,N_9280);
and U10254 (N_10254,N_9404,N_9563);
and U10255 (N_10255,N_9585,N_9521);
and U10256 (N_10256,N_9601,N_9716);
or U10257 (N_10257,N_9225,N_9087);
xnor U10258 (N_10258,N_9708,N_9711);
or U10259 (N_10259,N_9675,N_9636);
or U10260 (N_10260,N_9486,N_9335);
and U10261 (N_10261,N_9643,N_9722);
or U10262 (N_10262,N_9535,N_9720);
nand U10263 (N_10263,N_9025,N_9444);
xnor U10264 (N_10264,N_9374,N_9187);
xnor U10265 (N_10265,N_9081,N_9170);
xor U10266 (N_10266,N_9491,N_9703);
nand U10267 (N_10267,N_9422,N_9110);
and U10268 (N_10268,N_9047,N_9068);
nor U10269 (N_10269,N_9416,N_9098);
nand U10270 (N_10270,N_9486,N_9209);
nor U10271 (N_10271,N_9530,N_9156);
nor U10272 (N_10272,N_9623,N_9102);
or U10273 (N_10273,N_9169,N_9277);
and U10274 (N_10274,N_9546,N_9137);
xnor U10275 (N_10275,N_9223,N_9585);
nand U10276 (N_10276,N_9344,N_9459);
nor U10277 (N_10277,N_9314,N_9159);
and U10278 (N_10278,N_9025,N_9467);
and U10279 (N_10279,N_9283,N_9678);
xnor U10280 (N_10280,N_9467,N_9069);
and U10281 (N_10281,N_9170,N_9146);
xor U10282 (N_10282,N_9640,N_9335);
and U10283 (N_10283,N_9199,N_9163);
nor U10284 (N_10284,N_9377,N_9337);
nand U10285 (N_10285,N_9265,N_9343);
and U10286 (N_10286,N_9411,N_9061);
or U10287 (N_10287,N_9424,N_9337);
or U10288 (N_10288,N_9231,N_9389);
nand U10289 (N_10289,N_9462,N_9681);
xor U10290 (N_10290,N_9366,N_9570);
nand U10291 (N_10291,N_9358,N_9406);
and U10292 (N_10292,N_9143,N_9594);
nand U10293 (N_10293,N_9454,N_9558);
xnor U10294 (N_10294,N_9260,N_9383);
or U10295 (N_10295,N_9554,N_9108);
nor U10296 (N_10296,N_9299,N_9296);
nand U10297 (N_10297,N_9294,N_9176);
nor U10298 (N_10298,N_9391,N_9329);
or U10299 (N_10299,N_9555,N_9339);
and U10300 (N_10300,N_9475,N_9207);
or U10301 (N_10301,N_9227,N_9090);
nand U10302 (N_10302,N_9636,N_9314);
nand U10303 (N_10303,N_9427,N_9550);
nor U10304 (N_10304,N_9412,N_9392);
or U10305 (N_10305,N_9350,N_9592);
nand U10306 (N_10306,N_9271,N_9557);
xor U10307 (N_10307,N_9157,N_9343);
xor U10308 (N_10308,N_9681,N_9374);
xnor U10309 (N_10309,N_9151,N_9387);
xnor U10310 (N_10310,N_9432,N_9193);
xnor U10311 (N_10311,N_9244,N_9426);
or U10312 (N_10312,N_9387,N_9169);
or U10313 (N_10313,N_9027,N_9686);
nand U10314 (N_10314,N_9094,N_9647);
and U10315 (N_10315,N_9659,N_9164);
nand U10316 (N_10316,N_9246,N_9360);
and U10317 (N_10317,N_9458,N_9628);
or U10318 (N_10318,N_9698,N_9182);
and U10319 (N_10319,N_9746,N_9190);
or U10320 (N_10320,N_9341,N_9290);
xor U10321 (N_10321,N_9425,N_9667);
nor U10322 (N_10322,N_9284,N_9397);
nor U10323 (N_10323,N_9677,N_9673);
nor U10324 (N_10324,N_9299,N_9670);
nor U10325 (N_10325,N_9085,N_9459);
xnor U10326 (N_10326,N_9672,N_9565);
nand U10327 (N_10327,N_9142,N_9621);
nor U10328 (N_10328,N_9600,N_9675);
and U10329 (N_10329,N_9376,N_9422);
nand U10330 (N_10330,N_9274,N_9113);
nand U10331 (N_10331,N_9609,N_9042);
nor U10332 (N_10332,N_9531,N_9665);
nand U10333 (N_10333,N_9743,N_9146);
nand U10334 (N_10334,N_9692,N_9422);
nand U10335 (N_10335,N_9369,N_9093);
or U10336 (N_10336,N_9564,N_9674);
nand U10337 (N_10337,N_9592,N_9630);
xor U10338 (N_10338,N_9696,N_9729);
nand U10339 (N_10339,N_9334,N_9167);
xnor U10340 (N_10340,N_9100,N_9297);
nor U10341 (N_10341,N_9244,N_9164);
nand U10342 (N_10342,N_9434,N_9304);
and U10343 (N_10343,N_9047,N_9086);
nor U10344 (N_10344,N_9304,N_9545);
or U10345 (N_10345,N_9037,N_9227);
nand U10346 (N_10346,N_9628,N_9188);
or U10347 (N_10347,N_9643,N_9114);
nand U10348 (N_10348,N_9349,N_9232);
xor U10349 (N_10349,N_9523,N_9406);
xnor U10350 (N_10350,N_9523,N_9173);
or U10351 (N_10351,N_9507,N_9538);
and U10352 (N_10352,N_9710,N_9283);
or U10353 (N_10353,N_9164,N_9499);
xnor U10354 (N_10354,N_9204,N_9579);
or U10355 (N_10355,N_9197,N_9690);
nand U10356 (N_10356,N_9312,N_9119);
or U10357 (N_10357,N_9414,N_9706);
and U10358 (N_10358,N_9598,N_9592);
and U10359 (N_10359,N_9375,N_9251);
and U10360 (N_10360,N_9410,N_9082);
nor U10361 (N_10361,N_9347,N_9741);
xnor U10362 (N_10362,N_9622,N_9625);
and U10363 (N_10363,N_9412,N_9037);
xnor U10364 (N_10364,N_9641,N_9184);
xnor U10365 (N_10365,N_9409,N_9120);
and U10366 (N_10366,N_9468,N_9383);
xnor U10367 (N_10367,N_9375,N_9264);
nand U10368 (N_10368,N_9185,N_9603);
nand U10369 (N_10369,N_9616,N_9548);
and U10370 (N_10370,N_9135,N_9059);
nor U10371 (N_10371,N_9036,N_9522);
or U10372 (N_10372,N_9494,N_9720);
nor U10373 (N_10373,N_9381,N_9472);
nor U10374 (N_10374,N_9306,N_9718);
xnor U10375 (N_10375,N_9018,N_9698);
xor U10376 (N_10376,N_9238,N_9258);
or U10377 (N_10377,N_9598,N_9280);
nor U10378 (N_10378,N_9119,N_9020);
nor U10379 (N_10379,N_9181,N_9273);
nor U10380 (N_10380,N_9482,N_9084);
nor U10381 (N_10381,N_9289,N_9676);
xor U10382 (N_10382,N_9099,N_9207);
or U10383 (N_10383,N_9573,N_9380);
or U10384 (N_10384,N_9347,N_9531);
nor U10385 (N_10385,N_9465,N_9390);
xor U10386 (N_10386,N_9648,N_9618);
or U10387 (N_10387,N_9148,N_9194);
and U10388 (N_10388,N_9155,N_9647);
xor U10389 (N_10389,N_9076,N_9560);
xnor U10390 (N_10390,N_9135,N_9464);
xor U10391 (N_10391,N_9227,N_9408);
xnor U10392 (N_10392,N_9679,N_9749);
xnor U10393 (N_10393,N_9257,N_9332);
nand U10394 (N_10394,N_9735,N_9439);
and U10395 (N_10395,N_9675,N_9369);
and U10396 (N_10396,N_9289,N_9229);
and U10397 (N_10397,N_9374,N_9526);
nor U10398 (N_10398,N_9534,N_9137);
nand U10399 (N_10399,N_9719,N_9720);
xor U10400 (N_10400,N_9664,N_9718);
or U10401 (N_10401,N_9093,N_9691);
nand U10402 (N_10402,N_9531,N_9717);
or U10403 (N_10403,N_9713,N_9324);
xor U10404 (N_10404,N_9567,N_9729);
and U10405 (N_10405,N_9061,N_9425);
nand U10406 (N_10406,N_9303,N_9389);
nand U10407 (N_10407,N_9174,N_9276);
nand U10408 (N_10408,N_9385,N_9393);
nor U10409 (N_10409,N_9703,N_9706);
xnor U10410 (N_10410,N_9482,N_9687);
and U10411 (N_10411,N_9027,N_9236);
nand U10412 (N_10412,N_9253,N_9704);
nand U10413 (N_10413,N_9238,N_9534);
nand U10414 (N_10414,N_9397,N_9444);
or U10415 (N_10415,N_9702,N_9185);
nand U10416 (N_10416,N_9330,N_9429);
nand U10417 (N_10417,N_9499,N_9039);
nor U10418 (N_10418,N_9446,N_9599);
or U10419 (N_10419,N_9023,N_9390);
nand U10420 (N_10420,N_9337,N_9131);
or U10421 (N_10421,N_9026,N_9373);
nor U10422 (N_10422,N_9169,N_9439);
xnor U10423 (N_10423,N_9412,N_9680);
and U10424 (N_10424,N_9566,N_9408);
or U10425 (N_10425,N_9700,N_9005);
or U10426 (N_10426,N_9173,N_9133);
and U10427 (N_10427,N_9240,N_9394);
or U10428 (N_10428,N_9278,N_9370);
or U10429 (N_10429,N_9295,N_9682);
nand U10430 (N_10430,N_9096,N_9566);
nor U10431 (N_10431,N_9634,N_9340);
and U10432 (N_10432,N_9088,N_9569);
xor U10433 (N_10433,N_9644,N_9039);
or U10434 (N_10434,N_9269,N_9200);
nand U10435 (N_10435,N_9687,N_9282);
xor U10436 (N_10436,N_9253,N_9161);
xor U10437 (N_10437,N_9607,N_9158);
nor U10438 (N_10438,N_9315,N_9231);
nand U10439 (N_10439,N_9091,N_9040);
xor U10440 (N_10440,N_9497,N_9469);
or U10441 (N_10441,N_9195,N_9510);
nor U10442 (N_10442,N_9090,N_9230);
and U10443 (N_10443,N_9265,N_9542);
or U10444 (N_10444,N_9247,N_9686);
nor U10445 (N_10445,N_9403,N_9629);
nor U10446 (N_10446,N_9379,N_9266);
nand U10447 (N_10447,N_9605,N_9397);
nand U10448 (N_10448,N_9388,N_9134);
nor U10449 (N_10449,N_9711,N_9324);
or U10450 (N_10450,N_9724,N_9266);
nand U10451 (N_10451,N_9255,N_9482);
nor U10452 (N_10452,N_9033,N_9321);
nand U10453 (N_10453,N_9099,N_9669);
or U10454 (N_10454,N_9230,N_9435);
or U10455 (N_10455,N_9243,N_9594);
nor U10456 (N_10456,N_9526,N_9664);
nor U10457 (N_10457,N_9051,N_9587);
nor U10458 (N_10458,N_9125,N_9276);
or U10459 (N_10459,N_9236,N_9241);
nand U10460 (N_10460,N_9315,N_9485);
and U10461 (N_10461,N_9482,N_9258);
nand U10462 (N_10462,N_9639,N_9561);
nor U10463 (N_10463,N_9459,N_9534);
xnor U10464 (N_10464,N_9121,N_9615);
nor U10465 (N_10465,N_9121,N_9570);
nand U10466 (N_10466,N_9252,N_9520);
or U10467 (N_10467,N_9721,N_9352);
nor U10468 (N_10468,N_9603,N_9639);
nand U10469 (N_10469,N_9248,N_9613);
xnor U10470 (N_10470,N_9410,N_9369);
nor U10471 (N_10471,N_9748,N_9603);
nor U10472 (N_10472,N_9246,N_9602);
xor U10473 (N_10473,N_9152,N_9449);
nand U10474 (N_10474,N_9380,N_9625);
nor U10475 (N_10475,N_9250,N_9670);
xnor U10476 (N_10476,N_9056,N_9041);
and U10477 (N_10477,N_9085,N_9045);
nand U10478 (N_10478,N_9336,N_9365);
nand U10479 (N_10479,N_9545,N_9085);
nand U10480 (N_10480,N_9689,N_9120);
and U10481 (N_10481,N_9222,N_9598);
and U10482 (N_10482,N_9120,N_9043);
nor U10483 (N_10483,N_9434,N_9139);
nand U10484 (N_10484,N_9129,N_9004);
xor U10485 (N_10485,N_9691,N_9646);
nand U10486 (N_10486,N_9041,N_9718);
nor U10487 (N_10487,N_9594,N_9160);
xnor U10488 (N_10488,N_9650,N_9520);
nand U10489 (N_10489,N_9466,N_9507);
and U10490 (N_10490,N_9296,N_9252);
nand U10491 (N_10491,N_9429,N_9195);
or U10492 (N_10492,N_9513,N_9195);
xnor U10493 (N_10493,N_9214,N_9093);
and U10494 (N_10494,N_9708,N_9109);
and U10495 (N_10495,N_9193,N_9615);
nor U10496 (N_10496,N_9525,N_9014);
xnor U10497 (N_10497,N_9404,N_9098);
or U10498 (N_10498,N_9048,N_9391);
nand U10499 (N_10499,N_9691,N_9699);
nand U10500 (N_10500,N_9883,N_10200);
xnor U10501 (N_10501,N_9989,N_10280);
or U10502 (N_10502,N_10185,N_10124);
and U10503 (N_10503,N_10442,N_10339);
nor U10504 (N_10504,N_10343,N_10108);
nand U10505 (N_10505,N_10315,N_10444);
and U10506 (N_10506,N_9938,N_10173);
nor U10507 (N_10507,N_10325,N_9875);
or U10508 (N_10508,N_9904,N_9873);
xor U10509 (N_10509,N_10311,N_9854);
nand U10510 (N_10510,N_9998,N_9830);
nor U10511 (N_10511,N_10133,N_9850);
or U10512 (N_10512,N_9943,N_10475);
nor U10513 (N_10513,N_10372,N_10143);
or U10514 (N_10514,N_10091,N_10050);
xnor U10515 (N_10515,N_10429,N_10430);
nand U10516 (N_10516,N_10121,N_10090);
nor U10517 (N_10517,N_10456,N_9800);
nand U10518 (N_10518,N_10150,N_10135);
xor U10519 (N_10519,N_10335,N_10453);
or U10520 (N_10520,N_9769,N_10345);
nor U10521 (N_10521,N_10243,N_9765);
and U10522 (N_10522,N_9892,N_9999);
nor U10523 (N_10523,N_10228,N_9864);
or U10524 (N_10524,N_10419,N_10403);
and U10525 (N_10525,N_10418,N_10162);
or U10526 (N_10526,N_10235,N_10136);
nand U10527 (N_10527,N_10175,N_9823);
xor U10528 (N_10528,N_10066,N_9751);
or U10529 (N_10529,N_9799,N_9960);
and U10530 (N_10530,N_9896,N_10396);
nand U10531 (N_10531,N_10320,N_10313);
nand U10532 (N_10532,N_10354,N_10151);
nor U10533 (N_10533,N_10349,N_10237);
or U10534 (N_10534,N_10160,N_10476);
xnor U10535 (N_10535,N_10045,N_9819);
or U10536 (N_10536,N_10131,N_10473);
nor U10537 (N_10537,N_9940,N_9956);
nand U10538 (N_10538,N_9847,N_10415);
nor U10539 (N_10539,N_10125,N_10461);
xnor U10540 (N_10540,N_10348,N_9821);
xnor U10541 (N_10541,N_10364,N_9889);
nor U10542 (N_10542,N_10431,N_10283);
nand U10543 (N_10543,N_10405,N_9959);
nand U10544 (N_10544,N_10267,N_9764);
xnor U10545 (N_10545,N_10326,N_9796);
and U10546 (N_10546,N_10103,N_9802);
and U10547 (N_10547,N_9907,N_9891);
nand U10548 (N_10548,N_10174,N_10384);
nor U10549 (N_10549,N_10460,N_9981);
nor U10550 (N_10550,N_9818,N_10255);
or U10551 (N_10551,N_10044,N_10229);
nand U10552 (N_10552,N_10035,N_10296);
and U10553 (N_10553,N_9951,N_9795);
nor U10554 (N_10554,N_9852,N_9817);
xnor U10555 (N_10555,N_9857,N_10117);
nand U10556 (N_10556,N_10282,N_10164);
and U10557 (N_10557,N_10240,N_10203);
and U10558 (N_10558,N_10299,N_9978);
nand U10559 (N_10559,N_10012,N_9969);
xor U10560 (N_10560,N_10395,N_10141);
nor U10561 (N_10561,N_10491,N_10201);
and U10562 (N_10562,N_9828,N_9897);
xnor U10563 (N_10563,N_10365,N_10382);
and U10564 (N_10564,N_10184,N_10060);
xor U10565 (N_10565,N_10191,N_9779);
and U10566 (N_10566,N_10104,N_9901);
nand U10567 (N_10567,N_10197,N_10290);
or U10568 (N_10568,N_10347,N_9871);
nand U10569 (N_10569,N_10061,N_10353);
xnor U10570 (N_10570,N_10195,N_9895);
nor U10571 (N_10571,N_9813,N_10176);
nor U10572 (N_10572,N_10079,N_9804);
or U10573 (N_10573,N_9816,N_9899);
nand U10574 (N_10574,N_10161,N_10234);
nor U10575 (N_10575,N_9803,N_10378);
xor U10576 (N_10576,N_10149,N_10084);
nand U10577 (N_10577,N_10190,N_10294);
nand U10578 (N_10578,N_10186,N_9964);
nand U10579 (N_10579,N_10206,N_10020);
nor U10580 (N_10580,N_10011,N_10192);
or U10581 (N_10581,N_9851,N_10497);
nor U10582 (N_10582,N_9842,N_10328);
and U10583 (N_10583,N_9811,N_9945);
and U10584 (N_10584,N_10379,N_10029);
xor U10585 (N_10585,N_10427,N_10134);
nand U10586 (N_10586,N_9988,N_10163);
nor U10587 (N_10587,N_9877,N_10227);
nand U10588 (N_10588,N_9972,N_10244);
nand U10589 (N_10589,N_10356,N_10248);
and U10590 (N_10590,N_9844,N_9922);
nor U10591 (N_10591,N_10252,N_9924);
and U10592 (N_10592,N_9954,N_9880);
xnor U10593 (N_10593,N_10441,N_9784);
nand U10594 (N_10594,N_9782,N_10447);
or U10595 (N_10595,N_9771,N_10152);
nor U10596 (N_10596,N_10231,N_10038);
xor U10597 (N_10597,N_10346,N_10119);
xor U10598 (N_10598,N_10073,N_10309);
or U10599 (N_10599,N_9820,N_10445);
xor U10600 (N_10600,N_10097,N_10170);
nand U10601 (N_10601,N_10211,N_10145);
nand U10602 (N_10602,N_10049,N_10128);
or U10603 (N_10603,N_10452,N_10142);
nand U10604 (N_10604,N_9787,N_9831);
and U10605 (N_10605,N_10178,N_9843);
nor U10606 (N_10606,N_9867,N_10218);
and U10607 (N_10607,N_9773,N_10426);
and U10608 (N_10608,N_9991,N_10017);
xor U10609 (N_10609,N_10433,N_10024);
or U10610 (N_10610,N_10193,N_9866);
or U10611 (N_10611,N_9761,N_10407);
nand U10612 (N_10612,N_9996,N_10261);
nor U10613 (N_10613,N_10048,N_10167);
or U10614 (N_10614,N_10479,N_10494);
nor U10615 (N_10615,N_10392,N_10490);
and U10616 (N_10616,N_10391,N_9947);
xnor U10617 (N_10617,N_9993,N_10041);
nor U10618 (N_10618,N_10398,N_9815);
nand U10619 (N_10619,N_10249,N_9965);
or U10620 (N_10620,N_10068,N_9801);
and U10621 (N_10621,N_10139,N_10324);
nand U10622 (N_10622,N_10010,N_10153);
or U10623 (N_10623,N_10300,N_10291);
and U10624 (N_10624,N_9810,N_10110);
or U10625 (N_10625,N_9797,N_10417);
xnor U10626 (N_10626,N_9832,N_10375);
nand U10627 (N_10627,N_10387,N_10388);
nand U10628 (N_10628,N_10102,N_10069);
nand U10629 (N_10629,N_9794,N_10113);
or U10630 (N_10630,N_9923,N_10308);
and U10631 (N_10631,N_10159,N_10306);
and U10632 (N_10632,N_10363,N_10223);
and U10633 (N_10633,N_9992,N_10230);
and U10634 (N_10634,N_10389,N_10368);
xnor U10635 (N_10635,N_10006,N_10487);
or U10636 (N_10636,N_10137,N_9903);
and U10637 (N_10637,N_9775,N_10087);
nand U10638 (N_10638,N_9848,N_10123);
or U10639 (N_10639,N_9925,N_9882);
or U10640 (N_10640,N_9872,N_10086);
nand U10641 (N_10641,N_10478,N_10138);
xnor U10642 (N_10642,N_10471,N_9911);
nor U10643 (N_10643,N_10007,N_10242);
or U10644 (N_10644,N_10014,N_9772);
xnor U10645 (N_10645,N_10495,N_9939);
nor U10646 (N_10646,N_10381,N_9783);
or U10647 (N_10647,N_10366,N_10472);
nand U10648 (N_10648,N_10156,N_10120);
xor U10649 (N_10649,N_10101,N_9929);
nand U10650 (N_10650,N_10221,N_9827);
xor U10651 (N_10651,N_10093,N_10115);
or U10652 (N_10652,N_10224,N_10344);
or U10653 (N_10653,N_10266,N_10030);
and U10654 (N_10654,N_9862,N_9760);
nand U10655 (N_10655,N_10168,N_10371);
xnor U10656 (N_10656,N_10199,N_10043);
and U10657 (N_10657,N_9807,N_10004);
xor U10658 (N_10658,N_10358,N_9789);
and U10659 (N_10659,N_9752,N_9825);
or U10660 (N_10660,N_10361,N_9754);
xor U10661 (N_10661,N_10039,N_10287);
or U10662 (N_10662,N_9997,N_10023);
xor U10663 (N_10663,N_9905,N_10385);
xnor U10664 (N_10664,N_10263,N_10466);
nor U10665 (N_10665,N_9791,N_10307);
nand U10666 (N_10666,N_10336,N_10327);
or U10667 (N_10667,N_9890,N_9868);
nand U10668 (N_10668,N_9987,N_10028);
xnor U10669 (N_10669,N_9906,N_9898);
nand U10670 (N_10670,N_10107,N_9888);
nand U10671 (N_10671,N_10303,N_10081);
nand U10672 (N_10672,N_10155,N_10122);
xor U10673 (N_10673,N_10496,N_10067);
nand U10674 (N_10674,N_10063,N_10411);
nand U10675 (N_10675,N_10250,N_10438);
nand U10676 (N_10676,N_10443,N_9946);
or U10677 (N_10677,N_10077,N_9753);
or U10678 (N_10678,N_10446,N_10436);
xnor U10679 (N_10679,N_10292,N_10009);
nor U10680 (N_10680,N_9930,N_9927);
xnor U10681 (N_10681,N_10390,N_10027);
and U10682 (N_10682,N_10312,N_10106);
nor U10683 (N_10683,N_10359,N_10148);
and U10684 (N_10684,N_9975,N_9756);
or U10685 (N_10685,N_10402,N_9958);
xnor U10686 (N_10686,N_10099,N_9759);
nor U10687 (N_10687,N_10207,N_10220);
nand U10688 (N_10688,N_10051,N_9837);
nor U10689 (N_10689,N_10275,N_10321);
and U10690 (N_10690,N_10377,N_9912);
xor U10691 (N_10691,N_10253,N_10268);
and U10692 (N_10692,N_9824,N_9928);
nor U10693 (N_10693,N_10485,N_10474);
nor U10694 (N_10694,N_10406,N_10373);
xnor U10695 (N_10695,N_10219,N_10065);
xnor U10696 (N_10696,N_10208,N_10042);
nor U10697 (N_10697,N_9983,N_10092);
or U10698 (N_10698,N_10053,N_10468);
or U10699 (N_10699,N_9786,N_9962);
nand U10700 (N_10700,N_10214,N_9944);
or U10701 (N_10701,N_10022,N_10074);
and U10702 (N_10702,N_9841,N_10037);
and U10703 (N_10703,N_9846,N_10424);
or U10704 (N_10704,N_9974,N_10129);
nand U10705 (N_10705,N_9835,N_10238);
xnor U10706 (N_10706,N_10305,N_10459);
nand U10707 (N_10707,N_10058,N_10034);
and U10708 (N_10708,N_10181,N_10467);
and U10709 (N_10709,N_9840,N_9879);
or U10710 (N_10710,N_10260,N_10409);
or U10711 (N_10711,N_10054,N_9984);
xnor U10712 (N_10712,N_10357,N_10055);
xnor U10713 (N_10713,N_10286,N_9781);
xor U10714 (N_10714,N_10188,N_9986);
or U10715 (N_10715,N_9788,N_10257);
xnor U10716 (N_10716,N_10413,N_9919);
nand U10717 (N_10717,N_10450,N_10410);
or U10718 (N_10718,N_10075,N_9878);
or U10719 (N_10719,N_10408,N_10481);
or U10720 (N_10720,N_9806,N_10013);
xor U10721 (N_10721,N_9778,N_10322);
nand U10722 (N_10722,N_10350,N_10165);
nand U10723 (N_10723,N_10241,N_10019);
nor U10724 (N_10724,N_10435,N_10177);
nand U10725 (N_10725,N_9913,N_10222);
nor U10726 (N_10726,N_10302,N_10140);
nor U10727 (N_10727,N_10293,N_10032);
and U10728 (N_10728,N_9853,N_9900);
xnor U10729 (N_10729,N_9766,N_10209);
or U10730 (N_10730,N_10018,N_10454);
or U10731 (N_10731,N_10338,N_10130);
and U10732 (N_10732,N_10329,N_10289);
nor U10733 (N_10733,N_10215,N_10341);
or U10734 (N_10734,N_10298,N_9793);
or U10735 (N_10735,N_9833,N_9948);
nand U10736 (N_10736,N_10171,N_10047);
nor U10737 (N_10737,N_9910,N_10166);
xor U10738 (N_10738,N_9822,N_9750);
or U10739 (N_10739,N_9834,N_10132);
xnor U10740 (N_10740,N_10146,N_10493);
nand U10741 (N_10741,N_9968,N_10112);
and U10742 (N_10742,N_10273,N_10265);
nand U10743 (N_10743,N_10380,N_9870);
nand U10744 (N_10744,N_10455,N_9836);
nor U10745 (N_10745,N_10025,N_9957);
xnor U10746 (N_10746,N_10272,N_10182);
xor U10747 (N_10747,N_10310,N_9770);
nor U10748 (N_10748,N_9942,N_10469);
xor U10749 (N_10749,N_9926,N_9776);
nand U10750 (N_10750,N_9894,N_10434);
or U10751 (N_10751,N_10276,N_10154);
or U10752 (N_10752,N_9861,N_10016);
nor U10753 (N_10753,N_10204,N_9829);
nor U10754 (N_10754,N_10334,N_10369);
and U10755 (N_10755,N_10072,N_9885);
nor U10756 (N_10756,N_10367,N_9990);
and U10757 (N_10757,N_10439,N_10233);
and U10758 (N_10758,N_10111,N_9921);
or U10759 (N_10759,N_9982,N_9994);
xor U10760 (N_10760,N_9808,N_10499);
nand U10761 (N_10761,N_10394,N_10202);
or U10762 (N_10762,N_10180,N_10089);
and U10763 (N_10763,N_10437,N_9767);
nand U10764 (N_10764,N_10096,N_9839);
nand U10765 (N_10765,N_9845,N_10082);
and U10766 (N_10766,N_9869,N_10210);
nand U10767 (N_10767,N_10217,N_10008);
nor U10768 (N_10768,N_10330,N_10465);
xnor U10769 (N_10769,N_10458,N_10127);
nor U10770 (N_10770,N_10064,N_10340);
and U10771 (N_10771,N_9953,N_10251);
or U10772 (N_10772,N_10337,N_9961);
nor U10773 (N_10773,N_10071,N_9995);
xnor U10774 (N_10774,N_9774,N_10301);
xnor U10775 (N_10775,N_9763,N_10374);
nand U10776 (N_10776,N_10126,N_9812);
xor U10777 (N_10777,N_9952,N_10351);
xor U10778 (N_10778,N_10259,N_10040);
nand U10779 (N_10779,N_9935,N_10318);
xor U10780 (N_10780,N_10271,N_10057);
xor U10781 (N_10781,N_10056,N_9790);
nor U10782 (N_10782,N_10488,N_9884);
and U10783 (N_10783,N_10059,N_10297);
nand U10784 (N_10784,N_10036,N_10278);
nor U10785 (N_10785,N_10383,N_10236);
and U10786 (N_10786,N_9967,N_10046);
or U10787 (N_10787,N_9963,N_10205);
xor U10788 (N_10788,N_10212,N_10246);
nor U10789 (N_10789,N_9886,N_10393);
nor U10790 (N_10790,N_9932,N_10225);
xnor U10791 (N_10791,N_10247,N_9863);
or U10792 (N_10792,N_9934,N_10425);
or U10793 (N_10793,N_10331,N_9874);
and U10794 (N_10794,N_10031,N_9809);
and U10795 (N_10795,N_9971,N_10109);
xor U10796 (N_10796,N_9918,N_10457);
and U10797 (N_10797,N_9893,N_9858);
nor U10798 (N_10798,N_10464,N_10015);
xor U10799 (N_10799,N_10095,N_10187);
nand U10800 (N_10800,N_10486,N_10021);
and U10801 (N_10801,N_10470,N_10232);
and U10802 (N_10802,N_10342,N_10480);
nor U10803 (N_10803,N_10094,N_9950);
xnor U10804 (N_10804,N_10428,N_10269);
or U10805 (N_10805,N_9976,N_10404);
xnor U10806 (N_10806,N_10304,N_10362);
nor U10807 (N_10807,N_10370,N_10001);
and U10808 (N_10808,N_10158,N_10194);
nand U10809 (N_10809,N_9936,N_10451);
xor U10810 (N_10810,N_10105,N_10264);
nand U10811 (N_10811,N_9762,N_10005);
or U10812 (N_10812,N_10295,N_10003);
nand U10813 (N_10813,N_9785,N_9920);
or U10814 (N_10814,N_10198,N_9859);
nor U10815 (N_10815,N_10277,N_10245);
xor U10816 (N_10816,N_10423,N_9856);
nand U10817 (N_10817,N_10098,N_9915);
and U10818 (N_10818,N_9973,N_10449);
nor U10819 (N_10819,N_10477,N_9792);
nor U10820 (N_10820,N_10400,N_9805);
and U10821 (N_10821,N_10114,N_10397);
nand U10822 (N_10822,N_10157,N_9909);
nand U10823 (N_10823,N_10033,N_10213);
nand U10824 (N_10824,N_10483,N_10189);
xor U10825 (N_10825,N_10262,N_10216);
or U10826 (N_10826,N_9931,N_10002);
nor U10827 (N_10827,N_10323,N_10448);
or U10828 (N_10828,N_9876,N_10416);
nor U10829 (N_10829,N_10078,N_9768);
nand U10830 (N_10830,N_9955,N_9966);
or U10831 (N_10831,N_10279,N_9758);
or U10832 (N_10832,N_10281,N_10412);
xor U10833 (N_10833,N_9979,N_10144);
or U10834 (N_10834,N_10088,N_10258);
and U10835 (N_10835,N_9937,N_9881);
nor U10836 (N_10836,N_10026,N_10355);
or U10837 (N_10837,N_10314,N_10254);
or U10838 (N_10838,N_10256,N_10116);
nand U10839 (N_10839,N_9977,N_10274);
nor U10840 (N_10840,N_10000,N_10076);
nand U10841 (N_10841,N_10360,N_9902);
and U10842 (N_10842,N_10432,N_10463);
or U10843 (N_10843,N_9941,N_9777);
and U10844 (N_10844,N_10179,N_10062);
nor U10845 (N_10845,N_9887,N_10482);
nand U10846 (N_10846,N_9757,N_9933);
xnor U10847 (N_10847,N_10352,N_10376);
nand U10848 (N_10848,N_10440,N_10462);
nand U10849 (N_10849,N_9860,N_10332);
and U10850 (N_10850,N_10316,N_9916);
xor U10851 (N_10851,N_9970,N_10319);
nor U10852 (N_10852,N_9908,N_10085);
and U10853 (N_10853,N_10489,N_10118);
xnor U10854 (N_10854,N_10288,N_10420);
nor U10855 (N_10855,N_9949,N_10421);
and U10856 (N_10856,N_9826,N_10492);
and U10857 (N_10857,N_9865,N_10414);
nand U10858 (N_10858,N_10172,N_9980);
xnor U10859 (N_10859,N_10270,N_10169);
nand U10860 (N_10860,N_9985,N_10484);
and U10861 (N_10861,N_10498,N_10083);
nor U10862 (N_10862,N_10052,N_9838);
xor U10863 (N_10863,N_10422,N_9855);
nand U10864 (N_10864,N_10399,N_10100);
nor U10865 (N_10865,N_10285,N_10386);
or U10866 (N_10866,N_10284,N_10239);
xor U10867 (N_10867,N_10317,N_10226);
nand U10868 (N_10868,N_10070,N_9798);
and U10869 (N_10869,N_9780,N_10401);
and U10870 (N_10870,N_9914,N_9755);
nor U10871 (N_10871,N_9814,N_10080);
or U10872 (N_10872,N_10196,N_9917);
and U10873 (N_10873,N_10333,N_9849);
and U10874 (N_10874,N_10147,N_10183);
nor U10875 (N_10875,N_10224,N_10208);
nor U10876 (N_10876,N_10434,N_10196);
xor U10877 (N_10877,N_9760,N_10490);
and U10878 (N_10878,N_10283,N_9775);
xor U10879 (N_10879,N_9987,N_10363);
and U10880 (N_10880,N_10205,N_10015);
nor U10881 (N_10881,N_10295,N_9752);
xnor U10882 (N_10882,N_10322,N_10136);
xor U10883 (N_10883,N_10481,N_10309);
nand U10884 (N_10884,N_10183,N_9882);
nor U10885 (N_10885,N_9767,N_10376);
nand U10886 (N_10886,N_10021,N_10372);
nor U10887 (N_10887,N_10115,N_10314);
xnor U10888 (N_10888,N_9836,N_9900);
and U10889 (N_10889,N_10032,N_10022);
and U10890 (N_10890,N_10448,N_9867);
or U10891 (N_10891,N_10382,N_10029);
xnor U10892 (N_10892,N_10389,N_10470);
nand U10893 (N_10893,N_10199,N_10103);
and U10894 (N_10894,N_10336,N_10319);
nor U10895 (N_10895,N_9982,N_10281);
nand U10896 (N_10896,N_10300,N_9924);
or U10897 (N_10897,N_10355,N_10005);
nor U10898 (N_10898,N_9802,N_10436);
and U10899 (N_10899,N_10313,N_9891);
nor U10900 (N_10900,N_10403,N_10133);
xor U10901 (N_10901,N_10360,N_9919);
or U10902 (N_10902,N_9979,N_9900);
nor U10903 (N_10903,N_9921,N_9905);
nand U10904 (N_10904,N_9985,N_9912);
and U10905 (N_10905,N_10153,N_10173);
nand U10906 (N_10906,N_10403,N_10241);
and U10907 (N_10907,N_10166,N_9897);
nand U10908 (N_10908,N_9902,N_10232);
and U10909 (N_10909,N_10165,N_9856);
or U10910 (N_10910,N_9835,N_9796);
or U10911 (N_10911,N_9939,N_9801);
or U10912 (N_10912,N_9876,N_9799);
nor U10913 (N_10913,N_10321,N_10242);
and U10914 (N_10914,N_10056,N_10354);
xnor U10915 (N_10915,N_9866,N_10143);
nor U10916 (N_10916,N_10055,N_9830);
or U10917 (N_10917,N_10390,N_10402);
or U10918 (N_10918,N_10412,N_9863);
nand U10919 (N_10919,N_10394,N_9840);
or U10920 (N_10920,N_9916,N_10095);
xnor U10921 (N_10921,N_10230,N_10270);
and U10922 (N_10922,N_10474,N_9802);
xnor U10923 (N_10923,N_9962,N_9815);
and U10924 (N_10924,N_9955,N_10414);
nand U10925 (N_10925,N_10342,N_10291);
nand U10926 (N_10926,N_10221,N_10311);
nor U10927 (N_10927,N_10038,N_9846);
and U10928 (N_10928,N_10218,N_10375);
nor U10929 (N_10929,N_10114,N_10199);
nand U10930 (N_10930,N_9835,N_9964);
xnor U10931 (N_10931,N_10388,N_9907);
nand U10932 (N_10932,N_9795,N_10349);
or U10933 (N_10933,N_10199,N_10063);
or U10934 (N_10934,N_10223,N_10117);
nand U10935 (N_10935,N_10248,N_10307);
and U10936 (N_10936,N_10308,N_10061);
nor U10937 (N_10937,N_10391,N_10420);
and U10938 (N_10938,N_9787,N_10160);
and U10939 (N_10939,N_10432,N_10401);
xor U10940 (N_10940,N_10363,N_10043);
or U10941 (N_10941,N_10093,N_9756);
nand U10942 (N_10942,N_10188,N_10268);
or U10943 (N_10943,N_10416,N_10184);
xnor U10944 (N_10944,N_10143,N_10371);
xnor U10945 (N_10945,N_9890,N_10408);
nor U10946 (N_10946,N_10465,N_10141);
and U10947 (N_10947,N_9821,N_10333);
and U10948 (N_10948,N_10098,N_10046);
and U10949 (N_10949,N_9905,N_10064);
nand U10950 (N_10950,N_10277,N_10113);
or U10951 (N_10951,N_9859,N_10116);
nand U10952 (N_10952,N_10100,N_10239);
xnor U10953 (N_10953,N_10198,N_10406);
nand U10954 (N_10954,N_10094,N_10057);
xnor U10955 (N_10955,N_10143,N_10359);
and U10956 (N_10956,N_9813,N_10455);
or U10957 (N_10957,N_9946,N_10111);
nand U10958 (N_10958,N_10180,N_10330);
nand U10959 (N_10959,N_10414,N_9824);
nand U10960 (N_10960,N_9916,N_10263);
nor U10961 (N_10961,N_10114,N_9893);
or U10962 (N_10962,N_10210,N_10116);
or U10963 (N_10963,N_10252,N_10346);
nand U10964 (N_10964,N_9976,N_10455);
nand U10965 (N_10965,N_10293,N_10071);
nand U10966 (N_10966,N_9838,N_10496);
xor U10967 (N_10967,N_10299,N_10139);
xnor U10968 (N_10968,N_9930,N_10204);
xor U10969 (N_10969,N_9896,N_10185);
nor U10970 (N_10970,N_9933,N_10430);
or U10971 (N_10971,N_9791,N_10300);
xor U10972 (N_10972,N_10483,N_9818);
and U10973 (N_10973,N_10156,N_10343);
and U10974 (N_10974,N_9923,N_9949);
nor U10975 (N_10975,N_9861,N_9885);
and U10976 (N_10976,N_10337,N_9920);
and U10977 (N_10977,N_9994,N_10405);
nand U10978 (N_10978,N_9814,N_10126);
xnor U10979 (N_10979,N_10429,N_9914);
and U10980 (N_10980,N_10162,N_10157);
or U10981 (N_10981,N_9813,N_10412);
or U10982 (N_10982,N_10190,N_10392);
nor U10983 (N_10983,N_10121,N_9858);
nor U10984 (N_10984,N_10477,N_10037);
or U10985 (N_10985,N_10435,N_10336);
and U10986 (N_10986,N_10408,N_10052);
or U10987 (N_10987,N_10216,N_9784);
nor U10988 (N_10988,N_10215,N_9911);
nor U10989 (N_10989,N_10146,N_9881);
xor U10990 (N_10990,N_9922,N_10496);
and U10991 (N_10991,N_9756,N_10324);
or U10992 (N_10992,N_9758,N_10180);
nor U10993 (N_10993,N_9992,N_10089);
nor U10994 (N_10994,N_10176,N_10199);
nand U10995 (N_10995,N_9907,N_10282);
and U10996 (N_10996,N_10422,N_9935);
and U10997 (N_10997,N_10030,N_9795);
xnor U10998 (N_10998,N_10140,N_9974);
nand U10999 (N_10999,N_10443,N_9782);
and U11000 (N_11000,N_10207,N_10119);
and U11001 (N_11001,N_9889,N_10086);
and U11002 (N_11002,N_9987,N_10418);
xnor U11003 (N_11003,N_10308,N_10012);
and U11004 (N_11004,N_10319,N_10203);
nor U11005 (N_11005,N_9962,N_10126);
nor U11006 (N_11006,N_10385,N_9916);
nor U11007 (N_11007,N_10333,N_10484);
nand U11008 (N_11008,N_10413,N_10205);
xor U11009 (N_11009,N_10405,N_10380);
nor U11010 (N_11010,N_9768,N_10437);
nand U11011 (N_11011,N_9983,N_9974);
nand U11012 (N_11012,N_10002,N_9879);
nor U11013 (N_11013,N_9835,N_9901);
or U11014 (N_11014,N_9754,N_10002);
or U11015 (N_11015,N_9822,N_9790);
or U11016 (N_11016,N_9788,N_10433);
nor U11017 (N_11017,N_10383,N_10476);
nor U11018 (N_11018,N_9952,N_10359);
xor U11019 (N_11019,N_10133,N_9864);
and U11020 (N_11020,N_9811,N_10037);
nor U11021 (N_11021,N_9784,N_10372);
xor U11022 (N_11022,N_10180,N_9762);
xor U11023 (N_11023,N_9954,N_10413);
nand U11024 (N_11024,N_10038,N_10105);
xor U11025 (N_11025,N_9762,N_10285);
nand U11026 (N_11026,N_10255,N_9816);
or U11027 (N_11027,N_10420,N_10123);
nor U11028 (N_11028,N_9816,N_10258);
xnor U11029 (N_11029,N_9890,N_9901);
or U11030 (N_11030,N_10191,N_10426);
or U11031 (N_11031,N_10221,N_10204);
nand U11032 (N_11032,N_10194,N_9855);
nand U11033 (N_11033,N_10495,N_10313);
or U11034 (N_11034,N_9762,N_9904);
or U11035 (N_11035,N_10202,N_9837);
nor U11036 (N_11036,N_10187,N_9965);
and U11037 (N_11037,N_10455,N_9756);
nand U11038 (N_11038,N_10341,N_10352);
or U11039 (N_11039,N_10285,N_10390);
nor U11040 (N_11040,N_9935,N_10484);
and U11041 (N_11041,N_9856,N_10131);
nand U11042 (N_11042,N_10252,N_9896);
and U11043 (N_11043,N_9819,N_10451);
xor U11044 (N_11044,N_10023,N_9931);
and U11045 (N_11045,N_10004,N_9833);
nor U11046 (N_11046,N_10097,N_10079);
nand U11047 (N_11047,N_10338,N_10389);
and U11048 (N_11048,N_10450,N_10483);
xor U11049 (N_11049,N_10077,N_10151);
or U11050 (N_11050,N_10236,N_9785);
nor U11051 (N_11051,N_10075,N_9958);
nor U11052 (N_11052,N_10194,N_10057);
and U11053 (N_11053,N_10197,N_9885);
nor U11054 (N_11054,N_10484,N_10055);
xnor U11055 (N_11055,N_10049,N_10346);
and U11056 (N_11056,N_10139,N_9911);
xnor U11057 (N_11057,N_10408,N_10372);
and U11058 (N_11058,N_9804,N_10452);
or U11059 (N_11059,N_9844,N_10333);
or U11060 (N_11060,N_10205,N_9899);
or U11061 (N_11061,N_10101,N_10153);
nor U11062 (N_11062,N_10246,N_9812);
and U11063 (N_11063,N_10107,N_9873);
and U11064 (N_11064,N_10445,N_10319);
nand U11065 (N_11065,N_10328,N_9992);
xnor U11066 (N_11066,N_10429,N_10190);
and U11067 (N_11067,N_9947,N_10169);
nor U11068 (N_11068,N_9800,N_10109);
nand U11069 (N_11069,N_10112,N_9888);
nand U11070 (N_11070,N_10278,N_9906);
or U11071 (N_11071,N_10264,N_9771);
nand U11072 (N_11072,N_9982,N_10304);
nor U11073 (N_11073,N_10126,N_10186);
and U11074 (N_11074,N_10087,N_10487);
xor U11075 (N_11075,N_9987,N_10214);
nand U11076 (N_11076,N_9893,N_10148);
or U11077 (N_11077,N_9848,N_10096);
nor U11078 (N_11078,N_10343,N_10181);
nor U11079 (N_11079,N_9878,N_10134);
nor U11080 (N_11080,N_10356,N_9765);
and U11081 (N_11081,N_10360,N_9834);
nand U11082 (N_11082,N_9802,N_10347);
or U11083 (N_11083,N_9961,N_10093);
nand U11084 (N_11084,N_10322,N_10137);
or U11085 (N_11085,N_10448,N_9883);
nor U11086 (N_11086,N_10082,N_9855);
or U11087 (N_11087,N_10449,N_10408);
nand U11088 (N_11088,N_10332,N_10052);
nor U11089 (N_11089,N_10490,N_10330);
nor U11090 (N_11090,N_9909,N_9977);
xor U11091 (N_11091,N_10418,N_9862);
and U11092 (N_11092,N_10390,N_9783);
or U11093 (N_11093,N_9983,N_10463);
xor U11094 (N_11094,N_10216,N_10290);
and U11095 (N_11095,N_10145,N_10004);
nor U11096 (N_11096,N_10434,N_9775);
xor U11097 (N_11097,N_10277,N_10255);
or U11098 (N_11098,N_9956,N_10206);
and U11099 (N_11099,N_10396,N_9998);
xnor U11100 (N_11100,N_10239,N_10408);
nand U11101 (N_11101,N_10384,N_10314);
or U11102 (N_11102,N_10413,N_10154);
nand U11103 (N_11103,N_10034,N_10186);
nand U11104 (N_11104,N_9810,N_9853);
nor U11105 (N_11105,N_9820,N_9830);
and U11106 (N_11106,N_10416,N_10300);
nor U11107 (N_11107,N_10390,N_10244);
xor U11108 (N_11108,N_10067,N_10149);
xor U11109 (N_11109,N_10340,N_10155);
nand U11110 (N_11110,N_10148,N_9971);
nor U11111 (N_11111,N_10007,N_9985);
or U11112 (N_11112,N_10102,N_10061);
nor U11113 (N_11113,N_10476,N_9912);
xor U11114 (N_11114,N_10070,N_10473);
and U11115 (N_11115,N_9775,N_10040);
and U11116 (N_11116,N_10195,N_9832);
and U11117 (N_11117,N_10462,N_9946);
nor U11118 (N_11118,N_9822,N_9996);
xor U11119 (N_11119,N_9813,N_10221);
and U11120 (N_11120,N_10019,N_10434);
xnor U11121 (N_11121,N_10099,N_10469);
and U11122 (N_11122,N_10234,N_10380);
nand U11123 (N_11123,N_10456,N_10220);
or U11124 (N_11124,N_10133,N_10177);
nor U11125 (N_11125,N_10196,N_10182);
nor U11126 (N_11126,N_10294,N_10387);
nor U11127 (N_11127,N_10340,N_9775);
nor U11128 (N_11128,N_9892,N_10189);
nand U11129 (N_11129,N_9981,N_10164);
and U11130 (N_11130,N_9975,N_9967);
and U11131 (N_11131,N_10205,N_10273);
and U11132 (N_11132,N_10286,N_9988);
and U11133 (N_11133,N_9762,N_9792);
xnor U11134 (N_11134,N_10100,N_9964);
nor U11135 (N_11135,N_10010,N_10070);
xnor U11136 (N_11136,N_9835,N_9963);
or U11137 (N_11137,N_10143,N_9793);
nand U11138 (N_11138,N_10350,N_10303);
or U11139 (N_11139,N_9779,N_10453);
nor U11140 (N_11140,N_9986,N_9779);
and U11141 (N_11141,N_10372,N_10210);
or U11142 (N_11142,N_9775,N_10203);
and U11143 (N_11143,N_9979,N_10274);
xnor U11144 (N_11144,N_10433,N_10302);
nor U11145 (N_11145,N_10059,N_10384);
or U11146 (N_11146,N_10024,N_9753);
or U11147 (N_11147,N_10218,N_9948);
and U11148 (N_11148,N_10285,N_10025);
xor U11149 (N_11149,N_9952,N_10129);
nand U11150 (N_11150,N_9814,N_10468);
or U11151 (N_11151,N_10239,N_9938);
and U11152 (N_11152,N_10208,N_10128);
and U11153 (N_11153,N_10101,N_10066);
nor U11154 (N_11154,N_10242,N_10011);
nor U11155 (N_11155,N_10446,N_10424);
nor U11156 (N_11156,N_10098,N_10224);
xnor U11157 (N_11157,N_10364,N_10360);
and U11158 (N_11158,N_10327,N_9938);
nor U11159 (N_11159,N_9969,N_9953);
or U11160 (N_11160,N_10230,N_10433);
nand U11161 (N_11161,N_10164,N_9876);
nor U11162 (N_11162,N_10415,N_10126);
and U11163 (N_11163,N_10206,N_9960);
and U11164 (N_11164,N_10127,N_10367);
xnor U11165 (N_11165,N_9864,N_9879);
or U11166 (N_11166,N_9953,N_10002);
or U11167 (N_11167,N_10159,N_9948);
nand U11168 (N_11168,N_10456,N_10266);
or U11169 (N_11169,N_10116,N_10160);
xnor U11170 (N_11170,N_9752,N_10435);
nand U11171 (N_11171,N_10205,N_9946);
and U11172 (N_11172,N_10175,N_10496);
or U11173 (N_11173,N_9887,N_10396);
xor U11174 (N_11174,N_10324,N_10132);
and U11175 (N_11175,N_10036,N_10125);
xor U11176 (N_11176,N_9774,N_10448);
nand U11177 (N_11177,N_9834,N_10374);
or U11178 (N_11178,N_10329,N_10044);
nand U11179 (N_11179,N_10455,N_10445);
and U11180 (N_11180,N_9765,N_10395);
or U11181 (N_11181,N_9890,N_10325);
nand U11182 (N_11182,N_9932,N_9987);
nand U11183 (N_11183,N_9986,N_10299);
nand U11184 (N_11184,N_10267,N_10006);
nand U11185 (N_11185,N_9880,N_10060);
nor U11186 (N_11186,N_10327,N_9826);
nand U11187 (N_11187,N_10127,N_10499);
or U11188 (N_11188,N_9980,N_10166);
and U11189 (N_11189,N_10178,N_10061);
or U11190 (N_11190,N_10347,N_10276);
and U11191 (N_11191,N_9928,N_9802);
or U11192 (N_11192,N_10436,N_9780);
nand U11193 (N_11193,N_10409,N_9961);
and U11194 (N_11194,N_10011,N_10375);
or U11195 (N_11195,N_9756,N_10026);
or U11196 (N_11196,N_9767,N_10460);
or U11197 (N_11197,N_10436,N_10163);
xnor U11198 (N_11198,N_9906,N_10388);
nor U11199 (N_11199,N_9845,N_9932);
nor U11200 (N_11200,N_10355,N_10313);
nor U11201 (N_11201,N_10191,N_10000);
or U11202 (N_11202,N_10223,N_10284);
or U11203 (N_11203,N_10434,N_9824);
and U11204 (N_11204,N_9857,N_10049);
xor U11205 (N_11205,N_9890,N_9902);
and U11206 (N_11206,N_10019,N_10300);
nand U11207 (N_11207,N_10159,N_10263);
nor U11208 (N_11208,N_10366,N_10097);
or U11209 (N_11209,N_10154,N_9951);
nand U11210 (N_11210,N_10255,N_9881);
nand U11211 (N_11211,N_10135,N_10088);
nor U11212 (N_11212,N_10477,N_9762);
nor U11213 (N_11213,N_9891,N_10298);
xnor U11214 (N_11214,N_9949,N_10022);
nor U11215 (N_11215,N_10405,N_9870);
nand U11216 (N_11216,N_10032,N_9828);
nand U11217 (N_11217,N_10051,N_10387);
xnor U11218 (N_11218,N_10142,N_10167);
nor U11219 (N_11219,N_10035,N_10363);
or U11220 (N_11220,N_9779,N_9926);
and U11221 (N_11221,N_10474,N_10230);
nor U11222 (N_11222,N_10049,N_10247);
nor U11223 (N_11223,N_9827,N_10268);
nor U11224 (N_11224,N_10175,N_10026);
nand U11225 (N_11225,N_9772,N_9787);
and U11226 (N_11226,N_10371,N_9819);
nand U11227 (N_11227,N_9813,N_10230);
xnor U11228 (N_11228,N_10438,N_10124);
or U11229 (N_11229,N_10087,N_10350);
nand U11230 (N_11230,N_9998,N_10174);
nand U11231 (N_11231,N_10467,N_9947);
and U11232 (N_11232,N_10376,N_9903);
or U11233 (N_11233,N_10043,N_9913);
nor U11234 (N_11234,N_10236,N_9761);
and U11235 (N_11235,N_10421,N_10044);
nor U11236 (N_11236,N_10298,N_9878);
nor U11237 (N_11237,N_10353,N_10459);
xnor U11238 (N_11238,N_10040,N_10008);
xnor U11239 (N_11239,N_9878,N_9908);
or U11240 (N_11240,N_10045,N_9974);
nor U11241 (N_11241,N_9782,N_9830);
and U11242 (N_11242,N_10277,N_10156);
nor U11243 (N_11243,N_10184,N_10010);
nor U11244 (N_11244,N_9938,N_9901);
nand U11245 (N_11245,N_10194,N_10210);
or U11246 (N_11246,N_10026,N_9964);
nor U11247 (N_11247,N_10352,N_10405);
nor U11248 (N_11248,N_10451,N_10471);
or U11249 (N_11249,N_10118,N_10460);
or U11250 (N_11250,N_10537,N_10779);
nor U11251 (N_11251,N_10816,N_10514);
and U11252 (N_11252,N_11013,N_10679);
nor U11253 (N_11253,N_11208,N_11155);
xnor U11254 (N_11254,N_10631,N_11140);
xnor U11255 (N_11255,N_10682,N_11084);
nand U11256 (N_11256,N_10750,N_11211);
nand U11257 (N_11257,N_10529,N_10548);
or U11258 (N_11258,N_10600,N_10835);
or U11259 (N_11259,N_10871,N_11100);
or U11260 (N_11260,N_10730,N_10734);
nor U11261 (N_11261,N_10878,N_11225);
nor U11262 (N_11262,N_10795,N_11164);
nor U11263 (N_11263,N_11056,N_10638);
xor U11264 (N_11264,N_10508,N_10846);
or U11265 (N_11265,N_10655,N_10982);
xnor U11266 (N_11266,N_11103,N_10998);
or U11267 (N_11267,N_10891,N_10762);
nand U11268 (N_11268,N_10761,N_10554);
and U11269 (N_11269,N_10993,N_10789);
or U11270 (N_11270,N_11047,N_10593);
and U11271 (N_11271,N_11133,N_11132);
xor U11272 (N_11272,N_10768,N_10776);
nor U11273 (N_11273,N_10944,N_10851);
and U11274 (N_11274,N_10536,N_11038);
nor U11275 (N_11275,N_10524,N_11186);
and U11276 (N_11276,N_10943,N_10757);
nand U11277 (N_11277,N_10644,N_10756);
nand U11278 (N_11278,N_11070,N_10958);
or U11279 (N_11279,N_10510,N_10842);
or U11280 (N_11280,N_11147,N_11049);
and U11281 (N_11281,N_11030,N_10935);
and U11282 (N_11282,N_10528,N_10926);
nor U11283 (N_11283,N_10705,N_11096);
or U11284 (N_11284,N_11042,N_11152);
xor U11285 (N_11285,N_11019,N_11207);
nor U11286 (N_11286,N_11245,N_11205);
nor U11287 (N_11287,N_10879,N_11102);
xor U11288 (N_11288,N_10589,N_10966);
nor U11289 (N_11289,N_10830,N_10639);
nand U11290 (N_11290,N_10530,N_10526);
and U11291 (N_11291,N_10857,N_11117);
nor U11292 (N_11292,N_10573,N_11003);
xor U11293 (N_11293,N_11137,N_10659);
or U11294 (N_11294,N_10901,N_10582);
nor U11295 (N_11295,N_11144,N_11112);
nor U11296 (N_11296,N_10911,N_11203);
and U11297 (N_11297,N_11009,N_10781);
and U11298 (N_11298,N_10610,N_11165);
and U11299 (N_11299,N_11162,N_10736);
nand U11300 (N_11300,N_11005,N_10652);
nor U11301 (N_11301,N_10597,N_11215);
xor U11302 (N_11302,N_11166,N_10615);
or U11303 (N_11303,N_11174,N_11247);
xnor U11304 (N_11304,N_10803,N_10534);
nand U11305 (N_11305,N_10562,N_10905);
or U11306 (N_11306,N_10619,N_10825);
xor U11307 (N_11307,N_10604,N_10745);
xnor U11308 (N_11308,N_10625,N_11143);
nand U11309 (N_11309,N_10581,N_10856);
nor U11310 (N_11310,N_11039,N_11237);
nand U11311 (N_11311,N_10599,N_10695);
and U11312 (N_11312,N_10633,N_10792);
and U11313 (N_11313,N_11241,N_10650);
or U11314 (N_11314,N_11122,N_11190);
xnor U11315 (N_11315,N_11016,N_10778);
xnor U11316 (N_11316,N_11017,N_10668);
nand U11317 (N_11317,N_11057,N_10544);
xor U11318 (N_11318,N_10831,N_10986);
or U11319 (N_11319,N_11108,N_10811);
xnor U11320 (N_11320,N_11189,N_10643);
nand U11321 (N_11321,N_10653,N_10937);
nor U11322 (N_11322,N_11249,N_10721);
nor U11323 (N_11323,N_10671,N_10635);
nor U11324 (N_11324,N_11218,N_10620);
or U11325 (N_11325,N_10931,N_11236);
nand U11326 (N_11326,N_11136,N_11200);
and U11327 (N_11327,N_10664,N_10894);
xor U11328 (N_11328,N_10665,N_11101);
or U11329 (N_11329,N_10836,N_11078);
nand U11330 (N_11330,N_11120,N_10896);
xor U11331 (N_11331,N_10543,N_11075);
nand U11332 (N_11332,N_10838,N_10691);
nand U11333 (N_11333,N_10787,N_11223);
xnor U11334 (N_11334,N_11015,N_10661);
xnor U11335 (N_11335,N_10670,N_10719);
or U11336 (N_11336,N_11074,N_10833);
nor U11337 (N_11337,N_10511,N_10929);
xnor U11338 (N_11338,N_11014,N_10553);
nor U11339 (N_11339,N_10991,N_10922);
nand U11340 (N_11340,N_10626,N_11028);
nand U11341 (N_11341,N_10797,N_10907);
or U11342 (N_11342,N_11179,N_10961);
nor U11343 (N_11343,N_11068,N_10782);
and U11344 (N_11344,N_10595,N_10527);
nor U11345 (N_11345,N_11182,N_10977);
xnor U11346 (N_11346,N_11077,N_10748);
or U11347 (N_11347,N_11149,N_10662);
nand U11348 (N_11348,N_11163,N_10974);
and U11349 (N_11349,N_10747,N_10590);
nor U11350 (N_11350,N_10686,N_10868);
and U11351 (N_11351,N_10788,N_10746);
and U11352 (N_11352,N_10583,N_11002);
xnor U11353 (N_11353,N_10801,N_10802);
or U11354 (N_11354,N_10711,N_10568);
nor U11355 (N_11355,N_11181,N_10699);
or U11356 (N_11356,N_10873,N_10696);
nor U11357 (N_11357,N_10587,N_11107);
nand U11358 (N_11358,N_11011,N_10983);
xor U11359 (N_11359,N_11041,N_10975);
nand U11360 (N_11360,N_10909,N_10557);
nand U11361 (N_11361,N_10503,N_10718);
and U11362 (N_11362,N_11008,N_10767);
nor U11363 (N_11363,N_10965,N_10794);
nand U11364 (N_11364,N_11021,N_10790);
nor U11365 (N_11365,N_10641,N_10906);
or U11366 (N_11366,N_10743,N_10613);
or U11367 (N_11367,N_10507,N_10985);
or U11368 (N_11368,N_11206,N_10561);
xnor U11369 (N_11369,N_10737,N_10884);
and U11370 (N_11370,N_10576,N_10675);
xnor U11371 (N_11371,N_10855,N_10706);
or U11372 (N_11372,N_10899,N_10577);
or U11373 (N_11373,N_10988,N_10770);
nor U11374 (N_11374,N_10956,N_10708);
or U11375 (N_11375,N_10924,N_10948);
nor U11376 (N_11376,N_11201,N_10598);
nor U11377 (N_11377,N_11234,N_10775);
or U11378 (N_11378,N_11157,N_10952);
or U11379 (N_11379,N_10919,N_10550);
and U11380 (N_11380,N_10940,N_10783);
and U11381 (N_11381,N_10932,N_10877);
xnor U11382 (N_11382,N_10515,N_10996);
or U11383 (N_11383,N_10531,N_10785);
nor U11384 (N_11384,N_11048,N_11188);
nand U11385 (N_11385,N_11058,N_10826);
nor U11386 (N_11386,N_10841,N_11081);
nand U11387 (N_11387,N_11083,N_10869);
xnor U11388 (N_11388,N_10552,N_10588);
or U11389 (N_11389,N_10642,N_10513);
nor U11390 (N_11390,N_10602,N_11145);
xor U11391 (N_11391,N_10637,N_10569);
nor U11392 (N_11392,N_10607,N_10606);
nor U11393 (N_11393,N_10880,N_10547);
xnor U11394 (N_11394,N_10621,N_10798);
xor U11395 (N_11395,N_10640,N_10964);
nor U11396 (N_11396,N_11035,N_11171);
or U11397 (N_11397,N_10727,N_10847);
and U11398 (N_11398,N_11138,N_10815);
nand U11399 (N_11399,N_10731,N_10611);
xor U11400 (N_11400,N_11125,N_11060);
nor U11401 (N_11401,N_11046,N_10697);
or U11402 (N_11402,N_11061,N_10751);
nor U11403 (N_11403,N_11160,N_10729);
and U11404 (N_11404,N_10674,N_10654);
or U11405 (N_11405,N_11178,N_11045);
nand U11406 (N_11406,N_11097,N_11246);
or U11407 (N_11407,N_11092,N_10647);
nor U11408 (N_11408,N_11232,N_10912);
and U11409 (N_11409,N_11240,N_10567);
or U11410 (N_11410,N_10518,N_11220);
nor U11411 (N_11411,N_10834,N_10810);
and U11412 (N_11412,N_11183,N_10804);
and U11413 (N_11413,N_10564,N_10592);
nor U11414 (N_11414,N_11036,N_11071);
and U11415 (N_11415,N_10942,N_11131);
xor U11416 (N_11416,N_10915,N_10819);
nor U11417 (N_11417,N_10735,N_11216);
nand U11418 (N_11418,N_10954,N_10506);
or U11419 (N_11419,N_10990,N_11175);
and U11420 (N_11420,N_11053,N_11198);
nand U11421 (N_11421,N_10934,N_10591);
xnor U11422 (N_11422,N_10973,N_10728);
and U11423 (N_11423,N_10765,N_10571);
nor U11424 (N_11424,N_10663,N_10887);
nand U11425 (N_11425,N_10546,N_10755);
and U11426 (N_11426,N_10800,N_11033);
or U11427 (N_11427,N_10987,N_11034);
nor U11428 (N_11428,N_10533,N_10744);
or U11429 (N_11429,N_10519,N_11230);
nor U11430 (N_11430,N_10829,N_10549);
nor U11431 (N_11431,N_11177,N_10870);
and U11432 (N_11432,N_10839,N_10875);
nand U11433 (N_11433,N_10651,N_11135);
and U11434 (N_11434,N_10914,N_11202);
xor U11435 (N_11435,N_11024,N_11025);
and U11436 (N_11436,N_10694,N_10740);
and U11437 (N_11437,N_10951,N_10683);
nor U11438 (N_11438,N_10898,N_10558);
nor U11439 (N_11439,N_10722,N_10703);
nor U11440 (N_11440,N_10876,N_11228);
or U11441 (N_11441,N_10648,N_11079);
nand U11442 (N_11442,N_11080,N_10823);
nand U11443 (N_11443,N_11116,N_10525);
or U11444 (N_11444,N_10749,N_10888);
or U11445 (N_11445,N_10962,N_10886);
nor U11446 (N_11446,N_10786,N_11156);
and U11447 (N_11447,N_10676,N_10720);
nor U11448 (N_11448,N_10502,N_11055);
and U11449 (N_11449,N_11209,N_11187);
or U11450 (N_11450,N_11054,N_11065);
and U11451 (N_11451,N_10628,N_11172);
nor U11452 (N_11452,N_10849,N_11180);
nor U11453 (N_11453,N_10960,N_11159);
nor U11454 (N_11454,N_10704,N_10978);
and U11455 (N_11455,N_10805,N_11128);
xor U11456 (N_11456,N_10541,N_10759);
or U11457 (N_11457,N_10578,N_11212);
nor U11458 (N_11458,N_11020,N_11231);
and U11459 (N_11459,N_10936,N_10707);
xor U11460 (N_11460,N_10723,N_10684);
nand U11461 (N_11461,N_10585,N_11010);
nor U11462 (N_11462,N_10902,N_11006);
xor U11463 (N_11463,N_10716,N_10563);
nand U11464 (N_11464,N_11063,N_10555);
and U11465 (N_11465,N_11085,N_10596);
or U11466 (N_11466,N_11098,N_10520);
xor U11467 (N_11467,N_10672,N_11022);
nand U11468 (N_11468,N_10574,N_11153);
nand U11469 (N_11469,N_11073,N_10687);
and U11470 (N_11470,N_11104,N_10614);
nor U11471 (N_11471,N_10752,N_10840);
or U11472 (N_11472,N_10813,N_11219);
nor U11473 (N_11473,N_10881,N_10617);
nor U11474 (N_11474,N_11114,N_11026);
nor U11475 (N_11475,N_10997,N_10742);
nand U11476 (N_11476,N_10758,N_10680);
nand U11477 (N_11477,N_10714,N_10764);
nand U11478 (N_11478,N_10913,N_10636);
nand U11479 (N_11479,N_10538,N_10889);
and U11480 (N_11480,N_11027,N_10732);
xor U11481 (N_11481,N_10681,N_11062);
nand U11482 (N_11482,N_11233,N_11076);
and U11483 (N_11483,N_10853,N_10715);
xor U11484 (N_11484,N_11109,N_10709);
nand U11485 (N_11485,N_11093,N_11210);
and U11486 (N_11486,N_11023,N_10504);
and U11487 (N_11487,N_10817,N_10771);
and U11488 (N_11488,N_11118,N_11185);
and U11489 (N_11489,N_10698,N_10989);
or U11490 (N_11490,N_10918,N_11032);
xor U11491 (N_11491,N_11224,N_10540);
xor U11492 (N_11492,N_10843,N_10917);
or U11493 (N_11493,N_11069,N_11126);
nor U11494 (N_11494,N_11094,N_11227);
nand U11495 (N_11495,N_11151,N_11127);
nand U11496 (N_11496,N_10972,N_11168);
or U11497 (N_11497,N_10669,N_10949);
xor U11498 (N_11498,N_11139,N_10941);
and U11499 (N_11499,N_10678,N_10809);
or U11500 (N_11500,N_11242,N_11130);
nor U11501 (N_11501,N_11222,N_10814);
and U11502 (N_11502,N_10923,N_10624);
nor U11503 (N_11503,N_10575,N_11043);
xor U11504 (N_11504,N_11018,N_10505);
xor U11505 (N_11505,N_11052,N_10791);
or U11506 (N_11506,N_11088,N_10844);
nand U11507 (N_11507,N_10892,N_10710);
or U11508 (N_11508,N_10845,N_11197);
or U11509 (N_11509,N_10850,N_10947);
and U11510 (N_11510,N_10657,N_11244);
xnor U11511 (N_11511,N_10971,N_10897);
nor U11512 (N_11512,N_11192,N_10821);
nor U11513 (N_11513,N_10629,N_10772);
nor U11514 (N_11514,N_10632,N_10572);
nand U11515 (N_11515,N_11099,N_10793);
nor U11516 (N_11516,N_11167,N_10930);
nand U11517 (N_11517,N_11150,N_10612);
and U11518 (N_11518,N_10967,N_10559);
or U11519 (N_11519,N_11204,N_11115);
or U11520 (N_11520,N_10953,N_11106);
and U11521 (N_11521,N_10532,N_11148);
nand U11522 (N_11522,N_11044,N_10908);
nor U11523 (N_11523,N_11105,N_10760);
nor U11524 (N_11524,N_11217,N_10666);
or U11525 (N_11525,N_10827,N_10784);
or U11526 (N_11526,N_10777,N_10579);
xnor U11527 (N_11527,N_10565,N_11194);
nor U11528 (N_11528,N_11064,N_11141);
and U11529 (N_11529,N_10645,N_10904);
nand U11530 (N_11530,N_10713,N_10859);
xor U11531 (N_11531,N_10866,N_10566);
or U11532 (N_11532,N_10660,N_10594);
or U11533 (N_11533,N_10910,N_10808);
and U11534 (N_11534,N_10861,N_11191);
nor U11535 (N_11535,N_10959,N_10939);
xor U11536 (N_11536,N_11124,N_11243);
nor U11537 (N_11537,N_10501,N_10979);
and U11538 (N_11538,N_10616,N_10700);
nand U11539 (N_11539,N_10509,N_10516);
xor U11540 (N_11540,N_11170,N_10885);
nor U11541 (N_11541,N_10535,N_11195);
or U11542 (N_11542,N_10928,N_11111);
nor U11543 (N_11543,N_10521,N_10837);
or U11544 (N_11544,N_10824,N_10981);
nor U11545 (N_11545,N_10754,N_10539);
nor U11546 (N_11546,N_11091,N_10980);
xnor U11547 (N_11547,N_11196,N_10946);
and U11548 (N_11548,N_10848,N_10689);
and U11549 (N_11549,N_10916,N_11029);
and U11550 (N_11550,N_11066,N_10522);
or U11551 (N_11551,N_10938,N_11113);
or U11552 (N_11552,N_10864,N_10551);
nand U11553 (N_11553,N_11226,N_10560);
nand U11554 (N_11554,N_11040,N_10608);
xnor U11555 (N_11555,N_10634,N_10806);
or U11556 (N_11556,N_10500,N_10725);
xor U11557 (N_11557,N_10656,N_10933);
xor U11558 (N_11558,N_10970,N_10976);
xor U11559 (N_11559,N_10992,N_11004);
xor U11560 (N_11560,N_10601,N_11095);
nor U11561 (N_11561,N_11199,N_10584);
or U11562 (N_11562,N_11221,N_10984);
nand U11563 (N_11563,N_10556,N_11072);
nand U11564 (N_11564,N_10822,N_11007);
nand U11565 (N_11565,N_10812,N_10920);
nand U11566 (N_11566,N_10692,N_11051);
xnor U11567 (N_11567,N_10832,N_11213);
or U11568 (N_11568,N_11142,N_10753);
nand U11569 (N_11569,N_10605,N_11176);
nor U11570 (N_11570,N_10945,N_11000);
and U11571 (N_11571,N_10673,N_10733);
xnor U11572 (N_11572,N_11087,N_10724);
or U11573 (N_11573,N_10677,N_10603);
nand U11574 (N_11574,N_11067,N_10852);
nand U11575 (N_11575,N_10623,N_10622);
xnor U11576 (N_11576,N_10649,N_11119);
xor U11577 (N_11577,N_11193,N_11173);
xnor U11578 (N_11578,N_11012,N_11214);
nand U11579 (N_11579,N_10701,N_11146);
xor U11580 (N_11580,N_10890,N_10712);
or U11581 (N_11581,N_10872,N_10925);
xnor U11582 (N_11582,N_10658,N_10921);
nor U11583 (N_11583,N_10627,N_11134);
xor U11584 (N_11584,N_11184,N_10586);
nor U11585 (N_11585,N_10769,N_10667);
or U11586 (N_11586,N_10895,N_10865);
and U11587 (N_11587,N_10862,N_10517);
and U11588 (N_11588,N_10994,N_10854);
nor U11589 (N_11589,N_11082,N_10618);
nor U11590 (N_11590,N_10512,N_10799);
nor U11591 (N_11591,N_10726,N_11059);
xnor U11592 (N_11592,N_10867,N_10766);
nor U11593 (N_11593,N_10950,N_11248);
nor U11594 (N_11594,N_10763,N_10820);
xnor U11595 (N_11595,N_10999,N_11129);
or U11596 (N_11596,N_11086,N_10828);
or U11597 (N_11597,N_10690,N_10955);
or U11598 (N_11598,N_11229,N_10969);
and U11599 (N_11599,N_11089,N_10796);
or U11600 (N_11600,N_10882,N_11169);
nand U11601 (N_11601,N_11121,N_11158);
and U11602 (N_11602,N_10646,N_10883);
and U11603 (N_11603,N_11123,N_10860);
or U11604 (N_11604,N_10580,N_10702);
nand U11605 (N_11605,N_11161,N_11050);
and U11606 (N_11606,N_10739,N_11090);
nor U11607 (N_11607,N_11238,N_10780);
and U11608 (N_11608,N_10900,N_11031);
and U11609 (N_11609,N_10693,N_10963);
or U11610 (N_11610,N_11154,N_10863);
xnor U11611 (N_11611,N_10807,N_10927);
nor U11612 (N_11612,N_11235,N_10630);
nand U11613 (N_11613,N_11239,N_10874);
xor U11614 (N_11614,N_10858,N_11001);
or U11615 (N_11615,N_10818,N_10685);
nor U11616 (N_11616,N_11037,N_10523);
or U11617 (N_11617,N_10688,N_10957);
nor U11618 (N_11618,N_10968,N_10570);
xor U11619 (N_11619,N_11110,N_10773);
nand U11620 (N_11620,N_10545,N_10995);
nand U11621 (N_11621,N_10903,N_10893);
nand U11622 (N_11622,N_10609,N_10774);
and U11623 (N_11623,N_10741,N_10542);
and U11624 (N_11624,N_10717,N_10738);
or U11625 (N_11625,N_10748,N_10817);
or U11626 (N_11626,N_11089,N_10975);
xnor U11627 (N_11627,N_11221,N_10526);
nand U11628 (N_11628,N_10609,N_11111);
or U11629 (N_11629,N_10668,N_10623);
or U11630 (N_11630,N_11014,N_10805);
and U11631 (N_11631,N_10674,N_10613);
or U11632 (N_11632,N_11087,N_10635);
and U11633 (N_11633,N_10518,N_10787);
or U11634 (N_11634,N_11007,N_10820);
and U11635 (N_11635,N_11044,N_11205);
or U11636 (N_11636,N_11041,N_11089);
or U11637 (N_11637,N_10856,N_11226);
or U11638 (N_11638,N_11139,N_10891);
nor U11639 (N_11639,N_10770,N_10833);
nand U11640 (N_11640,N_11074,N_10692);
xnor U11641 (N_11641,N_10939,N_10781);
xnor U11642 (N_11642,N_11140,N_10551);
and U11643 (N_11643,N_11158,N_10570);
nor U11644 (N_11644,N_10863,N_10919);
nor U11645 (N_11645,N_11103,N_10991);
or U11646 (N_11646,N_10862,N_11216);
and U11647 (N_11647,N_10931,N_11232);
and U11648 (N_11648,N_10943,N_11249);
and U11649 (N_11649,N_11002,N_10651);
and U11650 (N_11650,N_10800,N_11101);
or U11651 (N_11651,N_10665,N_11188);
xnor U11652 (N_11652,N_11015,N_10666);
and U11653 (N_11653,N_10663,N_11040);
or U11654 (N_11654,N_10621,N_10727);
or U11655 (N_11655,N_11145,N_11123);
xor U11656 (N_11656,N_10761,N_10962);
nand U11657 (N_11657,N_11100,N_10761);
and U11658 (N_11658,N_10940,N_11042);
nand U11659 (N_11659,N_11249,N_11068);
and U11660 (N_11660,N_10951,N_10784);
or U11661 (N_11661,N_10843,N_11027);
nand U11662 (N_11662,N_10739,N_10998);
xor U11663 (N_11663,N_11127,N_10728);
or U11664 (N_11664,N_10648,N_11148);
nand U11665 (N_11665,N_10525,N_11227);
nor U11666 (N_11666,N_10833,N_10788);
xor U11667 (N_11667,N_10927,N_11115);
nor U11668 (N_11668,N_10503,N_10925);
nor U11669 (N_11669,N_10664,N_11219);
xnor U11670 (N_11670,N_11177,N_10687);
nand U11671 (N_11671,N_10634,N_10940);
nor U11672 (N_11672,N_10929,N_11023);
nor U11673 (N_11673,N_10851,N_10971);
xor U11674 (N_11674,N_10927,N_10515);
or U11675 (N_11675,N_11190,N_10627);
nor U11676 (N_11676,N_10511,N_10654);
nor U11677 (N_11677,N_10503,N_10767);
nor U11678 (N_11678,N_10560,N_10973);
nor U11679 (N_11679,N_10684,N_10847);
nand U11680 (N_11680,N_11144,N_10707);
or U11681 (N_11681,N_10517,N_10568);
nand U11682 (N_11682,N_10607,N_10910);
xor U11683 (N_11683,N_10917,N_10904);
or U11684 (N_11684,N_10642,N_11190);
xor U11685 (N_11685,N_10563,N_10944);
nand U11686 (N_11686,N_10793,N_10680);
and U11687 (N_11687,N_10712,N_10619);
nor U11688 (N_11688,N_10767,N_10527);
or U11689 (N_11689,N_11200,N_10673);
and U11690 (N_11690,N_10900,N_10752);
and U11691 (N_11691,N_10745,N_10939);
nand U11692 (N_11692,N_10956,N_11057);
and U11693 (N_11693,N_10639,N_10593);
and U11694 (N_11694,N_10804,N_10691);
or U11695 (N_11695,N_11024,N_10892);
xor U11696 (N_11696,N_10893,N_10995);
nand U11697 (N_11697,N_10988,N_11037);
xor U11698 (N_11698,N_10822,N_10925);
nor U11699 (N_11699,N_10974,N_11188);
or U11700 (N_11700,N_11120,N_11005);
and U11701 (N_11701,N_10955,N_11018);
and U11702 (N_11702,N_11094,N_10737);
xnor U11703 (N_11703,N_11168,N_10876);
or U11704 (N_11704,N_11176,N_10715);
xor U11705 (N_11705,N_11189,N_10712);
and U11706 (N_11706,N_10955,N_10566);
or U11707 (N_11707,N_11170,N_10514);
or U11708 (N_11708,N_11017,N_10536);
nor U11709 (N_11709,N_10817,N_10891);
xnor U11710 (N_11710,N_10514,N_11008);
nand U11711 (N_11711,N_10826,N_10915);
and U11712 (N_11712,N_10836,N_10975);
nor U11713 (N_11713,N_11082,N_11239);
and U11714 (N_11714,N_11248,N_10872);
or U11715 (N_11715,N_10513,N_10826);
or U11716 (N_11716,N_11185,N_10563);
nand U11717 (N_11717,N_10848,N_11229);
nand U11718 (N_11718,N_11157,N_11220);
nor U11719 (N_11719,N_10584,N_10996);
nand U11720 (N_11720,N_11157,N_10684);
xnor U11721 (N_11721,N_10567,N_11125);
or U11722 (N_11722,N_10882,N_10689);
and U11723 (N_11723,N_10579,N_10990);
xnor U11724 (N_11724,N_10826,N_10571);
xor U11725 (N_11725,N_11116,N_10744);
or U11726 (N_11726,N_10734,N_11136);
and U11727 (N_11727,N_10573,N_11111);
xnor U11728 (N_11728,N_10636,N_10533);
or U11729 (N_11729,N_10835,N_10730);
or U11730 (N_11730,N_10815,N_10627);
nand U11731 (N_11731,N_10564,N_10670);
nor U11732 (N_11732,N_10700,N_10702);
xnor U11733 (N_11733,N_10877,N_11123);
xnor U11734 (N_11734,N_10780,N_10685);
xor U11735 (N_11735,N_10513,N_11102);
nand U11736 (N_11736,N_11134,N_10800);
nor U11737 (N_11737,N_10909,N_10692);
or U11738 (N_11738,N_10918,N_10966);
xor U11739 (N_11739,N_11228,N_10551);
nor U11740 (N_11740,N_10724,N_11107);
and U11741 (N_11741,N_10670,N_11145);
xnor U11742 (N_11742,N_10605,N_10773);
and U11743 (N_11743,N_10549,N_11215);
or U11744 (N_11744,N_10525,N_10631);
xor U11745 (N_11745,N_11161,N_10756);
or U11746 (N_11746,N_11174,N_10901);
and U11747 (N_11747,N_10793,N_11243);
xnor U11748 (N_11748,N_10578,N_11113);
xnor U11749 (N_11749,N_11002,N_10500);
and U11750 (N_11750,N_11236,N_11243);
xnor U11751 (N_11751,N_10880,N_11098);
nor U11752 (N_11752,N_11170,N_11240);
and U11753 (N_11753,N_10999,N_10891);
nand U11754 (N_11754,N_10619,N_11247);
xor U11755 (N_11755,N_10644,N_10918);
and U11756 (N_11756,N_10776,N_10622);
and U11757 (N_11757,N_10831,N_11085);
xnor U11758 (N_11758,N_10820,N_10709);
nor U11759 (N_11759,N_11212,N_11241);
or U11760 (N_11760,N_11007,N_10601);
xnor U11761 (N_11761,N_10952,N_10946);
nand U11762 (N_11762,N_11066,N_11175);
xnor U11763 (N_11763,N_10624,N_10784);
nand U11764 (N_11764,N_10839,N_10929);
nand U11765 (N_11765,N_11067,N_10708);
or U11766 (N_11766,N_11124,N_11180);
or U11767 (N_11767,N_11230,N_10611);
or U11768 (N_11768,N_10723,N_11199);
or U11769 (N_11769,N_10802,N_10923);
nand U11770 (N_11770,N_10723,N_10976);
xor U11771 (N_11771,N_11229,N_10648);
or U11772 (N_11772,N_10811,N_10558);
nand U11773 (N_11773,N_10881,N_10654);
xor U11774 (N_11774,N_10567,N_11076);
nand U11775 (N_11775,N_10957,N_10983);
or U11776 (N_11776,N_11084,N_10887);
nand U11777 (N_11777,N_10877,N_11020);
nand U11778 (N_11778,N_10539,N_11058);
and U11779 (N_11779,N_10816,N_11074);
nand U11780 (N_11780,N_10924,N_10849);
xnor U11781 (N_11781,N_10625,N_10620);
nor U11782 (N_11782,N_10823,N_11150);
nand U11783 (N_11783,N_10640,N_10974);
nand U11784 (N_11784,N_10908,N_11010);
or U11785 (N_11785,N_10851,N_10763);
and U11786 (N_11786,N_10774,N_10980);
nand U11787 (N_11787,N_10554,N_10975);
and U11788 (N_11788,N_10939,N_10704);
and U11789 (N_11789,N_10983,N_10730);
nand U11790 (N_11790,N_10720,N_10651);
or U11791 (N_11791,N_10559,N_10925);
nand U11792 (N_11792,N_10855,N_10928);
xor U11793 (N_11793,N_10786,N_10751);
nand U11794 (N_11794,N_10870,N_11103);
xnor U11795 (N_11795,N_10524,N_10874);
nor U11796 (N_11796,N_11239,N_10771);
xor U11797 (N_11797,N_10600,N_11175);
xnor U11798 (N_11798,N_10708,N_10634);
nor U11799 (N_11799,N_10996,N_10563);
and U11800 (N_11800,N_11101,N_10534);
and U11801 (N_11801,N_11138,N_10604);
and U11802 (N_11802,N_10775,N_10619);
and U11803 (N_11803,N_11247,N_10677);
and U11804 (N_11804,N_10961,N_11152);
or U11805 (N_11805,N_10713,N_10921);
nand U11806 (N_11806,N_11204,N_10790);
xnor U11807 (N_11807,N_10633,N_11114);
nand U11808 (N_11808,N_11030,N_10553);
or U11809 (N_11809,N_10741,N_10636);
xor U11810 (N_11810,N_10906,N_11061);
and U11811 (N_11811,N_11145,N_10659);
nor U11812 (N_11812,N_11034,N_10670);
nand U11813 (N_11813,N_10892,N_11041);
and U11814 (N_11814,N_10898,N_11241);
or U11815 (N_11815,N_11124,N_10936);
or U11816 (N_11816,N_10798,N_10943);
or U11817 (N_11817,N_10895,N_10617);
nand U11818 (N_11818,N_10965,N_10795);
and U11819 (N_11819,N_11024,N_10693);
nand U11820 (N_11820,N_11044,N_10523);
nor U11821 (N_11821,N_11218,N_10513);
xor U11822 (N_11822,N_10733,N_10942);
nand U11823 (N_11823,N_11077,N_10927);
nand U11824 (N_11824,N_10856,N_10664);
and U11825 (N_11825,N_10996,N_10695);
and U11826 (N_11826,N_10920,N_10720);
xnor U11827 (N_11827,N_11206,N_10900);
xnor U11828 (N_11828,N_11122,N_10656);
or U11829 (N_11829,N_10757,N_10913);
and U11830 (N_11830,N_10580,N_10525);
nand U11831 (N_11831,N_10536,N_10735);
or U11832 (N_11832,N_10897,N_10856);
nand U11833 (N_11833,N_11131,N_11149);
or U11834 (N_11834,N_10660,N_11137);
nand U11835 (N_11835,N_11136,N_10872);
nand U11836 (N_11836,N_10704,N_10747);
nor U11837 (N_11837,N_10538,N_10933);
xnor U11838 (N_11838,N_10567,N_10746);
and U11839 (N_11839,N_10673,N_11221);
or U11840 (N_11840,N_10653,N_10743);
nand U11841 (N_11841,N_10973,N_10985);
or U11842 (N_11842,N_11082,N_10907);
and U11843 (N_11843,N_10648,N_10578);
or U11844 (N_11844,N_11214,N_10676);
xnor U11845 (N_11845,N_11094,N_10857);
nor U11846 (N_11846,N_11144,N_10847);
nor U11847 (N_11847,N_10602,N_11095);
nor U11848 (N_11848,N_10902,N_11197);
xnor U11849 (N_11849,N_11038,N_10907);
or U11850 (N_11850,N_10995,N_10972);
nand U11851 (N_11851,N_10720,N_11200);
nand U11852 (N_11852,N_10825,N_11191);
and U11853 (N_11853,N_10900,N_10947);
xor U11854 (N_11854,N_10911,N_11133);
nor U11855 (N_11855,N_11183,N_11081);
xnor U11856 (N_11856,N_11024,N_10970);
and U11857 (N_11857,N_11045,N_11176);
or U11858 (N_11858,N_11205,N_10834);
xor U11859 (N_11859,N_10533,N_10518);
nor U11860 (N_11860,N_11073,N_10875);
nand U11861 (N_11861,N_11071,N_11031);
nand U11862 (N_11862,N_10822,N_10923);
nand U11863 (N_11863,N_11032,N_11183);
nand U11864 (N_11864,N_11029,N_10669);
and U11865 (N_11865,N_10690,N_10871);
nand U11866 (N_11866,N_10626,N_11178);
or U11867 (N_11867,N_10810,N_10935);
nand U11868 (N_11868,N_11214,N_11117);
nand U11869 (N_11869,N_10669,N_10991);
xnor U11870 (N_11870,N_11006,N_10951);
and U11871 (N_11871,N_10818,N_10541);
nor U11872 (N_11872,N_10745,N_10557);
nand U11873 (N_11873,N_10871,N_10718);
nand U11874 (N_11874,N_11086,N_11036);
nor U11875 (N_11875,N_10524,N_11120);
or U11876 (N_11876,N_10947,N_10866);
nor U11877 (N_11877,N_11249,N_11085);
and U11878 (N_11878,N_10796,N_10738);
nor U11879 (N_11879,N_10583,N_10516);
and U11880 (N_11880,N_10844,N_11171);
and U11881 (N_11881,N_11066,N_10712);
nor U11882 (N_11882,N_11035,N_10806);
or U11883 (N_11883,N_10889,N_10848);
xnor U11884 (N_11884,N_11060,N_10982);
nor U11885 (N_11885,N_10762,N_10830);
nand U11886 (N_11886,N_10885,N_10665);
and U11887 (N_11887,N_10758,N_11023);
nand U11888 (N_11888,N_10731,N_10683);
nand U11889 (N_11889,N_11244,N_10734);
nand U11890 (N_11890,N_11013,N_11100);
nand U11891 (N_11891,N_10768,N_10767);
nor U11892 (N_11892,N_11180,N_10633);
nor U11893 (N_11893,N_11201,N_10837);
and U11894 (N_11894,N_11048,N_10555);
or U11895 (N_11895,N_10863,N_10948);
xor U11896 (N_11896,N_10813,N_11004);
and U11897 (N_11897,N_10955,N_11084);
xor U11898 (N_11898,N_11017,N_11021);
or U11899 (N_11899,N_10661,N_10919);
nor U11900 (N_11900,N_11130,N_10676);
or U11901 (N_11901,N_11077,N_11129);
nand U11902 (N_11902,N_10943,N_11159);
nand U11903 (N_11903,N_11242,N_10556);
nor U11904 (N_11904,N_10599,N_11137);
xnor U11905 (N_11905,N_11164,N_11249);
nand U11906 (N_11906,N_11062,N_10911);
nor U11907 (N_11907,N_10706,N_11030);
nand U11908 (N_11908,N_11125,N_10563);
nor U11909 (N_11909,N_10740,N_11023);
nor U11910 (N_11910,N_11189,N_10775);
or U11911 (N_11911,N_10596,N_11059);
nand U11912 (N_11912,N_10630,N_10878);
xnor U11913 (N_11913,N_10577,N_11020);
xor U11914 (N_11914,N_10975,N_10870);
nand U11915 (N_11915,N_10704,N_10636);
and U11916 (N_11916,N_10983,N_11008);
and U11917 (N_11917,N_10788,N_11016);
nor U11918 (N_11918,N_10659,N_10720);
xnor U11919 (N_11919,N_10796,N_10525);
nand U11920 (N_11920,N_10854,N_10762);
nor U11921 (N_11921,N_10749,N_10771);
and U11922 (N_11922,N_11155,N_10951);
xnor U11923 (N_11923,N_11182,N_10556);
or U11924 (N_11924,N_10919,N_10912);
xor U11925 (N_11925,N_10802,N_10880);
or U11926 (N_11926,N_10957,N_10541);
and U11927 (N_11927,N_10825,N_11035);
or U11928 (N_11928,N_10949,N_10634);
xnor U11929 (N_11929,N_10896,N_10668);
nor U11930 (N_11930,N_10929,N_10596);
or U11931 (N_11931,N_10630,N_10676);
and U11932 (N_11932,N_11139,N_10580);
xor U11933 (N_11933,N_10988,N_10735);
and U11934 (N_11934,N_11238,N_10688);
xor U11935 (N_11935,N_10679,N_10623);
xor U11936 (N_11936,N_10697,N_11208);
xnor U11937 (N_11937,N_10762,N_10886);
nand U11938 (N_11938,N_10756,N_11065);
nor U11939 (N_11939,N_11003,N_10583);
xor U11940 (N_11940,N_11202,N_10606);
nand U11941 (N_11941,N_10739,N_11187);
nand U11942 (N_11942,N_10597,N_10893);
nand U11943 (N_11943,N_11234,N_10716);
or U11944 (N_11944,N_11200,N_10683);
and U11945 (N_11945,N_10754,N_10674);
and U11946 (N_11946,N_10989,N_11054);
nor U11947 (N_11947,N_11224,N_10737);
or U11948 (N_11948,N_10665,N_11200);
xnor U11949 (N_11949,N_10992,N_11110);
nand U11950 (N_11950,N_10535,N_10588);
nand U11951 (N_11951,N_10898,N_10748);
or U11952 (N_11952,N_10967,N_10622);
nor U11953 (N_11953,N_10634,N_10611);
and U11954 (N_11954,N_10787,N_10635);
xnor U11955 (N_11955,N_10872,N_10504);
and U11956 (N_11956,N_10858,N_10562);
nor U11957 (N_11957,N_10984,N_10718);
or U11958 (N_11958,N_11164,N_10953);
xor U11959 (N_11959,N_10891,N_10924);
or U11960 (N_11960,N_10811,N_11043);
xnor U11961 (N_11961,N_11059,N_10826);
and U11962 (N_11962,N_10549,N_10823);
nor U11963 (N_11963,N_10938,N_11207);
nor U11964 (N_11964,N_10567,N_11067);
xor U11965 (N_11965,N_10716,N_10740);
xnor U11966 (N_11966,N_10851,N_10653);
xnor U11967 (N_11967,N_10930,N_11104);
or U11968 (N_11968,N_11123,N_10525);
nand U11969 (N_11969,N_10682,N_10500);
and U11970 (N_11970,N_11197,N_10683);
and U11971 (N_11971,N_10697,N_10691);
nor U11972 (N_11972,N_11089,N_10915);
xnor U11973 (N_11973,N_11216,N_11088);
nor U11974 (N_11974,N_10677,N_11006);
xnor U11975 (N_11975,N_10800,N_11215);
or U11976 (N_11976,N_10833,N_10823);
or U11977 (N_11977,N_10592,N_10993);
and U11978 (N_11978,N_11240,N_10558);
and U11979 (N_11979,N_11020,N_10754);
xnor U11980 (N_11980,N_10659,N_11030);
xor U11981 (N_11981,N_11008,N_11177);
nand U11982 (N_11982,N_10667,N_11122);
and U11983 (N_11983,N_11051,N_11168);
or U11984 (N_11984,N_11131,N_10596);
or U11985 (N_11985,N_10911,N_10756);
nand U11986 (N_11986,N_10798,N_10747);
or U11987 (N_11987,N_11204,N_11213);
and U11988 (N_11988,N_11199,N_10885);
or U11989 (N_11989,N_10765,N_10566);
nand U11990 (N_11990,N_11011,N_10812);
xnor U11991 (N_11991,N_10969,N_11076);
and U11992 (N_11992,N_10972,N_10585);
or U11993 (N_11993,N_11194,N_10548);
and U11994 (N_11994,N_10724,N_11156);
nor U11995 (N_11995,N_11203,N_10703);
nand U11996 (N_11996,N_10999,N_10585);
and U11997 (N_11997,N_10832,N_11134);
nand U11998 (N_11998,N_10609,N_10844);
xnor U11999 (N_11999,N_10639,N_11208);
xnor U12000 (N_12000,N_11323,N_11258);
nor U12001 (N_12001,N_11932,N_11480);
xor U12002 (N_12002,N_11803,N_11705);
or U12003 (N_12003,N_11368,N_11523);
nor U12004 (N_12004,N_11844,N_11808);
nand U12005 (N_12005,N_11863,N_11336);
nor U12006 (N_12006,N_11382,N_11913);
and U12007 (N_12007,N_11327,N_11373);
nor U12008 (N_12008,N_11536,N_11745);
and U12009 (N_12009,N_11305,N_11629);
or U12010 (N_12010,N_11527,N_11814);
xor U12011 (N_12011,N_11748,N_11701);
nor U12012 (N_12012,N_11810,N_11770);
xor U12013 (N_12013,N_11857,N_11849);
nand U12014 (N_12014,N_11537,N_11736);
and U12015 (N_12015,N_11321,N_11965);
xnor U12016 (N_12016,N_11641,N_11337);
and U12017 (N_12017,N_11504,N_11391);
nand U12018 (N_12018,N_11372,N_11667);
or U12019 (N_12019,N_11998,N_11474);
nand U12020 (N_12020,N_11503,N_11779);
nor U12021 (N_12021,N_11912,N_11395);
nand U12022 (N_12022,N_11466,N_11429);
nand U12023 (N_12023,N_11737,N_11587);
or U12024 (N_12024,N_11813,N_11573);
and U12025 (N_12025,N_11762,N_11680);
nor U12026 (N_12026,N_11432,N_11982);
nor U12027 (N_12027,N_11401,N_11659);
xnor U12028 (N_12028,N_11823,N_11377);
or U12029 (N_12029,N_11329,N_11684);
or U12030 (N_12030,N_11797,N_11665);
nor U12031 (N_12031,N_11826,N_11981);
and U12032 (N_12032,N_11679,N_11974);
nand U12033 (N_12033,N_11361,N_11984);
and U12034 (N_12034,N_11458,N_11456);
nor U12035 (N_12035,N_11549,N_11371);
xnor U12036 (N_12036,N_11742,N_11953);
or U12037 (N_12037,N_11709,N_11482);
or U12038 (N_12038,N_11552,N_11827);
or U12039 (N_12039,N_11695,N_11563);
and U12040 (N_12040,N_11443,N_11653);
and U12041 (N_12041,N_11557,N_11265);
nor U12042 (N_12042,N_11835,N_11686);
xnor U12043 (N_12043,N_11764,N_11402);
nand U12044 (N_12044,N_11362,N_11383);
and U12045 (N_12045,N_11817,N_11483);
xor U12046 (N_12046,N_11427,N_11714);
or U12047 (N_12047,N_11741,N_11809);
nand U12048 (N_12048,N_11546,N_11767);
nand U12049 (N_12049,N_11850,N_11479);
xnor U12050 (N_12050,N_11822,N_11528);
nand U12051 (N_12051,N_11880,N_11409);
xor U12052 (N_12052,N_11387,N_11284);
or U12053 (N_12053,N_11920,N_11936);
nand U12054 (N_12054,N_11304,N_11992);
xnor U12055 (N_12055,N_11398,N_11644);
and U12056 (N_12056,N_11423,N_11875);
or U12057 (N_12057,N_11971,N_11494);
or U12058 (N_12058,N_11800,N_11859);
nor U12059 (N_12059,N_11670,N_11340);
nor U12060 (N_12060,N_11935,N_11300);
and U12061 (N_12061,N_11869,N_11365);
xnor U12062 (N_12062,N_11961,N_11307);
and U12063 (N_12063,N_11472,N_11820);
nand U12064 (N_12064,N_11638,N_11554);
or U12065 (N_12065,N_11261,N_11375);
xor U12066 (N_12066,N_11440,N_11821);
and U12067 (N_12067,N_11862,N_11513);
nand U12068 (N_12068,N_11853,N_11671);
xor U12069 (N_12069,N_11654,N_11461);
or U12070 (N_12070,N_11757,N_11646);
and U12071 (N_12071,N_11811,N_11279);
and U12072 (N_12072,N_11778,N_11914);
nor U12073 (N_12073,N_11302,N_11297);
or U12074 (N_12074,N_11393,N_11635);
xnor U12075 (N_12075,N_11611,N_11343);
nor U12076 (N_12076,N_11866,N_11656);
xnor U12077 (N_12077,N_11595,N_11309);
nor U12078 (N_12078,N_11711,N_11367);
and U12079 (N_12079,N_11754,N_11454);
nand U12080 (N_12080,N_11785,N_11311);
or U12081 (N_12081,N_11521,N_11255);
xnor U12082 (N_12082,N_11379,N_11675);
or U12083 (N_12083,N_11975,N_11290);
xor U12084 (N_12084,N_11649,N_11418);
nor U12085 (N_12085,N_11389,N_11796);
and U12086 (N_12086,N_11586,N_11958);
and U12087 (N_12087,N_11723,N_11506);
and U12088 (N_12088,N_11435,N_11882);
nor U12089 (N_12089,N_11699,N_11366);
or U12090 (N_12090,N_11792,N_11353);
and U12091 (N_12091,N_11783,N_11488);
nor U12092 (N_12092,N_11970,N_11782);
xnor U12093 (N_12093,N_11918,N_11788);
xnor U12094 (N_12094,N_11385,N_11747);
nor U12095 (N_12095,N_11446,N_11415);
nor U12096 (N_12096,N_11816,N_11344);
or U12097 (N_12097,N_11658,N_11606);
nand U12098 (N_12098,N_11685,N_11678);
and U12099 (N_12099,N_11356,N_11316);
and U12100 (N_12100,N_11358,N_11845);
nand U12101 (N_12101,N_11901,N_11477);
nor U12102 (N_12102,N_11760,N_11565);
and U12103 (N_12103,N_11614,N_11569);
or U12104 (N_12104,N_11713,N_11990);
or U12105 (N_12105,N_11887,N_11275);
xnor U12106 (N_12106,N_11496,N_11765);
or U12107 (N_12107,N_11396,N_11904);
or U12108 (N_12108,N_11906,N_11433);
and U12109 (N_12109,N_11553,N_11514);
xor U12110 (N_12110,N_11610,N_11408);
and U12111 (N_12111,N_11335,N_11497);
or U12112 (N_12112,N_11453,N_11956);
xnor U12113 (N_12113,N_11399,N_11286);
or U12114 (N_12114,N_11436,N_11855);
xnor U12115 (N_12115,N_11802,N_11299);
nand U12116 (N_12116,N_11681,N_11314);
nand U12117 (N_12117,N_11459,N_11331);
or U12118 (N_12118,N_11651,N_11350);
and U12119 (N_12119,N_11473,N_11541);
or U12120 (N_12120,N_11605,N_11627);
or U12121 (N_12121,N_11643,N_11942);
and U12122 (N_12122,N_11596,N_11465);
xor U12123 (N_12123,N_11831,N_11621);
and U12124 (N_12124,N_11292,N_11842);
nor U12125 (N_12125,N_11438,N_11317);
nand U12126 (N_12126,N_11938,N_11493);
or U12127 (N_12127,N_11896,N_11425);
nand U12128 (N_12128,N_11355,N_11381);
nand U12129 (N_12129,N_11420,N_11652);
nand U12130 (N_12130,N_11897,N_11457);
nor U12131 (N_12131,N_11374,N_11444);
and U12132 (N_12132,N_11698,N_11588);
or U12133 (N_12133,N_11294,N_11403);
and U12134 (N_12134,N_11895,N_11445);
or U12135 (N_12135,N_11417,N_11999);
xnor U12136 (N_12136,N_11848,N_11660);
and U12137 (N_12137,N_11922,N_11577);
nand U12138 (N_12138,N_11806,N_11475);
and U12139 (N_12139,N_11828,N_11648);
or U12140 (N_12140,N_11793,N_11930);
nor U12141 (N_12141,N_11568,N_11966);
nand U12142 (N_12142,N_11532,N_11950);
xnor U12143 (N_12143,N_11907,N_11538);
nand U12144 (N_12144,N_11271,N_11666);
nand U12145 (N_12145,N_11771,N_11562);
and U12146 (N_12146,N_11941,N_11676);
and U12147 (N_12147,N_11609,N_11949);
or U12148 (N_12148,N_11738,N_11910);
or U12149 (N_12149,N_11430,N_11750);
xor U12150 (N_12150,N_11500,N_11392);
and U12151 (N_12151,N_11283,N_11661);
xnor U12152 (N_12152,N_11636,N_11566);
nand U12153 (N_12153,N_11925,N_11468);
and U12154 (N_12154,N_11945,N_11341);
nor U12155 (N_12155,N_11968,N_11702);
and U12156 (N_12156,N_11773,N_11751);
nand U12157 (N_12157,N_11268,N_11753);
xnor U12158 (N_12158,N_11871,N_11662);
and U12159 (N_12159,N_11919,N_11404);
and U12160 (N_12160,N_11623,N_11732);
and U12161 (N_12161,N_11967,N_11634);
xor U12162 (N_12162,N_11406,N_11986);
xor U12163 (N_12163,N_11510,N_11301);
and U12164 (N_12164,N_11916,N_11450);
xor U12165 (N_12165,N_11664,N_11567);
or U12166 (N_12166,N_11893,N_11775);
or U12167 (N_12167,N_11560,N_11891);
nand U12168 (N_12168,N_11583,N_11884);
nor U12169 (N_12169,N_11630,N_11960);
xor U12170 (N_12170,N_11766,N_11346);
nand U12171 (N_12171,N_11861,N_11318);
nand U12172 (N_12172,N_11807,N_11498);
and U12173 (N_12173,N_11668,N_11278);
xor U12174 (N_12174,N_11428,N_11674);
nor U12175 (N_12175,N_11511,N_11692);
nand U12176 (N_12176,N_11997,N_11501);
xor U12177 (N_12177,N_11939,N_11281);
nor U12178 (N_12178,N_11755,N_11943);
or U12179 (N_12179,N_11288,N_11424);
xnor U12180 (N_12180,N_11703,N_11449);
xor U12181 (N_12181,N_11535,N_11502);
or U12182 (N_12182,N_11551,N_11499);
or U12183 (N_12183,N_11599,N_11731);
and U12184 (N_12184,N_11548,N_11915);
nand U12185 (N_12185,N_11865,N_11619);
and U12186 (N_12186,N_11710,N_11704);
nand U12187 (N_12187,N_11856,N_11386);
nand U12188 (N_12188,N_11898,N_11786);
and U12189 (N_12189,N_11780,N_11957);
nor U12190 (N_12190,N_11825,N_11364);
nand U12191 (N_12191,N_11917,N_11412);
and U12192 (N_12192,N_11378,N_11927);
nand U12193 (N_12193,N_11273,N_11544);
nor U12194 (N_12194,N_11252,N_11830);
nand U12195 (N_12195,N_11534,N_11794);
and U12196 (N_12196,N_11717,N_11892);
or U12197 (N_12197,N_11376,N_11791);
nand U12198 (N_12198,N_11603,N_11860);
nor U12199 (N_12199,N_11929,N_11540);
or U12200 (N_12200,N_11285,N_11463);
or U12201 (N_12201,N_11733,N_11706);
xnor U12202 (N_12202,N_11481,N_11334);
and U12203 (N_12203,N_11324,N_11602);
nand U12204 (N_12204,N_11962,N_11905);
nor U12205 (N_12205,N_11784,N_11987);
and U12206 (N_12206,N_11952,N_11909);
nor U12207 (N_12207,N_11526,N_11642);
xnor U12208 (N_12208,N_11618,N_11476);
and U12209 (N_12209,N_11947,N_11734);
nor U12210 (N_12210,N_11405,N_11508);
xnor U12211 (N_12211,N_11868,N_11263);
xor U12212 (N_12212,N_11448,N_11416);
nor U12213 (N_12213,N_11533,N_11253);
and U12214 (N_12214,N_11854,N_11798);
nand U12215 (N_12215,N_11529,N_11359);
xnor U12216 (N_12216,N_11616,N_11647);
or U12217 (N_12217,N_11840,N_11715);
xor U12218 (N_12218,N_11325,N_11490);
nand U12219 (N_12219,N_11617,N_11951);
nand U12220 (N_12220,N_11312,N_11873);
nor U12221 (N_12221,N_11581,N_11274);
xnor U12222 (N_12222,N_11296,N_11759);
xnor U12223 (N_12223,N_11597,N_11883);
nand U12224 (N_12224,N_11574,N_11524);
and U12225 (N_12225,N_11894,N_11491);
or U12226 (N_12226,N_11633,N_11819);
nor U12227 (N_12227,N_11315,N_11555);
nand U12228 (N_12228,N_11460,N_11697);
or U12229 (N_12229,N_11937,N_11721);
and U12230 (N_12230,N_11600,N_11262);
nand U12231 (N_12231,N_11872,N_11495);
nor U12232 (N_12232,N_11579,N_11888);
nor U12233 (N_12233,N_11516,N_11801);
or U12234 (N_12234,N_11545,N_11347);
and U12235 (N_12235,N_11972,N_11696);
and U12236 (N_12236,N_11351,N_11812);
xnor U12237 (N_12237,N_11934,N_11266);
nand U12238 (N_12238,N_11257,N_11303);
nor U12239 (N_12239,N_11963,N_11471);
xor U12240 (N_12240,N_11357,N_11923);
nor U12241 (N_12241,N_11889,N_11615);
nor U12242 (N_12242,N_11608,N_11580);
and U12243 (N_12243,N_11576,N_11272);
nand U12244 (N_12244,N_11735,N_11763);
or U12245 (N_12245,N_11774,N_11585);
and U12246 (N_12246,N_11756,N_11640);
nand U12247 (N_12247,N_11726,N_11991);
or U12248 (N_12248,N_11470,N_11989);
nor U12249 (N_12249,N_11776,N_11598);
xor U12250 (N_12250,N_11354,N_11531);
or U12251 (N_12251,N_11622,N_11486);
nor U12252 (N_12252,N_11712,N_11276);
nor U12253 (N_12253,N_11464,N_11570);
or U12254 (N_12254,N_11690,N_11841);
xnor U12255 (N_12255,N_11694,N_11795);
nor U12256 (N_12256,N_11940,N_11442);
or U12257 (N_12257,N_11988,N_11632);
and U12258 (N_12258,N_11979,N_11421);
or U12259 (N_12259,N_11289,N_11881);
nor U12260 (N_12260,N_11899,N_11250);
xor U12261 (N_12261,N_11769,N_11677);
or U12262 (N_12262,N_11522,N_11559);
nand U12263 (N_12263,N_11264,N_11360);
or U12264 (N_12264,N_11964,N_11969);
and U12265 (N_12265,N_11384,N_11693);
xnor U12266 (N_12266,N_11411,N_11295);
xnor U12267 (N_12267,N_11320,N_11267);
or U12268 (N_12268,N_11650,N_11837);
nand U12269 (N_12269,N_11370,N_11847);
nand U12270 (N_12270,N_11900,N_11328);
nor U12271 (N_12271,N_11903,N_11380);
or U12272 (N_12272,N_11270,N_11319);
nand U12273 (N_12273,N_11864,N_11489);
xnor U12274 (N_12274,N_11928,N_11781);
xnor U12275 (N_12275,N_11743,N_11310);
or U12276 (N_12276,N_11832,N_11575);
xor U12277 (N_12277,N_11836,N_11985);
xor U12278 (N_12278,N_11948,N_11592);
and U12279 (N_12279,N_11422,N_11749);
xor U12280 (N_12280,N_11407,N_11876);
xnor U12281 (N_12281,N_11911,N_11571);
or U12282 (N_12282,N_11682,N_11607);
nand U12283 (N_12283,N_11363,N_11419);
or U12284 (N_12284,N_11879,N_11455);
nor U12285 (N_12285,N_11451,N_11724);
nor U12286 (N_12286,N_11672,N_11761);
and U12287 (N_12287,N_11515,N_11637);
or U12288 (N_12288,N_11687,N_11447);
xnor U12289 (N_12289,N_11833,N_11700);
and U12290 (N_12290,N_11890,N_11768);
nand U12291 (N_12291,N_11517,N_11519);
nand U12292 (N_12292,N_11729,N_11254);
nor U12293 (N_12293,N_11777,N_11342);
nor U12294 (N_12294,N_11558,N_11469);
and U12295 (N_12295,N_11613,N_11744);
nand U12296 (N_12296,N_11485,N_11931);
nor U12297 (N_12297,N_11716,N_11867);
nor U12298 (N_12298,N_11954,N_11369);
and U12299 (N_12299,N_11955,N_11878);
nand U12300 (N_12300,N_11484,N_11708);
nand U12301 (N_12301,N_11413,N_11400);
nand U12302 (N_12302,N_11722,N_11345);
or U12303 (N_12303,N_11707,N_11604);
xor U12304 (N_12304,N_11787,N_11338);
and U12305 (N_12305,N_11397,N_11348);
xor U12306 (N_12306,N_11944,N_11730);
nor U12307 (N_12307,N_11655,N_11505);
xnor U12308 (N_12308,N_11790,N_11556);
or U12309 (N_12309,N_11691,N_11886);
nand U12310 (N_12310,N_11333,N_11752);
or U12311 (N_12311,N_11933,N_11799);
xor U12312 (N_12312,N_11349,N_11322);
nor U12313 (N_12313,N_11902,N_11657);
nand U12314 (N_12314,N_11829,N_11631);
nor U12315 (N_12315,N_11584,N_11530);
or U12316 (N_12316,N_11725,N_11578);
nand U12317 (N_12317,N_11256,N_11959);
and U12318 (N_12318,N_11547,N_11539);
or U12319 (N_12319,N_11824,N_11414);
or U12320 (N_12320,N_11946,N_11926);
nand U12321 (N_12321,N_11572,N_11280);
nor U12322 (N_12322,N_11976,N_11260);
and U12323 (N_12323,N_11620,N_11719);
and U12324 (N_12324,N_11720,N_11628);
nand U12325 (N_12325,N_11426,N_11512);
nand U12326 (N_12326,N_11439,N_11805);
nand U12327 (N_12327,N_11478,N_11851);
or U12328 (N_12328,N_11282,N_11924);
xor U12329 (N_12329,N_11983,N_11308);
nor U12330 (N_12330,N_11591,N_11718);
and U12331 (N_12331,N_11739,N_11452);
and U12332 (N_12332,N_11689,N_11789);
nor U12333 (N_12333,N_11838,N_11277);
nand U12334 (N_12334,N_11441,N_11639);
nor U12335 (N_12335,N_11434,N_11727);
nor U12336 (N_12336,N_11688,N_11994);
or U12337 (N_12337,N_11728,N_11673);
and U12338 (N_12338,N_11259,N_11908);
nor U12339 (N_12339,N_11542,N_11870);
and U12340 (N_12340,N_11846,N_11564);
nand U12341 (N_12341,N_11758,N_11525);
nand U12342 (N_12342,N_11394,N_11978);
nor U12343 (N_12343,N_11293,N_11996);
or U12344 (N_12344,N_11973,N_11582);
nor U12345 (N_12345,N_11645,N_11507);
and U12346 (N_12346,N_11431,N_11269);
xor U12347 (N_12347,N_11518,N_11462);
and U12348 (N_12348,N_11818,N_11326);
and U12349 (N_12349,N_11993,N_11625);
nor U12350 (N_12350,N_11663,N_11746);
or U12351 (N_12351,N_11388,N_11858);
and U12352 (N_12352,N_11980,N_11291);
or U12353 (N_12353,N_11287,N_11492);
nand U12354 (N_12354,N_11339,N_11885);
nand U12355 (N_12355,N_11487,N_11330);
and U12356 (N_12356,N_11669,N_11815);
nand U12357 (N_12357,N_11977,N_11594);
nor U12358 (N_12358,N_11740,N_11589);
and U12359 (N_12359,N_11352,N_11520);
nand U12360 (N_12360,N_11306,N_11839);
or U12361 (N_12361,N_11590,N_11772);
and U12362 (N_12362,N_11509,N_11626);
xnor U12363 (N_12363,N_11877,N_11410);
and U12364 (N_12364,N_11804,N_11390);
or U12365 (N_12365,N_11843,N_11298);
xor U12366 (N_12366,N_11624,N_11874);
and U12367 (N_12367,N_11467,N_11251);
nand U12368 (N_12368,N_11995,N_11313);
nand U12369 (N_12369,N_11601,N_11921);
nor U12370 (N_12370,N_11612,N_11543);
or U12371 (N_12371,N_11332,N_11437);
and U12372 (N_12372,N_11561,N_11550);
and U12373 (N_12373,N_11683,N_11593);
xnor U12374 (N_12374,N_11834,N_11852);
nand U12375 (N_12375,N_11763,N_11836);
xor U12376 (N_12376,N_11974,N_11968);
nor U12377 (N_12377,N_11469,N_11435);
xor U12378 (N_12378,N_11954,N_11807);
or U12379 (N_12379,N_11801,N_11951);
or U12380 (N_12380,N_11565,N_11839);
nand U12381 (N_12381,N_11875,N_11361);
nand U12382 (N_12382,N_11261,N_11380);
and U12383 (N_12383,N_11284,N_11625);
and U12384 (N_12384,N_11984,N_11833);
nand U12385 (N_12385,N_11906,N_11444);
nand U12386 (N_12386,N_11660,N_11680);
and U12387 (N_12387,N_11358,N_11686);
and U12388 (N_12388,N_11270,N_11800);
xor U12389 (N_12389,N_11809,N_11974);
xnor U12390 (N_12390,N_11438,N_11781);
nand U12391 (N_12391,N_11973,N_11967);
nor U12392 (N_12392,N_11278,N_11339);
xor U12393 (N_12393,N_11622,N_11497);
xnor U12394 (N_12394,N_11763,N_11407);
or U12395 (N_12395,N_11904,N_11666);
and U12396 (N_12396,N_11537,N_11823);
nor U12397 (N_12397,N_11377,N_11884);
or U12398 (N_12398,N_11552,N_11683);
xnor U12399 (N_12399,N_11342,N_11341);
nand U12400 (N_12400,N_11319,N_11874);
or U12401 (N_12401,N_11590,N_11297);
nand U12402 (N_12402,N_11554,N_11890);
or U12403 (N_12403,N_11690,N_11691);
and U12404 (N_12404,N_11662,N_11261);
nand U12405 (N_12405,N_11763,N_11527);
or U12406 (N_12406,N_11967,N_11490);
and U12407 (N_12407,N_11794,N_11543);
xnor U12408 (N_12408,N_11312,N_11926);
nand U12409 (N_12409,N_11774,N_11470);
xor U12410 (N_12410,N_11590,N_11400);
nor U12411 (N_12411,N_11617,N_11517);
and U12412 (N_12412,N_11349,N_11589);
xnor U12413 (N_12413,N_11307,N_11991);
and U12414 (N_12414,N_11316,N_11976);
nand U12415 (N_12415,N_11907,N_11656);
and U12416 (N_12416,N_11358,N_11768);
nand U12417 (N_12417,N_11649,N_11431);
nor U12418 (N_12418,N_11594,N_11889);
xor U12419 (N_12419,N_11931,N_11744);
nor U12420 (N_12420,N_11795,N_11673);
xor U12421 (N_12421,N_11367,N_11616);
and U12422 (N_12422,N_11702,N_11262);
nor U12423 (N_12423,N_11770,N_11321);
nor U12424 (N_12424,N_11444,N_11360);
or U12425 (N_12425,N_11397,N_11932);
nand U12426 (N_12426,N_11469,N_11899);
or U12427 (N_12427,N_11695,N_11662);
nand U12428 (N_12428,N_11309,N_11351);
nor U12429 (N_12429,N_11688,N_11262);
nor U12430 (N_12430,N_11619,N_11372);
nor U12431 (N_12431,N_11668,N_11583);
and U12432 (N_12432,N_11547,N_11585);
or U12433 (N_12433,N_11625,N_11692);
and U12434 (N_12434,N_11582,N_11616);
xor U12435 (N_12435,N_11509,N_11684);
nand U12436 (N_12436,N_11999,N_11542);
and U12437 (N_12437,N_11749,N_11419);
xnor U12438 (N_12438,N_11535,N_11762);
nand U12439 (N_12439,N_11293,N_11383);
or U12440 (N_12440,N_11884,N_11414);
xnor U12441 (N_12441,N_11350,N_11525);
nand U12442 (N_12442,N_11315,N_11289);
or U12443 (N_12443,N_11871,N_11663);
and U12444 (N_12444,N_11433,N_11647);
and U12445 (N_12445,N_11375,N_11407);
or U12446 (N_12446,N_11496,N_11746);
xnor U12447 (N_12447,N_11277,N_11938);
xnor U12448 (N_12448,N_11471,N_11789);
nor U12449 (N_12449,N_11830,N_11658);
and U12450 (N_12450,N_11578,N_11543);
nor U12451 (N_12451,N_11385,N_11906);
nor U12452 (N_12452,N_11522,N_11907);
and U12453 (N_12453,N_11589,N_11427);
or U12454 (N_12454,N_11788,N_11529);
or U12455 (N_12455,N_11514,N_11438);
nor U12456 (N_12456,N_11327,N_11786);
or U12457 (N_12457,N_11673,N_11444);
or U12458 (N_12458,N_11527,N_11910);
and U12459 (N_12459,N_11603,N_11729);
xor U12460 (N_12460,N_11859,N_11732);
xnor U12461 (N_12461,N_11631,N_11950);
or U12462 (N_12462,N_11731,N_11531);
or U12463 (N_12463,N_11544,N_11772);
nor U12464 (N_12464,N_11445,N_11673);
nor U12465 (N_12465,N_11283,N_11593);
nor U12466 (N_12466,N_11586,N_11785);
nand U12467 (N_12467,N_11916,N_11358);
nor U12468 (N_12468,N_11454,N_11946);
or U12469 (N_12469,N_11533,N_11815);
xnor U12470 (N_12470,N_11657,N_11385);
nand U12471 (N_12471,N_11979,N_11441);
or U12472 (N_12472,N_11393,N_11912);
xor U12473 (N_12473,N_11872,N_11832);
nand U12474 (N_12474,N_11879,N_11597);
and U12475 (N_12475,N_11262,N_11358);
or U12476 (N_12476,N_11589,N_11412);
nor U12477 (N_12477,N_11832,N_11270);
and U12478 (N_12478,N_11929,N_11385);
nor U12479 (N_12479,N_11667,N_11665);
xor U12480 (N_12480,N_11582,N_11490);
or U12481 (N_12481,N_11621,N_11594);
or U12482 (N_12482,N_11310,N_11727);
nor U12483 (N_12483,N_11250,N_11814);
nand U12484 (N_12484,N_11916,N_11477);
and U12485 (N_12485,N_11319,N_11385);
nand U12486 (N_12486,N_11782,N_11743);
and U12487 (N_12487,N_11882,N_11848);
nor U12488 (N_12488,N_11920,N_11900);
xor U12489 (N_12489,N_11288,N_11477);
and U12490 (N_12490,N_11345,N_11335);
nor U12491 (N_12491,N_11634,N_11934);
nor U12492 (N_12492,N_11890,N_11687);
xor U12493 (N_12493,N_11796,N_11441);
nand U12494 (N_12494,N_11729,N_11997);
and U12495 (N_12495,N_11670,N_11378);
or U12496 (N_12496,N_11839,N_11939);
nor U12497 (N_12497,N_11639,N_11529);
nor U12498 (N_12498,N_11637,N_11915);
nor U12499 (N_12499,N_11724,N_11398);
nand U12500 (N_12500,N_11364,N_11387);
and U12501 (N_12501,N_11554,N_11954);
nand U12502 (N_12502,N_11686,N_11544);
nor U12503 (N_12503,N_11441,N_11702);
and U12504 (N_12504,N_11725,N_11745);
nand U12505 (N_12505,N_11310,N_11583);
xnor U12506 (N_12506,N_11764,N_11477);
nor U12507 (N_12507,N_11356,N_11652);
nand U12508 (N_12508,N_11368,N_11623);
nand U12509 (N_12509,N_11423,N_11950);
or U12510 (N_12510,N_11823,N_11477);
nor U12511 (N_12511,N_11615,N_11938);
nor U12512 (N_12512,N_11565,N_11304);
nand U12513 (N_12513,N_11605,N_11989);
and U12514 (N_12514,N_11933,N_11930);
nor U12515 (N_12515,N_11722,N_11426);
or U12516 (N_12516,N_11682,N_11646);
and U12517 (N_12517,N_11278,N_11509);
and U12518 (N_12518,N_11277,N_11936);
nor U12519 (N_12519,N_11483,N_11708);
xnor U12520 (N_12520,N_11537,N_11425);
nand U12521 (N_12521,N_11293,N_11554);
xor U12522 (N_12522,N_11361,N_11961);
nand U12523 (N_12523,N_11871,N_11973);
xnor U12524 (N_12524,N_11729,N_11745);
nand U12525 (N_12525,N_11662,N_11828);
nor U12526 (N_12526,N_11907,N_11354);
or U12527 (N_12527,N_11566,N_11715);
or U12528 (N_12528,N_11769,N_11378);
or U12529 (N_12529,N_11935,N_11828);
or U12530 (N_12530,N_11952,N_11783);
xnor U12531 (N_12531,N_11496,N_11458);
nor U12532 (N_12532,N_11945,N_11895);
or U12533 (N_12533,N_11445,N_11392);
nand U12534 (N_12534,N_11955,N_11840);
and U12535 (N_12535,N_11936,N_11466);
nor U12536 (N_12536,N_11955,N_11995);
xnor U12537 (N_12537,N_11948,N_11949);
and U12538 (N_12538,N_11373,N_11887);
xor U12539 (N_12539,N_11556,N_11513);
nor U12540 (N_12540,N_11306,N_11599);
nor U12541 (N_12541,N_11579,N_11963);
xor U12542 (N_12542,N_11885,N_11769);
nor U12543 (N_12543,N_11662,N_11617);
xnor U12544 (N_12544,N_11266,N_11662);
nand U12545 (N_12545,N_11724,N_11519);
xnor U12546 (N_12546,N_11536,N_11942);
nor U12547 (N_12547,N_11658,N_11512);
nand U12548 (N_12548,N_11325,N_11601);
nand U12549 (N_12549,N_11555,N_11356);
nor U12550 (N_12550,N_11971,N_11304);
xnor U12551 (N_12551,N_11894,N_11587);
nand U12552 (N_12552,N_11255,N_11802);
and U12553 (N_12553,N_11603,N_11765);
nand U12554 (N_12554,N_11577,N_11951);
xor U12555 (N_12555,N_11509,N_11886);
nor U12556 (N_12556,N_11677,N_11628);
or U12557 (N_12557,N_11294,N_11535);
xnor U12558 (N_12558,N_11289,N_11297);
nor U12559 (N_12559,N_11687,N_11521);
xor U12560 (N_12560,N_11644,N_11737);
and U12561 (N_12561,N_11585,N_11387);
and U12562 (N_12562,N_11859,N_11337);
nor U12563 (N_12563,N_11851,N_11923);
nor U12564 (N_12564,N_11855,N_11492);
or U12565 (N_12565,N_11305,N_11412);
and U12566 (N_12566,N_11393,N_11990);
and U12567 (N_12567,N_11787,N_11348);
and U12568 (N_12568,N_11363,N_11394);
xor U12569 (N_12569,N_11411,N_11263);
xor U12570 (N_12570,N_11337,N_11253);
or U12571 (N_12571,N_11472,N_11325);
xor U12572 (N_12572,N_11385,N_11612);
xnor U12573 (N_12573,N_11600,N_11506);
and U12574 (N_12574,N_11620,N_11587);
and U12575 (N_12575,N_11709,N_11862);
xnor U12576 (N_12576,N_11470,N_11609);
xor U12577 (N_12577,N_11861,N_11612);
or U12578 (N_12578,N_11354,N_11494);
or U12579 (N_12579,N_11525,N_11589);
nand U12580 (N_12580,N_11647,N_11589);
and U12581 (N_12581,N_11849,N_11459);
nand U12582 (N_12582,N_11302,N_11495);
and U12583 (N_12583,N_11505,N_11557);
and U12584 (N_12584,N_11743,N_11990);
or U12585 (N_12585,N_11918,N_11925);
nand U12586 (N_12586,N_11786,N_11793);
or U12587 (N_12587,N_11865,N_11958);
nand U12588 (N_12588,N_11366,N_11473);
and U12589 (N_12589,N_11846,N_11642);
nand U12590 (N_12590,N_11528,N_11500);
nand U12591 (N_12591,N_11690,N_11810);
nor U12592 (N_12592,N_11966,N_11336);
xor U12593 (N_12593,N_11957,N_11755);
nor U12594 (N_12594,N_11330,N_11594);
nor U12595 (N_12595,N_11718,N_11826);
or U12596 (N_12596,N_11587,N_11705);
nand U12597 (N_12597,N_11749,N_11882);
xnor U12598 (N_12598,N_11924,N_11761);
or U12599 (N_12599,N_11666,N_11309);
and U12600 (N_12600,N_11978,N_11930);
nand U12601 (N_12601,N_11905,N_11256);
or U12602 (N_12602,N_11517,N_11507);
and U12603 (N_12603,N_11649,N_11458);
and U12604 (N_12604,N_11458,N_11348);
or U12605 (N_12605,N_11389,N_11655);
or U12606 (N_12606,N_11865,N_11327);
nand U12607 (N_12607,N_11269,N_11328);
nand U12608 (N_12608,N_11308,N_11751);
and U12609 (N_12609,N_11874,N_11574);
and U12610 (N_12610,N_11927,N_11769);
or U12611 (N_12611,N_11714,N_11389);
and U12612 (N_12612,N_11530,N_11917);
or U12613 (N_12613,N_11346,N_11417);
nand U12614 (N_12614,N_11975,N_11623);
and U12615 (N_12615,N_11545,N_11360);
or U12616 (N_12616,N_11318,N_11450);
xnor U12617 (N_12617,N_11760,N_11856);
or U12618 (N_12618,N_11865,N_11972);
nand U12619 (N_12619,N_11641,N_11406);
nand U12620 (N_12620,N_11675,N_11571);
and U12621 (N_12621,N_11322,N_11495);
and U12622 (N_12622,N_11863,N_11928);
or U12623 (N_12623,N_11669,N_11889);
xor U12624 (N_12624,N_11377,N_11389);
and U12625 (N_12625,N_11824,N_11566);
nor U12626 (N_12626,N_11806,N_11852);
or U12627 (N_12627,N_11504,N_11759);
xor U12628 (N_12628,N_11717,N_11646);
nand U12629 (N_12629,N_11970,N_11951);
or U12630 (N_12630,N_11895,N_11846);
nor U12631 (N_12631,N_11365,N_11265);
and U12632 (N_12632,N_11371,N_11788);
and U12633 (N_12633,N_11993,N_11936);
xnor U12634 (N_12634,N_11671,N_11532);
or U12635 (N_12635,N_11297,N_11632);
or U12636 (N_12636,N_11915,N_11413);
or U12637 (N_12637,N_11506,N_11517);
xnor U12638 (N_12638,N_11863,N_11415);
nor U12639 (N_12639,N_11404,N_11997);
and U12640 (N_12640,N_11848,N_11693);
or U12641 (N_12641,N_11990,N_11696);
xor U12642 (N_12642,N_11455,N_11775);
xnor U12643 (N_12643,N_11746,N_11478);
and U12644 (N_12644,N_11913,N_11553);
or U12645 (N_12645,N_11374,N_11893);
nand U12646 (N_12646,N_11923,N_11687);
xor U12647 (N_12647,N_11616,N_11397);
xnor U12648 (N_12648,N_11618,N_11852);
nand U12649 (N_12649,N_11686,N_11517);
xor U12650 (N_12650,N_11743,N_11512);
xnor U12651 (N_12651,N_11453,N_11534);
and U12652 (N_12652,N_11262,N_11562);
nand U12653 (N_12653,N_11992,N_11370);
xor U12654 (N_12654,N_11803,N_11860);
xor U12655 (N_12655,N_11923,N_11926);
xor U12656 (N_12656,N_11581,N_11525);
nand U12657 (N_12657,N_11982,N_11538);
xnor U12658 (N_12658,N_11478,N_11459);
nor U12659 (N_12659,N_11670,N_11919);
and U12660 (N_12660,N_11639,N_11635);
nand U12661 (N_12661,N_11250,N_11404);
and U12662 (N_12662,N_11560,N_11471);
nor U12663 (N_12663,N_11889,N_11679);
nand U12664 (N_12664,N_11372,N_11565);
nor U12665 (N_12665,N_11933,N_11985);
nand U12666 (N_12666,N_11900,N_11957);
or U12667 (N_12667,N_11609,N_11308);
or U12668 (N_12668,N_11519,N_11296);
and U12669 (N_12669,N_11781,N_11654);
nand U12670 (N_12670,N_11835,N_11634);
nand U12671 (N_12671,N_11766,N_11859);
nand U12672 (N_12672,N_11878,N_11267);
nand U12673 (N_12673,N_11360,N_11466);
nor U12674 (N_12674,N_11280,N_11916);
and U12675 (N_12675,N_11540,N_11270);
nand U12676 (N_12676,N_11632,N_11920);
nand U12677 (N_12677,N_11753,N_11504);
or U12678 (N_12678,N_11552,N_11285);
xor U12679 (N_12679,N_11555,N_11277);
nand U12680 (N_12680,N_11984,N_11878);
and U12681 (N_12681,N_11631,N_11780);
xnor U12682 (N_12682,N_11510,N_11967);
and U12683 (N_12683,N_11257,N_11734);
nand U12684 (N_12684,N_11349,N_11265);
nor U12685 (N_12685,N_11302,N_11393);
and U12686 (N_12686,N_11711,N_11991);
or U12687 (N_12687,N_11677,N_11624);
nand U12688 (N_12688,N_11680,N_11833);
or U12689 (N_12689,N_11299,N_11744);
nor U12690 (N_12690,N_11470,N_11416);
or U12691 (N_12691,N_11539,N_11477);
or U12692 (N_12692,N_11883,N_11254);
and U12693 (N_12693,N_11455,N_11304);
nor U12694 (N_12694,N_11784,N_11577);
xor U12695 (N_12695,N_11743,N_11783);
xnor U12696 (N_12696,N_11413,N_11395);
and U12697 (N_12697,N_11422,N_11556);
nor U12698 (N_12698,N_11389,N_11689);
or U12699 (N_12699,N_11548,N_11827);
and U12700 (N_12700,N_11697,N_11913);
or U12701 (N_12701,N_11438,N_11262);
and U12702 (N_12702,N_11763,N_11761);
nor U12703 (N_12703,N_11947,N_11483);
and U12704 (N_12704,N_11997,N_11936);
nand U12705 (N_12705,N_11781,N_11546);
or U12706 (N_12706,N_11617,N_11832);
nor U12707 (N_12707,N_11447,N_11357);
nand U12708 (N_12708,N_11842,N_11339);
and U12709 (N_12709,N_11964,N_11538);
and U12710 (N_12710,N_11877,N_11281);
xnor U12711 (N_12711,N_11260,N_11285);
nand U12712 (N_12712,N_11700,N_11593);
or U12713 (N_12713,N_11408,N_11329);
xor U12714 (N_12714,N_11895,N_11989);
or U12715 (N_12715,N_11570,N_11352);
nor U12716 (N_12716,N_11584,N_11311);
nor U12717 (N_12717,N_11675,N_11725);
nand U12718 (N_12718,N_11908,N_11759);
xnor U12719 (N_12719,N_11360,N_11935);
or U12720 (N_12720,N_11628,N_11638);
and U12721 (N_12721,N_11354,N_11550);
nand U12722 (N_12722,N_11318,N_11464);
nor U12723 (N_12723,N_11581,N_11932);
and U12724 (N_12724,N_11807,N_11294);
nand U12725 (N_12725,N_11984,N_11842);
or U12726 (N_12726,N_11840,N_11849);
nor U12727 (N_12727,N_11970,N_11325);
nor U12728 (N_12728,N_11807,N_11760);
and U12729 (N_12729,N_11455,N_11415);
xnor U12730 (N_12730,N_11691,N_11631);
and U12731 (N_12731,N_11805,N_11347);
xnor U12732 (N_12732,N_11803,N_11904);
and U12733 (N_12733,N_11265,N_11308);
nand U12734 (N_12734,N_11554,N_11778);
and U12735 (N_12735,N_11387,N_11306);
nand U12736 (N_12736,N_11719,N_11490);
or U12737 (N_12737,N_11463,N_11423);
xor U12738 (N_12738,N_11635,N_11687);
nor U12739 (N_12739,N_11419,N_11477);
xnor U12740 (N_12740,N_11378,N_11574);
and U12741 (N_12741,N_11633,N_11905);
and U12742 (N_12742,N_11899,N_11365);
xor U12743 (N_12743,N_11892,N_11697);
xnor U12744 (N_12744,N_11272,N_11493);
and U12745 (N_12745,N_11315,N_11936);
and U12746 (N_12746,N_11994,N_11897);
or U12747 (N_12747,N_11350,N_11699);
or U12748 (N_12748,N_11985,N_11298);
or U12749 (N_12749,N_11839,N_11570);
nor U12750 (N_12750,N_12743,N_12699);
nand U12751 (N_12751,N_12302,N_12073);
nand U12752 (N_12752,N_12039,N_12217);
and U12753 (N_12753,N_12234,N_12350);
nor U12754 (N_12754,N_12293,N_12229);
nand U12755 (N_12755,N_12109,N_12540);
nand U12756 (N_12756,N_12210,N_12047);
and U12757 (N_12757,N_12211,N_12006);
and U12758 (N_12758,N_12444,N_12209);
or U12759 (N_12759,N_12377,N_12333);
nor U12760 (N_12760,N_12405,N_12521);
xor U12761 (N_12761,N_12393,N_12711);
nor U12762 (N_12762,N_12583,N_12306);
nor U12763 (N_12763,N_12403,N_12335);
xnor U12764 (N_12764,N_12121,N_12471);
and U12765 (N_12765,N_12387,N_12218);
xnor U12766 (N_12766,N_12451,N_12247);
and U12767 (N_12767,N_12475,N_12362);
nor U12768 (N_12768,N_12119,N_12627);
xor U12769 (N_12769,N_12677,N_12465);
nand U12770 (N_12770,N_12093,N_12733);
nor U12771 (N_12771,N_12037,N_12505);
nor U12772 (N_12772,N_12597,N_12500);
and U12773 (N_12773,N_12022,N_12185);
nand U12774 (N_12774,N_12285,N_12042);
nor U12775 (N_12775,N_12352,N_12686);
nand U12776 (N_12776,N_12226,N_12263);
and U12777 (N_12777,N_12025,N_12246);
xnor U12778 (N_12778,N_12545,N_12590);
nand U12779 (N_12779,N_12360,N_12174);
nand U12780 (N_12780,N_12466,N_12469);
or U12781 (N_12781,N_12598,N_12072);
and U12782 (N_12782,N_12001,N_12323);
nor U12783 (N_12783,N_12150,N_12230);
or U12784 (N_12784,N_12573,N_12083);
xor U12785 (N_12785,N_12404,N_12544);
or U12786 (N_12786,N_12433,N_12515);
nand U12787 (N_12787,N_12248,N_12354);
xnor U12788 (N_12788,N_12558,N_12554);
xnor U12789 (N_12789,N_12443,N_12303);
or U12790 (N_12790,N_12024,N_12700);
xnor U12791 (N_12791,N_12696,N_12049);
xnor U12792 (N_12792,N_12084,N_12113);
and U12793 (N_12793,N_12068,N_12679);
or U12794 (N_12794,N_12088,N_12522);
nand U12795 (N_12795,N_12675,N_12565);
nand U12796 (N_12796,N_12551,N_12114);
nand U12797 (N_12797,N_12177,N_12528);
or U12798 (N_12798,N_12026,N_12144);
nand U12799 (N_12799,N_12625,N_12574);
nor U12800 (N_12800,N_12513,N_12474);
nand U12801 (N_12801,N_12007,N_12043);
and U12802 (N_12802,N_12529,N_12227);
xor U12803 (N_12803,N_12348,N_12734);
xor U12804 (N_12804,N_12407,N_12721);
nor U12805 (N_12805,N_12657,N_12607);
nand U12806 (N_12806,N_12301,N_12324);
and U12807 (N_12807,N_12608,N_12311);
and U12808 (N_12808,N_12029,N_12391);
xnor U12809 (N_12809,N_12682,N_12669);
and U12810 (N_12810,N_12347,N_12603);
nor U12811 (N_12811,N_12196,N_12138);
nand U12812 (N_12812,N_12532,N_12718);
nand U12813 (N_12813,N_12313,N_12535);
xnor U12814 (N_12814,N_12320,N_12673);
or U12815 (N_12815,N_12631,N_12260);
or U12816 (N_12816,N_12566,N_12117);
nor U12817 (N_12817,N_12648,N_12108);
nor U12818 (N_12818,N_12462,N_12291);
nor U12819 (N_12819,N_12413,N_12666);
or U12820 (N_12820,N_12330,N_12292);
and U12821 (N_12821,N_12056,N_12110);
xnor U12822 (N_12822,N_12103,N_12261);
nor U12823 (N_12823,N_12112,N_12204);
nor U12824 (N_12824,N_12099,N_12132);
nand U12825 (N_12825,N_12621,N_12325);
or U12826 (N_12826,N_12687,N_12271);
and U12827 (N_12827,N_12460,N_12123);
or U12828 (N_12828,N_12539,N_12432);
nor U12829 (N_12829,N_12438,N_12568);
and U12830 (N_12830,N_12251,N_12375);
and U12831 (N_12831,N_12312,N_12082);
nand U12832 (N_12832,N_12690,N_12710);
nand U12833 (N_12833,N_12168,N_12319);
xor U12834 (N_12834,N_12611,N_12105);
or U12835 (N_12835,N_12041,N_12388);
nor U12836 (N_12836,N_12592,N_12050);
xor U12837 (N_12837,N_12536,N_12698);
and U12838 (N_12838,N_12215,N_12078);
xnor U12839 (N_12839,N_12013,N_12664);
and U12840 (N_12840,N_12694,N_12149);
nor U12841 (N_12841,N_12200,N_12076);
and U12842 (N_12842,N_12672,N_12428);
xnor U12843 (N_12843,N_12142,N_12612);
or U12844 (N_12844,N_12137,N_12647);
xor U12845 (N_12845,N_12283,N_12418);
nor U12846 (N_12846,N_12747,N_12392);
nor U12847 (N_12847,N_12705,N_12649);
nand U12848 (N_12848,N_12178,N_12289);
xor U12849 (N_12849,N_12616,N_12715);
nor U12850 (N_12850,N_12118,N_12000);
xnor U12851 (N_12851,N_12512,N_12359);
nor U12852 (N_12852,N_12395,N_12693);
and U12853 (N_12853,N_12337,N_12183);
nor U12854 (N_12854,N_12031,N_12599);
or U12855 (N_12855,N_12345,N_12125);
and U12856 (N_12856,N_12156,N_12678);
nor U12857 (N_12857,N_12129,N_12635);
nand U12858 (N_12858,N_12508,N_12424);
nand U12859 (N_12859,N_12151,N_12143);
and U12860 (N_12860,N_12579,N_12652);
nand U12861 (N_12861,N_12446,N_12439);
or U12862 (N_12862,N_12070,N_12258);
nor U12863 (N_12863,N_12336,N_12563);
or U12864 (N_12864,N_12224,N_12268);
and U12865 (N_12865,N_12662,N_12382);
nor U12866 (N_12866,N_12610,N_12576);
or U12867 (N_12867,N_12706,N_12442);
nand U12868 (N_12868,N_12243,N_12427);
nor U12869 (N_12869,N_12018,N_12537);
and U12870 (N_12870,N_12282,N_12133);
xor U12871 (N_12871,N_12477,N_12735);
nand U12872 (N_12872,N_12380,N_12334);
nor U12873 (N_12873,N_12327,N_12638);
nand U12874 (N_12874,N_12180,N_12572);
or U12875 (N_12875,N_12300,N_12250);
xor U12876 (N_12876,N_12594,N_12437);
nand U12877 (N_12877,N_12371,N_12464);
or U12878 (N_12878,N_12501,N_12378);
nor U12879 (N_12879,N_12684,N_12159);
nor U12880 (N_12880,N_12434,N_12061);
and U12881 (N_12881,N_12090,N_12309);
and U12882 (N_12882,N_12569,N_12527);
nand U12883 (N_12883,N_12738,N_12317);
or U12884 (N_12884,N_12278,N_12096);
nand U12885 (N_12885,N_12517,N_12134);
nor U12886 (N_12886,N_12550,N_12379);
nor U12887 (N_12887,N_12152,N_12228);
or U12888 (N_12888,N_12267,N_12122);
nand U12889 (N_12889,N_12467,N_12028);
nor U12890 (N_12890,N_12717,N_12339);
or U12891 (N_12891,N_12255,N_12578);
nor U12892 (N_12892,N_12615,N_12280);
nand U12893 (N_12893,N_12493,N_12128);
xor U12894 (N_12894,N_12491,N_12340);
xnor U12895 (N_12895,N_12081,N_12441);
nand U12896 (N_12896,N_12729,N_12507);
and U12897 (N_12897,N_12514,N_12184);
nor U12898 (N_12898,N_12744,N_12044);
nand U12899 (N_12899,N_12447,N_12641);
or U12900 (N_12900,N_12027,N_12533);
nand U12901 (N_12901,N_12148,N_12127);
nor U12902 (N_12902,N_12486,N_12269);
nand U12903 (N_12903,N_12499,N_12020);
xor U12904 (N_12904,N_12086,N_12012);
nand U12905 (N_12905,N_12587,N_12170);
and U12906 (N_12906,N_12046,N_12213);
and U12907 (N_12907,N_12483,N_12737);
and U12908 (N_12908,N_12470,N_12741);
and U12909 (N_12909,N_12235,N_12487);
nor U12910 (N_12910,N_12498,N_12604);
and U12911 (N_12911,N_12653,N_12725);
or U12912 (N_12912,N_12383,N_12193);
and U12913 (N_12913,N_12160,N_12634);
or U12914 (N_12914,N_12208,N_12098);
or U12915 (N_12915,N_12723,N_12497);
nor U12916 (N_12916,N_12365,N_12236);
and U12917 (N_12917,N_12089,N_12473);
and U12918 (N_12918,N_12021,N_12338);
nor U12919 (N_12919,N_12692,N_12212);
xnor U12920 (N_12920,N_12015,N_12195);
nand U12921 (N_12921,N_12531,N_12102);
or U12922 (N_12922,N_12273,N_12461);
and U12923 (N_12923,N_12010,N_12452);
nor U12924 (N_12924,N_12600,N_12552);
or U12925 (N_12925,N_12488,N_12351);
nor U12926 (N_12926,N_12035,N_12019);
xnor U12927 (N_12927,N_12368,N_12586);
xnor U12928 (N_12928,N_12701,N_12660);
and U12929 (N_12929,N_12238,N_12186);
nand U12930 (N_12930,N_12175,N_12511);
nor U12931 (N_12931,N_12131,N_12490);
or U12932 (N_12932,N_12179,N_12708);
nand U12933 (N_12933,N_12277,N_12748);
nand U12934 (N_12934,N_12310,N_12298);
nor U12935 (N_12935,N_12326,N_12582);
nand U12936 (N_12936,N_12626,N_12116);
nand U12937 (N_12937,N_12704,N_12410);
nor U12938 (N_12938,N_12617,N_12166);
and U12939 (N_12939,N_12328,N_12085);
xnor U12940 (N_12940,N_12346,N_12058);
and U12941 (N_12941,N_12571,N_12014);
nor U12942 (N_12942,N_12613,N_12290);
nor U12943 (N_12943,N_12394,N_12004);
and U12944 (N_12944,N_12420,N_12087);
nand U12945 (N_12945,N_12547,N_12079);
nand U12946 (N_12946,N_12130,N_12454);
nor U12947 (N_12947,N_12104,N_12373);
or U12948 (N_12948,N_12609,N_12264);
and U12949 (N_12949,N_12445,N_12644);
xnor U12950 (N_12950,N_12640,N_12065);
xnor U12951 (N_12951,N_12423,N_12633);
and U12952 (N_12952,N_12581,N_12139);
nor U12953 (N_12953,N_12074,N_12398);
and U12954 (N_12954,N_12624,N_12100);
or U12955 (N_12955,N_12199,N_12396);
nor U12956 (N_12956,N_12376,N_12695);
and U12957 (N_12957,N_12596,N_12489);
xnor U12958 (N_12958,N_12421,N_12182);
nand U12959 (N_12959,N_12530,N_12426);
xor U12960 (N_12960,N_12448,N_12045);
nor U12961 (N_12961,N_12730,N_12069);
and U12962 (N_12962,N_12555,N_12153);
xnor U12963 (N_12963,N_12431,N_12343);
or U12964 (N_12964,N_12745,N_12189);
nand U12965 (N_12965,N_12585,N_12270);
nor U12966 (N_12966,N_12389,N_12342);
nand U12967 (N_12967,N_12632,N_12667);
or U12968 (N_12968,N_12494,N_12147);
xnor U12969 (N_12969,N_12075,N_12402);
or U12970 (N_12970,N_12746,N_12449);
nand U12971 (N_12971,N_12220,N_12457);
xor U12972 (N_12972,N_12157,N_12059);
nor U12973 (N_12973,N_12367,N_12057);
and U12974 (N_12974,N_12164,N_12223);
or U12975 (N_12975,N_12242,N_12203);
nor U12976 (N_12976,N_12299,N_12111);
nand U12977 (N_12977,N_12141,N_12409);
nand U12978 (N_12978,N_12106,N_12369);
and U12979 (N_12979,N_12017,N_12120);
nand U12980 (N_12980,N_12526,N_12510);
nand U12981 (N_12981,N_12202,N_12400);
and U12982 (N_12982,N_12496,N_12425);
and U12983 (N_12983,N_12214,N_12048);
or U12984 (N_12984,N_12637,N_12005);
nand U12985 (N_12985,N_12331,N_12385);
nand U12986 (N_12986,N_12749,N_12262);
xor U12987 (N_12987,N_12219,N_12205);
or U12988 (N_12988,N_12559,N_12194);
xnor U12989 (N_12989,N_12655,N_12685);
nor U12990 (N_12990,N_12249,N_12524);
xnor U12991 (N_12991,N_12008,N_12736);
and U12992 (N_12992,N_12016,N_12557);
nand U12993 (N_12993,N_12456,N_12658);
xor U12994 (N_12994,N_12714,N_12286);
xor U12995 (N_12995,N_12661,N_12622);
xnor U12996 (N_12996,N_12288,N_12188);
nand U12997 (N_12997,N_12479,N_12689);
xor U12998 (N_12998,N_12623,N_12266);
or U12999 (N_12999,N_12358,N_12198);
and U13000 (N_13000,N_12158,N_12115);
or U13001 (N_13001,N_12315,N_12284);
nor U13002 (N_13002,N_12314,N_12002);
or U13003 (N_13003,N_12009,N_12727);
or U13004 (N_13004,N_12620,N_12304);
xor U13005 (N_13005,N_12408,N_12419);
xor U13006 (N_13006,N_12032,N_12584);
nor U13007 (N_13007,N_12197,N_12502);
or U13008 (N_13008,N_12639,N_12201);
and U13009 (N_13009,N_12216,N_12478);
xor U13010 (N_13010,N_12053,N_12406);
and U13011 (N_13011,N_12023,N_12161);
nor U13012 (N_13012,N_12276,N_12646);
nand U13013 (N_13013,N_12232,N_12172);
nor U13014 (N_13014,N_12556,N_12011);
nand U13015 (N_13015,N_12066,N_12476);
nand U13016 (N_13016,N_12668,N_12656);
or U13017 (N_13017,N_12650,N_12651);
and U13018 (N_13018,N_12372,N_12254);
nor U13019 (N_13019,N_12239,N_12308);
nand U13020 (N_13020,N_12003,N_12485);
or U13021 (N_13021,N_12724,N_12728);
nor U13022 (N_13022,N_12726,N_12401);
nand U13023 (N_13023,N_12034,N_12480);
nand U13024 (N_13024,N_12676,N_12732);
or U13025 (N_13025,N_12541,N_12589);
and U13026 (N_13026,N_12481,N_12455);
xor U13027 (N_13027,N_12173,N_12674);
or U13028 (N_13028,N_12356,N_12274);
xnor U13029 (N_13029,N_12548,N_12165);
xor U13030 (N_13030,N_12305,N_12739);
nand U13031 (N_13031,N_12560,N_12107);
nor U13032 (N_13032,N_12145,N_12519);
and U13033 (N_13033,N_12422,N_12095);
and U13034 (N_13034,N_12484,N_12630);
nand U13035 (N_13035,N_12436,N_12091);
nand U13036 (N_13036,N_12221,N_12344);
nand U13037 (N_13037,N_12691,N_12176);
or U13038 (N_13038,N_12171,N_12450);
nor U13039 (N_13039,N_12731,N_12440);
nor U13040 (N_13040,N_12570,N_12222);
xnor U13041 (N_13041,N_12071,N_12534);
and U13042 (N_13042,N_12719,N_12683);
nor U13043 (N_13043,N_12275,N_12062);
and U13044 (N_13044,N_12740,N_12191);
or U13045 (N_13045,N_12458,N_12033);
or U13046 (N_13046,N_12580,N_12094);
nor U13047 (N_13047,N_12453,N_12244);
nor U13048 (N_13048,N_12355,N_12716);
nand U13049 (N_13049,N_12169,N_12468);
nor U13050 (N_13050,N_12417,N_12629);
and U13051 (N_13051,N_12561,N_12546);
or U13052 (N_13052,N_12318,N_12231);
or U13053 (N_13053,N_12601,N_12593);
or U13054 (N_13054,N_12187,N_12642);
nor U13055 (N_13055,N_12643,N_12038);
or U13056 (N_13056,N_12588,N_12245);
nor U13057 (N_13057,N_12154,N_12595);
nand U13058 (N_13058,N_12329,N_12415);
or U13059 (N_13059,N_12272,N_12386);
or U13060 (N_13060,N_12543,N_12294);
or U13061 (N_13061,N_12688,N_12163);
xor U13062 (N_13062,N_12390,N_12472);
and U13063 (N_13063,N_12397,N_12167);
xnor U13064 (N_13064,N_12506,N_12628);
and U13065 (N_13065,N_12322,N_12363);
xor U13066 (N_13066,N_12060,N_12126);
nor U13067 (N_13067,N_12567,N_12602);
or U13068 (N_13068,N_12703,N_12562);
nand U13069 (N_13069,N_12697,N_12575);
or U13070 (N_13070,N_12670,N_12720);
nor U13071 (N_13071,N_12645,N_12349);
nor U13072 (N_13072,N_12665,N_12067);
nand U13073 (N_13073,N_12155,N_12279);
or U13074 (N_13074,N_12542,N_12492);
xnor U13075 (N_13075,N_12619,N_12052);
or U13076 (N_13076,N_12495,N_12518);
and U13077 (N_13077,N_12430,N_12136);
and U13078 (N_13078,N_12549,N_12092);
nand U13079 (N_13079,N_12503,N_12281);
or U13080 (N_13080,N_12520,N_12654);
xnor U13081 (N_13081,N_12124,N_12206);
nor U13082 (N_13082,N_12553,N_12680);
xor U13083 (N_13083,N_12463,N_12722);
and U13084 (N_13084,N_12399,N_12538);
or U13085 (N_13085,N_12591,N_12414);
or U13086 (N_13086,N_12207,N_12162);
or U13087 (N_13087,N_12101,N_12055);
nand U13088 (N_13088,N_12190,N_12181);
xnor U13089 (N_13089,N_12051,N_12435);
nor U13090 (N_13090,N_12077,N_12225);
and U13091 (N_13091,N_12357,N_12707);
or U13092 (N_13092,N_12671,N_12659);
and U13093 (N_13093,N_12287,N_12080);
nand U13094 (N_13094,N_12416,N_12482);
xor U13095 (N_13095,N_12636,N_12516);
nand U13096 (N_13096,N_12509,N_12064);
nand U13097 (N_13097,N_12564,N_12040);
xnor U13098 (N_13098,N_12713,N_12321);
nand U13099 (N_13099,N_12332,N_12297);
nand U13100 (N_13100,N_12361,N_12237);
and U13101 (N_13101,N_12257,N_12146);
or U13102 (N_13102,N_12241,N_12135);
xnor U13103 (N_13103,N_12742,N_12429);
nand U13104 (N_13104,N_12381,N_12233);
and U13105 (N_13105,N_12140,N_12256);
nor U13106 (N_13106,N_12030,N_12364);
nand U13107 (N_13107,N_12097,N_12252);
or U13108 (N_13108,N_12709,N_12504);
and U13109 (N_13109,N_12353,N_12605);
and U13110 (N_13110,N_12054,N_12525);
and U13111 (N_13111,N_12618,N_12307);
nor U13112 (N_13112,N_12192,N_12036);
nor U13113 (N_13113,N_12384,N_12370);
and U13114 (N_13114,N_12240,N_12681);
xnor U13115 (N_13115,N_12341,N_12316);
nor U13116 (N_13116,N_12296,N_12663);
nor U13117 (N_13117,N_12265,N_12412);
and U13118 (N_13118,N_12259,N_12614);
nand U13119 (N_13119,N_12523,N_12374);
or U13120 (N_13120,N_12063,N_12606);
or U13121 (N_13121,N_12411,N_12702);
and U13122 (N_13122,N_12712,N_12459);
nor U13123 (N_13123,N_12366,N_12253);
xor U13124 (N_13124,N_12577,N_12295);
nor U13125 (N_13125,N_12604,N_12079);
xnor U13126 (N_13126,N_12465,N_12298);
nor U13127 (N_13127,N_12239,N_12539);
and U13128 (N_13128,N_12702,N_12082);
nor U13129 (N_13129,N_12096,N_12619);
or U13130 (N_13130,N_12343,N_12377);
or U13131 (N_13131,N_12552,N_12388);
xnor U13132 (N_13132,N_12581,N_12471);
nor U13133 (N_13133,N_12258,N_12318);
xnor U13134 (N_13134,N_12166,N_12602);
nand U13135 (N_13135,N_12424,N_12270);
xor U13136 (N_13136,N_12561,N_12016);
and U13137 (N_13137,N_12678,N_12467);
nor U13138 (N_13138,N_12271,N_12556);
or U13139 (N_13139,N_12156,N_12397);
xnor U13140 (N_13140,N_12110,N_12376);
or U13141 (N_13141,N_12571,N_12200);
xor U13142 (N_13142,N_12216,N_12645);
or U13143 (N_13143,N_12682,N_12713);
xor U13144 (N_13144,N_12550,N_12067);
or U13145 (N_13145,N_12682,N_12569);
or U13146 (N_13146,N_12465,N_12062);
nor U13147 (N_13147,N_12353,N_12542);
xnor U13148 (N_13148,N_12366,N_12673);
nor U13149 (N_13149,N_12260,N_12593);
nor U13150 (N_13150,N_12597,N_12128);
xnor U13151 (N_13151,N_12560,N_12174);
nand U13152 (N_13152,N_12664,N_12598);
nor U13153 (N_13153,N_12436,N_12057);
nor U13154 (N_13154,N_12617,N_12632);
and U13155 (N_13155,N_12739,N_12114);
xnor U13156 (N_13156,N_12614,N_12347);
or U13157 (N_13157,N_12716,N_12114);
or U13158 (N_13158,N_12537,N_12181);
nor U13159 (N_13159,N_12199,N_12133);
nand U13160 (N_13160,N_12354,N_12405);
or U13161 (N_13161,N_12523,N_12539);
nand U13162 (N_13162,N_12128,N_12236);
xor U13163 (N_13163,N_12128,N_12111);
xor U13164 (N_13164,N_12339,N_12184);
xor U13165 (N_13165,N_12264,N_12652);
nand U13166 (N_13166,N_12451,N_12387);
nor U13167 (N_13167,N_12325,N_12199);
or U13168 (N_13168,N_12322,N_12038);
or U13169 (N_13169,N_12188,N_12457);
or U13170 (N_13170,N_12313,N_12728);
nor U13171 (N_13171,N_12564,N_12168);
xor U13172 (N_13172,N_12311,N_12321);
and U13173 (N_13173,N_12238,N_12386);
nor U13174 (N_13174,N_12384,N_12017);
nand U13175 (N_13175,N_12281,N_12483);
nor U13176 (N_13176,N_12574,N_12469);
nand U13177 (N_13177,N_12390,N_12669);
and U13178 (N_13178,N_12651,N_12657);
xor U13179 (N_13179,N_12110,N_12329);
or U13180 (N_13180,N_12649,N_12520);
xor U13181 (N_13181,N_12266,N_12067);
nand U13182 (N_13182,N_12004,N_12736);
or U13183 (N_13183,N_12369,N_12033);
xor U13184 (N_13184,N_12373,N_12263);
xor U13185 (N_13185,N_12716,N_12172);
xnor U13186 (N_13186,N_12455,N_12673);
nor U13187 (N_13187,N_12431,N_12051);
xnor U13188 (N_13188,N_12713,N_12324);
nand U13189 (N_13189,N_12661,N_12573);
or U13190 (N_13190,N_12068,N_12593);
nand U13191 (N_13191,N_12029,N_12032);
or U13192 (N_13192,N_12131,N_12271);
xor U13193 (N_13193,N_12245,N_12643);
nand U13194 (N_13194,N_12669,N_12552);
or U13195 (N_13195,N_12362,N_12005);
nand U13196 (N_13196,N_12304,N_12176);
nor U13197 (N_13197,N_12150,N_12110);
nand U13198 (N_13198,N_12398,N_12127);
and U13199 (N_13199,N_12202,N_12038);
nand U13200 (N_13200,N_12591,N_12552);
and U13201 (N_13201,N_12118,N_12643);
xnor U13202 (N_13202,N_12512,N_12577);
or U13203 (N_13203,N_12308,N_12101);
nand U13204 (N_13204,N_12604,N_12198);
and U13205 (N_13205,N_12659,N_12406);
nand U13206 (N_13206,N_12591,N_12507);
nor U13207 (N_13207,N_12589,N_12263);
and U13208 (N_13208,N_12637,N_12184);
and U13209 (N_13209,N_12504,N_12578);
or U13210 (N_13210,N_12033,N_12456);
or U13211 (N_13211,N_12515,N_12742);
or U13212 (N_13212,N_12079,N_12055);
xnor U13213 (N_13213,N_12254,N_12493);
xor U13214 (N_13214,N_12427,N_12419);
and U13215 (N_13215,N_12435,N_12513);
nor U13216 (N_13216,N_12691,N_12511);
nand U13217 (N_13217,N_12109,N_12509);
nor U13218 (N_13218,N_12467,N_12580);
and U13219 (N_13219,N_12085,N_12007);
xor U13220 (N_13220,N_12446,N_12745);
xnor U13221 (N_13221,N_12192,N_12003);
or U13222 (N_13222,N_12654,N_12161);
nand U13223 (N_13223,N_12517,N_12280);
or U13224 (N_13224,N_12502,N_12627);
xnor U13225 (N_13225,N_12417,N_12552);
or U13226 (N_13226,N_12167,N_12347);
or U13227 (N_13227,N_12024,N_12590);
xor U13228 (N_13228,N_12102,N_12084);
nor U13229 (N_13229,N_12261,N_12427);
nand U13230 (N_13230,N_12733,N_12479);
nand U13231 (N_13231,N_12473,N_12279);
xnor U13232 (N_13232,N_12501,N_12656);
nor U13233 (N_13233,N_12048,N_12724);
nor U13234 (N_13234,N_12000,N_12293);
and U13235 (N_13235,N_12273,N_12483);
or U13236 (N_13236,N_12399,N_12687);
nor U13237 (N_13237,N_12408,N_12251);
and U13238 (N_13238,N_12396,N_12251);
nor U13239 (N_13239,N_12536,N_12528);
and U13240 (N_13240,N_12625,N_12595);
nand U13241 (N_13241,N_12525,N_12144);
xor U13242 (N_13242,N_12053,N_12133);
or U13243 (N_13243,N_12585,N_12403);
nand U13244 (N_13244,N_12584,N_12072);
nand U13245 (N_13245,N_12266,N_12188);
nor U13246 (N_13246,N_12092,N_12196);
nand U13247 (N_13247,N_12035,N_12433);
xor U13248 (N_13248,N_12387,N_12345);
xnor U13249 (N_13249,N_12352,N_12254);
xnor U13250 (N_13250,N_12728,N_12351);
nand U13251 (N_13251,N_12147,N_12453);
and U13252 (N_13252,N_12480,N_12247);
and U13253 (N_13253,N_12603,N_12419);
xnor U13254 (N_13254,N_12585,N_12728);
nand U13255 (N_13255,N_12025,N_12727);
and U13256 (N_13256,N_12669,N_12024);
nor U13257 (N_13257,N_12668,N_12438);
nand U13258 (N_13258,N_12028,N_12408);
nand U13259 (N_13259,N_12093,N_12653);
xnor U13260 (N_13260,N_12549,N_12294);
xor U13261 (N_13261,N_12089,N_12467);
xor U13262 (N_13262,N_12312,N_12042);
or U13263 (N_13263,N_12177,N_12386);
xor U13264 (N_13264,N_12685,N_12668);
nor U13265 (N_13265,N_12156,N_12539);
nand U13266 (N_13266,N_12366,N_12402);
xor U13267 (N_13267,N_12547,N_12191);
nor U13268 (N_13268,N_12193,N_12462);
xnor U13269 (N_13269,N_12093,N_12458);
nand U13270 (N_13270,N_12184,N_12402);
xor U13271 (N_13271,N_12233,N_12417);
nand U13272 (N_13272,N_12642,N_12695);
and U13273 (N_13273,N_12689,N_12558);
nand U13274 (N_13274,N_12126,N_12417);
or U13275 (N_13275,N_12487,N_12234);
nand U13276 (N_13276,N_12236,N_12320);
nor U13277 (N_13277,N_12551,N_12357);
or U13278 (N_13278,N_12620,N_12485);
and U13279 (N_13279,N_12569,N_12174);
xor U13280 (N_13280,N_12284,N_12598);
nand U13281 (N_13281,N_12012,N_12746);
nor U13282 (N_13282,N_12361,N_12393);
nor U13283 (N_13283,N_12362,N_12026);
or U13284 (N_13284,N_12056,N_12294);
or U13285 (N_13285,N_12255,N_12315);
nor U13286 (N_13286,N_12395,N_12240);
nor U13287 (N_13287,N_12130,N_12735);
nand U13288 (N_13288,N_12075,N_12557);
or U13289 (N_13289,N_12174,N_12168);
nand U13290 (N_13290,N_12055,N_12536);
xor U13291 (N_13291,N_12356,N_12472);
or U13292 (N_13292,N_12033,N_12466);
nor U13293 (N_13293,N_12188,N_12270);
xor U13294 (N_13294,N_12264,N_12238);
nor U13295 (N_13295,N_12588,N_12393);
nor U13296 (N_13296,N_12565,N_12292);
and U13297 (N_13297,N_12320,N_12258);
and U13298 (N_13298,N_12023,N_12234);
and U13299 (N_13299,N_12077,N_12617);
nor U13300 (N_13300,N_12366,N_12020);
and U13301 (N_13301,N_12727,N_12520);
nor U13302 (N_13302,N_12692,N_12562);
or U13303 (N_13303,N_12698,N_12320);
and U13304 (N_13304,N_12056,N_12084);
nand U13305 (N_13305,N_12113,N_12669);
nor U13306 (N_13306,N_12480,N_12713);
or U13307 (N_13307,N_12327,N_12159);
nor U13308 (N_13308,N_12509,N_12575);
nand U13309 (N_13309,N_12705,N_12153);
or U13310 (N_13310,N_12183,N_12239);
nor U13311 (N_13311,N_12402,N_12745);
nand U13312 (N_13312,N_12072,N_12540);
xnor U13313 (N_13313,N_12644,N_12061);
or U13314 (N_13314,N_12443,N_12723);
or U13315 (N_13315,N_12655,N_12398);
nor U13316 (N_13316,N_12092,N_12681);
or U13317 (N_13317,N_12551,N_12078);
nor U13318 (N_13318,N_12104,N_12048);
nor U13319 (N_13319,N_12714,N_12023);
nor U13320 (N_13320,N_12432,N_12689);
and U13321 (N_13321,N_12155,N_12470);
or U13322 (N_13322,N_12062,N_12178);
nand U13323 (N_13323,N_12495,N_12583);
xnor U13324 (N_13324,N_12225,N_12253);
nor U13325 (N_13325,N_12734,N_12653);
or U13326 (N_13326,N_12648,N_12621);
nor U13327 (N_13327,N_12545,N_12259);
xor U13328 (N_13328,N_12392,N_12225);
nand U13329 (N_13329,N_12654,N_12221);
nor U13330 (N_13330,N_12704,N_12155);
xnor U13331 (N_13331,N_12429,N_12433);
xnor U13332 (N_13332,N_12749,N_12186);
xor U13333 (N_13333,N_12008,N_12177);
or U13334 (N_13334,N_12353,N_12392);
or U13335 (N_13335,N_12457,N_12285);
nor U13336 (N_13336,N_12371,N_12274);
or U13337 (N_13337,N_12512,N_12605);
xor U13338 (N_13338,N_12042,N_12561);
nor U13339 (N_13339,N_12576,N_12489);
or U13340 (N_13340,N_12179,N_12469);
and U13341 (N_13341,N_12106,N_12453);
and U13342 (N_13342,N_12738,N_12350);
and U13343 (N_13343,N_12624,N_12424);
nor U13344 (N_13344,N_12063,N_12521);
nand U13345 (N_13345,N_12280,N_12294);
and U13346 (N_13346,N_12633,N_12583);
and U13347 (N_13347,N_12440,N_12049);
nand U13348 (N_13348,N_12173,N_12031);
nand U13349 (N_13349,N_12252,N_12444);
and U13350 (N_13350,N_12091,N_12693);
nand U13351 (N_13351,N_12743,N_12561);
nor U13352 (N_13352,N_12531,N_12272);
nand U13353 (N_13353,N_12530,N_12505);
nand U13354 (N_13354,N_12736,N_12278);
or U13355 (N_13355,N_12208,N_12497);
or U13356 (N_13356,N_12463,N_12659);
nand U13357 (N_13357,N_12060,N_12597);
xnor U13358 (N_13358,N_12731,N_12373);
nor U13359 (N_13359,N_12192,N_12051);
and U13360 (N_13360,N_12034,N_12097);
and U13361 (N_13361,N_12596,N_12261);
xor U13362 (N_13362,N_12603,N_12194);
nand U13363 (N_13363,N_12309,N_12151);
xnor U13364 (N_13364,N_12529,N_12654);
nor U13365 (N_13365,N_12232,N_12136);
nand U13366 (N_13366,N_12602,N_12664);
xor U13367 (N_13367,N_12403,N_12065);
and U13368 (N_13368,N_12170,N_12306);
and U13369 (N_13369,N_12682,N_12079);
and U13370 (N_13370,N_12574,N_12656);
xnor U13371 (N_13371,N_12135,N_12352);
nor U13372 (N_13372,N_12157,N_12203);
or U13373 (N_13373,N_12412,N_12610);
or U13374 (N_13374,N_12473,N_12465);
and U13375 (N_13375,N_12491,N_12089);
xnor U13376 (N_13376,N_12262,N_12194);
nor U13377 (N_13377,N_12149,N_12021);
and U13378 (N_13378,N_12004,N_12316);
or U13379 (N_13379,N_12332,N_12519);
nand U13380 (N_13380,N_12125,N_12334);
or U13381 (N_13381,N_12192,N_12523);
and U13382 (N_13382,N_12151,N_12173);
nor U13383 (N_13383,N_12426,N_12556);
or U13384 (N_13384,N_12628,N_12522);
xnor U13385 (N_13385,N_12246,N_12569);
nand U13386 (N_13386,N_12170,N_12533);
nand U13387 (N_13387,N_12476,N_12620);
and U13388 (N_13388,N_12147,N_12627);
nand U13389 (N_13389,N_12003,N_12033);
and U13390 (N_13390,N_12738,N_12082);
xnor U13391 (N_13391,N_12117,N_12703);
xnor U13392 (N_13392,N_12732,N_12348);
nand U13393 (N_13393,N_12080,N_12356);
xor U13394 (N_13394,N_12086,N_12220);
and U13395 (N_13395,N_12455,N_12594);
nor U13396 (N_13396,N_12381,N_12341);
nand U13397 (N_13397,N_12080,N_12491);
nand U13398 (N_13398,N_12470,N_12010);
or U13399 (N_13399,N_12580,N_12726);
nand U13400 (N_13400,N_12661,N_12529);
nand U13401 (N_13401,N_12294,N_12146);
and U13402 (N_13402,N_12184,N_12597);
nand U13403 (N_13403,N_12256,N_12616);
nand U13404 (N_13404,N_12544,N_12183);
xor U13405 (N_13405,N_12695,N_12632);
or U13406 (N_13406,N_12627,N_12547);
xor U13407 (N_13407,N_12074,N_12245);
and U13408 (N_13408,N_12427,N_12625);
or U13409 (N_13409,N_12017,N_12029);
and U13410 (N_13410,N_12723,N_12301);
nor U13411 (N_13411,N_12260,N_12555);
nand U13412 (N_13412,N_12682,N_12491);
nand U13413 (N_13413,N_12681,N_12193);
nand U13414 (N_13414,N_12068,N_12271);
xnor U13415 (N_13415,N_12603,N_12396);
or U13416 (N_13416,N_12588,N_12167);
and U13417 (N_13417,N_12596,N_12621);
and U13418 (N_13418,N_12095,N_12213);
or U13419 (N_13419,N_12298,N_12137);
nand U13420 (N_13420,N_12393,N_12555);
or U13421 (N_13421,N_12612,N_12560);
nand U13422 (N_13422,N_12531,N_12454);
or U13423 (N_13423,N_12517,N_12039);
nand U13424 (N_13424,N_12652,N_12238);
or U13425 (N_13425,N_12323,N_12235);
or U13426 (N_13426,N_12531,N_12602);
nor U13427 (N_13427,N_12223,N_12326);
nor U13428 (N_13428,N_12182,N_12348);
and U13429 (N_13429,N_12045,N_12176);
xor U13430 (N_13430,N_12598,N_12391);
or U13431 (N_13431,N_12385,N_12013);
or U13432 (N_13432,N_12733,N_12689);
nor U13433 (N_13433,N_12084,N_12127);
and U13434 (N_13434,N_12305,N_12524);
nand U13435 (N_13435,N_12685,N_12002);
or U13436 (N_13436,N_12426,N_12709);
nand U13437 (N_13437,N_12637,N_12629);
or U13438 (N_13438,N_12550,N_12573);
and U13439 (N_13439,N_12585,N_12183);
nor U13440 (N_13440,N_12342,N_12250);
nand U13441 (N_13441,N_12261,N_12667);
and U13442 (N_13442,N_12565,N_12501);
xnor U13443 (N_13443,N_12131,N_12187);
and U13444 (N_13444,N_12075,N_12500);
nor U13445 (N_13445,N_12017,N_12531);
xnor U13446 (N_13446,N_12458,N_12396);
or U13447 (N_13447,N_12673,N_12127);
nor U13448 (N_13448,N_12056,N_12650);
nand U13449 (N_13449,N_12158,N_12205);
nor U13450 (N_13450,N_12299,N_12551);
nor U13451 (N_13451,N_12738,N_12258);
nand U13452 (N_13452,N_12262,N_12589);
or U13453 (N_13453,N_12100,N_12003);
nand U13454 (N_13454,N_12501,N_12029);
or U13455 (N_13455,N_12277,N_12188);
nand U13456 (N_13456,N_12045,N_12477);
nor U13457 (N_13457,N_12298,N_12096);
nand U13458 (N_13458,N_12226,N_12276);
or U13459 (N_13459,N_12014,N_12180);
xnor U13460 (N_13460,N_12352,N_12474);
and U13461 (N_13461,N_12492,N_12217);
nor U13462 (N_13462,N_12172,N_12348);
and U13463 (N_13463,N_12248,N_12549);
nor U13464 (N_13464,N_12406,N_12061);
or U13465 (N_13465,N_12509,N_12002);
and U13466 (N_13466,N_12498,N_12292);
xor U13467 (N_13467,N_12690,N_12640);
xor U13468 (N_13468,N_12653,N_12194);
nand U13469 (N_13469,N_12683,N_12481);
or U13470 (N_13470,N_12480,N_12532);
or U13471 (N_13471,N_12174,N_12273);
nand U13472 (N_13472,N_12499,N_12366);
and U13473 (N_13473,N_12261,N_12132);
xnor U13474 (N_13474,N_12391,N_12581);
and U13475 (N_13475,N_12180,N_12134);
and U13476 (N_13476,N_12532,N_12437);
nand U13477 (N_13477,N_12016,N_12401);
xnor U13478 (N_13478,N_12413,N_12389);
xor U13479 (N_13479,N_12428,N_12693);
and U13480 (N_13480,N_12577,N_12681);
xor U13481 (N_13481,N_12555,N_12635);
and U13482 (N_13482,N_12423,N_12226);
and U13483 (N_13483,N_12634,N_12102);
nor U13484 (N_13484,N_12016,N_12690);
nor U13485 (N_13485,N_12002,N_12514);
nor U13486 (N_13486,N_12477,N_12743);
and U13487 (N_13487,N_12510,N_12709);
or U13488 (N_13488,N_12584,N_12696);
nor U13489 (N_13489,N_12007,N_12439);
xnor U13490 (N_13490,N_12508,N_12580);
nor U13491 (N_13491,N_12246,N_12064);
nand U13492 (N_13492,N_12677,N_12628);
xor U13493 (N_13493,N_12430,N_12392);
or U13494 (N_13494,N_12290,N_12133);
nand U13495 (N_13495,N_12299,N_12631);
nor U13496 (N_13496,N_12119,N_12531);
and U13497 (N_13497,N_12107,N_12208);
and U13498 (N_13498,N_12313,N_12492);
nor U13499 (N_13499,N_12292,N_12220);
xor U13500 (N_13500,N_13414,N_12908);
and U13501 (N_13501,N_12839,N_12847);
or U13502 (N_13502,N_13081,N_13492);
xor U13503 (N_13503,N_12900,N_13082);
or U13504 (N_13504,N_13441,N_13011);
nand U13505 (N_13505,N_13243,N_13387);
or U13506 (N_13506,N_13267,N_13286);
and U13507 (N_13507,N_13303,N_13352);
xor U13508 (N_13508,N_12957,N_12833);
xor U13509 (N_13509,N_13177,N_13094);
nor U13510 (N_13510,N_13043,N_13460);
xor U13511 (N_13511,N_12815,N_13151);
and U13512 (N_13512,N_12841,N_13042);
xor U13513 (N_13513,N_13284,N_13401);
xnor U13514 (N_13514,N_13174,N_13224);
nand U13515 (N_13515,N_13464,N_13411);
xor U13516 (N_13516,N_13100,N_13426);
nor U13517 (N_13517,N_13214,N_12765);
nor U13518 (N_13518,N_12934,N_12972);
or U13519 (N_13519,N_13476,N_13375);
nor U13520 (N_13520,N_12905,N_12946);
or U13521 (N_13521,N_13415,N_12901);
nand U13522 (N_13522,N_13465,N_13257);
and U13523 (N_13523,N_13144,N_13193);
xnor U13524 (N_13524,N_13312,N_13106);
and U13525 (N_13525,N_13205,N_13156);
and U13526 (N_13526,N_13485,N_12903);
and U13527 (N_13527,N_12964,N_12912);
nand U13528 (N_13528,N_13330,N_12853);
or U13529 (N_13529,N_13201,N_12759);
nor U13530 (N_13530,N_13351,N_13064);
xnor U13531 (N_13531,N_12933,N_13425);
nand U13532 (N_13532,N_12857,N_13198);
nand U13533 (N_13533,N_12860,N_13127);
nor U13534 (N_13534,N_12898,N_13489);
xor U13535 (N_13535,N_12862,N_13037);
and U13536 (N_13536,N_13095,N_13114);
nor U13537 (N_13537,N_13435,N_13110);
nand U13538 (N_13538,N_13399,N_13164);
xor U13539 (N_13539,N_12775,N_12866);
or U13540 (N_13540,N_13305,N_13413);
xor U13541 (N_13541,N_13368,N_13188);
nand U13542 (N_13542,N_13341,N_13204);
and U13543 (N_13543,N_13402,N_13310);
nor U13544 (N_13544,N_13072,N_13221);
or U13545 (N_13545,N_13484,N_13486);
nand U13546 (N_13546,N_12940,N_13113);
xor U13547 (N_13547,N_13480,N_12921);
nand U13548 (N_13548,N_13124,N_12819);
and U13549 (N_13549,N_12896,N_13481);
and U13550 (N_13550,N_13051,N_13248);
and U13551 (N_13551,N_13382,N_13390);
and U13552 (N_13552,N_12965,N_13207);
and U13553 (N_13553,N_13115,N_13394);
nor U13554 (N_13554,N_13142,N_13308);
nand U13555 (N_13555,N_12913,N_13009);
nor U13556 (N_13556,N_13470,N_12872);
nand U13557 (N_13557,N_13007,N_13107);
nand U13558 (N_13558,N_13105,N_12973);
nand U13559 (N_13559,N_12968,N_13377);
nor U13560 (N_13560,N_13167,N_13398);
nand U13561 (N_13561,N_12779,N_13266);
xnor U13562 (N_13562,N_13227,N_13317);
xor U13563 (N_13563,N_13490,N_13309);
nand U13564 (N_13564,N_13443,N_13208);
nand U13565 (N_13565,N_13469,N_12832);
xnor U13566 (N_13566,N_12978,N_12825);
nand U13567 (N_13567,N_13463,N_13274);
and U13568 (N_13568,N_12971,N_13129);
or U13569 (N_13569,N_13391,N_12774);
nor U13570 (N_13570,N_13288,N_13392);
nor U13571 (N_13571,N_13001,N_13334);
and U13572 (N_13572,N_13218,N_13119);
and U13573 (N_13573,N_13272,N_12776);
or U13574 (N_13574,N_12751,N_13249);
and U13575 (N_13575,N_12920,N_13121);
xor U13576 (N_13576,N_13353,N_12999);
xnor U13577 (N_13577,N_13191,N_12889);
or U13578 (N_13578,N_12991,N_13455);
nand U13579 (N_13579,N_13373,N_12918);
xor U13580 (N_13580,N_12909,N_13196);
or U13581 (N_13581,N_13275,N_13062);
nand U13582 (N_13582,N_13233,N_12880);
and U13583 (N_13583,N_13182,N_13141);
xor U13584 (N_13584,N_12958,N_13098);
and U13585 (N_13585,N_13152,N_12855);
nand U13586 (N_13586,N_13299,N_13349);
or U13587 (N_13587,N_13298,N_13245);
nand U13588 (N_13588,N_13319,N_12788);
and U13589 (N_13589,N_12888,N_13358);
nor U13590 (N_13590,N_12840,N_12810);
nand U13591 (N_13591,N_12783,N_13383);
and U13592 (N_13592,N_13168,N_12930);
nor U13593 (N_13593,N_13421,N_13423);
xnor U13594 (N_13594,N_13154,N_13217);
nor U13595 (N_13595,N_13035,N_12809);
nor U13596 (N_13596,N_13070,N_12984);
or U13597 (N_13597,N_12952,N_12950);
nor U13598 (N_13598,N_12975,N_12969);
nand U13599 (N_13599,N_12789,N_13462);
and U13600 (N_13600,N_12791,N_13241);
and U13601 (N_13601,N_13451,N_13483);
nand U13602 (N_13602,N_12937,N_12773);
or U13603 (N_13603,N_13041,N_13192);
xor U13604 (N_13604,N_12769,N_13270);
xor U13605 (N_13605,N_12797,N_13091);
nor U13606 (N_13606,N_13102,N_13161);
and U13607 (N_13607,N_12931,N_13336);
or U13608 (N_13608,N_13276,N_13406);
and U13609 (N_13609,N_12895,N_13316);
nand U13610 (N_13610,N_13172,N_13295);
and U13611 (N_13611,N_12928,N_13005);
or U13612 (N_13612,N_13326,N_12959);
nand U13613 (N_13613,N_12761,N_13291);
or U13614 (N_13614,N_13194,N_12807);
xnor U13615 (N_13615,N_13003,N_13021);
or U13616 (N_13616,N_12942,N_12846);
or U13617 (N_13617,N_12793,N_13246);
or U13618 (N_13618,N_13431,N_12827);
xor U13619 (N_13619,N_12836,N_13340);
nand U13620 (N_13620,N_13211,N_13123);
nor U13621 (N_13621,N_13120,N_12814);
and U13622 (N_13622,N_13439,N_12987);
and U13623 (N_13623,N_13150,N_13364);
nor U13624 (N_13624,N_13499,N_12886);
xor U13625 (N_13625,N_12870,N_12760);
or U13626 (N_13626,N_13418,N_12763);
and U13627 (N_13627,N_13342,N_12954);
and U13628 (N_13628,N_13496,N_12838);
nor U13629 (N_13629,N_12976,N_13006);
nand U13630 (N_13630,N_13442,N_13149);
nor U13631 (N_13631,N_13103,N_12925);
or U13632 (N_13632,N_13494,N_13283);
or U13633 (N_13633,N_13016,N_12885);
xor U13634 (N_13634,N_13446,N_13086);
or U13635 (N_13635,N_12842,N_12963);
nor U13636 (N_13636,N_13289,N_12906);
nor U13637 (N_13637,N_12828,N_13153);
nand U13638 (N_13638,N_13117,N_13228);
nor U13639 (N_13639,N_13200,N_13139);
nand U13640 (N_13640,N_13143,N_13017);
nand U13641 (N_13641,N_13447,N_13047);
xor U13642 (N_13642,N_13449,N_13077);
xor U13643 (N_13643,N_13058,N_12758);
and U13644 (N_13644,N_13277,N_13067);
or U13645 (N_13645,N_12997,N_12831);
and U13646 (N_13646,N_13432,N_13090);
xor U13647 (N_13647,N_13258,N_13032);
or U13648 (N_13648,N_12877,N_13155);
nor U13649 (N_13649,N_12803,N_13474);
or U13650 (N_13650,N_12935,N_12891);
nor U13651 (N_13651,N_13050,N_13213);
or U13652 (N_13652,N_13126,N_12943);
or U13653 (N_13653,N_12820,N_13203);
nor U13654 (N_13654,N_12923,N_13018);
nand U13655 (N_13655,N_13458,N_12786);
nand U13656 (N_13656,N_12936,N_13345);
nor U13657 (N_13657,N_13456,N_13491);
nand U13658 (N_13658,N_13222,N_13410);
and U13659 (N_13659,N_13256,N_13393);
xnor U13660 (N_13660,N_13220,N_13014);
nor U13661 (N_13661,N_12869,N_12829);
nand U13662 (N_13662,N_12823,N_12874);
and U13663 (N_13663,N_13362,N_12953);
or U13664 (N_13664,N_13029,N_12985);
nand U13665 (N_13665,N_12893,N_12939);
nand U13666 (N_13666,N_13122,N_12995);
nor U13667 (N_13667,N_13273,N_13053);
and U13668 (N_13668,N_13135,N_13173);
and U13669 (N_13669,N_13263,N_12911);
nor U13670 (N_13670,N_13428,N_13370);
xnor U13671 (N_13671,N_13287,N_13015);
or U13672 (N_13672,N_13031,N_13417);
nor U13673 (N_13673,N_13337,N_13332);
or U13674 (N_13674,N_12910,N_13379);
and U13675 (N_13675,N_13453,N_13374);
and U13676 (N_13676,N_13049,N_13381);
and U13677 (N_13677,N_13092,N_13136);
or U13678 (N_13678,N_13012,N_13473);
or U13679 (N_13679,N_12899,N_13422);
xor U13680 (N_13680,N_12945,N_12979);
xor U13681 (N_13681,N_12816,N_12917);
nor U13682 (N_13682,N_13323,N_13259);
and U13683 (N_13683,N_13096,N_12817);
and U13684 (N_13684,N_13322,N_12998);
or U13685 (N_13685,N_13075,N_13089);
nand U13686 (N_13686,N_12805,N_13229);
nand U13687 (N_13687,N_13230,N_13297);
nand U13688 (N_13688,N_13268,N_13147);
nor U13689 (N_13689,N_13450,N_13157);
nand U13690 (N_13690,N_13396,N_12983);
and U13691 (N_13691,N_12851,N_13118);
nor U13692 (N_13692,N_13159,N_13290);
nand U13693 (N_13693,N_12882,N_13372);
and U13694 (N_13694,N_13242,N_13493);
and U13695 (N_13695,N_13216,N_13088);
and U13696 (N_13696,N_13479,N_13388);
nand U13697 (N_13697,N_12941,N_13355);
nor U13698 (N_13698,N_13344,N_13125);
nor U13699 (N_13699,N_13137,N_12753);
or U13700 (N_13700,N_13285,N_13033);
nand U13701 (N_13701,N_12990,N_12951);
nand U13702 (N_13702,N_13302,N_13335);
and U13703 (N_13703,N_12854,N_13386);
nand U13704 (N_13704,N_13461,N_13408);
and U13705 (N_13705,N_13130,N_12821);
and U13706 (N_13706,N_12927,N_12777);
nor U13707 (N_13707,N_13027,N_13145);
or U13708 (N_13708,N_13436,N_13024);
nand U13709 (N_13709,N_12986,N_12795);
xnor U13710 (N_13710,N_13467,N_13178);
or U13711 (N_13711,N_13262,N_12892);
xnor U13712 (N_13712,N_13348,N_13293);
and U13713 (N_13713,N_13099,N_13071);
xor U13714 (N_13714,N_12926,N_13325);
xor U13715 (N_13715,N_13260,N_13294);
xor U13716 (N_13716,N_12770,N_12919);
or U13717 (N_13717,N_12792,N_13186);
or U13718 (N_13718,N_12755,N_13400);
nor U13719 (N_13719,N_13101,N_13165);
xor U13720 (N_13720,N_13300,N_12980);
and U13721 (N_13721,N_12808,N_12822);
xor U13722 (N_13722,N_13281,N_12812);
or U13723 (N_13723,N_12782,N_13472);
xnor U13724 (N_13724,N_13429,N_13189);
nor U13725 (N_13725,N_13002,N_13466);
or U13726 (N_13726,N_12904,N_13199);
xor U13727 (N_13727,N_13251,N_13269);
nor U13728 (N_13728,N_13320,N_12757);
xor U13729 (N_13729,N_12837,N_13104);
nor U13730 (N_13730,N_13360,N_13111);
nor U13731 (N_13731,N_13057,N_12982);
nand U13732 (N_13732,N_13440,N_13482);
xnor U13733 (N_13733,N_12859,N_13069);
or U13734 (N_13734,N_13225,N_13219);
nand U13735 (N_13735,N_13244,N_12844);
nor U13736 (N_13736,N_13404,N_13039);
nand U13737 (N_13737,N_12806,N_13314);
nor U13738 (N_13738,N_12868,N_13471);
xor U13739 (N_13739,N_12852,N_12752);
nand U13740 (N_13740,N_12944,N_13066);
nor U13741 (N_13741,N_12875,N_12798);
xnor U13742 (N_13742,N_12989,N_12813);
nand U13743 (N_13743,N_13389,N_12878);
or U13744 (N_13744,N_13056,N_13495);
and U13745 (N_13745,N_13369,N_12916);
xnor U13746 (N_13746,N_12861,N_13055);
xor U13747 (N_13747,N_13347,N_13022);
or U13748 (N_13748,N_12938,N_13183);
xnor U13749 (N_13749,N_13475,N_13231);
xnor U13750 (N_13750,N_12960,N_12858);
xor U13751 (N_13751,N_12994,N_12849);
xnor U13752 (N_13752,N_13264,N_13040);
nand U13753 (N_13753,N_13457,N_13255);
and U13754 (N_13754,N_13052,N_13278);
or U13755 (N_13755,N_13197,N_12830);
nor U13756 (N_13756,N_13282,N_13328);
nor U13757 (N_13757,N_13063,N_13010);
and U13758 (N_13758,N_12800,N_13280);
or U13759 (N_13759,N_12996,N_13146);
and U13760 (N_13760,N_13138,N_12756);
xor U13761 (N_13761,N_12887,N_12780);
or U13762 (N_13762,N_13030,N_13215);
nand U13763 (N_13763,N_13020,N_12826);
or U13764 (N_13764,N_12949,N_13301);
or U13765 (N_13765,N_12845,N_12867);
or U13766 (N_13766,N_13430,N_12790);
nand U13767 (N_13767,N_13433,N_13148);
nor U13768 (N_13768,N_12824,N_12915);
or U13769 (N_13769,N_13023,N_13468);
xnor U13770 (N_13770,N_13498,N_13307);
or U13771 (N_13771,N_13079,N_12929);
xnor U13772 (N_13772,N_13250,N_13253);
xor U13773 (N_13773,N_13419,N_13327);
nand U13774 (N_13774,N_13279,N_12865);
and U13775 (N_13775,N_13085,N_13160);
nand U13776 (N_13776,N_12932,N_13363);
or U13777 (N_13777,N_13254,N_12766);
nor U13778 (N_13778,N_13292,N_13179);
nor U13779 (N_13779,N_13008,N_12835);
nor U13780 (N_13780,N_13026,N_13065);
or U13781 (N_13781,N_12796,N_13271);
nand U13782 (N_13782,N_12881,N_13420);
nor U13783 (N_13783,N_13108,N_13346);
or U13784 (N_13784,N_13180,N_12768);
or U13785 (N_13785,N_13331,N_13190);
xnor U13786 (N_13786,N_13350,N_12811);
or U13787 (N_13787,N_13166,N_12962);
nor U13788 (N_13788,N_13234,N_13434);
and U13789 (N_13789,N_12981,N_13185);
nand U13790 (N_13790,N_13397,N_12974);
or U13791 (N_13791,N_12977,N_13184);
nor U13792 (N_13792,N_12988,N_12754);
or U13793 (N_13793,N_12778,N_12956);
or U13794 (N_13794,N_13338,N_13444);
xnor U13795 (N_13795,N_13044,N_13036);
nand U13796 (N_13796,N_12948,N_13078);
nor U13797 (N_13797,N_13409,N_12802);
xor U13798 (N_13798,N_13376,N_13318);
nor U13799 (N_13799,N_12947,N_13131);
or U13800 (N_13800,N_12794,N_13361);
xor U13801 (N_13801,N_13306,N_13210);
and U13802 (N_13802,N_13170,N_13236);
nand U13803 (N_13803,N_13296,N_13437);
nor U13804 (N_13804,N_12764,N_12873);
or U13805 (N_13805,N_13232,N_12784);
and U13806 (N_13806,N_13163,N_13424);
nand U13807 (N_13807,N_13416,N_13004);
or U13808 (N_13808,N_13261,N_12902);
nor U13809 (N_13809,N_13343,N_12863);
xor U13810 (N_13810,N_13202,N_13384);
and U13811 (N_13811,N_13097,N_13116);
and U13812 (N_13812,N_13240,N_13304);
or U13813 (N_13813,N_13265,N_13158);
nor U13814 (N_13814,N_13354,N_13380);
nand U13815 (N_13815,N_13046,N_12785);
nand U13816 (N_13816,N_13084,N_13324);
or U13817 (N_13817,N_13054,N_13074);
xor U13818 (N_13818,N_12804,N_13371);
xnor U13819 (N_13819,N_13237,N_13239);
nand U13820 (N_13820,N_12907,N_12879);
and U13821 (N_13821,N_12883,N_13329);
or U13822 (N_13822,N_13477,N_13187);
nor U13823 (N_13823,N_13412,N_13445);
and U13824 (N_13824,N_13478,N_13365);
and U13825 (N_13825,N_13176,N_13073);
or U13826 (N_13826,N_13034,N_12922);
xnor U13827 (N_13827,N_13226,N_13385);
or U13828 (N_13828,N_13252,N_13367);
xor U13829 (N_13829,N_12762,N_13315);
nand U13830 (N_13830,N_12993,N_13321);
or U13831 (N_13831,N_13212,N_13452);
and U13832 (N_13832,N_13128,N_13025);
nand U13833 (N_13833,N_13311,N_13038);
nand U13834 (N_13834,N_13497,N_13366);
nor U13835 (N_13835,N_13169,N_13112);
or U13836 (N_13836,N_13171,N_12955);
and U13837 (N_13837,N_13060,N_12850);
and U13838 (N_13838,N_13235,N_13209);
nor U13839 (N_13839,N_12914,N_13048);
nor U13840 (N_13840,N_12961,N_13175);
or U13841 (N_13841,N_12924,N_13333);
xor U13842 (N_13842,N_12848,N_12897);
or U13843 (N_13843,N_12871,N_13378);
or U13844 (N_13844,N_13133,N_13162);
and U13845 (N_13845,N_13488,N_13356);
xor U13846 (N_13846,N_13028,N_13313);
and U13847 (N_13847,N_12970,N_12787);
or U13848 (N_13848,N_12834,N_13438);
and U13849 (N_13849,N_12781,N_13206);
xor U13850 (N_13850,N_12801,N_13405);
or U13851 (N_13851,N_13407,N_12799);
nor U13852 (N_13852,N_12856,N_12771);
or U13853 (N_13853,N_13247,N_13195);
and U13854 (N_13854,N_12884,N_12767);
and U13855 (N_13855,N_13223,N_13083);
and U13856 (N_13856,N_13181,N_13087);
nand U13857 (N_13857,N_12876,N_13403);
or U13858 (N_13858,N_13013,N_12992);
and U13859 (N_13859,N_12750,N_13448);
and U13860 (N_13860,N_13045,N_13000);
or U13861 (N_13861,N_13140,N_12818);
and U13862 (N_13862,N_13059,N_13395);
nor U13863 (N_13863,N_12864,N_13109);
xor U13864 (N_13864,N_13238,N_13339);
and U13865 (N_13865,N_12894,N_13487);
nand U13866 (N_13866,N_12966,N_13068);
or U13867 (N_13867,N_13061,N_12967);
xor U13868 (N_13868,N_12772,N_13357);
nor U13869 (N_13869,N_13076,N_13132);
or U13870 (N_13870,N_12843,N_13454);
xor U13871 (N_13871,N_13427,N_13459);
nor U13872 (N_13872,N_13080,N_13359);
or U13873 (N_13873,N_13134,N_13093);
nand U13874 (N_13874,N_12890,N_13019);
and U13875 (N_13875,N_13106,N_12783);
and U13876 (N_13876,N_12918,N_13172);
xnor U13877 (N_13877,N_13368,N_13079);
nor U13878 (N_13878,N_12894,N_13110);
nand U13879 (N_13879,N_13227,N_13008);
nor U13880 (N_13880,N_13313,N_13172);
or U13881 (N_13881,N_13134,N_13002);
nand U13882 (N_13882,N_13448,N_13047);
xor U13883 (N_13883,N_13350,N_13094);
or U13884 (N_13884,N_13483,N_13095);
nor U13885 (N_13885,N_12886,N_12759);
xor U13886 (N_13886,N_12919,N_13304);
nand U13887 (N_13887,N_13429,N_13240);
and U13888 (N_13888,N_13199,N_13009);
or U13889 (N_13889,N_13153,N_13343);
nor U13890 (N_13890,N_13407,N_13297);
nand U13891 (N_13891,N_12970,N_12912);
and U13892 (N_13892,N_12919,N_13446);
xor U13893 (N_13893,N_13344,N_13074);
xnor U13894 (N_13894,N_13151,N_13130);
xor U13895 (N_13895,N_13278,N_13410);
or U13896 (N_13896,N_12845,N_13437);
nand U13897 (N_13897,N_12850,N_13012);
nand U13898 (N_13898,N_12929,N_13031);
and U13899 (N_13899,N_13257,N_13428);
and U13900 (N_13900,N_13316,N_13471);
and U13901 (N_13901,N_13168,N_13292);
xor U13902 (N_13902,N_13407,N_13179);
nand U13903 (N_13903,N_13327,N_12780);
or U13904 (N_13904,N_13475,N_12811);
nor U13905 (N_13905,N_13132,N_13470);
and U13906 (N_13906,N_12803,N_12970);
and U13907 (N_13907,N_13057,N_12776);
xnor U13908 (N_13908,N_13317,N_13391);
and U13909 (N_13909,N_13257,N_13351);
nand U13910 (N_13910,N_13484,N_12947);
or U13911 (N_13911,N_12865,N_13456);
nor U13912 (N_13912,N_12944,N_13278);
nand U13913 (N_13913,N_13079,N_12828);
nor U13914 (N_13914,N_13316,N_13158);
or U13915 (N_13915,N_13264,N_12826);
or U13916 (N_13916,N_13436,N_12975);
and U13917 (N_13917,N_13465,N_13323);
xnor U13918 (N_13918,N_13176,N_13248);
xor U13919 (N_13919,N_13224,N_13063);
nor U13920 (N_13920,N_12849,N_12871);
nand U13921 (N_13921,N_13472,N_13231);
xor U13922 (N_13922,N_12954,N_12824);
nand U13923 (N_13923,N_13153,N_12922);
or U13924 (N_13924,N_13239,N_12920);
xnor U13925 (N_13925,N_13406,N_13164);
xnor U13926 (N_13926,N_13147,N_12883);
nor U13927 (N_13927,N_13168,N_12831);
nand U13928 (N_13928,N_13122,N_13281);
nand U13929 (N_13929,N_12956,N_13041);
xnor U13930 (N_13930,N_13264,N_12922);
or U13931 (N_13931,N_13384,N_12843);
xnor U13932 (N_13932,N_13424,N_13253);
xor U13933 (N_13933,N_13110,N_13461);
or U13934 (N_13934,N_12865,N_12913);
xnor U13935 (N_13935,N_12978,N_12863);
xnor U13936 (N_13936,N_12765,N_13061);
nor U13937 (N_13937,N_13336,N_12834);
nand U13938 (N_13938,N_12857,N_13393);
nor U13939 (N_13939,N_12824,N_13445);
xor U13940 (N_13940,N_12922,N_13454);
xnor U13941 (N_13941,N_13011,N_13356);
or U13942 (N_13942,N_12959,N_13210);
or U13943 (N_13943,N_12924,N_13403);
nor U13944 (N_13944,N_13021,N_13467);
xor U13945 (N_13945,N_12917,N_12852);
nor U13946 (N_13946,N_13120,N_13069);
xnor U13947 (N_13947,N_12824,N_13080);
nand U13948 (N_13948,N_13461,N_13227);
xnor U13949 (N_13949,N_13185,N_13146);
nor U13950 (N_13950,N_12835,N_13446);
xnor U13951 (N_13951,N_12992,N_13139);
and U13952 (N_13952,N_13027,N_13495);
xnor U13953 (N_13953,N_13253,N_12864);
xor U13954 (N_13954,N_13139,N_13374);
or U13955 (N_13955,N_13312,N_12825);
nand U13956 (N_13956,N_13265,N_13471);
nor U13957 (N_13957,N_12892,N_13112);
xnor U13958 (N_13958,N_12834,N_12836);
nor U13959 (N_13959,N_13317,N_12884);
and U13960 (N_13960,N_13273,N_13103);
nand U13961 (N_13961,N_12764,N_13409);
nor U13962 (N_13962,N_13023,N_12888);
nor U13963 (N_13963,N_13435,N_13073);
nand U13964 (N_13964,N_13431,N_13443);
or U13965 (N_13965,N_13439,N_12931);
nand U13966 (N_13966,N_13206,N_12921);
xnor U13967 (N_13967,N_13412,N_13340);
nand U13968 (N_13968,N_13342,N_13199);
or U13969 (N_13969,N_13441,N_13488);
and U13970 (N_13970,N_12978,N_13257);
nand U13971 (N_13971,N_12777,N_13396);
nor U13972 (N_13972,N_13321,N_13000);
nor U13973 (N_13973,N_13231,N_12978);
nand U13974 (N_13974,N_13216,N_13391);
xor U13975 (N_13975,N_12862,N_12968);
nand U13976 (N_13976,N_13230,N_12929);
or U13977 (N_13977,N_13091,N_13396);
and U13978 (N_13978,N_13171,N_13483);
nand U13979 (N_13979,N_13034,N_13065);
or U13980 (N_13980,N_12967,N_12903);
nand U13981 (N_13981,N_12991,N_13061);
xnor U13982 (N_13982,N_13025,N_13455);
and U13983 (N_13983,N_12907,N_12928);
nor U13984 (N_13984,N_12824,N_13263);
nor U13985 (N_13985,N_13224,N_12929);
and U13986 (N_13986,N_13121,N_13284);
xor U13987 (N_13987,N_12828,N_13154);
nand U13988 (N_13988,N_12987,N_13264);
nor U13989 (N_13989,N_13101,N_13074);
xnor U13990 (N_13990,N_12787,N_13473);
and U13991 (N_13991,N_12987,N_13209);
and U13992 (N_13992,N_13275,N_13098);
and U13993 (N_13993,N_13232,N_13467);
or U13994 (N_13994,N_13309,N_12911);
or U13995 (N_13995,N_13206,N_12987);
xor U13996 (N_13996,N_13366,N_12795);
and U13997 (N_13997,N_13478,N_13086);
or U13998 (N_13998,N_13471,N_13226);
xnor U13999 (N_13999,N_12823,N_13301);
nor U14000 (N_14000,N_13217,N_13224);
or U14001 (N_14001,N_13190,N_13152);
nand U14002 (N_14002,N_12866,N_12922);
or U14003 (N_14003,N_13425,N_13141);
and U14004 (N_14004,N_13398,N_13193);
or U14005 (N_14005,N_12873,N_13039);
and U14006 (N_14006,N_12972,N_13356);
nor U14007 (N_14007,N_13360,N_13447);
and U14008 (N_14008,N_13252,N_13030);
xnor U14009 (N_14009,N_13090,N_12879);
or U14010 (N_14010,N_13471,N_12997);
xor U14011 (N_14011,N_13306,N_12985);
nand U14012 (N_14012,N_13300,N_12958);
or U14013 (N_14013,N_13377,N_13045);
xnor U14014 (N_14014,N_13250,N_13121);
and U14015 (N_14015,N_13262,N_12784);
nand U14016 (N_14016,N_12870,N_13414);
or U14017 (N_14017,N_13110,N_12892);
nand U14018 (N_14018,N_12939,N_12855);
nor U14019 (N_14019,N_13233,N_13366);
and U14020 (N_14020,N_12774,N_13292);
xor U14021 (N_14021,N_13150,N_13010);
xor U14022 (N_14022,N_13114,N_13356);
xor U14023 (N_14023,N_13100,N_13466);
nand U14024 (N_14024,N_13161,N_13290);
xnor U14025 (N_14025,N_13319,N_13019);
nor U14026 (N_14026,N_13382,N_13212);
xnor U14027 (N_14027,N_13148,N_13103);
or U14028 (N_14028,N_12962,N_12973);
or U14029 (N_14029,N_12804,N_13418);
xor U14030 (N_14030,N_13363,N_12905);
and U14031 (N_14031,N_13262,N_13074);
or U14032 (N_14032,N_13064,N_13428);
or U14033 (N_14033,N_13435,N_13404);
and U14034 (N_14034,N_12984,N_13355);
xor U14035 (N_14035,N_12779,N_13403);
or U14036 (N_14036,N_13476,N_13078);
nand U14037 (N_14037,N_13188,N_12783);
or U14038 (N_14038,N_13373,N_13456);
nand U14039 (N_14039,N_13146,N_13103);
xnor U14040 (N_14040,N_12859,N_13177);
xnor U14041 (N_14041,N_12876,N_12994);
xnor U14042 (N_14042,N_13016,N_13192);
and U14043 (N_14043,N_13111,N_12972);
xnor U14044 (N_14044,N_13385,N_13459);
xnor U14045 (N_14045,N_12886,N_12889);
nand U14046 (N_14046,N_13395,N_12897);
and U14047 (N_14047,N_13424,N_13154);
or U14048 (N_14048,N_12795,N_12966);
nand U14049 (N_14049,N_13341,N_12777);
and U14050 (N_14050,N_13308,N_12968);
and U14051 (N_14051,N_13003,N_13328);
xor U14052 (N_14052,N_13232,N_13247);
nor U14053 (N_14053,N_13325,N_13305);
xor U14054 (N_14054,N_13495,N_13435);
or U14055 (N_14055,N_12868,N_12989);
nand U14056 (N_14056,N_13014,N_13001);
nand U14057 (N_14057,N_13107,N_13160);
and U14058 (N_14058,N_13279,N_13410);
xnor U14059 (N_14059,N_13202,N_12822);
nor U14060 (N_14060,N_12975,N_13108);
nor U14061 (N_14061,N_12754,N_12985);
xor U14062 (N_14062,N_13140,N_13380);
xnor U14063 (N_14063,N_13120,N_13452);
xor U14064 (N_14064,N_12780,N_13367);
nand U14065 (N_14065,N_13167,N_13322);
nor U14066 (N_14066,N_13233,N_13408);
nand U14067 (N_14067,N_12967,N_13227);
xor U14068 (N_14068,N_12915,N_13014);
or U14069 (N_14069,N_13357,N_13419);
nand U14070 (N_14070,N_13320,N_13476);
nor U14071 (N_14071,N_13129,N_12849);
or U14072 (N_14072,N_12999,N_13259);
xor U14073 (N_14073,N_13055,N_13443);
xor U14074 (N_14074,N_12976,N_12891);
nand U14075 (N_14075,N_13468,N_12907);
or U14076 (N_14076,N_13348,N_12789);
or U14077 (N_14077,N_13138,N_13158);
xnor U14078 (N_14078,N_13234,N_12834);
and U14079 (N_14079,N_13426,N_13442);
or U14080 (N_14080,N_13263,N_13472);
or U14081 (N_14081,N_13316,N_13095);
or U14082 (N_14082,N_13445,N_13491);
or U14083 (N_14083,N_13103,N_12809);
nor U14084 (N_14084,N_13035,N_13483);
and U14085 (N_14085,N_12884,N_13102);
or U14086 (N_14086,N_13135,N_12944);
or U14087 (N_14087,N_12849,N_12822);
xor U14088 (N_14088,N_13092,N_13122);
and U14089 (N_14089,N_12848,N_13398);
or U14090 (N_14090,N_12977,N_13480);
xor U14091 (N_14091,N_13314,N_12796);
xnor U14092 (N_14092,N_13286,N_12839);
and U14093 (N_14093,N_13029,N_13148);
or U14094 (N_14094,N_12882,N_13283);
nor U14095 (N_14095,N_12967,N_13047);
or U14096 (N_14096,N_13206,N_12977);
or U14097 (N_14097,N_13094,N_13171);
or U14098 (N_14098,N_12761,N_13375);
nand U14099 (N_14099,N_13385,N_12879);
and U14100 (N_14100,N_13227,N_13232);
and U14101 (N_14101,N_12752,N_13062);
or U14102 (N_14102,N_13492,N_13326);
nand U14103 (N_14103,N_12814,N_12855);
and U14104 (N_14104,N_13324,N_13222);
and U14105 (N_14105,N_12939,N_12771);
and U14106 (N_14106,N_12985,N_13076);
nor U14107 (N_14107,N_13464,N_13475);
and U14108 (N_14108,N_12787,N_13004);
nand U14109 (N_14109,N_12974,N_12913);
xor U14110 (N_14110,N_13375,N_13289);
and U14111 (N_14111,N_12810,N_12890);
nand U14112 (N_14112,N_13033,N_13301);
nor U14113 (N_14113,N_12754,N_13262);
xnor U14114 (N_14114,N_13181,N_12848);
nand U14115 (N_14115,N_13154,N_13179);
or U14116 (N_14116,N_13322,N_13497);
and U14117 (N_14117,N_13036,N_12978);
and U14118 (N_14118,N_13246,N_13320);
or U14119 (N_14119,N_12844,N_13070);
and U14120 (N_14120,N_13088,N_13084);
or U14121 (N_14121,N_13189,N_12943);
xnor U14122 (N_14122,N_13134,N_13205);
xnor U14123 (N_14123,N_13191,N_12882);
and U14124 (N_14124,N_12770,N_12828);
and U14125 (N_14125,N_12915,N_12939);
nor U14126 (N_14126,N_12801,N_13325);
and U14127 (N_14127,N_13489,N_12865);
xnor U14128 (N_14128,N_13493,N_13433);
nand U14129 (N_14129,N_13341,N_13495);
or U14130 (N_14130,N_13377,N_13439);
nand U14131 (N_14131,N_13481,N_12765);
xnor U14132 (N_14132,N_13491,N_13159);
xnor U14133 (N_14133,N_13096,N_13499);
xor U14134 (N_14134,N_13216,N_13276);
xor U14135 (N_14135,N_13421,N_13179);
xnor U14136 (N_14136,N_13000,N_13224);
nor U14137 (N_14137,N_12801,N_12985);
or U14138 (N_14138,N_12973,N_13090);
and U14139 (N_14139,N_13491,N_12828);
nor U14140 (N_14140,N_12821,N_13163);
and U14141 (N_14141,N_13041,N_13059);
and U14142 (N_14142,N_13479,N_12753);
and U14143 (N_14143,N_12992,N_13015);
or U14144 (N_14144,N_13057,N_13015);
and U14145 (N_14145,N_13071,N_13243);
nand U14146 (N_14146,N_12838,N_13210);
nor U14147 (N_14147,N_12794,N_13484);
nor U14148 (N_14148,N_13001,N_13422);
nor U14149 (N_14149,N_13060,N_13175);
and U14150 (N_14150,N_12791,N_13089);
xnor U14151 (N_14151,N_13482,N_13265);
nand U14152 (N_14152,N_13318,N_13176);
nor U14153 (N_14153,N_13128,N_13483);
and U14154 (N_14154,N_13221,N_13250);
or U14155 (N_14155,N_13073,N_13175);
nand U14156 (N_14156,N_13192,N_13083);
or U14157 (N_14157,N_13321,N_12778);
nor U14158 (N_14158,N_13000,N_12798);
xor U14159 (N_14159,N_13237,N_12975);
and U14160 (N_14160,N_13208,N_13480);
nor U14161 (N_14161,N_13166,N_13050);
xor U14162 (N_14162,N_13278,N_13215);
and U14163 (N_14163,N_12918,N_13395);
nor U14164 (N_14164,N_12822,N_13495);
xor U14165 (N_14165,N_12763,N_13489);
or U14166 (N_14166,N_12952,N_12951);
or U14167 (N_14167,N_13365,N_12872);
xnor U14168 (N_14168,N_13336,N_12955);
and U14169 (N_14169,N_13247,N_13464);
nor U14170 (N_14170,N_12930,N_13228);
xnor U14171 (N_14171,N_13281,N_13476);
nand U14172 (N_14172,N_13368,N_13155);
nand U14173 (N_14173,N_12884,N_13187);
xor U14174 (N_14174,N_13137,N_12756);
nor U14175 (N_14175,N_13424,N_12897);
xor U14176 (N_14176,N_12907,N_13357);
xnor U14177 (N_14177,N_13179,N_12898);
xnor U14178 (N_14178,N_13175,N_13013);
nor U14179 (N_14179,N_13012,N_13128);
nor U14180 (N_14180,N_13253,N_13272);
and U14181 (N_14181,N_12825,N_13478);
nand U14182 (N_14182,N_13161,N_13160);
or U14183 (N_14183,N_13160,N_13129);
and U14184 (N_14184,N_13151,N_13210);
and U14185 (N_14185,N_12861,N_12942);
or U14186 (N_14186,N_13154,N_13481);
and U14187 (N_14187,N_13239,N_13265);
nor U14188 (N_14188,N_13253,N_12764);
or U14189 (N_14189,N_12798,N_12909);
xor U14190 (N_14190,N_13491,N_12939);
nor U14191 (N_14191,N_13448,N_13131);
and U14192 (N_14192,N_12973,N_12886);
nor U14193 (N_14193,N_13322,N_13418);
and U14194 (N_14194,N_12804,N_13489);
nand U14195 (N_14195,N_13155,N_12761);
nor U14196 (N_14196,N_13192,N_13193);
or U14197 (N_14197,N_12883,N_12969);
xor U14198 (N_14198,N_13053,N_13476);
or U14199 (N_14199,N_13498,N_13164);
xnor U14200 (N_14200,N_13371,N_12880);
nor U14201 (N_14201,N_12863,N_13368);
or U14202 (N_14202,N_13481,N_13345);
nand U14203 (N_14203,N_13292,N_13285);
and U14204 (N_14204,N_13133,N_13060);
xnor U14205 (N_14205,N_13377,N_12972);
and U14206 (N_14206,N_13343,N_13436);
and U14207 (N_14207,N_13388,N_13486);
xor U14208 (N_14208,N_13233,N_12859);
or U14209 (N_14209,N_13426,N_13187);
xor U14210 (N_14210,N_12870,N_13208);
nor U14211 (N_14211,N_13102,N_12761);
nand U14212 (N_14212,N_13099,N_13332);
nor U14213 (N_14213,N_12750,N_13195);
nor U14214 (N_14214,N_13007,N_12774);
nor U14215 (N_14215,N_13147,N_12995);
and U14216 (N_14216,N_12832,N_13288);
xnor U14217 (N_14217,N_13326,N_12854);
xnor U14218 (N_14218,N_13473,N_13180);
nand U14219 (N_14219,N_13142,N_13397);
nor U14220 (N_14220,N_13136,N_13215);
xnor U14221 (N_14221,N_13149,N_12942);
nand U14222 (N_14222,N_13434,N_13006);
nor U14223 (N_14223,N_13055,N_13007);
nor U14224 (N_14224,N_13342,N_12863);
nor U14225 (N_14225,N_13327,N_12792);
nor U14226 (N_14226,N_13223,N_13009);
nor U14227 (N_14227,N_12881,N_13035);
nand U14228 (N_14228,N_13466,N_12796);
or U14229 (N_14229,N_13478,N_12829);
and U14230 (N_14230,N_12778,N_12924);
or U14231 (N_14231,N_12822,N_12772);
and U14232 (N_14232,N_13482,N_13042);
nor U14233 (N_14233,N_12845,N_12959);
nor U14234 (N_14234,N_12884,N_13342);
xor U14235 (N_14235,N_13113,N_13242);
nor U14236 (N_14236,N_13252,N_12752);
and U14237 (N_14237,N_13285,N_12970);
xor U14238 (N_14238,N_12944,N_13330);
and U14239 (N_14239,N_13252,N_13282);
and U14240 (N_14240,N_13024,N_13180);
or U14241 (N_14241,N_13031,N_13471);
and U14242 (N_14242,N_13225,N_13279);
xor U14243 (N_14243,N_13450,N_13159);
nand U14244 (N_14244,N_12993,N_13239);
nor U14245 (N_14245,N_12751,N_13453);
xor U14246 (N_14246,N_13432,N_13213);
nand U14247 (N_14247,N_12945,N_13365);
xnor U14248 (N_14248,N_13481,N_13299);
xor U14249 (N_14249,N_12805,N_12915);
nor U14250 (N_14250,N_13566,N_13959);
xnor U14251 (N_14251,N_13558,N_13816);
xnor U14252 (N_14252,N_14191,N_13638);
nand U14253 (N_14253,N_14056,N_14164);
nand U14254 (N_14254,N_14016,N_13739);
xor U14255 (N_14255,N_13673,N_13832);
nand U14256 (N_14256,N_14059,N_13946);
or U14257 (N_14257,N_13622,N_14020);
or U14258 (N_14258,N_13679,N_14000);
xnor U14259 (N_14259,N_14105,N_14229);
xor U14260 (N_14260,N_13817,N_13740);
nor U14261 (N_14261,N_13874,N_14092);
xor U14262 (N_14262,N_13981,N_13974);
xnor U14263 (N_14263,N_13624,N_13991);
nor U14264 (N_14264,N_14017,N_13630);
nand U14265 (N_14265,N_13797,N_14209);
nand U14266 (N_14266,N_14051,N_13831);
and U14267 (N_14267,N_14176,N_13579);
or U14268 (N_14268,N_13815,N_14024);
and U14269 (N_14269,N_14023,N_13954);
or U14270 (N_14270,N_13888,N_14230);
nand U14271 (N_14271,N_13572,N_13507);
nand U14272 (N_14272,N_13601,N_13556);
or U14273 (N_14273,N_13890,N_13899);
or U14274 (N_14274,N_14211,N_14037);
or U14275 (N_14275,N_13736,N_13654);
and U14276 (N_14276,N_13957,N_14066);
nor U14277 (N_14277,N_13674,N_13509);
xor U14278 (N_14278,N_13830,N_13903);
nand U14279 (N_14279,N_13933,N_13748);
nor U14280 (N_14280,N_13966,N_13887);
xnor U14281 (N_14281,N_13685,N_14188);
or U14282 (N_14282,N_13517,N_13500);
and U14283 (N_14283,N_13828,N_13606);
or U14284 (N_14284,N_13620,N_13561);
nand U14285 (N_14285,N_13574,N_13687);
or U14286 (N_14286,N_13709,N_13503);
nand U14287 (N_14287,N_13531,N_13608);
xnor U14288 (N_14288,N_13690,N_13875);
or U14289 (N_14289,N_13548,N_13914);
and U14290 (N_14290,N_13962,N_14005);
nand U14291 (N_14291,N_13502,N_13861);
nand U14292 (N_14292,N_14027,N_14062);
nor U14293 (N_14293,N_14243,N_13523);
or U14294 (N_14294,N_13961,N_14232);
xor U14295 (N_14295,N_13824,N_13636);
or U14296 (N_14296,N_13960,N_13650);
nand U14297 (N_14297,N_13508,N_13879);
nand U14298 (N_14298,N_13759,N_13807);
nor U14299 (N_14299,N_13805,N_13818);
xor U14300 (N_14300,N_13973,N_14126);
or U14301 (N_14301,N_14123,N_13592);
and U14302 (N_14302,N_13617,N_13868);
and U14303 (N_14303,N_14124,N_13684);
xor U14304 (N_14304,N_13677,N_13696);
and U14305 (N_14305,N_14200,N_13920);
or U14306 (N_14306,N_13651,N_14151);
nor U14307 (N_14307,N_13848,N_14057);
or U14308 (N_14308,N_13589,N_14085);
and U14309 (N_14309,N_14247,N_14028);
or U14310 (N_14310,N_13770,N_13796);
nor U14311 (N_14311,N_13999,N_13757);
or U14312 (N_14312,N_14179,N_14212);
and U14313 (N_14313,N_13747,N_13664);
xor U14314 (N_14314,N_13794,N_13778);
xnor U14315 (N_14315,N_14014,N_13814);
nor U14316 (N_14316,N_13541,N_13937);
or U14317 (N_14317,N_13777,N_13542);
or U14318 (N_14318,N_14128,N_14141);
and U14319 (N_14319,N_14181,N_14069);
nand U14320 (N_14320,N_13925,N_13774);
nor U14321 (N_14321,N_13915,N_13595);
nand U14322 (N_14322,N_13922,N_13626);
or U14323 (N_14323,N_13604,N_14204);
nand U14324 (N_14324,N_13825,N_14030);
xnor U14325 (N_14325,N_14121,N_14127);
and U14326 (N_14326,N_13569,N_13993);
xor U14327 (N_14327,N_13853,N_14091);
nor U14328 (N_14328,N_13940,N_14042);
and U14329 (N_14329,N_14155,N_13844);
and U14330 (N_14330,N_14072,N_13893);
xor U14331 (N_14331,N_14180,N_13938);
and U14332 (N_14332,N_14118,N_14029);
nand U14333 (N_14333,N_14008,N_13694);
and U14334 (N_14334,N_14087,N_13667);
nand U14335 (N_14335,N_13970,N_13886);
and U14336 (N_14336,N_14183,N_13926);
or U14337 (N_14337,N_13640,N_14142);
nor U14338 (N_14338,N_13733,N_13917);
nor U14339 (N_14339,N_14018,N_13958);
xnor U14340 (N_14340,N_13758,N_14046);
nor U14341 (N_14341,N_14048,N_14224);
xor U14342 (N_14342,N_14119,N_13826);
nor U14343 (N_14343,N_13929,N_13632);
nand U14344 (N_14344,N_13905,N_14113);
or U14345 (N_14345,N_13785,N_14074);
xnor U14346 (N_14346,N_14114,N_13851);
xnor U14347 (N_14347,N_14090,N_13704);
xnor U14348 (N_14348,N_14136,N_13633);
nor U14349 (N_14349,N_13554,N_13935);
nor U14350 (N_14350,N_14182,N_13551);
nor U14351 (N_14351,N_13896,N_13615);
or U14352 (N_14352,N_13819,N_13560);
and U14353 (N_14353,N_14089,N_13707);
xnor U14354 (N_14354,N_14117,N_14001);
and U14355 (N_14355,N_13616,N_14153);
or U14356 (N_14356,N_13901,N_13878);
nand U14357 (N_14357,N_13576,N_13977);
nor U14358 (N_14358,N_14236,N_13555);
nor U14359 (N_14359,N_13725,N_13869);
and U14360 (N_14360,N_13575,N_13994);
nand U14361 (N_14361,N_13522,N_14055);
or U14362 (N_14362,N_14221,N_13742);
xor U14363 (N_14363,N_13990,N_13543);
xnor U14364 (N_14364,N_13989,N_13649);
nor U14365 (N_14365,N_13688,N_13600);
nor U14366 (N_14366,N_14079,N_14120);
or U14367 (N_14367,N_14190,N_14194);
nand U14368 (N_14368,N_13978,N_13516);
and U14369 (N_14369,N_13867,N_13565);
xor U14370 (N_14370,N_14208,N_13609);
or U14371 (N_14371,N_14013,N_14039);
or U14372 (N_14372,N_13773,N_13614);
or U14373 (N_14373,N_13505,N_13941);
xnor U14374 (N_14374,N_13792,N_13950);
xnor U14375 (N_14375,N_13806,N_13699);
and U14376 (N_14376,N_13676,N_14009);
xnor U14377 (N_14377,N_13908,N_13968);
nor U14378 (N_14378,N_13672,N_13976);
nand U14379 (N_14379,N_13822,N_14060);
or U14380 (N_14380,N_14148,N_13501);
nand U14381 (N_14381,N_13544,N_13618);
and U14382 (N_14382,N_14154,N_13741);
nand U14383 (N_14383,N_13997,N_13812);
nand U14384 (N_14384,N_13534,N_13919);
nand U14385 (N_14385,N_13971,N_14094);
xnor U14386 (N_14386,N_14096,N_14196);
nand U14387 (N_14387,N_13536,N_13652);
nand U14388 (N_14388,N_14054,N_13889);
nand U14389 (N_14389,N_13563,N_14082);
or U14390 (N_14390,N_13708,N_13979);
nand U14391 (N_14391,N_13537,N_13559);
xor U14392 (N_14392,N_13882,N_13586);
xnor U14393 (N_14393,N_13698,N_13921);
nor U14394 (N_14394,N_14184,N_13755);
or U14395 (N_14395,N_14093,N_14244);
xnor U14396 (N_14396,N_13634,N_14246);
nor U14397 (N_14397,N_13644,N_13891);
and U14398 (N_14398,N_13827,N_14203);
and U14399 (N_14399,N_13945,N_13530);
and U14400 (N_14400,N_13539,N_14041);
xnor U14401 (N_14401,N_13573,N_13710);
xnor U14402 (N_14402,N_14097,N_13843);
or U14403 (N_14403,N_14234,N_14088);
xnor U14404 (N_14404,N_13720,N_13647);
or U14405 (N_14405,N_13716,N_13728);
and U14406 (N_14406,N_13602,N_13907);
and U14407 (N_14407,N_13860,N_13801);
or U14408 (N_14408,N_14077,N_13847);
and U14409 (N_14409,N_14165,N_13553);
or U14410 (N_14410,N_13972,N_14162);
or U14411 (N_14411,N_13768,N_13924);
or U14412 (N_14412,N_14242,N_13852);
and U14413 (N_14413,N_14132,N_14135);
nand U14414 (N_14414,N_14158,N_14193);
nor U14415 (N_14415,N_13823,N_13700);
and U14416 (N_14416,N_13939,N_14167);
or U14417 (N_14417,N_13841,N_14207);
and U14418 (N_14418,N_14248,N_13686);
xnor U14419 (N_14419,N_14219,N_13656);
and U14420 (N_14420,N_13766,N_14226);
or U14421 (N_14421,N_13749,N_13964);
nor U14422 (N_14422,N_13776,N_13745);
xor U14423 (N_14423,N_13629,N_14107);
xor U14424 (N_14424,N_13913,N_13786);
xor U14425 (N_14425,N_14171,N_13675);
xor U14426 (N_14426,N_13975,N_14173);
nor U14427 (N_14427,N_13857,N_13625);
xor U14428 (N_14428,N_13721,N_13809);
xnor U14429 (N_14429,N_14061,N_13948);
nor U14430 (N_14430,N_14198,N_14239);
or U14431 (N_14431,N_13840,N_13582);
xnor U14432 (N_14432,N_13528,N_13884);
nand U14433 (N_14433,N_13876,N_14220);
or U14434 (N_14434,N_13692,N_14241);
nand U14435 (N_14435,N_13691,N_14098);
and U14436 (N_14436,N_14021,N_14227);
xnor U14437 (N_14437,N_13779,N_13932);
nor U14438 (N_14438,N_14011,N_14063);
nor U14439 (N_14439,N_13538,N_13859);
xor U14440 (N_14440,N_14228,N_13750);
or U14441 (N_14441,N_14245,N_13943);
nor U14442 (N_14442,N_14073,N_13682);
and U14443 (N_14443,N_13872,N_13506);
xor U14444 (N_14444,N_13969,N_14214);
nand U14445 (N_14445,N_14007,N_13552);
xnor U14446 (N_14446,N_13645,N_13525);
nor U14447 (N_14447,N_13599,N_14215);
nand U14448 (N_14448,N_13845,N_13753);
and U14449 (N_14449,N_14022,N_13655);
nand U14450 (N_14450,N_14110,N_14015);
nand U14451 (N_14451,N_13570,N_13928);
or U14452 (N_14452,N_13646,N_13562);
nand U14453 (N_14453,N_13722,N_14177);
nand U14454 (N_14454,N_13787,N_14139);
or U14455 (N_14455,N_13767,N_13577);
or U14456 (N_14456,N_13963,N_14064);
nand U14457 (N_14457,N_13607,N_13892);
and U14458 (N_14458,N_13871,N_13810);
nand U14459 (N_14459,N_13947,N_14010);
xor U14460 (N_14460,N_13723,N_13870);
xnor U14461 (N_14461,N_14157,N_14160);
xnor U14462 (N_14462,N_13992,N_14086);
nand U14463 (N_14463,N_13578,N_13836);
and U14464 (N_14464,N_14033,N_13695);
nor U14465 (N_14465,N_13714,N_13762);
or U14466 (N_14466,N_13746,N_13628);
and U14467 (N_14467,N_13521,N_13858);
nor U14468 (N_14468,N_14003,N_14159);
xor U14469 (N_14469,N_14161,N_13621);
and U14470 (N_14470,N_13631,N_13862);
and U14471 (N_14471,N_14144,N_13916);
nor U14472 (N_14472,N_14216,N_13581);
and U14473 (N_14473,N_14076,N_13658);
nor U14474 (N_14474,N_13951,N_14031);
or U14475 (N_14475,N_13511,N_14099);
or U14476 (N_14476,N_14134,N_14233);
or U14477 (N_14477,N_13513,N_14125);
nand U14478 (N_14478,N_13846,N_14217);
xor U14479 (N_14479,N_13729,N_13590);
nor U14480 (N_14480,N_13838,N_14104);
nand U14481 (N_14481,N_13895,N_13769);
or U14482 (N_14482,N_13781,N_13930);
and U14483 (N_14483,N_14240,N_13744);
and U14484 (N_14484,N_13789,N_14034);
or U14485 (N_14485,N_13512,N_13584);
nand U14486 (N_14486,N_14108,N_14019);
nand U14487 (N_14487,N_14084,N_13980);
or U14488 (N_14488,N_13603,N_13567);
nand U14489 (N_14489,N_13995,N_14035);
xnor U14490 (N_14490,N_13751,N_13591);
nor U14491 (N_14491,N_13705,N_13661);
nor U14492 (N_14492,N_13952,N_13526);
or U14493 (N_14493,N_14249,N_14111);
xnor U14494 (N_14494,N_13648,N_13585);
nand U14495 (N_14495,N_13670,N_13835);
nand U14496 (N_14496,N_14213,N_13571);
nand U14497 (N_14497,N_14202,N_14185);
or U14498 (N_14498,N_13524,N_13983);
or U14499 (N_14499,N_13518,N_13985);
or U14500 (N_14500,N_14145,N_14053);
nand U14501 (N_14501,N_14186,N_13965);
nand U14502 (N_14502,N_13550,N_13911);
or U14503 (N_14503,N_13760,N_13732);
xnor U14504 (N_14504,N_13927,N_14235);
or U14505 (N_14505,N_13623,N_13735);
nand U14506 (N_14506,N_13904,N_13738);
or U14507 (N_14507,N_14174,N_13934);
or U14508 (N_14508,N_13715,N_13906);
and U14509 (N_14509,N_13529,N_13821);
nand U14510 (N_14510,N_13653,N_13793);
and U14511 (N_14511,N_13663,N_13597);
nand U14512 (N_14512,N_13545,N_13701);
xnor U14513 (N_14513,N_13535,N_14080);
xor U14514 (N_14514,N_13737,N_13880);
and U14515 (N_14515,N_13942,N_13568);
nor U14516 (N_14516,N_14223,N_14137);
or U14517 (N_14517,N_13804,N_14065);
and U14518 (N_14518,N_13829,N_13593);
xor U14519 (N_14519,N_14058,N_14050);
nor U14520 (N_14520,N_13894,N_13706);
and U14521 (N_14521,N_13772,N_14101);
and U14522 (N_14522,N_14036,N_14070);
and U14523 (N_14523,N_13956,N_13923);
or U14524 (N_14524,N_13689,N_13743);
or U14525 (N_14525,N_14081,N_13811);
nand U14526 (N_14526,N_13849,N_14040);
nand U14527 (N_14527,N_13864,N_13885);
nand U14528 (N_14528,N_14140,N_13863);
or U14529 (N_14529,N_14044,N_14143);
nor U14530 (N_14530,N_13866,N_13782);
or U14531 (N_14531,N_14047,N_14131);
xnor U14532 (N_14532,N_13795,N_14049);
or U14533 (N_14533,N_13788,N_13660);
or U14534 (N_14534,N_14197,N_13842);
xnor U14535 (N_14535,N_14149,N_13662);
nor U14536 (N_14536,N_14002,N_13987);
xnor U14537 (N_14537,N_13909,N_13612);
and U14538 (N_14538,N_13703,N_13659);
or U14539 (N_14539,N_13873,N_14163);
xnor U14540 (N_14540,N_13900,N_14170);
and U14541 (N_14541,N_14147,N_13883);
xor U14542 (N_14542,N_13754,N_14201);
and U14543 (N_14543,N_14195,N_14205);
nand U14544 (N_14544,N_14178,N_13711);
and U14545 (N_14545,N_13726,N_13763);
xor U14546 (N_14546,N_13641,N_14192);
nor U14547 (N_14547,N_13731,N_14032);
and U14548 (N_14548,N_14115,N_13955);
or U14549 (N_14549,N_13802,N_13588);
and U14550 (N_14550,N_13799,N_13771);
xor U14551 (N_14551,N_13504,N_14109);
xnor U14552 (N_14552,N_14199,N_13697);
nand U14553 (N_14553,N_14025,N_13519);
or U14554 (N_14554,N_14075,N_13637);
or U14555 (N_14555,N_14172,N_13761);
nor U14556 (N_14556,N_14006,N_13800);
nor U14557 (N_14557,N_13587,N_14100);
xor U14558 (N_14558,N_14038,N_13520);
nand U14559 (N_14559,N_13533,N_13657);
or U14560 (N_14560,N_14106,N_14146);
nand U14561 (N_14561,N_13752,N_13865);
and U14562 (N_14562,N_13912,N_13627);
nand U14563 (N_14563,N_13730,N_14102);
and U14564 (N_14564,N_13635,N_13798);
xnor U14565 (N_14565,N_14133,N_13727);
nand U14566 (N_14566,N_13510,N_13967);
xor U14567 (N_14567,N_13944,N_13918);
nand U14568 (N_14568,N_14103,N_13718);
nor U14569 (N_14569,N_13639,N_13557);
xor U14570 (N_14570,N_13693,N_14130);
or U14571 (N_14571,N_13514,N_13642);
or U14572 (N_14572,N_13953,N_13936);
xnor U14573 (N_14573,N_13619,N_13702);
or U14574 (N_14574,N_14004,N_13820);
xnor U14575 (N_14575,N_14067,N_13666);
or U14576 (N_14576,N_13643,N_13610);
nor U14577 (N_14577,N_13765,N_13680);
or U14578 (N_14578,N_13515,N_13813);
or U14579 (N_14579,N_13540,N_13668);
nor U14580 (N_14580,N_13596,N_14138);
xor U14581 (N_14581,N_13605,N_14166);
or U14582 (N_14582,N_13877,N_13583);
or U14583 (N_14583,N_13764,N_14112);
and U14584 (N_14584,N_13665,N_13756);
xnor U14585 (N_14585,N_14210,N_13681);
or U14586 (N_14586,N_14129,N_13855);
nand U14587 (N_14587,N_14225,N_13910);
nand U14588 (N_14588,N_13784,N_14237);
or U14589 (N_14589,N_14222,N_13898);
or U14590 (N_14590,N_14083,N_14238);
nor U14591 (N_14591,N_13717,N_13881);
nor U14592 (N_14592,N_13594,N_13897);
nor U14593 (N_14593,N_13532,N_13931);
or U14594 (N_14594,N_13683,N_13850);
and U14595 (N_14595,N_13549,N_13986);
nand U14596 (N_14596,N_13724,N_13803);
or U14597 (N_14597,N_14045,N_14012);
and U14598 (N_14598,N_13837,N_14078);
xor U14599 (N_14599,N_13834,N_13854);
or U14600 (N_14600,N_13713,N_13808);
or U14601 (N_14601,N_13839,N_13791);
or U14602 (N_14602,N_13671,N_14052);
xor U14603 (N_14603,N_13982,N_14150);
nand U14604 (N_14604,N_13984,N_14175);
nor U14605 (N_14605,N_13856,N_14168);
nand U14606 (N_14606,N_13783,N_14068);
xor U14607 (N_14607,N_13564,N_13902);
xnor U14608 (N_14608,N_14043,N_14206);
or U14609 (N_14609,N_13712,N_14071);
nor U14610 (N_14610,N_14187,N_13775);
and U14611 (N_14611,N_14026,N_13598);
and U14612 (N_14612,N_14116,N_13998);
nor U14613 (N_14613,N_13580,N_13546);
and U14614 (N_14614,N_13719,N_14152);
or U14615 (N_14615,N_13988,N_13949);
xor U14616 (N_14616,N_14095,N_14231);
or U14617 (N_14617,N_14189,N_14169);
and U14618 (N_14618,N_13527,N_14122);
nor U14619 (N_14619,N_13547,N_14156);
nor U14620 (N_14620,N_13833,N_13790);
and U14621 (N_14621,N_13669,N_14218);
xor U14622 (N_14622,N_13613,N_13734);
xnor U14623 (N_14623,N_13678,N_13996);
xnor U14624 (N_14624,N_13611,N_13780);
and U14625 (N_14625,N_13592,N_13909);
nor U14626 (N_14626,N_13531,N_14138);
nand U14627 (N_14627,N_14160,N_14174);
nor U14628 (N_14628,N_14095,N_13558);
xnor U14629 (N_14629,N_13958,N_14091);
nor U14630 (N_14630,N_13649,N_13985);
nand U14631 (N_14631,N_13647,N_13533);
nor U14632 (N_14632,N_13517,N_13926);
nor U14633 (N_14633,N_13975,N_14004);
nand U14634 (N_14634,N_14181,N_14109);
or U14635 (N_14635,N_13582,N_13527);
xor U14636 (N_14636,N_14056,N_13508);
nor U14637 (N_14637,N_13872,N_14140);
and U14638 (N_14638,N_13816,N_13852);
and U14639 (N_14639,N_13507,N_14226);
nand U14640 (N_14640,N_14102,N_14238);
nor U14641 (N_14641,N_14201,N_14073);
nand U14642 (N_14642,N_14220,N_13513);
nor U14643 (N_14643,N_13877,N_13655);
nor U14644 (N_14644,N_13965,N_14181);
xnor U14645 (N_14645,N_13524,N_13505);
or U14646 (N_14646,N_14120,N_13551);
xnor U14647 (N_14647,N_13944,N_13934);
and U14648 (N_14648,N_13806,N_14092);
and U14649 (N_14649,N_13633,N_13646);
nand U14650 (N_14650,N_14181,N_13768);
or U14651 (N_14651,N_13600,N_13554);
and U14652 (N_14652,N_14115,N_13632);
or U14653 (N_14653,N_14032,N_14040);
nand U14654 (N_14654,N_13626,N_13629);
nor U14655 (N_14655,N_13700,N_13719);
and U14656 (N_14656,N_14023,N_13931);
nor U14657 (N_14657,N_14028,N_13690);
nand U14658 (N_14658,N_13845,N_14084);
nand U14659 (N_14659,N_13575,N_13741);
xor U14660 (N_14660,N_14178,N_14045);
and U14661 (N_14661,N_13736,N_13820);
nand U14662 (N_14662,N_14151,N_13506);
and U14663 (N_14663,N_13674,N_14136);
and U14664 (N_14664,N_13620,N_13825);
or U14665 (N_14665,N_14222,N_14223);
nand U14666 (N_14666,N_14100,N_13685);
or U14667 (N_14667,N_13711,N_14050);
nand U14668 (N_14668,N_14164,N_14005);
xor U14669 (N_14669,N_13738,N_13627);
nand U14670 (N_14670,N_13805,N_14028);
xnor U14671 (N_14671,N_13502,N_14112);
and U14672 (N_14672,N_13966,N_14084);
xor U14673 (N_14673,N_13879,N_14203);
and U14674 (N_14674,N_13917,N_13924);
nor U14675 (N_14675,N_13770,N_13760);
nand U14676 (N_14676,N_13653,N_13556);
or U14677 (N_14677,N_14057,N_14083);
nand U14678 (N_14678,N_13824,N_13526);
nand U14679 (N_14679,N_14076,N_13725);
and U14680 (N_14680,N_13944,N_13672);
or U14681 (N_14681,N_13957,N_13593);
and U14682 (N_14682,N_13902,N_13678);
xnor U14683 (N_14683,N_13885,N_13963);
and U14684 (N_14684,N_13527,N_13593);
nand U14685 (N_14685,N_13918,N_14238);
and U14686 (N_14686,N_13585,N_14115);
or U14687 (N_14687,N_13798,N_14049);
or U14688 (N_14688,N_13570,N_13589);
xor U14689 (N_14689,N_13654,N_13693);
nor U14690 (N_14690,N_14017,N_13568);
nor U14691 (N_14691,N_13785,N_13637);
nand U14692 (N_14692,N_13671,N_14158);
and U14693 (N_14693,N_14151,N_14066);
and U14694 (N_14694,N_13630,N_14056);
or U14695 (N_14695,N_14000,N_13959);
xor U14696 (N_14696,N_14246,N_13764);
and U14697 (N_14697,N_14043,N_14090);
nand U14698 (N_14698,N_13578,N_13767);
xnor U14699 (N_14699,N_13971,N_13721);
or U14700 (N_14700,N_13760,N_14235);
xor U14701 (N_14701,N_13782,N_14039);
and U14702 (N_14702,N_14183,N_13976);
xor U14703 (N_14703,N_13860,N_14166);
nor U14704 (N_14704,N_13682,N_13627);
xnor U14705 (N_14705,N_14157,N_13695);
nand U14706 (N_14706,N_13522,N_13618);
or U14707 (N_14707,N_14226,N_14016);
xor U14708 (N_14708,N_13821,N_14003);
nor U14709 (N_14709,N_13635,N_14182);
xnor U14710 (N_14710,N_13810,N_14063);
nor U14711 (N_14711,N_14130,N_13690);
or U14712 (N_14712,N_14248,N_13982);
nand U14713 (N_14713,N_13964,N_14086);
nor U14714 (N_14714,N_13642,N_13927);
or U14715 (N_14715,N_13833,N_14197);
or U14716 (N_14716,N_13583,N_14081);
xor U14717 (N_14717,N_14226,N_13612);
nor U14718 (N_14718,N_13920,N_14095);
or U14719 (N_14719,N_13618,N_14103);
xnor U14720 (N_14720,N_13576,N_13899);
and U14721 (N_14721,N_14192,N_14195);
and U14722 (N_14722,N_13684,N_14049);
nand U14723 (N_14723,N_14079,N_14132);
and U14724 (N_14724,N_13690,N_14204);
xor U14725 (N_14725,N_13583,N_14178);
and U14726 (N_14726,N_14115,N_13688);
nand U14727 (N_14727,N_13929,N_14178);
nor U14728 (N_14728,N_13896,N_13705);
xnor U14729 (N_14729,N_14214,N_14008);
or U14730 (N_14730,N_13656,N_13997);
or U14731 (N_14731,N_13689,N_13814);
nor U14732 (N_14732,N_13922,N_13782);
nor U14733 (N_14733,N_13713,N_14121);
or U14734 (N_14734,N_14026,N_14093);
and U14735 (N_14735,N_13580,N_14229);
nand U14736 (N_14736,N_13978,N_13779);
xor U14737 (N_14737,N_13992,N_13673);
or U14738 (N_14738,N_14076,N_13945);
nand U14739 (N_14739,N_13629,N_14113);
nor U14740 (N_14740,N_13878,N_14067);
and U14741 (N_14741,N_13823,N_13749);
or U14742 (N_14742,N_13729,N_13675);
nand U14743 (N_14743,N_13657,N_14203);
nand U14744 (N_14744,N_13507,N_13576);
nor U14745 (N_14745,N_14093,N_13576);
and U14746 (N_14746,N_13515,N_13760);
or U14747 (N_14747,N_14108,N_13968);
nor U14748 (N_14748,N_13709,N_13890);
or U14749 (N_14749,N_14091,N_13877);
nor U14750 (N_14750,N_13967,N_13541);
xor U14751 (N_14751,N_14042,N_13760);
and U14752 (N_14752,N_13917,N_13528);
and U14753 (N_14753,N_13896,N_13988);
nand U14754 (N_14754,N_13594,N_13548);
and U14755 (N_14755,N_13858,N_14022);
nor U14756 (N_14756,N_13647,N_13563);
xor U14757 (N_14757,N_13967,N_13537);
or U14758 (N_14758,N_13945,N_13991);
nand U14759 (N_14759,N_13720,N_13713);
xor U14760 (N_14760,N_13973,N_13595);
xnor U14761 (N_14761,N_14081,N_13939);
nor U14762 (N_14762,N_13752,N_14072);
or U14763 (N_14763,N_13975,N_13700);
or U14764 (N_14764,N_14031,N_14113);
xor U14765 (N_14765,N_13708,N_14110);
and U14766 (N_14766,N_13735,N_13578);
and U14767 (N_14767,N_13553,N_13827);
xnor U14768 (N_14768,N_13950,N_14237);
nand U14769 (N_14769,N_13731,N_14089);
nand U14770 (N_14770,N_14220,N_13719);
nand U14771 (N_14771,N_14182,N_14156);
or U14772 (N_14772,N_13948,N_13678);
and U14773 (N_14773,N_13714,N_13927);
nor U14774 (N_14774,N_14107,N_13565);
nand U14775 (N_14775,N_13852,N_13548);
nor U14776 (N_14776,N_14163,N_13959);
nand U14777 (N_14777,N_13777,N_13524);
nand U14778 (N_14778,N_14050,N_14179);
nand U14779 (N_14779,N_14168,N_13530);
and U14780 (N_14780,N_13822,N_13642);
xnor U14781 (N_14781,N_13567,N_13849);
xor U14782 (N_14782,N_13820,N_13833);
nand U14783 (N_14783,N_13706,N_13546);
nand U14784 (N_14784,N_13869,N_13621);
and U14785 (N_14785,N_13628,N_14074);
nand U14786 (N_14786,N_13934,N_14117);
nand U14787 (N_14787,N_13980,N_13750);
nand U14788 (N_14788,N_13627,N_14020);
or U14789 (N_14789,N_13571,N_13549);
nor U14790 (N_14790,N_14021,N_14188);
or U14791 (N_14791,N_14081,N_14098);
and U14792 (N_14792,N_14240,N_13913);
and U14793 (N_14793,N_13968,N_13673);
and U14794 (N_14794,N_13838,N_13579);
nand U14795 (N_14795,N_14095,N_13584);
and U14796 (N_14796,N_13509,N_14043);
or U14797 (N_14797,N_14027,N_13912);
nor U14798 (N_14798,N_14168,N_13836);
or U14799 (N_14799,N_13525,N_13648);
or U14800 (N_14800,N_13616,N_13747);
or U14801 (N_14801,N_14036,N_13553);
and U14802 (N_14802,N_13615,N_13553);
or U14803 (N_14803,N_13670,N_13940);
nand U14804 (N_14804,N_13520,N_14112);
or U14805 (N_14805,N_14006,N_13714);
nor U14806 (N_14806,N_13782,N_14084);
xor U14807 (N_14807,N_14204,N_13721);
or U14808 (N_14808,N_13993,N_14205);
or U14809 (N_14809,N_13585,N_14177);
nand U14810 (N_14810,N_13623,N_13949);
nand U14811 (N_14811,N_13597,N_13631);
xor U14812 (N_14812,N_13999,N_13980);
nand U14813 (N_14813,N_14011,N_13710);
nor U14814 (N_14814,N_13933,N_14100);
xor U14815 (N_14815,N_13912,N_13741);
or U14816 (N_14816,N_13688,N_14086);
nor U14817 (N_14817,N_13701,N_13873);
xnor U14818 (N_14818,N_13934,N_13504);
and U14819 (N_14819,N_13631,N_13652);
nor U14820 (N_14820,N_14181,N_14205);
nand U14821 (N_14821,N_13853,N_13717);
or U14822 (N_14822,N_13556,N_13510);
or U14823 (N_14823,N_14129,N_14218);
and U14824 (N_14824,N_13503,N_13719);
nor U14825 (N_14825,N_13882,N_14106);
and U14826 (N_14826,N_14134,N_13917);
xor U14827 (N_14827,N_14149,N_14152);
and U14828 (N_14828,N_14045,N_13741);
nand U14829 (N_14829,N_14203,N_13752);
or U14830 (N_14830,N_13964,N_13823);
nor U14831 (N_14831,N_13702,N_13916);
and U14832 (N_14832,N_14226,N_13615);
nor U14833 (N_14833,N_13857,N_13995);
nand U14834 (N_14834,N_13870,N_14224);
nand U14835 (N_14835,N_13515,N_13739);
xnor U14836 (N_14836,N_13840,N_13679);
or U14837 (N_14837,N_13715,N_14218);
nand U14838 (N_14838,N_13933,N_13723);
or U14839 (N_14839,N_14187,N_14057);
nor U14840 (N_14840,N_14230,N_14203);
or U14841 (N_14841,N_13656,N_14089);
xnor U14842 (N_14842,N_14090,N_14012);
nor U14843 (N_14843,N_14178,N_13986);
and U14844 (N_14844,N_13551,N_13517);
or U14845 (N_14845,N_14118,N_13807);
and U14846 (N_14846,N_13844,N_13526);
xor U14847 (N_14847,N_13664,N_14153);
and U14848 (N_14848,N_14145,N_13742);
xor U14849 (N_14849,N_13612,N_13514);
and U14850 (N_14850,N_13915,N_13663);
nor U14851 (N_14851,N_14030,N_13908);
xor U14852 (N_14852,N_13704,N_13642);
or U14853 (N_14853,N_13886,N_14009);
xnor U14854 (N_14854,N_13572,N_13925);
and U14855 (N_14855,N_13935,N_13898);
nor U14856 (N_14856,N_13529,N_13923);
xor U14857 (N_14857,N_13804,N_13660);
nor U14858 (N_14858,N_13898,N_13716);
nor U14859 (N_14859,N_14111,N_13787);
or U14860 (N_14860,N_13717,N_14037);
and U14861 (N_14861,N_13800,N_13602);
nor U14862 (N_14862,N_14070,N_14015);
xor U14863 (N_14863,N_13634,N_14218);
nor U14864 (N_14864,N_13540,N_13544);
nor U14865 (N_14865,N_13526,N_13854);
xnor U14866 (N_14866,N_13514,N_13806);
nor U14867 (N_14867,N_13944,N_13793);
xnor U14868 (N_14868,N_14213,N_13527);
nor U14869 (N_14869,N_13983,N_13741);
nor U14870 (N_14870,N_13836,N_13977);
nand U14871 (N_14871,N_13913,N_13966);
or U14872 (N_14872,N_14213,N_13793);
and U14873 (N_14873,N_13612,N_14018);
and U14874 (N_14874,N_13596,N_14119);
nor U14875 (N_14875,N_14126,N_13588);
nand U14876 (N_14876,N_13563,N_13529);
nor U14877 (N_14877,N_13763,N_13513);
xor U14878 (N_14878,N_14024,N_13918);
nand U14879 (N_14879,N_13772,N_13676);
or U14880 (N_14880,N_13521,N_13954);
or U14881 (N_14881,N_14208,N_14067);
xnor U14882 (N_14882,N_13850,N_13547);
nor U14883 (N_14883,N_13693,N_13562);
nor U14884 (N_14884,N_13852,N_14067);
nor U14885 (N_14885,N_13630,N_13834);
nor U14886 (N_14886,N_13730,N_13961);
nand U14887 (N_14887,N_13960,N_13584);
xor U14888 (N_14888,N_13500,N_13607);
or U14889 (N_14889,N_13644,N_14192);
and U14890 (N_14890,N_13742,N_14047);
nor U14891 (N_14891,N_13652,N_14182);
and U14892 (N_14892,N_13654,N_14063);
nor U14893 (N_14893,N_13502,N_13860);
nor U14894 (N_14894,N_14223,N_13957);
and U14895 (N_14895,N_13958,N_14195);
xor U14896 (N_14896,N_13631,N_14168);
nand U14897 (N_14897,N_14176,N_14132);
xor U14898 (N_14898,N_14031,N_13839);
nand U14899 (N_14899,N_13537,N_13724);
and U14900 (N_14900,N_13535,N_13647);
and U14901 (N_14901,N_14033,N_14052);
and U14902 (N_14902,N_14001,N_13647);
and U14903 (N_14903,N_14203,N_13826);
xor U14904 (N_14904,N_14074,N_13654);
and U14905 (N_14905,N_14171,N_13583);
and U14906 (N_14906,N_13542,N_13712);
nand U14907 (N_14907,N_13602,N_13788);
nand U14908 (N_14908,N_13587,N_13927);
nand U14909 (N_14909,N_13812,N_13773);
and U14910 (N_14910,N_14161,N_13894);
nor U14911 (N_14911,N_13675,N_13900);
or U14912 (N_14912,N_13519,N_14119);
and U14913 (N_14913,N_13522,N_13933);
nor U14914 (N_14914,N_14024,N_13946);
xnor U14915 (N_14915,N_14146,N_13565);
nor U14916 (N_14916,N_13769,N_13966);
or U14917 (N_14917,N_14215,N_14085);
nand U14918 (N_14918,N_13690,N_14173);
or U14919 (N_14919,N_13891,N_14210);
xor U14920 (N_14920,N_14121,N_14176);
nor U14921 (N_14921,N_14242,N_13809);
nand U14922 (N_14922,N_13859,N_14163);
xor U14923 (N_14923,N_13810,N_13821);
xnor U14924 (N_14924,N_13633,N_13790);
xor U14925 (N_14925,N_14056,N_13741);
nand U14926 (N_14926,N_13928,N_13683);
nand U14927 (N_14927,N_13774,N_14119);
and U14928 (N_14928,N_14020,N_13914);
and U14929 (N_14929,N_13961,N_14152);
nand U14930 (N_14930,N_13517,N_14010);
and U14931 (N_14931,N_13814,N_14209);
xor U14932 (N_14932,N_14100,N_13610);
xor U14933 (N_14933,N_13837,N_13596);
or U14934 (N_14934,N_13600,N_13579);
nand U14935 (N_14935,N_14165,N_13929);
nor U14936 (N_14936,N_13515,N_13900);
xor U14937 (N_14937,N_13785,N_13726);
and U14938 (N_14938,N_14061,N_13875);
nor U14939 (N_14939,N_14121,N_13819);
nand U14940 (N_14940,N_13624,N_13833);
nand U14941 (N_14941,N_13963,N_13653);
nor U14942 (N_14942,N_13748,N_13712);
xor U14943 (N_14943,N_13658,N_13871);
nand U14944 (N_14944,N_13768,N_13767);
and U14945 (N_14945,N_14091,N_14148);
nand U14946 (N_14946,N_14070,N_14193);
xor U14947 (N_14947,N_13744,N_14035);
nand U14948 (N_14948,N_14070,N_14182);
xor U14949 (N_14949,N_13647,N_13678);
and U14950 (N_14950,N_14194,N_13546);
nand U14951 (N_14951,N_13812,N_13658);
nand U14952 (N_14952,N_13707,N_13801);
and U14953 (N_14953,N_13839,N_13653);
xor U14954 (N_14954,N_13566,N_14096);
xor U14955 (N_14955,N_14131,N_13675);
xor U14956 (N_14956,N_13550,N_13523);
or U14957 (N_14957,N_14020,N_14010);
nand U14958 (N_14958,N_13563,N_14059);
or U14959 (N_14959,N_14032,N_13886);
or U14960 (N_14960,N_14026,N_14124);
nor U14961 (N_14961,N_13952,N_13734);
xor U14962 (N_14962,N_13787,N_13969);
xnor U14963 (N_14963,N_13570,N_14211);
or U14964 (N_14964,N_13639,N_14022);
nand U14965 (N_14965,N_13964,N_14111);
or U14966 (N_14966,N_13519,N_14008);
or U14967 (N_14967,N_13886,N_13983);
or U14968 (N_14968,N_13522,N_13896);
xor U14969 (N_14969,N_13742,N_14112);
xnor U14970 (N_14970,N_13905,N_13948);
xor U14971 (N_14971,N_14111,N_14202);
and U14972 (N_14972,N_13942,N_13636);
nor U14973 (N_14973,N_13825,N_14218);
or U14974 (N_14974,N_14201,N_13661);
and U14975 (N_14975,N_13605,N_13633);
and U14976 (N_14976,N_13539,N_14049);
xnor U14977 (N_14977,N_13664,N_13571);
nand U14978 (N_14978,N_13771,N_13940);
and U14979 (N_14979,N_13652,N_13612);
nand U14980 (N_14980,N_13594,N_14214);
or U14981 (N_14981,N_14013,N_13913);
xnor U14982 (N_14982,N_13594,N_13572);
or U14983 (N_14983,N_14145,N_14173);
or U14984 (N_14984,N_13577,N_14248);
nand U14985 (N_14985,N_13706,N_13774);
or U14986 (N_14986,N_13563,N_13501);
or U14987 (N_14987,N_13863,N_13596);
and U14988 (N_14988,N_13736,N_13744);
nor U14989 (N_14989,N_13878,N_14152);
and U14990 (N_14990,N_13814,N_14211);
xor U14991 (N_14991,N_13807,N_14135);
xor U14992 (N_14992,N_13513,N_13707);
nand U14993 (N_14993,N_13528,N_14180);
or U14994 (N_14994,N_13754,N_13601);
nand U14995 (N_14995,N_13738,N_14170);
nor U14996 (N_14996,N_14052,N_13708);
xnor U14997 (N_14997,N_14238,N_14123);
nand U14998 (N_14998,N_14038,N_14016);
xor U14999 (N_14999,N_14053,N_13817);
xnor UO_0 (O_0,N_14542,N_14556);
nand UO_1 (O_1,N_14665,N_14694);
nand UO_2 (O_2,N_14641,N_14440);
or UO_3 (O_3,N_14916,N_14298);
nor UO_4 (O_4,N_14423,N_14264);
or UO_5 (O_5,N_14553,N_14319);
nor UO_6 (O_6,N_14770,N_14984);
xor UO_7 (O_7,N_14502,N_14890);
or UO_8 (O_8,N_14882,N_14708);
xnor UO_9 (O_9,N_14924,N_14449);
nor UO_10 (O_10,N_14596,N_14413);
nand UO_11 (O_11,N_14383,N_14995);
or UO_12 (O_12,N_14853,N_14799);
or UO_13 (O_13,N_14583,N_14565);
and UO_14 (O_14,N_14636,N_14490);
xor UO_15 (O_15,N_14633,N_14331);
or UO_16 (O_16,N_14758,N_14558);
nand UO_17 (O_17,N_14524,N_14399);
nand UO_18 (O_18,N_14482,N_14888);
nand UO_19 (O_19,N_14274,N_14554);
nand UO_20 (O_20,N_14541,N_14921);
and UO_21 (O_21,N_14766,N_14481);
nor UO_22 (O_22,N_14914,N_14687);
xor UO_23 (O_23,N_14631,N_14259);
xor UO_24 (O_24,N_14785,N_14326);
or UO_25 (O_25,N_14877,N_14963);
or UO_26 (O_26,N_14266,N_14838);
or UO_27 (O_27,N_14858,N_14437);
nor UO_28 (O_28,N_14485,N_14262);
and UO_29 (O_29,N_14508,N_14709);
nor UO_30 (O_30,N_14342,N_14599);
nor UO_31 (O_31,N_14892,N_14464);
or UO_32 (O_32,N_14957,N_14864);
xnor UO_33 (O_33,N_14945,N_14487);
or UO_34 (O_34,N_14412,N_14279);
and UO_35 (O_35,N_14462,N_14947);
or UO_36 (O_36,N_14314,N_14704);
or UO_37 (O_37,N_14680,N_14375);
nand UO_38 (O_38,N_14675,N_14801);
nand UO_39 (O_39,N_14357,N_14926);
and UO_40 (O_40,N_14610,N_14251);
nor UO_41 (O_41,N_14579,N_14951);
nor UO_42 (O_42,N_14880,N_14370);
and UO_43 (O_43,N_14460,N_14682);
nand UO_44 (O_44,N_14563,N_14564);
xor UO_45 (O_45,N_14250,N_14330);
nand UO_46 (O_46,N_14852,N_14691);
xor UO_47 (O_47,N_14513,N_14588);
and UO_48 (O_48,N_14639,N_14949);
xor UO_49 (O_49,N_14561,N_14846);
nand UO_50 (O_50,N_14891,N_14574);
xnor UO_51 (O_51,N_14716,N_14897);
nand UO_52 (O_52,N_14611,N_14403);
xnor UO_53 (O_53,N_14782,N_14476);
nand UO_54 (O_54,N_14387,N_14982);
nor UO_55 (O_55,N_14968,N_14965);
xor UO_56 (O_56,N_14505,N_14277);
nor UO_57 (O_57,N_14337,N_14724);
nor UO_58 (O_58,N_14964,N_14350);
nor UO_59 (O_59,N_14759,N_14878);
nor UO_60 (O_60,N_14769,N_14281);
xnor UO_61 (O_61,N_14261,N_14934);
and UO_62 (O_62,N_14318,N_14991);
or UO_63 (O_63,N_14567,N_14378);
nor UO_64 (O_64,N_14754,N_14252);
nand UO_65 (O_65,N_14349,N_14922);
nor UO_66 (O_66,N_14276,N_14933);
nand UO_67 (O_67,N_14278,N_14551);
nand UO_68 (O_68,N_14421,N_14500);
or UO_69 (O_69,N_14900,N_14819);
xnor UO_70 (O_70,N_14550,N_14268);
nand UO_71 (O_71,N_14428,N_14534);
and UO_72 (O_72,N_14712,N_14334);
nand UO_73 (O_73,N_14673,N_14685);
or UO_74 (O_74,N_14750,N_14339);
and UO_75 (O_75,N_14745,N_14803);
nand UO_76 (O_76,N_14400,N_14340);
nor UO_77 (O_77,N_14828,N_14280);
and UO_78 (O_78,N_14355,N_14875);
nor UO_79 (O_79,N_14929,N_14736);
nand UO_80 (O_80,N_14742,N_14402);
and UO_81 (O_81,N_14919,N_14970);
or UO_82 (O_82,N_14771,N_14453);
nand UO_83 (O_83,N_14604,N_14265);
nand UO_84 (O_84,N_14452,N_14931);
xor UO_85 (O_85,N_14672,N_14966);
or UO_86 (O_86,N_14836,N_14284);
and UO_87 (O_87,N_14637,N_14824);
nand UO_88 (O_88,N_14841,N_14523);
xor UO_89 (O_89,N_14371,N_14729);
or UO_90 (O_90,N_14868,N_14384);
nand UO_91 (O_91,N_14696,N_14862);
and UO_92 (O_92,N_14415,N_14952);
nor UO_93 (O_93,N_14789,N_14308);
nor UO_94 (O_94,N_14743,N_14559);
xnor UO_95 (O_95,N_14393,N_14478);
nand UO_96 (O_96,N_14796,N_14869);
xnor UO_97 (O_97,N_14444,N_14661);
nand UO_98 (O_98,N_14320,N_14812);
xnor UO_99 (O_99,N_14755,N_14999);
and UO_100 (O_100,N_14938,N_14411);
or UO_101 (O_101,N_14373,N_14312);
xnor UO_102 (O_102,N_14871,N_14809);
or UO_103 (O_103,N_14840,N_14630);
or UO_104 (O_104,N_14867,N_14917);
xnor UO_105 (O_105,N_14904,N_14735);
nand UO_106 (O_106,N_14446,N_14823);
or UO_107 (O_107,N_14733,N_14529);
nor UO_108 (O_108,N_14580,N_14613);
xor UO_109 (O_109,N_14748,N_14351);
or UO_110 (O_110,N_14686,N_14315);
xnor UO_111 (O_111,N_14594,N_14407);
nor UO_112 (O_112,N_14689,N_14555);
nor UO_113 (O_113,N_14872,N_14722);
xor UO_114 (O_114,N_14540,N_14532);
xor UO_115 (O_115,N_14698,N_14323);
xor UO_116 (O_116,N_14959,N_14333);
nor UO_117 (O_117,N_14292,N_14723);
nand UO_118 (O_118,N_14707,N_14902);
or UO_119 (O_119,N_14635,N_14971);
nand UO_120 (O_120,N_14394,N_14692);
nor UO_121 (O_121,N_14644,N_14480);
and UO_122 (O_122,N_14918,N_14396);
xor UO_123 (O_123,N_14688,N_14911);
or UO_124 (O_124,N_14424,N_14659);
or UO_125 (O_125,N_14622,N_14417);
or UO_126 (O_126,N_14710,N_14512);
nand UO_127 (O_127,N_14730,N_14625);
or UO_128 (O_128,N_14653,N_14587);
nor UO_129 (O_129,N_14711,N_14619);
nand UO_130 (O_130,N_14458,N_14632);
or UO_131 (O_131,N_14270,N_14360);
and UO_132 (O_132,N_14560,N_14607);
xnor UO_133 (O_133,N_14740,N_14905);
nor UO_134 (O_134,N_14954,N_14527);
xnor UO_135 (O_135,N_14294,N_14649);
nand UO_136 (O_136,N_14996,N_14346);
nor UO_137 (O_137,N_14465,N_14570);
nand UO_138 (O_138,N_14648,N_14420);
or UO_139 (O_139,N_14662,N_14806);
and UO_140 (O_140,N_14794,N_14805);
nand UO_141 (O_141,N_14489,N_14863);
or UO_142 (O_142,N_14398,N_14498);
and UO_143 (O_143,N_14706,N_14848);
and UO_144 (O_144,N_14908,N_14376);
xnor UO_145 (O_145,N_14448,N_14557);
and UO_146 (O_146,N_14749,N_14666);
nand UO_147 (O_147,N_14395,N_14426);
nand UO_148 (O_148,N_14486,N_14545);
xor UO_149 (O_149,N_14844,N_14255);
and UO_150 (O_150,N_14516,N_14324);
xor UO_151 (O_151,N_14416,N_14501);
nor UO_152 (O_152,N_14504,N_14650);
nand UO_153 (O_153,N_14263,N_14721);
or UO_154 (O_154,N_14483,N_14693);
nor UO_155 (O_155,N_14998,N_14569);
xnor UO_156 (O_156,N_14859,N_14920);
and UO_157 (O_157,N_14296,N_14906);
xor UO_158 (O_158,N_14623,N_14760);
and UO_159 (O_159,N_14930,N_14629);
nand UO_160 (O_160,N_14592,N_14356);
or UO_161 (O_161,N_14311,N_14443);
nand UO_162 (O_162,N_14329,N_14595);
xnor UO_163 (O_163,N_14492,N_14690);
nand UO_164 (O_164,N_14850,N_14804);
nor UO_165 (O_165,N_14295,N_14621);
xnor UO_166 (O_166,N_14586,N_14600);
and UO_167 (O_167,N_14883,N_14461);
nand UO_168 (O_168,N_14969,N_14992);
nand UO_169 (O_169,N_14361,N_14454);
nor UO_170 (O_170,N_14435,N_14386);
nor UO_171 (O_171,N_14896,N_14566);
xnor UO_172 (O_172,N_14624,N_14466);
nor UO_173 (O_173,N_14946,N_14471);
nor UO_174 (O_174,N_14885,N_14327);
and UO_175 (O_175,N_14705,N_14839);
xor UO_176 (O_176,N_14288,N_14404);
and UO_177 (O_177,N_14347,N_14354);
xnor UO_178 (O_178,N_14937,N_14577);
and UO_179 (O_179,N_14652,N_14479);
or UO_180 (O_180,N_14656,N_14677);
or UO_181 (O_181,N_14293,N_14974);
nand UO_182 (O_182,N_14562,N_14581);
nor UO_183 (O_183,N_14683,N_14681);
nand UO_184 (O_184,N_14713,N_14870);
and UO_185 (O_185,N_14747,N_14299);
nand UO_186 (O_186,N_14283,N_14301);
nor UO_187 (O_187,N_14651,N_14257);
xor UO_188 (O_188,N_14978,N_14663);
xor UO_189 (O_189,N_14338,N_14522);
xor UO_190 (O_190,N_14432,N_14985);
and UO_191 (O_191,N_14741,N_14436);
nor UO_192 (O_192,N_14539,N_14856);
or UO_193 (O_193,N_14365,N_14544);
nor UO_194 (O_194,N_14936,N_14297);
nor UO_195 (O_195,N_14406,N_14389);
nor UO_196 (O_196,N_14793,N_14660);
xor UO_197 (O_197,N_14367,N_14700);
nor UO_198 (O_198,N_14955,N_14752);
or UO_199 (O_199,N_14605,N_14484);
nor UO_200 (O_200,N_14585,N_14874);
nand UO_201 (O_201,N_14463,N_14470);
and UO_202 (O_202,N_14341,N_14753);
nor UO_203 (O_203,N_14617,N_14849);
and UO_204 (O_204,N_14667,N_14986);
and UO_205 (O_205,N_14517,N_14571);
xnor UO_206 (O_206,N_14441,N_14515);
xor UO_207 (O_207,N_14438,N_14835);
nor UO_208 (O_208,N_14409,N_14887);
nor UO_209 (O_209,N_14668,N_14410);
or UO_210 (O_210,N_14684,N_14451);
xnor UO_211 (O_211,N_14598,N_14772);
nand UO_212 (O_212,N_14302,N_14290);
xor UO_213 (O_213,N_14788,N_14953);
xnor UO_214 (O_214,N_14495,N_14943);
and UO_215 (O_215,N_14510,N_14275);
xor UO_216 (O_216,N_14431,N_14855);
and UO_217 (O_217,N_14348,N_14382);
nor UO_218 (O_218,N_14552,N_14972);
nor UO_219 (O_219,N_14285,N_14695);
and UO_220 (O_220,N_14989,N_14572);
or UO_221 (O_221,N_14427,N_14608);
nand UO_222 (O_222,N_14286,N_14520);
and UO_223 (O_223,N_14603,N_14895);
nand UO_224 (O_224,N_14702,N_14537);
and UO_225 (O_225,N_14976,N_14575);
and UO_226 (O_226,N_14763,N_14303);
nor UO_227 (O_227,N_14674,N_14948);
xnor UO_228 (O_228,N_14925,N_14573);
or UO_229 (O_229,N_14457,N_14634);
nor UO_230 (O_230,N_14519,N_14780);
xor UO_231 (O_231,N_14352,N_14894);
nor UO_232 (O_232,N_14739,N_14815);
nor UO_233 (O_233,N_14843,N_14783);
or UO_234 (O_234,N_14291,N_14851);
nor UO_235 (O_235,N_14313,N_14734);
nor UO_236 (O_236,N_14973,N_14678);
xor UO_237 (O_237,N_14792,N_14363);
or UO_238 (O_238,N_14514,N_14493);
and UO_239 (O_239,N_14774,N_14576);
xor UO_240 (O_240,N_14939,N_14533);
and UO_241 (O_241,N_14791,N_14993);
and UO_242 (O_242,N_14385,N_14761);
nor UO_243 (O_243,N_14322,N_14518);
nand UO_244 (O_244,N_14615,N_14956);
nor UO_245 (O_245,N_14807,N_14456);
nand UO_246 (O_246,N_14756,N_14548);
nand UO_247 (O_247,N_14781,N_14343);
and UO_248 (O_248,N_14467,N_14353);
xor UO_249 (O_249,N_14601,N_14697);
nor UO_250 (O_250,N_14627,N_14638);
nor UO_251 (O_251,N_14990,N_14810);
or UO_252 (O_252,N_14475,N_14818);
and UO_253 (O_253,N_14256,N_14907);
and UO_254 (O_254,N_14988,N_14776);
nand UO_255 (O_255,N_14271,N_14831);
nand UO_256 (O_256,N_14857,N_14310);
nand UO_257 (O_257,N_14531,N_14307);
nand UO_258 (O_258,N_14287,N_14549);
and UO_259 (O_259,N_14765,N_14726);
and UO_260 (O_260,N_14983,N_14751);
nand UO_261 (O_261,N_14606,N_14808);
nor UO_262 (O_262,N_14344,N_14414);
nor UO_263 (O_263,N_14521,N_14827);
or UO_264 (O_264,N_14737,N_14811);
xor UO_265 (O_265,N_14787,N_14506);
and UO_266 (O_266,N_14718,N_14260);
and UO_267 (O_267,N_14813,N_14701);
nor UO_268 (O_268,N_14817,N_14738);
xor UO_269 (O_269,N_14655,N_14829);
nor UO_270 (O_270,N_14790,N_14732);
and UO_271 (O_271,N_14826,N_14477);
nand UO_272 (O_272,N_14507,N_14590);
nand UO_273 (O_273,N_14731,N_14884);
and UO_274 (O_274,N_14720,N_14474);
nor UO_275 (O_275,N_14499,N_14496);
xor UO_276 (O_276,N_14703,N_14802);
xor UO_277 (O_277,N_14860,N_14616);
and UO_278 (O_278,N_14380,N_14401);
or UO_279 (O_279,N_14762,N_14670);
and UO_280 (O_280,N_14913,N_14997);
xnor UO_281 (O_281,N_14372,N_14643);
nand UO_282 (O_282,N_14535,N_14669);
nor UO_283 (O_283,N_14422,N_14779);
xor UO_284 (O_284,N_14795,N_14980);
nand UO_285 (O_285,N_14910,N_14321);
and UO_286 (O_286,N_14775,N_14744);
nor UO_287 (O_287,N_14473,N_14254);
or UO_288 (O_288,N_14854,N_14899);
nor UO_289 (O_289,N_14935,N_14447);
nor UO_290 (O_290,N_14364,N_14543);
xnor UO_291 (O_291,N_14469,N_14253);
and UO_292 (O_292,N_14830,N_14317);
xnor UO_293 (O_293,N_14358,N_14958);
and UO_294 (O_294,N_14994,N_14797);
xor UO_295 (O_295,N_14306,N_14778);
or UO_296 (O_296,N_14433,N_14391);
nand UO_297 (O_297,N_14784,N_14430);
xnor UO_298 (O_298,N_14960,N_14408);
xor UO_299 (O_299,N_14273,N_14881);
nand UO_300 (O_300,N_14923,N_14834);
xor UO_301 (O_301,N_14379,N_14397);
and UO_302 (O_302,N_14450,N_14578);
nor UO_303 (O_303,N_14614,N_14981);
nor UO_304 (O_304,N_14491,N_14717);
xnor UO_305 (O_305,N_14975,N_14366);
nor UO_306 (O_306,N_14377,N_14488);
nand UO_307 (O_307,N_14773,N_14511);
nor UO_308 (O_308,N_14272,N_14626);
nor UO_309 (O_309,N_14679,N_14865);
and UO_310 (O_310,N_14419,N_14786);
nand UO_311 (O_311,N_14445,N_14258);
xnor UO_312 (O_312,N_14359,N_14332);
and UO_313 (O_313,N_14584,N_14942);
xor UO_314 (O_314,N_14442,N_14876);
or UO_315 (O_315,N_14645,N_14825);
nand UO_316 (O_316,N_14374,N_14950);
or UO_317 (O_317,N_14757,N_14530);
nand UO_318 (O_318,N_14612,N_14597);
or UO_319 (O_319,N_14434,N_14335);
nand UO_320 (O_320,N_14593,N_14336);
xor UO_321 (O_321,N_14676,N_14833);
nor UO_322 (O_322,N_14628,N_14368);
xnor UO_323 (O_323,N_14715,N_14889);
xnor UO_324 (O_324,N_14468,N_14509);
nand UO_325 (O_325,N_14699,N_14439);
and UO_326 (O_326,N_14962,N_14901);
nand UO_327 (O_327,N_14746,N_14664);
and UO_328 (O_328,N_14903,N_14714);
xnor UO_329 (O_329,N_14886,N_14362);
xnor UO_330 (O_330,N_14609,N_14820);
nor UO_331 (O_331,N_14728,N_14832);
nand UO_332 (O_332,N_14912,N_14381);
nor UO_333 (O_333,N_14842,N_14642);
nor UO_334 (O_334,N_14282,N_14525);
xor UO_335 (O_335,N_14671,N_14316);
nand UO_336 (O_336,N_14909,N_14987);
nor UO_337 (O_337,N_14602,N_14503);
xor UO_338 (O_338,N_14618,N_14289);
nand UO_339 (O_339,N_14494,N_14429);
and UO_340 (O_340,N_14547,N_14657);
nor UO_341 (O_341,N_14879,N_14944);
xor UO_342 (O_342,N_14837,N_14658);
or UO_343 (O_343,N_14405,N_14455);
and UO_344 (O_344,N_14768,N_14979);
nor UO_345 (O_345,N_14767,N_14727);
xor UO_346 (O_346,N_14418,N_14928);
xor UO_347 (O_347,N_14941,N_14345);
and UO_348 (O_348,N_14568,N_14725);
or UO_349 (O_349,N_14269,N_14816);
nor UO_350 (O_350,N_14764,N_14873);
xnor UO_351 (O_351,N_14425,N_14961);
nor UO_352 (O_352,N_14369,N_14647);
xor UO_353 (O_353,N_14915,N_14528);
and UO_354 (O_354,N_14459,N_14967);
xnor UO_355 (O_355,N_14821,N_14392);
xor UO_356 (O_356,N_14497,N_14893);
nor UO_357 (O_357,N_14390,N_14546);
nand UO_358 (O_358,N_14305,N_14814);
nor UO_359 (O_359,N_14526,N_14845);
xnor UO_360 (O_360,N_14654,N_14719);
xnor UO_361 (O_361,N_14822,N_14300);
nand UO_362 (O_362,N_14898,N_14325);
and UO_363 (O_363,N_14589,N_14536);
xnor UO_364 (O_364,N_14861,N_14932);
and UO_365 (O_365,N_14847,N_14646);
or UO_366 (O_366,N_14472,N_14328);
nand UO_367 (O_367,N_14309,N_14777);
and UO_368 (O_368,N_14977,N_14620);
nor UO_369 (O_369,N_14940,N_14640);
or UO_370 (O_370,N_14800,N_14591);
xnor UO_371 (O_371,N_14927,N_14304);
and UO_372 (O_372,N_14582,N_14538);
and UO_373 (O_373,N_14388,N_14866);
or UO_374 (O_374,N_14267,N_14798);
xor UO_375 (O_375,N_14664,N_14805);
xnor UO_376 (O_376,N_14795,N_14428);
nor UO_377 (O_377,N_14393,N_14879);
nand UO_378 (O_378,N_14974,N_14933);
xnor UO_379 (O_379,N_14657,N_14708);
nand UO_380 (O_380,N_14457,N_14843);
nand UO_381 (O_381,N_14673,N_14479);
xor UO_382 (O_382,N_14352,N_14556);
xnor UO_383 (O_383,N_14856,N_14870);
or UO_384 (O_384,N_14296,N_14397);
nor UO_385 (O_385,N_14510,N_14687);
or UO_386 (O_386,N_14361,N_14908);
xnor UO_387 (O_387,N_14403,N_14628);
nor UO_388 (O_388,N_14530,N_14444);
xor UO_389 (O_389,N_14882,N_14435);
or UO_390 (O_390,N_14997,N_14569);
nor UO_391 (O_391,N_14935,N_14765);
nand UO_392 (O_392,N_14250,N_14838);
and UO_393 (O_393,N_14653,N_14552);
or UO_394 (O_394,N_14956,N_14664);
and UO_395 (O_395,N_14368,N_14646);
xor UO_396 (O_396,N_14768,N_14967);
nor UO_397 (O_397,N_14950,N_14784);
and UO_398 (O_398,N_14390,N_14955);
or UO_399 (O_399,N_14870,N_14573);
nand UO_400 (O_400,N_14380,N_14654);
nand UO_401 (O_401,N_14587,N_14300);
nand UO_402 (O_402,N_14970,N_14279);
or UO_403 (O_403,N_14765,N_14617);
nand UO_404 (O_404,N_14387,N_14354);
nand UO_405 (O_405,N_14282,N_14552);
xor UO_406 (O_406,N_14745,N_14705);
or UO_407 (O_407,N_14673,N_14884);
nand UO_408 (O_408,N_14726,N_14775);
and UO_409 (O_409,N_14582,N_14729);
or UO_410 (O_410,N_14993,N_14796);
and UO_411 (O_411,N_14255,N_14842);
or UO_412 (O_412,N_14405,N_14313);
nand UO_413 (O_413,N_14362,N_14861);
nand UO_414 (O_414,N_14818,N_14693);
and UO_415 (O_415,N_14758,N_14848);
or UO_416 (O_416,N_14764,N_14598);
and UO_417 (O_417,N_14855,N_14964);
and UO_418 (O_418,N_14563,N_14780);
xnor UO_419 (O_419,N_14408,N_14896);
xor UO_420 (O_420,N_14580,N_14434);
nand UO_421 (O_421,N_14467,N_14301);
nand UO_422 (O_422,N_14317,N_14624);
or UO_423 (O_423,N_14360,N_14851);
nand UO_424 (O_424,N_14468,N_14972);
xnor UO_425 (O_425,N_14384,N_14412);
xor UO_426 (O_426,N_14699,N_14307);
and UO_427 (O_427,N_14818,N_14961);
nor UO_428 (O_428,N_14908,N_14297);
nand UO_429 (O_429,N_14641,N_14900);
nor UO_430 (O_430,N_14398,N_14992);
and UO_431 (O_431,N_14630,N_14616);
nand UO_432 (O_432,N_14801,N_14677);
nor UO_433 (O_433,N_14347,N_14583);
nor UO_434 (O_434,N_14313,N_14294);
xnor UO_435 (O_435,N_14931,N_14500);
nor UO_436 (O_436,N_14450,N_14308);
or UO_437 (O_437,N_14606,N_14682);
or UO_438 (O_438,N_14576,N_14495);
nand UO_439 (O_439,N_14758,N_14363);
nor UO_440 (O_440,N_14893,N_14648);
nand UO_441 (O_441,N_14471,N_14624);
and UO_442 (O_442,N_14714,N_14608);
nor UO_443 (O_443,N_14711,N_14944);
nand UO_444 (O_444,N_14421,N_14579);
and UO_445 (O_445,N_14913,N_14798);
and UO_446 (O_446,N_14715,N_14906);
nand UO_447 (O_447,N_14579,N_14623);
or UO_448 (O_448,N_14733,N_14361);
and UO_449 (O_449,N_14587,N_14721);
nand UO_450 (O_450,N_14726,N_14874);
or UO_451 (O_451,N_14806,N_14671);
nor UO_452 (O_452,N_14866,N_14501);
nor UO_453 (O_453,N_14527,N_14502);
nand UO_454 (O_454,N_14299,N_14341);
or UO_455 (O_455,N_14471,N_14450);
nor UO_456 (O_456,N_14661,N_14311);
and UO_457 (O_457,N_14609,N_14346);
or UO_458 (O_458,N_14766,N_14420);
nand UO_459 (O_459,N_14964,N_14989);
xnor UO_460 (O_460,N_14624,N_14329);
nor UO_461 (O_461,N_14773,N_14796);
nand UO_462 (O_462,N_14747,N_14499);
or UO_463 (O_463,N_14270,N_14738);
and UO_464 (O_464,N_14269,N_14541);
or UO_465 (O_465,N_14744,N_14872);
and UO_466 (O_466,N_14818,N_14965);
nor UO_467 (O_467,N_14736,N_14658);
nand UO_468 (O_468,N_14442,N_14494);
nor UO_469 (O_469,N_14263,N_14367);
nor UO_470 (O_470,N_14474,N_14500);
or UO_471 (O_471,N_14846,N_14535);
xor UO_472 (O_472,N_14574,N_14445);
or UO_473 (O_473,N_14871,N_14722);
nand UO_474 (O_474,N_14396,N_14282);
xnor UO_475 (O_475,N_14388,N_14627);
nor UO_476 (O_476,N_14307,N_14741);
and UO_477 (O_477,N_14496,N_14743);
nand UO_478 (O_478,N_14913,N_14518);
nor UO_479 (O_479,N_14792,N_14615);
and UO_480 (O_480,N_14369,N_14955);
nor UO_481 (O_481,N_14417,N_14857);
xor UO_482 (O_482,N_14427,N_14951);
xnor UO_483 (O_483,N_14520,N_14744);
and UO_484 (O_484,N_14764,N_14590);
nand UO_485 (O_485,N_14965,N_14650);
and UO_486 (O_486,N_14367,N_14309);
xor UO_487 (O_487,N_14791,N_14638);
and UO_488 (O_488,N_14432,N_14568);
xnor UO_489 (O_489,N_14550,N_14433);
and UO_490 (O_490,N_14781,N_14890);
nand UO_491 (O_491,N_14789,N_14637);
nand UO_492 (O_492,N_14976,N_14419);
nand UO_493 (O_493,N_14978,N_14264);
xor UO_494 (O_494,N_14579,N_14279);
and UO_495 (O_495,N_14879,N_14363);
or UO_496 (O_496,N_14280,N_14910);
xor UO_497 (O_497,N_14535,N_14717);
nand UO_498 (O_498,N_14707,N_14872);
xnor UO_499 (O_499,N_14945,N_14299);
nand UO_500 (O_500,N_14365,N_14904);
nor UO_501 (O_501,N_14935,N_14436);
or UO_502 (O_502,N_14793,N_14573);
xor UO_503 (O_503,N_14748,N_14259);
xnor UO_504 (O_504,N_14392,N_14716);
nor UO_505 (O_505,N_14293,N_14987);
or UO_506 (O_506,N_14771,N_14475);
or UO_507 (O_507,N_14377,N_14999);
nand UO_508 (O_508,N_14656,N_14384);
or UO_509 (O_509,N_14562,N_14444);
or UO_510 (O_510,N_14698,N_14724);
nor UO_511 (O_511,N_14358,N_14478);
xnor UO_512 (O_512,N_14789,N_14404);
nand UO_513 (O_513,N_14520,N_14901);
or UO_514 (O_514,N_14581,N_14398);
nand UO_515 (O_515,N_14377,N_14753);
nand UO_516 (O_516,N_14751,N_14732);
xnor UO_517 (O_517,N_14367,N_14821);
nand UO_518 (O_518,N_14668,N_14835);
nand UO_519 (O_519,N_14254,N_14969);
nor UO_520 (O_520,N_14941,N_14319);
xnor UO_521 (O_521,N_14631,N_14544);
nand UO_522 (O_522,N_14708,N_14891);
nor UO_523 (O_523,N_14842,N_14997);
nor UO_524 (O_524,N_14636,N_14641);
nand UO_525 (O_525,N_14673,N_14625);
or UO_526 (O_526,N_14480,N_14814);
xor UO_527 (O_527,N_14727,N_14901);
or UO_528 (O_528,N_14896,N_14980);
nand UO_529 (O_529,N_14773,N_14805);
xor UO_530 (O_530,N_14772,N_14479);
xnor UO_531 (O_531,N_14372,N_14550);
xor UO_532 (O_532,N_14599,N_14519);
nor UO_533 (O_533,N_14995,N_14927);
nor UO_534 (O_534,N_14457,N_14301);
nor UO_535 (O_535,N_14701,N_14839);
xor UO_536 (O_536,N_14539,N_14304);
nor UO_537 (O_537,N_14433,N_14825);
xor UO_538 (O_538,N_14945,N_14624);
or UO_539 (O_539,N_14257,N_14459);
xor UO_540 (O_540,N_14417,N_14438);
nand UO_541 (O_541,N_14281,N_14922);
xnor UO_542 (O_542,N_14262,N_14861);
or UO_543 (O_543,N_14726,N_14673);
nor UO_544 (O_544,N_14812,N_14736);
or UO_545 (O_545,N_14572,N_14361);
nand UO_546 (O_546,N_14650,N_14971);
and UO_547 (O_547,N_14628,N_14514);
and UO_548 (O_548,N_14510,N_14644);
or UO_549 (O_549,N_14250,N_14507);
and UO_550 (O_550,N_14578,N_14453);
nor UO_551 (O_551,N_14586,N_14306);
nand UO_552 (O_552,N_14399,N_14591);
xnor UO_553 (O_553,N_14558,N_14997);
nand UO_554 (O_554,N_14400,N_14399);
nor UO_555 (O_555,N_14793,N_14657);
and UO_556 (O_556,N_14623,N_14913);
and UO_557 (O_557,N_14994,N_14897);
xor UO_558 (O_558,N_14391,N_14444);
and UO_559 (O_559,N_14444,N_14308);
xnor UO_560 (O_560,N_14285,N_14913);
xor UO_561 (O_561,N_14744,N_14567);
or UO_562 (O_562,N_14359,N_14294);
nand UO_563 (O_563,N_14601,N_14825);
and UO_564 (O_564,N_14272,N_14306);
xor UO_565 (O_565,N_14828,N_14877);
or UO_566 (O_566,N_14924,N_14969);
and UO_567 (O_567,N_14419,N_14545);
nor UO_568 (O_568,N_14560,N_14713);
xnor UO_569 (O_569,N_14936,N_14568);
or UO_570 (O_570,N_14292,N_14645);
xnor UO_571 (O_571,N_14479,N_14954);
and UO_572 (O_572,N_14851,N_14957);
nand UO_573 (O_573,N_14809,N_14601);
nand UO_574 (O_574,N_14991,N_14480);
or UO_575 (O_575,N_14455,N_14540);
nand UO_576 (O_576,N_14732,N_14305);
or UO_577 (O_577,N_14740,N_14689);
and UO_578 (O_578,N_14747,N_14510);
and UO_579 (O_579,N_14348,N_14251);
xor UO_580 (O_580,N_14930,N_14861);
and UO_581 (O_581,N_14922,N_14465);
or UO_582 (O_582,N_14789,N_14802);
nand UO_583 (O_583,N_14721,N_14606);
or UO_584 (O_584,N_14707,N_14548);
nand UO_585 (O_585,N_14845,N_14278);
nand UO_586 (O_586,N_14935,N_14486);
or UO_587 (O_587,N_14348,N_14608);
xor UO_588 (O_588,N_14592,N_14545);
nand UO_589 (O_589,N_14815,N_14853);
and UO_590 (O_590,N_14354,N_14599);
or UO_591 (O_591,N_14688,N_14485);
nor UO_592 (O_592,N_14832,N_14658);
nand UO_593 (O_593,N_14855,N_14263);
nor UO_594 (O_594,N_14665,N_14977);
nor UO_595 (O_595,N_14663,N_14833);
nand UO_596 (O_596,N_14459,N_14295);
and UO_597 (O_597,N_14743,N_14259);
and UO_598 (O_598,N_14285,N_14557);
xor UO_599 (O_599,N_14588,N_14984);
nor UO_600 (O_600,N_14685,N_14554);
xor UO_601 (O_601,N_14526,N_14757);
or UO_602 (O_602,N_14767,N_14800);
nand UO_603 (O_603,N_14275,N_14712);
nand UO_604 (O_604,N_14804,N_14911);
nand UO_605 (O_605,N_14765,N_14536);
and UO_606 (O_606,N_14823,N_14607);
nand UO_607 (O_607,N_14920,N_14648);
or UO_608 (O_608,N_14405,N_14604);
and UO_609 (O_609,N_14428,N_14365);
nor UO_610 (O_610,N_14809,N_14528);
nand UO_611 (O_611,N_14334,N_14543);
nand UO_612 (O_612,N_14496,N_14699);
or UO_613 (O_613,N_14294,N_14741);
or UO_614 (O_614,N_14555,N_14368);
or UO_615 (O_615,N_14682,N_14332);
and UO_616 (O_616,N_14279,N_14540);
and UO_617 (O_617,N_14389,N_14758);
and UO_618 (O_618,N_14781,N_14917);
nand UO_619 (O_619,N_14905,N_14445);
and UO_620 (O_620,N_14872,N_14506);
and UO_621 (O_621,N_14486,N_14374);
or UO_622 (O_622,N_14908,N_14329);
or UO_623 (O_623,N_14424,N_14786);
xor UO_624 (O_624,N_14430,N_14849);
nor UO_625 (O_625,N_14774,N_14612);
nand UO_626 (O_626,N_14388,N_14651);
or UO_627 (O_627,N_14378,N_14847);
and UO_628 (O_628,N_14318,N_14979);
and UO_629 (O_629,N_14972,N_14364);
nor UO_630 (O_630,N_14589,N_14775);
nor UO_631 (O_631,N_14554,N_14504);
nand UO_632 (O_632,N_14939,N_14384);
or UO_633 (O_633,N_14784,N_14645);
nand UO_634 (O_634,N_14792,N_14355);
xor UO_635 (O_635,N_14434,N_14426);
xor UO_636 (O_636,N_14987,N_14470);
xnor UO_637 (O_637,N_14918,N_14527);
nand UO_638 (O_638,N_14359,N_14745);
nand UO_639 (O_639,N_14549,N_14672);
nor UO_640 (O_640,N_14730,N_14619);
nand UO_641 (O_641,N_14503,N_14843);
nor UO_642 (O_642,N_14269,N_14286);
xnor UO_643 (O_643,N_14541,N_14965);
or UO_644 (O_644,N_14989,N_14563);
nand UO_645 (O_645,N_14773,N_14312);
nor UO_646 (O_646,N_14479,N_14758);
nand UO_647 (O_647,N_14349,N_14666);
xnor UO_648 (O_648,N_14384,N_14696);
or UO_649 (O_649,N_14566,N_14959);
xor UO_650 (O_650,N_14501,N_14891);
or UO_651 (O_651,N_14678,N_14836);
or UO_652 (O_652,N_14349,N_14283);
and UO_653 (O_653,N_14846,N_14328);
or UO_654 (O_654,N_14337,N_14286);
xnor UO_655 (O_655,N_14347,N_14546);
xnor UO_656 (O_656,N_14851,N_14483);
xor UO_657 (O_657,N_14815,N_14385);
nor UO_658 (O_658,N_14437,N_14549);
and UO_659 (O_659,N_14601,N_14786);
and UO_660 (O_660,N_14719,N_14774);
nand UO_661 (O_661,N_14319,N_14966);
or UO_662 (O_662,N_14785,N_14722);
nor UO_663 (O_663,N_14967,N_14501);
and UO_664 (O_664,N_14434,N_14481);
xnor UO_665 (O_665,N_14348,N_14729);
or UO_666 (O_666,N_14371,N_14310);
and UO_667 (O_667,N_14556,N_14625);
nor UO_668 (O_668,N_14285,N_14401);
or UO_669 (O_669,N_14876,N_14413);
nor UO_670 (O_670,N_14916,N_14269);
and UO_671 (O_671,N_14370,N_14732);
or UO_672 (O_672,N_14814,N_14823);
nand UO_673 (O_673,N_14645,N_14867);
and UO_674 (O_674,N_14600,N_14467);
nor UO_675 (O_675,N_14337,N_14769);
and UO_676 (O_676,N_14981,N_14432);
or UO_677 (O_677,N_14293,N_14278);
nand UO_678 (O_678,N_14946,N_14391);
and UO_679 (O_679,N_14643,N_14612);
nand UO_680 (O_680,N_14531,N_14588);
or UO_681 (O_681,N_14435,N_14566);
or UO_682 (O_682,N_14259,N_14664);
and UO_683 (O_683,N_14931,N_14812);
nor UO_684 (O_684,N_14370,N_14945);
and UO_685 (O_685,N_14562,N_14513);
xor UO_686 (O_686,N_14485,N_14720);
nand UO_687 (O_687,N_14576,N_14949);
nand UO_688 (O_688,N_14611,N_14738);
nor UO_689 (O_689,N_14931,N_14429);
xor UO_690 (O_690,N_14348,N_14424);
or UO_691 (O_691,N_14664,N_14385);
nand UO_692 (O_692,N_14686,N_14633);
xnor UO_693 (O_693,N_14384,N_14768);
nor UO_694 (O_694,N_14401,N_14827);
or UO_695 (O_695,N_14559,N_14615);
and UO_696 (O_696,N_14911,N_14815);
and UO_697 (O_697,N_14435,N_14562);
and UO_698 (O_698,N_14939,N_14727);
nand UO_699 (O_699,N_14503,N_14894);
nor UO_700 (O_700,N_14756,N_14941);
xor UO_701 (O_701,N_14833,N_14796);
or UO_702 (O_702,N_14757,N_14500);
xor UO_703 (O_703,N_14607,N_14567);
nand UO_704 (O_704,N_14613,N_14651);
or UO_705 (O_705,N_14878,N_14842);
nor UO_706 (O_706,N_14673,N_14974);
and UO_707 (O_707,N_14800,N_14663);
and UO_708 (O_708,N_14329,N_14625);
nand UO_709 (O_709,N_14482,N_14417);
xnor UO_710 (O_710,N_14637,N_14964);
and UO_711 (O_711,N_14466,N_14757);
xor UO_712 (O_712,N_14681,N_14264);
nor UO_713 (O_713,N_14868,N_14620);
or UO_714 (O_714,N_14553,N_14633);
xnor UO_715 (O_715,N_14609,N_14753);
nor UO_716 (O_716,N_14663,N_14587);
and UO_717 (O_717,N_14425,N_14918);
xor UO_718 (O_718,N_14303,N_14845);
nor UO_719 (O_719,N_14544,N_14747);
or UO_720 (O_720,N_14490,N_14820);
xnor UO_721 (O_721,N_14993,N_14980);
or UO_722 (O_722,N_14880,N_14513);
xnor UO_723 (O_723,N_14516,N_14466);
nand UO_724 (O_724,N_14346,N_14872);
xor UO_725 (O_725,N_14274,N_14888);
and UO_726 (O_726,N_14620,N_14592);
xor UO_727 (O_727,N_14725,N_14705);
and UO_728 (O_728,N_14262,N_14518);
nand UO_729 (O_729,N_14265,N_14959);
and UO_730 (O_730,N_14848,N_14594);
nor UO_731 (O_731,N_14279,N_14852);
and UO_732 (O_732,N_14556,N_14371);
nor UO_733 (O_733,N_14690,N_14865);
and UO_734 (O_734,N_14794,N_14620);
nor UO_735 (O_735,N_14793,N_14499);
nor UO_736 (O_736,N_14673,N_14309);
or UO_737 (O_737,N_14664,N_14787);
or UO_738 (O_738,N_14964,N_14991);
or UO_739 (O_739,N_14514,N_14263);
nand UO_740 (O_740,N_14848,N_14843);
xor UO_741 (O_741,N_14782,N_14702);
or UO_742 (O_742,N_14459,N_14724);
or UO_743 (O_743,N_14444,N_14815);
xnor UO_744 (O_744,N_14843,N_14759);
and UO_745 (O_745,N_14636,N_14520);
or UO_746 (O_746,N_14464,N_14424);
nand UO_747 (O_747,N_14456,N_14824);
xnor UO_748 (O_748,N_14314,N_14702);
nor UO_749 (O_749,N_14395,N_14337);
nor UO_750 (O_750,N_14562,N_14442);
xnor UO_751 (O_751,N_14603,N_14994);
nand UO_752 (O_752,N_14354,N_14517);
nor UO_753 (O_753,N_14875,N_14493);
and UO_754 (O_754,N_14526,N_14675);
or UO_755 (O_755,N_14473,N_14260);
or UO_756 (O_756,N_14422,N_14916);
xnor UO_757 (O_757,N_14313,N_14488);
nor UO_758 (O_758,N_14537,N_14692);
or UO_759 (O_759,N_14396,N_14578);
nand UO_760 (O_760,N_14572,N_14553);
or UO_761 (O_761,N_14317,N_14320);
xnor UO_762 (O_762,N_14440,N_14689);
nand UO_763 (O_763,N_14542,N_14598);
xnor UO_764 (O_764,N_14499,N_14478);
nand UO_765 (O_765,N_14893,N_14444);
nor UO_766 (O_766,N_14468,N_14638);
or UO_767 (O_767,N_14713,N_14397);
nor UO_768 (O_768,N_14276,N_14409);
xor UO_769 (O_769,N_14575,N_14337);
nand UO_770 (O_770,N_14462,N_14512);
and UO_771 (O_771,N_14652,N_14847);
nor UO_772 (O_772,N_14654,N_14444);
and UO_773 (O_773,N_14437,N_14927);
and UO_774 (O_774,N_14617,N_14812);
nand UO_775 (O_775,N_14284,N_14583);
xor UO_776 (O_776,N_14575,N_14703);
nand UO_777 (O_777,N_14387,N_14398);
and UO_778 (O_778,N_14916,N_14903);
and UO_779 (O_779,N_14428,N_14921);
and UO_780 (O_780,N_14669,N_14305);
xor UO_781 (O_781,N_14269,N_14764);
xor UO_782 (O_782,N_14359,N_14981);
nor UO_783 (O_783,N_14407,N_14721);
nand UO_784 (O_784,N_14679,N_14439);
and UO_785 (O_785,N_14341,N_14636);
and UO_786 (O_786,N_14917,N_14530);
nand UO_787 (O_787,N_14797,N_14925);
and UO_788 (O_788,N_14358,N_14525);
xor UO_789 (O_789,N_14778,N_14331);
and UO_790 (O_790,N_14442,N_14701);
or UO_791 (O_791,N_14681,N_14288);
nand UO_792 (O_792,N_14453,N_14423);
or UO_793 (O_793,N_14751,N_14611);
and UO_794 (O_794,N_14469,N_14339);
or UO_795 (O_795,N_14971,N_14398);
and UO_796 (O_796,N_14777,N_14522);
nor UO_797 (O_797,N_14665,N_14469);
or UO_798 (O_798,N_14504,N_14730);
xnor UO_799 (O_799,N_14689,N_14263);
nand UO_800 (O_800,N_14905,N_14269);
nand UO_801 (O_801,N_14296,N_14451);
or UO_802 (O_802,N_14478,N_14446);
xnor UO_803 (O_803,N_14891,N_14366);
nand UO_804 (O_804,N_14320,N_14761);
nand UO_805 (O_805,N_14394,N_14710);
nand UO_806 (O_806,N_14724,N_14281);
and UO_807 (O_807,N_14917,N_14581);
nand UO_808 (O_808,N_14585,N_14619);
nand UO_809 (O_809,N_14677,N_14968);
xnor UO_810 (O_810,N_14419,N_14843);
nand UO_811 (O_811,N_14632,N_14808);
nand UO_812 (O_812,N_14853,N_14330);
nor UO_813 (O_813,N_14372,N_14914);
and UO_814 (O_814,N_14329,N_14366);
or UO_815 (O_815,N_14647,N_14366);
nor UO_816 (O_816,N_14525,N_14786);
nor UO_817 (O_817,N_14881,N_14854);
xor UO_818 (O_818,N_14313,N_14654);
or UO_819 (O_819,N_14300,N_14871);
xnor UO_820 (O_820,N_14471,N_14499);
xor UO_821 (O_821,N_14821,N_14429);
xor UO_822 (O_822,N_14623,N_14607);
nand UO_823 (O_823,N_14323,N_14424);
and UO_824 (O_824,N_14505,N_14373);
xor UO_825 (O_825,N_14593,N_14962);
nor UO_826 (O_826,N_14480,N_14294);
or UO_827 (O_827,N_14830,N_14411);
or UO_828 (O_828,N_14840,N_14304);
and UO_829 (O_829,N_14950,N_14660);
and UO_830 (O_830,N_14930,N_14788);
nand UO_831 (O_831,N_14714,N_14400);
nand UO_832 (O_832,N_14522,N_14939);
nor UO_833 (O_833,N_14391,N_14542);
or UO_834 (O_834,N_14659,N_14739);
and UO_835 (O_835,N_14708,N_14416);
or UO_836 (O_836,N_14265,N_14387);
or UO_837 (O_837,N_14549,N_14496);
nand UO_838 (O_838,N_14884,N_14857);
xnor UO_839 (O_839,N_14756,N_14671);
or UO_840 (O_840,N_14924,N_14434);
nor UO_841 (O_841,N_14909,N_14309);
or UO_842 (O_842,N_14399,N_14918);
and UO_843 (O_843,N_14458,N_14387);
nand UO_844 (O_844,N_14605,N_14905);
or UO_845 (O_845,N_14874,N_14398);
nor UO_846 (O_846,N_14865,N_14533);
or UO_847 (O_847,N_14706,N_14452);
xor UO_848 (O_848,N_14668,N_14323);
nor UO_849 (O_849,N_14870,N_14438);
xnor UO_850 (O_850,N_14331,N_14657);
nand UO_851 (O_851,N_14712,N_14439);
nand UO_852 (O_852,N_14490,N_14438);
nand UO_853 (O_853,N_14442,N_14437);
nand UO_854 (O_854,N_14606,N_14521);
xor UO_855 (O_855,N_14558,N_14590);
nand UO_856 (O_856,N_14650,N_14947);
nand UO_857 (O_857,N_14376,N_14987);
xor UO_858 (O_858,N_14779,N_14378);
and UO_859 (O_859,N_14667,N_14273);
and UO_860 (O_860,N_14272,N_14782);
xor UO_861 (O_861,N_14333,N_14416);
nor UO_862 (O_862,N_14521,N_14344);
and UO_863 (O_863,N_14274,N_14948);
or UO_864 (O_864,N_14316,N_14966);
nor UO_865 (O_865,N_14282,N_14292);
nand UO_866 (O_866,N_14602,N_14710);
nand UO_867 (O_867,N_14747,N_14284);
nor UO_868 (O_868,N_14658,N_14787);
xor UO_869 (O_869,N_14800,N_14503);
xor UO_870 (O_870,N_14441,N_14364);
or UO_871 (O_871,N_14291,N_14335);
nor UO_872 (O_872,N_14497,N_14455);
nand UO_873 (O_873,N_14391,N_14528);
xnor UO_874 (O_874,N_14885,N_14657);
xnor UO_875 (O_875,N_14386,N_14264);
nand UO_876 (O_876,N_14744,N_14496);
nand UO_877 (O_877,N_14445,N_14893);
and UO_878 (O_878,N_14366,N_14926);
nand UO_879 (O_879,N_14699,N_14849);
and UO_880 (O_880,N_14261,N_14671);
nor UO_881 (O_881,N_14333,N_14362);
or UO_882 (O_882,N_14747,N_14945);
nor UO_883 (O_883,N_14650,N_14430);
and UO_884 (O_884,N_14395,N_14475);
nor UO_885 (O_885,N_14937,N_14835);
or UO_886 (O_886,N_14925,N_14658);
nand UO_887 (O_887,N_14425,N_14585);
xor UO_888 (O_888,N_14891,N_14881);
and UO_889 (O_889,N_14932,N_14752);
nand UO_890 (O_890,N_14511,N_14714);
xor UO_891 (O_891,N_14949,N_14495);
xnor UO_892 (O_892,N_14309,N_14456);
or UO_893 (O_893,N_14549,N_14595);
nor UO_894 (O_894,N_14822,N_14430);
nand UO_895 (O_895,N_14758,N_14417);
and UO_896 (O_896,N_14275,N_14603);
xnor UO_897 (O_897,N_14303,N_14599);
nor UO_898 (O_898,N_14288,N_14375);
nor UO_899 (O_899,N_14930,N_14324);
nor UO_900 (O_900,N_14990,N_14301);
nand UO_901 (O_901,N_14624,N_14664);
or UO_902 (O_902,N_14483,N_14485);
xor UO_903 (O_903,N_14866,N_14255);
xnor UO_904 (O_904,N_14454,N_14788);
and UO_905 (O_905,N_14939,N_14600);
or UO_906 (O_906,N_14820,N_14761);
nand UO_907 (O_907,N_14252,N_14699);
and UO_908 (O_908,N_14713,N_14742);
or UO_909 (O_909,N_14761,N_14393);
nor UO_910 (O_910,N_14388,N_14447);
nor UO_911 (O_911,N_14370,N_14901);
nand UO_912 (O_912,N_14618,N_14351);
nand UO_913 (O_913,N_14498,N_14779);
nor UO_914 (O_914,N_14410,N_14993);
or UO_915 (O_915,N_14470,N_14909);
nand UO_916 (O_916,N_14402,N_14276);
xnor UO_917 (O_917,N_14256,N_14742);
and UO_918 (O_918,N_14912,N_14671);
xor UO_919 (O_919,N_14906,N_14635);
nor UO_920 (O_920,N_14622,N_14326);
or UO_921 (O_921,N_14252,N_14721);
and UO_922 (O_922,N_14385,N_14359);
or UO_923 (O_923,N_14667,N_14856);
nand UO_924 (O_924,N_14858,N_14904);
and UO_925 (O_925,N_14315,N_14440);
xor UO_926 (O_926,N_14513,N_14868);
xnor UO_927 (O_927,N_14950,N_14597);
and UO_928 (O_928,N_14490,N_14478);
or UO_929 (O_929,N_14858,N_14363);
xnor UO_930 (O_930,N_14701,N_14560);
or UO_931 (O_931,N_14630,N_14409);
and UO_932 (O_932,N_14302,N_14534);
nand UO_933 (O_933,N_14939,N_14360);
or UO_934 (O_934,N_14959,N_14770);
nor UO_935 (O_935,N_14400,N_14334);
nor UO_936 (O_936,N_14634,N_14375);
or UO_937 (O_937,N_14354,N_14761);
and UO_938 (O_938,N_14644,N_14746);
or UO_939 (O_939,N_14696,N_14755);
or UO_940 (O_940,N_14928,N_14690);
nand UO_941 (O_941,N_14319,N_14842);
xor UO_942 (O_942,N_14735,N_14263);
nand UO_943 (O_943,N_14937,N_14884);
nor UO_944 (O_944,N_14710,N_14307);
or UO_945 (O_945,N_14921,N_14535);
or UO_946 (O_946,N_14339,N_14351);
xnor UO_947 (O_947,N_14942,N_14434);
or UO_948 (O_948,N_14591,N_14376);
or UO_949 (O_949,N_14618,N_14982);
and UO_950 (O_950,N_14457,N_14362);
or UO_951 (O_951,N_14804,N_14734);
and UO_952 (O_952,N_14930,N_14541);
and UO_953 (O_953,N_14951,N_14648);
xor UO_954 (O_954,N_14803,N_14595);
xor UO_955 (O_955,N_14628,N_14256);
nor UO_956 (O_956,N_14862,N_14494);
or UO_957 (O_957,N_14252,N_14410);
nor UO_958 (O_958,N_14782,N_14775);
or UO_959 (O_959,N_14515,N_14853);
or UO_960 (O_960,N_14653,N_14743);
nand UO_961 (O_961,N_14868,N_14341);
nor UO_962 (O_962,N_14251,N_14972);
nor UO_963 (O_963,N_14715,N_14840);
and UO_964 (O_964,N_14739,N_14273);
and UO_965 (O_965,N_14949,N_14630);
nand UO_966 (O_966,N_14836,N_14360);
nor UO_967 (O_967,N_14994,N_14385);
nand UO_968 (O_968,N_14327,N_14994);
or UO_969 (O_969,N_14547,N_14255);
xnor UO_970 (O_970,N_14536,N_14942);
nand UO_971 (O_971,N_14731,N_14954);
xor UO_972 (O_972,N_14323,N_14787);
and UO_973 (O_973,N_14580,N_14390);
and UO_974 (O_974,N_14412,N_14861);
or UO_975 (O_975,N_14392,N_14455);
nand UO_976 (O_976,N_14373,N_14496);
xnor UO_977 (O_977,N_14687,N_14284);
xnor UO_978 (O_978,N_14732,N_14639);
and UO_979 (O_979,N_14839,N_14442);
and UO_980 (O_980,N_14355,N_14755);
and UO_981 (O_981,N_14797,N_14765);
xnor UO_982 (O_982,N_14309,N_14895);
nand UO_983 (O_983,N_14324,N_14374);
nor UO_984 (O_984,N_14715,N_14796);
nand UO_985 (O_985,N_14913,N_14276);
xnor UO_986 (O_986,N_14571,N_14935);
xor UO_987 (O_987,N_14828,N_14288);
xor UO_988 (O_988,N_14504,N_14572);
nor UO_989 (O_989,N_14447,N_14777);
nand UO_990 (O_990,N_14791,N_14424);
xor UO_991 (O_991,N_14533,N_14291);
or UO_992 (O_992,N_14945,N_14929);
or UO_993 (O_993,N_14381,N_14548);
nor UO_994 (O_994,N_14477,N_14409);
nand UO_995 (O_995,N_14484,N_14780);
and UO_996 (O_996,N_14946,N_14380);
or UO_997 (O_997,N_14627,N_14482);
nand UO_998 (O_998,N_14723,N_14260);
nor UO_999 (O_999,N_14703,N_14373);
or UO_1000 (O_1000,N_14595,N_14981);
nor UO_1001 (O_1001,N_14476,N_14955);
or UO_1002 (O_1002,N_14879,N_14517);
nand UO_1003 (O_1003,N_14678,N_14363);
nand UO_1004 (O_1004,N_14305,N_14807);
and UO_1005 (O_1005,N_14462,N_14367);
nand UO_1006 (O_1006,N_14346,N_14456);
xnor UO_1007 (O_1007,N_14735,N_14952);
xnor UO_1008 (O_1008,N_14879,N_14531);
or UO_1009 (O_1009,N_14775,N_14391);
nor UO_1010 (O_1010,N_14319,N_14831);
xor UO_1011 (O_1011,N_14548,N_14413);
nor UO_1012 (O_1012,N_14696,N_14628);
xor UO_1013 (O_1013,N_14582,N_14322);
xor UO_1014 (O_1014,N_14333,N_14280);
xor UO_1015 (O_1015,N_14333,N_14526);
nor UO_1016 (O_1016,N_14983,N_14428);
nand UO_1017 (O_1017,N_14321,N_14564);
nor UO_1018 (O_1018,N_14480,N_14860);
xor UO_1019 (O_1019,N_14742,N_14421);
and UO_1020 (O_1020,N_14548,N_14509);
and UO_1021 (O_1021,N_14719,N_14313);
nor UO_1022 (O_1022,N_14672,N_14907);
nor UO_1023 (O_1023,N_14533,N_14563);
or UO_1024 (O_1024,N_14461,N_14303);
or UO_1025 (O_1025,N_14888,N_14485);
and UO_1026 (O_1026,N_14702,N_14811);
and UO_1027 (O_1027,N_14946,N_14948);
or UO_1028 (O_1028,N_14513,N_14673);
xnor UO_1029 (O_1029,N_14907,N_14310);
and UO_1030 (O_1030,N_14277,N_14462);
nor UO_1031 (O_1031,N_14810,N_14449);
xnor UO_1032 (O_1032,N_14961,N_14308);
and UO_1033 (O_1033,N_14787,N_14406);
and UO_1034 (O_1034,N_14290,N_14944);
and UO_1035 (O_1035,N_14647,N_14878);
nand UO_1036 (O_1036,N_14314,N_14518);
and UO_1037 (O_1037,N_14818,N_14756);
nor UO_1038 (O_1038,N_14339,N_14927);
nor UO_1039 (O_1039,N_14802,N_14756);
nand UO_1040 (O_1040,N_14872,N_14788);
and UO_1041 (O_1041,N_14768,N_14473);
nor UO_1042 (O_1042,N_14938,N_14656);
or UO_1043 (O_1043,N_14497,N_14891);
xnor UO_1044 (O_1044,N_14412,N_14417);
nand UO_1045 (O_1045,N_14517,N_14993);
or UO_1046 (O_1046,N_14251,N_14984);
or UO_1047 (O_1047,N_14696,N_14898);
xor UO_1048 (O_1048,N_14591,N_14576);
or UO_1049 (O_1049,N_14681,N_14525);
or UO_1050 (O_1050,N_14513,N_14300);
nor UO_1051 (O_1051,N_14466,N_14493);
or UO_1052 (O_1052,N_14374,N_14272);
nand UO_1053 (O_1053,N_14911,N_14953);
or UO_1054 (O_1054,N_14459,N_14253);
and UO_1055 (O_1055,N_14533,N_14735);
nand UO_1056 (O_1056,N_14251,N_14373);
and UO_1057 (O_1057,N_14772,N_14744);
nand UO_1058 (O_1058,N_14821,N_14690);
xor UO_1059 (O_1059,N_14849,N_14921);
xor UO_1060 (O_1060,N_14880,N_14439);
nand UO_1061 (O_1061,N_14920,N_14368);
nand UO_1062 (O_1062,N_14508,N_14351);
and UO_1063 (O_1063,N_14855,N_14646);
nor UO_1064 (O_1064,N_14916,N_14595);
nor UO_1065 (O_1065,N_14800,N_14460);
or UO_1066 (O_1066,N_14784,N_14813);
or UO_1067 (O_1067,N_14673,N_14723);
nor UO_1068 (O_1068,N_14572,N_14458);
nor UO_1069 (O_1069,N_14741,N_14369);
nor UO_1070 (O_1070,N_14420,N_14781);
and UO_1071 (O_1071,N_14577,N_14790);
nand UO_1072 (O_1072,N_14822,N_14714);
or UO_1073 (O_1073,N_14537,N_14280);
nor UO_1074 (O_1074,N_14930,N_14587);
and UO_1075 (O_1075,N_14614,N_14523);
nand UO_1076 (O_1076,N_14685,N_14459);
nand UO_1077 (O_1077,N_14451,N_14371);
or UO_1078 (O_1078,N_14270,N_14505);
or UO_1079 (O_1079,N_14508,N_14511);
nand UO_1080 (O_1080,N_14538,N_14409);
nand UO_1081 (O_1081,N_14863,N_14991);
and UO_1082 (O_1082,N_14971,N_14556);
nor UO_1083 (O_1083,N_14269,N_14824);
nand UO_1084 (O_1084,N_14615,N_14337);
nand UO_1085 (O_1085,N_14774,N_14459);
or UO_1086 (O_1086,N_14680,N_14263);
xnor UO_1087 (O_1087,N_14876,N_14529);
nor UO_1088 (O_1088,N_14766,N_14533);
nand UO_1089 (O_1089,N_14921,N_14612);
nand UO_1090 (O_1090,N_14399,N_14989);
and UO_1091 (O_1091,N_14903,N_14985);
nor UO_1092 (O_1092,N_14523,N_14377);
and UO_1093 (O_1093,N_14376,N_14344);
nand UO_1094 (O_1094,N_14855,N_14584);
nand UO_1095 (O_1095,N_14472,N_14862);
or UO_1096 (O_1096,N_14364,N_14486);
and UO_1097 (O_1097,N_14435,N_14906);
nor UO_1098 (O_1098,N_14316,N_14280);
nand UO_1099 (O_1099,N_14296,N_14624);
or UO_1100 (O_1100,N_14501,N_14699);
or UO_1101 (O_1101,N_14498,N_14786);
and UO_1102 (O_1102,N_14499,N_14261);
and UO_1103 (O_1103,N_14926,N_14678);
or UO_1104 (O_1104,N_14632,N_14276);
nand UO_1105 (O_1105,N_14884,N_14409);
nand UO_1106 (O_1106,N_14961,N_14874);
or UO_1107 (O_1107,N_14457,N_14384);
and UO_1108 (O_1108,N_14997,N_14665);
nor UO_1109 (O_1109,N_14714,N_14394);
nor UO_1110 (O_1110,N_14531,N_14537);
nor UO_1111 (O_1111,N_14436,N_14600);
nor UO_1112 (O_1112,N_14317,N_14696);
or UO_1113 (O_1113,N_14469,N_14759);
nor UO_1114 (O_1114,N_14631,N_14935);
xor UO_1115 (O_1115,N_14646,N_14280);
xnor UO_1116 (O_1116,N_14907,N_14454);
nor UO_1117 (O_1117,N_14871,N_14579);
or UO_1118 (O_1118,N_14932,N_14941);
or UO_1119 (O_1119,N_14572,N_14390);
nand UO_1120 (O_1120,N_14293,N_14809);
or UO_1121 (O_1121,N_14307,N_14612);
and UO_1122 (O_1122,N_14649,N_14354);
xnor UO_1123 (O_1123,N_14451,N_14523);
xor UO_1124 (O_1124,N_14760,N_14557);
xor UO_1125 (O_1125,N_14895,N_14498);
nand UO_1126 (O_1126,N_14633,N_14350);
and UO_1127 (O_1127,N_14348,N_14257);
nand UO_1128 (O_1128,N_14547,N_14957);
nand UO_1129 (O_1129,N_14902,N_14463);
xor UO_1130 (O_1130,N_14306,N_14484);
and UO_1131 (O_1131,N_14451,N_14390);
or UO_1132 (O_1132,N_14552,N_14530);
and UO_1133 (O_1133,N_14985,N_14409);
nand UO_1134 (O_1134,N_14846,N_14549);
nand UO_1135 (O_1135,N_14273,N_14821);
nand UO_1136 (O_1136,N_14388,N_14565);
xor UO_1137 (O_1137,N_14733,N_14270);
xnor UO_1138 (O_1138,N_14855,N_14628);
or UO_1139 (O_1139,N_14399,N_14932);
or UO_1140 (O_1140,N_14440,N_14680);
nand UO_1141 (O_1141,N_14977,N_14697);
nor UO_1142 (O_1142,N_14543,N_14456);
nor UO_1143 (O_1143,N_14541,N_14919);
nor UO_1144 (O_1144,N_14834,N_14350);
and UO_1145 (O_1145,N_14676,N_14445);
nor UO_1146 (O_1146,N_14762,N_14381);
nor UO_1147 (O_1147,N_14994,N_14370);
or UO_1148 (O_1148,N_14670,N_14479);
xor UO_1149 (O_1149,N_14274,N_14739);
or UO_1150 (O_1150,N_14638,N_14978);
xnor UO_1151 (O_1151,N_14348,N_14589);
xnor UO_1152 (O_1152,N_14953,N_14320);
xnor UO_1153 (O_1153,N_14902,N_14401);
nand UO_1154 (O_1154,N_14546,N_14705);
nand UO_1155 (O_1155,N_14553,N_14518);
and UO_1156 (O_1156,N_14917,N_14894);
or UO_1157 (O_1157,N_14560,N_14347);
nand UO_1158 (O_1158,N_14927,N_14348);
xor UO_1159 (O_1159,N_14734,N_14690);
xor UO_1160 (O_1160,N_14336,N_14949);
and UO_1161 (O_1161,N_14635,N_14790);
xor UO_1162 (O_1162,N_14459,N_14378);
or UO_1163 (O_1163,N_14646,N_14539);
nand UO_1164 (O_1164,N_14695,N_14889);
and UO_1165 (O_1165,N_14967,N_14390);
nor UO_1166 (O_1166,N_14392,N_14619);
or UO_1167 (O_1167,N_14568,N_14652);
and UO_1168 (O_1168,N_14718,N_14941);
or UO_1169 (O_1169,N_14847,N_14498);
nand UO_1170 (O_1170,N_14483,N_14635);
nand UO_1171 (O_1171,N_14681,N_14769);
or UO_1172 (O_1172,N_14970,N_14601);
nor UO_1173 (O_1173,N_14334,N_14564);
nor UO_1174 (O_1174,N_14362,N_14801);
nand UO_1175 (O_1175,N_14285,N_14748);
xnor UO_1176 (O_1176,N_14630,N_14344);
xor UO_1177 (O_1177,N_14356,N_14301);
and UO_1178 (O_1178,N_14626,N_14612);
or UO_1179 (O_1179,N_14719,N_14696);
nor UO_1180 (O_1180,N_14360,N_14492);
nand UO_1181 (O_1181,N_14271,N_14485);
nand UO_1182 (O_1182,N_14392,N_14833);
or UO_1183 (O_1183,N_14481,N_14845);
nor UO_1184 (O_1184,N_14443,N_14608);
and UO_1185 (O_1185,N_14375,N_14633);
nand UO_1186 (O_1186,N_14921,N_14407);
and UO_1187 (O_1187,N_14934,N_14594);
or UO_1188 (O_1188,N_14827,N_14508);
xnor UO_1189 (O_1189,N_14796,N_14620);
nor UO_1190 (O_1190,N_14923,N_14974);
xnor UO_1191 (O_1191,N_14937,N_14692);
or UO_1192 (O_1192,N_14403,N_14552);
nor UO_1193 (O_1193,N_14718,N_14996);
and UO_1194 (O_1194,N_14772,N_14588);
and UO_1195 (O_1195,N_14946,N_14770);
xnor UO_1196 (O_1196,N_14258,N_14844);
xnor UO_1197 (O_1197,N_14805,N_14346);
or UO_1198 (O_1198,N_14675,N_14895);
nor UO_1199 (O_1199,N_14329,N_14775);
xor UO_1200 (O_1200,N_14770,N_14653);
xor UO_1201 (O_1201,N_14441,N_14788);
or UO_1202 (O_1202,N_14286,N_14404);
nand UO_1203 (O_1203,N_14558,N_14630);
xor UO_1204 (O_1204,N_14896,N_14695);
nor UO_1205 (O_1205,N_14418,N_14938);
nor UO_1206 (O_1206,N_14539,N_14779);
xnor UO_1207 (O_1207,N_14671,N_14624);
and UO_1208 (O_1208,N_14403,N_14584);
and UO_1209 (O_1209,N_14918,N_14468);
or UO_1210 (O_1210,N_14253,N_14904);
nor UO_1211 (O_1211,N_14752,N_14302);
or UO_1212 (O_1212,N_14430,N_14351);
nand UO_1213 (O_1213,N_14758,N_14258);
and UO_1214 (O_1214,N_14529,N_14572);
and UO_1215 (O_1215,N_14594,N_14401);
and UO_1216 (O_1216,N_14521,N_14363);
xnor UO_1217 (O_1217,N_14889,N_14646);
or UO_1218 (O_1218,N_14783,N_14647);
xor UO_1219 (O_1219,N_14853,N_14406);
xnor UO_1220 (O_1220,N_14533,N_14340);
or UO_1221 (O_1221,N_14568,N_14547);
xor UO_1222 (O_1222,N_14972,N_14300);
xnor UO_1223 (O_1223,N_14491,N_14441);
and UO_1224 (O_1224,N_14471,N_14986);
nor UO_1225 (O_1225,N_14304,N_14604);
or UO_1226 (O_1226,N_14968,N_14311);
and UO_1227 (O_1227,N_14399,N_14820);
or UO_1228 (O_1228,N_14956,N_14489);
xor UO_1229 (O_1229,N_14557,N_14845);
or UO_1230 (O_1230,N_14379,N_14775);
nand UO_1231 (O_1231,N_14796,N_14451);
and UO_1232 (O_1232,N_14867,N_14961);
nand UO_1233 (O_1233,N_14357,N_14740);
and UO_1234 (O_1234,N_14504,N_14536);
or UO_1235 (O_1235,N_14935,N_14574);
or UO_1236 (O_1236,N_14868,N_14325);
xnor UO_1237 (O_1237,N_14371,N_14828);
or UO_1238 (O_1238,N_14749,N_14641);
or UO_1239 (O_1239,N_14692,N_14440);
nand UO_1240 (O_1240,N_14722,N_14814);
or UO_1241 (O_1241,N_14379,N_14792);
and UO_1242 (O_1242,N_14577,N_14823);
or UO_1243 (O_1243,N_14977,N_14810);
or UO_1244 (O_1244,N_14362,N_14848);
xor UO_1245 (O_1245,N_14366,N_14853);
xnor UO_1246 (O_1246,N_14295,N_14938);
or UO_1247 (O_1247,N_14259,N_14285);
nand UO_1248 (O_1248,N_14483,N_14779);
xor UO_1249 (O_1249,N_14389,N_14900);
xnor UO_1250 (O_1250,N_14513,N_14934);
nand UO_1251 (O_1251,N_14530,N_14942);
nand UO_1252 (O_1252,N_14772,N_14620);
nor UO_1253 (O_1253,N_14788,N_14821);
or UO_1254 (O_1254,N_14944,N_14840);
nand UO_1255 (O_1255,N_14545,N_14461);
and UO_1256 (O_1256,N_14447,N_14629);
or UO_1257 (O_1257,N_14731,N_14319);
and UO_1258 (O_1258,N_14503,N_14340);
xnor UO_1259 (O_1259,N_14996,N_14253);
nand UO_1260 (O_1260,N_14639,N_14597);
nand UO_1261 (O_1261,N_14355,N_14585);
nand UO_1262 (O_1262,N_14423,N_14502);
and UO_1263 (O_1263,N_14815,N_14602);
nand UO_1264 (O_1264,N_14559,N_14560);
nor UO_1265 (O_1265,N_14953,N_14430);
nor UO_1266 (O_1266,N_14617,N_14272);
and UO_1267 (O_1267,N_14525,N_14615);
or UO_1268 (O_1268,N_14283,N_14298);
nand UO_1269 (O_1269,N_14612,N_14769);
or UO_1270 (O_1270,N_14966,N_14938);
nor UO_1271 (O_1271,N_14369,N_14846);
and UO_1272 (O_1272,N_14738,N_14835);
and UO_1273 (O_1273,N_14710,N_14980);
or UO_1274 (O_1274,N_14591,N_14666);
or UO_1275 (O_1275,N_14923,N_14331);
nand UO_1276 (O_1276,N_14527,N_14904);
or UO_1277 (O_1277,N_14603,N_14841);
and UO_1278 (O_1278,N_14306,N_14749);
and UO_1279 (O_1279,N_14314,N_14499);
and UO_1280 (O_1280,N_14984,N_14627);
nand UO_1281 (O_1281,N_14333,N_14505);
nand UO_1282 (O_1282,N_14641,N_14740);
and UO_1283 (O_1283,N_14477,N_14708);
or UO_1284 (O_1284,N_14409,N_14929);
and UO_1285 (O_1285,N_14877,N_14865);
or UO_1286 (O_1286,N_14641,N_14795);
xor UO_1287 (O_1287,N_14374,N_14909);
or UO_1288 (O_1288,N_14632,N_14596);
nor UO_1289 (O_1289,N_14574,N_14266);
nor UO_1290 (O_1290,N_14495,N_14666);
nand UO_1291 (O_1291,N_14576,N_14424);
nand UO_1292 (O_1292,N_14269,N_14621);
nand UO_1293 (O_1293,N_14604,N_14664);
xnor UO_1294 (O_1294,N_14954,N_14959);
or UO_1295 (O_1295,N_14865,N_14301);
and UO_1296 (O_1296,N_14987,N_14997);
or UO_1297 (O_1297,N_14959,N_14846);
or UO_1298 (O_1298,N_14499,N_14285);
nand UO_1299 (O_1299,N_14850,N_14975);
nand UO_1300 (O_1300,N_14911,N_14463);
nand UO_1301 (O_1301,N_14791,N_14764);
nand UO_1302 (O_1302,N_14519,N_14677);
xnor UO_1303 (O_1303,N_14630,N_14868);
nand UO_1304 (O_1304,N_14943,N_14307);
or UO_1305 (O_1305,N_14836,N_14698);
nand UO_1306 (O_1306,N_14709,N_14500);
or UO_1307 (O_1307,N_14481,N_14761);
and UO_1308 (O_1308,N_14672,N_14368);
nand UO_1309 (O_1309,N_14579,N_14605);
and UO_1310 (O_1310,N_14558,N_14632);
or UO_1311 (O_1311,N_14812,N_14830);
and UO_1312 (O_1312,N_14607,N_14712);
and UO_1313 (O_1313,N_14856,N_14556);
or UO_1314 (O_1314,N_14722,N_14948);
or UO_1315 (O_1315,N_14532,N_14457);
nor UO_1316 (O_1316,N_14996,N_14606);
nand UO_1317 (O_1317,N_14998,N_14812);
or UO_1318 (O_1318,N_14549,N_14999);
nand UO_1319 (O_1319,N_14866,N_14863);
nand UO_1320 (O_1320,N_14361,N_14870);
and UO_1321 (O_1321,N_14835,N_14398);
nand UO_1322 (O_1322,N_14940,N_14693);
xnor UO_1323 (O_1323,N_14408,N_14981);
nor UO_1324 (O_1324,N_14644,N_14615);
and UO_1325 (O_1325,N_14540,N_14942);
nor UO_1326 (O_1326,N_14518,N_14503);
or UO_1327 (O_1327,N_14907,N_14531);
nor UO_1328 (O_1328,N_14523,N_14635);
nand UO_1329 (O_1329,N_14906,N_14340);
nand UO_1330 (O_1330,N_14501,N_14596);
nand UO_1331 (O_1331,N_14885,N_14978);
nand UO_1332 (O_1332,N_14343,N_14790);
xnor UO_1333 (O_1333,N_14577,N_14821);
nand UO_1334 (O_1334,N_14745,N_14878);
or UO_1335 (O_1335,N_14966,N_14774);
xnor UO_1336 (O_1336,N_14256,N_14461);
xor UO_1337 (O_1337,N_14496,N_14798);
and UO_1338 (O_1338,N_14919,N_14892);
xnor UO_1339 (O_1339,N_14636,N_14349);
xnor UO_1340 (O_1340,N_14257,N_14691);
xor UO_1341 (O_1341,N_14691,N_14419);
or UO_1342 (O_1342,N_14656,N_14839);
xnor UO_1343 (O_1343,N_14754,N_14388);
or UO_1344 (O_1344,N_14863,N_14793);
and UO_1345 (O_1345,N_14709,N_14446);
nor UO_1346 (O_1346,N_14451,N_14705);
nor UO_1347 (O_1347,N_14549,N_14625);
or UO_1348 (O_1348,N_14867,N_14306);
nor UO_1349 (O_1349,N_14987,N_14901);
xnor UO_1350 (O_1350,N_14366,N_14887);
nor UO_1351 (O_1351,N_14295,N_14268);
xor UO_1352 (O_1352,N_14422,N_14666);
and UO_1353 (O_1353,N_14320,N_14586);
or UO_1354 (O_1354,N_14940,N_14498);
nand UO_1355 (O_1355,N_14344,N_14940);
nor UO_1356 (O_1356,N_14396,N_14586);
and UO_1357 (O_1357,N_14716,N_14905);
nor UO_1358 (O_1358,N_14482,N_14328);
nor UO_1359 (O_1359,N_14712,N_14909);
or UO_1360 (O_1360,N_14707,N_14905);
or UO_1361 (O_1361,N_14737,N_14545);
or UO_1362 (O_1362,N_14845,N_14812);
nand UO_1363 (O_1363,N_14537,N_14814);
or UO_1364 (O_1364,N_14723,N_14512);
xor UO_1365 (O_1365,N_14567,N_14765);
and UO_1366 (O_1366,N_14932,N_14905);
xor UO_1367 (O_1367,N_14659,N_14410);
xnor UO_1368 (O_1368,N_14803,N_14928);
or UO_1369 (O_1369,N_14586,N_14565);
and UO_1370 (O_1370,N_14944,N_14830);
xor UO_1371 (O_1371,N_14607,N_14945);
nor UO_1372 (O_1372,N_14977,N_14822);
or UO_1373 (O_1373,N_14873,N_14832);
nand UO_1374 (O_1374,N_14265,N_14699);
and UO_1375 (O_1375,N_14377,N_14797);
and UO_1376 (O_1376,N_14638,N_14948);
or UO_1377 (O_1377,N_14441,N_14998);
nand UO_1378 (O_1378,N_14599,N_14880);
nand UO_1379 (O_1379,N_14523,N_14469);
nand UO_1380 (O_1380,N_14955,N_14842);
xnor UO_1381 (O_1381,N_14722,N_14854);
or UO_1382 (O_1382,N_14616,N_14614);
nor UO_1383 (O_1383,N_14864,N_14816);
and UO_1384 (O_1384,N_14413,N_14394);
xor UO_1385 (O_1385,N_14957,N_14368);
or UO_1386 (O_1386,N_14773,N_14438);
and UO_1387 (O_1387,N_14660,N_14749);
and UO_1388 (O_1388,N_14966,N_14704);
nand UO_1389 (O_1389,N_14896,N_14655);
nor UO_1390 (O_1390,N_14560,N_14578);
nor UO_1391 (O_1391,N_14788,N_14420);
nor UO_1392 (O_1392,N_14657,N_14960);
xor UO_1393 (O_1393,N_14764,N_14266);
nand UO_1394 (O_1394,N_14560,N_14811);
or UO_1395 (O_1395,N_14895,N_14298);
and UO_1396 (O_1396,N_14587,N_14280);
nand UO_1397 (O_1397,N_14426,N_14269);
xnor UO_1398 (O_1398,N_14385,N_14981);
nand UO_1399 (O_1399,N_14756,N_14400);
nand UO_1400 (O_1400,N_14337,N_14268);
nor UO_1401 (O_1401,N_14722,N_14587);
and UO_1402 (O_1402,N_14725,N_14383);
xor UO_1403 (O_1403,N_14616,N_14417);
and UO_1404 (O_1404,N_14929,N_14960);
nor UO_1405 (O_1405,N_14829,N_14742);
xnor UO_1406 (O_1406,N_14530,N_14970);
or UO_1407 (O_1407,N_14998,N_14944);
and UO_1408 (O_1408,N_14458,N_14867);
or UO_1409 (O_1409,N_14318,N_14502);
or UO_1410 (O_1410,N_14484,N_14338);
or UO_1411 (O_1411,N_14462,N_14785);
and UO_1412 (O_1412,N_14858,N_14452);
and UO_1413 (O_1413,N_14934,N_14698);
or UO_1414 (O_1414,N_14270,N_14601);
and UO_1415 (O_1415,N_14840,N_14973);
and UO_1416 (O_1416,N_14715,N_14874);
nand UO_1417 (O_1417,N_14910,N_14333);
and UO_1418 (O_1418,N_14754,N_14626);
nor UO_1419 (O_1419,N_14589,N_14394);
and UO_1420 (O_1420,N_14675,N_14372);
xor UO_1421 (O_1421,N_14670,N_14994);
nand UO_1422 (O_1422,N_14710,N_14659);
nor UO_1423 (O_1423,N_14842,N_14487);
or UO_1424 (O_1424,N_14354,N_14258);
and UO_1425 (O_1425,N_14619,N_14360);
nor UO_1426 (O_1426,N_14731,N_14470);
and UO_1427 (O_1427,N_14362,N_14846);
nand UO_1428 (O_1428,N_14519,N_14970);
and UO_1429 (O_1429,N_14585,N_14640);
nor UO_1430 (O_1430,N_14883,N_14399);
or UO_1431 (O_1431,N_14478,N_14252);
nor UO_1432 (O_1432,N_14584,N_14857);
xor UO_1433 (O_1433,N_14656,N_14481);
xnor UO_1434 (O_1434,N_14531,N_14853);
and UO_1435 (O_1435,N_14512,N_14412);
xnor UO_1436 (O_1436,N_14925,N_14259);
nand UO_1437 (O_1437,N_14419,N_14400);
and UO_1438 (O_1438,N_14570,N_14887);
xor UO_1439 (O_1439,N_14634,N_14250);
xor UO_1440 (O_1440,N_14664,N_14751);
xnor UO_1441 (O_1441,N_14986,N_14745);
nor UO_1442 (O_1442,N_14434,N_14651);
or UO_1443 (O_1443,N_14289,N_14702);
nand UO_1444 (O_1444,N_14608,N_14350);
or UO_1445 (O_1445,N_14674,N_14814);
nor UO_1446 (O_1446,N_14579,N_14943);
nor UO_1447 (O_1447,N_14373,N_14635);
or UO_1448 (O_1448,N_14340,N_14506);
nand UO_1449 (O_1449,N_14763,N_14437);
or UO_1450 (O_1450,N_14605,N_14658);
xnor UO_1451 (O_1451,N_14462,N_14378);
or UO_1452 (O_1452,N_14268,N_14402);
nor UO_1453 (O_1453,N_14316,N_14636);
nor UO_1454 (O_1454,N_14328,N_14490);
xnor UO_1455 (O_1455,N_14445,N_14417);
and UO_1456 (O_1456,N_14334,N_14818);
and UO_1457 (O_1457,N_14784,N_14531);
or UO_1458 (O_1458,N_14339,N_14424);
xnor UO_1459 (O_1459,N_14748,N_14606);
nor UO_1460 (O_1460,N_14443,N_14902);
and UO_1461 (O_1461,N_14921,N_14453);
or UO_1462 (O_1462,N_14863,N_14338);
nand UO_1463 (O_1463,N_14418,N_14425);
nand UO_1464 (O_1464,N_14985,N_14690);
or UO_1465 (O_1465,N_14867,N_14436);
and UO_1466 (O_1466,N_14757,N_14771);
nand UO_1467 (O_1467,N_14713,N_14991);
xor UO_1468 (O_1468,N_14723,N_14717);
nand UO_1469 (O_1469,N_14470,N_14498);
xnor UO_1470 (O_1470,N_14704,N_14940);
nand UO_1471 (O_1471,N_14531,N_14991);
and UO_1472 (O_1472,N_14398,N_14597);
nand UO_1473 (O_1473,N_14678,N_14834);
xor UO_1474 (O_1474,N_14442,N_14834);
nand UO_1475 (O_1475,N_14726,N_14288);
nor UO_1476 (O_1476,N_14342,N_14254);
xnor UO_1477 (O_1477,N_14417,N_14408);
xor UO_1478 (O_1478,N_14419,N_14713);
and UO_1479 (O_1479,N_14691,N_14824);
and UO_1480 (O_1480,N_14530,N_14688);
xor UO_1481 (O_1481,N_14952,N_14605);
and UO_1482 (O_1482,N_14317,N_14339);
nor UO_1483 (O_1483,N_14936,N_14443);
and UO_1484 (O_1484,N_14742,N_14827);
nor UO_1485 (O_1485,N_14677,N_14272);
nand UO_1486 (O_1486,N_14308,N_14732);
xnor UO_1487 (O_1487,N_14952,N_14549);
and UO_1488 (O_1488,N_14431,N_14684);
nor UO_1489 (O_1489,N_14341,N_14533);
nand UO_1490 (O_1490,N_14729,N_14291);
xnor UO_1491 (O_1491,N_14259,N_14592);
or UO_1492 (O_1492,N_14358,N_14728);
xor UO_1493 (O_1493,N_14975,N_14411);
or UO_1494 (O_1494,N_14291,N_14318);
xor UO_1495 (O_1495,N_14444,N_14257);
xor UO_1496 (O_1496,N_14714,N_14620);
nand UO_1497 (O_1497,N_14652,N_14718);
or UO_1498 (O_1498,N_14931,N_14691);
and UO_1499 (O_1499,N_14803,N_14783);
and UO_1500 (O_1500,N_14963,N_14700);
nor UO_1501 (O_1501,N_14733,N_14900);
xnor UO_1502 (O_1502,N_14446,N_14812);
or UO_1503 (O_1503,N_14862,N_14617);
and UO_1504 (O_1504,N_14845,N_14666);
and UO_1505 (O_1505,N_14282,N_14519);
xnor UO_1506 (O_1506,N_14876,N_14438);
nand UO_1507 (O_1507,N_14434,N_14686);
xor UO_1508 (O_1508,N_14523,N_14644);
nor UO_1509 (O_1509,N_14496,N_14996);
or UO_1510 (O_1510,N_14472,N_14994);
or UO_1511 (O_1511,N_14713,N_14838);
and UO_1512 (O_1512,N_14489,N_14891);
xnor UO_1513 (O_1513,N_14391,N_14820);
or UO_1514 (O_1514,N_14423,N_14858);
or UO_1515 (O_1515,N_14328,N_14517);
xnor UO_1516 (O_1516,N_14263,N_14922);
and UO_1517 (O_1517,N_14767,N_14810);
and UO_1518 (O_1518,N_14616,N_14593);
xnor UO_1519 (O_1519,N_14382,N_14942);
or UO_1520 (O_1520,N_14533,N_14522);
xnor UO_1521 (O_1521,N_14910,N_14285);
or UO_1522 (O_1522,N_14288,N_14862);
nor UO_1523 (O_1523,N_14806,N_14850);
nand UO_1524 (O_1524,N_14732,N_14668);
or UO_1525 (O_1525,N_14413,N_14953);
nand UO_1526 (O_1526,N_14298,N_14738);
or UO_1527 (O_1527,N_14515,N_14329);
and UO_1528 (O_1528,N_14488,N_14810);
nand UO_1529 (O_1529,N_14534,N_14470);
xor UO_1530 (O_1530,N_14461,N_14774);
nand UO_1531 (O_1531,N_14605,N_14762);
xnor UO_1532 (O_1532,N_14538,N_14408);
nand UO_1533 (O_1533,N_14530,N_14455);
nor UO_1534 (O_1534,N_14686,N_14269);
xor UO_1535 (O_1535,N_14617,N_14427);
and UO_1536 (O_1536,N_14365,N_14536);
and UO_1537 (O_1537,N_14429,N_14697);
xor UO_1538 (O_1538,N_14657,N_14626);
xor UO_1539 (O_1539,N_14789,N_14427);
nor UO_1540 (O_1540,N_14300,N_14776);
or UO_1541 (O_1541,N_14704,N_14609);
xnor UO_1542 (O_1542,N_14832,N_14793);
or UO_1543 (O_1543,N_14340,N_14505);
nor UO_1544 (O_1544,N_14827,N_14879);
and UO_1545 (O_1545,N_14509,N_14402);
nand UO_1546 (O_1546,N_14875,N_14702);
nand UO_1547 (O_1547,N_14553,N_14428);
nor UO_1548 (O_1548,N_14795,N_14525);
nor UO_1549 (O_1549,N_14906,N_14819);
nor UO_1550 (O_1550,N_14887,N_14637);
and UO_1551 (O_1551,N_14826,N_14550);
nor UO_1552 (O_1552,N_14968,N_14935);
nor UO_1553 (O_1553,N_14747,N_14915);
nor UO_1554 (O_1554,N_14400,N_14530);
xnor UO_1555 (O_1555,N_14342,N_14597);
nand UO_1556 (O_1556,N_14421,N_14862);
xor UO_1557 (O_1557,N_14477,N_14343);
nand UO_1558 (O_1558,N_14454,N_14404);
nor UO_1559 (O_1559,N_14759,N_14600);
or UO_1560 (O_1560,N_14636,N_14351);
xor UO_1561 (O_1561,N_14659,N_14716);
nor UO_1562 (O_1562,N_14566,N_14655);
nor UO_1563 (O_1563,N_14854,N_14261);
xnor UO_1564 (O_1564,N_14311,N_14598);
xnor UO_1565 (O_1565,N_14933,N_14354);
xnor UO_1566 (O_1566,N_14777,N_14439);
xor UO_1567 (O_1567,N_14994,N_14926);
nor UO_1568 (O_1568,N_14602,N_14596);
xnor UO_1569 (O_1569,N_14537,N_14871);
xor UO_1570 (O_1570,N_14663,N_14669);
or UO_1571 (O_1571,N_14587,N_14640);
xnor UO_1572 (O_1572,N_14649,N_14409);
xor UO_1573 (O_1573,N_14709,N_14538);
and UO_1574 (O_1574,N_14679,N_14252);
or UO_1575 (O_1575,N_14939,N_14883);
nand UO_1576 (O_1576,N_14372,N_14267);
nand UO_1577 (O_1577,N_14810,N_14713);
or UO_1578 (O_1578,N_14954,N_14906);
and UO_1579 (O_1579,N_14333,N_14318);
or UO_1580 (O_1580,N_14764,N_14531);
or UO_1581 (O_1581,N_14685,N_14697);
and UO_1582 (O_1582,N_14507,N_14574);
and UO_1583 (O_1583,N_14959,N_14979);
and UO_1584 (O_1584,N_14864,N_14822);
or UO_1585 (O_1585,N_14826,N_14832);
nand UO_1586 (O_1586,N_14548,N_14556);
and UO_1587 (O_1587,N_14689,N_14417);
or UO_1588 (O_1588,N_14422,N_14624);
nor UO_1589 (O_1589,N_14388,N_14773);
nor UO_1590 (O_1590,N_14868,N_14687);
and UO_1591 (O_1591,N_14751,N_14826);
nand UO_1592 (O_1592,N_14678,N_14545);
nand UO_1593 (O_1593,N_14333,N_14408);
or UO_1594 (O_1594,N_14295,N_14477);
nand UO_1595 (O_1595,N_14881,N_14929);
nand UO_1596 (O_1596,N_14938,N_14258);
nor UO_1597 (O_1597,N_14571,N_14462);
xnor UO_1598 (O_1598,N_14965,N_14785);
nor UO_1599 (O_1599,N_14579,N_14551);
and UO_1600 (O_1600,N_14600,N_14549);
or UO_1601 (O_1601,N_14605,N_14313);
xor UO_1602 (O_1602,N_14922,N_14880);
and UO_1603 (O_1603,N_14874,N_14631);
xor UO_1604 (O_1604,N_14808,N_14489);
and UO_1605 (O_1605,N_14346,N_14930);
xor UO_1606 (O_1606,N_14607,N_14972);
or UO_1607 (O_1607,N_14972,N_14747);
nand UO_1608 (O_1608,N_14276,N_14540);
nor UO_1609 (O_1609,N_14480,N_14416);
and UO_1610 (O_1610,N_14978,N_14353);
xor UO_1611 (O_1611,N_14519,N_14735);
xor UO_1612 (O_1612,N_14268,N_14655);
and UO_1613 (O_1613,N_14945,N_14432);
xnor UO_1614 (O_1614,N_14656,N_14475);
or UO_1615 (O_1615,N_14412,N_14798);
nand UO_1616 (O_1616,N_14462,N_14615);
nand UO_1617 (O_1617,N_14495,N_14322);
xor UO_1618 (O_1618,N_14925,N_14404);
nor UO_1619 (O_1619,N_14303,N_14312);
nand UO_1620 (O_1620,N_14661,N_14846);
xnor UO_1621 (O_1621,N_14855,N_14299);
nand UO_1622 (O_1622,N_14346,N_14605);
nor UO_1623 (O_1623,N_14908,N_14341);
nand UO_1624 (O_1624,N_14290,N_14684);
xor UO_1625 (O_1625,N_14919,N_14658);
nor UO_1626 (O_1626,N_14319,N_14514);
xor UO_1627 (O_1627,N_14950,N_14836);
or UO_1628 (O_1628,N_14314,N_14390);
or UO_1629 (O_1629,N_14441,N_14826);
or UO_1630 (O_1630,N_14838,N_14761);
nor UO_1631 (O_1631,N_14814,N_14712);
or UO_1632 (O_1632,N_14825,N_14910);
and UO_1633 (O_1633,N_14595,N_14961);
and UO_1634 (O_1634,N_14828,N_14672);
and UO_1635 (O_1635,N_14274,N_14931);
and UO_1636 (O_1636,N_14952,N_14272);
nor UO_1637 (O_1637,N_14572,N_14560);
or UO_1638 (O_1638,N_14675,N_14932);
nor UO_1639 (O_1639,N_14396,N_14816);
xnor UO_1640 (O_1640,N_14839,N_14868);
or UO_1641 (O_1641,N_14494,N_14468);
xnor UO_1642 (O_1642,N_14296,N_14283);
nand UO_1643 (O_1643,N_14334,N_14594);
nand UO_1644 (O_1644,N_14413,N_14692);
nand UO_1645 (O_1645,N_14399,N_14836);
and UO_1646 (O_1646,N_14679,N_14447);
nand UO_1647 (O_1647,N_14379,N_14732);
xnor UO_1648 (O_1648,N_14865,N_14478);
or UO_1649 (O_1649,N_14891,N_14642);
nand UO_1650 (O_1650,N_14846,N_14740);
nand UO_1651 (O_1651,N_14616,N_14294);
or UO_1652 (O_1652,N_14379,N_14762);
or UO_1653 (O_1653,N_14380,N_14277);
nand UO_1654 (O_1654,N_14439,N_14751);
nor UO_1655 (O_1655,N_14497,N_14689);
xnor UO_1656 (O_1656,N_14721,N_14895);
or UO_1657 (O_1657,N_14496,N_14763);
xnor UO_1658 (O_1658,N_14912,N_14552);
or UO_1659 (O_1659,N_14554,N_14476);
nor UO_1660 (O_1660,N_14582,N_14467);
and UO_1661 (O_1661,N_14522,N_14439);
and UO_1662 (O_1662,N_14304,N_14791);
xor UO_1663 (O_1663,N_14573,N_14504);
xor UO_1664 (O_1664,N_14816,N_14593);
or UO_1665 (O_1665,N_14344,N_14882);
nor UO_1666 (O_1666,N_14768,N_14513);
nor UO_1667 (O_1667,N_14482,N_14425);
and UO_1668 (O_1668,N_14445,N_14498);
or UO_1669 (O_1669,N_14272,N_14805);
xnor UO_1670 (O_1670,N_14621,N_14866);
and UO_1671 (O_1671,N_14484,N_14830);
nand UO_1672 (O_1672,N_14439,N_14539);
xor UO_1673 (O_1673,N_14683,N_14483);
nor UO_1674 (O_1674,N_14793,N_14394);
nor UO_1675 (O_1675,N_14477,N_14656);
and UO_1676 (O_1676,N_14438,N_14489);
nor UO_1677 (O_1677,N_14423,N_14743);
and UO_1678 (O_1678,N_14977,N_14329);
or UO_1679 (O_1679,N_14567,N_14796);
nand UO_1680 (O_1680,N_14574,N_14265);
or UO_1681 (O_1681,N_14855,N_14721);
and UO_1682 (O_1682,N_14704,N_14293);
or UO_1683 (O_1683,N_14607,N_14472);
nor UO_1684 (O_1684,N_14753,N_14494);
nand UO_1685 (O_1685,N_14857,N_14784);
nor UO_1686 (O_1686,N_14764,N_14662);
or UO_1687 (O_1687,N_14464,N_14268);
xor UO_1688 (O_1688,N_14537,N_14716);
and UO_1689 (O_1689,N_14942,N_14351);
nor UO_1690 (O_1690,N_14945,N_14401);
xor UO_1691 (O_1691,N_14716,N_14935);
nand UO_1692 (O_1692,N_14441,N_14822);
nor UO_1693 (O_1693,N_14882,N_14586);
xnor UO_1694 (O_1694,N_14515,N_14364);
or UO_1695 (O_1695,N_14573,N_14849);
xnor UO_1696 (O_1696,N_14795,N_14650);
nor UO_1697 (O_1697,N_14672,N_14696);
or UO_1698 (O_1698,N_14411,N_14933);
or UO_1699 (O_1699,N_14766,N_14996);
nand UO_1700 (O_1700,N_14734,N_14756);
and UO_1701 (O_1701,N_14932,N_14337);
nor UO_1702 (O_1702,N_14991,N_14994);
nor UO_1703 (O_1703,N_14802,N_14481);
or UO_1704 (O_1704,N_14371,N_14667);
nor UO_1705 (O_1705,N_14480,N_14462);
and UO_1706 (O_1706,N_14840,N_14756);
nand UO_1707 (O_1707,N_14567,N_14706);
or UO_1708 (O_1708,N_14341,N_14333);
or UO_1709 (O_1709,N_14825,N_14890);
xor UO_1710 (O_1710,N_14546,N_14437);
and UO_1711 (O_1711,N_14345,N_14580);
nor UO_1712 (O_1712,N_14500,N_14400);
and UO_1713 (O_1713,N_14668,N_14738);
and UO_1714 (O_1714,N_14519,N_14386);
nand UO_1715 (O_1715,N_14544,N_14306);
nor UO_1716 (O_1716,N_14567,N_14666);
nand UO_1717 (O_1717,N_14716,N_14817);
nand UO_1718 (O_1718,N_14856,N_14572);
or UO_1719 (O_1719,N_14786,N_14316);
and UO_1720 (O_1720,N_14490,N_14703);
nand UO_1721 (O_1721,N_14706,N_14653);
or UO_1722 (O_1722,N_14646,N_14953);
nand UO_1723 (O_1723,N_14351,N_14656);
and UO_1724 (O_1724,N_14492,N_14966);
nand UO_1725 (O_1725,N_14638,N_14378);
nand UO_1726 (O_1726,N_14505,N_14394);
nor UO_1727 (O_1727,N_14833,N_14932);
xnor UO_1728 (O_1728,N_14605,N_14981);
and UO_1729 (O_1729,N_14617,N_14265);
or UO_1730 (O_1730,N_14255,N_14832);
xnor UO_1731 (O_1731,N_14406,N_14908);
nor UO_1732 (O_1732,N_14344,N_14455);
xor UO_1733 (O_1733,N_14831,N_14579);
nand UO_1734 (O_1734,N_14779,N_14715);
nor UO_1735 (O_1735,N_14584,N_14560);
or UO_1736 (O_1736,N_14345,N_14553);
nand UO_1737 (O_1737,N_14313,N_14880);
nand UO_1738 (O_1738,N_14380,N_14749);
and UO_1739 (O_1739,N_14589,N_14449);
xor UO_1740 (O_1740,N_14951,N_14497);
nor UO_1741 (O_1741,N_14877,N_14883);
and UO_1742 (O_1742,N_14739,N_14254);
and UO_1743 (O_1743,N_14582,N_14280);
xor UO_1744 (O_1744,N_14345,N_14461);
nand UO_1745 (O_1745,N_14280,N_14642);
xor UO_1746 (O_1746,N_14707,N_14580);
nor UO_1747 (O_1747,N_14453,N_14820);
and UO_1748 (O_1748,N_14748,N_14332);
nand UO_1749 (O_1749,N_14346,N_14809);
and UO_1750 (O_1750,N_14828,N_14319);
and UO_1751 (O_1751,N_14719,N_14358);
or UO_1752 (O_1752,N_14250,N_14367);
nor UO_1753 (O_1753,N_14737,N_14817);
xnor UO_1754 (O_1754,N_14690,N_14585);
or UO_1755 (O_1755,N_14508,N_14362);
and UO_1756 (O_1756,N_14344,N_14751);
and UO_1757 (O_1757,N_14531,N_14272);
and UO_1758 (O_1758,N_14385,N_14417);
xnor UO_1759 (O_1759,N_14721,N_14369);
xnor UO_1760 (O_1760,N_14273,N_14603);
and UO_1761 (O_1761,N_14283,N_14818);
nor UO_1762 (O_1762,N_14296,N_14445);
and UO_1763 (O_1763,N_14455,N_14300);
or UO_1764 (O_1764,N_14272,N_14621);
xor UO_1765 (O_1765,N_14674,N_14928);
and UO_1766 (O_1766,N_14758,N_14497);
or UO_1767 (O_1767,N_14780,N_14767);
nor UO_1768 (O_1768,N_14312,N_14642);
and UO_1769 (O_1769,N_14950,N_14424);
nor UO_1770 (O_1770,N_14973,N_14568);
xnor UO_1771 (O_1771,N_14449,N_14538);
nor UO_1772 (O_1772,N_14808,N_14464);
or UO_1773 (O_1773,N_14902,N_14490);
nor UO_1774 (O_1774,N_14765,N_14341);
or UO_1775 (O_1775,N_14321,N_14952);
nand UO_1776 (O_1776,N_14552,N_14656);
or UO_1777 (O_1777,N_14665,N_14828);
xnor UO_1778 (O_1778,N_14996,N_14433);
or UO_1779 (O_1779,N_14381,N_14542);
nor UO_1780 (O_1780,N_14510,N_14494);
nand UO_1781 (O_1781,N_14305,N_14278);
nand UO_1782 (O_1782,N_14468,N_14463);
xor UO_1783 (O_1783,N_14422,N_14615);
or UO_1784 (O_1784,N_14685,N_14735);
and UO_1785 (O_1785,N_14472,N_14752);
nor UO_1786 (O_1786,N_14346,N_14945);
and UO_1787 (O_1787,N_14299,N_14480);
nor UO_1788 (O_1788,N_14432,N_14542);
nand UO_1789 (O_1789,N_14758,N_14855);
xnor UO_1790 (O_1790,N_14849,N_14561);
and UO_1791 (O_1791,N_14536,N_14508);
nor UO_1792 (O_1792,N_14335,N_14484);
xor UO_1793 (O_1793,N_14261,N_14988);
nor UO_1794 (O_1794,N_14374,N_14724);
or UO_1795 (O_1795,N_14951,N_14805);
nand UO_1796 (O_1796,N_14293,N_14687);
nand UO_1797 (O_1797,N_14745,N_14852);
nor UO_1798 (O_1798,N_14628,N_14973);
nor UO_1799 (O_1799,N_14597,N_14334);
nand UO_1800 (O_1800,N_14605,N_14939);
nor UO_1801 (O_1801,N_14426,N_14432);
and UO_1802 (O_1802,N_14606,N_14908);
or UO_1803 (O_1803,N_14303,N_14447);
nand UO_1804 (O_1804,N_14472,N_14938);
nand UO_1805 (O_1805,N_14881,N_14413);
nor UO_1806 (O_1806,N_14891,N_14600);
nor UO_1807 (O_1807,N_14559,N_14679);
nor UO_1808 (O_1808,N_14981,N_14777);
or UO_1809 (O_1809,N_14978,N_14610);
and UO_1810 (O_1810,N_14864,N_14522);
nand UO_1811 (O_1811,N_14307,N_14250);
nand UO_1812 (O_1812,N_14717,N_14983);
and UO_1813 (O_1813,N_14642,N_14816);
or UO_1814 (O_1814,N_14595,N_14574);
nand UO_1815 (O_1815,N_14622,N_14830);
and UO_1816 (O_1816,N_14932,N_14714);
and UO_1817 (O_1817,N_14462,N_14362);
xor UO_1818 (O_1818,N_14607,N_14332);
nor UO_1819 (O_1819,N_14938,N_14546);
or UO_1820 (O_1820,N_14973,N_14683);
or UO_1821 (O_1821,N_14909,N_14601);
nand UO_1822 (O_1822,N_14741,N_14485);
nor UO_1823 (O_1823,N_14625,N_14848);
and UO_1824 (O_1824,N_14603,N_14622);
and UO_1825 (O_1825,N_14523,N_14776);
nor UO_1826 (O_1826,N_14272,N_14565);
xnor UO_1827 (O_1827,N_14903,N_14812);
nor UO_1828 (O_1828,N_14715,N_14275);
and UO_1829 (O_1829,N_14495,N_14596);
xnor UO_1830 (O_1830,N_14882,N_14359);
or UO_1831 (O_1831,N_14960,N_14443);
and UO_1832 (O_1832,N_14891,N_14474);
nand UO_1833 (O_1833,N_14564,N_14662);
and UO_1834 (O_1834,N_14747,N_14309);
nand UO_1835 (O_1835,N_14431,N_14908);
nor UO_1836 (O_1836,N_14702,N_14868);
and UO_1837 (O_1837,N_14922,N_14757);
and UO_1838 (O_1838,N_14284,N_14473);
and UO_1839 (O_1839,N_14719,N_14928);
nor UO_1840 (O_1840,N_14269,N_14577);
nand UO_1841 (O_1841,N_14455,N_14737);
and UO_1842 (O_1842,N_14936,N_14255);
and UO_1843 (O_1843,N_14489,N_14953);
and UO_1844 (O_1844,N_14911,N_14771);
and UO_1845 (O_1845,N_14908,N_14595);
xnor UO_1846 (O_1846,N_14838,N_14903);
nand UO_1847 (O_1847,N_14694,N_14720);
or UO_1848 (O_1848,N_14870,N_14388);
nand UO_1849 (O_1849,N_14464,N_14942);
xnor UO_1850 (O_1850,N_14722,N_14922);
or UO_1851 (O_1851,N_14938,N_14302);
and UO_1852 (O_1852,N_14591,N_14443);
nor UO_1853 (O_1853,N_14574,N_14842);
and UO_1854 (O_1854,N_14879,N_14769);
nor UO_1855 (O_1855,N_14911,N_14587);
and UO_1856 (O_1856,N_14848,N_14745);
and UO_1857 (O_1857,N_14817,N_14413);
and UO_1858 (O_1858,N_14645,N_14665);
xnor UO_1859 (O_1859,N_14755,N_14437);
xor UO_1860 (O_1860,N_14925,N_14298);
and UO_1861 (O_1861,N_14562,N_14333);
or UO_1862 (O_1862,N_14443,N_14876);
or UO_1863 (O_1863,N_14898,N_14408);
or UO_1864 (O_1864,N_14850,N_14637);
nand UO_1865 (O_1865,N_14925,N_14935);
or UO_1866 (O_1866,N_14913,N_14747);
xnor UO_1867 (O_1867,N_14754,N_14337);
nand UO_1868 (O_1868,N_14330,N_14903);
nand UO_1869 (O_1869,N_14865,N_14782);
and UO_1870 (O_1870,N_14466,N_14291);
or UO_1871 (O_1871,N_14911,N_14726);
xor UO_1872 (O_1872,N_14518,N_14263);
nand UO_1873 (O_1873,N_14760,N_14406);
nor UO_1874 (O_1874,N_14918,N_14298);
nand UO_1875 (O_1875,N_14846,N_14376);
or UO_1876 (O_1876,N_14755,N_14872);
or UO_1877 (O_1877,N_14767,N_14782);
or UO_1878 (O_1878,N_14377,N_14597);
and UO_1879 (O_1879,N_14636,N_14909);
or UO_1880 (O_1880,N_14469,N_14691);
nand UO_1881 (O_1881,N_14785,N_14440);
and UO_1882 (O_1882,N_14916,N_14744);
or UO_1883 (O_1883,N_14501,N_14499);
nor UO_1884 (O_1884,N_14616,N_14782);
nand UO_1885 (O_1885,N_14762,N_14430);
nand UO_1886 (O_1886,N_14410,N_14301);
and UO_1887 (O_1887,N_14918,N_14293);
nor UO_1888 (O_1888,N_14325,N_14948);
xor UO_1889 (O_1889,N_14694,N_14553);
xor UO_1890 (O_1890,N_14724,N_14557);
nor UO_1891 (O_1891,N_14673,N_14300);
xor UO_1892 (O_1892,N_14970,N_14469);
or UO_1893 (O_1893,N_14885,N_14858);
and UO_1894 (O_1894,N_14534,N_14911);
and UO_1895 (O_1895,N_14917,N_14676);
xor UO_1896 (O_1896,N_14282,N_14862);
nor UO_1897 (O_1897,N_14828,N_14960);
and UO_1898 (O_1898,N_14408,N_14534);
nand UO_1899 (O_1899,N_14458,N_14600);
nand UO_1900 (O_1900,N_14727,N_14758);
nand UO_1901 (O_1901,N_14826,N_14739);
nand UO_1902 (O_1902,N_14258,N_14428);
xnor UO_1903 (O_1903,N_14544,N_14854);
xnor UO_1904 (O_1904,N_14516,N_14535);
nor UO_1905 (O_1905,N_14840,N_14578);
or UO_1906 (O_1906,N_14483,N_14906);
nor UO_1907 (O_1907,N_14629,N_14680);
xnor UO_1908 (O_1908,N_14418,N_14257);
or UO_1909 (O_1909,N_14524,N_14698);
nand UO_1910 (O_1910,N_14308,N_14632);
and UO_1911 (O_1911,N_14906,N_14784);
xnor UO_1912 (O_1912,N_14498,N_14893);
xor UO_1913 (O_1913,N_14537,N_14723);
nand UO_1914 (O_1914,N_14984,N_14277);
nor UO_1915 (O_1915,N_14720,N_14265);
xnor UO_1916 (O_1916,N_14256,N_14795);
and UO_1917 (O_1917,N_14301,N_14758);
xnor UO_1918 (O_1918,N_14428,N_14377);
nand UO_1919 (O_1919,N_14421,N_14385);
nand UO_1920 (O_1920,N_14996,N_14587);
nor UO_1921 (O_1921,N_14360,N_14628);
nor UO_1922 (O_1922,N_14761,N_14841);
nor UO_1923 (O_1923,N_14643,N_14619);
nand UO_1924 (O_1924,N_14289,N_14617);
and UO_1925 (O_1925,N_14705,N_14363);
nand UO_1926 (O_1926,N_14342,N_14872);
nor UO_1927 (O_1927,N_14281,N_14725);
or UO_1928 (O_1928,N_14679,N_14808);
nand UO_1929 (O_1929,N_14634,N_14762);
and UO_1930 (O_1930,N_14354,N_14270);
nor UO_1931 (O_1931,N_14338,N_14368);
or UO_1932 (O_1932,N_14457,N_14370);
or UO_1933 (O_1933,N_14980,N_14354);
xor UO_1934 (O_1934,N_14417,N_14290);
nand UO_1935 (O_1935,N_14522,N_14376);
xnor UO_1936 (O_1936,N_14952,N_14946);
nor UO_1937 (O_1937,N_14522,N_14290);
and UO_1938 (O_1938,N_14934,N_14525);
xor UO_1939 (O_1939,N_14379,N_14604);
xor UO_1940 (O_1940,N_14740,N_14542);
and UO_1941 (O_1941,N_14827,N_14278);
xnor UO_1942 (O_1942,N_14686,N_14428);
nor UO_1943 (O_1943,N_14676,N_14388);
or UO_1944 (O_1944,N_14460,N_14968);
nor UO_1945 (O_1945,N_14815,N_14436);
xnor UO_1946 (O_1946,N_14254,N_14713);
nand UO_1947 (O_1947,N_14831,N_14419);
nand UO_1948 (O_1948,N_14603,N_14283);
nand UO_1949 (O_1949,N_14629,N_14578);
nor UO_1950 (O_1950,N_14811,N_14320);
xor UO_1951 (O_1951,N_14873,N_14953);
nand UO_1952 (O_1952,N_14746,N_14378);
xor UO_1953 (O_1953,N_14598,N_14415);
nand UO_1954 (O_1954,N_14712,N_14793);
nand UO_1955 (O_1955,N_14503,N_14494);
nor UO_1956 (O_1956,N_14849,N_14858);
xor UO_1957 (O_1957,N_14344,N_14441);
xor UO_1958 (O_1958,N_14975,N_14597);
and UO_1959 (O_1959,N_14625,N_14719);
and UO_1960 (O_1960,N_14539,N_14715);
nor UO_1961 (O_1961,N_14920,N_14484);
nor UO_1962 (O_1962,N_14585,N_14716);
nand UO_1963 (O_1963,N_14845,N_14455);
nand UO_1964 (O_1964,N_14610,N_14392);
or UO_1965 (O_1965,N_14658,N_14727);
xnor UO_1966 (O_1966,N_14851,N_14675);
nor UO_1967 (O_1967,N_14749,N_14255);
nand UO_1968 (O_1968,N_14769,N_14954);
nor UO_1969 (O_1969,N_14537,N_14589);
nor UO_1970 (O_1970,N_14739,N_14866);
xnor UO_1971 (O_1971,N_14285,N_14324);
nand UO_1972 (O_1972,N_14664,N_14373);
and UO_1973 (O_1973,N_14311,N_14738);
nor UO_1974 (O_1974,N_14762,N_14777);
or UO_1975 (O_1975,N_14275,N_14572);
or UO_1976 (O_1976,N_14518,N_14671);
xor UO_1977 (O_1977,N_14953,N_14585);
nor UO_1978 (O_1978,N_14904,N_14305);
nor UO_1979 (O_1979,N_14410,N_14638);
and UO_1980 (O_1980,N_14268,N_14865);
and UO_1981 (O_1981,N_14793,N_14429);
nor UO_1982 (O_1982,N_14538,N_14689);
xnor UO_1983 (O_1983,N_14425,N_14964);
nand UO_1984 (O_1984,N_14261,N_14912);
and UO_1985 (O_1985,N_14745,N_14650);
or UO_1986 (O_1986,N_14474,N_14400);
and UO_1987 (O_1987,N_14265,N_14750);
nor UO_1988 (O_1988,N_14927,N_14426);
nor UO_1989 (O_1989,N_14533,N_14737);
nor UO_1990 (O_1990,N_14880,N_14545);
and UO_1991 (O_1991,N_14685,N_14894);
xor UO_1992 (O_1992,N_14390,N_14868);
and UO_1993 (O_1993,N_14698,N_14332);
nor UO_1994 (O_1994,N_14367,N_14356);
nor UO_1995 (O_1995,N_14368,N_14836);
and UO_1996 (O_1996,N_14858,N_14871);
nand UO_1997 (O_1997,N_14465,N_14568);
or UO_1998 (O_1998,N_14391,N_14734);
or UO_1999 (O_1999,N_14429,N_14916);
endmodule