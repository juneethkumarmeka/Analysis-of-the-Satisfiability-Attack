module basic_500_3000_500_15_levels_5xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
xnor U0 (N_0,In_356,In_298);
nor U1 (N_1,In_184,In_52);
nand U2 (N_2,In_339,In_312);
and U3 (N_3,In_334,In_486);
and U4 (N_4,In_131,In_388);
or U5 (N_5,In_324,In_418);
or U6 (N_6,In_8,In_327);
nor U7 (N_7,In_168,In_101);
or U8 (N_8,In_423,In_147);
xor U9 (N_9,In_203,In_217);
xor U10 (N_10,In_17,In_54);
or U11 (N_11,In_460,In_129);
or U12 (N_12,In_474,In_408);
nand U13 (N_13,In_58,In_482);
or U14 (N_14,In_372,In_228);
nor U15 (N_15,In_336,In_459);
or U16 (N_16,In_133,In_94);
nor U17 (N_17,In_452,In_28);
nand U18 (N_18,In_303,In_247);
nor U19 (N_19,In_427,In_497);
nor U20 (N_20,In_79,In_330);
and U21 (N_21,In_83,In_103);
and U22 (N_22,In_78,In_57);
xor U23 (N_23,In_439,In_390);
nand U24 (N_24,In_405,In_358);
xor U25 (N_25,In_496,In_499);
or U26 (N_26,In_267,In_242);
nand U27 (N_27,In_127,In_430);
nor U28 (N_28,In_498,In_323);
xor U29 (N_29,In_74,In_111);
nor U30 (N_30,In_266,In_332);
nor U31 (N_31,In_462,In_260);
or U32 (N_32,In_273,In_268);
nand U33 (N_33,In_185,In_441);
nand U34 (N_34,In_89,In_92);
nor U35 (N_35,In_422,In_21);
or U36 (N_36,In_443,In_55);
or U37 (N_37,In_475,In_47);
nand U38 (N_38,In_48,In_15);
and U39 (N_39,In_425,In_46);
or U40 (N_40,In_3,In_331);
or U41 (N_41,In_467,In_299);
nand U42 (N_42,In_181,In_428);
or U43 (N_43,In_387,In_230);
nand U44 (N_44,In_108,In_357);
nor U45 (N_45,In_189,In_162);
nor U46 (N_46,In_302,In_346);
nand U47 (N_47,In_60,In_16);
nor U48 (N_48,In_176,In_179);
or U49 (N_49,In_286,In_288);
or U50 (N_50,In_300,In_106);
nor U51 (N_51,In_420,In_442);
and U52 (N_52,In_464,In_237);
nor U53 (N_53,In_436,In_151);
nand U54 (N_54,In_326,In_257);
or U55 (N_55,In_367,In_297);
or U56 (N_56,In_274,In_248);
or U57 (N_57,In_278,In_112);
xor U58 (N_58,In_39,In_1);
or U59 (N_59,In_161,In_457);
and U60 (N_60,In_276,In_333);
or U61 (N_61,In_170,In_22);
nand U62 (N_62,In_322,In_148);
nand U63 (N_63,In_338,In_56);
nor U64 (N_64,In_279,In_448);
nand U65 (N_65,In_403,In_280);
or U66 (N_66,In_262,In_310);
and U67 (N_67,In_251,In_195);
nand U68 (N_68,In_292,In_153);
nor U69 (N_69,In_289,In_488);
nor U70 (N_70,In_171,In_377);
and U71 (N_71,In_281,In_156);
nor U72 (N_72,In_212,In_354);
nand U73 (N_73,In_159,In_183);
xor U74 (N_74,In_205,In_490);
nor U75 (N_75,In_117,In_264);
or U76 (N_76,In_100,In_296);
or U77 (N_77,In_27,In_398);
nand U78 (N_78,In_187,In_23);
nand U79 (N_79,In_72,In_191);
nor U80 (N_80,In_199,In_107);
nor U81 (N_81,In_360,In_366);
nor U82 (N_82,In_59,In_68);
or U83 (N_83,In_419,In_210);
nand U84 (N_84,In_362,In_487);
nor U85 (N_85,In_82,In_105);
nand U86 (N_86,In_400,In_456);
and U87 (N_87,In_320,In_53);
and U88 (N_88,In_136,In_383);
or U89 (N_89,In_18,In_227);
or U90 (N_90,In_144,In_402);
or U91 (N_91,In_468,In_244);
nand U92 (N_92,In_328,In_365);
nand U93 (N_93,In_149,In_114);
xor U94 (N_94,In_359,In_392);
and U95 (N_95,In_97,In_122);
or U96 (N_96,In_69,In_174);
and U97 (N_97,In_65,In_253);
or U98 (N_98,In_50,In_382);
and U99 (N_99,In_344,In_313);
xnor U100 (N_100,In_222,In_413);
nand U101 (N_101,In_77,In_325);
nor U102 (N_102,In_173,In_36);
xnor U103 (N_103,In_235,In_369);
and U104 (N_104,In_182,In_216);
or U105 (N_105,In_88,In_43);
nor U106 (N_106,In_7,In_469);
nand U107 (N_107,In_113,In_252);
nand U108 (N_108,In_305,In_416);
nand U109 (N_109,In_33,In_283);
and U110 (N_110,In_435,In_411);
nor U111 (N_111,In_86,In_353);
nand U112 (N_112,In_142,In_209);
or U113 (N_113,In_479,In_407);
nor U114 (N_114,In_141,In_316);
nand U115 (N_115,In_215,In_306);
or U116 (N_116,In_478,In_396);
nor U117 (N_117,In_98,In_14);
nor U118 (N_118,In_219,In_90);
nand U119 (N_119,In_317,In_66);
or U120 (N_120,In_269,In_348);
nor U121 (N_121,In_431,In_424);
xnor U122 (N_122,In_393,In_34);
and U123 (N_123,In_473,In_485);
and U124 (N_124,In_211,In_406);
nor U125 (N_125,In_221,In_437);
xnor U126 (N_126,In_109,In_342);
nor U127 (N_127,In_355,In_453);
nor U128 (N_128,In_275,In_410);
nand U129 (N_129,In_2,In_287);
and U130 (N_130,In_73,In_5);
or U131 (N_131,In_493,In_120);
nor U132 (N_132,In_255,In_294);
and U133 (N_133,In_449,In_96);
nor U134 (N_134,In_125,In_186);
and U135 (N_135,In_471,In_373);
or U136 (N_136,In_91,In_350);
and U137 (N_137,In_138,In_225);
nand U138 (N_138,In_261,In_236);
or U139 (N_139,In_207,In_495);
and U140 (N_140,In_232,In_139);
and U141 (N_141,In_38,In_87);
nor U142 (N_142,In_384,In_140);
nor U143 (N_143,In_24,In_51);
nor U144 (N_144,In_128,In_29);
and U145 (N_145,In_318,In_399);
nand U146 (N_146,In_351,In_391);
nor U147 (N_147,In_12,In_284);
and U148 (N_148,In_220,In_61);
nand U149 (N_149,In_9,In_238);
and U150 (N_150,In_172,In_433);
nand U151 (N_151,In_308,In_285);
nand U152 (N_152,In_0,In_206);
or U153 (N_153,In_63,In_379);
xor U154 (N_154,In_67,In_152);
and U155 (N_155,In_218,In_470);
and U156 (N_156,In_45,In_415);
nand U157 (N_157,In_190,In_163);
or U158 (N_158,In_81,In_31);
xnor U159 (N_159,In_314,In_463);
nor U160 (N_160,In_116,In_135);
and U161 (N_161,In_447,In_193);
or U162 (N_162,In_432,In_145);
and U163 (N_163,In_95,In_231);
and U164 (N_164,In_201,In_71);
and U165 (N_165,In_226,In_434);
or U166 (N_166,In_394,In_385);
and U167 (N_167,In_480,In_123);
nor U168 (N_168,In_102,In_481);
or U169 (N_169,In_343,In_341);
and U170 (N_170,In_64,In_154);
xor U171 (N_171,In_370,In_223);
and U172 (N_172,In_401,In_241);
nand U173 (N_173,In_389,In_349);
and U174 (N_174,In_380,In_375);
or U175 (N_175,In_282,In_438);
nand U176 (N_176,In_62,In_99);
and U177 (N_177,In_492,In_472);
nor U178 (N_178,In_397,In_352);
nor U179 (N_179,In_254,In_118);
and U180 (N_180,In_315,In_291);
and U181 (N_181,In_304,In_178);
or U182 (N_182,In_426,In_249);
or U183 (N_183,In_451,In_155);
nor U184 (N_184,In_44,In_455);
nand U185 (N_185,In_126,In_445);
and U186 (N_186,In_263,In_440);
and U187 (N_187,In_35,In_6);
and U188 (N_188,In_409,In_85);
xnor U189 (N_189,In_265,In_192);
nor U190 (N_190,In_250,In_293);
nor U191 (N_191,In_477,In_75);
or U192 (N_192,In_272,In_446);
and U193 (N_193,In_200,In_347);
or U194 (N_194,In_42,In_76);
nor U195 (N_195,In_361,In_10);
nand U196 (N_196,In_41,In_11);
nor U197 (N_197,In_158,In_466);
nor U198 (N_198,In_414,In_40);
nand U199 (N_199,In_202,In_124);
and U200 (N_200,N_159,N_88);
or U201 (N_201,N_4,N_53);
nand U202 (N_202,N_139,N_151);
nor U203 (N_203,N_98,N_155);
or U204 (N_204,N_142,In_93);
nand U205 (N_205,N_149,N_71);
nor U206 (N_206,N_190,In_25);
xnor U207 (N_207,In_157,In_119);
nand U208 (N_208,In_484,N_126);
nor U209 (N_209,N_94,N_189);
or U210 (N_210,N_154,N_19);
or U211 (N_211,In_290,In_70);
nand U212 (N_212,In_461,In_319);
or U213 (N_213,N_10,N_109);
and U214 (N_214,N_186,In_115);
nor U215 (N_215,In_167,N_177);
nor U216 (N_216,N_34,In_386);
nand U217 (N_217,N_167,N_22);
and U218 (N_218,N_163,N_116);
nand U219 (N_219,N_67,N_134);
and U220 (N_220,N_74,N_188);
xnor U221 (N_221,In_374,N_73);
nor U222 (N_222,In_329,N_30);
nand U223 (N_223,In_246,In_340);
and U224 (N_224,In_37,N_122);
or U225 (N_225,N_172,N_64);
and U226 (N_226,In_134,N_45);
and U227 (N_227,N_183,N_147);
nand U228 (N_228,In_160,N_160);
and U229 (N_229,N_86,N_3);
nand U230 (N_230,N_108,In_234);
nand U231 (N_231,N_33,N_6);
or U232 (N_232,N_2,N_136);
nand U233 (N_233,N_131,N_96);
or U234 (N_234,N_46,In_270);
xor U235 (N_235,In_130,N_125);
and U236 (N_236,In_309,N_79);
or U237 (N_237,N_91,N_114);
and U238 (N_238,N_23,N_120);
xor U239 (N_239,In_110,N_7);
nor U240 (N_240,N_55,In_32);
and U241 (N_241,N_168,N_1);
or U242 (N_242,N_41,N_145);
or U243 (N_243,In_494,In_104);
nand U244 (N_244,N_141,In_213);
xor U245 (N_245,N_138,In_233);
or U246 (N_246,In_80,N_127);
or U247 (N_247,N_24,N_47);
nor U248 (N_248,N_105,In_150);
or U249 (N_249,In_295,In_454);
and U250 (N_250,N_31,N_146);
or U251 (N_251,N_161,N_42);
nor U252 (N_252,In_49,N_51);
or U253 (N_253,N_121,In_224);
xor U254 (N_254,N_171,N_28);
nor U255 (N_255,N_78,N_11);
nor U256 (N_256,N_198,In_164);
nor U257 (N_257,N_16,N_100);
and U258 (N_258,In_121,N_104);
and U259 (N_259,N_187,In_30);
nor U260 (N_260,N_194,In_245);
or U261 (N_261,In_364,N_92);
and U262 (N_262,N_152,N_140);
nand U263 (N_263,N_153,In_277);
and U264 (N_264,N_148,N_95);
nor U265 (N_265,N_93,N_62);
nand U266 (N_266,In_476,N_65);
nand U267 (N_267,N_5,N_80);
and U268 (N_268,N_169,N_43);
or U269 (N_269,In_271,In_483);
nor U270 (N_270,N_44,N_110);
nor U271 (N_271,N_90,In_395);
and U272 (N_272,N_132,N_192);
and U273 (N_273,In_465,In_458);
and U274 (N_274,N_124,N_14);
nor U275 (N_275,N_99,In_229);
or U276 (N_276,N_36,N_29);
and U277 (N_277,In_132,N_27);
nor U278 (N_278,N_25,N_191);
nor U279 (N_279,N_48,N_184);
or U280 (N_280,N_37,N_97);
and U281 (N_281,In_450,N_103);
nor U282 (N_282,N_50,In_301);
nand U283 (N_283,In_165,N_178);
or U284 (N_284,In_180,N_83);
nor U285 (N_285,N_150,In_13);
nand U286 (N_286,In_20,N_54);
or U287 (N_287,N_199,N_69);
or U288 (N_288,N_196,N_182);
and U289 (N_289,N_72,In_321);
xnor U290 (N_290,In_258,N_123);
or U291 (N_291,In_204,N_61);
nand U292 (N_292,N_0,N_8);
nand U293 (N_293,N_176,N_157);
xor U294 (N_294,In_198,In_166);
or U295 (N_295,N_52,N_17);
and U296 (N_296,N_174,N_133);
and U297 (N_297,N_195,N_49);
nor U298 (N_298,In_137,N_68);
nor U299 (N_299,N_89,N_39);
nor U300 (N_300,N_156,In_84);
nand U301 (N_301,In_381,In_26);
or U302 (N_302,N_143,N_185);
nor U303 (N_303,In_337,N_179);
or U304 (N_304,N_107,In_240);
nand U305 (N_305,N_76,In_491);
nand U306 (N_306,In_239,N_102);
or U307 (N_307,N_21,N_12);
xnor U308 (N_308,N_18,N_181);
nor U309 (N_309,In_311,In_412);
nor U310 (N_310,In_194,N_193);
and U311 (N_311,In_421,N_85);
and U312 (N_312,In_363,In_376);
nor U313 (N_313,In_378,N_197);
or U314 (N_314,N_111,N_135);
nand U315 (N_315,N_40,In_175);
and U316 (N_316,In_256,N_9);
nand U317 (N_317,N_26,In_196);
and U318 (N_318,N_101,In_214);
nor U319 (N_319,In_146,In_335);
nor U320 (N_320,In_208,N_115);
or U321 (N_321,N_15,In_345);
and U322 (N_322,In_188,In_243);
and U323 (N_323,In_404,N_84);
nand U324 (N_324,In_417,N_180);
or U325 (N_325,N_60,In_371);
or U326 (N_326,N_56,N_112);
nor U327 (N_327,N_81,N_166);
nand U328 (N_328,N_106,N_66);
nand U329 (N_329,N_164,N_35);
nand U330 (N_330,In_143,N_165);
nand U331 (N_331,N_128,N_58);
or U332 (N_332,N_170,N_119);
nor U333 (N_333,N_175,In_259);
or U334 (N_334,N_70,N_32);
and U335 (N_335,In_177,In_429);
and U336 (N_336,In_19,N_57);
nand U337 (N_337,N_87,N_59);
nand U338 (N_338,N_82,N_113);
or U339 (N_339,N_158,N_144);
and U340 (N_340,N_162,N_77);
and U341 (N_341,N_75,In_489);
or U342 (N_342,N_117,N_129);
or U343 (N_343,N_137,N_38);
nor U344 (N_344,N_130,N_63);
nand U345 (N_345,N_118,In_169);
and U346 (N_346,N_13,In_4);
nor U347 (N_347,N_173,In_307);
nor U348 (N_348,In_444,In_197);
or U349 (N_349,In_368,N_20);
nand U350 (N_350,In_246,In_258);
nand U351 (N_351,In_246,N_113);
and U352 (N_352,N_25,N_14);
or U353 (N_353,N_60,In_368);
or U354 (N_354,N_19,N_196);
nand U355 (N_355,N_102,N_161);
nand U356 (N_356,In_197,N_48);
nor U357 (N_357,In_240,N_96);
nor U358 (N_358,In_197,N_195);
nand U359 (N_359,N_102,N_61);
nand U360 (N_360,In_204,N_113);
and U361 (N_361,In_194,In_412);
and U362 (N_362,N_74,In_157);
or U363 (N_363,In_417,N_67);
or U364 (N_364,In_484,N_46);
and U365 (N_365,N_31,N_7);
nand U366 (N_366,N_139,N_161);
nor U367 (N_367,N_185,N_55);
or U368 (N_368,In_240,N_180);
nand U369 (N_369,N_162,N_181);
and U370 (N_370,N_103,In_198);
nor U371 (N_371,N_148,N_106);
nand U372 (N_372,In_177,In_49);
xor U373 (N_373,N_27,In_277);
or U374 (N_374,In_143,N_153);
nand U375 (N_375,N_180,N_152);
nor U376 (N_376,N_149,N_171);
and U377 (N_377,In_417,N_118);
nor U378 (N_378,N_10,N_7);
nand U379 (N_379,N_29,In_26);
and U380 (N_380,N_80,N_162);
or U381 (N_381,N_17,In_381);
nor U382 (N_382,In_321,In_180);
or U383 (N_383,N_17,In_164);
xor U384 (N_384,In_483,N_99);
or U385 (N_385,N_75,N_192);
or U386 (N_386,In_364,N_21);
nand U387 (N_387,N_25,N_34);
xnor U388 (N_388,N_105,N_19);
and U389 (N_389,N_78,N_63);
or U390 (N_390,In_489,N_131);
nor U391 (N_391,N_23,N_48);
nor U392 (N_392,In_245,N_184);
nand U393 (N_393,In_150,N_86);
nand U394 (N_394,In_19,N_77);
and U395 (N_395,N_95,In_164);
nand U396 (N_396,In_150,In_319);
nand U397 (N_397,In_245,N_50);
and U398 (N_398,In_180,In_188);
nand U399 (N_399,N_24,N_41);
xor U400 (N_400,N_352,N_249);
and U401 (N_401,N_212,N_285);
or U402 (N_402,N_290,N_349);
or U403 (N_403,N_390,N_354);
or U404 (N_404,N_235,N_399);
xnor U405 (N_405,N_307,N_293);
or U406 (N_406,N_364,N_221);
nand U407 (N_407,N_381,N_328);
and U408 (N_408,N_276,N_264);
or U409 (N_409,N_296,N_347);
nor U410 (N_410,N_256,N_389);
or U411 (N_411,N_394,N_391);
nor U412 (N_412,N_286,N_335);
and U413 (N_413,N_227,N_216);
nand U414 (N_414,N_214,N_243);
xnor U415 (N_415,N_304,N_244);
and U416 (N_416,N_311,N_254);
nand U417 (N_417,N_386,N_383);
nand U418 (N_418,N_396,N_261);
nor U419 (N_419,N_213,N_255);
or U420 (N_420,N_269,N_232);
nand U421 (N_421,N_226,N_313);
or U422 (N_422,N_340,N_306);
xnor U423 (N_423,N_294,N_375);
or U424 (N_424,N_208,N_250);
nor U425 (N_425,N_362,N_372);
xnor U426 (N_426,N_329,N_283);
or U427 (N_427,N_267,N_268);
nor U428 (N_428,N_280,N_397);
nand U429 (N_429,N_339,N_305);
nand U430 (N_430,N_272,N_238);
nor U431 (N_431,N_299,N_271);
nor U432 (N_432,N_218,N_277);
nor U433 (N_433,N_225,N_263);
nand U434 (N_434,N_374,N_346);
and U435 (N_435,N_316,N_382);
nor U436 (N_436,N_317,N_330);
or U437 (N_437,N_247,N_262);
xnor U438 (N_438,N_358,N_302);
nand U439 (N_439,N_231,N_334);
or U440 (N_440,N_395,N_361);
or U441 (N_441,N_266,N_228);
xor U442 (N_442,N_363,N_204);
nor U443 (N_443,N_245,N_303);
nor U444 (N_444,N_275,N_259);
or U445 (N_445,N_200,N_357);
xnor U446 (N_446,N_336,N_265);
nand U447 (N_447,N_327,N_350);
or U448 (N_448,N_209,N_332);
nor U449 (N_449,N_278,N_234);
nor U450 (N_450,N_322,N_260);
nand U451 (N_451,N_388,N_312);
nor U452 (N_452,N_337,N_369);
or U453 (N_453,N_201,N_343);
xnor U454 (N_454,N_242,N_351);
or U455 (N_455,N_370,N_325);
nor U456 (N_456,N_233,N_241);
or U457 (N_457,N_368,N_373);
nor U458 (N_458,N_309,N_331);
nand U459 (N_459,N_392,N_291);
or U460 (N_460,N_282,N_314);
nand U461 (N_461,N_378,N_203);
or U462 (N_462,N_205,N_252);
and U463 (N_463,N_365,N_310);
nor U464 (N_464,N_297,N_207);
nor U465 (N_465,N_359,N_230);
nand U466 (N_466,N_236,N_279);
xor U467 (N_467,N_300,N_251);
and U468 (N_468,N_217,N_211);
and U469 (N_469,N_287,N_206);
nand U470 (N_470,N_248,N_356);
xor U471 (N_471,N_239,N_215);
nand U472 (N_472,N_284,N_274);
or U473 (N_473,N_376,N_289);
nand U474 (N_474,N_301,N_341);
nand U475 (N_475,N_387,N_342);
xnor U476 (N_476,N_367,N_393);
or U477 (N_477,N_281,N_348);
nand U478 (N_478,N_324,N_344);
nand U479 (N_479,N_253,N_377);
nand U480 (N_480,N_292,N_321);
and U481 (N_481,N_288,N_224);
and U482 (N_482,N_338,N_308);
nand U483 (N_483,N_219,N_246);
and U484 (N_484,N_371,N_223);
nand U485 (N_485,N_240,N_366);
or U486 (N_486,N_353,N_323);
nand U487 (N_487,N_318,N_345);
nand U488 (N_488,N_385,N_270);
and U489 (N_489,N_319,N_222);
nor U490 (N_490,N_295,N_220);
and U491 (N_491,N_320,N_379);
nand U492 (N_492,N_229,N_355);
nand U493 (N_493,N_298,N_360);
or U494 (N_494,N_326,N_398);
nand U495 (N_495,N_333,N_380);
nor U496 (N_496,N_384,N_237);
and U497 (N_497,N_202,N_315);
or U498 (N_498,N_273,N_257);
and U499 (N_499,N_258,N_210);
nand U500 (N_500,N_369,N_298);
nor U501 (N_501,N_305,N_396);
and U502 (N_502,N_339,N_260);
nor U503 (N_503,N_243,N_295);
nand U504 (N_504,N_228,N_389);
or U505 (N_505,N_314,N_392);
nand U506 (N_506,N_263,N_248);
nand U507 (N_507,N_319,N_256);
or U508 (N_508,N_209,N_236);
nand U509 (N_509,N_324,N_201);
nand U510 (N_510,N_240,N_361);
nand U511 (N_511,N_365,N_223);
xor U512 (N_512,N_297,N_315);
nor U513 (N_513,N_307,N_347);
xnor U514 (N_514,N_245,N_383);
and U515 (N_515,N_269,N_315);
or U516 (N_516,N_382,N_200);
or U517 (N_517,N_342,N_284);
and U518 (N_518,N_386,N_235);
nor U519 (N_519,N_272,N_245);
nor U520 (N_520,N_282,N_380);
nor U521 (N_521,N_261,N_302);
xnor U522 (N_522,N_201,N_392);
nor U523 (N_523,N_210,N_387);
or U524 (N_524,N_278,N_306);
and U525 (N_525,N_273,N_224);
or U526 (N_526,N_229,N_341);
and U527 (N_527,N_327,N_303);
xnor U528 (N_528,N_363,N_333);
xnor U529 (N_529,N_377,N_316);
nor U530 (N_530,N_347,N_355);
nor U531 (N_531,N_283,N_342);
xor U532 (N_532,N_309,N_378);
nor U533 (N_533,N_265,N_389);
or U534 (N_534,N_272,N_332);
and U535 (N_535,N_216,N_342);
xnor U536 (N_536,N_261,N_264);
nor U537 (N_537,N_200,N_298);
or U538 (N_538,N_274,N_244);
or U539 (N_539,N_296,N_361);
xnor U540 (N_540,N_385,N_248);
nor U541 (N_541,N_352,N_339);
or U542 (N_542,N_397,N_369);
or U543 (N_543,N_340,N_298);
and U544 (N_544,N_279,N_384);
and U545 (N_545,N_210,N_367);
and U546 (N_546,N_249,N_221);
and U547 (N_547,N_299,N_361);
or U548 (N_548,N_395,N_378);
or U549 (N_549,N_377,N_349);
nor U550 (N_550,N_295,N_237);
xnor U551 (N_551,N_342,N_393);
or U552 (N_552,N_248,N_204);
nand U553 (N_553,N_274,N_326);
nand U554 (N_554,N_329,N_337);
or U555 (N_555,N_331,N_379);
and U556 (N_556,N_240,N_388);
nor U557 (N_557,N_388,N_209);
or U558 (N_558,N_370,N_280);
and U559 (N_559,N_383,N_212);
or U560 (N_560,N_269,N_300);
nand U561 (N_561,N_204,N_380);
nand U562 (N_562,N_316,N_229);
nand U563 (N_563,N_299,N_259);
and U564 (N_564,N_300,N_239);
or U565 (N_565,N_317,N_236);
and U566 (N_566,N_294,N_384);
xnor U567 (N_567,N_252,N_317);
nand U568 (N_568,N_290,N_315);
xnor U569 (N_569,N_359,N_207);
nand U570 (N_570,N_241,N_216);
nor U571 (N_571,N_243,N_339);
or U572 (N_572,N_395,N_344);
nand U573 (N_573,N_321,N_388);
or U574 (N_574,N_357,N_348);
nand U575 (N_575,N_329,N_231);
and U576 (N_576,N_336,N_270);
nor U577 (N_577,N_297,N_351);
and U578 (N_578,N_333,N_283);
xor U579 (N_579,N_270,N_210);
or U580 (N_580,N_335,N_324);
or U581 (N_581,N_302,N_253);
and U582 (N_582,N_315,N_204);
and U583 (N_583,N_230,N_310);
nand U584 (N_584,N_244,N_260);
nor U585 (N_585,N_211,N_276);
nor U586 (N_586,N_305,N_306);
nand U587 (N_587,N_390,N_229);
and U588 (N_588,N_205,N_227);
xnor U589 (N_589,N_225,N_353);
nor U590 (N_590,N_334,N_267);
nand U591 (N_591,N_324,N_309);
nor U592 (N_592,N_331,N_211);
nand U593 (N_593,N_215,N_344);
and U594 (N_594,N_344,N_245);
nand U595 (N_595,N_201,N_243);
and U596 (N_596,N_375,N_234);
nor U597 (N_597,N_284,N_206);
or U598 (N_598,N_376,N_367);
xnor U599 (N_599,N_392,N_296);
and U600 (N_600,N_548,N_403);
xnor U601 (N_601,N_420,N_534);
nor U602 (N_602,N_536,N_439);
nand U603 (N_603,N_452,N_437);
or U604 (N_604,N_570,N_527);
and U605 (N_605,N_412,N_554);
or U606 (N_606,N_423,N_443);
and U607 (N_607,N_572,N_427);
nor U608 (N_608,N_475,N_540);
or U609 (N_609,N_477,N_598);
nand U610 (N_610,N_448,N_532);
and U611 (N_611,N_469,N_556);
nor U612 (N_612,N_509,N_595);
nand U613 (N_613,N_511,N_487);
and U614 (N_614,N_472,N_596);
and U615 (N_615,N_408,N_464);
or U616 (N_616,N_560,N_411);
nor U617 (N_617,N_497,N_587);
and U618 (N_618,N_459,N_529);
nor U619 (N_619,N_454,N_599);
and U620 (N_620,N_440,N_582);
and U621 (N_621,N_467,N_405);
and U622 (N_622,N_549,N_425);
and U623 (N_623,N_579,N_471);
or U624 (N_624,N_493,N_580);
and U625 (N_625,N_531,N_483);
or U626 (N_626,N_577,N_555);
nand U627 (N_627,N_465,N_495);
xor U628 (N_628,N_508,N_557);
and U629 (N_629,N_571,N_462);
and U630 (N_630,N_450,N_490);
nor U631 (N_631,N_586,N_568);
xor U632 (N_632,N_401,N_442);
and U633 (N_633,N_461,N_575);
or U634 (N_634,N_515,N_498);
and U635 (N_635,N_521,N_516);
nor U636 (N_636,N_589,N_518);
nor U637 (N_637,N_410,N_447);
or U638 (N_638,N_417,N_441);
and U639 (N_639,N_507,N_496);
nand U640 (N_640,N_583,N_431);
nor U641 (N_641,N_550,N_510);
and U642 (N_642,N_470,N_415);
or U643 (N_643,N_504,N_546);
nand U644 (N_644,N_514,N_416);
and U645 (N_645,N_499,N_422);
and U646 (N_646,N_519,N_530);
and U647 (N_647,N_578,N_528);
xnor U648 (N_648,N_526,N_562);
and U649 (N_649,N_481,N_432);
nor U650 (N_650,N_478,N_535);
xnor U651 (N_651,N_500,N_429);
or U652 (N_652,N_491,N_473);
or U653 (N_653,N_406,N_503);
nor U654 (N_654,N_485,N_466);
and U655 (N_655,N_463,N_559);
nor U656 (N_656,N_482,N_565);
nand U657 (N_657,N_494,N_553);
and U658 (N_658,N_538,N_492);
and U659 (N_659,N_460,N_576);
and U660 (N_660,N_409,N_480);
or U661 (N_661,N_505,N_543);
or U662 (N_662,N_573,N_435);
nand U663 (N_663,N_592,N_407);
or U664 (N_664,N_542,N_414);
nor U665 (N_665,N_418,N_545);
nor U666 (N_666,N_523,N_588);
xnor U667 (N_667,N_541,N_413);
nor U668 (N_668,N_436,N_458);
nand U669 (N_669,N_426,N_591);
and U670 (N_670,N_486,N_584);
nor U671 (N_671,N_438,N_502);
or U672 (N_672,N_456,N_501);
nand U673 (N_673,N_424,N_563);
or U674 (N_674,N_446,N_561);
and U675 (N_675,N_451,N_537);
xnor U676 (N_676,N_569,N_551);
nor U677 (N_677,N_457,N_402);
nand U678 (N_678,N_547,N_558);
and U679 (N_679,N_566,N_590);
or U680 (N_680,N_585,N_479);
nand U681 (N_681,N_581,N_444);
nand U682 (N_682,N_524,N_525);
nor U683 (N_683,N_544,N_453);
xnor U684 (N_684,N_489,N_419);
xor U685 (N_685,N_533,N_434);
nand U686 (N_686,N_512,N_400);
and U687 (N_687,N_513,N_404);
nor U688 (N_688,N_539,N_506);
and U689 (N_689,N_567,N_474);
nand U690 (N_690,N_484,N_597);
and U691 (N_691,N_564,N_593);
xnor U692 (N_692,N_552,N_428);
nand U693 (N_693,N_449,N_574);
nand U694 (N_694,N_433,N_594);
nand U695 (N_695,N_455,N_430);
nand U696 (N_696,N_445,N_488);
nand U697 (N_697,N_421,N_522);
nand U698 (N_698,N_476,N_468);
xnor U699 (N_699,N_517,N_520);
or U700 (N_700,N_569,N_552);
xnor U701 (N_701,N_530,N_534);
nor U702 (N_702,N_407,N_524);
nand U703 (N_703,N_507,N_568);
or U704 (N_704,N_446,N_588);
nand U705 (N_705,N_407,N_576);
xor U706 (N_706,N_595,N_479);
or U707 (N_707,N_526,N_542);
and U708 (N_708,N_494,N_523);
nand U709 (N_709,N_490,N_448);
nand U710 (N_710,N_581,N_556);
or U711 (N_711,N_524,N_505);
or U712 (N_712,N_597,N_475);
and U713 (N_713,N_592,N_472);
nand U714 (N_714,N_509,N_450);
nor U715 (N_715,N_404,N_464);
xor U716 (N_716,N_512,N_452);
and U717 (N_717,N_466,N_543);
nand U718 (N_718,N_442,N_489);
nand U719 (N_719,N_435,N_414);
or U720 (N_720,N_585,N_513);
xnor U721 (N_721,N_577,N_467);
or U722 (N_722,N_453,N_485);
or U723 (N_723,N_568,N_559);
or U724 (N_724,N_552,N_486);
xnor U725 (N_725,N_486,N_429);
nor U726 (N_726,N_441,N_531);
nor U727 (N_727,N_585,N_453);
nor U728 (N_728,N_402,N_515);
or U729 (N_729,N_558,N_594);
nor U730 (N_730,N_508,N_531);
and U731 (N_731,N_454,N_547);
nand U732 (N_732,N_596,N_564);
and U733 (N_733,N_573,N_544);
nand U734 (N_734,N_450,N_571);
nor U735 (N_735,N_471,N_497);
xnor U736 (N_736,N_513,N_570);
and U737 (N_737,N_453,N_507);
and U738 (N_738,N_479,N_488);
nand U739 (N_739,N_405,N_568);
xnor U740 (N_740,N_570,N_430);
or U741 (N_741,N_594,N_412);
nor U742 (N_742,N_540,N_457);
nor U743 (N_743,N_427,N_543);
and U744 (N_744,N_540,N_415);
nor U745 (N_745,N_575,N_537);
nand U746 (N_746,N_473,N_436);
and U747 (N_747,N_505,N_453);
nand U748 (N_748,N_548,N_472);
or U749 (N_749,N_482,N_406);
or U750 (N_750,N_470,N_474);
nor U751 (N_751,N_500,N_478);
xnor U752 (N_752,N_537,N_566);
and U753 (N_753,N_441,N_447);
nand U754 (N_754,N_585,N_593);
or U755 (N_755,N_414,N_588);
xnor U756 (N_756,N_449,N_576);
nor U757 (N_757,N_542,N_499);
nor U758 (N_758,N_424,N_411);
nor U759 (N_759,N_551,N_492);
nand U760 (N_760,N_570,N_424);
nor U761 (N_761,N_490,N_469);
and U762 (N_762,N_401,N_428);
nand U763 (N_763,N_477,N_419);
or U764 (N_764,N_490,N_496);
nand U765 (N_765,N_546,N_596);
nor U766 (N_766,N_548,N_431);
nor U767 (N_767,N_522,N_545);
and U768 (N_768,N_428,N_420);
nand U769 (N_769,N_422,N_463);
nand U770 (N_770,N_457,N_563);
or U771 (N_771,N_447,N_418);
and U772 (N_772,N_437,N_528);
nor U773 (N_773,N_566,N_455);
nor U774 (N_774,N_434,N_459);
or U775 (N_775,N_575,N_536);
nand U776 (N_776,N_414,N_497);
or U777 (N_777,N_448,N_476);
or U778 (N_778,N_529,N_402);
nand U779 (N_779,N_404,N_425);
and U780 (N_780,N_530,N_441);
nor U781 (N_781,N_530,N_483);
or U782 (N_782,N_452,N_491);
nor U783 (N_783,N_446,N_430);
or U784 (N_784,N_426,N_551);
and U785 (N_785,N_461,N_595);
or U786 (N_786,N_552,N_438);
and U787 (N_787,N_493,N_503);
and U788 (N_788,N_455,N_402);
nand U789 (N_789,N_428,N_458);
and U790 (N_790,N_433,N_460);
and U791 (N_791,N_452,N_595);
or U792 (N_792,N_591,N_404);
nand U793 (N_793,N_519,N_584);
xnor U794 (N_794,N_588,N_402);
nand U795 (N_795,N_563,N_499);
and U796 (N_796,N_519,N_552);
xor U797 (N_797,N_544,N_596);
or U798 (N_798,N_472,N_483);
nor U799 (N_799,N_441,N_516);
and U800 (N_800,N_791,N_638);
and U801 (N_801,N_769,N_735);
nand U802 (N_802,N_622,N_651);
nand U803 (N_803,N_716,N_632);
or U804 (N_804,N_705,N_694);
nor U805 (N_805,N_657,N_715);
or U806 (N_806,N_780,N_695);
nor U807 (N_807,N_661,N_795);
nand U808 (N_808,N_720,N_699);
nor U809 (N_809,N_667,N_686);
or U810 (N_810,N_617,N_765);
and U811 (N_811,N_644,N_603);
nor U812 (N_812,N_739,N_799);
xnor U813 (N_813,N_797,N_776);
and U814 (N_814,N_748,N_728);
nand U815 (N_815,N_727,N_767);
and U816 (N_816,N_677,N_750);
and U817 (N_817,N_740,N_680);
nand U818 (N_818,N_764,N_691);
or U819 (N_819,N_736,N_630);
nand U820 (N_820,N_761,N_796);
or U821 (N_821,N_604,N_743);
xor U822 (N_822,N_708,N_671);
xnor U823 (N_823,N_723,N_774);
or U824 (N_824,N_659,N_607);
or U825 (N_825,N_656,N_712);
nor U826 (N_826,N_713,N_654);
nor U827 (N_827,N_717,N_792);
and U828 (N_828,N_786,N_672);
and U829 (N_829,N_729,N_665);
nand U830 (N_830,N_726,N_741);
nor U831 (N_831,N_624,N_790);
nand U832 (N_832,N_636,N_692);
nand U833 (N_833,N_766,N_777);
nor U834 (N_834,N_730,N_754);
xor U835 (N_835,N_623,N_641);
nand U836 (N_836,N_643,N_785);
nor U837 (N_837,N_683,N_724);
or U838 (N_838,N_646,N_778);
nand U839 (N_839,N_605,N_600);
nor U840 (N_840,N_771,N_666);
or U841 (N_841,N_752,N_634);
nor U842 (N_842,N_744,N_710);
and U843 (N_843,N_745,N_709);
or U844 (N_844,N_658,N_606);
nand U845 (N_845,N_633,N_673);
or U846 (N_846,N_649,N_775);
nor U847 (N_847,N_627,N_770);
nor U848 (N_848,N_763,N_663);
or U849 (N_849,N_642,N_782);
nand U850 (N_850,N_609,N_664);
or U851 (N_851,N_614,N_722);
or U852 (N_852,N_616,N_697);
and U853 (N_853,N_685,N_731);
nor U854 (N_854,N_732,N_718);
xor U855 (N_855,N_700,N_652);
and U856 (N_856,N_682,N_681);
or U857 (N_857,N_612,N_679);
or U858 (N_858,N_655,N_719);
and U859 (N_859,N_758,N_611);
nor U860 (N_860,N_690,N_647);
nand U861 (N_861,N_615,N_674);
or U862 (N_862,N_794,N_737);
nand U863 (N_863,N_779,N_698);
nand U864 (N_864,N_601,N_798);
nand U865 (N_865,N_773,N_760);
or U866 (N_866,N_704,N_693);
and U867 (N_867,N_668,N_689);
nor U868 (N_868,N_688,N_670);
or U869 (N_869,N_755,N_703);
and U870 (N_870,N_687,N_621);
and U871 (N_871,N_628,N_706);
and U872 (N_872,N_620,N_678);
nor U873 (N_873,N_640,N_759);
or U874 (N_874,N_619,N_618);
or U875 (N_875,N_707,N_742);
nor U876 (N_876,N_684,N_753);
nand U877 (N_877,N_631,N_783);
nand U878 (N_878,N_746,N_721);
nand U879 (N_879,N_669,N_676);
and U880 (N_880,N_714,N_762);
nand U881 (N_881,N_751,N_639);
and U882 (N_882,N_756,N_701);
nor U883 (N_883,N_608,N_787);
or U884 (N_884,N_747,N_725);
nand U885 (N_885,N_650,N_602);
nand U886 (N_886,N_757,N_772);
nor U887 (N_887,N_696,N_734);
nand U888 (N_888,N_660,N_784);
nand U889 (N_889,N_788,N_702);
or U890 (N_890,N_738,N_626);
nand U891 (N_891,N_653,N_637);
xor U892 (N_892,N_635,N_648);
nand U893 (N_893,N_613,N_610);
nor U894 (N_894,N_749,N_733);
nand U895 (N_895,N_789,N_711);
nand U896 (N_896,N_793,N_768);
and U897 (N_897,N_645,N_625);
or U898 (N_898,N_781,N_675);
nor U899 (N_899,N_662,N_629);
or U900 (N_900,N_610,N_634);
and U901 (N_901,N_758,N_775);
or U902 (N_902,N_792,N_655);
nand U903 (N_903,N_794,N_665);
nor U904 (N_904,N_664,N_779);
nor U905 (N_905,N_627,N_707);
or U906 (N_906,N_617,N_639);
nor U907 (N_907,N_789,N_649);
or U908 (N_908,N_669,N_779);
nand U909 (N_909,N_664,N_784);
nand U910 (N_910,N_638,N_737);
and U911 (N_911,N_743,N_693);
or U912 (N_912,N_781,N_604);
nand U913 (N_913,N_614,N_747);
and U914 (N_914,N_712,N_622);
nand U915 (N_915,N_640,N_714);
nor U916 (N_916,N_725,N_649);
and U917 (N_917,N_650,N_784);
xor U918 (N_918,N_709,N_728);
and U919 (N_919,N_625,N_680);
or U920 (N_920,N_692,N_702);
or U921 (N_921,N_756,N_709);
nor U922 (N_922,N_629,N_709);
xnor U923 (N_923,N_622,N_678);
nand U924 (N_924,N_680,N_663);
nor U925 (N_925,N_799,N_771);
or U926 (N_926,N_603,N_762);
xor U927 (N_927,N_768,N_697);
nor U928 (N_928,N_715,N_701);
or U929 (N_929,N_786,N_605);
nor U930 (N_930,N_744,N_684);
nor U931 (N_931,N_799,N_607);
nand U932 (N_932,N_702,N_682);
and U933 (N_933,N_697,N_663);
or U934 (N_934,N_790,N_698);
and U935 (N_935,N_723,N_741);
nand U936 (N_936,N_790,N_674);
nor U937 (N_937,N_690,N_747);
or U938 (N_938,N_692,N_612);
or U939 (N_939,N_736,N_754);
nand U940 (N_940,N_671,N_747);
nand U941 (N_941,N_782,N_696);
xnor U942 (N_942,N_714,N_708);
and U943 (N_943,N_739,N_613);
nand U944 (N_944,N_604,N_628);
or U945 (N_945,N_613,N_669);
nor U946 (N_946,N_794,N_749);
and U947 (N_947,N_603,N_674);
nor U948 (N_948,N_638,N_607);
nand U949 (N_949,N_635,N_691);
nand U950 (N_950,N_644,N_655);
nor U951 (N_951,N_683,N_620);
xnor U952 (N_952,N_658,N_748);
nand U953 (N_953,N_681,N_779);
and U954 (N_954,N_626,N_646);
xor U955 (N_955,N_621,N_787);
nand U956 (N_956,N_773,N_658);
or U957 (N_957,N_653,N_783);
or U958 (N_958,N_741,N_722);
nand U959 (N_959,N_657,N_731);
or U960 (N_960,N_673,N_774);
or U961 (N_961,N_719,N_622);
nand U962 (N_962,N_704,N_790);
or U963 (N_963,N_672,N_679);
nand U964 (N_964,N_723,N_648);
nor U965 (N_965,N_790,N_693);
nor U966 (N_966,N_682,N_699);
nand U967 (N_967,N_730,N_628);
and U968 (N_968,N_607,N_600);
nor U969 (N_969,N_683,N_656);
and U970 (N_970,N_700,N_786);
nor U971 (N_971,N_663,N_619);
nand U972 (N_972,N_618,N_794);
nand U973 (N_973,N_629,N_620);
or U974 (N_974,N_710,N_772);
and U975 (N_975,N_600,N_715);
and U976 (N_976,N_692,N_780);
xnor U977 (N_977,N_771,N_755);
or U978 (N_978,N_767,N_774);
nand U979 (N_979,N_698,N_602);
nand U980 (N_980,N_694,N_723);
or U981 (N_981,N_686,N_611);
or U982 (N_982,N_722,N_625);
or U983 (N_983,N_671,N_797);
and U984 (N_984,N_789,N_687);
and U985 (N_985,N_626,N_653);
and U986 (N_986,N_688,N_623);
or U987 (N_987,N_768,N_759);
and U988 (N_988,N_770,N_611);
and U989 (N_989,N_639,N_750);
or U990 (N_990,N_650,N_655);
xor U991 (N_991,N_759,N_746);
nand U992 (N_992,N_770,N_636);
nor U993 (N_993,N_654,N_710);
and U994 (N_994,N_740,N_690);
nor U995 (N_995,N_607,N_626);
and U996 (N_996,N_685,N_763);
or U997 (N_997,N_730,N_681);
and U998 (N_998,N_651,N_718);
xnor U999 (N_999,N_678,N_636);
or U1000 (N_1000,N_968,N_928);
or U1001 (N_1001,N_874,N_865);
nand U1002 (N_1002,N_831,N_976);
nor U1003 (N_1003,N_929,N_923);
or U1004 (N_1004,N_944,N_950);
and U1005 (N_1005,N_999,N_926);
nor U1006 (N_1006,N_821,N_924);
or U1007 (N_1007,N_801,N_900);
nor U1008 (N_1008,N_855,N_982);
xnor U1009 (N_1009,N_869,N_861);
nand U1010 (N_1010,N_803,N_812);
nor U1011 (N_1011,N_827,N_818);
and U1012 (N_1012,N_959,N_931);
and U1013 (N_1013,N_962,N_935);
or U1014 (N_1014,N_909,N_899);
or U1015 (N_1015,N_977,N_895);
nand U1016 (N_1016,N_989,N_860);
nand U1017 (N_1017,N_859,N_811);
or U1018 (N_1018,N_921,N_836);
nor U1019 (N_1019,N_823,N_802);
or U1020 (N_1020,N_878,N_907);
or U1021 (N_1021,N_835,N_971);
or U1022 (N_1022,N_882,N_883);
nand U1023 (N_1023,N_941,N_894);
nor U1024 (N_1024,N_996,N_911);
nand U1025 (N_1025,N_912,N_884);
nor U1026 (N_1026,N_913,N_978);
nor U1027 (N_1027,N_858,N_958);
and U1028 (N_1028,N_800,N_914);
nand U1029 (N_1029,N_833,N_892);
or U1030 (N_1030,N_871,N_816);
xnor U1031 (N_1031,N_842,N_930);
or U1032 (N_1032,N_893,N_973);
and U1033 (N_1033,N_870,N_969);
or U1034 (N_1034,N_872,N_938);
or U1035 (N_1035,N_937,N_805);
or U1036 (N_1036,N_980,N_824);
and U1037 (N_1037,N_820,N_804);
and U1038 (N_1038,N_873,N_844);
and U1039 (N_1039,N_970,N_916);
nor U1040 (N_1040,N_940,N_843);
and U1041 (N_1041,N_849,N_898);
nand U1042 (N_1042,N_840,N_974);
nor U1043 (N_1043,N_954,N_987);
nor U1044 (N_1044,N_890,N_879);
nand U1045 (N_1045,N_828,N_813);
or U1046 (N_1046,N_953,N_922);
or U1047 (N_1047,N_965,N_903);
or U1048 (N_1048,N_846,N_994);
nor U1049 (N_1049,N_910,N_942);
or U1050 (N_1050,N_990,N_939);
nand U1051 (N_1051,N_806,N_866);
nor U1052 (N_1052,N_839,N_966);
xnor U1053 (N_1053,N_815,N_810);
nand U1054 (N_1054,N_837,N_850);
xor U1055 (N_1055,N_972,N_960);
nor U1056 (N_1056,N_887,N_863);
xor U1057 (N_1057,N_988,N_955);
or U1058 (N_1058,N_975,N_829);
or U1059 (N_1059,N_952,N_830);
xor U1060 (N_1060,N_908,N_864);
or U1061 (N_1061,N_933,N_904);
nand U1062 (N_1062,N_891,N_979);
or U1063 (N_1063,N_917,N_932);
xnor U1064 (N_1064,N_985,N_817);
or U1065 (N_1065,N_814,N_983);
nor U1066 (N_1066,N_888,N_832);
or U1067 (N_1067,N_822,N_880);
xnor U1068 (N_1068,N_902,N_957);
and U1069 (N_1069,N_877,N_851);
or U1070 (N_1070,N_881,N_834);
nand U1071 (N_1071,N_826,N_915);
or U1072 (N_1072,N_862,N_934);
or U1073 (N_1073,N_956,N_897);
nand U1074 (N_1074,N_868,N_901);
nand U1075 (N_1075,N_946,N_998);
xor U1076 (N_1076,N_925,N_951);
nor U1077 (N_1077,N_905,N_986);
or U1078 (N_1078,N_992,N_876);
or U1079 (N_1079,N_857,N_867);
nand U1080 (N_1080,N_809,N_807);
and U1081 (N_1081,N_886,N_981);
or U1082 (N_1082,N_918,N_943);
nor U1083 (N_1083,N_995,N_964);
nor U1084 (N_1084,N_991,N_838);
nor U1085 (N_1085,N_949,N_945);
nand U1086 (N_1086,N_885,N_967);
xnor U1087 (N_1087,N_853,N_852);
nor U1088 (N_1088,N_896,N_845);
and U1089 (N_1089,N_825,N_906);
nor U1090 (N_1090,N_947,N_963);
or U1091 (N_1091,N_848,N_808);
xor U1092 (N_1092,N_847,N_920);
nand U1093 (N_1093,N_997,N_993);
or U1094 (N_1094,N_854,N_927);
or U1095 (N_1095,N_948,N_841);
or U1096 (N_1096,N_936,N_984);
nor U1097 (N_1097,N_961,N_875);
and U1098 (N_1098,N_919,N_889);
and U1099 (N_1099,N_819,N_856);
nand U1100 (N_1100,N_862,N_851);
nand U1101 (N_1101,N_918,N_885);
or U1102 (N_1102,N_973,N_999);
nand U1103 (N_1103,N_834,N_913);
nand U1104 (N_1104,N_925,N_823);
nor U1105 (N_1105,N_924,N_801);
and U1106 (N_1106,N_983,N_836);
and U1107 (N_1107,N_840,N_846);
and U1108 (N_1108,N_909,N_876);
nand U1109 (N_1109,N_945,N_963);
and U1110 (N_1110,N_837,N_932);
nor U1111 (N_1111,N_933,N_838);
or U1112 (N_1112,N_839,N_993);
and U1113 (N_1113,N_892,N_807);
or U1114 (N_1114,N_974,N_870);
nor U1115 (N_1115,N_952,N_810);
xor U1116 (N_1116,N_967,N_964);
and U1117 (N_1117,N_823,N_851);
nor U1118 (N_1118,N_989,N_936);
nand U1119 (N_1119,N_906,N_969);
nand U1120 (N_1120,N_872,N_936);
nand U1121 (N_1121,N_878,N_982);
xor U1122 (N_1122,N_831,N_881);
or U1123 (N_1123,N_926,N_893);
and U1124 (N_1124,N_910,N_824);
and U1125 (N_1125,N_929,N_841);
or U1126 (N_1126,N_970,N_972);
and U1127 (N_1127,N_826,N_855);
xnor U1128 (N_1128,N_987,N_831);
nand U1129 (N_1129,N_946,N_899);
nand U1130 (N_1130,N_853,N_991);
or U1131 (N_1131,N_940,N_840);
and U1132 (N_1132,N_947,N_810);
nand U1133 (N_1133,N_935,N_863);
and U1134 (N_1134,N_996,N_821);
nand U1135 (N_1135,N_802,N_860);
nand U1136 (N_1136,N_873,N_882);
xnor U1137 (N_1137,N_900,N_983);
and U1138 (N_1138,N_943,N_979);
nand U1139 (N_1139,N_825,N_967);
and U1140 (N_1140,N_845,N_914);
xnor U1141 (N_1141,N_841,N_818);
nand U1142 (N_1142,N_807,N_812);
or U1143 (N_1143,N_910,N_975);
and U1144 (N_1144,N_833,N_827);
or U1145 (N_1145,N_802,N_903);
nand U1146 (N_1146,N_981,N_820);
nand U1147 (N_1147,N_879,N_931);
or U1148 (N_1148,N_971,N_853);
nand U1149 (N_1149,N_844,N_933);
or U1150 (N_1150,N_828,N_874);
nor U1151 (N_1151,N_822,N_831);
and U1152 (N_1152,N_965,N_845);
xor U1153 (N_1153,N_800,N_926);
xor U1154 (N_1154,N_846,N_959);
nor U1155 (N_1155,N_959,N_801);
or U1156 (N_1156,N_808,N_866);
xor U1157 (N_1157,N_809,N_910);
or U1158 (N_1158,N_912,N_843);
nand U1159 (N_1159,N_810,N_983);
nand U1160 (N_1160,N_928,N_880);
or U1161 (N_1161,N_999,N_988);
nor U1162 (N_1162,N_823,N_880);
or U1163 (N_1163,N_903,N_848);
xor U1164 (N_1164,N_812,N_988);
and U1165 (N_1165,N_905,N_832);
or U1166 (N_1166,N_932,N_891);
and U1167 (N_1167,N_909,N_845);
and U1168 (N_1168,N_978,N_927);
or U1169 (N_1169,N_950,N_831);
or U1170 (N_1170,N_970,N_831);
nor U1171 (N_1171,N_863,N_817);
nand U1172 (N_1172,N_919,N_992);
xnor U1173 (N_1173,N_929,N_997);
or U1174 (N_1174,N_905,N_926);
nand U1175 (N_1175,N_987,N_908);
nand U1176 (N_1176,N_857,N_879);
xor U1177 (N_1177,N_945,N_887);
nor U1178 (N_1178,N_864,N_859);
nand U1179 (N_1179,N_877,N_916);
and U1180 (N_1180,N_826,N_801);
and U1181 (N_1181,N_978,N_856);
or U1182 (N_1182,N_851,N_885);
or U1183 (N_1183,N_942,N_806);
nand U1184 (N_1184,N_858,N_825);
nor U1185 (N_1185,N_965,N_881);
nor U1186 (N_1186,N_931,N_812);
xor U1187 (N_1187,N_894,N_883);
and U1188 (N_1188,N_971,N_973);
nor U1189 (N_1189,N_986,N_893);
and U1190 (N_1190,N_874,N_902);
nand U1191 (N_1191,N_953,N_813);
and U1192 (N_1192,N_826,N_899);
and U1193 (N_1193,N_971,N_883);
nand U1194 (N_1194,N_937,N_833);
nand U1195 (N_1195,N_824,N_946);
and U1196 (N_1196,N_801,N_858);
or U1197 (N_1197,N_969,N_820);
nand U1198 (N_1198,N_984,N_822);
nor U1199 (N_1199,N_818,N_994);
nor U1200 (N_1200,N_1167,N_1072);
or U1201 (N_1201,N_1008,N_1050);
xnor U1202 (N_1202,N_1099,N_1006);
nor U1203 (N_1203,N_1005,N_1137);
or U1204 (N_1204,N_1158,N_1120);
nand U1205 (N_1205,N_1035,N_1121);
or U1206 (N_1206,N_1108,N_1040);
nor U1207 (N_1207,N_1066,N_1053);
xor U1208 (N_1208,N_1179,N_1028);
and U1209 (N_1209,N_1161,N_1139);
nand U1210 (N_1210,N_1188,N_1110);
nand U1211 (N_1211,N_1123,N_1021);
and U1212 (N_1212,N_1163,N_1029);
xor U1213 (N_1213,N_1063,N_1159);
nor U1214 (N_1214,N_1178,N_1140);
and U1215 (N_1215,N_1141,N_1046);
nand U1216 (N_1216,N_1007,N_1042);
or U1217 (N_1217,N_1152,N_1142);
xor U1218 (N_1218,N_1086,N_1165);
nand U1219 (N_1219,N_1034,N_1043);
nand U1220 (N_1220,N_1032,N_1192);
xnor U1221 (N_1221,N_1122,N_1181);
nand U1222 (N_1222,N_1020,N_1107);
and U1223 (N_1223,N_1138,N_1109);
nor U1224 (N_1224,N_1155,N_1001);
and U1225 (N_1225,N_1124,N_1134);
nand U1226 (N_1226,N_1060,N_1116);
nand U1227 (N_1227,N_1030,N_1149);
or U1228 (N_1228,N_1111,N_1198);
nor U1229 (N_1229,N_1164,N_1081);
or U1230 (N_1230,N_1176,N_1027);
or U1231 (N_1231,N_1002,N_1000);
nor U1232 (N_1232,N_1076,N_1173);
and U1233 (N_1233,N_1003,N_1051);
and U1234 (N_1234,N_1045,N_1112);
and U1235 (N_1235,N_1048,N_1185);
xnor U1236 (N_1236,N_1041,N_1074);
or U1237 (N_1237,N_1044,N_1170);
and U1238 (N_1238,N_1118,N_1059);
or U1239 (N_1239,N_1154,N_1102);
nor U1240 (N_1240,N_1071,N_1146);
nor U1241 (N_1241,N_1077,N_1147);
nor U1242 (N_1242,N_1054,N_1017);
xnor U1243 (N_1243,N_1068,N_1130);
nand U1244 (N_1244,N_1153,N_1101);
or U1245 (N_1245,N_1083,N_1055);
and U1246 (N_1246,N_1150,N_1022);
nand U1247 (N_1247,N_1065,N_1199);
and U1248 (N_1248,N_1169,N_1145);
xor U1249 (N_1249,N_1049,N_1067);
nand U1250 (N_1250,N_1160,N_1015);
or U1251 (N_1251,N_1119,N_1057);
xnor U1252 (N_1252,N_1174,N_1196);
nand U1253 (N_1253,N_1187,N_1105);
nand U1254 (N_1254,N_1190,N_1082);
nor U1255 (N_1255,N_1016,N_1106);
nor U1256 (N_1256,N_1056,N_1189);
and U1257 (N_1257,N_1125,N_1097);
or U1258 (N_1258,N_1127,N_1186);
and U1259 (N_1259,N_1151,N_1004);
nand U1260 (N_1260,N_1148,N_1114);
and U1261 (N_1261,N_1024,N_1088);
xnor U1262 (N_1262,N_1031,N_1070);
nand U1263 (N_1263,N_1009,N_1047);
and U1264 (N_1264,N_1085,N_1019);
or U1265 (N_1265,N_1166,N_1018);
nand U1266 (N_1266,N_1144,N_1033);
nor U1267 (N_1267,N_1132,N_1096);
and U1268 (N_1268,N_1094,N_1104);
xor U1269 (N_1269,N_1010,N_1194);
or U1270 (N_1270,N_1103,N_1162);
nand U1271 (N_1271,N_1091,N_1013);
xnor U1272 (N_1272,N_1180,N_1089);
or U1273 (N_1273,N_1090,N_1037);
or U1274 (N_1274,N_1168,N_1062);
and U1275 (N_1275,N_1095,N_1156);
and U1276 (N_1276,N_1079,N_1084);
and U1277 (N_1277,N_1080,N_1026);
and U1278 (N_1278,N_1171,N_1075);
or U1279 (N_1279,N_1184,N_1183);
and U1280 (N_1280,N_1117,N_1175);
nor U1281 (N_1281,N_1023,N_1133);
and U1282 (N_1282,N_1135,N_1038);
and U1283 (N_1283,N_1113,N_1087);
or U1284 (N_1284,N_1128,N_1011);
nand U1285 (N_1285,N_1131,N_1098);
or U1286 (N_1286,N_1025,N_1126);
nand U1287 (N_1287,N_1039,N_1191);
and U1288 (N_1288,N_1193,N_1078);
nor U1289 (N_1289,N_1182,N_1073);
nand U1290 (N_1290,N_1143,N_1014);
nand U1291 (N_1291,N_1115,N_1012);
or U1292 (N_1292,N_1197,N_1157);
and U1293 (N_1293,N_1129,N_1093);
and U1294 (N_1294,N_1069,N_1172);
nor U1295 (N_1295,N_1036,N_1136);
nand U1296 (N_1296,N_1100,N_1061);
and U1297 (N_1297,N_1177,N_1058);
or U1298 (N_1298,N_1064,N_1195);
xnor U1299 (N_1299,N_1092,N_1052);
and U1300 (N_1300,N_1035,N_1161);
nand U1301 (N_1301,N_1174,N_1027);
and U1302 (N_1302,N_1133,N_1038);
nor U1303 (N_1303,N_1162,N_1038);
nor U1304 (N_1304,N_1114,N_1095);
and U1305 (N_1305,N_1082,N_1023);
and U1306 (N_1306,N_1186,N_1152);
or U1307 (N_1307,N_1065,N_1095);
xor U1308 (N_1308,N_1061,N_1164);
xor U1309 (N_1309,N_1065,N_1020);
nor U1310 (N_1310,N_1191,N_1008);
or U1311 (N_1311,N_1038,N_1086);
xnor U1312 (N_1312,N_1113,N_1189);
nor U1313 (N_1313,N_1043,N_1164);
nor U1314 (N_1314,N_1144,N_1006);
and U1315 (N_1315,N_1068,N_1035);
or U1316 (N_1316,N_1135,N_1054);
nand U1317 (N_1317,N_1135,N_1096);
nand U1318 (N_1318,N_1155,N_1161);
nand U1319 (N_1319,N_1089,N_1030);
nand U1320 (N_1320,N_1123,N_1000);
nor U1321 (N_1321,N_1182,N_1175);
nor U1322 (N_1322,N_1019,N_1018);
and U1323 (N_1323,N_1187,N_1127);
xnor U1324 (N_1324,N_1178,N_1037);
nand U1325 (N_1325,N_1145,N_1056);
nand U1326 (N_1326,N_1060,N_1127);
or U1327 (N_1327,N_1007,N_1020);
nand U1328 (N_1328,N_1193,N_1095);
nand U1329 (N_1329,N_1032,N_1005);
nor U1330 (N_1330,N_1023,N_1157);
nor U1331 (N_1331,N_1081,N_1109);
and U1332 (N_1332,N_1188,N_1026);
or U1333 (N_1333,N_1070,N_1034);
nor U1334 (N_1334,N_1108,N_1116);
xnor U1335 (N_1335,N_1120,N_1109);
and U1336 (N_1336,N_1033,N_1087);
and U1337 (N_1337,N_1105,N_1107);
nand U1338 (N_1338,N_1050,N_1185);
or U1339 (N_1339,N_1029,N_1035);
nor U1340 (N_1340,N_1014,N_1039);
nand U1341 (N_1341,N_1131,N_1062);
nor U1342 (N_1342,N_1154,N_1151);
and U1343 (N_1343,N_1063,N_1045);
nor U1344 (N_1344,N_1052,N_1061);
or U1345 (N_1345,N_1191,N_1091);
and U1346 (N_1346,N_1053,N_1062);
or U1347 (N_1347,N_1119,N_1136);
or U1348 (N_1348,N_1166,N_1058);
and U1349 (N_1349,N_1057,N_1126);
nand U1350 (N_1350,N_1054,N_1092);
and U1351 (N_1351,N_1044,N_1006);
nand U1352 (N_1352,N_1064,N_1179);
nor U1353 (N_1353,N_1097,N_1079);
and U1354 (N_1354,N_1033,N_1052);
nand U1355 (N_1355,N_1142,N_1144);
xor U1356 (N_1356,N_1168,N_1152);
nand U1357 (N_1357,N_1055,N_1101);
nor U1358 (N_1358,N_1092,N_1085);
nand U1359 (N_1359,N_1048,N_1153);
and U1360 (N_1360,N_1112,N_1082);
nand U1361 (N_1361,N_1000,N_1191);
or U1362 (N_1362,N_1104,N_1081);
xnor U1363 (N_1363,N_1013,N_1189);
and U1364 (N_1364,N_1085,N_1014);
and U1365 (N_1365,N_1184,N_1071);
or U1366 (N_1366,N_1072,N_1089);
nand U1367 (N_1367,N_1052,N_1004);
nand U1368 (N_1368,N_1071,N_1141);
nor U1369 (N_1369,N_1003,N_1056);
nor U1370 (N_1370,N_1015,N_1074);
or U1371 (N_1371,N_1186,N_1047);
and U1372 (N_1372,N_1162,N_1042);
or U1373 (N_1373,N_1063,N_1177);
and U1374 (N_1374,N_1029,N_1167);
or U1375 (N_1375,N_1139,N_1010);
or U1376 (N_1376,N_1162,N_1086);
nor U1377 (N_1377,N_1196,N_1028);
or U1378 (N_1378,N_1146,N_1191);
or U1379 (N_1379,N_1169,N_1099);
and U1380 (N_1380,N_1006,N_1187);
or U1381 (N_1381,N_1131,N_1138);
nor U1382 (N_1382,N_1100,N_1092);
xor U1383 (N_1383,N_1183,N_1000);
and U1384 (N_1384,N_1170,N_1002);
and U1385 (N_1385,N_1089,N_1071);
nand U1386 (N_1386,N_1022,N_1007);
and U1387 (N_1387,N_1192,N_1128);
and U1388 (N_1388,N_1134,N_1162);
nand U1389 (N_1389,N_1185,N_1055);
nor U1390 (N_1390,N_1158,N_1065);
nor U1391 (N_1391,N_1029,N_1050);
or U1392 (N_1392,N_1044,N_1175);
nand U1393 (N_1393,N_1146,N_1078);
nor U1394 (N_1394,N_1134,N_1139);
xor U1395 (N_1395,N_1001,N_1064);
nand U1396 (N_1396,N_1176,N_1114);
nand U1397 (N_1397,N_1030,N_1082);
xor U1398 (N_1398,N_1183,N_1160);
xnor U1399 (N_1399,N_1025,N_1028);
or U1400 (N_1400,N_1321,N_1202);
nor U1401 (N_1401,N_1285,N_1263);
nand U1402 (N_1402,N_1262,N_1255);
nor U1403 (N_1403,N_1300,N_1247);
nand U1404 (N_1404,N_1391,N_1258);
nand U1405 (N_1405,N_1370,N_1346);
nor U1406 (N_1406,N_1312,N_1292);
nor U1407 (N_1407,N_1315,N_1338);
nor U1408 (N_1408,N_1318,N_1343);
or U1409 (N_1409,N_1261,N_1331);
nor U1410 (N_1410,N_1365,N_1214);
or U1411 (N_1411,N_1220,N_1369);
and U1412 (N_1412,N_1244,N_1273);
nor U1413 (N_1413,N_1265,N_1274);
nor U1414 (N_1414,N_1355,N_1394);
nand U1415 (N_1415,N_1211,N_1282);
xor U1416 (N_1416,N_1382,N_1390);
nand U1417 (N_1417,N_1309,N_1381);
and U1418 (N_1418,N_1277,N_1208);
and U1419 (N_1419,N_1298,N_1389);
and U1420 (N_1420,N_1250,N_1397);
nand U1421 (N_1421,N_1399,N_1325);
or U1422 (N_1422,N_1260,N_1347);
or U1423 (N_1423,N_1305,N_1266);
nand U1424 (N_1424,N_1246,N_1368);
nor U1425 (N_1425,N_1254,N_1230);
and U1426 (N_1426,N_1334,N_1323);
nand U1427 (N_1427,N_1367,N_1299);
nand U1428 (N_1428,N_1294,N_1398);
nor U1429 (N_1429,N_1395,N_1359);
nor U1430 (N_1430,N_1336,N_1295);
xnor U1431 (N_1431,N_1339,N_1362);
or U1432 (N_1432,N_1233,N_1332);
nand U1433 (N_1433,N_1342,N_1311);
nor U1434 (N_1434,N_1363,N_1242);
nor U1435 (N_1435,N_1303,N_1205);
and U1436 (N_1436,N_1270,N_1241);
and U1437 (N_1437,N_1322,N_1240);
or U1438 (N_1438,N_1326,N_1231);
nand U1439 (N_1439,N_1200,N_1207);
and U1440 (N_1440,N_1340,N_1224);
nand U1441 (N_1441,N_1380,N_1375);
or U1442 (N_1442,N_1223,N_1267);
or U1443 (N_1443,N_1280,N_1210);
or U1444 (N_1444,N_1324,N_1269);
and U1445 (N_1445,N_1320,N_1335);
or U1446 (N_1446,N_1286,N_1313);
and U1447 (N_1447,N_1228,N_1287);
and U1448 (N_1448,N_1349,N_1253);
nor U1449 (N_1449,N_1352,N_1364);
xnor U1450 (N_1450,N_1328,N_1226);
nand U1451 (N_1451,N_1354,N_1212);
or U1452 (N_1452,N_1351,N_1206);
nand U1453 (N_1453,N_1304,N_1310);
xor U1454 (N_1454,N_1215,N_1371);
xnor U1455 (N_1455,N_1275,N_1234);
nor U1456 (N_1456,N_1290,N_1232);
and U1457 (N_1457,N_1203,N_1376);
nand U1458 (N_1458,N_1393,N_1356);
nand U1459 (N_1459,N_1392,N_1219);
xor U1460 (N_1460,N_1385,N_1296);
xnor U1461 (N_1461,N_1317,N_1308);
and U1462 (N_1462,N_1307,N_1252);
xor U1463 (N_1463,N_1276,N_1378);
and U1464 (N_1464,N_1377,N_1222);
and U1465 (N_1465,N_1288,N_1204);
or U1466 (N_1466,N_1278,N_1256);
or U1467 (N_1467,N_1345,N_1396);
or U1468 (N_1468,N_1379,N_1357);
and U1469 (N_1469,N_1279,N_1384);
nand U1470 (N_1470,N_1386,N_1209);
xor U1471 (N_1471,N_1201,N_1330);
or U1472 (N_1472,N_1237,N_1239);
nand U1473 (N_1473,N_1344,N_1217);
nor U1474 (N_1474,N_1358,N_1301);
and U1475 (N_1475,N_1272,N_1293);
and U1476 (N_1476,N_1302,N_1264);
nor U1477 (N_1477,N_1248,N_1283);
nand U1478 (N_1478,N_1341,N_1225);
nor U1479 (N_1479,N_1337,N_1383);
nand U1480 (N_1480,N_1271,N_1243);
nand U1481 (N_1481,N_1251,N_1227);
nor U1482 (N_1482,N_1350,N_1327);
nand U1483 (N_1483,N_1216,N_1316);
nand U1484 (N_1484,N_1235,N_1249);
nor U1485 (N_1485,N_1297,N_1218);
nand U1486 (N_1486,N_1361,N_1306);
or U1487 (N_1487,N_1333,N_1329);
or U1488 (N_1488,N_1229,N_1289);
nand U1489 (N_1489,N_1372,N_1257);
nand U1490 (N_1490,N_1213,N_1259);
nand U1491 (N_1491,N_1281,N_1221);
nor U1492 (N_1492,N_1360,N_1387);
and U1493 (N_1493,N_1319,N_1268);
and U1494 (N_1494,N_1291,N_1236);
or U1495 (N_1495,N_1245,N_1388);
nor U1496 (N_1496,N_1374,N_1366);
nor U1497 (N_1497,N_1314,N_1353);
nand U1498 (N_1498,N_1284,N_1238);
nor U1499 (N_1499,N_1348,N_1373);
or U1500 (N_1500,N_1200,N_1248);
or U1501 (N_1501,N_1300,N_1288);
nor U1502 (N_1502,N_1234,N_1209);
nand U1503 (N_1503,N_1380,N_1291);
and U1504 (N_1504,N_1337,N_1220);
or U1505 (N_1505,N_1305,N_1291);
or U1506 (N_1506,N_1292,N_1337);
or U1507 (N_1507,N_1256,N_1296);
nor U1508 (N_1508,N_1251,N_1253);
nor U1509 (N_1509,N_1391,N_1378);
nand U1510 (N_1510,N_1205,N_1345);
or U1511 (N_1511,N_1367,N_1398);
and U1512 (N_1512,N_1236,N_1265);
nor U1513 (N_1513,N_1279,N_1331);
and U1514 (N_1514,N_1344,N_1277);
nor U1515 (N_1515,N_1296,N_1359);
nor U1516 (N_1516,N_1336,N_1275);
or U1517 (N_1517,N_1212,N_1238);
and U1518 (N_1518,N_1261,N_1235);
or U1519 (N_1519,N_1245,N_1369);
or U1520 (N_1520,N_1201,N_1302);
nand U1521 (N_1521,N_1393,N_1286);
nand U1522 (N_1522,N_1263,N_1238);
nand U1523 (N_1523,N_1248,N_1319);
nor U1524 (N_1524,N_1389,N_1290);
and U1525 (N_1525,N_1209,N_1372);
nand U1526 (N_1526,N_1285,N_1245);
xor U1527 (N_1527,N_1336,N_1254);
xnor U1528 (N_1528,N_1365,N_1207);
nor U1529 (N_1529,N_1225,N_1348);
nand U1530 (N_1530,N_1294,N_1354);
nand U1531 (N_1531,N_1266,N_1213);
nor U1532 (N_1532,N_1204,N_1290);
and U1533 (N_1533,N_1219,N_1290);
nand U1534 (N_1534,N_1334,N_1315);
or U1535 (N_1535,N_1316,N_1375);
xnor U1536 (N_1536,N_1220,N_1353);
xnor U1537 (N_1537,N_1334,N_1264);
or U1538 (N_1538,N_1324,N_1268);
nand U1539 (N_1539,N_1240,N_1272);
nand U1540 (N_1540,N_1258,N_1283);
nor U1541 (N_1541,N_1217,N_1296);
xor U1542 (N_1542,N_1335,N_1247);
nor U1543 (N_1543,N_1208,N_1338);
xnor U1544 (N_1544,N_1389,N_1293);
nand U1545 (N_1545,N_1305,N_1315);
and U1546 (N_1546,N_1300,N_1334);
nor U1547 (N_1547,N_1283,N_1252);
and U1548 (N_1548,N_1289,N_1334);
nand U1549 (N_1549,N_1315,N_1286);
and U1550 (N_1550,N_1236,N_1286);
nor U1551 (N_1551,N_1313,N_1314);
or U1552 (N_1552,N_1393,N_1216);
or U1553 (N_1553,N_1256,N_1367);
nand U1554 (N_1554,N_1390,N_1325);
nor U1555 (N_1555,N_1354,N_1225);
nor U1556 (N_1556,N_1299,N_1232);
nor U1557 (N_1557,N_1217,N_1321);
and U1558 (N_1558,N_1290,N_1206);
and U1559 (N_1559,N_1370,N_1296);
and U1560 (N_1560,N_1244,N_1301);
nand U1561 (N_1561,N_1231,N_1362);
or U1562 (N_1562,N_1251,N_1371);
nand U1563 (N_1563,N_1366,N_1222);
nand U1564 (N_1564,N_1214,N_1357);
or U1565 (N_1565,N_1385,N_1337);
nand U1566 (N_1566,N_1326,N_1244);
and U1567 (N_1567,N_1268,N_1282);
and U1568 (N_1568,N_1287,N_1293);
nor U1569 (N_1569,N_1291,N_1320);
and U1570 (N_1570,N_1253,N_1330);
nand U1571 (N_1571,N_1305,N_1221);
and U1572 (N_1572,N_1396,N_1265);
nor U1573 (N_1573,N_1370,N_1263);
nor U1574 (N_1574,N_1237,N_1243);
nor U1575 (N_1575,N_1350,N_1238);
or U1576 (N_1576,N_1216,N_1341);
or U1577 (N_1577,N_1304,N_1217);
and U1578 (N_1578,N_1331,N_1247);
and U1579 (N_1579,N_1225,N_1340);
and U1580 (N_1580,N_1385,N_1307);
nand U1581 (N_1581,N_1219,N_1307);
xor U1582 (N_1582,N_1258,N_1204);
or U1583 (N_1583,N_1352,N_1241);
nor U1584 (N_1584,N_1250,N_1367);
or U1585 (N_1585,N_1348,N_1218);
and U1586 (N_1586,N_1359,N_1362);
or U1587 (N_1587,N_1224,N_1368);
or U1588 (N_1588,N_1346,N_1290);
nor U1589 (N_1589,N_1387,N_1382);
nand U1590 (N_1590,N_1263,N_1272);
and U1591 (N_1591,N_1395,N_1220);
nand U1592 (N_1592,N_1365,N_1324);
or U1593 (N_1593,N_1262,N_1387);
nor U1594 (N_1594,N_1312,N_1315);
and U1595 (N_1595,N_1305,N_1383);
or U1596 (N_1596,N_1235,N_1287);
and U1597 (N_1597,N_1340,N_1349);
nor U1598 (N_1598,N_1267,N_1230);
nand U1599 (N_1599,N_1215,N_1294);
xor U1600 (N_1600,N_1575,N_1472);
or U1601 (N_1601,N_1520,N_1581);
and U1602 (N_1602,N_1462,N_1523);
nand U1603 (N_1603,N_1522,N_1423);
nor U1604 (N_1604,N_1555,N_1441);
and U1605 (N_1605,N_1454,N_1558);
nor U1606 (N_1606,N_1533,N_1501);
and U1607 (N_1607,N_1570,N_1557);
or U1608 (N_1608,N_1416,N_1587);
nand U1609 (N_1609,N_1420,N_1574);
nand U1610 (N_1610,N_1552,N_1485);
and U1611 (N_1611,N_1455,N_1521);
nand U1612 (N_1612,N_1537,N_1516);
and U1613 (N_1613,N_1413,N_1504);
or U1614 (N_1614,N_1493,N_1494);
and U1615 (N_1615,N_1426,N_1512);
nand U1616 (N_1616,N_1590,N_1573);
and U1617 (N_1617,N_1432,N_1459);
xor U1618 (N_1618,N_1466,N_1442);
and U1619 (N_1619,N_1473,N_1599);
and U1620 (N_1620,N_1528,N_1408);
or U1621 (N_1621,N_1484,N_1475);
and U1622 (N_1622,N_1540,N_1443);
and U1623 (N_1623,N_1583,N_1439);
nand U1624 (N_1624,N_1465,N_1591);
or U1625 (N_1625,N_1553,N_1593);
xor U1626 (N_1626,N_1433,N_1403);
or U1627 (N_1627,N_1436,N_1489);
xor U1628 (N_1628,N_1476,N_1486);
nor U1629 (N_1629,N_1487,N_1507);
nor U1630 (N_1630,N_1513,N_1542);
or U1631 (N_1631,N_1425,N_1526);
or U1632 (N_1632,N_1519,N_1577);
nor U1633 (N_1633,N_1479,N_1409);
or U1634 (N_1634,N_1497,N_1500);
nor U1635 (N_1635,N_1576,N_1527);
nor U1636 (N_1636,N_1406,N_1562);
nor U1637 (N_1637,N_1578,N_1586);
nor U1638 (N_1638,N_1453,N_1598);
and U1639 (N_1639,N_1474,N_1518);
nand U1640 (N_1640,N_1596,N_1414);
or U1641 (N_1641,N_1421,N_1588);
or U1642 (N_1642,N_1410,N_1511);
or U1643 (N_1643,N_1402,N_1450);
and U1644 (N_1644,N_1452,N_1424);
and U1645 (N_1645,N_1422,N_1415);
nand U1646 (N_1646,N_1505,N_1571);
nor U1647 (N_1647,N_1449,N_1546);
or U1648 (N_1648,N_1404,N_1429);
and U1649 (N_1649,N_1490,N_1503);
nor U1650 (N_1650,N_1529,N_1531);
and U1651 (N_1651,N_1594,N_1534);
xnor U1652 (N_1652,N_1483,N_1556);
nand U1653 (N_1653,N_1464,N_1440);
nor U1654 (N_1654,N_1538,N_1417);
xnor U1655 (N_1655,N_1400,N_1480);
nor U1656 (N_1656,N_1515,N_1477);
nand U1657 (N_1657,N_1506,N_1547);
nor U1658 (N_1658,N_1458,N_1580);
nor U1659 (N_1659,N_1498,N_1549);
xor U1660 (N_1660,N_1446,N_1456);
and U1661 (N_1661,N_1524,N_1595);
or U1662 (N_1662,N_1569,N_1457);
and U1663 (N_1663,N_1563,N_1509);
nand U1664 (N_1664,N_1438,N_1469);
or U1665 (N_1665,N_1514,N_1565);
and U1666 (N_1666,N_1428,N_1418);
nor U1667 (N_1667,N_1496,N_1585);
xnor U1668 (N_1668,N_1460,N_1427);
nand U1669 (N_1669,N_1434,N_1437);
nor U1670 (N_1670,N_1405,N_1589);
or U1671 (N_1671,N_1544,N_1510);
xor U1672 (N_1672,N_1541,N_1543);
or U1673 (N_1673,N_1582,N_1592);
and U1674 (N_1674,N_1502,N_1597);
nor U1675 (N_1675,N_1564,N_1431);
nand U1676 (N_1676,N_1584,N_1430);
or U1677 (N_1677,N_1447,N_1419);
or U1678 (N_1678,N_1461,N_1435);
nor U1679 (N_1679,N_1470,N_1579);
nand U1680 (N_1680,N_1401,N_1567);
or U1681 (N_1681,N_1482,N_1445);
and U1682 (N_1682,N_1451,N_1532);
xor U1683 (N_1683,N_1478,N_1535);
nor U1684 (N_1684,N_1491,N_1554);
or U1685 (N_1685,N_1467,N_1551);
and U1686 (N_1686,N_1572,N_1463);
and U1687 (N_1687,N_1561,N_1550);
nor U1688 (N_1688,N_1488,N_1495);
and U1689 (N_1689,N_1545,N_1499);
nand U1690 (N_1690,N_1412,N_1411);
or U1691 (N_1691,N_1448,N_1530);
nor U1692 (N_1692,N_1536,N_1471);
nor U1693 (N_1693,N_1508,N_1566);
and U1694 (N_1694,N_1517,N_1468);
and U1695 (N_1695,N_1444,N_1525);
or U1696 (N_1696,N_1481,N_1568);
nor U1697 (N_1697,N_1559,N_1560);
and U1698 (N_1698,N_1407,N_1492);
nand U1699 (N_1699,N_1548,N_1539);
nor U1700 (N_1700,N_1507,N_1430);
nor U1701 (N_1701,N_1527,N_1459);
nor U1702 (N_1702,N_1411,N_1497);
xnor U1703 (N_1703,N_1539,N_1440);
and U1704 (N_1704,N_1536,N_1503);
nor U1705 (N_1705,N_1532,N_1456);
and U1706 (N_1706,N_1474,N_1538);
and U1707 (N_1707,N_1552,N_1491);
or U1708 (N_1708,N_1569,N_1498);
nand U1709 (N_1709,N_1596,N_1500);
nand U1710 (N_1710,N_1534,N_1558);
or U1711 (N_1711,N_1492,N_1421);
xnor U1712 (N_1712,N_1506,N_1494);
xnor U1713 (N_1713,N_1586,N_1559);
or U1714 (N_1714,N_1585,N_1512);
nor U1715 (N_1715,N_1520,N_1555);
nor U1716 (N_1716,N_1512,N_1565);
or U1717 (N_1717,N_1540,N_1565);
nand U1718 (N_1718,N_1523,N_1548);
and U1719 (N_1719,N_1544,N_1582);
nor U1720 (N_1720,N_1598,N_1471);
nand U1721 (N_1721,N_1455,N_1585);
nor U1722 (N_1722,N_1594,N_1464);
nand U1723 (N_1723,N_1578,N_1415);
nor U1724 (N_1724,N_1409,N_1595);
nand U1725 (N_1725,N_1448,N_1547);
and U1726 (N_1726,N_1476,N_1496);
nor U1727 (N_1727,N_1499,N_1523);
nor U1728 (N_1728,N_1410,N_1498);
nand U1729 (N_1729,N_1544,N_1580);
xnor U1730 (N_1730,N_1587,N_1420);
and U1731 (N_1731,N_1497,N_1585);
or U1732 (N_1732,N_1536,N_1492);
nor U1733 (N_1733,N_1404,N_1555);
nand U1734 (N_1734,N_1464,N_1563);
nor U1735 (N_1735,N_1541,N_1575);
nand U1736 (N_1736,N_1569,N_1535);
xor U1737 (N_1737,N_1415,N_1557);
nor U1738 (N_1738,N_1516,N_1594);
or U1739 (N_1739,N_1457,N_1483);
or U1740 (N_1740,N_1425,N_1586);
nor U1741 (N_1741,N_1413,N_1410);
xnor U1742 (N_1742,N_1587,N_1472);
and U1743 (N_1743,N_1407,N_1454);
nand U1744 (N_1744,N_1513,N_1528);
nor U1745 (N_1745,N_1493,N_1486);
nand U1746 (N_1746,N_1428,N_1415);
and U1747 (N_1747,N_1476,N_1479);
nand U1748 (N_1748,N_1403,N_1461);
or U1749 (N_1749,N_1405,N_1402);
or U1750 (N_1750,N_1519,N_1576);
and U1751 (N_1751,N_1559,N_1451);
nor U1752 (N_1752,N_1485,N_1519);
nand U1753 (N_1753,N_1599,N_1545);
nor U1754 (N_1754,N_1469,N_1585);
and U1755 (N_1755,N_1467,N_1577);
and U1756 (N_1756,N_1539,N_1518);
nand U1757 (N_1757,N_1597,N_1573);
xnor U1758 (N_1758,N_1442,N_1480);
xor U1759 (N_1759,N_1564,N_1490);
and U1760 (N_1760,N_1414,N_1562);
or U1761 (N_1761,N_1460,N_1465);
xor U1762 (N_1762,N_1598,N_1424);
nor U1763 (N_1763,N_1486,N_1467);
or U1764 (N_1764,N_1458,N_1548);
or U1765 (N_1765,N_1489,N_1542);
nand U1766 (N_1766,N_1547,N_1519);
or U1767 (N_1767,N_1539,N_1561);
nand U1768 (N_1768,N_1452,N_1579);
xor U1769 (N_1769,N_1421,N_1433);
xnor U1770 (N_1770,N_1599,N_1489);
nand U1771 (N_1771,N_1451,N_1452);
and U1772 (N_1772,N_1449,N_1571);
nand U1773 (N_1773,N_1573,N_1436);
nand U1774 (N_1774,N_1409,N_1499);
nor U1775 (N_1775,N_1531,N_1536);
and U1776 (N_1776,N_1406,N_1418);
nand U1777 (N_1777,N_1417,N_1518);
or U1778 (N_1778,N_1563,N_1517);
or U1779 (N_1779,N_1423,N_1563);
or U1780 (N_1780,N_1547,N_1512);
xor U1781 (N_1781,N_1519,N_1410);
nand U1782 (N_1782,N_1569,N_1597);
xnor U1783 (N_1783,N_1446,N_1485);
nand U1784 (N_1784,N_1542,N_1432);
nor U1785 (N_1785,N_1450,N_1474);
or U1786 (N_1786,N_1455,N_1506);
xnor U1787 (N_1787,N_1565,N_1482);
nand U1788 (N_1788,N_1477,N_1461);
and U1789 (N_1789,N_1450,N_1596);
or U1790 (N_1790,N_1458,N_1575);
nand U1791 (N_1791,N_1498,N_1519);
nor U1792 (N_1792,N_1467,N_1478);
nand U1793 (N_1793,N_1467,N_1534);
and U1794 (N_1794,N_1457,N_1464);
or U1795 (N_1795,N_1518,N_1467);
nand U1796 (N_1796,N_1530,N_1527);
nand U1797 (N_1797,N_1425,N_1583);
or U1798 (N_1798,N_1560,N_1509);
nor U1799 (N_1799,N_1431,N_1522);
xnor U1800 (N_1800,N_1747,N_1662);
or U1801 (N_1801,N_1731,N_1792);
nand U1802 (N_1802,N_1742,N_1766);
or U1803 (N_1803,N_1713,N_1611);
or U1804 (N_1804,N_1651,N_1667);
nand U1805 (N_1805,N_1695,N_1761);
and U1806 (N_1806,N_1697,N_1607);
and U1807 (N_1807,N_1724,N_1729);
and U1808 (N_1808,N_1613,N_1615);
nand U1809 (N_1809,N_1682,N_1633);
nand U1810 (N_1810,N_1640,N_1658);
and U1811 (N_1811,N_1636,N_1602);
nand U1812 (N_1812,N_1637,N_1630);
nand U1813 (N_1813,N_1641,N_1702);
or U1814 (N_1814,N_1670,N_1751);
nor U1815 (N_1815,N_1764,N_1683);
nor U1816 (N_1816,N_1616,N_1688);
nand U1817 (N_1817,N_1782,N_1626);
nor U1818 (N_1818,N_1696,N_1623);
nor U1819 (N_1819,N_1609,N_1786);
nand U1820 (N_1820,N_1760,N_1690);
nand U1821 (N_1821,N_1627,N_1663);
nand U1822 (N_1822,N_1680,N_1705);
and U1823 (N_1823,N_1784,N_1620);
or U1824 (N_1824,N_1716,N_1733);
or U1825 (N_1825,N_1614,N_1675);
or U1826 (N_1826,N_1700,N_1628);
or U1827 (N_1827,N_1785,N_1650);
nand U1828 (N_1828,N_1798,N_1619);
nor U1829 (N_1829,N_1701,N_1715);
nor U1830 (N_1830,N_1765,N_1612);
or U1831 (N_1831,N_1600,N_1684);
and U1832 (N_1832,N_1638,N_1718);
and U1833 (N_1833,N_1744,N_1754);
xnor U1834 (N_1834,N_1787,N_1645);
nand U1835 (N_1835,N_1677,N_1624);
nor U1836 (N_1836,N_1767,N_1686);
or U1837 (N_1837,N_1692,N_1743);
nor U1838 (N_1838,N_1691,N_1618);
and U1839 (N_1839,N_1750,N_1622);
nor U1840 (N_1840,N_1741,N_1625);
nand U1841 (N_1841,N_1610,N_1781);
nand U1842 (N_1842,N_1770,N_1749);
and U1843 (N_1843,N_1657,N_1779);
and U1844 (N_1844,N_1711,N_1788);
nand U1845 (N_1845,N_1714,N_1706);
and U1846 (N_1846,N_1685,N_1634);
and U1847 (N_1847,N_1762,N_1694);
nor U1848 (N_1848,N_1717,N_1709);
nor U1849 (N_1849,N_1608,N_1652);
or U1850 (N_1850,N_1757,N_1719);
nor U1851 (N_1851,N_1643,N_1725);
xnor U1852 (N_1852,N_1649,N_1654);
nand U1853 (N_1853,N_1606,N_1659);
nor U1854 (N_1854,N_1726,N_1796);
nand U1855 (N_1855,N_1740,N_1669);
nor U1856 (N_1856,N_1672,N_1720);
nand U1857 (N_1857,N_1664,N_1648);
nor U1858 (N_1858,N_1708,N_1689);
nand U1859 (N_1859,N_1769,N_1723);
nand U1860 (N_1860,N_1727,N_1738);
and U1861 (N_1861,N_1730,N_1674);
nor U1862 (N_1862,N_1763,N_1722);
and U1863 (N_1863,N_1794,N_1797);
or U1864 (N_1864,N_1776,N_1728);
and U1865 (N_1865,N_1777,N_1656);
nand U1866 (N_1866,N_1789,N_1721);
nor U1867 (N_1867,N_1737,N_1793);
nand U1868 (N_1868,N_1790,N_1681);
nand U1869 (N_1869,N_1768,N_1687);
nor U1870 (N_1870,N_1707,N_1629);
nand U1871 (N_1871,N_1679,N_1621);
xor U1872 (N_1872,N_1712,N_1732);
or U1873 (N_1873,N_1710,N_1780);
nand U1874 (N_1874,N_1791,N_1774);
or U1875 (N_1875,N_1693,N_1673);
and U1876 (N_1876,N_1655,N_1631);
nand U1877 (N_1877,N_1660,N_1603);
and U1878 (N_1878,N_1604,N_1703);
and U1879 (N_1879,N_1799,N_1783);
and U1880 (N_1880,N_1632,N_1605);
nor U1881 (N_1881,N_1601,N_1676);
xor U1882 (N_1882,N_1739,N_1678);
nand U1883 (N_1883,N_1736,N_1661);
or U1884 (N_1884,N_1745,N_1665);
nor U1885 (N_1885,N_1735,N_1753);
or U1886 (N_1886,N_1759,N_1746);
and U1887 (N_1887,N_1772,N_1647);
and U1888 (N_1888,N_1756,N_1795);
nor U1889 (N_1889,N_1644,N_1699);
nor U1890 (N_1890,N_1671,N_1646);
xor U1891 (N_1891,N_1653,N_1748);
nor U1892 (N_1892,N_1778,N_1775);
nand U1893 (N_1893,N_1773,N_1771);
nand U1894 (N_1894,N_1635,N_1668);
xnor U1895 (N_1895,N_1639,N_1617);
nand U1896 (N_1896,N_1704,N_1734);
xor U1897 (N_1897,N_1758,N_1666);
nand U1898 (N_1898,N_1752,N_1642);
nand U1899 (N_1899,N_1698,N_1755);
or U1900 (N_1900,N_1752,N_1705);
and U1901 (N_1901,N_1698,N_1784);
xor U1902 (N_1902,N_1743,N_1751);
and U1903 (N_1903,N_1718,N_1704);
or U1904 (N_1904,N_1611,N_1663);
or U1905 (N_1905,N_1603,N_1787);
nor U1906 (N_1906,N_1778,N_1787);
and U1907 (N_1907,N_1671,N_1796);
or U1908 (N_1908,N_1761,N_1650);
or U1909 (N_1909,N_1716,N_1784);
nand U1910 (N_1910,N_1630,N_1625);
nor U1911 (N_1911,N_1642,N_1674);
or U1912 (N_1912,N_1609,N_1602);
xor U1913 (N_1913,N_1739,N_1686);
or U1914 (N_1914,N_1783,N_1724);
or U1915 (N_1915,N_1746,N_1711);
nand U1916 (N_1916,N_1661,N_1632);
or U1917 (N_1917,N_1771,N_1665);
or U1918 (N_1918,N_1647,N_1604);
nor U1919 (N_1919,N_1794,N_1791);
and U1920 (N_1920,N_1616,N_1610);
nand U1921 (N_1921,N_1782,N_1622);
nor U1922 (N_1922,N_1688,N_1681);
xor U1923 (N_1923,N_1600,N_1622);
nor U1924 (N_1924,N_1619,N_1765);
nor U1925 (N_1925,N_1758,N_1769);
or U1926 (N_1926,N_1683,N_1699);
nand U1927 (N_1927,N_1774,N_1743);
nand U1928 (N_1928,N_1646,N_1732);
and U1929 (N_1929,N_1679,N_1666);
nor U1930 (N_1930,N_1766,N_1633);
or U1931 (N_1931,N_1604,N_1756);
nor U1932 (N_1932,N_1600,N_1771);
or U1933 (N_1933,N_1770,N_1720);
nand U1934 (N_1934,N_1639,N_1792);
nor U1935 (N_1935,N_1624,N_1667);
xor U1936 (N_1936,N_1725,N_1705);
or U1937 (N_1937,N_1786,N_1671);
or U1938 (N_1938,N_1700,N_1606);
and U1939 (N_1939,N_1649,N_1751);
nor U1940 (N_1940,N_1744,N_1799);
or U1941 (N_1941,N_1619,N_1651);
nor U1942 (N_1942,N_1770,N_1768);
nor U1943 (N_1943,N_1605,N_1650);
nor U1944 (N_1944,N_1636,N_1635);
and U1945 (N_1945,N_1657,N_1682);
nand U1946 (N_1946,N_1600,N_1774);
nor U1947 (N_1947,N_1748,N_1753);
or U1948 (N_1948,N_1749,N_1742);
and U1949 (N_1949,N_1628,N_1618);
nand U1950 (N_1950,N_1649,N_1784);
nor U1951 (N_1951,N_1786,N_1627);
and U1952 (N_1952,N_1600,N_1645);
nand U1953 (N_1953,N_1676,N_1638);
nor U1954 (N_1954,N_1615,N_1766);
xor U1955 (N_1955,N_1670,N_1756);
and U1956 (N_1956,N_1776,N_1723);
and U1957 (N_1957,N_1725,N_1771);
or U1958 (N_1958,N_1685,N_1691);
and U1959 (N_1959,N_1624,N_1646);
and U1960 (N_1960,N_1742,N_1693);
nand U1961 (N_1961,N_1731,N_1729);
and U1962 (N_1962,N_1619,N_1604);
nand U1963 (N_1963,N_1609,N_1667);
nand U1964 (N_1964,N_1725,N_1745);
nor U1965 (N_1965,N_1610,N_1648);
nor U1966 (N_1966,N_1799,N_1787);
and U1967 (N_1967,N_1681,N_1764);
or U1968 (N_1968,N_1784,N_1799);
or U1969 (N_1969,N_1703,N_1624);
nand U1970 (N_1970,N_1667,N_1632);
or U1971 (N_1971,N_1715,N_1618);
nand U1972 (N_1972,N_1690,N_1784);
nor U1973 (N_1973,N_1629,N_1725);
nor U1974 (N_1974,N_1764,N_1657);
nor U1975 (N_1975,N_1772,N_1649);
nand U1976 (N_1976,N_1640,N_1691);
or U1977 (N_1977,N_1624,N_1761);
nand U1978 (N_1978,N_1654,N_1614);
nor U1979 (N_1979,N_1776,N_1623);
or U1980 (N_1980,N_1605,N_1633);
and U1981 (N_1981,N_1647,N_1678);
xor U1982 (N_1982,N_1691,N_1787);
nand U1983 (N_1983,N_1718,N_1758);
nand U1984 (N_1984,N_1633,N_1760);
or U1985 (N_1985,N_1649,N_1663);
and U1986 (N_1986,N_1735,N_1733);
nand U1987 (N_1987,N_1674,N_1685);
nand U1988 (N_1988,N_1662,N_1797);
and U1989 (N_1989,N_1789,N_1736);
xnor U1990 (N_1990,N_1635,N_1723);
nor U1991 (N_1991,N_1768,N_1634);
and U1992 (N_1992,N_1789,N_1607);
nor U1993 (N_1993,N_1761,N_1753);
xnor U1994 (N_1994,N_1622,N_1653);
nor U1995 (N_1995,N_1690,N_1646);
nand U1996 (N_1996,N_1764,N_1640);
nor U1997 (N_1997,N_1618,N_1600);
or U1998 (N_1998,N_1732,N_1673);
nand U1999 (N_1999,N_1709,N_1726);
and U2000 (N_2000,N_1821,N_1800);
nor U2001 (N_2001,N_1868,N_1844);
nor U2002 (N_2002,N_1923,N_1955);
or U2003 (N_2003,N_1948,N_1896);
or U2004 (N_2004,N_1976,N_1910);
or U2005 (N_2005,N_1820,N_1853);
nor U2006 (N_2006,N_1890,N_1857);
nor U2007 (N_2007,N_1850,N_1939);
or U2008 (N_2008,N_1845,N_1804);
nand U2009 (N_2009,N_1993,N_1994);
or U2010 (N_2010,N_1876,N_1995);
or U2011 (N_2011,N_1919,N_1989);
xor U2012 (N_2012,N_1847,N_1832);
and U2013 (N_2013,N_1894,N_1892);
or U2014 (N_2014,N_1932,N_1897);
xor U2015 (N_2015,N_1867,N_1831);
or U2016 (N_2016,N_1991,N_1858);
and U2017 (N_2017,N_1814,N_1986);
and U2018 (N_2018,N_1801,N_1851);
nor U2019 (N_2019,N_1980,N_1972);
nor U2020 (N_2020,N_1975,N_1998);
or U2021 (N_2021,N_1946,N_1865);
nor U2022 (N_2022,N_1913,N_1860);
or U2023 (N_2023,N_1862,N_1873);
and U2024 (N_2024,N_1840,N_1914);
and U2025 (N_2025,N_1916,N_1958);
and U2026 (N_2026,N_1981,N_1918);
nand U2027 (N_2027,N_1816,N_1978);
nand U2028 (N_2028,N_1930,N_1999);
nor U2029 (N_2029,N_1852,N_1912);
nor U2030 (N_2030,N_1979,N_1909);
nor U2031 (N_2031,N_1951,N_1870);
or U2032 (N_2032,N_1974,N_1927);
nand U2033 (N_2033,N_1812,N_1882);
nor U2034 (N_2034,N_1817,N_1823);
nand U2035 (N_2035,N_1849,N_1936);
or U2036 (N_2036,N_1956,N_1926);
or U2037 (N_2037,N_1921,N_1963);
or U2038 (N_2038,N_1997,N_1872);
or U2039 (N_2039,N_1925,N_1859);
and U2040 (N_2040,N_1992,N_1911);
or U2041 (N_2041,N_1815,N_1960);
nor U2042 (N_2042,N_1808,N_1887);
xnor U2043 (N_2043,N_1842,N_1837);
nand U2044 (N_2044,N_1973,N_1889);
and U2045 (N_2045,N_1818,N_1953);
or U2046 (N_2046,N_1898,N_1891);
or U2047 (N_2047,N_1968,N_1877);
and U2048 (N_2048,N_1826,N_1869);
and U2049 (N_2049,N_1985,N_1871);
and U2050 (N_2050,N_1964,N_1824);
and U2051 (N_2051,N_1938,N_1878);
nand U2052 (N_2052,N_1929,N_1885);
nand U2053 (N_2053,N_1966,N_1880);
and U2054 (N_2054,N_1848,N_1983);
and U2055 (N_2055,N_1883,N_1841);
and U2056 (N_2056,N_1987,N_1901);
and U2057 (N_2057,N_1811,N_1954);
xor U2058 (N_2058,N_1990,N_1805);
and U2059 (N_2059,N_1947,N_1866);
and U2060 (N_2060,N_1984,N_1933);
nor U2061 (N_2061,N_1982,N_1917);
nor U2062 (N_2062,N_1920,N_1949);
or U2063 (N_2063,N_1843,N_1950);
nand U2064 (N_2064,N_1996,N_1810);
or U2065 (N_2065,N_1830,N_1846);
nand U2066 (N_2066,N_1904,N_1806);
and U2067 (N_2067,N_1944,N_1934);
and U2068 (N_2068,N_1855,N_1822);
nor U2069 (N_2069,N_1902,N_1819);
nand U2070 (N_2070,N_1893,N_1977);
or U2071 (N_2071,N_1961,N_1856);
nor U2072 (N_2072,N_1924,N_1864);
nand U2073 (N_2073,N_1807,N_1967);
xnor U2074 (N_2074,N_1942,N_1861);
nor U2075 (N_2075,N_1915,N_1941);
xor U2076 (N_2076,N_1881,N_1971);
nor U2077 (N_2077,N_1969,N_1906);
and U2078 (N_2078,N_1863,N_1884);
and U2079 (N_2079,N_1952,N_1833);
or U2080 (N_2080,N_1888,N_1827);
and U2081 (N_2081,N_1922,N_1879);
nand U2082 (N_2082,N_1935,N_1854);
nor U2083 (N_2083,N_1962,N_1931);
xor U2084 (N_2084,N_1813,N_1943);
and U2085 (N_2085,N_1828,N_1945);
nand U2086 (N_2086,N_1940,N_1803);
and U2087 (N_2087,N_1829,N_1886);
nor U2088 (N_2088,N_1928,N_1937);
nand U2089 (N_2089,N_1957,N_1908);
or U2090 (N_2090,N_1905,N_1839);
and U2091 (N_2091,N_1834,N_1874);
xor U2092 (N_2092,N_1802,N_1970);
nor U2093 (N_2093,N_1836,N_1959);
or U2094 (N_2094,N_1835,N_1965);
and U2095 (N_2095,N_1899,N_1809);
and U2096 (N_2096,N_1825,N_1838);
nand U2097 (N_2097,N_1988,N_1900);
nand U2098 (N_2098,N_1907,N_1903);
or U2099 (N_2099,N_1895,N_1875);
nand U2100 (N_2100,N_1934,N_1973);
nand U2101 (N_2101,N_1950,N_1897);
or U2102 (N_2102,N_1924,N_1827);
xnor U2103 (N_2103,N_1966,N_1846);
nor U2104 (N_2104,N_1981,N_1980);
or U2105 (N_2105,N_1908,N_1934);
or U2106 (N_2106,N_1849,N_1959);
and U2107 (N_2107,N_1823,N_1948);
and U2108 (N_2108,N_1817,N_1832);
or U2109 (N_2109,N_1969,N_1840);
or U2110 (N_2110,N_1966,N_1929);
and U2111 (N_2111,N_1801,N_1908);
and U2112 (N_2112,N_1990,N_1856);
or U2113 (N_2113,N_1948,N_1821);
nor U2114 (N_2114,N_1803,N_1814);
nand U2115 (N_2115,N_1816,N_1905);
nor U2116 (N_2116,N_1948,N_1809);
or U2117 (N_2117,N_1985,N_1957);
and U2118 (N_2118,N_1916,N_1952);
nand U2119 (N_2119,N_1945,N_1841);
and U2120 (N_2120,N_1940,N_1953);
nand U2121 (N_2121,N_1976,N_1860);
and U2122 (N_2122,N_1811,N_1993);
nor U2123 (N_2123,N_1804,N_1898);
nand U2124 (N_2124,N_1856,N_1988);
nor U2125 (N_2125,N_1989,N_1906);
nor U2126 (N_2126,N_1961,N_1872);
and U2127 (N_2127,N_1984,N_1915);
nand U2128 (N_2128,N_1855,N_1838);
nand U2129 (N_2129,N_1879,N_1805);
and U2130 (N_2130,N_1988,N_1803);
xor U2131 (N_2131,N_1942,N_1847);
nor U2132 (N_2132,N_1995,N_1832);
nand U2133 (N_2133,N_1923,N_1914);
xor U2134 (N_2134,N_1824,N_1986);
nand U2135 (N_2135,N_1903,N_1808);
nand U2136 (N_2136,N_1819,N_1953);
and U2137 (N_2137,N_1929,N_1999);
nand U2138 (N_2138,N_1927,N_1878);
or U2139 (N_2139,N_1910,N_1836);
nand U2140 (N_2140,N_1859,N_1953);
and U2141 (N_2141,N_1851,N_1889);
nor U2142 (N_2142,N_1981,N_1828);
nor U2143 (N_2143,N_1865,N_1953);
or U2144 (N_2144,N_1968,N_1972);
nor U2145 (N_2145,N_1960,N_1902);
or U2146 (N_2146,N_1825,N_1860);
nor U2147 (N_2147,N_1841,N_1902);
and U2148 (N_2148,N_1965,N_1824);
or U2149 (N_2149,N_1950,N_1982);
or U2150 (N_2150,N_1884,N_1822);
nor U2151 (N_2151,N_1967,N_1932);
or U2152 (N_2152,N_1848,N_1939);
nand U2153 (N_2153,N_1940,N_1827);
or U2154 (N_2154,N_1817,N_1826);
nor U2155 (N_2155,N_1917,N_1928);
nand U2156 (N_2156,N_1851,N_1805);
nor U2157 (N_2157,N_1828,N_1963);
nand U2158 (N_2158,N_1862,N_1906);
nand U2159 (N_2159,N_1844,N_1867);
and U2160 (N_2160,N_1805,N_1827);
or U2161 (N_2161,N_1924,N_1921);
and U2162 (N_2162,N_1804,N_1988);
or U2163 (N_2163,N_1989,N_1963);
nor U2164 (N_2164,N_1877,N_1864);
xor U2165 (N_2165,N_1960,N_1941);
and U2166 (N_2166,N_1884,N_1996);
xnor U2167 (N_2167,N_1971,N_1927);
xnor U2168 (N_2168,N_1966,N_1967);
nor U2169 (N_2169,N_1817,N_1974);
nand U2170 (N_2170,N_1915,N_1865);
nor U2171 (N_2171,N_1908,N_1941);
or U2172 (N_2172,N_1958,N_1831);
or U2173 (N_2173,N_1995,N_1865);
nor U2174 (N_2174,N_1944,N_1933);
nor U2175 (N_2175,N_1883,N_1815);
nand U2176 (N_2176,N_1826,N_1909);
xnor U2177 (N_2177,N_1840,N_1849);
nand U2178 (N_2178,N_1826,N_1999);
or U2179 (N_2179,N_1853,N_1962);
nor U2180 (N_2180,N_1948,N_1832);
nor U2181 (N_2181,N_1893,N_1829);
nand U2182 (N_2182,N_1868,N_1943);
nor U2183 (N_2183,N_1972,N_1811);
nor U2184 (N_2184,N_1850,N_1919);
or U2185 (N_2185,N_1930,N_1991);
xor U2186 (N_2186,N_1820,N_1849);
nor U2187 (N_2187,N_1808,N_1892);
nand U2188 (N_2188,N_1908,N_1915);
xnor U2189 (N_2189,N_1856,N_1942);
or U2190 (N_2190,N_1810,N_1821);
or U2191 (N_2191,N_1925,N_1840);
and U2192 (N_2192,N_1990,N_1898);
xor U2193 (N_2193,N_1948,N_1819);
nor U2194 (N_2194,N_1911,N_1941);
or U2195 (N_2195,N_1933,N_1887);
nor U2196 (N_2196,N_1862,N_1941);
xor U2197 (N_2197,N_1854,N_1995);
nand U2198 (N_2198,N_1800,N_1870);
and U2199 (N_2199,N_1962,N_1923);
nor U2200 (N_2200,N_2151,N_2082);
and U2201 (N_2201,N_2016,N_2083);
and U2202 (N_2202,N_2110,N_2167);
nand U2203 (N_2203,N_2153,N_2126);
nand U2204 (N_2204,N_2028,N_2152);
or U2205 (N_2205,N_2145,N_2056);
and U2206 (N_2206,N_2094,N_2074);
nor U2207 (N_2207,N_2177,N_2007);
or U2208 (N_2208,N_2164,N_2147);
nor U2209 (N_2209,N_2143,N_2071);
nor U2210 (N_2210,N_2024,N_2085);
nor U2211 (N_2211,N_2178,N_2127);
xnor U2212 (N_2212,N_2122,N_2189);
xnor U2213 (N_2213,N_2069,N_2109);
and U2214 (N_2214,N_2101,N_2188);
nand U2215 (N_2215,N_2044,N_2176);
nand U2216 (N_2216,N_2031,N_2088);
and U2217 (N_2217,N_2046,N_2013);
xor U2218 (N_2218,N_2198,N_2113);
xor U2219 (N_2219,N_2165,N_2142);
and U2220 (N_2220,N_2196,N_2084);
nand U2221 (N_2221,N_2146,N_2135);
and U2222 (N_2222,N_2186,N_2040);
and U2223 (N_2223,N_2193,N_2050);
and U2224 (N_2224,N_2080,N_2158);
xnor U2225 (N_2225,N_2062,N_2053);
or U2226 (N_2226,N_2096,N_2163);
or U2227 (N_2227,N_2022,N_2175);
xor U2228 (N_2228,N_2144,N_2138);
nand U2229 (N_2229,N_2045,N_2025);
and U2230 (N_2230,N_2059,N_2141);
and U2231 (N_2231,N_2011,N_2006);
or U2232 (N_2232,N_2012,N_2047);
nor U2233 (N_2233,N_2041,N_2105);
nand U2234 (N_2234,N_2015,N_2183);
nand U2235 (N_2235,N_2184,N_2019);
and U2236 (N_2236,N_2108,N_2095);
nand U2237 (N_2237,N_2150,N_2001);
xnor U2238 (N_2238,N_2195,N_2063);
and U2239 (N_2239,N_2037,N_2118);
nor U2240 (N_2240,N_2087,N_2107);
xnor U2241 (N_2241,N_2170,N_2034);
or U2242 (N_2242,N_2199,N_2134);
and U2243 (N_2243,N_2078,N_2171);
nor U2244 (N_2244,N_2111,N_2077);
or U2245 (N_2245,N_2136,N_2021);
and U2246 (N_2246,N_2039,N_2194);
and U2247 (N_2247,N_2174,N_2057);
nand U2248 (N_2248,N_2058,N_2002);
nand U2249 (N_2249,N_2156,N_2020);
xnor U2250 (N_2250,N_2067,N_2098);
and U2251 (N_2251,N_2173,N_2003);
nand U2252 (N_2252,N_2191,N_2115);
nand U2253 (N_2253,N_2090,N_2159);
or U2254 (N_2254,N_2099,N_2154);
nand U2255 (N_2255,N_2155,N_2157);
and U2256 (N_2256,N_2131,N_2097);
and U2257 (N_2257,N_2168,N_2180);
and U2258 (N_2258,N_2181,N_2149);
nor U2259 (N_2259,N_2075,N_2102);
and U2260 (N_2260,N_2124,N_2120);
and U2261 (N_2261,N_2166,N_2086);
or U2262 (N_2262,N_2051,N_2119);
nor U2263 (N_2263,N_2192,N_2000);
nor U2264 (N_2264,N_2065,N_2029);
xnor U2265 (N_2265,N_2161,N_2018);
nor U2266 (N_2266,N_2140,N_2005);
or U2267 (N_2267,N_2017,N_2103);
nand U2268 (N_2268,N_2060,N_2148);
nand U2269 (N_2269,N_2117,N_2190);
or U2270 (N_2270,N_2010,N_2089);
nor U2271 (N_2271,N_2133,N_2100);
and U2272 (N_2272,N_2023,N_2076);
or U2273 (N_2273,N_2123,N_2014);
nand U2274 (N_2274,N_2137,N_2032);
or U2275 (N_2275,N_2081,N_2172);
xnor U2276 (N_2276,N_2061,N_2038);
nor U2277 (N_2277,N_2129,N_2197);
or U2278 (N_2278,N_2116,N_2008);
nand U2279 (N_2279,N_2030,N_2027);
and U2280 (N_2280,N_2066,N_2091);
nor U2281 (N_2281,N_2182,N_2125);
xor U2282 (N_2282,N_2064,N_2072);
nor U2283 (N_2283,N_2049,N_2162);
and U2284 (N_2284,N_2187,N_2112);
nand U2285 (N_2285,N_2121,N_2160);
or U2286 (N_2286,N_2004,N_2054);
or U2287 (N_2287,N_2128,N_2033);
and U2288 (N_2288,N_2042,N_2026);
nor U2289 (N_2289,N_2179,N_2055);
and U2290 (N_2290,N_2130,N_2092);
nor U2291 (N_2291,N_2106,N_2132);
xnor U2292 (N_2292,N_2009,N_2052);
nand U2293 (N_2293,N_2104,N_2043);
nand U2294 (N_2294,N_2114,N_2036);
and U2295 (N_2295,N_2048,N_2185);
or U2296 (N_2296,N_2169,N_2139);
nor U2297 (N_2297,N_2073,N_2035);
nand U2298 (N_2298,N_2068,N_2070);
nand U2299 (N_2299,N_2093,N_2079);
and U2300 (N_2300,N_2033,N_2048);
or U2301 (N_2301,N_2073,N_2165);
nand U2302 (N_2302,N_2019,N_2118);
nand U2303 (N_2303,N_2001,N_2063);
or U2304 (N_2304,N_2147,N_2101);
nand U2305 (N_2305,N_2019,N_2078);
or U2306 (N_2306,N_2179,N_2119);
and U2307 (N_2307,N_2140,N_2132);
nand U2308 (N_2308,N_2166,N_2000);
or U2309 (N_2309,N_2029,N_2191);
or U2310 (N_2310,N_2150,N_2102);
nand U2311 (N_2311,N_2108,N_2097);
and U2312 (N_2312,N_2088,N_2112);
nor U2313 (N_2313,N_2154,N_2107);
nand U2314 (N_2314,N_2103,N_2003);
or U2315 (N_2315,N_2051,N_2055);
nor U2316 (N_2316,N_2102,N_2117);
or U2317 (N_2317,N_2158,N_2007);
xnor U2318 (N_2318,N_2194,N_2032);
nor U2319 (N_2319,N_2005,N_2085);
nand U2320 (N_2320,N_2078,N_2083);
and U2321 (N_2321,N_2015,N_2180);
xnor U2322 (N_2322,N_2111,N_2025);
or U2323 (N_2323,N_2008,N_2040);
nand U2324 (N_2324,N_2161,N_2090);
and U2325 (N_2325,N_2078,N_2097);
xnor U2326 (N_2326,N_2185,N_2023);
nand U2327 (N_2327,N_2144,N_2048);
nand U2328 (N_2328,N_2141,N_2007);
nand U2329 (N_2329,N_2036,N_2155);
nand U2330 (N_2330,N_2168,N_2008);
nor U2331 (N_2331,N_2087,N_2171);
or U2332 (N_2332,N_2114,N_2086);
nor U2333 (N_2333,N_2154,N_2171);
and U2334 (N_2334,N_2046,N_2038);
and U2335 (N_2335,N_2109,N_2126);
or U2336 (N_2336,N_2148,N_2174);
and U2337 (N_2337,N_2143,N_2028);
nand U2338 (N_2338,N_2111,N_2038);
xnor U2339 (N_2339,N_2097,N_2185);
nor U2340 (N_2340,N_2087,N_2172);
nor U2341 (N_2341,N_2176,N_2107);
or U2342 (N_2342,N_2025,N_2078);
and U2343 (N_2343,N_2068,N_2181);
nand U2344 (N_2344,N_2110,N_2022);
nand U2345 (N_2345,N_2016,N_2111);
xnor U2346 (N_2346,N_2097,N_2018);
nand U2347 (N_2347,N_2052,N_2187);
or U2348 (N_2348,N_2143,N_2037);
and U2349 (N_2349,N_2185,N_2031);
nor U2350 (N_2350,N_2158,N_2028);
xnor U2351 (N_2351,N_2071,N_2187);
and U2352 (N_2352,N_2186,N_2020);
nand U2353 (N_2353,N_2056,N_2037);
and U2354 (N_2354,N_2150,N_2005);
and U2355 (N_2355,N_2195,N_2054);
nand U2356 (N_2356,N_2111,N_2182);
nand U2357 (N_2357,N_2121,N_2151);
and U2358 (N_2358,N_2001,N_2184);
or U2359 (N_2359,N_2014,N_2018);
and U2360 (N_2360,N_2131,N_2196);
nand U2361 (N_2361,N_2137,N_2094);
and U2362 (N_2362,N_2157,N_2045);
nor U2363 (N_2363,N_2110,N_2088);
nor U2364 (N_2364,N_2137,N_2189);
nor U2365 (N_2365,N_2124,N_2073);
xor U2366 (N_2366,N_2170,N_2158);
or U2367 (N_2367,N_2047,N_2035);
nor U2368 (N_2368,N_2068,N_2147);
nor U2369 (N_2369,N_2026,N_2170);
nand U2370 (N_2370,N_2053,N_2076);
or U2371 (N_2371,N_2008,N_2169);
xor U2372 (N_2372,N_2035,N_2044);
or U2373 (N_2373,N_2131,N_2084);
xor U2374 (N_2374,N_2082,N_2023);
nand U2375 (N_2375,N_2000,N_2183);
nor U2376 (N_2376,N_2030,N_2139);
nand U2377 (N_2377,N_2051,N_2167);
xnor U2378 (N_2378,N_2012,N_2144);
or U2379 (N_2379,N_2168,N_2078);
nor U2380 (N_2380,N_2095,N_2002);
xnor U2381 (N_2381,N_2012,N_2197);
nand U2382 (N_2382,N_2028,N_2001);
nand U2383 (N_2383,N_2020,N_2154);
or U2384 (N_2384,N_2076,N_2072);
nor U2385 (N_2385,N_2140,N_2091);
nor U2386 (N_2386,N_2161,N_2097);
or U2387 (N_2387,N_2039,N_2074);
and U2388 (N_2388,N_2085,N_2037);
nor U2389 (N_2389,N_2188,N_2033);
nor U2390 (N_2390,N_2021,N_2152);
nor U2391 (N_2391,N_2101,N_2010);
nand U2392 (N_2392,N_2150,N_2033);
or U2393 (N_2393,N_2172,N_2038);
and U2394 (N_2394,N_2061,N_2125);
and U2395 (N_2395,N_2100,N_2081);
xor U2396 (N_2396,N_2072,N_2002);
and U2397 (N_2397,N_2089,N_2121);
nor U2398 (N_2398,N_2075,N_2177);
and U2399 (N_2399,N_2071,N_2064);
or U2400 (N_2400,N_2335,N_2354);
or U2401 (N_2401,N_2246,N_2261);
and U2402 (N_2402,N_2289,N_2371);
nor U2403 (N_2403,N_2391,N_2216);
xnor U2404 (N_2404,N_2217,N_2324);
xnor U2405 (N_2405,N_2293,N_2303);
or U2406 (N_2406,N_2247,N_2239);
and U2407 (N_2407,N_2250,N_2292);
and U2408 (N_2408,N_2279,N_2361);
xnor U2409 (N_2409,N_2213,N_2257);
and U2410 (N_2410,N_2284,N_2226);
and U2411 (N_2411,N_2328,N_2351);
or U2412 (N_2412,N_2388,N_2294);
nand U2413 (N_2413,N_2364,N_2270);
nand U2414 (N_2414,N_2368,N_2278);
and U2415 (N_2415,N_2398,N_2314);
and U2416 (N_2416,N_2206,N_2382);
and U2417 (N_2417,N_2343,N_2298);
or U2418 (N_2418,N_2297,N_2287);
or U2419 (N_2419,N_2262,N_2258);
nand U2420 (N_2420,N_2367,N_2353);
nor U2421 (N_2421,N_2394,N_2393);
or U2422 (N_2422,N_2363,N_2295);
and U2423 (N_2423,N_2340,N_2265);
nor U2424 (N_2424,N_2319,N_2268);
nand U2425 (N_2425,N_2288,N_2224);
and U2426 (N_2426,N_2307,N_2330);
or U2427 (N_2427,N_2241,N_2357);
and U2428 (N_2428,N_2329,N_2325);
xnor U2429 (N_2429,N_2286,N_2327);
or U2430 (N_2430,N_2267,N_2221);
xor U2431 (N_2431,N_2338,N_2304);
xor U2432 (N_2432,N_2211,N_2225);
and U2433 (N_2433,N_2390,N_2399);
nor U2434 (N_2434,N_2299,N_2263);
nand U2435 (N_2435,N_2227,N_2240);
nand U2436 (N_2436,N_2296,N_2210);
and U2437 (N_2437,N_2312,N_2272);
or U2438 (N_2438,N_2385,N_2396);
or U2439 (N_2439,N_2311,N_2315);
nor U2440 (N_2440,N_2281,N_2362);
nor U2441 (N_2441,N_2233,N_2234);
nor U2442 (N_2442,N_2342,N_2229);
and U2443 (N_2443,N_2280,N_2337);
nand U2444 (N_2444,N_2208,N_2242);
nor U2445 (N_2445,N_2231,N_2223);
xnor U2446 (N_2446,N_2245,N_2238);
xor U2447 (N_2447,N_2259,N_2379);
and U2448 (N_2448,N_2256,N_2318);
or U2449 (N_2449,N_2222,N_2277);
nor U2450 (N_2450,N_2260,N_2341);
xnor U2451 (N_2451,N_2271,N_2283);
or U2452 (N_2452,N_2269,N_2360);
and U2453 (N_2453,N_2290,N_2285);
xor U2454 (N_2454,N_2384,N_2321);
and U2455 (N_2455,N_2306,N_2346);
or U2456 (N_2456,N_2202,N_2282);
nand U2457 (N_2457,N_2235,N_2365);
nand U2458 (N_2458,N_2331,N_2322);
xor U2459 (N_2459,N_2344,N_2317);
nor U2460 (N_2460,N_2205,N_2326);
nand U2461 (N_2461,N_2214,N_2301);
nand U2462 (N_2462,N_2300,N_2236);
nor U2463 (N_2463,N_2266,N_2249);
and U2464 (N_2464,N_2219,N_2203);
or U2465 (N_2465,N_2308,N_2358);
nor U2466 (N_2466,N_2370,N_2392);
nand U2467 (N_2467,N_2252,N_2209);
nand U2468 (N_2468,N_2276,N_2383);
nor U2469 (N_2469,N_2200,N_2355);
and U2470 (N_2470,N_2380,N_2359);
or U2471 (N_2471,N_2352,N_2377);
nor U2472 (N_2472,N_2372,N_2356);
nor U2473 (N_2473,N_2373,N_2204);
nor U2474 (N_2474,N_2323,N_2349);
xor U2475 (N_2475,N_2248,N_2395);
nor U2476 (N_2476,N_2339,N_2369);
nand U2477 (N_2477,N_2273,N_2305);
nor U2478 (N_2478,N_2378,N_2264);
nor U2479 (N_2479,N_2386,N_2251);
and U2480 (N_2480,N_2255,N_2389);
nor U2481 (N_2481,N_2244,N_2253);
or U2482 (N_2482,N_2345,N_2347);
nor U2483 (N_2483,N_2201,N_2228);
or U2484 (N_2484,N_2275,N_2207);
xnor U2485 (N_2485,N_2215,N_2336);
nor U2486 (N_2486,N_2332,N_2237);
nor U2487 (N_2487,N_2374,N_2291);
nand U2488 (N_2488,N_2309,N_2220);
nand U2489 (N_2489,N_2274,N_2218);
xor U2490 (N_2490,N_2313,N_2334);
nor U2491 (N_2491,N_2302,N_2254);
or U2492 (N_2492,N_2375,N_2381);
nor U2493 (N_2493,N_2243,N_2310);
nor U2494 (N_2494,N_2348,N_2230);
or U2495 (N_2495,N_2376,N_2320);
or U2496 (N_2496,N_2333,N_2366);
or U2497 (N_2497,N_2316,N_2232);
or U2498 (N_2498,N_2397,N_2350);
or U2499 (N_2499,N_2387,N_2212);
and U2500 (N_2500,N_2292,N_2389);
or U2501 (N_2501,N_2256,N_2353);
nor U2502 (N_2502,N_2257,N_2375);
or U2503 (N_2503,N_2257,N_2285);
or U2504 (N_2504,N_2329,N_2362);
nand U2505 (N_2505,N_2290,N_2259);
nor U2506 (N_2506,N_2319,N_2241);
nor U2507 (N_2507,N_2323,N_2363);
or U2508 (N_2508,N_2357,N_2254);
nor U2509 (N_2509,N_2399,N_2331);
xor U2510 (N_2510,N_2342,N_2244);
nor U2511 (N_2511,N_2331,N_2342);
nor U2512 (N_2512,N_2397,N_2282);
nand U2513 (N_2513,N_2249,N_2242);
nor U2514 (N_2514,N_2291,N_2369);
xnor U2515 (N_2515,N_2228,N_2248);
nand U2516 (N_2516,N_2336,N_2255);
or U2517 (N_2517,N_2348,N_2309);
and U2518 (N_2518,N_2390,N_2244);
and U2519 (N_2519,N_2278,N_2339);
or U2520 (N_2520,N_2347,N_2281);
and U2521 (N_2521,N_2240,N_2311);
nand U2522 (N_2522,N_2203,N_2200);
or U2523 (N_2523,N_2248,N_2275);
and U2524 (N_2524,N_2218,N_2370);
nand U2525 (N_2525,N_2268,N_2332);
nor U2526 (N_2526,N_2267,N_2332);
nor U2527 (N_2527,N_2317,N_2353);
nand U2528 (N_2528,N_2219,N_2265);
or U2529 (N_2529,N_2318,N_2290);
or U2530 (N_2530,N_2213,N_2347);
or U2531 (N_2531,N_2360,N_2246);
nand U2532 (N_2532,N_2319,N_2286);
and U2533 (N_2533,N_2291,N_2354);
nand U2534 (N_2534,N_2342,N_2307);
or U2535 (N_2535,N_2342,N_2224);
xor U2536 (N_2536,N_2212,N_2316);
or U2537 (N_2537,N_2230,N_2383);
nor U2538 (N_2538,N_2384,N_2385);
or U2539 (N_2539,N_2294,N_2364);
nor U2540 (N_2540,N_2379,N_2326);
nor U2541 (N_2541,N_2327,N_2205);
nand U2542 (N_2542,N_2390,N_2386);
nor U2543 (N_2543,N_2389,N_2390);
or U2544 (N_2544,N_2397,N_2295);
or U2545 (N_2545,N_2251,N_2277);
nor U2546 (N_2546,N_2246,N_2301);
nor U2547 (N_2547,N_2399,N_2364);
nand U2548 (N_2548,N_2368,N_2212);
or U2549 (N_2549,N_2387,N_2257);
nor U2550 (N_2550,N_2337,N_2237);
and U2551 (N_2551,N_2248,N_2390);
nand U2552 (N_2552,N_2360,N_2332);
and U2553 (N_2553,N_2333,N_2292);
or U2554 (N_2554,N_2209,N_2290);
or U2555 (N_2555,N_2386,N_2374);
xor U2556 (N_2556,N_2359,N_2379);
xnor U2557 (N_2557,N_2306,N_2243);
nor U2558 (N_2558,N_2206,N_2351);
nand U2559 (N_2559,N_2374,N_2262);
or U2560 (N_2560,N_2265,N_2292);
nand U2561 (N_2561,N_2251,N_2222);
nand U2562 (N_2562,N_2275,N_2292);
and U2563 (N_2563,N_2211,N_2285);
nor U2564 (N_2564,N_2266,N_2338);
nand U2565 (N_2565,N_2372,N_2243);
and U2566 (N_2566,N_2234,N_2246);
nor U2567 (N_2567,N_2218,N_2305);
and U2568 (N_2568,N_2375,N_2356);
nand U2569 (N_2569,N_2237,N_2296);
nand U2570 (N_2570,N_2377,N_2247);
or U2571 (N_2571,N_2334,N_2244);
xnor U2572 (N_2572,N_2255,N_2270);
nand U2573 (N_2573,N_2276,N_2258);
nand U2574 (N_2574,N_2335,N_2374);
nor U2575 (N_2575,N_2320,N_2336);
or U2576 (N_2576,N_2216,N_2330);
and U2577 (N_2577,N_2351,N_2242);
and U2578 (N_2578,N_2251,N_2273);
xnor U2579 (N_2579,N_2251,N_2393);
and U2580 (N_2580,N_2328,N_2391);
or U2581 (N_2581,N_2395,N_2275);
nor U2582 (N_2582,N_2241,N_2341);
and U2583 (N_2583,N_2318,N_2250);
or U2584 (N_2584,N_2331,N_2262);
nand U2585 (N_2585,N_2257,N_2266);
nand U2586 (N_2586,N_2249,N_2394);
and U2587 (N_2587,N_2271,N_2363);
or U2588 (N_2588,N_2323,N_2345);
or U2589 (N_2589,N_2310,N_2301);
or U2590 (N_2590,N_2325,N_2356);
nand U2591 (N_2591,N_2258,N_2385);
nor U2592 (N_2592,N_2205,N_2266);
nand U2593 (N_2593,N_2264,N_2381);
nor U2594 (N_2594,N_2223,N_2382);
nand U2595 (N_2595,N_2389,N_2220);
nand U2596 (N_2596,N_2281,N_2236);
nor U2597 (N_2597,N_2211,N_2385);
or U2598 (N_2598,N_2312,N_2389);
or U2599 (N_2599,N_2238,N_2259);
or U2600 (N_2600,N_2535,N_2437);
or U2601 (N_2601,N_2495,N_2599);
and U2602 (N_2602,N_2428,N_2520);
or U2603 (N_2603,N_2540,N_2410);
nand U2604 (N_2604,N_2567,N_2444);
nor U2605 (N_2605,N_2522,N_2560);
nor U2606 (N_2606,N_2562,N_2506);
and U2607 (N_2607,N_2486,N_2431);
or U2608 (N_2608,N_2504,N_2448);
nand U2609 (N_2609,N_2490,N_2566);
or U2610 (N_2610,N_2581,N_2571);
or U2611 (N_2611,N_2467,N_2422);
and U2612 (N_2612,N_2469,N_2425);
or U2613 (N_2613,N_2528,N_2510);
nor U2614 (N_2614,N_2589,N_2430);
nor U2615 (N_2615,N_2439,N_2508);
and U2616 (N_2616,N_2434,N_2572);
and U2617 (N_2617,N_2468,N_2565);
nand U2618 (N_2618,N_2505,N_2408);
or U2619 (N_2619,N_2512,N_2597);
nand U2620 (N_2620,N_2554,N_2543);
and U2621 (N_2621,N_2534,N_2471);
or U2622 (N_2622,N_2523,N_2484);
nand U2623 (N_2623,N_2474,N_2545);
nor U2624 (N_2624,N_2438,N_2558);
nand U2625 (N_2625,N_2532,N_2501);
and U2626 (N_2626,N_2524,N_2582);
and U2627 (N_2627,N_2452,N_2514);
and U2628 (N_2628,N_2577,N_2497);
nand U2629 (N_2629,N_2449,N_2480);
xor U2630 (N_2630,N_2406,N_2450);
or U2631 (N_2631,N_2461,N_2433);
and U2632 (N_2632,N_2479,N_2441);
nor U2633 (N_2633,N_2592,N_2584);
xnor U2634 (N_2634,N_2455,N_2503);
and U2635 (N_2635,N_2412,N_2570);
nand U2636 (N_2636,N_2550,N_2487);
nor U2637 (N_2637,N_2458,N_2456);
nor U2638 (N_2638,N_2411,N_2556);
and U2639 (N_2639,N_2546,N_2473);
or U2640 (N_2640,N_2518,N_2419);
nand U2641 (N_2641,N_2579,N_2553);
xnor U2642 (N_2642,N_2541,N_2521);
and U2643 (N_2643,N_2472,N_2516);
or U2644 (N_2644,N_2513,N_2594);
or U2645 (N_2645,N_2586,N_2475);
nor U2646 (N_2646,N_2426,N_2561);
nor U2647 (N_2647,N_2563,N_2493);
nor U2648 (N_2648,N_2407,N_2537);
and U2649 (N_2649,N_2440,N_2421);
nand U2650 (N_2650,N_2445,N_2574);
and U2651 (N_2651,N_2551,N_2402);
nand U2652 (N_2652,N_2557,N_2464);
nand U2653 (N_2653,N_2466,N_2446);
and U2654 (N_2654,N_2416,N_2498);
nand U2655 (N_2655,N_2559,N_2596);
nand U2656 (N_2656,N_2588,N_2488);
nor U2657 (N_2657,N_2519,N_2485);
nand U2658 (N_2658,N_2568,N_2401);
xor U2659 (N_2659,N_2549,N_2511);
nand U2660 (N_2660,N_2529,N_2470);
xnor U2661 (N_2661,N_2492,N_2536);
nor U2662 (N_2662,N_2400,N_2491);
nand U2663 (N_2663,N_2526,N_2443);
xor U2664 (N_2664,N_2564,N_2531);
or U2665 (N_2665,N_2548,N_2442);
nor U2666 (N_2666,N_2575,N_2447);
xor U2667 (N_2667,N_2593,N_2457);
nand U2668 (N_2668,N_2569,N_2598);
nor U2669 (N_2669,N_2417,N_2555);
and U2670 (N_2670,N_2415,N_2414);
and U2671 (N_2671,N_2478,N_2404);
nor U2672 (N_2672,N_2576,N_2538);
nand U2673 (N_2673,N_2420,N_2580);
nor U2674 (N_2674,N_2547,N_2403);
xor U2675 (N_2675,N_2413,N_2517);
and U2676 (N_2676,N_2573,N_2423);
nor U2677 (N_2677,N_2482,N_2583);
or U2678 (N_2678,N_2489,N_2496);
or U2679 (N_2679,N_2515,N_2544);
nand U2680 (N_2680,N_2435,N_2451);
nand U2681 (N_2681,N_2585,N_2483);
or U2682 (N_2682,N_2499,N_2595);
nor U2683 (N_2683,N_2481,N_2542);
nand U2684 (N_2684,N_2530,N_2500);
or U2685 (N_2685,N_2591,N_2525);
or U2686 (N_2686,N_2460,N_2587);
or U2687 (N_2687,N_2527,N_2432);
xor U2688 (N_2688,N_2476,N_2436);
and U2689 (N_2689,N_2429,N_2509);
nand U2690 (N_2690,N_2507,N_2424);
and U2691 (N_2691,N_2477,N_2552);
nor U2692 (N_2692,N_2590,N_2494);
or U2693 (N_2693,N_2459,N_2453);
or U2694 (N_2694,N_2409,N_2533);
and U2695 (N_2695,N_2502,N_2462);
and U2696 (N_2696,N_2454,N_2418);
xor U2697 (N_2697,N_2465,N_2427);
nand U2698 (N_2698,N_2578,N_2463);
nand U2699 (N_2699,N_2405,N_2539);
or U2700 (N_2700,N_2563,N_2575);
and U2701 (N_2701,N_2560,N_2462);
or U2702 (N_2702,N_2595,N_2425);
nand U2703 (N_2703,N_2572,N_2576);
xor U2704 (N_2704,N_2457,N_2461);
and U2705 (N_2705,N_2546,N_2586);
and U2706 (N_2706,N_2519,N_2561);
or U2707 (N_2707,N_2530,N_2454);
nand U2708 (N_2708,N_2539,N_2510);
or U2709 (N_2709,N_2484,N_2413);
nand U2710 (N_2710,N_2532,N_2567);
and U2711 (N_2711,N_2596,N_2527);
nand U2712 (N_2712,N_2599,N_2591);
and U2713 (N_2713,N_2416,N_2417);
or U2714 (N_2714,N_2452,N_2505);
nand U2715 (N_2715,N_2509,N_2440);
and U2716 (N_2716,N_2592,N_2425);
nand U2717 (N_2717,N_2598,N_2469);
xnor U2718 (N_2718,N_2474,N_2515);
xnor U2719 (N_2719,N_2417,N_2561);
and U2720 (N_2720,N_2544,N_2464);
or U2721 (N_2721,N_2530,N_2595);
nor U2722 (N_2722,N_2574,N_2462);
or U2723 (N_2723,N_2584,N_2484);
nor U2724 (N_2724,N_2495,N_2509);
xnor U2725 (N_2725,N_2488,N_2508);
and U2726 (N_2726,N_2431,N_2529);
nand U2727 (N_2727,N_2478,N_2461);
and U2728 (N_2728,N_2557,N_2515);
or U2729 (N_2729,N_2460,N_2434);
nor U2730 (N_2730,N_2576,N_2455);
or U2731 (N_2731,N_2459,N_2436);
or U2732 (N_2732,N_2447,N_2581);
nand U2733 (N_2733,N_2476,N_2514);
or U2734 (N_2734,N_2564,N_2483);
xor U2735 (N_2735,N_2462,N_2588);
and U2736 (N_2736,N_2584,N_2558);
and U2737 (N_2737,N_2590,N_2545);
nand U2738 (N_2738,N_2480,N_2494);
and U2739 (N_2739,N_2536,N_2524);
xor U2740 (N_2740,N_2542,N_2430);
and U2741 (N_2741,N_2586,N_2408);
or U2742 (N_2742,N_2519,N_2455);
and U2743 (N_2743,N_2591,N_2446);
xor U2744 (N_2744,N_2496,N_2549);
nand U2745 (N_2745,N_2568,N_2570);
and U2746 (N_2746,N_2545,N_2440);
and U2747 (N_2747,N_2479,N_2537);
nand U2748 (N_2748,N_2514,N_2408);
nand U2749 (N_2749,N_2424,N_2536);
and U2750 (N_2750,N_2477,N_2409);
or U2751 (N_2751,N_2488,N_2512);
and U2752 (N_2752,N_2535,N_2466);
nor U2753 (N_2753,N_2472,N_2596);
nor U2754 (N_2754,N_2592,N_2475);
nor U2755 (N_2755,N_2520,N_2488);
nor U2756 (N_2756,N_2400,N_2410);
nand U2757 (N_2757,N_2412,N_2567);
nor U2758 (N_2758,N_2424,N_2454);
nor U2759 (N_2759,N_2474,N_2572);
and U2760 (N_2760,N_2443,N_2571);
or U2761 (N_2761,N_2426,N_2491);
and U2762 (N_2762,N_2533,N_2559);
nor U2763 (N_2763,N_2537,N_2508);
and U2764 (N_2764,N_2451,N_2480);
or U2765 (N_2765,N_2498,N_2435);
xnor U2766 (N_2766,N_2437,N_2400);
or U2767 (N_2767,N_2496,N_2467);
nor U2768 (N_2768,N_2527,N_2445);
nand U2769 (N_2769,N_2494,N_2455);
xnor U2770 (N_2770,N_2495,N_2411);
xnor U2771 (N_2771,N_2593,N_2559);
nor U2772 (N_2772,N_2593,N_2568);
nand U2773 (N_2773,N_2537,N_2505);
nor U2774 (N_2774,N_2469,N_2405);
nand U2775 (N_2775,N_2434,N_2549);
nand U2776 (N_2776,N_2570,N_2464);
or U2777 (N_2777,N_2563,N_2509);
nor U2778 (N_2778,N_2522,N_2411);
and U2779 (N_2779,N_2463,N_2410);
nand U2780 (N_2780,N_2447,N_2466);
nor U2781 (N_2781,N_2521,N_2442);
nand U2782 (N_2782,N_2556,N_2517);
nor U2783 (N_2783,N_2559,N_2450);
or U2784 (N_2784,N_2534,N_2598);
and U2785 (N_2785,N_2508,N_2464);
nor U2786 (N_2786,N_2438,N_2546);
xnor U2787 (N_2787,N_2551,N_2565);
nand U2788 (N_2788,N_2541,N_2478);
nand U2789 (N_2789,N_2489,N_2402);
and U2790 (N_2790,N_2549,N_2536);
nor U2791 (N_2791,N_2566,N_2573);
nand U2792 (N_2792,N_2411,N_2447);
nand U2793 (N_2793,N_2558,N_2569);
nor U2794 (N_2794,N_2542,N_2575);
and U2795 (N_2795,N_2409,N_2404);
and U2796 (N_2796,N_2419,N_2557);
or U2797 (N_2797,N_2493,N_2595);
or U2798 (N_2798,N_2591,N_2549);
or U2799 (N_2799,N_2467,N_2523);
and U2800 (N_2800,N_2648,N_2745);
or U2801 (N_2801,N_2667,N_2716);
and U2802 (N_2802,N_2755,N_2732);
or U2803 (N_2803,N_2734,N_2616);
xor U2804 (N_2804,N_2737,N_2624);
and U2805 (N_2805,N_2660,N_2721);
and U2806 (N_2806,N_2680,N_2780);
and U2807 (N_2807,N_2735,N_2795);
and U2808 (N_2808,N_2677,N_2672);
nor U2809 (N_2809,N_2767,N_2772);
nor U2810 (N_2810,N_2607,N_2654);
and U2811 (N_2811,N_2738,N_2704);
nor U2812 (N_2812,N_2712,N_2752);
nand U2813 (N_2813,N_2696,N_2643);
nand U2814 (N_2814,N_2601,N_2797);
nor U2815 (N_2815,N_2622,N_2720);
nor U2816 (N_2816,N_2662,N_2671);
nor U2817 (N_2817,N_2787,N_2663);
or U2818 (N_2818,N_2640,N_2610);
and U2819 (N_2819,N_2685,N_2706);
nor U2820 (N_2820,N_2681,N_2626);
nor U2821 (N_2821,N_2705,N_2708);
nor U2822 (N_2822,N_2764,N_2757);
nor U2823 (N_2823,N_2623,N_2760);
or U2824 (N_2824,N_2698,N_2781);
nor U2825 (N_2825,N_2744,N_2668);
xnor U2826 (N_2826,N_2687,N_2665);
nor U2827 (N_2827,N_2620,N_2730);
or U2828 (N_2828,N_2666,N_2639);
nor U2829 (N_2829,N_2707,N_2604);
nand U2830 (N_2830,N_2766,N_2630);
nor U2831 (N_2831,N_2790,N_2778);
nand U2832 (N_2832,N_2633,N_2670);
nand U2833 (N_2833,N_2742,N_2776);
and U2834 (N_2834,N_2692,N_2765);
nand U2835 (N_2835,N_2618,N_2740);
nand U2836 (N_2836,N_2756,N_2689);
or U2837 (N_2837,N_2650,N_2678);
nand U2838 (N_2838,N_2613,N_2686);
and U2839 (N_2839,N_2651,N_2750);
and U2840 (N_2840,N_2621,N_2612);
or U2841 (N_2841,N_2653,N_2729);
nand U2842 (N_2842,N_2602,N_2658);
and U2843 (N_2843,N_2784,N_2635);
nand U2844 (N_2844,N_2632,N_2655);
xnor U2845 (N_2845,N_2701,N_2773);
or U2846 (N_2846,N_2726,N_2682);
and U2847 (N_2847,N_2777,N_2673);
or U2848 (N_2848,N_2679,N_2657);
and U2849 (N_2849,N_2649,N_2774);
nor U2850 (N_2850,N_2748,N_2600);
or U2851 (N_2851,N_2770,N_2644);
nor U2852 (N_2852,N_2746,N_2683);
xor U2853 (N_2853,N_2609,N_2637);
xnor U2854 (N_2854,N_2669,N_2747);
or U2855 (N_2855,N_2647,N_2611);
or U2856 (N_2856,N_2792,N_2645);
or U2857 (N_2857,N_2783,N_2661);
nor U2858 (N_2858,N_2631,N_2606);
nor U2859 (N_2859,N_2718,N_2785);
and U2860 (N_2860,N_2711,N_2736);
and U2861 (N_2861,N_2775,N_2675);
and U2862 (N_2862,N_2768,N_2674);
nand U2863 (N_2863,N_2779,N_2771);
or U2864 (N_2864,N_2652,N_2793);
nand U2865 (N_2865,N_2743,N_2782);
nand U2866 (N_2866,N_2724,N_2614);
nand U2867 (N_2867,N_2625,N_2641);
nand U2868 (N_2868,N_2751,N_2753);
and U2869 (N_2869,N_2754,N_2731);
nand U2870 (N_2870,N_2634,N_2638);
and U2871 (N_2871,N_2700,N_2722);
or U2872 (N_2872,N_2761,N_2791);
or U2873 (N_2873,N_2615,N_2628);
nor U2874 (N_2874,N_2688,N_2741);
or U2875 (N_2875,N_2699,N_2789);
nor U2876 (N_2876,N_2759,N_2715);
and U2877 (N_2877,N_2691,N_2646);
xnor U2878 (N_2878,N_2725,N_2684);
xor U2879 (N_2879,N_2642,N_2723);
or U2880 (N_2880,N_2702,N_2786);
or U2881 (N_2881,N_2627,N_2664);
nor U2882 (N_2882,N_2656,N_2629);
and U2883 (N_2883,N_2758,N_2690);
and U2884 (N_2884,N_2798,N_2727);
nand U2885 (N_2885,N_2703,N_2709);
nor U2886 (N_2886,N_2769,N_2695);
or U2887 (N_2887,N_2693,N_2619);
and U2888 (N_2888,N_2788,N_2717);
and U2889 (N_2889,N_2794,N_2659);
or U2890 (N_2890,N_2739,N_2636);
nor U2891 (N_2891,N_2676,N_2697);
and U2892 (N_2892,N_2714,N_2719);
nor U2893 (N_2893,N_2733,N_2617);
and U2894 (N_2894,N_2605,N_2796);
nand U2895 (N_2895,N_2713,N_2749);
nand U2896 (N_2896,N_2763,N_2710);
and U2897 (N_2897,N_2694,N_2603);
or U2898 (N_2898,N_2762,N_2799);
nand U2899 (N_2899,N_2728,N_2608);
xor U2900 (N_2900,N_2672,N_2706);
or U2901 (N_2901,N_2702,N_2699);
and U2902 (N_2902,N_2621,N_2678);
nand U2903 (N_2903,N_2608,N_2631);
and U2904 (N_2904,N_2756,N_2776);
or U2905 (N_2905,N_2710,N_2656);
or U2906 (N_2906,N_2797,N_2749);
or U2907 (N_2907,N_2704,N_2694);
or U2908 (N_2908,N_2721,N_2799);
xnor U2909 (N_2909,N_2630,N_2634);
nand U2910 (N_2910,N_2678,N_2676);
and U2911 (N_2911,N_2719,N_2779);
xor U2912 (N_2912,N_2674,N_2734);
or U2913 (N_2913,N_2695,N_2721);
nand U2914 (N_2914,N_2612,N_2758);
and U2915 (N_2915,N_2696,N_2637);
or U2916 (N_2916,N_2711,N_2721);
and U2917 (N_2917,N_2732,N_2741);
or U2918 (N_2918,N_2785,N_2641);
nor U2919 (N_2919,N_2772,N_2761);
and U2920 (N_2920,N_2625,N_2603);
or U2921 (N_2921,N_2648,N_2708);
nand U2922 (N_2922,N_2768,N_2792);
nor U2923 (N_2923,N_2633,N_2695);
nand U2924 (N_2924,N_2736,N_2690);
and U2925 (N_2925,N_2693,N_2709);
or U2926 (N_2926,N_2603,N_2624);
nand U2927 (N_2927,N_2725,N_2746);
nand U2928 (N_2928,N_2649,N_2700);
nor U2929 (N_2929,N_2706,N_2799);
or U2930 (N_2930,N_2711,N_2792);
or U2931 (N_2931,N_2634,N_2631);
and U2932 (N_2932,N_2719,N_2602);
nand U2933 (N_2933,N_2796,N_2752);
and U2934 (N_2934,N_2658,N_2747);
and U2935 (N_2935,N_2736,N_2666);
xor U2936 (N_2936,N_2793,N_2763);
and U2937 (N_2937,N_2790,N_2735);
or U2938 (N_2938,N_2725,N_2765);
and U2939 (N_2939,N_2755,N_2716);
and U2940 (N_2940,N_2657,N_2713);
xnor U2941 (N_2941,N_2697,N_2753);
or U2942 (N_2942,N_2694,N_2786);
nand U2943 (N_2943,N_2747,N_2731);
or U2944 (N_2944,N_2794,N_2604);
or U2945 (N_2945,N_2649,N_2664);
nand U2946 (N_2946,N_2603,N_2702);
and U2947 (N_2947,N_2605,N_2628);
nor U2948 (N_2948,N_2600,N_2703);
and U2949 (N_2949,N_2671,N_2767);
nand U2950 (N_2950,N_2778,N_2604);
nor U2951 (N_2951,N_2717,N_2610);
nand U2952 (N_2952,N_2705,N_2613);
or U2953 (N_2953,N_2750,N_2690);
xor U2954 (N_2954,N_2622,N_2740);
nand U2955 (N_2955,N_2604,N_2639);
nor U2956 (N_2956,N_2732,N_2750);
nand U2957 (N_2957,N_2600,N_2737);
and U2958 (N_2958,N_2630,N_2610);
nor U2959 (N_2959,N_2665,N_2736);
and U2960 (N_2960,N_2646,N_2771);
nand U2961 (N_2961,N_2674,N_2711);
nor U2962 (N_2962,N_2751,N_2611);
nand U2963 (N_2963,N_2739,N_2744);
nand U2964 (N_2964,N_2698,N_2747);
and U2965 (N_2965,N_2736,N_2629);
and U2966 (N_2966,N_2746,N_2775);
and U2967 (N_2967,N_2726,N_2629);
and U2968 (N_2968,N_2701,N_2702);
nor U2969 (N_2969,N_2777,N_2705);
nor U2970 (N_2970,N_2776,N_2602);
and U2971 (N_2971,N_2760,N_2656);
nor U2972 (N_2972,N_2683,N_2730);
and U2973 (N_2973,N_2667,N_2740);
or U2974 (N_2974,N_2721,N_2680);
or U2975 (N_2975,N_2729,N_2663);
nor U2976 (N_2976,N_2687,N_2728);
or U2977 (N_2977,N_2693,N_2792);
nand U2978 (N_2978,N_2794,N_2688);
or U2979 (N_2979,N_2606,N_2715);
xor U2980 (N_2980,N_2601,N_2754);
xor U2981 (N_2981,N_2624,N_2756);
and U2982 (N_2982,N_2794,N_2748);
nand U2983 (N_2983,N_2725,N_2666);
nand U2984 (N_2984,N_2725,N_2659);
xor U2985 (N_2985,N_2792,N_2745);
nand U2986 (N_2986,N_2728,N_2767);
nand U2987 (N_2987,N_2670,N_2733);
nand U2988 (N_2988,N_2629,N_2767);
xor U2989 (N_2989,N_2724,N_2607);
nor U2990 (N_2990,N_2657,N_2663);
or U2991 (N_2991,N_2635,N_2658);
and U2992 (N_2992,N_2681,N_2651);
nor U2993 (N_2993,N_2676,N_2601);
or U2994 (N_2994,N_2623,N_2626);
nor U2995 (N_2995,N_2722,N_2621);
nor U2996 (N_2996,N_2633,N_2788);
and U2997 (N_2997,N_2652,N_2759);
nor U2998 (N_2998,N_2644,N_2692);
nand U2999 (N_2999,N_2706,N_2668);
xor UO_0 (O_0,N_2954,N_2974);
or UO_1 (O_1,N_2846,N_2953);
and UO_2 (O_2,N_2961,N_2951);
nand UO_3 (O_3,N_2870,N_2872);
nor UO_4 (O_4,N_2925,N_2835);
nand UO_5 (O_5,N_2917,N_2841);
nor UO_6 (O_6,N_2970,N_2826);
nor UO_7 (O_7,N_2918,N_2849);
nor UO_8 (O_8,N_2831,N_2855);
nor UO_9 (O_9,N_2968,N_2994);
nor UO_10 (O_10,N_2866,N_2914);
nor UO_11 (O_11,N_2889,N_2860);
or UO_12 (O_12,N_2875,N_2977);
xnor UO_13 (O_13,N_2880,N_2833);
nand UO_14 (O_14,N_2922,N_2899);
nand UO_15 (O_15,N_2989,N_2896);
nor UO_16 (O_16,N_2828,N_2965);
and UO_17 (O_17,N_2991,N_2827);
nand UO_18 (O_18,N_2853,N_2840);
nor UO_19 (O_19,N_2924,N_2947);
and UO_20 (O_20,N_2877,N_2851);
or UO_21 (O_21,N_2990,N_2992);
nand UO_22 (O_22,N_2843,N_2823);
or UO_23 (O_23,N_2937,N_2803);
and UO_24 (O_24,N_2816,N_2883);
nand UO_25 (O_25,N_2832,N_2969);
and UO_26 (O_26,N_2857,N_2871);
xor UO_27 (O_27,N_2962,N_2993);
xnor UO_28 (O_28,N_2876,N_2967);
nor UO_29 (O_29,N_2834,N_2906);
xor UO_30 (O_30,N_2988,N_2932);
and UO_31 (O_31,N_2824,N_2890);
and UO_32 (O_32,N_2931,N_2808);
xor UO_33 (O_33,N_2907,N_2905);
and UO_34 (O_34,N_2984,N_2972);
or UO_35 (O_35,N_2874,N_2812);
or UO_36 (O_36,N_2956,N_2935);
and UO_37 (O_37,N_2921,N_2926);
and UO_38 (O_38,N_2838,N_2893);
and UO_39 (O_39,N_2818,N_2847);
nand UO_40 (O_40,N_2882,N_2983);
or UO_41 (O_41,N_2911,N_2930);
nand UO_42 (O_42,N_2819,N_2825);
nor UO_43 (O_43,N_2986,N_2806);
or UO_44 (O_44,N_2815,N_2813);
nand UO_45 (O_45,N_2894,N_2901);
nand UO_46 (O_46,N_2941,N_2801);
nand UO_47 (O_47,N_2936,N_2904);
and UO_48 (O_48,N_2879,N_2915);
and UO_49 (O_49,N_2942,N_2892);
nor UO_50 (O_50,N_2946,N_2934);
or UO_51 (O_51,N_2839,N_2928);
nor UO_52 (O_52,N_2809,N_2878);
and UO_53 (O_53,N_2869,N_2981);
or UO_54 (O_54,N_2944,N_2980);
nand UO_55 (O_55,N_2881,N_2837);
nor UO_56 (O_56,N_2927,N_2933);
nor UO_57 (O_57,N_2845,N_2976);
and UO_58 (O_58,N_2820,N_2959);
xnor UO_59 (O_59,N_2999,N_2957);
or UO_60 (O_60,N_2802,N_2913);
nor UO_61 (O_61,N_2908,N_2963);
or UO_62 (O_62,N_2960,N_2919);
and UO_63 (O_63,N_2997,N_2856);
nand UO_64 (O_64,N_2995,N_2854);
and UO_65 (O_65,N_2943,N_2861);
xnor UO_66 (O_66,N_2949,N_2897);
and UO_67 (O_67,N_2821,N_2966);
and UO_68 (O_68,N_2916,N_2829);
or UO_69 (O_69,N_2863,N_2848);
nor UO_70 (O_70,N_2945,N_2805);
nand UO_71 (O_71,N_2964,N_2888);
nand UO_72 (O_72,N_2887,N_2804);
nor UO_73 (O_73,N_2939,N_2902);
nand UO_74 (O_74,N_2973,N_2891);
nor UO_75 (O_75,N_2884,N_2865);
nor UO_76 (O_76,N_2955,N_2830);
nor UO_77 (O_77,N_2862,N_2822);
and UO_78 (O_78,N_2998,N_2859);
and UO_79 (O_79,N_2950,N_2885);
nand UO_80 (O_80,N_2858,N_2910);
or UO_81 (O_81,N_2920,N_2900);
or UO_82 (O_82,N_2873,N_2886);
nor UO_83 (O_83,N_2912,N_2923);
nand UO_84 (O_84,N_2985,N_2842);
or UO_85 (O_85,N_2810,N_2817);
nor UO_86 (O_86,N_2929,N_2952);
nor UO_87 (O_87,N_2948,N_2807);
and UO_88 (O_88,N_2895,N_2975);
nor UO_89 (O_89,N_2938,N_2996);
xnor UO_90 (O_90,N_2867,N_2814);
nand UO_91 (O_91,N_2987,N_2850);
or UO_92 (O_92,N_2982,N_2844);
nor UO_93 (O_93,N_2958,N_2978);
and UO_94 (O_94,N_2909,N_2898);
nand UO_95 (O_95,N_2852,N_2868);
nor UO_96 (O_96,N_2800,N_2903);
and UO_97 (O_97,N_2979,N_2811);
or UO_98 (O_98,N_2864,N_2971);
or UO_99 (O_99,N_2940,N_2836);
or UO_100 (O_100,N_2921,N_2969);
nand UO_101 (O_101,N_2817,N_2932);
nor UO_102 (O_102,N_2873,N_2839);
nor UO_103 (O_103,N_2974,N_2865);
and UO_104 (O_104,N_2890,N_2884);
nand UO_105 (O_105,N_2830,N_2995);
and UO_106 (O_106,N_2892,N_2971);
or UO_107 (O_107,N_2900,N_2903);
xnor UO_108 (O_108,N_2905,N_2999);
and UO_109 (O_109,N_2955,N_2814);
or UO_110 (O_110,N_2811,N_2987);
or UO_111 (O_111,N_2894,N_2847);
xor UO_112 (O_112,N_2801,N_2936);
nand UO_113 (O_113,N_2861,N_2811);
nand UO_114 (O_114,N_2929,N_2964);
or UO_115 (O_115,N_2973,N_2995);
or UO_116 (O_116,N_2941,N_2884);
nand UO_117 (O_117,N_2817,N_2872);
and UO_118 (O_118,N_2897,N_2898);
nor UO_119 (O_119,N_2815,N_2853);
nand UO_120 (O_120,N_2831,N_2994);
and UO_121 (O_121,N_2870,N_2947);
xnor UO_122 (O_122,N_2820,N_2864);
and UO_123 (O_123,N_2890,N_2819);
nand UO_124 (O_124,N_2949,N_2889);
nand UO_125 (O_125,N_2837,N_2932);
xor UO_126 (O_126,N_2942,N_2976);
or UO_127 (O_127,N_2844,N_2821);
and UO_128 (O_128,N_2929,N_2979);
and UO_129 (O_129,N_2980,N_2995);
nor UO_130 (O_130,N_2940,N_2995);
nand UO_131 (O_131,N_2985,N_2922);
or UO_132 (O_132,N_2831,N_2841);
nand UO_133 (O_133,N_2861,N_2986);
and UO_134 (O_134,N_2885,N_2800);
nand UO_135 (O_135,N_2836,N_2942);
nor UO_136 (O_136,N_2862,N_2874);
nor UO_137 (O_137,N_2837,N_2920);
nor UO_138 (O_138,N_2866,N_2996);
nand UO_139 (O_139,N_2889,N_2947);
nand UO_140 (O_140,N_2910,N_2832);
or UO_141 (O_141,N_2925,N_2813);
or UO_142 (O_142,N_2870,N_2839);
and UO_143 (O_143,N_2812,N_2809);
or UO_144 (O_144,N_2927,N_2852);
nand UO_145 (O_145,N_2904,N_2992);
nand UO_146 (O_146,N_2929,N_2844);
xnor UO_147 (O_147,N_2929,N_2904);
or UO_148 (O_148,N_2825,N_2840);
nor UO_149 (O_149,N_2920,N_2952);
nor UO_150 (O_150,N_2914,N_2901);
and UO_151 (O_151,N_2840,N_2964);
and UO_152 (O_152,N_2923,N_2965);
nand UO_153 (O_153,N_2855,N_2923);
and UO_154 (O_154,N_2915,N_2887);
nor UO_155 (O_155,N_2991,N_2959);
and UO_156 (O_156,N_2843,N_2941);
and UO_157 (O_157,N_2988,N_2989);
and UO_158 (O_158,N_2902,N_2874);
nand UO_159 (O_159,N_2899,N_2855);
and UO_160 (O_160,N_2808,N_2864);
and UO_161 (O_161,N_2849,N_2884);
nand UO_162 (O_162,N_2907,N_2874);
or UO_163 (O_163,N_2919,N_2877);
and UO_164 (O_164,N_2859,N_2885);
nor UO_165 (O_165,N_2887,N_2979);
or UO_166 (O_166,N_2994,N_2987);
nor UO_167 (O_167,N_2848,N_2942);
and UO_168 (O_168,N_2875,N_2825);
nand UO_169 (O_169,N_2875,N_2839);
nand UO_170 (O_170,N_2870,N_2916);
nor UO_171 (O_171,N_2862,N_2948);
nand UO_172 (O_172,N_2991,N_2836);
nand UO_173 (O_173,N_2922,N_2936);
xor UO_174 (O_174,N_2820,N_2926);
and UO_175 (O_175,N_2986,N_2828);
nor UO_176 (O_176,N_2907,N_2925);
nor UO_177 (O_177,N_2822,N_2983);
nor UO_178 (O_178,N_2892,N_2863);
or UO_179 (O_179,N_2971,N_2958);
nor UO_180 (O_180,N_2895,N_2960);
or UO_181 (O_181,N_2984,N_2973);
nor UO_182 (O_182,N_2904,N_2975);
xnor UO_183 (O_183,N_2904,N_2804);
nand UO_184 (O_184,N_2991,N_2907);
nor UO_185 (O_185,N_2877,N_2976);
nor UO_186 (O_186,N_2916,N_2839);
and UO_187 (O_187,N_2955,N_2960);
xor UO_188 (O_188,N_2955,N_2928);
nor UO_189 (O_189,N_2832,N_2875);
or UO_190 (O_190,N_2851,N_2838);
xnor UO_191 (O_191,N_2977,N_2851);
nor UO_192 (O_192,N_2920,N_2983);
xor UO_193 (O_193,N_2848,N_2883);
nor UO_194 (O_194,N_2999,N_2839);
nand UO_195 (O_195,N_2950,N_2857);
nor UO_196 (O_196,N_2960,N_2900);
and UO_197 (O_197,N_2850,N_2923);
nand UO_198 (O_198,N_2807,N_2999);
nand UO_199 (O_199,N_2939,N_2879);
or UO_200 (O_200,N_2989,N_2977);
nor UO_201 (O_201,N_2910,N_2835);
nor UO_202 (O_202,N_2947,N_2825);
xor UO_203 (O_203,N_2836,N_2965);
and UO_204 (O_204,N_2939,N_2913);
nand UO_205 (O_205,N_2950,N_2957);
or UO_206 (O_206,N_2817,N_2954);
and UO_207 (O_207,N_2857,N_2899);
nor UO_208 (O_208,N_2963,N_2949);
nand UO_209 (O_209,N_2820,N_2997);
xnor UO_210 (O_210,N_2933,N_2952);
and UO_211 (O_211,N_2980,N_2843);
nor UO_212 (O_212,N_2918,N_2924);
and UO_213 (O_213,N_2898,N_2851);
xor UO_214 (O_214,N_2945,N_2845);
or UO_215 (O_215,N_2954,N_2921);
nor UO_216 (O_216,N_2976,N_2803);
nor UO_217 (O_217,N_2895,N_2846);
or UO_218 (O_218,N_2808,N_2857);
nand UO_219 (O_219,N_2980,N_2948);
nand UO_220 (O_220,N_2830,N_2871);
or UO_221 (O_221,N_2999,N_2831);
nor UO_222 (O_222,N_2800,N_2862);
and UO_223 (O_223,N_2852,N_2810);
nand UO_224 (O_224,N_2925,N_2822);
and UO_225 (O_225,N_2934,N_2944);
xor UO_226 (O_226,N_2897,N_2984);
nor UO_227 (O_227,N_2891,N_2959);
or UO_228 (O_228,N_2824,N_2983);
nor UO_229 (O_229,N_2818,N_2944);
or UO_230 (O_230,N_2903,N_2824);
nand UO_231 (O_231,N_2924,N_2864);
and UO_232 (O_232,N_2954,N_2842);
and UO_233 (O_233,N_2916,N_2866);
or UO_234 (O_234,N_2943,N_2955);
xnor UO_235 (O_235,N_2953,N_2971);
nand UO_236 (O_236,N_2958,N_2841);
or UO_237 (O_237,N_2950,N_2946);
or UO_238 (O_238,N_2935,N_2951);
and UO_239 (O_239,N_2994,N_2986);
nand UO_240 (O_240,N_2968,N_2898);
nor UO_241 (O_241,N_2812,N_2846);
and UO_242 (O_242,N_2986,N_2991);
and UO_243 (O_243,N_2853,N_2916);
or UO_244 (O_244,N_2853,N_2845);
and UO_245 (O_245,N_2820,N_2865);
nand UO_246 (O_246,N_2968,N_2842);
nand UO_247 (O_247,N_2831,N_2901);
nand UO_248 (O_248,N_2811,N_2866);
or UO_249 (O_249,N_2826,N_2880);
and UO_250 (O_250,N_2899,N_2926);
nand UO_251 (O_251,N_2824,N_2922);
or UO_252 (O_252,N_2969,N_2889);
xnor UO_253 (O_253,N_2880,N_2888);
or UO_254 (O_254,N_2992,N_2815);
nor UO_255 (O_255,N_2906,N_2855);
nand UO_256 (O_256,N_2849,N_2869);
nand UO_257 (O_257,N_2806,N_2888);
nand UO_258 (O_258,N_2827,N_2801);
and UO_259 (O_259,N_2904,N_2876);
nand UO_260 (O_260,N_2847,N_2947);
xnor UO_261 (O_261,N_2859,N_2974);
nor UO_262 (O_262,N_2976,N_2939);
or UO_263 (O_263,N_2897,N_2821);
nor UO_264 (O_264,N_2942,N_2983);
or UO_265 (O_265,N_2977,N_2879);
nor UO_266 (O_266,N_2947,N_2970);
or UO_267 (O_267,N_2832,N_2863);
nand UO_268 (O_268,N_2814,N_2894);
nand UO_269 (O_269,N_2904,N_2875);
or UO_270 (O_270,N_2950,N_2858);
or UO_271 (O_271,N_2838,N_2872);
nor UO_272 (O_272,N_2889,N_2885);
nand UO_273 (O_273,N_2822,N_2953);
and UO_274 (O_274,N_2824,N_2821);
nand UO_275 (O_275,N_2805,N_2803);
nand UO_276 (O_276,N_2925,N_2890);
nor UO_277 (O_277,N_2949,N_2945);
xor UO_278 (O_278,N_2819,N_2943);
nor UO_279 (O_279,N_2930,N_2828);
or UO_280 (O_280,N_2875,N_2870);
nand UO_281 (O_281,N_2812,N_2820);
nand UO_282 (O_282,N_2929,N_2842);
nor UO_283 (O_283,N_2922,N_2972);
and UO_284 (O_284,N_2882,N_2977);
and UO_285 (O_285,N_2862,N_2881);
and UO_286 (O_286,N_2964,N_2987);
nor UO_287 (O_287,N_2933,N_2919);
nand UO_288 (O_288,N_2970,N_2944);
or UO_289 (O_289,N_2986,N_2964);
nand UO_290 (O_290,N_2831,N_2938);
and UO_291 (O_291,N_2869,N_2809);
and UO_292 (O_292,N_2887,N_2968);
nand UO_293 (O_293,N_2980,N_2892);
nand UO_294 (O_294,N_2878,N_2817);
and UO_295 (O_295,N_2978,N_2957);
and UO_296 (O_296,N_2972,N_2876);
xnor UO_297 (O_297,N_2947,N_2984);
and UO_298 (O_298,N_2910,N_2880);
nor UO_299 (O_299,N_2872,N_2825);
nor UO_300 (O_300,N_2910,N_2992);
and UO_301 (O_301,N_2872,N_2816);
nor UO_302 (O_302,N_2943,N_2902);
nor UO_303 (O_303,N_2860,N_2834);
and UO_304 (O_304,N_2864,N_2977);
nand UO_305 (O_305,N_2984,N_2854);
nor UO_306 (O_306,N_2859,N_2994);
nand UO_307 (O_307,N_2827,N_2987);
nor UO_308 (O_308,N_2918,N_2820);
nor UO_309 (O_309,N_2822,N_2872);
xnor UO_310 (O_310,N_2954,N_2991);
xnor UO_311 (O_311,N_2802,N_2910);
nor UO_312 (O_312,N_2945,N_2916);
xnor UO_313 (O_313,N_2929,N_2874);
or UO_314 (O_314,N_2837,N_2925);
or UO_315 (O_315,N_2995,N_2984);
nand UO_316 (O_316,N_2885,N_2905);
nand UO_317 (O_317,N_2832,N_2874);
and UO_318 (O_318,N_2867,N_2859);
and UO_319 (O_319,N_2970,N_2808);
xnor UO_320 (O_320,N_2880,N_2855);
or UO_321 (O_321,N_2882,N_2952);
and UO_322 (O_322,N_2998,N_2830);
or UO_323 (O_323,N_2898,N_2825);
nor UO_324 (O_324,N_2966,N_2868);
or UO_325 (O_325,N_2900,N_2824);
or UO_326 (O_326,N_2800,N_2916);
nor UO_327 (O_327,N_2903,N_2819);
nand UO_328 (O_328,N_2873,N_2918);
nor UO_329 (O_329,N_2883,N_2927);
nand UO_330 (O_330,N_2822,N_2892);
nand UO_331 (O_331,N_2830,N_2835);
or UO_332 (O_332,N_2814,N_2857);
and UO_333 (O_333,N_2899,N_2928);
nand UO_334 (O_334,N_2856,N_2887);
or UO_335 (O_335,N_2896,N_2948);
or UO_336 (O_336,N_2989,N_2939);
nand UO_337 (O_337,N_2893,N_2809);
nor UO_338 (O_338,N_2855,N_2908);
nor UO_339 (O_339,N_2928,N_2903);
nor UO_340 (O_340,N_2929,N_2876);
or UO_341 (O_341,N_2877,N_2914);
nand UO_342 (O_342,N_2878,N_2983);
or UO_343 (O_343,N_2966,N_2804);
nor UO_344 (O_344,N_2838,N_2920);
nor UO_345 (O_345,N_2849,N_2802);
nand UO_346 (O_346,N_2827,N_2863);
and UO_347 (O_347,N_2900,N_2828);
xnor UO_348 (O_348,N_2966,N_2918);
nand UO_349 (O_349,N_2875,N_2989);
or UO_350 (O_350,N_2985,N_2837);
nand UO_351 (O_351,N_2829,N_2913);
nor UO_352 (O_352,N_2879,N_2882);
nand UO_353 (O_353,N_2906,N_2968);
nor UO_354 (O_354,N_2905,N_2887);
and UO_355 (O_355,N_2883,N_2838);
or UO_356 (O_356,N_2922,N_2813);
nand UO_357 (O_357,N_2831,N_2945);
nand UO_358 (O_358,N_2827,N_2867);
xnor UO_359 (O_359,N_2857,N_2901);
nor UO_360 (O_360,N_2898,N_2969);
nand UO_361 (O_361,N_2877,N_2905);
and UO_362 (O_362,N_2846,N_2932);
or UO_363 (O_363,N_2959,N_2882);
nand UO_364 (O_364,N_2997,N_2850);
or UO_365 (O_365,N_2868,N_2982);
or UO_366 (O_366,N_2803,N_2925);
nand UO_367 (O_367,N_2963,N_2897);
nor UO_368 (O_368,N_2801,N_2926);
nor UO_369 (O_369,N_2985,N_2953);
nand UO_370 (O_370,N_2828,N_2824);
nand UO_371 (O_371,N_2877,N_2816);
or UO_372 (O_372,N_2868,N_2948);
xnor UO_373 (O_373,N_2855,N_2910);
nand UO_374 (O_374,N_2931,N_2888);
and UO_375 (O_375,N_2849,N_2915);
nand UO_376 (O_376,N_2805,N_2833);
nor UO_377 (O_377,N_2954,N_2952);
and UO_378 (O_378,N_2880,N_2838);
and UO_379 (O_379,N_2859,N_2981);
and UO_380 (O_380,N_2940,N_2892);
nand UO_381 (O_381,N_2922,N_2843);
and UO_382 (O_382,N_2878,N_2992);
nand UO_383 (O_383,N_2869,N_2924);
and UO_384 (O_384,N_2865,N_2994);
and UO_385 (O_385,N_2862,N_2958);
or UO_386 (O_386,N_2849,N_2867);
or UO_387 (O_387,N_2841,N_2871);
nor UO_388 (O_388,N_2841,N_2915);
nand UO_389 (O_389,N_2871,N_2827);
nor UO_390 (O_390,N_2886,N_2920);
nor UO_391 (O_391,N_2816,N_2955);
nand UO_392 (O_392,N_2836,N_2875);
and UO_393 (O_393,N_2868,N_2900);
nor UO_394 (O_394,N_2833,N_2855);
or UO_395 (O_395,N_2808,N_2995);
nor UO_396 (O_396,N_2936,N_2895);
nor UO_397 (O_397,N_2905,N_2845);
nand UO_398 (O_398,N_2842,N_2918);
nand UO_399 (O_399,N_2996,N_2834);
nand UO_400 (O_400,N_2951,N_2994);
and UO_401 (O_401,N_2918,N_2906);
or UO_402 (O_402,N_2982,N_2919);
nor UO_403 (O_403,N_2937,N_2981);
nor UO_404 (O_404,N_2912,N_2981);
or UO_405 (O_405,N_2807,N_2874);
nor UO_406 (O_406,N_2863,N_2807);
or UO_407 (O_407,N_2875,N_2806);
nor UO_408 (O_408,N_2927,N_2907);
nand UO_409 (O_409,N_2955,N_2924);
xnor UO_410 (O_410,N_2998,N_2894);
nand UO_411 (O_411,N_2829,N_2848);
xor UO_412 (O_412,N_2869,N_2859);
nand UO_413 (O_413,N_2802,N_2946);
xor UO_414 (O_414,N_2930,N_2979);
nand UO_415 (O_415,N_2887,N_2980);
nor UO_416 (O_416,N_2908,N_2926);
and UO_417 (O_417,N_2903,N_2981);
and UO_418 (O_418,N_2928,N_2879);
or UO_419 (O_419,N_2909,N_2861);
nand UO_420 (O_420,N_2922,N_2915);
nor UO_421 (O_421,N_2954,N_2959);
nand UO_422 (O_422,N_2954,N_2830);
nor UO_423 (O_423,N_2809,N_2926);
xnor UO_424 (O_424,N_2873,N_2962);
xor UO_425 (O_425,N_2945,N_2819);
nand UO_426 (O_426,N_2910,N_2828);
nor UO_427 (O_427,N_2994,N_2852);
and UO_428 (O_428,N_2938,N_2961);
or UO_429 (O_429,N_2955,N_2882);
nor UO_430 (O_430,N_2910,N_2947);
or UO_431 (O_431,N_2945,N_2885);
nand UO_432 (O_432,N_2968,N_2911);
and UO_433 (O_433,N_2870,N_2949);
nand UO_434 (O_434,N_2826,N_2824);
and UO_435 (O_435,N_2916,N_2891);
and UO_436 (O_436,N_2819,N_2835);
nand UO_437 (O_437,N_2858,N_2868);
nand UO_438 (O_438,N_2810,N_2952);
and UO_439 (O_439,N_2869,N_2911);
xor UO_440 (O_440,N_2804,N_2816);
nor UO_441 (O_441,N_2860,N_2807);
nor UO_442 (O_442,N_2859,N_2925);
or UO_443 (O_443,N_2822,N_2963);
nand UO_444 (O_444,N_2837,N_2891);
nand UO_445 (O_445,N_2996,N_2840);
nand UO_446 (O_446,N_2978,N_2869);
xnor UO_447 (O_447,N_2870,N_2854);
or UO_448 (O_448,N_2898,N_2810);
or UO_449 (O_449,N_2990,N_2964);
nor UO_450 (O_450,N_2821,N_2973);
or UO_451 (O_451,N_2822,N_2964);
nor UO_452 (O_452,N_2882,N_2967);
or UO_453 (O_453,N_2951,N_2915);
nand UO_454 (O_454,N_2932,N_2863);
nor UO_455 (O_455,N_2942,N_2866);
and UO_456 (O_456,N_2941,N_2862);
nor UO_457 (O_457,N_2875,N_2951);
nand UO_458 (O_458,N_2833,N_2850);
or UO_459 (O_459,N_2935,N_2822);
nand UO_460 (O_460,N_2987,N_2826);
nor UO_461 (O_461,N_2914,N_2872);
or UO_462 (O_462,N_2980,N_2997);
and UO_463 (O_463,N_2807,N_2817);
nand UO_464 (O_464,N_2919,N_2904);
nor UO_465 (O_465,N_2886,N_2849);
or UO_466 (O_466,N_2892,N_2960);
nor UO_467 (O_467,N_2958,N_2951);
nand UO_468 (O_468,N_2930,N_2867);
nand UO_469 (O_469,N_2879,N_2899);
nand UO_470 (O_470,N_2899,N_2929);
or UO_471 (O_471,N_2882,N_2964);
nor UO_472 (O_472,N_2880,N_2921);
nor UO_473 (O_473,N_2893,N_2886);
nand UO_474 (O_474,N_2838,N_2925);
or UO_475 (O_475,N_2829,N_2926);
nor UO_476 (O_476,N_2823,N_2817);
nand UO_477 (O_477,N_2944,N_2865);
nor UO_478 (O_478,N_2826,N_2805);
nand UO_479 (O_479,N_2971,N_2983);
nor UO_480 (O_480,N_2869,N_2996);
nand UO_481 (O_481,N_2908,N_2824);
and UO_482 (O_482,N_2862,N_2810);
nor UO_483 (O_483,N_2848,N_2994);
and UO_484 (O_484,N_2964,N_2850);
nor UO_485 (O_485,N_2924,N_2968);
nand UO_486 (O_486,N_2947,N_2843);
and UO_487 (O_487,N_2935,N_2923);
nor UO_488 (O_488,N_2881,N_2908);
xnor UO_489 (O_489,N_2829,N_2915);
or UO_490 (O_490,N_2998,N_2852);
nor UO_491 (O_491,N_2894,N_2892);
or UO_492 (O_492,N_2921,N_2859);
and UO_493 (O_493,N_2934,N_2811);
nand UO_494 (O_494,N_2907,N_2911);
or UO_495 (O_495,N_2896,N_2868);
or UO_496 (O_496,N_2901,N_2937);
nor UO_497 (O_497,N_2954,N_2803);
or UO_498 (O_498,N_2935,N_2980);
or UO_499 (O_499,N_2862,N_2940);
endmodule