module basic_2500_25000_3000_20_levels_10xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_730,In_2093);
xnor U1 (N_1,In_1853,In_957);
nand U2 (N_2,In_838,In_2384);
nand U3 (N_3,In_2289,In_2269);
nand U4 (N_4,In_1497,In_293);
xor U5 (N_5,In_1982,In_791);
or U6 (N_6,In_2260,In_2121);
or U7 (N_7,In_1954,In_876);
or U8 (N_8,In_1513,In_1000);
and U9 (N_9,In_916,In_2191);
or U10 (N_10,In_1861,In_2494);
and U11 (N_11,In_1605,In_471);
nor U12 (N_12,In_1035,In_981);
xor U13 (N_13,In_1237,In_2087);
or U14 (N_14,In_1444,In_2450);
or U15 (N_15,In_1392,In_2466);
nor U16 (N_16,In_2412,In_105);
or U17 (N_17,In_1449,In_625);
or U18 (N_18,In_1330,In_1366);
xor U19 (N_19,In_1758,In_449);
xnor U20 (N_20,In_1396,In_1290);
and U21 (N_21,In_929,In_1895);
nand U22 (N_22,In_2428,In_1915);
nand U23 (N_23,In_6,In_15);
nand U24 (N_24,In_1477,In_773);
nand U25 (N_25,In_2148,In_2411);
nor U26 (N_26,In_588,In_1595);
nand U27 (N_27,In_1092,In_85);
nand U28 (N_28,In_968,In_1529);
nor U29 (N_29,In_1022,In_1610);
or U30 (N_30,In_1430,In_198);
nor U31 (N_31,In_1293,In_1421);
nand U32 (N_32,In_1768,In_1696);
xnor U33 (N_33,In_217,In_1206);
nand U34 (N_34,In_819,In_2048);
or U35 (N_35,In_1798,In_937);
nor U36 (N_36,In_828,In_2446);
or U37 (N_37,In_2056,In_1681);
nand U38 (N_38,In_2137,In_1727);
and U39 (N_39,In_1008,In_1918);
and U40 (N_40,In_794,In_1439);
or U41 (N_41,In_1787,In_770);
or U42 (N_42,In_1139,In_1380);
and U43 (N_43,In_716,In_1753);
xnor U44 (N_44,In_966,In_2439);
xnor U45 (N_45,In_970,In_1182);
nand U46 (N_46,In_1624,In_2051);
or U47 (N_47,In_2493,In_1950);
nand U48 (N_48,In_1199,In_721);
nand U49 (N_49,In_2266,In_501);
and U50 (N_50,In_2157,In_1908);
nand U51 (N_51,In_1188,In_2117);
xnor U52 (N_52,In_2455,In_1849);
and U53 (N_53,In_855,In_567);
and U54 (N_54,In_2331,In_2171);
or U55 (N_55,In_2255,In_2066);
nand U56 (N_56,In_1257,In_607);
xor U57 (N_57,In_1809,In_1086);
xnor U58 (N_58,In_1080,In_2488);
and U59 (N_59,In_1005,In_1431);
nor U60 (N_60,In_1572,In_591);
or U61 (N_61,In_1967,In_232);
nand U62 (N_62,In_175,In_1976);
xnor U63 (N_63,In_856,In_379);
nand U64 (N_64,In_2133,In_87);
nand U65 (N_65,In_1118,In_881);
or U66 (N_66,In_1952,In_1598);
or U67 (N_67,In_547,In_1304);
nor U68 (N_68,In_1576,In_1678);
xnor U69 (N_69,In_557,In_531);
nand U70 (N_70,In_1314,In_1644);
and U71 (N_71,In_247,In_639);
and U72 (N_72,In_2333,In_2403);
and U73 (N_73,In_1709,In_2473);
xnor U74 (N_74,In_0,In_1898);
or U75 (N_75,In_216,In_662);
and U76 (N_76,In_1484,In_1170);
nor U77 (N_77,In_1990,In_789);
and U78 (N_78,In_901,In_1723);
nand U79 (N_79,In_1207,In_2225);
or U80 (N_80,In_2363,In_1432);
nor U81 (N_81,In_2106,In_1362);
nand U82 (N_82,In_1567,In_315);
or U83 (N_83,In_713,In_1202);
or U84 (N_84,In_1817,In_1822);
nor U85 (N_85,In_2352,In_1784);
and U86 (N_86,In_324,In_1883);
nor U87 (N_87,In_294,In_7);
nor U88 (N_88,In_2485,In_1475);
xnor U89 (N_89,In_1355,In_892);
xor U90 (N_90,In_1397,In_173);
or U91 (N_91,In_400,In_1470);
and U92 (N_92,In_1042,In_960);
nand U93 (N_93,In_366,In_2313);
or U94 (N_94,In_709,In_1201);
or U95 (N_95,In_1391,In_825);
nor U96 (N_96,In_934,In_1276);
and U97 (N_97,In_243,In_803);
and U98 (N_98,In_367,In_1427);
nand U99 (N_99,In_1923,In_509);
or U100 (N_100,In_130,In_440);
xor U101 (N_101,In_1872,In_2110);
nand U102 (N_102,In_207,In_1090);
xnor U103 (N_103,In_2379,In_1532);
nand U104 (N_104,In_1603,In_2149);
nor U105 (N_105,In_1402,In_729);
xor U106 (N_106,In_463,In_1119);
xnor U107 (N_107,In_1543,In_86);
nor U108 (N_108,In_1596,In_2174);
or U109 (N_109,In_2319,In_536);
or U110 (N_110,In_484,In_561);
nor U111 (N_111,In_1937,In_678);
or U112 (N_112,In_1072,In_1867);
or U113 (N_113,In_555,In_944);
and U114 (N_114,In_907,In_654);
or U115 (N_115,In_1669,In_1810);
nor U116 (N_116,In_632,In_550);
nand U117 (N_117,In_717,In_138);
or U118 (N_118,In_2396,In_1030);
nand U119 (N_119,In_1450,In_1050);
and U120 (N_120,In_1300,In_2180);
nor U121 (N_121,In_2091,In_80);
or U122 (N_122,In_745,In_433);
nand U123 (N_123,In_1458,In_818);
nor U124 (N_124,In_487,In_287);
or U125 (N_125,In_1780,In_1085);
xor U126 (N_126,In_1194,In_759);
and U127 (N_127,In_749,In_1983);
nor U128 (N_128,In_1217,In_1562);
nor U129 (N_129,In_571,In_1944);
and U130 (N_130,In_1189,In_801);
nand U131 (N_131,In_784,In_2131);
nor U132 (N_132,In_1597,In_1679);
and U133 (N_133,In_1184,In_1826);
and U134 (N_134,In_734,In_1220);
xnor U135 (N_135,In_1551,In_768);
nand U136 (N_136,In_686,In_1100);
nand U137 (N_137,In_375,In_347);
nand U138 (N_138,In_940,In_1730);
or U139 (N_139,In_1645,In_1510);
xor U140 (N_140,In_2176,In_635);
nand U141 (N_141,In_354,In_1641);
xnor U142 (N_142,In_520,In_167);
xnor U143 (N_143,In_21,In_486);
nand U144 (N_144,In_2172,In_1691);
or U145 (N_145,In_1663,In_1344);
nor U146 (N_146,In_2429,In_905);
nand U147 (N_147,In_1233,In_1801);
nand U148 (N_148,In_787,In_200);
nand U149 (N_149,In_2454,In_2476);
or U150 (N_150,In_586,In_1120);
xor U151 (N_151,In_1420,In_58);
xor U152 (N_152,In_2491,In_2308);
and U153 (N_153,In_492,In_1246);
nor U154 (N_154,In_1660,In_1466);
xnor U155 (N_155,In_1770,In_1575);
and U156 (N_156,In_290,In_135);
xor U157 (N_157,In_1271,In_1451);
xnor U158 (N_158,In_2130,In_187);
nand U159 (N_159,In_1554,In_843);
nand U160 (N_160,In_2211,In_1882);
or U161 (N_161,In_2477,In_2281);
xor U162 (N_162,In_1150,In_2273);
nor U163 (N_163,In_785,In_1897);
and U164 (N_164,In_2479,In_1360);
nor U165 (N_165,In_141,In_128);
and U166 (N_166,In_1888,In_2055);
nor U167 (N_167,In_147,In_1067);
nor U168 (N_168,In_754,In_2298);
or U169 (N_169,In_2402,In_1253);
xnor U170 (N_170,In_2060,In_1694);
or U171 (N_171,In_932,In_1185);
and U172 (N_172,In_209,In_574);
nor U173 (N_173,In_1821,In_316);
nor U174 (N_174,In_652,In_2392);
or U175 (N_175,In_936,In_777);
xnor U176 (N_176,In_2008,In_958);
nand U177 (N_177,In_609,In_797);
or U178 (N_178,In_620,In_190);
xnor U179 (N_179,In_36,In_2230);
xnor U180 (N_180,In_2036,In_1692);
xnor U181 (N_181,In_942,In_597);
nand U182 (N_182,In_437,In_2290);
and U183 (N_183,In_1557,In_1178);
nand U184 (N_184,In_2090,In_655);
and U185 (N_185,In_1126,In_1365);
nand U186 (N_186,In_644,In_813);
and U187 (N_187,In_2199,In_2219);
xor U188 (N_188,In_2160,In_2336);
xor U189 (N_189,In_1547,In_604);
xnor U190 (N_190,In_599,In_1373);
nand U191 (N_191,In_2178,In_1445);
nor U192 (N_192,In_1070,In_42);
xnor U193 (N_193,In_2229,In_687);
nor U194 (N_194,In_672,In_1242);
xnor U195 (N_195,In_1634,In_1773);
or U196 (N_196,In_1713,In_723);
nand U197 (N_197,In_2404,In_1388);
nor U198 (N_198,In_1592,In_1599);
xor U199 (N_199,In_1416,In_2286);
nand U200 (N_200,In_535,In_2399);
xor U201 (N_201,In_2052,In_1863);
and U202 (N_202,In_1236,In_364);
and U203 (N_203,In_236,In_240);
nor U204 (N_204,In_1881,In_1827);
nor U205 (N_205,In_1788,In_1198);
nand U206 (N_206,In_62,In_757);
nand U207 (N_207,In_1407,In_827);
nand U208 (N_208,In_1132,In_746);
and U209 (N_209,In_707,In_2315);
or U210 (N_210,In_2419,In_904);
or U211 (N_211,In_30,In_808);
and U212 (N_212,In_1460,In_714);
and U213 (N_213,In_1374,In_1176);
nand U214 (N_214,In_1536,In_1270);
nor U215 (N_215,In_852,In_1633);
nor U216 (N_216,In_2226,In_155);
and U217 (N_217,In_2467,In_933);
and U218 (N_218,In_642,In_1196);
or U219 (N_219,In_1351,In_181);
nand U220 (N_220,In_1635,In_2294);
and U221 (N_221,In_342,In_946);
nor U222 (N_222,In_728,In_1101);
and U223 (N_223,In_2039,In_579);
nor U224 (N_224,In_1677,In_1117);
or U225 (N_225,In_1762,In_922);
xor U226 (N_226,In_1284,In_1103);
or U227 (N_227,In_1992,In_398);
nand U228 (N_228,In_1910,In_472);
or U229 (N_229,In_1089,In_2353);
or U230 (N_230,In_523,In_1155);
nand U231 (N_231,In_2385,In_204);
or U232 (N_232,In_2293,In_2258);
nor U233 (N_233,In_602,In_570);
nor U234 (N_234,In_1951,In_441);
or U235 (N_235,In_792,In_1682);
nor U236 (N_236,In_1511,In_959);
nand U237 (N_237,In_751,In_1856);
and U238 (N_238,In_1651,In_705);
nor U239 (N_239,In_956,In_1964);
and U240 (N_240,In_1507,In_1676);
or U241 (N_241,In_168,In_1854);
xnor U242 (N_242,In_1088,In_624);
and U243 (N_243,In_1157,In_118);
nand U244 (N_244,In_451,In_386);
xnor U245 (N_245,In_1746,In_2156);
xor U246 (N_246,In_582,In_2200);
and U247 (N_247,In_513,In_2212);
xnor U248 (N_248,In_887,In_798);
xnor U249 (N_249,In_1945,In_993);
nor U250 (N_250,In_1811,In_1429);
nand U251 (N_251,In_637,In_1131);
or U252 (N_252,In_421,In_1862);
or U253 (N_253,In_246,In_2128);
or U254 (N_254,In_1984,In_2074);
or U255 (N_255,In_1068,In_1311);
xor U256 (N_256,In_1286,In_51);
xor U257 (N_257,In_826,In_1903);
and U258 (N_258,In_1925,In_1779);
and U259 (N_259,In_1212,In_1516);
nand U260 (N_260,In_563,In_1037);
xnor U261 (N_261,In_722,In_185);
or U262 (N_262,In_2135,In_20);
nand U263 (N_263,In_1569,In_1098);
and U264 (N_264,In_1024,In_430);
xor U265 (N_265,In_2193,In_823);
and U266 (N_266,In_2481,In_2153);
or U267 (N_267,In_2065,In_1180);
xor U268 (N_268,In_2442,In_419);
and U269 (N_269,In_930,In_1369);
nand U270 (N_270,In_410,In_2018);
or U271 (N_271,In_339,In_23);
or U272 (N_272,In_2387,In_2007);
nor U273 (N_273,In_762,In_776);
nor U274 (N_274,In_132,In_2390);
or U275 (N_275,In_837,In_2031);
and U276 (N_276,In_1818,In_996);
or U277 (N_277,In_1031,In_1969);
xnor U278 (N_278,In_387,In_1277);
or U279 (N_279,In_683,In_47);
nand U280 (N_280,In_2283,In_2115);
xnor U281 (N_281,In_1805,In_595);
or U282 (N_282,In_2468,In_158);
or U283 (N_283,In_2068,In_1076);
or U284 (N_284,In_322,In_1461);
xor U285 (N_285,In_2146,In_2367);
and U286 (N_286,In_445,In_68);
nor U287 (N_287,In_202,In_2046);
nor U288 (N_288,In_1525,In_605);
and U289 (N_289,In_1454,In_61);
nor U290 (N_290,In_1312,In_159);
or U291 (N_291,In_1970,In_517);
nor U292 (N_292,In_1041,In_507);
nor U293 (N_293,In_2227,In_1517);
or U294 (N_294,In_12,In_1154);
or U295 (N_295,In_2444,In_1652);
xnor U296 (N_296,In_634,In_910);
nor U297 (N_297,In_2332,In_1193);
xor U298 (N_298,In_1671,In_1130);
xnor U299 (N_299,In_1621,In_438);
and U300 (N_300,In_2034,In_606);
xnor U301 (N_301,In_274,In_2001);
nor U302 (N_302,In_184,In_2010);
nor U303 (N_303,In_286,In_1791);
and U304 (N_304,In_1548,In_1695);
xor U305 (N_305,In_203,In_214);
and U306 (N_306,In_2122,In_182);
or U307 (N_307,In_1763,In_1754);
or U308 (N_308,In_1528,In_1716);
and U309 (N_309,In_1036,In_1542);
xnor U310 (N_310,In_598,In_296);
nor U311 (N_311,In_2158,In_779);
and U312 (N_312,In_650,In_1625);
xor U313 (N_313,In_911,In_1859);
or U314 (N_314,In_2424,In_2089);
or U315 (N_315,In_2220,In_1447);
nand U316 (N_316,In_412,In_2070);
or U317 (N_317,In_1640,In_564);
nor U318 (N_318,In_1729,In_2295);
nor U319 (N_319,In_2312,In_428);
or U320 (N_320,In_753,In_1462);
and U321 (N_321,In_2096,In_1422);
nand U322 (N_322,In_477,In_1636);
or U323 (N_323,In_763,In_1838);
or U324 (N_324,In_2116,In_1559);
and U325 (N_325,In_1264,In_804);
xnor U326 (N_326,In_2397,In_1174);
and U327 (N_327,In_1029,In_636);
or U328 (N_328,In_651,In_1852);
and U329 (N_329,In_962,In_473);
and U330 (N_330,In_991,In_300);
xor U331 (N_331,In_197,In_332);
or U332 (N_332,In_2100,In_373);
nor U333 (N_333,In_450,In_2103);
nor U334 (N_334,In_2271,In_551);
nor U335 (N_335,In_45,In_1408);
nor U336 (N_336,In_1111,In_1699);
nor U337 (N_337,In_120,In_1585);
nor U338 (N_338,In_392,In_875);
and U339 (N_339,In_1282,In_186);
nor U340 (N_340,In_1973,In_378);
xor U341 (N_341,In_583,In_82);
nor U342 (N_342,In_309,In_1382);
and U343 (N_343,In_1858,In_374);
xor U344 (N_344,In_1222,In_2002);
nor U345 (N_345,In_1501,In_1235);
or U346 (N_346,In_2022,In_1261);
or U347 (N_347,In_1329,In_2420);
or U348 (N_348,In_1425,In_589);
nor U349 (N_349,In_1323,In_2162);
nand U350 (N_350,In_1506,In_1229);
xor U351 (N_351,In_1994,In_1007);
nor U352 (N_352,In_920,In_245);
nand U353 (N_353,In_1978,In_1260);
and U354 (N_354,In_1527,In_385);
xor U355 (N_355,In_769,In_2321);
xor U356 (N_356,In_1776,In_201);
or U357 (N_357,In_1252,In_525);
xor U358 (N_358,In_171,In_1307);
nor U359 (N_359,In_326,In_593);
or U360 (N_360,In_1766,In_2080);
nand U361 (N_361,In_1590,In_967);
xnor U362 (N_362,In_357,In_772);
nor U363 (N_363,In_2040,In_1321);
and U364 (N_364,In_1411,In_1363);
nand U365 (N_365,In_2460,In_1110);
nor U366 (N_366,In_2086,In_2195);
and U367 (N_367,In_861,In_1656);
nand U368 (N_368,In_212,In_465);
and U369 (N_369,In_2084,In_1785);
nand U370 (N_370,In_9,In_299);
xor U371 (N_371,In_2126,In_2235);
xor U372 (N_372,In_1115,In_1144);
xor U373 (N_373,In_2447,In_2217);
and U374 (N_374,In_809,In_455);
xnor U375 (N_375,In_796,In_1463);
xnor U376 (N_376,In_680,In_1933);
nand U377 (N_377,In_663,In_1412);
nor U378 (N_378,In_850,In_1885);
xor U379 (N_379,In_1835,In_900);
nand U380 (N_380,In_2144,In_2453);
or U381 (N_381,In_912,In_310);
nand U382 (N_382,In_727,In_1141);
and U383 (N_383,In_1414,In_848);
nor U384 (N_384,In_1690,In_1325);
nor U385 (N_385,In_1761,In_1571);
xor U386 (N_386,In_14,In_1441);
nand U387 (N_387,In_562,In_2486);
xor U388 (N_388,In_1755,In_983);
or U389 (N_389,In_580,In_718);
xnor U390 (N_390,In_931,In_1152);
xor U391 (N_391,In_1712,In_1249);
or U392 (N_392,In_2240,In_1775);
xnor U393 (N_393,In_976,In_1191);
and U394 (N_394,In_495,In_546);
nand U395 (N_395,In_1424,In_2362);
or U396 (N_396,In_1192,In_1357);
nor U397 (N_397,In_1802,In_1032);
or U398 (N_398,In_2045,In_1148);
nand U399 (N_399,In_2306,In_867);
nor U400 (N_400,In_1341,In_1015);
xnor U401 (N_401,In_407,In_516);
xnor U402 (N_402,In_735,In_1409);
nor U403 (N_403,In_882,In_1689);
and U404 (N_404,In_880,In_1931);
or U405 (N_405,In_1108,In_1726);
and U406 (N_406,In_1541,In_1069);
nor U407 (N_407,In_2350,In_362);
nand U408 (N_408,In_205,In_331);
nand U409 (N_409,In_223,In_382);
xor U410 (N_410,In_1719,In_1018);
nand U411 (N_411,In_2497,In_1717);
nor U412 (N_412,In_953,In_2143);
nor U413 (N_413,In_950,In_681);
and U414 (N_414,In_90,In_2241);
xor U415 (N_415,In_2296,In_1778);
and U416 (N_416,In_60,In_2337);
and U417 (N_417,In_165,In_2139);
and U418 (N_418,In_1891,In_2369);
nand U419 (N_419,In_1673,In_1869);
or U420 (N_420,In_1946,In_1836);
nor U421 (N_421,In_16,In_712);
or U422 (N_422,In_1204,In_2138);
and U423 (N_423,In_774,In_519);
xor U424 (N_424,In_1019,In_1655);
nand U425 (N_425,In_1349,In_208);
nand U426 (N_426,In_1570,In_581);
nor U427 (N_427,In_914,In_657);
nor U428 (N_428,In_998,In_1887);
and U429 (N_429,In_619,In_824);
nor U430 (N_430,In_35,In_270);
xnor U431 (N_431,In_786,In_388);
xnor U432 (N_432,In_2417,In_1377);
or U433 (N_433,In_2147,In_54);
and U434 (N_434,In_391,In_2343);
xnor U435 (N_435,In_2111,In_1837);
nand U436 (N_436,In_1494,In_1828);
nor U437 (N_437,In_1829,In_732);
or U438 (N_438,In_1917,In_2216);
and U439 (N_439,In_1668,In_849);
xor U440 (N_440,In_24,In_847);
xnor U441 (N_441,In_1664,In_1467);
and U442 (N_442,In_886,In_2047);
and U443 (N_443,In_1880,In_1186);
nor U444 (N_444,In_1295,In_269);
and U445 (N_445,In_1254,In_2408);
nor U446 (N_446,In_1612,In_417);
nor U447 (N_447,In_73,In_1114);
or U448 (N_448,In_1748,In_1423);
nor U449 (N_449,In_1803,In_696);
or U450 (N_450,In_2004,In_2329);
nand U451 (N_451,In_1471,In_1386);
nor U452 (N_452,In_1745,In_2097);
xor U453 (N_453,In_67,In_2270);
nor U454 (N_454,In_615,In_514);
and U455 (N_455,In_954,In_1608);
or U456 (N_456,In_671,In_1760);
nor U457 (N_457,In_1884,In_2472);
xnor U458 (N_458,In_2243,In_1159);
and U459 (N_459,In_646,In_1986);
and U460 (N_460,In_1629,In_1740);
or U461 (N_461,In_1279,In_1767);
nand U462 (N_462,In_2347,In_2341);
or U463 (N_463,In_475,In_56);
or U464 (N_464,In_1701,In_2000);
nor U465 (N_465,In_2301,In_96);
nand U466 (N_466,In_2053,In_2185);
and U467 (N_467,In_949,In_853);
nand U468 (N_468,In_1303,In_1020);
nand U469 (N_469,In_690,In_2268);
or U470 (N_470,In_2380,In_502);
xnor U471 (N_471,In_89,In_2026);
nor U472 (N_472,In_1026,In_2335);
or U473 (N_473,In_1924,In_592);
nor U474 (N_474,In_1398,In_276);
nand U475 (N_475,In_1057,In_1419);
or U476 (N_476,In_1231,In_975);
and U477 (N_477,In_418,In_2025);
nor U478 (N_478,In_129,In_1685);
and U479 (N_479,In_2181,In_1346);
and U480 (N_480,In_104,In_1613);
and U481 (N_481,In_1298,In_255);
nor U482 (N_482,In_453,In_233);
xor U483 (N_483,In_578,In_832);
nand U484 (N_484,In_2448,In_1647);
or U485 (N_485,In_1082,In_272);
nor U486 (N_486,In_1919,In_1104);
nor U487 (N_487,In_126,In_1857);
nor U488 (N_488,In_1485,In_2482);
xor U489 (N_489,In_2431,In_542);
xnor U490 (N_490,In_37,In_1345);
and U491 (N_491,In_1340,In_2035);
or U492 (N_492,In_1975,In_1792);
nor U493 (N_493,In_1255,In_273);
nor U494 (N_494,In_1371,In_429);
and U495 (N_495,In_335,In_231);
and U496 (N_496,In_1631,In_151);
and U497 (N_497,In_267,In_2305);
nor U498 (N_498,In_2125,In_1581);
nand U499 (N_499,In_2438,In_1142);
nor U500 (N_500,In_1081,In_2006);
and U501 (N_501,In_280,In_610);
and U502 (N_502,In_896,In_2372);
xnor U503 (N_503,In_2334,In_764);
xor U504 (N_504,In_432,In_333);
or U505 (N_505,In_1797,In_1375);
nor U506 (N_506,In_1733,In_125);
and U507 (N_507,In_1239,In_658);
nand U508 (N_508,In_2490,In_1574);
or U509 (N_509,In_1800,In_1988);
nand U510 (N_510,In_482,In_2407);
xnor U511 (N_511,In_462,In_491);
xor U512 (N_512,In_793,In_2364);
xor U513 (N_513,In_76,In_1698);
and U514 (N_514,In_1045,In_1269);
nor U515 (N_515,In_1601,In_1209);
and U516 (N_516,In_219,In_1436);
nor U517 (N_517,In_2359,In_2284);
nand U518 (N_518,In_2127,In_113);
nor U519 (N_519,In_1509,In_2015);
xnor U520 (N_520,In_2071,In_1028);
nand U521 (N_521,In_164,In_2057);
nand U522 (N_522,In_1560,In_1285);
or U523 (N_523,In_1568,In_46);
xor U524 (N_524,In_1615,In_980);
or U525 (N_525,In_2291,In_854);
xor U526 (N_526,In_1400,In_2414);
nand U527 (N_527,In_1468,In_524);
nand U528 (N_528,In_1661,In_1224);
and U529 (N_529,In_2175,In_2023);
xnor U530 (N_530,In_1166,In_835);
xnor U531 (N_531,In_1245,In_2250);
nand U532 (N_532,In_122,In_211);
and U533 (N_533,In_2215,In_2099);
and U534 (N_534,In_747,In_2064);
and U535 (N_535,In_1384,In_2461);
and U536 (N_536,In_92,In_528);
or U537 (N_537,In_2457,In_1934);
nor U538 (N_538,In_404,In_238);
nand U539 (N_539,In_750,In_1834);
nand U540 (N_540,In_1850,In_601);
and U541 (N_541,In_2483,In_448);
or U542 (N_542,In_1228,In_1524);
xor U543 (N_543,In_1124,In_552);
nand U544 (N_544,In_995,In_341);
and U545 (N_545,In_1846,In_2277);
or U546 (N_546,In_183,In_1313);
or U547 (N_547,In_1515,In_2118);
nand U548 (N_548,In_788,In_1823);
nor U549 (N_549,In_565,In_1839);
nand U550 (N_550,In_613,In_169);
or U551 (N_551,In_2078,In_1957);
xnor U552 (N_552,In_2024,In_1387);
nand U553 (N_553,In_1530,In_1979);
and U554 (N_554,In_2032,In_1021);
or U555 (N_555,In_1134,In_1364);
nor U556 (N_556,In_2261,In_1038);
or U557 (N_557,In_1324,In_939);
nor U558 (N_558,In_1247,In_1265);
nor U559 (N_559,In_358,In_695);
nand U560 (N_560,In_1749,In_131);
xor U561 (N_561,In_268,In_1216);
or U562 (N_562,In_971,In_150);
nor U563 (N_563,In_2173,In_494);
xor U564 (N_564,In_668,In_1278);
xnor U565 (N_565,In_1614,In_845);
nand U566 (N_566,In_873,In_585);
nor U567 (N_567,In_2348,In_2119);
and U568 (N_568,In_41,In_526);
or U569 (N_569,In_2083,In_623);
or U570 (N_570,In_1503,In_74);
or U571 (N_571,In_806,In_196);
nand U572 (N_572,In_2108,In_925);
and U573 (N_573,In_178,In_2037);
and U574 (N_574,In_291,In_1338);
and U575 (N_575,In_1706,In_2027);
or U576 (N_576,In_1127,In_549);
xor U577 (N_577,In_1700,In_569);
or U578 (N_578,In_2206,In_1949);
or U579 (N_579,In_2205,In_1112);
or U580 (N_580,In_726,In_1972);
or U581 (N_581,In_402,In_1627);
nor U582 (N_582,In_1288,In_234);
nor U583 (N_583,In_1906,In_195);
nand U584 (N_584,In_145,In_742);
xnor U585 (N_585,In_371,In_281);
nand U586 (N_586,In_1459,In_1280);
nand U587 (N_587,In_1743,In_1626);
or U588 (N_588,In_174,In_612);
nand U589 (N_589,In_1123,In_2484);
or U590 (N_590,In_1381,In_1116);
nand U591 (N_591,In_1980,In_365);
and U592 (N_592,In_822,In_1167);
nand U593 (N_593,In_1405,In_679);
and U594 (N_594,In_2395,In_1133);
and U595 (N_595,In_2487,In_1063);
and U596 (N_596,In_2265,In_2280);
nand U597 (N_597,In_2011,In_1750);
nor U598 (N_598,In_458,In_1410);
xnor U599 (N_599,In_1563,In_684);
or U600 (N_600,In_1358,In_1318);
xor U601 (N_601,In_2340,In_1993);
and U602 (N_602,In_1208,In_1059);
and U603 (N_603,In_199,In_1145);
xnor U604 (N_604,In_989,In_1913);
nand U605 (N_605,In_737,In_1870);
or U606 (N_606,In_1866,In_1966);
and U607 (N_607,In_1947,In_2038);
or U608 (N_608,In_1244,In_1879);
nor U609 (N_609,In_1060,In_1079);
and U610 (N_610,In_1496,In_479);
or U611 (N_611,In_1697,In_102);
nand U612 (N_612,In_834,In_1877);
xor U613 (N_613,In_2236,In_1637);
and U614 (N_614,In_220,In_1606);
or U615 (N_615,In_2423,In_81);
and U616 (N_616,In_1806,In_31);
nor U617 (N_617,In_1956,In_1440);
xnor U618 (N_618,In_2349,In_1310);
and U619 (N_619,In_1508,In_222);
xnor U620 (N_620,In_65,In_1047);
and U621 (N_621,In_554,In_1437);
nand U622 (N_622,In_698,In_88);
xnor U623 (N_623,In_629,In_1138);
xnor U624 (N_624,In_461,In_2425);
nand U625 (N_625,In_748,In_256);
nand U626 (N_626,In_188,In_1922);
nand U627 (N_627,In_1686,In_846);
and U628 (N_628,In_2107,In_504);
nor U629 (N_629,In_1916,In_2492);
or U630 (N_630,In_643,In_693);
or U631 (N_631,In_1587,In_406);
nand U632 (N_632,In_1737,In_1958);
nor U633 (N_633,In_530,In_377);
xnor U634 (N_634,In_1830,In_144);
nor U635 (N_635,In_1544,In_1428);
nand U636 (N_636,In_2297,In_577);
and U637 (N_637,In_1981,In_1799);
nand U638 (N_638,In_2207,In_2426);
or U639 (N_639,In_2409,In_33);
xor U640 (N_640,In_2415,In_2279);
and U641 (N_641,In_1832,In_289);
or U642 (N_642,In_1315,In_978);
nand U643 (N_643,In_1275,In_1306);
nand U644 (N_644,In_2237,In_948);
nor U645 (N_645,In_1687,In_1495);
or U646 (N_646,In_997,In_221);
xnor U647 (N_647,In_638,In_1354);
and U648 (N_648,In_2094,In_2360);
and U649 (N_649,In_327,In_1378);
or U650 (N_650,In_363,In_1638);
nor U651 (N_651,In_2288,In_771);
and U652 (N_652,In_124,In_192);
xor U653 (N_653,In_489,In_943);
and U654 (N_654,In_2330,In_98);
nor U655 (N_655,In_301,In_308);
nor U656 (N_656,In_2105,In_1256);
xnor U657 (N_657,In_2318,In_1890);
nand U658 (N_658,In_1062,In_1456);
nand U659 (N_659,In_1406,In_194);
xnor U660 (N_660,In_2368,In_2194);
and U661 (N_661,In_618,In_1793);
or U662 (N_662,In_2475,In_878);
nand U663 (N_663,In_1181,In_2401);
and U664 (N_664,In_384,In_1789);
or U665 (N_665,In_1164,In_1049);
or U666 (N_666,In_870,In_866);
xnor U667 (N_667,In_1998,In_1017);
xnor U668 (N_668,In_1911,In_2310);
xnor U669 (N_669,In_235,In_2463);
nand U670 (N_670,In_1172,In_1291);
nand U671 (N_671,In_1896,In_2164);
or U672 (N_672,In_2264,In_2054);
or U673 (N_673,In_558,In_1955);
nand U674 (N_674,In_1971,In_84);
nand U675 (N_675,In_1977,In_1550);
or U676 (N_676,In_1938,In_162);
xor U677 (N_677,In_110,In_839);
and U678 (N_678,In_1808,In_394);
or U679 (N_679,In_1302,In_2304);
or U680 (N_680,In_2079,In_1845);
xnor U681 (N_681,In_2151,In_1125);
nor U682 (N_682,In_2406,In_669);
and U683 (N_683,In_2017,In_545);
or U684 (N_684,In_543,In_736);
nor U685 (N_685,In_2292,In_1960);
xnor U686 (N_686,In_1273,In_1289);
xnor U687 (N_687,In_1039,In_1443);
xor U688 (N_688,In_863,In_1985);
or U689 (N_689,In_2209,In_189);
xor U690 (N_690,In_2221,In_1140);
and U691 (N_691,In_778,In_468);
or U692 (N_692,In_1301,In_2242);
or U693 (N_693,In_1577,In_1874);
xor U694 (N_694,In_2400,In_2248);
xnor U695 (N_695,In_18,In_1526);
nor U696 (N_696,In_2275,In_1162);
nor U697 (N_697,In_2030,In_918);
xor U698 (N_698,In_2136,In_2092);
nand U699 (N_699,In_1073,In_1361);
and U700 (N_700,In_1452,In_1113);
xnor U701 (N_701,In_1643,In_2338);
or U702 (N_702,In_1091,In_1618);
nor U703 (N_703,In_161,In_1522);
or U704 (N_704,In_576,In_2109);
xnor U705 (N_705,In_1537,In_1317);
xnor U706 (N_706,In_1632,In_346);
nor U707 (N_707,In_1099,In_676);
xor U708 (N_708,In_1646,In_399);
nand U709 (N_709,In_1183,In_323);
nor U710 (N_710,In_1095,In_2365);
xor U711 (N_711,In_908,In_1751);
xnor U712 (N_712,In_836,In_2421);
xor U713 (N_713,In_2282,In_821);
and U714 (N_714,In_372,In_1804);
or U715 (N_715,In_1305,In_1446);
or U716 (N_716,In_869,In_1053);
nand U717 (N_717,In_359,In_1339);
nand U718 (N_718,In_2196,In_416);
or U719 (N_719,In_1210,In_1197);
or U720 (N_720,In_2062,In_2389);
or U721 (N_721,In_237,In_1078);
and U722 (N_722,In_2398,In_600);
xnor U723 (N_723,In_2358,In_446);
nand U724 (N_724,In_2,In_395);
and U725 (N_725,In_1335,In_389);
and U726 (N_726,In_889,In_2069);
xor U727 (N_727,In_938,In_560);
or U728 (N_728,In_2309,In_2316);
nand U729 (N_729,In_2182,In_1771);
nand U730 (N_730,In_1096,In_532);
or U731 (N_731,In_1014,In_295);
nor U732 (N_732,In_1813,In_1490);
nand U733 (N_733,In_2311,In_1653);
or U734 (N_734,In_329,In_622);
nand U735 (N_735,In_1061,In_1493);
and U736 (N_736,In_263,In_2391);
or U737 (N_737,In_807,In_1489);
xor U738 (N_738,In_1012,In_405);
or U739 (N_739,In_2187,In_411);
nand U740 (N_740,In_2123,In_1223);
xnor U741 (N_741,In_1795,In_1948);
xnor U742 (N_742,In_1520,In_587);
or U743 (N_743,In_206,In_1703);
and U744 (N_744,In_1179,In_229);
or U745 (N_745,In_631,In_874);
or U746 (N_746,In_328,In_820);
xnor U747 (N_747,In_1600,In_704);
xnor U748 (N_748,In_1153,In_1147);
or U749 (N_749,In_109,In_1442);
or U750 (N_750,In_390,In_459);
xor U751 (N_751,In_2183,In_177);
or U752 (N_752,In_1894,In_1267);
nand U753 (N_753,In_1649,In_575);
nand U754 (N_754,In_1940,In_888);
xor U755 (N_755,In_248,In_302);
or U756 (N_756,In_1630,In_1693);
nor U757 (N_757,In_176,In_193);
nor U758 (N_758,In_1001,In_2072);
or U759 (N_759,In_343,In_1054);
and U760 (N_760,In_2378,In_1772);
nor U761 (N_761,In_337,In_1077);
or U762 (N_762,In_408,In_2287);
and U763 (N_763,In_2049,In_464);
and U764 (N_764,In_691,In_952);
or U765 (N_765,In_2272,In_2188);
or U766 (N_766,In_511,In_752);
xnor U767 (N_767,In_1607,In_1292);
xnor U768 (N_768,In_817,In_2161);
nand U769 (N_769,In_945,In_114);
nand U770 (N_770,In_701,In_706);
nor U771 (N_771,In_2014,In_760);
or U772 (N_772,In_1052,In_1909);
nor U773 (N_773,In_720,In_883);
nand U774 (N_774,In_2393,In_1002);
nand U775 (N_775,In_877,In_2177);
and U776 (N_776,In_303,In_2198);
xnor U777 (N_777,In_1642,In_924);
xor U778 (N_778,In_739,In_1831);
or U779 (N_779,In_34,In_2451);
nor U780 (N_780,In_52,In_257);
nor U781 (N_781,In_1502,In_844);
or U782 (N_782,In_1383,In_627);
nand U783 (N_783,In_1921,In_556);
xor U784 (N_784,In_149,In_2422);
nor U785 (N_785,In_1221,In_1759);
and U786 (N_786,In_1287,In_478);
or U787 (N_787,In_566,In_1735);
and U788 (N_788,In_1434,In_1403);
nor U789 (N_789,In_1578,In_1777);
nand U790 (N_790,In_1240,In_1426);
and U791 (N_791,In_1582,In_1586);
and U792 (N_792,In_2452,In_2009);
xor U793 (N_793,In_811,In_360);
and U794 (N_794,In_515,In_731);
or U795 (N_795,In_344,In_941);
and U796 (N_796,In_860,In_483);
and U797 (N_797,In_136,In_2323);
xnor U798 (N_798,In_305,In_444);
or U799 (N_799,In_685,In_1003);
nor U800 (N_800,In_1274,In_1688);
nor U801 (N_801,In_538,In_381);
or U802 (N_802,In_2166,In_1790);
nor U803 (N_803,In_1670,In_647);
and U804 (N_804,In_228,In_743);
and U805 (N_805,In_66,In_1514);
and U806 (N_806,In_2134,In_1168);
or U807 (N_807,In_1342,In_738);
xnor U808 (N_808,In_436,In_802);
and U809 (N_809,In_833,In_1149);
nand U810 (N_810,In_2435,In_2307);
nor U811 (N_811,In_719,In_1109);
nor U812 (N_812,In_710,In_2189);
nand U813 (N_813,In_1200,In_935);
nor U814 (N_814,In_1889,In_44);
nor U815 (N_815,In_1591,In_977);
xnor U816 (N_816,In_413,In_1055);
or U817 (N_817,In_2098,In_673);
nor U818 (N_818,In_481,In_11);
and U819 (N_819,In_1177,In_1013);
or U820 (N_820,In_715,In_1628);
and U821 (N_821,In_891,In_2020);
nor U822 (N_822,In_1262,In_865);
and U823 (N_823,In_1234,In_1648);
nand U824 (N_824,In_2169,In_424);
xnor U825 (N_825,In_2170,In_476);
nand U826 (N_826,In_1558,In_972);
xor U827 (N_827,In_1333,In_2238);
nand U828 (N_828,In_1027,In_1394);
nand U829 (N_829,In_5,In_1564);
xnor U830 (N_830,In_667,In_1395);
nand U831 (N_831,In_951,In_1620);
xor U832 (N_832,In_1666,In_249);
nor U833 (N_833,In_902,In_1010);
nand U834 (N_834,In_1871,In_1565);
nor U835 (N_835,In_1736,In_1105);
and U836 (N_836,In_2019,In_275);
nand U837 (N_837,In_1720,In_2317);
nor U838 (N_838,In_1322,In_766);
nand U839 (N_839,In_955,In_1011);
nor U840 (N_840,In_2085,In_1533);
or U841 (N_841,In_349,In_994);
or U842 (N_842,In_1873,In_1593);
xor U843 (N_843,In_630,In_512);
or U844 (N_844,In_107,In_756);
nor U845 (N_845,In_670,In_22);
nand U846 (N_846,In_1294,In_2254);
or U847 (N_847,In_488,In_172);
or U848 (N_848,In_153,In_2325);
nor U849 (N_849,In_1987,In_2104);
nor U850 (N_850,In_313,In_1742);
xor U851 (N_851,In_703,In_1473);
nand U852 (N_852,In_1476,In_427);
nor U853 (N_853,In_447,In_1169);
and U854 (N_854,In_29,In_1190);
nor U855 (N_855,In_1886,In_1588);
and U856 (N_856,In_1662,In_1163);
nor U857 (N_857,In_800,In_1504);
nor U858 (N_858,In_1379,In_1211);
xnor U859 (N_859,In_77,In_2028);
xnor U860 (N_860,In_903,In_340);
and U861 (N_861,In_1996,In_2102);
nand U862 (N_862,In_1704,In_641);
xnor U863 (N_863,In_1491,In_2239);
or U864 (N_864,In_262,In_215);
nor U865 (N_865,In_1841,In_1143);
nor U866 (N_866,In_505,In_1935);
nor U867 (N_867,In_49,In_2322);
xnor U868 (N_868,In_140,In_1129);
or U869 (N_869,In_590,In_1561);
xnor U870 (N_870,In_1864,In_986);
xnor U871 (N_871,In_2058,In_617);
nor U872 (N_872,In_1106,In_682);
nand U873 (N_873,In_2462,In_2471);
or U874 (N_874,In_127,In_2464);
xor U875 (N_875,In_1710,In_851);
nand U876 (N_876,In_661,In_603);
and U877 (N_877,In_1083,In_139);
nand U878 (N_878,In_1714,In_529);
xor U879 (N_879,In_2042,In_2129);
nor U880 (N_880,In_974,In_499);
nor U881 (N_881,In_700,In_2299);
xor U882 (N_882,In_2458,In_659);
and U883 (N_883,In_319,In_288);
nor U884 (N_884,In_1929,In_1225);
nor U885 (N_885,In_1250,In_1500);
nor U886 (N_886,In_435,In_2405);
nand U887 (N_887,In_2480,In_1959);
nand U888 (N_888,In_2327,In_614);
nor U889 (N_889,In_1009,In_78);
and U890 (N_890,In_1187,In_2436);
nor U891 (N_891,In_1941,In_1328);
or U892 (N_892,In_442,In_1350);
nand U893 (N_893,In_160,In_352);
nor U894 (N_894,In_2345,In_50);
xor U895 (N_895,In_947,In_2355);
xor U896 (N_896,In_1097,In_1213);
or U897 (N_897,In_1161,In_1404);
nor U898 (N_898,In_656,In_2441);
and U899 (N_899,In_2465,In_1715);
xnor U900 (N_900,In_2346,In_1370);
and U901 (N_901,In_1936,In_1848);
and U902 (N_902,In_265,In_1492);
xor U903 (N_903,In_1546,In_452);
nor U904 (N_904,In_1151,In_1248);
nand U905 (N_905,In_1056,In_393);
xor U906 (N_906,In_2342,In_1622);
and U907 (N_907,In_969,In_999);
and U908 (N_908,In_261,In_1415);
nand U909 (N_909,In_2190,In_783);
xor U910 (N_910,In_1725,In_1336);
or U911 (N_911,In_100,In_1757);
or U912 (N_912,In_99,In_2274);
nand U913 (N_913,In_376,In_1158);
nand U914 (N_914,In_2314,In_304);
xnor U915 (N_915,In_1243,In_26);
or U916 (N_916,In_1368,In_1602);
nor U917 (N_917,In_831,In_2418);
and U918 (N_918,In_1043,In_2371);
nor U919 (N_919,In_253,In_2249);
nor U920 (N_920,In_163,In_1417);
or U921 (N_921,In_2192,In_71);
nor U922 (N_922,In_2383,In_906);
xnor U923 (N_923,In_1146,In_1556);
xnor U924 (N_924,In_830,In_608);
and U925 (N_925,In_1531,In_926);
or U926 (N_926,In_420,In_2285);
or U927 (N_927,In_1878,In_1584);
and U928 (N_928,In_1708,In_1995);
and U929 (N_929,In_2474,In_1926);
xnor U930 (N_930,In_2013,In_1722);
or U931 (N_931,In_1523,In_1991);
and U932 (N_932,In_982,In_1739);
or U933 (N_933,In_1974,In_1549);
and U934 (N_934,In_143,In_2114);
xnor U935 (N_935,In_1,In_1840);
or U936 (N_936,In_2082,In_244);
nand U937 (N_937,In_355,In_775);
and U938 (N_938,In_2263,In_119);
or U939 (N_939,In_653,In_345);
nand U940 (N_940,In_1390,In_1928);
and U941 (N_941,In_25,In_755);
and U942 (N_942,In_1901,In_1137);
xnor U943 (N_943,In_2101,In_250);
nand U944 (N_944,In_1481,In_893);
nor U945 (N_945,In_1389,In_121);
xor U946 (N_946,In_699,In_397);
nor U947 (N_947,In_1609,In_1136);
and U948 (N_948,In_2112,In_1327);
nor U949 (N_949,In_864,In_799);
xnor U950 (N_950,In_767,In_2073);
nor U951 (N_951,In_1156,In_500);
xnor U952 (N_952,In_1538,In_841);
nor U953 (N_953,In_1842,In_1457);
or U954 (N_954,In_2373,In_485);
xor U955 (N_955,In_2382,In_1238);
or U956 (N_956,In_2361,In_2344);
and U957 (N_957,In_474,In_688);
nand U958 (N_958,In_2253,In_170);
nor U959 (N_959,In_2459,In_1927);
nor U960 (N_960,In_1904,In_1320);
nand U961 (N_961,In_1258,In_1241);
or U962 (N_962,In_1820,In_633);
nor U963 (N_963,In_1907,In_356);
and U964 (N_964,In_858,In_1266);
and U965 (N_965,In_2152,In_2328);
nor U966 (N_966,In_534,In_1794);
and U967 (N_967,In_1353,In_325);
xnor U968 (N_968,In_2076,In_692);
xor U969 (N_969,In_961,In_1087);
or U970 (N_970,In_19,In_1774);
xor U971 (N_971,In_2388,In_781);
xnor U972 (N_972,In_2434,In_314);
or U973 (N_973,In_91,In_568);
and U974 (N_974,In_1953,In_1455);
nor U975 (N_975,In_927,In_426);
nor U976 (N_976,In_559,In_10);
xor U977 (N_977,In_1343,In_2186);
nand U978 (N_978,In_297,In_2075);
and U979 (N_979,In_490,In_1512);
xor U980 (N_980,In_334,In_649);
nor U981 (N_981,In_1968,In_2179);
nor U982 (N_982,In_2245,In_2208);
and U983 (N_983,In_1359,In_1332);
and U984 (N_984,In_27,In_1963);
nor U985 (N_985,In_320,In_112);
nand U986 (N_986,In_913,In_1965);
nand U987 (N_987,In_1438,In_815);
or U988 (N_988,In_2059,In_2223);
and U989 (N_989,In_857,In_338);
xnor U990 (N_990,In_279,In_43);
or U991 (N_991,In_2326,In_103);
nand U992 (N_992,In_2440,In_123);
and U993 (N_993,In_351,In_312);
or U994 (N_994,In_2204,In_2366);
nor U995 (N_995,In_1376,In_1555);
nor U996 (N_996,In_1711,In_596);
or U997 (N_997,In_1814,In_210);
and U998 (N_998,In_1534,In_1943);
and U999 (N_999,In_2356,In_990);
xor U1000 (N_1000,In_1942,In_1435);
and U1001 (N_1001,In_434,In_53);
xnor U1002 (N_1002,In_3,In_2067);
or U1003 (N_1003,In_2386,In_142);
nand U1004 (N_1004,In_537,In_28);
and U1005 (N_1005,In_1705,In_108);
nor U1006 (N_1006,In_2427,In_1075);
xor U1007 (N_1007,In_1281,In_2302);
nor U1008 (N_1008,In_1639,In_871);
or U1009 (N_1009,In_2489,In_284);
nor U1010 (N_1010,In_467,In_1372);
xor U1011 (N_1011,In_496,In_2381);
and U1012 (N_1012,In_1448,In_180);
xnor U1013 (N_1013,In_1121,In_1756);
and U1014 (N_1014,In_2168,In_1875);
or U1015 (N_1015,In_1483,In_64);
and U1016 (N_1016,In_1545,In_1084);
and U1017 (N_1017,In_553,In_814);
and U1018 (N_1018,In_1023,In_1299);
nand U1019 (N_1019,In_1283,In_573);
xor U1020 (N_1020,In_1319,In_702);
nor U1021 (N_1021,In_628,In_1782);
and U1022 (N_1022,In_1997,In_790);
nor U1023 (N_1023,In_1433,In_1352);
or U1024 (N_1024,In_1732,In_1684);
or U1025 (N_1025,In_979,In_829);
or U1026 (N_1026,In_758,In_2234);
nor U1027 (N_1027,In_225,In_116);
nor U1028 (N_1028,In_38,In_1583);
and U1029 (N_1029,In_1566,In_503);
xor U1030 (N_1030,In_1899,In_810);
nand U1031 (N_1031,In_498,In_1499);
nor U1032 (N_1032,In_1731,In_101);
and U1033 (N_1033,In_1876,In_2376);
or U1034 (N_1034,In_2141,In_2496);
nor U1035 (N_1035,In_1175,In_93);
nor U1036 (N_1036,In_1025,In_1553);
and U1037 (N_1037,In_1728,In_594);
or U1038 (N_1038,In_2120,In_1999);
nand U1039 (N_1039,In_1453,In_1348);
or U1040 (N_1040,In_2377,In_1465);
xor U1041 (N_1041,In_369,In_1227);
nand U1042 (N_1042,In_611,In_2339);
nand U1043 (N_1043,In_254,In_166);
and U1044 (N_1044,In_1296,In_963);
xor U1045 (N_1045,In_1654,In_1658);
nand U1046 (N_1046,In_1316,In_1930);
or U1047 (N_1047,In_2416,In_2394);
xor U1048 (N_1048,In_227,In_241);
xor U1049 (N_1049,In_1173,In_106);
nand U1050 (N_1050,In_1674,In_2061);
nand U1051 (N_1051,In_1657,In_761);
nand U1052 (N_1052,In_282,In_137);
or U1053 (N_1053,In_1718,In_1071);
nor U1054 (N_1054,In_1058,In_548);
or U1055 (N_1055,In_2228,In_1464);
nor U1056 (N_1056,In_277,In_1519);
or U1057 (N_1057,In_2095,In_2499);
and U1058 (N_1058,In_1171,In_1122);
xnor U1059 (N_1059,In_740,In_1094);
and U1060 (N_1060,In_2218,In_2088);
xnor U1061 (N_1061,In_1914,In_179);
or U1062 (N_1062,In_2300,In_317);
or U1063 (N_1063,In_1765,In_469);
nand U1064 (N_1064,In_780,In_1309);
xnor U1065 (N_1065,In_1165,In_156);
nor U1066 (N_1066,In_1472,In_985);
nor U1067 (N_1067,In_439,In_1263);
nand U1068 (N_1068,In_154,In_409);
and U1069 (N_1069,In_396,In_318);
or U1070 (N_1070,In_2231,In_1902);
nor U1071 (N_1071,In_111,In_923);
and U1072 (N_1072,In_2244,In_1594);
and U1073 (N_1073,In_1724,In_2222);
or U1074 (N_1074,In_765,In_59);
and U1075 (N_1075,In_733,In_330);
and U1076 (N_1076,In_689,In_1251);
nand U1077 (N_1077,In_884,In_348);
nor U1078 (N_1078,In_890,In_2145);
nand U1079 (N_1079,In_527,In_414);
nand U1080 (N_1080,In_258,In_616);
and U1081 (N_1081,In_2150,In_508);
nor U1082 (N_1082,In_510,In_1781);
or U1083 (N_1083,In_493,In_94);
nand U1084 (N_1084,In_39,In_897);
or U1085 (N_1085,In_711,In_2021);
or U1086 (N_1086,In_2433,In_1535);
nor U1087 (N_1087,In_55,In_368);
or U1088 (N_1088,In_2252,In_1905);
nor U1089 (N_1089,In_1619,In_242);
xnor U1090 (N_1090,In_1093,In_383);
and U1091 (N_1091,In_350,In_1932);
and U1092 (N_1092,In_1297,In_1675);
nand U1093 (N_1093,In_1589,In_915);
and U1094 (N_1094,In_917,In_1135);
xor U1095 (N_1095,In_2140,In_480);
nand U1096 (N_1096,In_872,In_2410);
and U1097 (N_1097,In_2259,In_1215);
nand U1098 (N_1098,In_230,In_1659);
or U1099 (N_1099,In_2077,In_1487);
nand U1100 (N_1100,In_1707,In_973);
nand U1101 (N_1101,In_1334,In_1051);
nand U1102 (N_1102,In_298,In_152);
nand U1103 (N_1103,In_191,In_584);
and U1104 (N_1104,In_457,In_266);
and U1105 (N_1105,In_665,In_988);
nor U1106 (N_1106,In_2354,In_2016);
nor U1107 (N_1107,In_674,In_213);
or U1108 (N_1108,In_133,In_2247);
nand U1109 (N_1109,In_1006,In_987);
or U1110 (N_1110,In_2184,In_1680);
nand U1111 (N_1111,In_1347,In_1764);
nor U1112 (N_1112,In_1552,In_518);
nor U1113 (N_1113,In_292,In_1912);
or U1114 (N_1114,In_1160,In_2202);
and U1115 (N_1115,In_1195,In_117);
or U1116 (N_1116,In_1868,In_2165);
nor U1117 (N_1117,In_885,In_259);
xnor U1118 (N_1118,In_1102,In_361);
nand U1119 (N_1119,In_522,In_1833);
or U1120 (N_1120,In_1851,In_1474);
and U1121 (N_1121,In_1308,In_1819);
xnor U1122 (N_1122,In_70,In_1040);
nor U1123 (N_1123,In_2278,In_2012);
nand U1124 (N_1124,In_307,In_2262);
nor U1125 (N_1125,In_898,In_1016);
nand U1126 (N_1126,In_2320,In_1900);
and U1127 (N_1127,In_2357,In_2449);
nor U1128 (N_1128,In_2154,In_470);
or U1129 (N_1129,In_260,In_965);
nand U1130 (N_1130,In_660,In_572);
and U1131 (N_1131,In_840,In_2370);
and U1132 (N_1132,In_1865,In_48);
or U1133 (N_1133,In_894,In_992);
nor U1134 (N_1134,In_1479,In_1539);
nor U1135 (N_1135,In_2142,In_1816);
and U1136 (N_1136,In_1226,In_2246);
nand U1137 (N_1137,In_1214,In_1044);
and U1138 (N_1138,In_744,In_32);
nand U1139 (N_1139,In_75,In_251);
nand U1140 (N_1140,In_1272,In_1331);
or U1141 (N_1141,In_17,In_842);
nand U1142 (N_1142,In_708,In_2203);
or U1143 (N_1143,In_95,In_1356);
nand U1144 (N_1144,In_456,In_640);
xnor U1145 (N_1145,In_2041,In_795);
nand U1146 (N_1146,In_2251,In_666);
xnor U1147 (N_1147,In_1418,In_805);
xor U1148 (N_1148,In_2063,In_2043);
xor U1149 (N_1149,In_1074,In_862);
or U1150 (N_1150,In_134,In_2224);
nand U1151 (N_1151,In_2303,In_2445);
and U1152 (N_1152,In_403,In_2005);
nand U1153 (N_1153,In_8,In_466);
nor U1154 (N_1154,In_2233,In_2257);
nand U1155 (N_1155,In_1989,In_1482);
or U1156 (N_1156,In_541,In_2232);
nand U1157 (N_1157,In_2478,In_401);
nor U1158 (N_1158,In_1623,In_521);
nor U1159 (N_1159,In_675,In_697);
nor U1160 (N_1160,In_868,In_1065);
and U1161 (N_1161,In_741,In_1004);
and U1162 (N_1162,In_725,In_1721);
or U1163 (N_1163,In_431,In_2029);
and U1164 (N_1164,In_1702,In_816);
nor U1165 (N_1165,In_812,In_306);
and U1166 (N_1166,In_97,In_271);
xnor U1167 (N_1167,In_1616,In_506);
or U1168 (N_1168,In_1844,In_1498);
and U1169 (N_1169,In_1752,In_2044);
and U1170 (N_1170,In_1573,In_1230);
nand U1171 (N_1171,In_1399,In_283);
and U1172 (N_1172,In_1367,In_336);
xnor U1173 (N_1173,In_1205,In_1034);
xor U1174 (N_1174,In_1393,In_148);
nor U1175 (N_1175,In_1401,In_40);
nor U1176 (N_1176,In_1738,In_239);
xor U1177 (N_1177,In_1812,In_1540);
and U1178 (N_1178,In_2470,In_423);
nand U1179 (N_1179,In_79,In_1521);
xor U1180 (N_1180,In_218,In_1961);
or U1181 (N_1181,In_2201,In_724);
nor U1182 (N_1182,In_984,In_2003);
or U1183 (N_1183,In_921,In_1815);
nor U1184 (N_1184,In_859,In_1939);
nor U1185 (N_1185,In_264,In_454);
xor U1186 (N_1186,In_1741,In_2213);
nand U1187 (N_1187,In_497,In_645);
xor U1188 (N_1188,In_1505,In_1769);
nand U1189 (N_1189,In_2324,In_63);
nand U1190 (N_1190,In_1219,In_909);
xnor U1191 (N_1191,In_1046,In_1847);
nand U1192 (N_1192,In_1218,In_1783);
nand U1193 (N_1193,In_1326,In_157);
and U1194 (N_1194,In_544,In_1048);
nor U1195 (N_1195,In_928,In_460);
nor U1196 (N_1196,In_1579,In_2351);
nand U1197 (N_1197,In_1268,In_1486);
nor U1198 (N_1198,In_1665,In_1385);
and U1199 (N_1199,In_278,In_2163);
and U1200 (N_1200,In_1066,In_1650);
nor U1201 (N_1201,In_353,In_677);
and U1202 (N_1202,In_964,In_1259);
nand U1203 (N_1203,In_899,In_1478);
nor U1204 (N_1204,In_1611,In_2159);
nand U1205 (N_1205,In_1796,In_2276);
nand U1206 (N_1206,In_415,In_1480);
or U1207 (N_1207,In_539,In_2495);
nor U1208 (N_1208,In_2124,In_782);
or U1209 (N_1209,In_1337,In_664);
nor U1210 (N_1210,In_1128,In_1855);
or U1211 (N_1211,In_1786,In_2437);
or U1212 (N_1212,In_2374,In_694);
nand U1213 (N_1213,In_115,In_648);
nand U1214 (N_1214,In_2167,In_1734);
and U1215 (N_1215,In_1672,In_2267);
and U1216 (N_1216,In_1744,In_2498);
nand U1217 (N_1217,In_1667,In_1892);
and U1218 (N_1218,In_1920,In_2132);
nor U1219 (N_1219,In_1604,In_1580);
and U1220 (N_1220,In_425,In_2113);
xnor U1221 (N_1221,In_83,In_380);
or U1222 (N_1222,In_311,In_626);
xor U1223 (N_1223,In_1518,In_1413);
and U1224 (N_1224,In_1107,In_57);
nor U1225 (N_1225,In_2256,In_1843);
or U1226 (N_1226,In_285,In_321);
or U1227 (N_1227,In_2050,In_2214);
and U1228 (N_1228,In_2413,In_1617);
or U1229 (N_1229,In_422,In_443);
xor U1230 (N_1230,In_1825,In_69);
xor U1231 (N_1231,In_252,In_621);
nand U1232 (N_1232,In_2432,In_2155);
xor U1233 (N_1233,In_226,In_1064);
and U1234 (N_1234,In_1807,In_1683);
nand U1235 (N_1235,In_1203,In_540);
or U1236 (N_1236,In_879,In_146);
nor U1237 (N_1237,In_2456,In_1488);
and U1238 (N_1238,In_1962,In_1747);
nor U1239 (N_1239,In_2430,In_1824);
and U1240 (N_1240,In_224,In_1033);
nand U1241 (N_1241,In_2197,In_1893);
and U1242 (N_1242,In_1469,In_370);
nor U1243 (N_1243,In_13,In_2081);
nor U1244 (N_1244,In_72,In_919);
nand U1245 (N_1245,In_2033,In_895);
xor U1246 (N_1246,In_2375,In_533);
or U1247 (N_1247,In_2443,In_4);
xor U1248 (N_1248,In_1232,In_2469);
xnor U1249 (N_1249,In_1860,In_2210);
xnor U1250 (N_1250,N_581,N_579);
nor U1251 (N_1251,N_738,N_677);
or U1252 (N_1252,N_343,N_815);
xnor U1253 (N_1253,N_486,N_1122);
nor U1254 (N_1254,N_707,N_1091);
or U1255 (N_1255,N_614,N_1143);
or U1256 (N_1256,N_862,N_850);
nand U1257 (N_1257,N_810,N_684);
nand U1258 (N_1258,N_542,N_555);
and U1259 (N_1259,N_252,N_726);
nand U1260 (N_1260,N_73,N_407);
nand U1261 (N_1261,N_488,N_364);
or U1262 (N_1262,N_601,N_247);
or U1263 (N_1263,N_1215,N_144);
xor U1264 (N_1264,N_433,N_122);
or U1265 (N_1265,N_953,N_1118);
and U1266 (N_1266,N_989,N_1181);
nand U1267 (N_1267,N_29,N_422);
nand U1268 (N_1268,N_728,N_33);
nand U1269 (N_1269,N_834,N_593);
and U1270 (N_1270,N_937,N_1115);
and U1271 (N_1271,N_316,N_213);
nand U1272 (N_1272,N_190,N_816);
nor U1273 (N_1273,N_468,N_870);
xor U1274 (N_1274,N_108,N_744);
xnor U1275 (N_1275,N_6,N_1145);
or U1276 (N_1276,N_775,N_991);
nand U1277 (N_1277,N_174,N_1157);
or U1278 (N_1278,N_1092,N_796);
nand U1279 (N_1279,N_175,N_809);
nand U1280 (N_1280,N_261,N_611);
or U1281 (N_1281,N_771,N_354);
or U1282 (N_1282,N_908,N_461);
nor U1283 (N_1283,N_1203,N_1242);
xnor U1284 (N_1284,N_403,N_968);
nor U1285 (N_1285,N_299,N_585);
xor U1286 (N_1286,N_1169,N_177);
and U1287 (N_1287,N_421,N_140);
nand U1288 (N_1288,N_903,N_892);
nor U1289 (N_1289,N_417,N_370);
or U1290 (N_1290,N_401,N_518);
nand U1291 (N_1291,N_376,N_921);
and U1292 (N_1292,N_179,N_764);
xnor U1293 (N_1293,N_625,N_1213);
and U1294 (N_1294,N_839,N_304);
nand U1295 (N_1295,N_363,N_99);
nor U1296 (N_1296,N_1241,N_676);
and U1297 (N_1297,N_694,N_1031);
nor U1298 (N_1298,N_1065,N_909);
and U1299 (N_1299,N_493,N_731);
nand U1300 (N_1300,N_1232,N_624);
xnor U1301 (N_1301,N_83,N_685);
nand U1302 (N_1302,N_754,N_896);
nor U1303 (N_1303,N_784,N_574);
nand U1304 (N_1304,N_180,N_788);
xor U1305 (N_1305,N_923,N_718);
nor U1306 (N_1306,N_498,N_920);
nor U1307 (N_1307,N_96,N_885);
nand U1308 (N_1308,N_380,N_1200);
xnor U1309 (N_1309,N_541,N_702);
nand U1310 (N_1310,N_291,N_1056);
or U1311 (N_1311,N_843,N_353);
nor U1312 (N_1312,N_1196,N_231);
nand U1313 (N_1313,N_860,N_214);
or U1314 (N_1314,N_183,N_564);
nand U1315 (N_1315,N_950,N_966);
nor U1316 (N_1316,N_910,N_698);
nand U1317 (N_1317,N_90,N_104);
nand U1318 (N_1318,N_75,N_1147);
or U1319 (N_1319,N_260,N_836);
nand U1320 (N_1320,N_272,N_878);
nor U1321 (N_1321,N_1030,N_1151);
nor U1322 (N_1322,N_833,N_230);
and U1323 (N_1323,N_1183,N_774);
and U1324 (N_1324,N_884,N_1063);
nor U1325 (N_1325,N_31,N_1037);
or U1326 (N_1326,N_761,N_1022);
nand U1327 (N_1327,N_598,N_1214);
nor U1328 (N_1328,N_510,N_650);
and U1329 (N_1329,N_263,N_543);
and U1330 (N_1330,N_168,N_1134);
xor U1331 (N_1331,N_164,N_476);
or U1332 (N_1332,N_1238,N_780);
and U1333 (N_1333,N_315,N_1139);
xnor U1334 (N_1334,N_1247,N_513);
nand U1335 (N_1335,N_462,N_1166);
nand U1336 (N_1336,N_1076,N_853);
nor U1337 (N_1337,N_922,N_1173);
and U1338 (N_1338,N_826,N_338);
nand U1339 (N_1339,N_596,N_975);
nand U1340 (N_1340,N_557,N_163);
xor U1341 (N_1341,N_1249,N_759);
xnor U1342 (N_1342,N_822,N_592);
or U1343 (N_1343,N_74,N_992);
and U1344 (N_1344,N_235,N_189);
or U1345 (N_1345,N_82,N_1088);
or U1346 (N_1346,N_1137,N_827);
nor U1347 (N_1347,N_730,N_340);
nor U1348 (N_1348,N_248,N_642);
or U1349 (N_1349,N_101,N_446);
or U1350 (N_1350,N_626,N_282);
xor U1351 (N_1351,N_872,N_1006);
and U1352 (N_1352,N_327,N_1226);
xor U1353 (N_1353,N_632,N_719);
or U1354 (N_1354,N_797,N_160);
xor U1355 (N_1355,N_724,N_1164);
nor U1356 (N_1356,N_32,N_11);
nor U1357 (N_1357,N_736,N_1175);
or U1358 (N_1358,N_1054,N_608);
nor U1359 (N_1359,N_1073,N_830);
nor U1360 (N_1360,N_553,N_695);
xor U1361 (N_1361,N_54,N_762);
and U1362 (N_1362,N_944,N_582);
or U1363 (N_1363,N_69,N_1028);
and U1364 (N_1364,N_609,N_118);
and U1365 (N_1365,N_960,N_652);
nand U1366 (N_1366,N_845,N_18);
xnor U1367 (N_1367,N_999,N_386);
xor U1368 (N_1368,N_151,N_628);
or U1369 (N_1369,N_317,N_929);
or U1370 (N_1370,N_52,N_986);
and U1371 (N_1371,N_1007,N_1075);
xnor U1372 (N_1372,N_215,N_755);
nand U1373 (N_1373,N_647,N_454);
nor U1374 (N_1374,N_634,N_977);
or U1375 (N_1375,N_237,N_1083);
and U1376 (N_1376,N_972,N_552);
nor U1377 (N_1377,N_107,N_331);
nor U1378 (N_1378,N_1052,N_259);
nor U1379 (N_1379,N_1219,N_1012);
nand U1380 (N_1380,N_587,N_886);
xor U1381 (N_1381,N_612,N_124);
and U1382 (N_1382,N_89,N_419);
nor U1383 (N_1383,N_741,N_1081);
or U1384 (N_1384,N_915,N_879);
or U1385 (N_1385,N_244,N_1032);
and U1386 (N_1386,N_645,N_1114);
or U1387 (N_1387,N_649,N_692);
or U1388 (N_1388,N_651,N_591);
or U1389 (N_1389,N_450,N_1230);
and U1390 (N_1390,N_727,N_105);
xor U1391 (N_1391,N_1191,N_371);
xnor U1392 (N_1392,N_390,N_538);
and U1393 (N_1393,N_1184,N_508);
xor U1394 (N_1394,N_98,N_389);
nand U1395 (N_1395,N_326,N_320);
or U1396 (N_1396,N_72,N_1246);
or U1397 (N_1397,N_722,N_1106);
xor U1398 (N_1398,N_982,N_324);
or U1399 (N_1399,N_673,N_657);
nor U1400 (N_1400,N_1104,N_152);
or U1401 (N_1401,N_911,N_249);
xor U1402 (N_1402,N_112,N_292);
xor U1403 (N_1403,N_418,N_137);
nor U1404 (N_1404,N_42,N_1228);
nand U1405 (N_1405,N_545,N_391);
or U1406 (N_1406,N_1180,N_1);
nor U1407 (N_1407,N_241,N_671);
nor U1408 (N_1408,N_198,N_372);
or U1409 (N_1409,N_696,N_1165);
xnor U1410 (N_1410,N_811,N_1149);
xor U1411 (N_1411,N_485,N_467);
nor U1412 (N_1412,N_1126,N_571);
nand U1413 (N_1413,N_414,N_1125);
or U1414 (N_1414,N_917,N_448);
and U1415 (N_1415,N_143,N_445);
nor U1416 (N_1416,N_630,N_184);
nand U1417 (N_1417,N_36,N_701);
nor U1418 (N_1418,N_904,N_495);
xor U1419 (N_1419,N_562,N_332);
nand U1420 (N_1420,N_225,N_50);
nand U1421 (N_1421,N_1023,N_37);
nand U1422 (N_1422,N_328,N_773);
and U1423 (N_1423,N_985,N_959);
nand U1424 (N_1424,N_279,N_740);
and U1425 (N_1425,N_998,N_1237);
or U1426 (N_1426,N_117,N_298);
and U1427 (N_1427,N_170,N_392);
nand U1428 (N_1428,N_1005,N_156);
nand U1429 (N_1429,N_23,N_206);
and U1430 (N_1430,N_1205,N_382);
nand U1431 (N_1431,N_1019,N_951);
nand U1432 (N_1432,N_477,N_120);
and U1433 (N_1433,N_690,N_114);
nor U1434 (N_1434,N_34,N_930);
xnor U1435 (N_1435,N_1148,N_66);
nor U1436 (N_1436,N_359,N_511);
nand U1437 (N_1437,N_1162,N_1103);
or U1438 (N_1438,N_396,N_8);
nand U1439 (N_1439,N_1211,N_801);
and U1440 (N_1440,N_110,N_700);
nor U1441 (N_1441,N_28,N_430);
or U1442 (N_1442,N_437,N_682);
nor U1443 (N_1443,N_173,N_566);
or U1444 (N_1444,N_621,N_907);
and U1445 (N_1445,N_303,N_852);
xor U1446 (N_1446,N_240,N_924);
nor U1447 (N_1447,N_519,N_182);
xor U1448 (N_1448,N_1108,N_265);
and U1449 (N_1449,N_308,N_132);
xnor U1450 (N_1450,N_505,N_1155);
nor U1451 (N_1451,N_936,N_1195);
nor U1452 (N_1452,N_293,N_940);
xor U1453 (N_1453,N_306,N_319);
xor U1454 (N_1454,N_1027,N_123);
xor U1455 (N_1455,N_1192,N_1220);
nand U1456 (N_1456,N_507,N_285);
nor U1457 (N_1457,N_341,N_1089);
or U1458 (N_1458,N_35,N_550);
and U1459 (N_1459,N_531,N_1085);
and U1460 (N_1460,N_424,N_350);
nor U1461 (N_1461,N_491,N_51);
nor U1462 (N_1462,N_721,N_674);
nor U1463 (N_1463,N_310,N_436);
nand U1464 (N_1464,N_1011,N_361);
xnor U1465 (N_1465,N_871,N_313);
and U1466 (N_1466,N_1024,N_1017);
or U1467 (N_1467,N_1188,N_116);
xnor U1468 (N_1468,N_578,N_1224);
or U1469 (N_1469,N_346,N_1047);
nand U1470 (N_1470,N_141,N_393);
nand U1471 (N_1471,N_374,N_606);
nand U1472 (N_1472,N_1045,N_239);
nand U1473 (N_1473,N_478,N_869);
nand U1474 (N_1474,N_544,N_1198);
and U1475 (N_1475,N_954,N_357);
nor U1476 (N_1476,N_296,N_136);
or U1477 (N_1477,N_356,N_1077);
or U1478 (N_1478,N_425,N_153);
and U1479 (N_1479,N_1185,N_25);
nand U1480 (N_1480,N_1153,N_381);
nand U1481 (N_1481,N_242,N_567);
or U1482 (N_1482,N_13,N_487);
or U1483 (N_1483,N_752,N_456);
or U1484 (N_1484,N_858,N_147);
nor U1485 (N_1485,N_1016,N_973);
and U1486 (N_1486,N_1001,N_5);
nand U1487 (N_1487,N_148,N_866);
nor U1488 (N_1488,N_238,N_791);
or U1489 (N_1489,N_45,N_49);
nor U1490 (N_1490,N_806,N_600);
nor U1491 (N_1491,N_406,N_334);
and U1492 (N_1492,N_535,N_271);
or U1493 (N_1493,N_415,N_464);
nor U1494 (N_1494,N_347,N_451);
or U1495 (N_1495,N_994,N_127);
nand U1496 (N_1496,N_828,N_349);
and U1497 (N_1497,N_720,N_281);
or U1498 (N_1498,N_536,N_1107);
nor U1499 (N_1499,N_12,N_155);
or U1500 (N_1500,N_1199,N_253);
and U1501 (N_1501,N_447,N_1218);
and U1502 (N_1502,N_800,N_662);
or U1503 (N_1503,N_221,N_440);
and U1504 (N_1504,N_947,N_528);
nand U1505 (N_1505,N_798,N_1204);
or U1506 (N_1506,N_1014,N_743);
nor U1507 (N_1507,N_365,N_438);
and U1508 (N_1508,N_474,N_765);
nor U1509 (N_1509,N_1060,N_1090);
nand U1510 (N_1510,N_1245,N_385);
or U1511 (N_1511,N_342,N_288);
nor U1512 (N_1512,N_67,N_1111);
nand U1513 (N_1513,N_945,N_683);
xnor U1514 (N_1514,N_678,N_1084);
nand U1515 (N_1515,N_368,N_713);
and U1516 (N_1516,N_805,N_680);
xor U1517 (N_1517,N_818,N_409);
and U1518 (N_1518,N_979,N_841);
nor U1519 (N_1519,N_369,N_514);
and U1520 (N_1520,N_348,N_16);
or U1521 (N_1521,N_1105,N_1057);
nand U1522 (N_1522,N_321,N_1174);
xnor U1523 (N_1523,N_355,N_877);
and U1524 (N_1524,N_274,N_126);
and U1525 (N_1525,N_494,N_501);
xnor U1526 (N_1526,N_1100,N_573);
nand U1527 (N_1527,N_1177,N_497);
xnor U1528 (N_1528,N_835,N_295);
or U1529 (N_1529,N_489,N_159);
nand U1530 (N_1530,N_337,N_1116);
and U1531 (N_1531,N_187,N_480);
or U1532 (N_1532,N_704,N_207);
xor U1533 (N_1533,N_14,N_161);
nand U1534 (N_1534,N_837,N_458);
and U1535 (N_1535,N_192,N_1070);
and U1536 (N_1536,N_185,N_842);
and U1537 (N_1537,N_1050,N_946);
or U1538 (N_1538,N_172,N_948);
xnor U1539 (N_1539,N_749,N_918);
nand U1540 (N_1540,N_7,N_873);
xor U1541 (N_1541,N_484,N_20);
nand U1542 (N_1542,N_1051,N_509);
or U1543 (N_1543,N_457,N_919);
or U1544 (N_1544,N_86,N_204);
and U1545 (N_1545,N_1038,N_202);
or U1546 (N_1546,N_831,N_128);
or U1547 (N_1547,N_776,N_932);
nor U1548 (N_1548,N_219,N_15);
nand U1549 (N_1549,N_935,N_167);
nand U1550 (N_1550,N_644,N_890);
or U1551 (N_1551,N_1248,N_974);
and U1552 (N_1552,N_969,N_233);
and U1553 (N_1553,N_595,N_746);
or U1554 (N_1554,N_849,N_635);
and U1555 (N_1555,N_268,N_1033);
nor U1556 (N_1556,N_1161,N_473);
or U1557 (N_1557,N_420,N_887);
nand U1558 (N_1558,N_119,N_53);
nor U1559 (N_1559,N_471,N_226);
xnor U1560 (N_1560,N_181,N_1129);
and U1561 (N_1561,N_532,N_848);
nor U1562 (N_1562,N_659,N_1216);
nor U1563 (N_1563,N_387,N_847);
nor U1564 (N_1564,N_68,N_675);
and U1565 (N_1565,N_335,N_648);
nand U1566 (N_1566,N_199,N_10);
nand U1567 (N_1567,N_1207,N_178);
or U1568 (N_1568,N_782,N_687);
xnor U1569 (N_1569,N_561,N_302);
nand U1570 (N_1570,N_914,N_60);
or U1571 (N_1571,N_522,N_270);
xnor U1572 (N_1572,N_669,N_193);
nand U1573 (N_1573,N_664,N_95);
or U1574 (N_1574,N_1233,N_732);
and U1575 (N_1575,N_1010,N_616);
or U1576 (N_1576,N_250,N_388);
nor U1577 (N_1577,N_266,N_705);
or U1578 (N_1578,N_459,N_875);
nor U1579 (N_1579,N_333,N_1101);
and U1580 (N_1580,N_547,N_435);
and U1581 (N_1581,N_100,N_410);
and U1582 (N_1582,N_269,N_971);
xor U1583 (N_1583,N_844,N_1206);
xnor U1584 (N_1584,N_408,N_1099);
or U1585 (N_1585,N_861,N_723);
and U1586 (N_1586,N_220,N_597);
xor U1587 (N_1587,N_1132,N_789);
and U1588 (N_1588,N_251,N_38);
xnor U1589 (N_1589,N_1035,N_623);
and U1590 (N_1590,N_1036,N_733);
nand U1591 (N_1591,N_820,N_577);
and U1592 (N_1592,N_627,N_526);
nand U1593 (N_1593,N_899,N_1102);
xor U1594 (N_1594,N_358,N_441);
nand U1595 (N_1595,N_1146,N_952);
and U1596 (N_1596,N_91,N_236);
or U1597 (N_1597,N_17,N_134);
nand U1598 (N_1598,N_452,N_146);
and U1599 (N_1599,N_786,N_209);
nand U1600 (N_1600,N_55,N_779);
or U1601 (N_1601,N_729,N_711);
nand U1602 (N_1602,N_305,N_162);
nand U1603 (N_1603,N_981,N_1141);
and U1604 (N_1604,N_617,N_1194);
xor U1605 (N_1605,N_758,N_139);
nor U1606 (N_1606,N_990,N_706);
or U1607 (N_1607,N_1080,N_255);
xor U1608 (N_1608,N_525,N_770);
xor U1609 (N_1609,N_400,N_294);
nand U1610 (N_1610,N_344,N_1098);
nor U1611 (N_1611,N_927,N_745);
nor U1612 (N_1612,N_1234,N_658);
and U1613 (N_1613,N_1117,N_483);
nor U1614 (N_1614,N_245,N_604);
or U1615 (N_1615,N_1078,N_186);
and U1616 (N_1616,N_829,N_1201);
nor U1617 (N_1617,N_336,N_130);
nand U1618 (N_1618,N_366,N_1178);
or U1619 (N_1619,N_121,N_618);
xor U1620 (N_1620,N_48,N_1133);
nor U1621 (N_1621,N_429,N_1061);
nor U1622 (N_1622,N_492,N_565);
nor U1623 (N_1623,N_643,N_1082);
and U1624 (N_1624,N_210,N_379);
nand U1625 (N_1625,N_62,N_449);
or U1626 (N_1626,N_515,N_817);
and U1627 (N_1627,N_902,N_859);
or U1628 (N_1628,N_113,N_276);
nand U1629 (N_1629,N_580,N_1158);
or U1630 (N_1630,N_330,N_699);
nor U1631 (N_1631,N_1168,N_1119);
xnor U1632 (N_1632,N_607,N_273);
nand U1633 (N_1633,N_666,N_1179);
or U1634 (N_1634,N_1172,N_1009);
xor U1635 (N_1635,N_637,N_443);
and U1636 (N_1636,N_619,N_560);
and U1637 (N_1637,N_257,N_1182);
or U1638 (N_1638,N_1240,N_194);
nor U1639 (N_1639,N_30,N_81);
xnor U1640 (N_1640,N_976,N_813);
nand U1641 (N_1641,N_1064,N_135);
nand U1642 (N_1642,N_444,N_748);
xnor U1643 (N_1643,N_1049,N_803);
nor U1644 (N_1644,N_229,N_176);
nor U1645 (N_1645,N_1140,N_405);
nor U1646 (N_1646,N_802,N_938);
nand U1647 (N_1647,N_322,N_523);
xnor U1648 (N_1648,N_778,N_21);
xor U1649 (N_1649,N_360,N_1044);
nor U1650 (N_1650,N_661,N_1187);
nor U1651 (N_1651,N_1208,N_1244);
nor U1652 (N_1652,N_1167,N_1041);
xnor U1653 (N_1653,N_466,N_216);
or U1654 (N_1654,N_39,N_27);
xnor U1655 (N_1655,N_165,N_962);
nand U1656 (N_1656,N_1002,N_70);
nor U1657 (N_1657,N_807,N_863);
or U1658 (N_1658,N_739,N_1095);
nor U1659 (N_1659,N_636,N_957);
nor U1660 (N_1660,N_825,N_463);
nor U1661 (N_1661,N_963,N_1212);
xor U1662 (N_1662,N_24,N_212);
and U1663 (N_1663,N_777,N_772);
xnor U1664 (N_1664,N_1110,N_1176);
nor U1665 (N_1665,N_1229,N_599);
xor U1666 (N_1666,N_943,N_1046);
nor U1667 (N_1667,N_329,N_399);
nand U1668 (N_1668,N_808,N_1068);
xnor U1669 (N_1669,N_679,N_1144);
nor U1670 (N_1670,N_256,N_898);
nand U1671 (N_1671,N_1015,N_769);
nor U1672 (N_1672,N_103,N_1039);
nand U1673 (N_1673,N_402,N_428);
nor U1674 (N_1674,N_693,N_783);
xnor U1675 (N_1675,N_865,N_812);
and U1676 (N_1676,N_93,N_1021);
xor U1677 (N_1677,N_1026,N_613);
nand U1678 (N_1678,N_715,N_667);
xor U1679 (N_1679,N_714,N_224);
xor U1680 (N_1680,N_1072,N_590);
and U1681 (N_1681,N_785,N_767);
nor U1682 (N_1682,N_1067,N_1113);
nor U1683 (N_1683,N_529,N_551);
nand U1684 (N_1684,N_925,N_314);
xor U1685 (N_1685,N_559,N_211);
or U1686 (N_1686,N_821,N_218);
and U1687 (N_1687,N_799,N_1152);
nor U1688 (N_1688,N_300,N_900);
and U1689 (N_1689,N_716,N_57);
nor U1690 (N_1690,N_1079,N_470);
or U1691 (N_1691,N_267,N_157);
xnor U1692 (N_1692,N_46,N_1042);
xor U1693 (N_1693,N_431,N_691);
nor U1694 (N_1694,N_854,N_94);
nand U1695 (N_1695,N_188,N_59);
xnor U1696 (N_1696,N_78,N_524);
xor U1697 (N_1697,N_232,N_790);
xor U1698 (N_1698,N_594,N_534);
and U1699 (N_1699,N_1135,N_1004);
nand U1700 (N_1700,N_620,N_115);
nand U1701 (N_1701,N_201,N_275);
or U1702 (N_1702,N_43,N_753);
nor U1703 (N_1703,N_913,N_1130);
nand U1704 (N_1704,N_109,N_92);
xnor U1705 (N_1705,N_373,N_196);
nand U1706 (N_1706,N_318,N_1048);
nor U1707 (N_1707,N_40,N_404);
and U1708 (N_1708,N_325,N_287);
nand U1709 (N_1709,N_56,N_301);
and U1710 (N_1710,N_965,N_222);
nand U1711 (N_1711,N_191,N_297);
or U1712 (N_1712,N_423,N_1223);
or U1713 (N_1713,N_416,N_1059);
and U1714 (N_1714,N_377,N_22);
nand U1715 (N_1715,N_610,N_154);
xnor U1716 (N_1716,N_670,N_88);
nand U1717 (N_1717,N_432,N_756);
and U1718 (N_1718,N_166,N_961);
nand U1719 (N_1719,N_516,N_984);
nor U1720 (N_1720,N_465,N_264);
nand U1721 (N_1721,N_537,N_768);
nor U1722 (N_1722,N_472,N_583);
or U1723 (N_1723,N_928,N_1074);
nor U1724 (N_1724,N_1124,N_970);
or U1725 (N_1725,N_996,N_427);
and U1726 (N_1726,N_540,N_978);
xor U1727 (N_1727,N_575,N_995);
or U1728 (N_1728,N_663,N_1150);
nor U1729 (N_1729,N_530,N_411);
xor U1730 (N_1730,N_686,N_26);
or U1731 (N_1731,N_1193,N_517);
nand U1732 (N_1732,N_895,N_362);
nand U1733 (N_1733,N_1121,N_85);
or U1734 (N_1734,N_106,N_169);
nor U1735 (N_1735,N_548,N_864);
nand U1736 (N_1736,N_983,N_129);
nand U1737 (N_1737,N_641,N_703);
nand U1738 (N_1738,N_1013,N_629);
nor U1739 (N_1739,N_1069,N_1000);
nand U1740 (N_1740,N_208,N_988);
nor U1741 (N_1741,N_9,N_640);
xnor U1742 (N_1742,N_747,N_1243);
xnor U1743 (N_1743,N_568,N_352);
nor U1744 (N_1744,N_1197,N_503);
nor U1745 (N_1745,N_1020,N_149);
nor U1746 (N_1746,N_967,N_793);
nor U1747 (N_1747,N_384,N_868);
or U1748 (N_1748,N_460,N_1210);
xor U1749 (N_1749,N_556,N_64);
nand U1750 (N_1750,N_77,N_905);
and U1751 (N_1751,N_760,N_993);
nor U1752 (N_1752,N_1171,N_312);
or U1753 (N_1753,N_906,N_912);
nor U1754 (N_1754,N_258,N_708);
nand U1755 (N_1755,N_781,N_111);
and U1756 (N_1756,N_717,N_655);
or U1757 (N_1757,N_897,N_1109);
xor U1758 (N_1758,N_874,N_546);
nor U1759 (N_1759,N_603,N_883);
and U1760 (N_1760,N_1040,N_709);
nor U1761 (N_1761,N_1222,N_1136);
and U1762 (N_1762,N_234,N_889);
and U1763 (N_1763,N_145,N_1055);
xnor U1764 (N_1764,N_855,N_413);
or U1765 (N_1765,N_665,N_856);
nand U1766 (N_1766,N_71,N_378);
nor U1767 (N_1767,N_931,N_1160);
xor U1768 (N_1768,N_725,N_997);
nor U1769 (N_1769,N_563,N_1018);
nor U1770 (N_1770,N_901,N_1120);
nand U1771 (N_1771,N_4,N_1159);
nand U1772 (N_1772,N_197,N_520);
nor U1773 (N_1773,N_787,N_277);
nor U1774 (N_1774,N_710,N_339);
xor U1775 (N_1775,N_615,N_794);
and U1776 (N_1776,N_949,N_737);
nor U1777 (N_1777,N_469,N_502);
xnor U1778 (N_1778,N_751,N_602);
and U1779 (N_1779,N_397,N_521);
nor U1780 (N_1780,N_734,N_47);
and U1781 (N_1781,N_65,N_284);
xor U1782 (N_1782,N_383,N_1123);
or U1783 (N_1783,N_576,N_639);
nand U1784 (N_1784,N_654,N_125);
nand U1785 (N_1785,N_980,N_496);
and U1786 (N_1786,N_394,N_1239);
nand U1787 (N_1787,N_804,N_1034);
or U1788 (N_1788,N_1127,N_0);
nand U1789 (N_1789,N_1094,N_857);
nand U1790 (N_1790,N_569,N_1087);
nor U1791 (N_1791,N_1170,N_819);
nand U1792 (N_1792,N_133,N_1062);
xnor U1793 (N_1793,N_1003,N_688);
nor U1794 (N_1794,N_792,N_309);
nor U1795 (N_1795,N_572,N_490);
nand U1796 (N_1796,N_1128,N_1043);
xor U1797 (N_1797,N_1227,N_823);
nand U1798 (N_1798,N_283,N_891);
xor U1799 (N_1799,N_171,N_881);
nand U1800 (N_1800,N_205,N_527);
xnor U1801 (N_1801,N_323,N_1221);
and U1802 (N_1802,N_504,N_712);
nor U1803 (N_1803,N_311,N_1202);
nand U1804 (N_1804,N_286,N_44);
nor U1805 (N_1805,N_243,N_1112);
xnor U1806 (N_1806,N_1008,N_1029);
xnor U1807 (N_1807,N_832,N_512);
and U1808 (N_1808,N_876,N_668);
xor U1809 (N_1809,N_638,N_646);
nand U1810 (N_1810,N_138,N_941);
nor U1811 (N_1811,N_1236,N_223);
nor U1812 (N_1812,N_442,N_475);
and U1813 (N_1813,N_846,N_1190);
nand U1814 (N_1814,N_412,N_750);
and U1815 (N_1815,N_814,N_766);
nor U1816 (N_1816,N_150,N_549);
nor U1817 (N_1817,N_1093,N_500);
and U1818 (N_1818,N_1217,N_3);
nand U1819 (N_1819,N_203,N_1163);
and U1820 (N_1820,N_942,N_453);
nor U1821 (N_1821,N_280,N_97);
and U1822 (N_1822,N_742,N_227);
xor U1823 (N_1823,N_76,N_228);
nor U1824 (N_1824,N_689,N_586);
or U1825 (N_1825,N_351,N_63);
or U1826 (N_1826,N_795,N_499);
or U1827 (N_1827,N_1071,N_633);
or U1828 (N_1828,N_345,N_838);
and U1829 (N_1829,N_41,N_1186);
or U1830 (N_1830,N_558,N_87);
nor U1831 (N_1831,N_939,N_735);
xor U1832 (N_1832,N_254,N_894);
nand U1833 (N_1833,N_672,N_80);
or U1834 (N_1834,N_1231,N_506);
nand U1835 (N_1835,N_697,N_955);
nor U1836 (N_1836,N_622,N_367);
nor U1837 (N_1837,N_455,N_882);
or U1838 (N_1838,N_1138,N_660);
or U1839 (N_1839,N_102,N_757);
or U1840 (N_1840,N_2,N_1154);
nor U1841 (N_1841,N_1209,N_58);
nand U1842 (N_1842,N_1189,N_653);
and U1843 (N_1843,N_398,N_375);
xnor U1844 (N_1844,N_926,N_1058);
or U1845 (N_1845,N_958,N_1086);
and U1846 (N_1846,N_289,N_142);
nand U1847 (N_1847,N_656,N_867);
and U1848 (N_1848,N_1131,N_158);
nand U1849 (N_1849,N_1142,N_290);
xor U1850 (N_1850,N_246,N_584);
or U1851 (N_1851,N_278,N_605);
xor U1852 (N_1852,N_79,N_763);
or U1853 (N_1853,N_840,N_61);
nand U1854 (N_1854,N_1225,N_934);
nand U1855 (N_1855,N_681,N_479);
or U1856 (N_1856,N_195,N_888);
nor U1857 (N_1857,N_916,N_824);
or U1858 (N_1858,N_893,N_131);
and U1859 (N_1859,N_1096,N_1066);
or U1860 (N_1860,N_439,N_987);
nor U1861 (N_1861,N_481,N_880);
xnor U1862 (N_1862,N_395,N_1097);
and U1863 (N_1863,N_482,N_1156);
and U1864 (N_1864,N_570,N_1235);
xnor U1865 (N_1865,N_84,N_631);
or U1866 (N_1866,N_19,N_933);
and U1867 (N_1867,N_589,N_588);
xnor U1868 (N_1868,N_851,N_200);
xnor U1869 (N_1869,N_1025,N_1053);
or U1870 (N_1870,N_533,N_434);
nor U1871 (N_1871,N_554,N_307);
or U1872 (N_1872,N_964,N_539);
nor U1873 (N_1873,N_217,N_956);
and U1874 (N_1874,N_426,N_262);
and U1875 (N_1875,N_166,N_580);
nand U1876 (N_1876,N_659,N_428);
nand U1877 (N_1877,N_762,N_1203);
nand U1878 (N_1878,N_437,N_1178);
xnor U1879 (N_1879,N_1208,N_857);
or U1880 (N_1880,N_189,N_546);
and U1881 (N_1881,N_65,N_1152);
nand U1882 (N_1882,N_954,N_664);
nor U1883 (N_1883,N_430,N_690);
nor U1884 (N_1884,N_651,N_1210);
or U1885 (N_1885,N_622,N_303);
nor U1886 (N_1886,N_267,N_1214);
nor U1887 (N_1887,N_478,N_656);
and U1888 (N_1888,N_197,N_843);
and U1889 (N_1889,N_325,N_612);
nor U1890 (N_1890,N_775,N_737);
nor U1891 (N_1891,N_1061,N_592);
nor U1892 (N_1892,N_762,N_450);
nand U1893 (N_1893,N_404,N_566);
nor U1894 (N_1894,N_796,N_277);
xnor U1895 (N_1895,N_576,N_692);
xor U1896 (N_1896,N_771,N_515);
xor U1897 (N_1897,N_1097,N_1096);
nor U1898 (N_1898,N_230,N_352);
nand U1899 (N_1899,N_520,N_639);
nor U1900 (N_1900,N_756,N_283);
or U1901 (N_1901,N_806,N_1199);
nor U1902 (N_1902,N_746,N_640);
nor U1903 (N_1903,N_265,N_1241);
and U1904 (N_1904,N_316,N_1151);
nand U1905 (N_1905,N_206,N_767);
xor U1906 (N_1906,N_32,N_147);
nand U1907 (N_1907,N_276,N_442);
or U1908 (N_1908,N_591,N_85);
and U1909 (N_1909,N_892,N_763);
nor U1910 (N_1910,N_855,N_587);
xnor U1911 (N_1911,N_229,N_991);
nor U1912 (N_1912,N_487,N_679);
xor U1913 (N_1913,N_981,N_170);
xor U1914 (N_1914,N_1163,N_840);
nand U1915 (N_1915,N_1246,N_370);
nand U1916 (N_1916,N_1223,N_1246);
nand U1917 (N_1917,N_613,N_989);
xor U1918 (N_1918,N_962,N_484);
or U1919 (N_1919,N_440,N_418);
or U1920 (N_1920,N_241,N_461);
and U1921 (N_1921,N_716,N_261);
xnor U1922 (N_1922,N_334,N_747);
and U1923 (N_1923,N_955,N_554);
and U1924 (N_1924,N_1242,N_1113);
and U1925 (N_1925,N_1091,N_41);
nand U1926 (N_1926,N_162,N_109);
nand U1927 (N_1927,N_38,N_284);
or U1928 (N_1928,N_452,N_395);
nor U1929 (N_1929,N_452,N_770);
and U1930 (N_1930,N_1195,N_682);
nor U1931 (N_1931,N_530,N_748);
or U1932 (N_1932,N_438,N_299);
and U1933 (N_1933,N_1083,N_1079);
and U1934 (N_1934,N_707,N_495);
and U1935 (N_1935,N_1017,N_239);
nand U1936 (N_1936,N_239,N_1067);
xnor U1937 (N_1937,N_101,N_1139);
or U1938 (N_1938,N_17,N_239);
nand U1939 (N_1939,N_433,N_773);
and U1940 (N_1940,N_1194,N_1073);
nand U1941 (N_1941,N_493,N_718);
nor U1942 (N_1942,N_966,N_195);
and U1943 (N_1943,N_70,N_700);
and U1944 (N_1944,N_599,N_1022);
and U1945 (N_1945,N_1216,N_1196);
and U1946 (N_1946,N_528,N_53);
and U1947 (N_1947,N_964,N_1190);
nand U1948 (N_1948,N_1113,N_386);
xnor U1949 (N_1949,N_1181,N_941);
nor U1950 (N_1950,N_763,N_110);
xnor U1951 (N_1951,N_256,N_84);
xor U1952 (N_1952,N_827,N_672);
nand U1953 (N_1953,N_909,N_997);
xor U1954 (N_1954,N_1104,N_447);
and U1955 (N_1955,N_447,N_599);
or U1956 (N_1956,N_1063,N_1176);
nand U1957 (N_1957,N_394,N_465);
nor U1958 (N_1958,N_877,N_607);
and U1959 (N_1959,N_355,N_126);
xor U1960 (N_1960,N_566,N_498);
and U1961 (N_1961,N_866,N_1012);
or U1962 (N_1962,N_377,N_638);
and U1963 (N_1963,N_416,N_394);
and U1964 (N_1964,N_1014,N_166);
xor U1965 (N_1965,N_406,N_958);
and U1966 (N_1966,N_1111,N_988);
and U1967 (N_1967,N_544,N_1074);
and U1968 (N_1968,N_683,N_71);
and U1969 (N_1969,N_576,N_764);
nor U1970 (N_1970,N_1018,N_49);
or U1971 (N_1971,N_1214,N_838);
xnor U1972 (N_1972,N_64,N_1047);
nand U1973 (N_1973,N_1216,N_716);
or U1974 (N_1974,N_246,N_465);
nor U1975 (N_1975,N_763,N_273);
nor U1976 (N_1976,N_104,N_693);
nand U1977 (N_1977,N_1119,N_785);
or U1978 (N_1978,N_1035,N_219);
nand U1979 (N_1979,N_504,N_688);
nor U1980 (N_1980,N_110,N_268);
or U1981 (N_1981,N_1194,N_587);
and U1982 (N_1982,N_784,N_236);
and U1983 (N_1983,N_165,N_542);
nand U1984 (N_1984,N_846,N_786);
and U1985 (N_1985,N_236,N_459);
nor U1986 (N_1986,N_889,N_643);
nand U1987 (N_1987,N_176,N_801);
nor U1988 (N_1988,N_1025,N_468);
and U1989 (N_1989,N_3,N_61);
or U1990 (N_1990,N_554,N_1212);
nand U1991 (N_1991,N_821,N_1207);
or U1992 (N_1992,N_1194,N_257);
nand U1993 (N_1993,N_263,N_343);
xor U1994 (N_1994,N_52,N_3);
nor U1995 (N_1995,N_680,N_1154);
nand U1996 (N_1996,N_1008,N_773);
nor U1997 (N_1997,N_377,N_488);
xor U1998 (N_1998,N_1083,N_849);
nand U1999 (N_1999,N_783,N_1208);
and U2000 (N_2000,N_555,N_13);
or U2001 (N_2001,N_884,N_765);
nor U2002 (N_2002,N_771,N_1117);
nor U2003 (N_2003,N_570,N_1179);
xnor U2004 (N_2004,N_220,N_1030);
and U2005 (N_2005,N_1248,N_893);
and U2006 (N_2006,N_339,N_1022);
or U2007 (N_2007,N_462,N_556);
and U2008 (N_2008,N_719,N_68);
xor U2009 (N_2009,N_31,N_1074);
nand U2010 (N_2010,N_201,N_477);
nor U2011 (N_2011,N_28,N_455);
or U2012 (N_2012,N_684,N_453);
and U2013 (N_2013,N_413,N_1158);
xnor U2014 (N_2014,N_187,N_640);
nor U2015 (N_2015,N_265,N_165);
or U2016 (N_2016,N_248,N_233);
nor U2017 (N_2017,N_109,N_457);
nor U2018 (N_2018,N_634,N_951);
nor U2019 (N_2019,N_264,N_1179);
xnor U2020 (N_2020,N_803,N_945);
nor U2021 (N_2021,N_669,N_564);
nand U2022 (N_2022,N_345,N_308);
nor U2023 (N_2023,N_1205,N_848);
nor U2024 (N_2024,N_1087,N_1076);
or U2025 (N_2025,N_1062,N_1219);
xnor U2026 (N_2026,N_32,N_1232);
xor U2027 (N_2027,N_755,N_829);
or U2028 (N_2028,N_253,N_1137);
or U2029 (N_2029,N_916,N_890);
and U2030 (N_2030,N_967,N_586);
nor U2031 (N_2031,N_1014,N_727);
xnor U2032 (N_2032,N_1231,N_571);
nor U2033 (N_2033,N_238,N_381);
or U2034 (N_2034,N_72,N_390);
or U2035 (N_2035,N_251,N_166);
nor U2036 (N_2036,N_1204,N_3);
or U2037 (N_2037,N_823,N_933);
or U2038 (N_2038,N_373,N_532);
nand U2039 (N_2039,N_545,N_1218);
nor U2040 (N_2040,N_216,N_320);
nand U2041 (N_2041,N_1019,N_802);
or U2042 (N_2042,N_1181,N_80);
nand U2043 (N_2043,N_498,N_595);
xnor U2044 (N_2044,N_379,N_15);
xor U2045 (N_2045,N_394,N_1052);
nand U2046 (N_2046,N_159,N_369);
or U2047 (N_2047,N_268,N_512);
xor U2048 (N_2048,N_686,N_477);
or U2049 (N_2049,N_645,N_374);
and U2050 (N_2050,N_351,N_441);
or U2051 (N_2051,N_42,N_1157);
or U2052 (N_2052,N_664,N_631);
or U2053 (N_2053,N_666,N_244);
xnor U2054 (N_2054,N_597,N_1047);
xor U2055 (N_2055,N_1046,N_183);
and U2056 (N_2056,N_189,N_905);
nor U2057 (N_2057,N_491,N_902);
nand U2058 (N_2058,N_53,N_744);
and U2059 (N_2059,N_446,N_1245);
and U2060 (N_2060,N_356,N_1234);
xor U2061 (N_2061,N_1018,N_933);
nor U2062 (N_2062,N_701,N_994);
nand U2063 (N_2063,N_1018,N_277);
xnor U2064 (N_2064,N_64,N_650);
or U2065 (N_2065,N_207,N_393);
xnor U2066 (N_2066,N_274,N_45);
nor U2067 (N_2067,N_221,N_467);
xnor U2068 (N_2068,N_1037,N_346);
xor U2069 (N_2069,N_669,N_786);
or U2070 (N_2070,N_40,N_233);
or U2071 (N_2071,N_944,N_1191);
xnor U2072 (N_2072,N_99,N_1046);
and U2073 (N_2073,N_15,N_455);
or U2074 (N_2074,N_287,N_59);
nor U2075 (N_2075,N_1044,N_286);
nor U2076 (N_2076,N_224,N_1151);
xor U2077 (N_2077,N_243,N_292);
xor U2078 (N_2078,N_179,N_444);
xnor U2079 (N_2079,N_807,N_49);
and U2080 (N_2080,N_687,N_10);
and U2081 (N_2081,N_1158,N_368);
or U2082 (N_2082,N_401,N_707);
nand U2083 (N_2083,N_901,N_891);
nor U2084 (N_2084,N_1059,N_105);
or U2085 (N_2085,N_1180,N_970);
nand U2086 (N_2086,N_915,N_225);
or U2087 (N_2087,N_315,N_484);
xnor U2088 (N_2088,N_1045,N_634);
or U2089 (N_2089,N_715,N_140);
and U2090 (N_2090,N_172,N_689);
nand U2091 (N_2091,N_268,N_75);
nor U2092 (N_2092,N_1127,N_490);
or U2093 (N_2093,N_613,N_1093);
or U2094 (N_2094,N_1019,N_965);
nand U2095 (N_2095,N_1236,N_559);
xnor U2096 (N_2096,N_185,N_980);
nor U2097 (N_2097,N_890,N_509);
nor U2098 (N_2098,N_1142,N_395);
nand U2099 (N_2099,N_359,N_560);
xor U2100 (N_2100,N_744,N_364);
nand U2101 (N_2101,N_703,N_193);
and U2102 (N_2102,N_250,N_282);
nor U2103 (N_2103,N_570,N_514);
or U2104 (N_2104,N_258,N_116);
xnor U2105 (N_2105,N_1056,N_1053);
nor U2106 (N_2106,N_598,N_27);
nor U2107 (N_2107,N_356,N_463);
or U2108 (N_2108,N_625,N_872);
or U2109 (N_2109,N_1054,N_49);
and U2110 (N_2110,N_830,N_1200);
and U2111 (N_2111,N_236,N_85);
nor U2112 (N_2112,N_707,N_36);
nor U2113 (N_2113,N_986,N_976);
or U2114 (N_2114,N_1094,N_102);
xnor U2115 (N_2115,N_731,N_342);
nand U2116 (N_2116,N_7,N_619);
nor U2117 (N_2117,N_924,N_289);
or U2118 (N_2118,N_27,N_448);
nand U2119 (N_2119,N_919,N_244);
and U2120 (N_2120,N_95,N_670);
and U2121 (N_2121,N_1099,N_1087);
and U2122 (N_2122,N_1087,N_1025);
nand U2123 (N_2123,N_156,N_744);
nand U2124 (N_2124,N_1070,N_777);
xor U2125 (N_2125,N_1075,N_1051);
xnor U2126 (N_2126,N_883,N_638);
or U2127 (N_2127,N_683,N_724);
and U2128 (N_2128,N_535,N_537);
xor U2129 (N_2129,N_61,N_94);
nor U2130 (N_2130,N_1034,N_918);
xnor U2131 (N_2131,N_516,N_1107);
or U2132 (N_2132,N_575,N_299);
or U2133 (N_2133,N_839,N_84);
nand U2134 (N_2134,N_369,N_1193);
and U2135 (N_2135,N_905,N_263);
xnor U2136 (N_2136,N_1203,N_28);
and U2137 (N_2137,N_1203,N_743);
or U2138 (N_2138,N_553,N_894);
xor U2139 (N_2139,N_673,N_1195);
xor U2140 (N_2140,N_510,N_726);
or U2141 (N_2141,N_261,N_347);
xnor U2142 (N_2142,N_1161,N_524);
and U2143 (N_2143,N_14,N_289);
xnor U2144 (N_2144,N_898,N_556);
nand U2145 (N_2145,N_98,N_419);
nor U2146 (N_2146,N_124,N_235);
nor U2147 (N_2147,N_650,N_1071);
nor U2148 (N_2148,N_755,N_852);
nor U2149 (N_2149,N_1193,N_42);
and U2150 (N_2150,N_671,N_232);
xnor U2151 (N_2151,N_689,N_697);
nor U2152 (N_2152,N_147,N_627);
and U2153 (N_2153,N_91,N_1128);
nand U2154 (N_2154,N_933,N_1151);
nor U2155 (N_2155,N_709,N_665);
nor U2156 (N_2156,N_713,N_373);
and U2157 (N_2157,N_494,N_215);
nand U2158 (N_2158,N_955,N_636);
and U2159 (N_2159,N_384,N_690);
xor U2160 (N_2160,N_715,N_227);
xor U2161 (N_2161,N_391,N_1058);
or U2162 (N_2162,N_564,N_886);
and U2163 (N_2163,N_483,N_683);
or U2164 (N_2164,N_385,N_602);
xnor U2165 (N_2165,N_416,N_1076);
and U2166 (N_2166,N_826,N_1184);
nand U2167 (N_2167,N_331,N_551);
xnor U2168 (N_2168,N_1151,N_495);
xor U2169 (N_2169,N_75,N_586);
xor U2170 (N_2170,N_141,N_326);
xor U2171 (N_2171,N_1239,N_785);
nor U2172 (N_2172,N_1043,N_627);
xnor U2173 (N_2173,N_418,N_667);
xnor U2174 (N_2174,N_160,N_785);
xor U2175 (N_2175,N_402,N_1056);
nor U2176 (N_2176,N_1229,N_304);
nand U2177 (N_2177,N_1098,N_166);
or U2178 (N_2178,N_892,N_1021);
xor U2179 (N_2179,N_270,N_449);
nand U2180 (N_2180,N_498,N_329);
nand U2181 (N_2181,N_460,N_401);
nand U2182 (N_2182,N_1211,N_1078);
or U2183 (N_2183,N_1219,N_626);
or U2184 (N_2184,N_96,N_29);
nand U2185 (N_2185,N_116,N_845);
nor U2186 (N_2186,N_69,N_111);
nor U2187 (N_2187,N_1199,N_667);
nand U2188 (N_2188,N_351,N_864);
nand U2189 (N_2189,N_1159,N_174);
xor U2190 (N_2190,N_558,N_778);
xnor U2191 (N_2191,N_615,N_885);
or U2192 (N_2192,N_128,N_1043);
xor U2193 (N_2193,N_1080,N_615);
xor U2194 (N_2194,N_376,N_142);
and U2195 (N_2195,N_898,N_34);
nand U2196 (N_2196,N_509,N_1095);
xnor U2197 (N_2197,N_885,N_779);
and U2198 (N_2198,N_42,N_932);
nor U2199 (N_2199,N_55,N_673);
xor U2200 (N_2200,N_1060,N_610);
xnor U2201 (N_2201,N_977,N_198);
and U2202 (N_2202,N_947,N_617);
nor U2203 (N_2203,N_285,N_409);
and U2204 (N_2204,N_438,N_423);
and U2205 (N_2205,N_509,N_839);
and U2206 (N_2206,N_855,N_376);
nor U2207 (N_2207,N_240,N_474);
and U2208 (N_2208,N_1109,N_395);
or U2209 (N_2209,N_819,N_582);
nor U2210 (N_2210,N_1224,N_1006);
nand U2211 (N_2211,N_185,N_677);
nand U2212 (N_2212,N_789,N_244);
xnor U2213 (N_2213,N_650,N_0);
or U2214 (N_2214,N_191,N_125);
xnor U2215 (N_2215,N_52,N_913);
nand U2216 (N_2216,N_1050,N_1030);
and U2217 (N_2217,N_394,N_97);
or U2218 (N_2218,N_765,N_785);
and U2219 (N_2219,N_1013,N_1240);
or U2220 (N_2220,N_932,N_850);
nand U2221 (N_2221,N_705,N_984);
or U2222 (N_2222,N_808,N_85);
nand U2223 (N_2223,N_758,N_1240);
and U2224 (N_2224,N_1130,N_86);
xor U2225 (N_2225,N_756,N_991);
and U2226 (N_2226,N_62,N_196);
nor U2227 (N_2227,N_519,N_1101);
xnor U2228 (N_2228,N_955,N_126);
and U2229 (N_2229,N_1043,N_303);
or U2230 (N_2230,N_101,N_952);
nand U2231 (N_2231,N_1244,N_785);
or U2232 (N_2232,N_373,N_267);
nor U2233 (N_2233,N_1047,N_604);
nor U2234 (N_2234,N_1000,N_677);
xnor U2235 (N_2235,N_21,N_99);
and U2236 (N_2236,N_981,N_876);
nor U2237 (N_2237,N_1075,N_27);
nand U2238 (N_2238,N_101,N_1108);
xnor U2239 (N_2239,N_739,N_604);
nand U2240 (N_2240,N_958,N_820);
nand U2241 (N_2241,N_527,N_563);
nor U2242 (N_2242,N_977,N_1074);
nand U2243 (N_2243,N_383,N_839);
or U2244 (N_2244,N_377,N_69);
or U2245 (N_2245,N_338,N_354);
nor U2246 (N_2246,N_389,N_397);
nor U2247 (N_2247,N_427,N_106);
nor U2248 (N_2248,N_312,N_545);
xor U2249 (N_2249,N_571,N_1129);
or U2250 (N_2250,N_1240,N_559);
xor U2251 (N_2251,N_1003,N_964);
xor U2252 (N_2252,N_1000,N_968);
or U2253 (N_2253,N_169,N_697);
or U2254 (N_2254,N_726,N_644);
and U2255 (N_2255,N_816,N_863);
or U2256 (N_2256,N_303,N_319);
and U2257 (N_2257,N_782,N_610);
nor U2258 (N_2258,N_431,N_474);
xnor U2259 (N_2259,N_361,N_81);
or U2260 (N_2260,N_1016,N_156);
and U2261 (N_2261,N_671,N_186);
nor U2262 (N_2262,N_1189,N_971);
nor U2263 (N_2263,N_131,N_862);
and U2264 (N_2264,N_182,N_1062);
and U2265 (N_2265,N_139,N_316);
or U2266 (N_2266,N_428,N_427);
or U2267 (N_2267,N_1168,N_465);
and U2268 (N_2268,N_483,N_711);
nor U2269 (N_2269,N_415,N_292);
xnor U2270 (N_2270,N_1008,N_1125);
and U2271 (N_2271,N_1173,N_1202);
and U2272 (N_2272,N_1176,N_40);
or U2273 (N_2273,N_796,N_1201);
and U2274 (N_2274,N_1153,N_1015);
xor U2275 (N_2275,N_578,N_725);
or U2276 (N_2276,N_423,N_742);
xnor U2277 (N_2277,N_160,N_1033);
or U2278 (N_2278,N_355,N_290);
and U2279 (N_2279,N_629,N_1149);
or U2280 (N_2280,N_27,N_475);
or U2281 (N_2281,N_681,N_726);
and U2282 (N_2282,N_1065,N_1105);
nand U2283 (N_2283,N_473,N_710);
nor U2284 (N_2284,N_1049,N_567);
and U2285 (N_2285,N_1118,N_973);
xnor U2286 (N_2286,N_135,N_732);
nand U2287 (N_2287,N_392,N_1134);
nand U2288 (N_2288,N_242,N_46);
nand U2289 (N_2289,N_463,N_108);
nor U2290 (N_2290,N_805,N_989);
nand U2291 (N_2291,N_566,N_299);
nor U2292 (N_2292,N_997,N_1043);
nor U2293 (N_2293,N_1173,N_1122);
nor U2294 (N_2294,N_150,N_538);
and U2295 (N_2295,N_1244,N_811);
and U2296 (N_2296,N_701,N_615);
nand U2297 (N_2297,N_131,N_896);
nand U2298 (N_2298,N_683,N_1188);
or U2299 (N_2299,N_925,N_1116);
or U2300 (N_2300,N_773,N_534);
nand U2301 (N_2301,N_407,N_1020);
xnor U2302 (N_2302,N_930,N_1224);
nor U2303 (N_2303,N_98,N_876);
xnor U2304 (N_2304,N_321,N_1004);
nand U2305 (N_2305,N_141,N_746);
nor U2306 (N_2306,N_1060,N_1220);
and U2307 (N_2307,N_892,N_1147);
and U2308 (N_2308,N_1200,N_1146);
nor U2309 (N_2309,N_732,N_1225);
or U2310 (N_2310,N_485,N_441);
xnor U2311 (N_2311,N_90,N_1177);
or U2312 (N_2312,N_465,N_1010);
or U2313 (N_2313,N_328,N_537);
or U2314 (N_2314,N_751,N_397);
nor U2315 (N_2315,N_669,N_88);
nand U2316 (N_2316,N_211,N_312);
xnor U2317 (N_2317,N_1117,N_111);
nor U2318 (N_2318,N_220,N_839);
and U2319 (N_2319,N_341,N_1121);
xor U2320 (N_2320,N_1142,N_1234);
nor U2321 (N_2321,N_898,N_427);
nor U2322 (N_2322,N_117,N_136);
xor U2323 (N_2323,N_35,N_258);
and U2324 (N_2324,N_673,N_45);
or U2325 (N_2325,N_1091,N_409);
xor U2326 (N_2326,N_197,N_683);
or U2327 (N_2327,N_1208,N_1144);
xor U2328 (N_2328,N_654,N_937);
xor U2329 (N_2329,N_631,N_483);
xnor U2330 (N_2330,N_908,N_120);
nand U2331 (N_2331,N_1246,N_1156);
or U2332 (N_2332,N_663,N_687);
or U2333 (N_2333,N_481,N_1148);
or U2334 (N_2334,N_1205,N_1007);
xor U2335 (N_2335,N_95,N_640);
and U2336 (N_2336,N_941,N_165);
or U2337 (N_2337,N_522,N_520);
or U2338 (N_2338,N_835,N_201);
xor U2339 (N_2339,N_924,N_463);
nand U2340 (N_2340,N_1237,N_476);
and U2341 (N_2341,N_1006,N_963);
nand U2342 (N_2342,N_362,N_465);
nand U2343 (N_2343,N_789,N_308);
nor U2344 (N_2344,N_741,N_528);
and U2345 (N_2345,N_1228,N_1077);
or U2346 (N_2346,N_396,N_362);
nor U2347 (N_2347,N_1146,N_338);
xnor U2348 (N_2348,N_366,N_526);
or U2349 (N_2349,N_1214,N_551);
xnor U2350 (N_2350,N_930,N_975);
or U2351 (N_2351,N_362,N_508);
xor U2352 (N_2352,N_479,N_439);
xnor U2353 (N_2353,N_1185,N_1167);
or U2354 (N_2354,N_1165,N_1024);
and U2355 (N_2355,N_950,N_703);
and U2356 (N_2356,N_517,N_598);
xnor U2357 (N_2357,N_1151,N_514);
nand U2358 (N_2358,N_736,N_824);
and U2359 (N_2359,N_536,N_517);
nor U2360 (N_2360,N_1,N_954);
xnor U2361 (N_2361,N_697,N_1081);
and U2362 (N_2362,N_756,N_351);
nand U2363 (N_2363,N_72,N_1056);
and U2364 (N_2364,N_455,N_767);
nand U2365 (N_2365,N_142,N_766);
nand U2366 (N_2366,N_148,N_695);
nand U2367 (N_2367,N_355,N_254);
nand U2368 (N_2368,N_4,N_1051);
xor U2369 (N_2369,N_1080,N_1163);
and U2370 (N_2370,N_606,N_1015);
or U2371 (N_2371,N_799,N_656);
nand U2372 (N_2372,N_1045,N_546);
nand U2373 (N_2373,N_508,N_643);
nand U2374 (N_2374,N_52,N_806);
nand U2375 (N_2375,N_838,N_1028);
or U2376 (N_2376,N_438,N_975);
or U2377 (N_2377,N_518,N_540);
nand U2378 (N_2378,N_461,N_526);
nor U2379 (N_2379,N_18,N_483);
nand U2380 (N_2380,N_613,N_1001);
nor U2381 (N_2381,N_144,N_833);
nor U2382 (N_2382,N_191,N_834);
or U2383 (N_2383,N_810,N_538);
or U2384 (N_2384,N_918,N_127);
xnor U2385 (N_2385,N_802,N_569);
nor U2386 (N_2386,N_332,N_802);
nor U2387 (N_2387,N_454,N_574);
nand U2388 (N_2388,N_9,N_24);
xor U2389 (N_2389,N_16,N_1135);
or U2390 (N_2390,N_1249,N_534);
or U2391 (N_2391,N_145,N_74);
or U2392 (N_2392,N_643,N_584);
nor U2393 (N_2393,N_76,N_736);
or U2394 (N_2394,N_677,N_452);
nor U2395 (N_2395,N_906,N_87);
nand U2396 (N_2396,N_566,N_589);
or U2397 (N_2397,N_665,N_1150);
xor U2398 (N_2398,N_965,N_469);
and U2399 (N_2399,N_667,N_304);
xnor U2400 (N_2400,N_752,N_310);
xnor U2401 (N_2401,N_602,N_135);
nor U2402 (N_2402,N_763,N_619);
or U2403 (N_2403,N_759,N_582);
nor U2404 (N_2404,N_687,N_261);
and U2405 (N_2405,N_429,N_518);
or U2406 (N_2406,N_697,N_991);
nand U2407 (N_2407,N_798,N_613);
xnor U2408 (N_2408,N_888,N_1063);
nor U2409 (N_2409,N_1174,N_1003);
xnor U2410 (N_2410,N_851,N_237);
nor U2411 (N_2411,N_943,N_753);
nor U2412 (N_2412,N_33,N_922);
or U2413 (N_2413,N_942,N_0);
nor U2414 (N_2414,N_678,N_95);
xnor U2415 (N_2415,N_1047,N_550);
nor U2416 (N_2416,N_819,N_488);
xnor U2417 (N_2417,N_127,N_1073);
xnor U2418 (N_2418,N_896,N_644);
and U2419 (N_2419,N_331,N_1165);
or U2420 (N_2420,N_1133,N_373);
xor U2421 (N_2421,N_714,N_238);
xnor U2422 (N_2422,N_277,N_1210);
and U2423 (N_2423,N_566,N_6);
and U2424 (N_2424,N_51,N_75);
nand U2425 (N_2425,N_1138,N_730);
nor U2426 (N_2426,N_943,N_55);
nor U2427 (N_2427,N_338,N_1192);
nand U2428 (N_2428,N_1003,N_1054);
nor U2429 (N_2429,N_926,N_789);
and U2430 (N_2430,N_595,N_1233);
xor U2431 (N_2431,N_396,N_1068);
xor U2432 (N_2432,N_817,N_342);
nand U2433 (N_2433,N_409,N_596);
or U2434 (N_2434,N_335,N_346);
and U2435 (N_2435,N_464,N_1167);
nand U2436 (N_2436,N_109,N_587);
nor U2437 (N_2437,N_1158,N_601);
nor U2438 (N_2438,N_770,N_22);
nor U2439 (N_2439,N_205,N_961);
and U2440 (N_2440,N_342,N_807);
nand U2441 (N_2441,N_582,N_1168);
nand U2442 (N_2442,N_155,N_974);
or U2443 (N_2443,N_79,N_48);
nor U2444 (N_2444,N_151,N_747);
or U2445 (N_2445,N_432,N_1030);
nor U2446 (N_2446,N_94,N_805);
xnor U2447 (N_2447,N_1087,N_900);
or U2448 (N_2448,N_442,N_839);
or U2449 (N_2449,N_574,N_989);
and U2450 (N_2450,N_524,N_604);
nand U2451 (N_2451,N_1085,N_246);
nor U2452 (N_2452,N_170,N_334);
xor U2453 (N_2453,N_1185,N_963);
or U2454 (N_2454,N_167,N_247);
or U2455 (N_2455,N_67,N_211);
nor U2456 (N_2456,N_861,N_707);
xnor U2457 (N_2457,N_845,N_602);
nand U2458 (N_2458,N_272,N_876);
and U2459 (N_2459,N_1076,N_1080);
nor U2460 (N_2460,N_617,N_749);
xor U2461 (N_2461,N_999,N_871);
nor U2462 (N_2462,N_1181,N_925);
nor U2463 (N_2463,N_409,N_223);
nor U2464 (N_2464,N_208,N_1010);
xnor U2465 (N_2465,N_7,N_1153);
nor U2466 (N_2466,N_1142,N_439);
and U2467 (N_2467,N_1225,N_731);
and U2468 (N_2468,N_474,N_249);
or U2469 (N_2469,N_1224,N_786);
and U2470 (N_2470,N_1139,N_104);
xor U2471 (N_2471,N_545,N_500);
xor U2472 (N_2472,N_1173,N_718);
xnor U2473 (N_2473,N_886,N_1140);
or U2474 (N_2474,N_794,N_456);
or U2475 (N_2475,N_14,N_599);
nor U2476 (N_2476,N_678,N_463);
or U2477 (N_2477,N_1034,N_784);
and U2478 (N_2478,N_307,N_498);
xnor U2479 (N_2479,N_702,N_358);
or U2480 (N_2480,N_87,N_1144);
and U2481 (N_2481,N_450,N_321);
nand U2482 (N_2482,N_357,N_311);
nand U2483 (N_2483,N_330,N_321);
and U2484 (N_2484,N_1153,N_1033);
xnor U2485 (N_2485,N_625,N_962);
or U2486 (N_2486,N_342,N_228);
or U2487 (N_2487,N_162,N_1167);
or U2488 (N_2488,N_899,N_803);
xor U2489 (N_2489,N_334,N_933);
or U2490 (N_2490,N_353,N_545);
xnor U2491 (N_2491,N_221,N_1149);
or U2492 (N_2492,N_796,N_476);
or U2493 (N_2493,N_26,N_786);
xor U2494 (N_2494,N_815,N_1204);
and U2495 (N_2495,N_1204,N_252);
or U2496 (N_2496,N_88,N_481);
nor U2497 (N_2497,N_1034,N_1126);
nor U2498 (N_2498,N_1243,N_7);
and U2499 (N_2499,N_521,N_221);
nor U2500 (N_2500,N_1855,N_1785);
and U2501 (N_2501,N_2379,N_2117);
xnor U2502 (N_2502,N_2472,N_2374);
and U2503 (N_2503,N_1517,N_1511);
nor U2504 (N_2504,N_1360,N_1483);
or U2505 (N_2505,N_2191,N_1663);
nor U2506 (N_2506,N_1425,N_2344);
nand U2507 (N_2507,N_1709,N_1794);
nand U2508 (N_2508,N_1610,N_1253);
or U2509 (N_2509,N_2373,N_1767);
xor U2510 (N_2510,N_1916,N_2488);
and U2511 (N_2511,N_1318,N_2314);
and U2512 (N_2512,N_2293,N_1774);
nor U2513 (N_2513,N_2402,N_1591);
nor U2514 (N_2514,N_2080,N_1841);
and U2515 (N_2515,N_1309,N_1843);
nor U2516 (N_2516,N_2031,N_1941);
nand U2517 (N_2517,N_1702,N_2214);
or U2518 (N_2518,N_2490,N_1406);
xnor U2519 (N_2519,N_1633,N_1716);
xnor U2520 (N_2520,N_1739,N_2285);
or U2521 (N_2521,N_1395,N_1749);
xor U2522 (N_2522,N_1825,N_2381);
xor U2523 (N_2523,N_2494,N_1305);
nor U2524 (N_2524,N_1846,N_1993);
or U2525 (N_2525,N_1355,N_1526);
xnor U2526 (N_2526,N_1752,N_1891);
xnor U2527 (N_2527,N_1530,N_2283);
and U2528 (N_2528,N_1604,N_2102);
nand U2529 (N_2529,N_2231,N_1995);
nor U2530 (N_2530,N_2313,N_2245);
nor U2531 (N_2531,N_1452,N_1595);
or U2532 (N_2532,N_1903,N_1271);
or U2533 (N_2533,N_1975,N_1555);
xor U2534 (N_2534,N_1323,N_2225);
or U2535 (N_2535,N_1438,N_1945);
or U2536 (N_2536,N_1850,N_1736);
nor U2537 (N_2537,N_1650,N_1653);
nor U2538 (N_2538,N_1811,N_2240);
xnor U2539 (N_2539,N_1701,N_1347);
and U2540 (N_2540,N_2461,N_2474);
xor U2541 (N_2541,N_1434,N_1432);
nor U2542 (N_2542,N_1992,N_1464);
xnor U2543 (N_2543,N_1605,N_2452);
and U2544 (N_2544,N_2052,N_1853);
xnor U2545 (N_2545,N_2294,N_1598);
or U2546 (N_2546,N_1957,N_1881);
xor U2547 (N_2547,N_1491,N_2471);
nand U2548 (N_2548,N_1256,N_1343);
nand U2549 (N_2549,N_1870,N_2105);
and U2550 (N_2550,N_2440,N_2441);
or U2551 (N_2551,N_1453,N_2423);
nand U2552 (N_2552,N_1563,N_1553);
and U2553 (N_2553,N_1960,N_2219);
and U2554 (N_2554,N_2264,N_2019);
nor U2555 (N_2555,N_2151,N_2376);
xnor U2556 (N_2556,N_2103,N_1704);
and U2557 (N_2557,N_1475,N_1354);
or U2558 (N_2558,N_1934,N_1978);
xor U2559 (N_2559,N_1759,N_2093);
and U2560 (N_2560,N_2449,N_2384);
nand U2561 (N_2561,N_2224,N_2171);
nor U2562 (N_2562,N_2128,N_1319);
xnor U2563 (N_2563,N_1766,N_1489);
nor U2564 (N_2564,N_1543,N_1775);
or U2565 (N_2565,N_1330,N_1478);
nor U2566 (N_2566,N_1665,N_2489);
and U2567 (N_2567,N_2247,N_1458);
nand U2568 (N_2568,N_1304,N_1872);
and U2569 (N_2569,N_2261,N_2020);
xor U2570 (N_2570,N_2324,N_2496);
nand U2571 (N_2571,N_1500,N_2346);
xnor U2572 (N_2572,N_2182,N_1282);
xor U2573 (N_2573,N_2258,N_2180);
and U2574 (N_2574,N_1910,N_1725);
xor U2575 (N_2575,N_1751,N_2465);
and U2576 (N_2576,N_2246,N_1279);
nand U2577 (N_2577,N_2401,N_1455);
nand U2578 (N_2578,N_1283,N_2140);
and U2579 (N_2579,N_2190,N_1567);
xor U2580 (N_2580,N_1422,N_1302);
xnor U2581 (N_2581,N_2403,N_1721);
nor U2582 (N_2582,N_2329,N_1871);
or U2583 (N_2583,N_2028,N_2322);
nor U2584 (N_2584,N_2234,N_1364);
and U2585 (N_2585,N_1274,N_1376);
nor U2586 (N_2586,N_1621,N_1815);
or U2587 (N_2587,N_1715,N_1833);
and U2588 (N_2588,N_1269,N_2493);
nor U2589 (N_2589,N_1280,N_2162);
and U2590 (N_2590,N_1415,N_1614);
nand U2591 (N_2591,N_1420,N_2364);
xor U2592 (N_2592,N_1680,N_1792);
or U2593 (N_2593,N_2183,N_1454);
and U2594 (N_2594,N_1911,N_2433);
or U2595 (N_2595,N_1669,N_2056);
nor U2596 (N_2596,N_1340,N_1706);
nand U2597 (N_2597,N_2492,N_2318);
and U2598 (N_2598,N_1925,N_2064);
and U2599 (N_2599,N_1533,N_2207);
nand U2600 (N_2600,N_1809,N_1735);
or U2601 (N_2601,N_1803,N_1732);
or U2602 (N_2602,N_2417,N_2091);
and U2603 (N_2603,N_2263,N_1996);
and U2604 (N_2604,N_1814,N_1922);
nand U2605 (N_2605,N_2340,N_1596);
and U2606 (N_2606,N_1450,N_2223);
or U2607 (N_2607,N_1674,N_1399);
and U2608 (N_2608,N_1789,N_1363);
xnor U2609 (N_2609,N_1413,N_2447);
or U2610 (N_2610,N_1700,N_1424);
xor U2611 (N_2611,N_1545,N_1398);
or U2612 (N_2612,N_1566,N_1358);
xnor U2613 (N_2613,N_2455,N_1710);
nor U2614 (N_2614,N_1968,N_2312);
nand U2615 (N_2615,N_2099,N_1310);
nor U2616 (N_2616,N_1394,N_1503);
xor U2617 (N_2617,N_1384,N_1969);
nand U2618 (N_2618,N_2420,N_2309);
or U2619 (N_2619,N_1582,N_2421);
nand U2620 (N_2620,N_1629,N_2107);
nand U2621 (N_2621,N_2173,N_1864);
nand U2622 (N_2622,N_2386,N_2157);
nor U2623 (N_2623,N_2327,N_1991);
or U2624 (N_2624,N_2053,N_2335);
nor U2625 (N_2625,N_2448,N_1559);
and U2626 (N_2626,N_2319,N_1908);
or U2627 (N_2627,N_1535,N_1327);
xor U2628 (N_2628,N_1942,N_2350);
or U2629 (N_2629,N_1324,N_1265);
xor U2630 (N_2630,N_2266,N_1976);
nand U2631 (N_2631,N_1805,N_1416);
nor U2632 (N_2632,N_1860,N_1727);
nor U2633 (N_2633,N_1408,N_1668);
or U2634 (N_2634,N_1959,N_2396);
nor U2635 (N_2635,N_1593,N_1608);
and U2636 (N_2636,N_1769,N_2252);
xor U2637 (N_2637,N_1580,N_2039);
and U2638 (N_2638,N_2229,N_2453);
nand U2639 (N_2639,N_2193,N_1733);
or U2640 (N_2640,N_1463,N_1381);
xnor U2641 (N_2641,N_2242,N_1666);
nand U2642 (N_2642,N_2317,N_1457);
or U2643 (N_2643,N_2291,N_1865);
and U2644 (N_2644,N_2348,N_1760);
xnor U2645 (N_2645,N_2431,N_2085);
nor U2646 (N_2646,N_1504,N_1697);
and U2647 (N_2647,N_2081,N_1400);
nand U2648 (N_2648,N_1849,N_1515);
or U2649 (N_2649,N_2389,N_2210);
nor U2650 (N_2650,N_2426,N_2310);
or U2651 (N_2651,N_1972,N_1869);
xor U2652 (N_2652,N_1722,N_2037);
nand U2653 (N_2653,N_2069,N_1788);
and U2654 (N_2654,N_1612,N_1404);
xor U2655 (N_2655,N_2347,N_2345);
and U2656 (N_2656,N_2259,N_1423);
xor U2657 (N_2657,N_1719,N_1387);
nor U2658 (N_2658,N_2476,N_1365);
and U2659 (N_2659,N_1393,N_1572);
and U2660 (N_2660,N_1795,N_1427);
nor U2661 (N_2661,N_1481,N_2236);
nor U2662 (N_2662,N_1714,N_1606);
or U2663 (N_2663,N_1664,N_2059);
xor U2664 (N_2664,N_1568,N_1800);
xor U2665 (N_2665,N_1461,N_1804);
or U2666 (N_2666,N_1409,N_1748);
and U2667 (N_2667,N_1966,N_1979);
xor U2668 (N_2668,N_1298,N_1963);
or U2669 (N_2669,N_2256,N_2362);
and U2670 (N_2670,N_2213,N_2311);
nand U2671 (N_2671,N_1254,N_1902);
and U2672 (N_2672,N_2485,N_1906);
and U2673 (N_2673,N_1385,N_2330);
nand U2674 (N_2674,N_1484,N_1578);
and U2675 (N_2675,N_1932,N_1962);
and U2676 (N_2676,N_1313,N_1923);
and U2677 (N_2677,N_2238,N_2243);
and U2678 (N_2678,N_1859,N_2170);
nand U2679 (N_2679,N_1885,N_1781);
nor U2680 (N_2680,N_2459,N_2155);
nand U2681 (N_2681,N_1410,N_1471);
nand U2682 (N_2682,N_1635,N_2016);
nand U2683 (N_2683,N_2068,N_1379);
or U2684 (N_2684,N_1625,N_1863);
nor U2685 (N_2685,N_2321,N_1981);
and U2686 (N_2686,N_2147,N_1440);
nor U2687 (N_2687,N_2135,N_1562);
nand U2688 (N_2688,N_1250,N_2209);
and U2689 (N_2689,N_1565,N_1643);
nor U2690 (N_2690,N_1389,N_1758);
xor U2691 (N_2691,N_2363,N_1574);
and U2692 (N_2692,N_2196,N_1514);
and U2693 (N_2693,N_1292,N_1487);
and U2694 (N_2694,N_1361,N_1268);
and U2695 (N_2695,N_1926,N_1971);
nor U2696 (N_2696,N_1301,N_2015);
nor U2697 (N_2697,N_1391,N_1854);
xnor U2698 (N_2698,N_1892,N_1429);
nand U2699 (N_2699,N_1592,N_1787);
or U2700 (N_2700,N_1616,N_1839);
nor U2701 (N_2701,N_1675,N_1777);
nand U2702 (N_2702,N_1488,N_1778);
xor U2703 (N_2703,N_2076,N_1428);
or U2704 (N_2704,N_1449,N_2220);
and U2705 (N_2705,N_1509,N_2048);
xnor U2706 (N_2706,N_2430,N_1480);
xor U2707 (N_2707,N_1636,N_1405);
nand U2708 (N_2708,N_2480,N_2148);
and U2709 (N_2709,N_2400,N_2161);
nor U2710 (N_2710,N_2275,N_1756);
nand U2711 (N_2711,N_2450,N_1289);
and U2712 (N_2712,N_2152,N_1901);
xnor U2713 (N_2713,N_2250,N_2030);
nor U2714 (N_2714,N_1768,N_1829);
and U2715 (N_2715,N_2290,N_1886);
nand U2716 (N_2716,N_1652,N_2111);
and U2717 (N_2717,N_1651,N_1366);
or U2718 (N_2718,N_2467,N_1508);
and U2719 (N_2719,N_1571,N_1920);
or U2720 (N_2720,N_2342,N_2334);
nand U2721 (N_2721,N_2123,N_1861);
and U2722 (N_2722,N_1974,N_1890);
or U2723 (N_2723,N_1492,N_2227);
nor U2724 (N_2724,N_2478,N_2139);
and U2725 (N_2725,N_1741,N_1382);
and U2726 (N_2726,N_1273,N_1842);
nand U2727 (N_2727,N_1808,N_1705);
and U2728 (N_2728,N_2274,N_1466);
xor U2729 (N_2729,N_2088,N_2338);
nand U2730 (N_2730,N_2078,N_2460);
nand U2731 (N_2731,N_1638,N_2253);
or U2732 (N_2732,N_2458,N_1513);
or U2733 (N_2733,N_1816,N_2305);
or U2734 (N_2734,N_2026,N_1634);
nand U2735 (N_2735,N_1882,N_1827);
nand U2736 (N_2736,N_1765,N_1998);
or U2737 (N_2737,N_1950,N_2277);
nor U2738 (N_2738,N_2462,N_1627);
and U2739 (N_2739,N_2415,N_1344);
xnor U2740 (N_2740,N_1388,N_1899);
or U2741 (N_2741,N_2142,N_2058);
or U2742 (N_2742,N_1443,N_1955);
and U2743 (N_2743,N_2042,N_1371);
nand U2744 (N_2744,N_2262,N_2286);
or U2745 (N_2745,N_1600,N_2438);
xnor U2746 (N_2746,N_2289,N_1284);
and U2747 (N_2747,N_1965,N_1505);
and U2748 (N_2748,N_1779,N_1826);
and U2749 (N_2749,N_2257,N_1683);
or U2750 (N_2750,N_2333,N_2370);
xor U2751 (N_2751,N_2216,N_2150);
and U2752 (N_2752,N_2138,N_1335);
xnor U2753 (N_2753,N_1818,N_1356);
nor U2754 (N_2754,N_1985,N_1331);
nand U2755 (N_2755,N_1522,N_1852);
or U2756 (N_2756,N_1496,N_1747);
nor U2757 (N_2757,N_1433,N_2040);
nand U2758 (N_2758,N_1694,N_1460);
xor U2759 (N_2759,N_2475,N_2297);
nand U2760 (N_2760,N_1938,N_1494);
and U2761 (N_2761,N_1677,N_1844);
or U2762 (N_2762,N_2255,N_2372);
or U2763 (N_2763,N_1397,N_1929);
xnor U2764 (N_2764,N_2482,N_1541);
xnor U2765 (N_2765,N_2398,N_2228);
nor U2766 (N_2766,N_1939,N_2116);
xor U2767 (N_2767,N_1332,N_1502);
nor U2768 (N_2768,N_1836,N_2375);
xor U2769 (N_2769,N_1306,N_1609);
nand U2770 (N_2770,N_1927,N_2188);
xnor U2771 (N_2771,N_2385,N_2292);
xnor U2772 (N_2772,N_2034,N_1479);
or U2773 (N_2773,N_2024,N_1984);
or U2774 (N_2774,N_2212,N_1977);
xnor U2775 (N_2775,N_2054,N_1790);
nand U2776 (N_2776,N_1953,N_2197);
or U2777 (N_2777,N_2481,N_1838);
and U2778 (N_2778,N_1924,N_2108);
xor U2779 (N_2779,N_2204,N_2248);
nor U2780 (N_2780,N_1730,N_1556);
xor U2781 (N_2781,N_2172,N_2136);
or U2782 (N_2782,N_2383,N_2442);
nand U2783 (N_2783,N_1898,N_1495);
nand U2784 (N_2784,N_1295,N_2166);
xnor U2785 (N_2785,N_2392,N_2284);
and U2786 (N_2786,N_1615,N_1510);
xor U2787 (N_2787,N_2164,N_1321);
or U2788 (N_2788,N_1696,N_2491);
nand U2789 (N_2789,N_2114,N_2226);
nor U2790 (N_2790,N_1619,N_2413);
xor U2791 (N_2791,N_1290,N_1695);
and U2792 (N_2792,N_1645,N_2023);
nand U2793 (N_2793,N_2466,N_1287);
xor U2794 (N_2794,N_2141,N_1396);
nor U2795 (N_2795,N_1518,N_1252);
nand U2796 (N_2796,N_1447,N_1528);
nand U2797 (N_2797,N_1681,N_1538);
nor U2798 (N_2798,N_1602,N_1678);
or U2799 (N_2799,N_2121,N_2487);
or U2800 (N_2800,N_1742,N_1812);
or U2801 (N_2801,N_1620,N_2267);
and U2802 (N_2802,N_1915,N_1921);
and U2803 (N_2803,N_1329,N_2165);
nand U2804 (N_2804,N_1367,N_1258);
and U2805 (N_2805,N_2143,N_1717);
nor U2806 (N_2806,N_1551,N_1300);
xor U2807 (N_2807,N_2418,N_2445);
nor U2808 (N_2808,N_2288,N_2051);
nand U2809 (N_2809,N_2282,N_1782);
or U2810 (N_2810,N_1499,N_1832);
nor U2811 (N_2811,N_1845,N_1958);
nor U2812 (N_2812,N_1316,N_1703);
xnor U2813 (N_2813,N_2395,N_1868);
or U2814 (N_2814,N_1362,N_1296);
or U2815 (N_2815,N_1904,N_1952);
and U2816 (N_2816,N_1589,N_1470);
and U2817 (N_2817,N_1866,N_2163);
and U2818 (N_2818,N_2167,N_2298);
nor U2819 (N_2819,N_1469,N_2404);
nor U2820 (N_2820,N_2281,N_1877);
or U2821 (N_2821,N_1713,N_1940);
nand U2822 (N_2822,N_1599,N_2178);
nor U2823 (N_2823,N_1293,N_1656);
nor U2824 (N_2824,N_1948,N_1412);
xnor U2825 (N_2825,N_2090,N_1835);
or U2826 (N_2826,N_1577,N_2184);
or U2827 (N_2827,N_1426,N_2195);
and U2828 (N_2828,N_1679,N_2014);
or U2829 (N_2829,N_2013,N_2098);
nand U2830 (N_2830,N_1328,N_1684);
nor U2831 (N_2831,N_1708,N_1506);
or U2832 (N_2832,N_2100,N_1720);
nand U2833 (N_2833,N_1383,N_1334);
nand U2834 (N_2834,N_1806,N_1338);
nand U2835 (N_2835,N_1576,N_2483);
nand U2836 (N_2836,N_1754,N_1848);
xnor U2837 (N_2837,N_1286,N_1264);
or U2838 (N_2838,N_2361,N_1659);
and U2839 (N_2839,N_2230,N_2018);
xor U2840 (N_2840,N_1617,N_1587);
nor U2841 (N_2841,N_1755,N_1688);
and U2842 (N_2842,N_2371,N_2295);
nand U2843 (N_2843,N_1346,N_1558);
or U2844 (N_2844,N_1983,N_1435);
nor U2845 (N_2845,N_2355,N_1607);
nor U2846 (N_2846,N_1847,N_2249);
or U2847 (N_2847,N_1575,N_1820);
and U2848 (N_2848,N_2454,N_2276);
xor U2849 (N_2849,N_2074,N_2301);
xor U2850 (N_2850,N_1990,N_2272);
and U2851 (N_2851,N_2307,N_1445);
nand U2852 (N_2852,N_2429,N_2200);
xnor U2853 (N_2853,N_1626,N_2129);
or U2854 (N_2854,N_2032,N_1879);
or U2855 (N_2855,N_1465,N_2206);
or U2856 (N_2856,N_1639,N_2125);
or U2857 (N_2857,N_1672,N_2235);
and U2858 (N_2858,N_2422,N_2096);
nor U2859 (N_2859,N_2092,N_1307);
and U2860 (N_2860,N_2038,N_1370);
or U2861 (N_2861,N_1707,N_2201);
or U2862 (N_2862,N_1547,N_2194);
nor U2863 (N_2863,N_1737,N_1402);
and U2864 (N_2864,N_1570,N_2222);
xnor U2865 (N_2865,N_1746,N_2145);
or U2866 (N_2866,N_2159,N_1947);
and U2867 (N_2867,N_2001,N_1339);
xor U2868 (N_2868,N_1336,N_1867);
or U2869 (N_2869,N_2218,N_2132);
nand U2870 (N_2870,N_2192,N_1771);
nand U2871 (N_2871,N_1546,N_1676);
or U2872 (N_2872,N_2268,N_2337);
nand U2873 (N_2873,N_2378,N_1851);
nand U2874 (N_2874,N_2470,N_1474);
or U2875 (N_2875,N_1999,N_1647);
or U2876 (N_2876,N_1618,N_2456);
nor U2877 (N_2877,N_1542,N_2414);
nand U2878 (N_2878,N_1997,N_2174);
or U2879 (N_2879,N_2003,N_2046);
xnor U2880 (N_2880,N_2144,N_2241);
nand U2881 (N_2881,N_1776,N_2208);
nand U2882 (N_2882,N_1276,N_2367);
and U2883 (N_2883,N_1482,N_1630);
and U2884 (N_2884,N_1642,N_1351);
nand U2885 (N_2885,N_2359,N_1586);
xnor U2886 (N_2886,N_1623,N_1900);
or U2887 (N_2887,N_1448,N_2017);
nor U2888 (N_2888,N_2067,N_1982);
nand U2889 (N_2889,N_1793,N_2041);
xor U2890 (N_2890,N_1281,N_1887);
nor U2891 (N_2891,N_1581,N_1529);
and U2892 (N_2892,N_1711,N_1521);
nand U2893 (N_2893,N_1931,N_2000);
or U2894 (N_2894,N_1516,N_1686);
or U2895 (N_2895,N_2073,N_1303);
and U2896 (N_2896,N_2412,N_1291);
nor U2897 (N_2897,N_1446,N_1320);
xor U2898 (N_2898,N_2341,N_1909);
nand U2899 (N_2899,N_1439,N_1796);
xor U2900 (N_2900,N_1731,N_1277);
and U2901 (N_2901,N_1342,N_2027);
xor U2902 (N_2902,N_2082,N_1267);
xor U2903 (N_2903,N_1401,N_1540);
nor U2904 (N_2904,N_2377,N_1662);
nand U2905 (N_2905,N_2211,N_1573);
nand U2906 (N_2906,N_1914,N_2233);
nand U2907 (N_2907,N_1956,N_1368);
nor U2908 (N_2908,N_1359,N_2217);
nand U2909 (N_2909,N_1584,N_2387);
nor U2910 (N_2910,N_1831,N_2469);
nand U2911 (N_2911,N_1744,N_1255);
nand U2912 (N_2912,N_2308,N_2036);
nand U2913 (N_2913,N_2432,N_2106);
nor U2914 (N_2914,N_2498,N_2354);
nand U2915 (N_2915,N_2176,N_2179);
nand U2916 (N_2916,N_1729,N_2109);
and U2917 (N_2917,N_1791,N_1403);
or U2918 (N_2918,N_1797,N_1322);
and U2919 (N_2919,N_1692,N_1660);
xor U2920 (N_2920,N_1987,N_1579);
and U2921 (N_2921,N_1810,N_1773);
or U2922 (N_2922,N_1257,N_1476);
xnor U2923 (N_2923,N_1337,N_1821);
or U2924 (N_2924,N_1601,N_1260);
xnor U2925 (N_2925,N_1333,N_2004);
nor U2926 (N_2926,N_1459,N_2203);
xnor U2927 (N_2927,N_2156,N_1745);
nand U2928 (N_2928,N_1341,N_1893);
nand U2929 (N_2929,N_1375,N_1317);
nor U2930 (N_2930,N_1813,N_2468);
or U2931 (N_2931,N_2443,N_1724);
or U2932 (N_2932,N_2060,N_1437);
xor U2933 (N_2933,N_2486,N_1685);
or U2934 (N_2934,N_2444,N_2205);
or U2935 (N_2935,N_2131,N_1726);
xor U2936 (N_2936,N_1928,N_1883);
and U2937 (N_2937,N_1876,N_1554);
or U2938 (N_2938,N_2049,N_2215);
nor U2939 (N_2939,N_1262,N_2065);
xor U2940 (N_2940,N_1691,N_1436);
xnor U2941 (N_2941,N_2437,N_2320);
xor U2942 (N_2942,N_2380,N_1392);
nand U2943 (N_2943,N_1350,N_1858);
xnor U2944 (N_2944,N_2446,N_1780);
xnor U2945 (N_2945,N_2104,N_2010);
nand U2946 (N_2946,N_1520,N_1613);
and U2947 (N_2947,N_1544,N_1661);
nor U2948 (N_2948,N_1986,N_1988);
or U2949 (N_2949,N_1989,N_2405);
nor U2950 (N_2950,N_1856,N_1837);
xnor U2951 (N_2951,N_1251,N_1548);
xnor U2952 (N_2952,N_1822,N_1477);
nand U2953 (N_2953,N_2356,N_1944);
xnor U2954 (N_2954,N_1583,N_2237);
nand U2955 (N_2955,N_1807,N_2025);
or U2956 (N_2956,N_1637,N_1772);
and U2957 (N_2957,N_2113,N_1297);
and U2958 (N_2958,N_1442,N_2279);
xor U2959 (N_2959,N_1456,N_2044);
nor U2960 (N_2960,N_2122,N_2185);
xnor U2961 (N_2961,N_2133,N_1386);
and U2962 (N_2962,N_1912,N_2352);
and U2963 (N_2963,N_1917,N_1897);
nor U2964 (N_2964,N_1486,N_1308);
nand U2965 (N_2965,N_2473,N_1585);
xor U2966 (N_2966,N_2047,N_1698);
and U2967 (N_2967,N_2271,N_2087);
nor U2968 (N_2968,N_1670,N_1930);
or U2969 (N_2969,N_1631,N_2477);
xnor U2970 (N_2970,N_1357,N_2351);
xor U2971 (N_2971,N_2254,N_1764);
and U2972 (N_2972,N_2177,N_2008);
nand U2973 (N_2973,N_2061,N_1873);
nor U2974 (N_2974,N_1770,N_2315);
and U2975 (N_2975,N_2336,N_1561);
nand U2976 (N_2976,N_1641,N_2126);
nor U2977 (N_2977,N_2436,N_1658);
and U2978 (N_2978,N_1430,N_2270);
and U2979 (N_2979,N_2495,N_2484);
and U2980 (N_2980,N_1532,N_2002);
and U2981 (N_2981,N_1786,N_2086);
nor U2982 (N_2982,N_2435,N_1830);
nor U2983 (N_2983,N_1970,N_1933);
nor U2984 (N_2984,N_1840,N_2296);
or U2985 (N_2985,N_1734,N_1946);
and U2986 (N_2986,N_1569,N_1936);
and U2987 (N_2987,N_2045,N_2006);
or U2988 (N_2988,N_2168,N_2110);
and U2989 (N_2989,N_1784,N_1373);
nand U2990 (N_2990,N_1594,N_2300);
nor U2991 (N_2991,N_1654,N_1418);
nor U2992 (N_2992,N_2434,N_1690);
nand U2993 (N_2993,N_1783,N_1951);
xnor U2994 (N_2994,N_1819,N_2382);
nand U2995 (N_2995,N_2075,N_2306);
and U2996 (N_2996,N_1644,N_1539);
nor U2997 (N_2997,N_2451,N_1523);
and U2998 (N_2998,N_2328,N_2186);
xor U2999 (N_2999,N_1728,N_2198);
nand U3000 (N_3000,N_1834,N_2332);
or U3001 (N_3001,N_1564,N_2079);
nor U3002 (N_3002,N_1501,N_1490);
nand U3003 (N_3003,N_2202,N_1549);
nand U3004 (N_3004,N_1473,N_1874);
xnor U3005 (N_3005,N_2033,N_2181);
and U3006 (N_3006,N_2011,N_1875);
or U3007 (N_3007,N_1750,N_2112);
xor U3008 (N_3008,N_2160,N_2084);
and U3009 (N_3009,N_1468,N_1689);
xor U3010 (N_3010,N_2369,N_1880);
xnor U3011 (N_3011,N_1884,N_1467);
and U3012 (N_3012,N_1693,N_1534);
and U3013 (N_3013,N_2158,N_2497);
xor U3014 (N_3014,N_1285,N_1802);
nand U3015 (N_3015,N_2043,N_2499);
nand U3016 (N_3016,N_1655,N_2119);
nand U3017 (N_3017,N_2457,N_1390);
nor U3018 (N_3018,N_2280,N_2394);
nand U3019 (N_3019,N_2137,N_2353);
or U3020 (N_3020,N_2419,N_1738);
nor U3021 (N_3021,N_2005,N_1524);
nor U3022 (N_3022,N_1753,N_2077);
and U3023 (N_3023,N_1611,N_2463);
nor U3024 (N_3024,N_2304,N_1640);
nor U3025 (N_3025,N_1557,N_1961);
nor U3026 (N_3026,N_2118,N_2428);
and U3027 (N_3027,N_2244,N_1312);
and U3028 (N_3028,N_1272,N_2007);
xnor U3029 (N_3029,N_1314,N_1421);
or U3030 (N_3030,N_1895,N_2349);
or U3031 (N_3031,N_1550,N_2175);
xor U3032 (N_3032,N_2366,N_2303);
and U3033 (N_3033,N_2149,N_2273);
xnor U3034 (N_3034,N_1949,N_2260);
or U3035 (N_3035,N_1414,N_1261);
nand U3036 (N_3036,N_1372,N_1954);
or U3037 (N_3037,N_2302,N_1374);
xnor U3038 (N_3038,N_2391,N_1407);
nand U3039 (N_3039,N_2397,N_2411);
nand U3040 (N_3040,N_1444,N_1943);
and U3041 (N_3041,N_1628,N_1646);
and U3042 (N_3042,N_2055,N_2094);
nor U3043 (N_3043,N_1671,N_2029);
nor U3044 (N_3044,N_1799,N_2406);
nand U3045 (N_3045,N_2278,N_1353);
nor U3046 (N_3046,N_1411,N_1377);
nor U3047 (N_3047,N_1512,N_2360);
xor U3048 (N_3048,N_1973,N_1462);
and U3049 (N_3049,N_1964,N_1485);
nor U3050 (N_3050,N_2127,N_1824);
xnor U3051 (N_3051,N_1419,N_2479);
nand U3052 (N_3052,N_1657,N_1649);
nor U3053 (N_3053,N_2022,N_1531);
xnor U3054 (N_3054,N_1507,N_2012);
nand U3055 (N_3055,N_2439,N_2101);
nand U3056 (N_3056,N_1537,N_2357);
or U3057 (N_3057,N_2390,N_2189);
nand U3058 (N_3058,N_1889,N_1299);
nor U3059 (N_3059,N_1967,N_1918);
nand U3060 (N_3060,N_2134,N_1560);
or U3061 (N_3061,N_1278,N_1823);
nand U3062 (N_3062,N_2407,N_1525);
nor U3063 (N_3063,N_1682,N_1913);
or U3064 (N_3064,N_2416,N_2325);
nor U3065 (N_3065,N_2187,N_1380);
nor U3066 (N_3066,N_2410,N_1896);
xor U3067 (N_3067,N_2062,N_2057);
nor U3068 (N_3068,N_2331,N_2388);
and U3069 (N_3069,N_1801,N_2070);
nand U3070 (N_3070,N_1743,N_1431);
and U3071 (N_3071,N_1994,N_2124);
or U3072 (N_3072,N_2154,N_1349);
xor U3073 (N_3073,N_1980,N_1937);
nand U3074 (N_3074,N_1687,N_2050);
or U3075 (N_3075,N_2316,N_1378);
xor U3076 (N_3076,N_1259,N_1632);
nand U3077 (N_3077,N_1266,N_2409);
nand U3078 (N_3078,N_2425,N_1315);
nand U3079 (N_3079,N_1498,N_1417);
nand U3080 (N_3080,N_2239,N_2097);
nor U3081 (N_3081,N_1270,N_1590);
nor U3082 (N_3082,N_1862,N_2343);
xor U3083 (N_3083,N_1624,N_1907);
xnor U3084 (N_3084,N_1311,N_2408);
nor U3085 (N_3085,N_1761,N_1763);
or U3086 (N_3086,N_1622,N_1597);
and U3087 (N_3087,N_1326,N_2130);
nor U3088 (N_3088,N_2063,N_2083);
and U3089 (N_3089,N_1648,N_2251);
xor U3090 (N_3090,N_1798,N_2399);
nand U3091 (N_3091,N_2232,N_2221);
and U3092 (N_3092,N_2095,N_1588);
or U3093 (N_3093,N_2146,N_1288);
or U3094 (N_3094,N_2424,N_2464);
xnor U3095 (N_3095,N_2021,N_1493);
and U3096 (N_3096,N_1828,N_1905);
nor U3097 (N_3097,N_2009,N_1536);
nor U3098 (N_3098,N_1919,N_2339);
or U3099 (N_3099,N_1935,N_1472);
nand U3100 (N_3100,N_1740,N_1552);
xnor U3101 (N_3101,N_1817,N_1369);
nor U3102 (N_3102,N_1894,N_2071);
and U3103 (N_3103,N_1527,N_2153);
xor U3104 (N_3104,N_1699,N_1667);
nand U3105 (N_3105,N_2299,N_2326);
and U3106 (N_3106,N_1352,N_1263);
nand U3107 (N_3107,N_2365,N_2393);
xnor U3108 (N_3108,N_1497,N_2368);
or U3109 (N_3109,N_2358,N_1451);
or U3110 (N_3110,N_2427,N_2120);
nand U3111 (N_3111,N_2265,N_2269);
nor U3112 (N_3112,N_1294,N_1348);
xnor U3113 (N_3113,N_1441,N_1519);
and U3114 (N_3114,N_1718,N_1325);
nand U3115 (N_3115,N_2072,N_1888);
nor U3116 (N_3116,N_2089,N_1723);
nand U3117 (N_3117,N_2199,N_2115);
and U3118 (N_3118,N_1603,N_1762);
nor U3119 (N_3119,N_1673,N_2323);
or U3120 (N_3120,N_1275,N_1857);
xor U3121 (N_3121,N_2169,N_1757);
xnor U3122 (N_3122,N_1712,N_2035);
nor U3123 (N_3123,N_2066,N_1878);
nand U3124 (N_3124,N_1345,N_2287);
or U3125 (N_3125,N_1484,N_1400);
xor U3126 (N_3126,N_1449,N_2395);
or U3127 (N_3127,N_1321,N_1947);
nand U3128 (N_3128,N_1558,N_1815);
and U3129 (N_3129,N_2304,N_2250);
or U3130 (N_3130,N_2160,N_1376);
nor U3131 (N_3131,N_1662,N_1381);
and U3132 (N_3132,N_1489,N_2393);
and U3133 (N_3133,N_1596,N_1962);
xor U3134 (N_3134,N_1770,N_1861);
or U3135 (N_3135,N_2179,N_1827);
xor U3136 (N_3136,N_1867,N_1475);
or U3137 (N_3137,N_1475,N_1486);
xnor U3138 (N_3138,N_2443,N_1733);
xor U3139 (N_3139,N_1378,N_2222);
xnor U3140 (N_3140,N_1901,N_1959);
nand U3141 (N_3141,N_2114,N_2070);
xnor U3142 (N_3142,N_1741,N_1381);
or U3143 (N_3143,N_1376,N_2085);
and U3144 (N_3144,N_2115,N_2172);
or U3145 (N_3145,N_1758,N_2243);
or U3146 (N_3146,N_2176,N_1394);
xnor U3147 (N_3147,N_1381,N_1435);
and U3148 (N_3148,N_1762,N_2183);
xor U3149 (N_3149,N_2398,N_1796);
nand U3150 (N_3150,N_2338,N_2154);
nand U3151 (N_3151,N_1959,N_1691);
nor U3152 (N_3152,N_1500,N_2252);
or U3153 (N_3153,N_1514,N_2135);
and U3154 (N_3154,N_2236,N_1362);
or U3155 (N_3155,N_1346,N_1426);
nor U3156 (N_3156,N_2372,N_1578);
and U3157 (N_3157,N_2230,N_1568);
nor U3158 (N_3158,N_1634,N_1358);
or U3159 (N_3159,N_1861,N_1884);
nor U3160 (N_3160,N_2482,N_2403);
nand U3161 (N_3161,N_2496,N_1585);
nand U3162 (N_3162,N_1969,N_1675);
and U3163 (N_3163,N_1295,N_2398);
nand U3164 (N_3164,N_2297,N_1915);
nand U3165 (N_3165,N_1799,N_1431);
and U3166 (N_3166,N_1636,N_2344);
nor U3167 (N_3167,N_1874,N_1405);
or U3168 (N_3168,N_2423,N_1278);
nor U3169 (N_3169,N_1768,N_1423);
xnor U3170 (N_3170,N_1730,N_1851);
nand U3171 (N_3171,N_2028,N_1362);
and U3172 (N_3172,N_2391,N_1434);
nor U3173 (N_3173,N_2337,N_1254);
and U3174 (N_3174,N_1264,N_1629);
or U3175 (N_3175,N_1702,N_2286);
and U3176 (N_3176,N_1350,N_2416);
nand U3177 (N_3177,N_1644,N_2292);
or U3178 (N_3178,N_1280,N_1730);
nand U3179 (N_3179,N_2006,N_1768);
xor U3180 (N_3180,N_2151,N_2388);
and U3181 (N_3181,N_2150,N_2302);
nand U3182 (N_3182,N_2218,N_1863);
and U3183 (N_3183,N_1497,N_2181);
or U3184 (N_3184,N_1349,N_2435);
nor U3185 (N_3185,N_2077,N_1335);
and U3186 (N_3186,N_1642,N_2016);
xnor U3187 (N_3187,N_1707,N_1313);
and U3188 (N_3188,N_1449,N_1828);
xnor U3189 (N_3189,N_1845,N_1734);
or U3190 (N_3190,N_1272,N_1498);
and U3191 (N_3191,N_1880,N_2167);
xor U3192 (N_3192,N_1684,N_2257);
and U3193 (N_3193,N_1361,N_2325);
or U3194 (N_3194,N_1465,N_2190);
and U3195 (N_3195,N_1548,N_2175);
and U3196 (N_3196,N_1397,N_2477);
nand U3197 (N_3197,N_2498,N_2241);
and U3198 (N_3198,N_1335,N_1869);
nor U3199 (N_3199,N_2144,N_1835);
nor U3200 (N_3200,N_1334,N_1910);
xor U3201 (N_3201,N_1310,N_1977);
xnor U3202 (N_3202,N_2264,N_1277);
nand U3203 (N_3203,N_1617,N_2394);
or U3204 (N_3204,N_1312,N_1804);
and U3205 (N_3205,N_1800,N_2147);
nand U3206 (N_3206,N_2225,N_1470);
nor U3207 (N_3207,N_2374,N_2018);
xnor U3208 (N_3208,N_1889,N_1435);
and U3209 (N_3209,N_1525,N_2358);
xnor U3210 (N_3210,N_1654,N_2389);
xnor U3211 (N_3211,N_1279,N_2482);
or U3212 (N_3212,N_2252,N_2257);
nand U3213 (N_3213,N_1442,N_1969);
nor U3214 (N_3214,N_2390,N_1565);
nor U3215 (N_3215,N_2255,N_1683);
and U3216 (N_3216,N_1855,N_1668);
xnor U3217 (N_3217,N_2024,N_2369);
xor U3218 (N_3218,N_2390,N_1436);
or U3219 (N_3219,N_2458,N_2354);
or U3220 (N_3220,N_2433,N_1536);
and U3221 (N_3221,N_1843,N_2072);
nand U3222 (N_3222,N_1917,N_1250);
nand U3223 (N_3223,N_2196,N_1836);
or U3224 (N_3224,N_2025,N_2138);
nand U3225 (N_3225,N_1796,N_2057);
nand U3226 (N_3226,N_2172,N_1705);
and U3227 (N_3227,N_2080,N_1781);
or U3228 (N_3228,N_2055,N_1455);
nor U3229 (N_3229,N_1259,N_2433);
nor U3230 (N_3230,N_2431,N_2121);
and U3231 (N_3231,N_1794,N_1798);
and U3232 (N_3232,N_1970,N_1376);
nand U3233 (N_3233,N_2183,N_1890);
or U3234 (N_3234,N_1686,N_1736);
nand U3235 (N_3235,N_1529,N_2356);
nand U3236 (N_3236,N_2127,N_1859);
and U3237 (N_3237,N_1872,N_1311);
xnor U3238 (N_3238,N_2316,N_1444);
or U3239 (N_3239,N_2470,N_1320);
or U3240 (N_3240,N_2216,N_2265);
nand U3241 (N_3241,N_2475,N_1386);
nor U3242 (N_3242,N_2170,N_2182);
and U3243 (N_3243,N_2206,N_1973);
xnor U3244 (N_3244,N_1372,N_1370);
xnor U3245 (N_3245,N_2226,N_2166);
and U3246 (N_3246,N_1949,N_1868);
and U3247 (N_3247,N_2095,N_1320);
and U3248 (N_3248,N_2028,N_1907);
xnor U3249 (N_3249,N_1635,N_1337);
and U3250 (N_3250,N_2127,N_2464);
and U3251 (N_3251,N_1916,N_1328);
nand U3252 (N_3252,N_1992,N_1539);
nand U3253 (N_3253,N_1859,N_2058);
nand U3254 (N_3254,N_2096,N_2209);
nor U3255 (N_3255,N_2352,N_1712);
or U3256 (N_3256,N_2089,N_1853);
nand U3257 (N_3257,N_1770,N_2483);
xnor U3258 (N_3258,N_1411,N_2173);
nor U3259 (N_3259,N_2047,N_2421);
and U3260 (N_3260,N_2306,N_2482);
nor U3261 (N_3261,N_2157,N_2056);
xor U3262 (N_3262,N_1725,N_2342);
and U3263 (N_3263,N_2377,N_1845);
and U3264 (N_3264,N_1677,N_2236);
xnor U3265 (N_3265,N_2233,N_1707);
xor U3266 (N_3266,N_1286,N_2268);
and U3267 (N_3267,N_1250,N_2122);
nand U3268 (N_3268,N_1291,N_1826);
or U3269 (N_3269,N_1357,N_1773);
or U3270 (N_3270,N_1472,N_2167);
nand U3271 (N_3271,N_2154,N_2353);
nand U3272 (N_3272,N_2167,N_1915);
nand U3273 (N_3273,N_1971,N_2490);
and U3274 (N_3274,N_1409,N_1922);
and U3275 (N_3275,N_1393,N_2142);
or U3276 (N_3276,N_1896,N_2499);
and U3277 (N_3277,N_1546,N_1881);
or U3278 (N_3278,N_1365,N_1345);
and U3279 (N_3279,N_1960,N_1475);
nand U3280 (N_3280,N_2451,N_1781);
and U3281 (N_3281,N_2325,N_1883);
xnor U3282 (N_3282,N_2367,N_2056);
or U3283 (N_3283,N_2259,N_1967);
and U3284 (N_3284,N_1578,N_2408);
nor U3285 (N_3285,N_2000,N_1776);
or U3286 (N_3286,N_2452,N_2036);
nor U3287 (N_3287,N_1706,N_2318);
or U3288 (N_3288,N_1416,N_1445);
nand U3289 (N_3289,N_1917,N_2084);
xor U3290 (N_3290,N_1909,N_1887);
nand U3291 (N_3291,N_1287,N_1443);
nand U3292 (N_3292,N_2271,N_1339);
nand U3293 (N_3293,N_1455,N_2299);
and U3294 (N_3294,N_2455,N_2062);
or U3295 (N_3295,N_2026,N_2408);
and U3296 (N_3296,N_2266,N_2204);
xor U3297 (N_3297,N_2084,N_1887);
and U3298 (N_3298,N_1351,N_1982);
xor U3299 (N_3299,N_2182,N_1945);
or U3300 (N_3300,N_1545,N_1733);
xor U3301 (N_3301,N_1320,N_2119);
nor U3302 (N_3302,N_1618,N_1409);
and U3303 (N_3303,N_2012,N_1436);
nand U3304 (N_3304,N_1386,N_2432);
and U3305 (N_3305,N_1996,N_1309);
nand U3306 (N_3306,N_1543,N_1386);
nor U3307 (N_3307,N_1363,N_1407);
nand U3308 (N_3308,N_1322,N_2110);
nand U3309 (N_3309,N_1791,N_1822);
or U3310 (N_3310,N_2165,N_1536);
and U3311 (N_3311,N_1355,N_1574);
xor U3312 (N_3312,N_1625,N_1288);
xnor U3313 (N_3313,N_1964,N_1472);
nand U3314 (N_3314,N_1336,N_1271);
or U3315 (N_3315,N_1953,N_1272);
xnor U3316 (N_3316,N_2030,N_2115);
xnor U3317 (N_3317,N_2333,N_2253);
nand U3318 (N_3318,N_1325,N_2115);
xnor U3319 (N_3319,N_2276,N_1635);
or U3320 (N_3320,N_1792,N_1979);
nand U3321 (N_3321,N_2086,N_1971);
nand U3322 (N_3322,N_1926,N_2099);
xnor U3323 (N_3323,N_2366,N_1669);
or U3324 (N_3324,N_2141,N_2110);
or U3325 (N_3325,N_1718,N_2067);
or U3326 (N_3326,N_1410,N_1297);
or U3327 (N_3327,N_1499,N_1795);
and U3328 (N_3328,N_1489,N_1604);
and U3329 (N_3329,N_1483,N_1288);
or U3330 (N_3330,N_1442,N_1759);
or U3331 (N_3331,N_1558,N_1838);
nor U3332 (N_3332,N_1254,N_1298);
or U3333 (N_3333,N_1746,N_1895);
or U3334 (N_3334,N_1905,N_1683);
or U3335 (N_3335,N_1792,N_2219);
xor U3336 (N_3336,N_1369,N_1720);
nand U3337 (N_3337,N_1640,N_1551);
or U3338 (N_3338,N_2496,N_1776);
or U3339 (N_3339,N_2374,N_2492);
or U3340 (N_3340,N_2017,N_2492);
nand U3341 (N_3341,N_2308,N_1439);
or U3342 (N_3342,N_1454,N_2175);
xor U3343 (N_3343,N_1806,N_2362);
nand U3344 (N_3344,N_2237,N_1866);
and U3345 (N_3345,N_2165,N_1603);
xnor U3346 (N_3346,N_1795,N_1679);
or U3347 (N_3347,N_1347,N_1737);
nand U3348 (N_3348,N_1358,N_2241);
nor U3349 (N_3349,N_2406,N_2337);
and U3350 (N_3350,N_2268,N_1273);
xor U3351 (N_3351,N_2158,N_2216);
xnor U3352 (N_3352,N_2391,N_1910);
xor U3353 (N_3353,N_1725,N_2025);
xnor U3354 (N_3354,N_1327,N_1497);
nor U3355 (N_3355,N_2336,N_1844);
xor U3356 (N_3356,N_1939,N_2337);
or U3357 (N_3357,N_2169,N_1452);
nor U3358 (N_3358,N_1572,N_2455);
xnor U3359 (N_3359,N_2382,N_1545);
nor U3360 (N_3360,N_2130,N_1481);
and U3361 (N_3361,N_1549,N_2349);
or U3362 (N_3362,N_1802,N_2248);
nand U3363 (N_3363,N_1537,N_1430);
nand U3364 (N_3364,N_1906,N_1929);
and U3365 (N_3365,N_2471,N_2187);
and U3366 (N_3366,N_1318,N_1271);
xor U3367 (N_3367,N_1385,N_2011);
or U3368 (N_3368,N_2391,N_2297);
nand U3369 (N_3369,N_1392,N_2021);
or U3370 (N_3370,N_1263,N_1711);
nand U3371 (N_3371,N_2388,N_1784);
and U3372 (N_3372,N_1723,N_2328);
nor U3373 (N_3373,N_1591,N_2111);
and U3374 (N_3374,N_2389,N_1274);
xor U3375 (N_3375,N_2448,N_1514);
and U3376 (N_3376,N_1675,N_1435);
nor U3377 (N_3377,N_1716,N_2068);
nand U3378 (N_3378,N_1544,N_1321);
nand U3379 (N_3379,N_1378,N_2256);
and U3380 (N_3380,N_1533,N_1495);
and U3381 (N_3381,N_2495,N_1903);
nand U3382 (N_3382,N_2274,N_1971);
xor U3383 (N_3383,N_2436,N_1289);
or U3384 (N_3384,N_1654,N_1517);
nand U3385 (N_3385,N_2025,N_2348);
or U3386 (N_3386,N_2267,N_2160);
nor U3387 (N_3387,N_2230,N_1391);
or U3388 (N_3388,N_1776,N_1701);
nand U3389 (N_3389,N_1391,N_2034);
and U3390 (N_3390,N_1626,N_1639);
and U3391 (N_3391,N_2253,N_2318);
xnor U3392 (N_3392,N_1523,N_1777);
nor U3393 (N_3393,N_1973,N_2375);
and U3394 (N_3394,N_1546,N_2483);
or U3395 (N_3395,N_2397,N_2178);
xor U3396 (N_3396,N_2301,N_1840);
nor U3397 (N_3397,N_2225,N_1465);
xor U3398 (N_3398,N_2056,N_1801);
xnor U3399 (N_3399,N_2492,N_2048);
and U3400 (N_3400,N_1773,N_1826);
xor U3401 (N_3401,N_1415,N_2436);
and U3402 (N_3402,N_2395,N_1250);
xnor U3403 (N_3403,N_1785,N_2126);
nor U3404 (N_3404,N_2365,N_2267);
xnor U3405 (N_3405,N_1793,N_2399);
or U3406 (N_3406,N_2363,N_2459);
nand U3407 (N_3407,N_1515,N_1348);
nand U3408 (N_3408,N_1256,N_1832);
nor U3409 (N_3409,N_1407,N_1787);
and U3410 (N_3410,N_2340,N_1602);
nor U3411 (N_3411,N_2308,N_1679);
nor U3412 (N_3412,N_2152,N_2011);
or U3413 (N_3413,N_1465,N_1609);
xor U3414 (N_3414,N_1288,N_2168);
and U3415 (N_3415,N_1255,N_1736);
and U3416 (N_3416,N_2356,N_1784);
nor U3417 (N_3417,N_1623,N_2075);
and U3418 (N_3418,N_2256,N_1799);
and U3419 (N_3419,N_1391,N_1386);
and U3420 (N_3420,N_1611,N_1752);
and U3421 (N_3421,N_2207,N_2153);
nor U3422 (N_3422,N_1581,N_1903);
xnor U3423 (N_3423,N_1549,N_2341);
xnor U3424 (N_3424,N_1251,N_2098);
nor U3425 (N_3425,N_2427,N_2251);
xor U3426 (N_3426,N_1559,N_2018);
nand U3427 (N_3427,N_1404,N_2097);
nor U3428 (N_3428,N_2281,N_1660);
nand U3429 (N_3429,N_1744,N_1601);
and U3430 (N_3430,N_2433,N_2052);
and U3431 (N_3431,N_1475,N_2156);
or U3432 (N_3432,N_2291,N_1874);
and U3433 (N_3433,N_2251,N_1871);
nand U3434 (N_3434,N_1913,N_1348);
xor U3435 (N_3435,N_1472,N_1990);
or U3436 (N_3436,N_2159,N_1461);
nor U3437 (N_3437,N_1522,N_1998);
or U3438 (N_3438,N_1323,N_2263);
nand U3439 (N_3439,N_2336,N_1934);
nor U3440 (N_3440,N_1935,N_2440);
or U3441 (N_3441,N_1363,N_1272);
and U3442 (N_3442,N_1568,N_1706);
xor U3443 (N_3443,N_1740,N_1367);
or U3444 (N_3444,N_2393,N_1801);
and U3445 (N_3445,N_1312,N_1943);
and U3446 (N_3446,N_2481,N_2059);
or U3447 (N_3447,N_1256,N_1488);
nand U3448 (N_3448,N_1850,N_2291);
or U3449 (N_3449,N_1624,N_1544);
or U3450 (N_3450,N_2044,N_1709);
nand U3451 (N_3451,N_1583,N_2364);
nor U3452 (N_3452,N_2135,N_1841);
xnor U3453 (N_3453,N_1612,N_1300);
or U3454 (N_3454,N_1853,N_2175);
nor U3455 (N_3455,N_2169,N_2278);
or U3456 (N_3456,N_2062,N_2476);
xnor U3457 (N_3457,N_1393,N_2235);
xnor U3458 (N_3458,N_1822,N_2325);
xor U3459 (N_3459,N_2497,N_1732);
nand U3460 (N_3460,N_1823,N_2039);
nand U3461 (N_3461,N_2377,N_2160);
nand U3462 (N_3462,N_2336,N_2090);
nand U3463 (N_3463,N_2336,N_1890);
nand U3464 (N_3464,N_2104,N_2149);
or U3465 (N_3465,N_2185,N_1966);
nor U3466 (N_3466,N_2243,N_1693);
and U3467 (N_3467,N_2434,N_1502);
xor U3468 (N_3468,N_1755,N_1645);
nand U3469 (N_3469,N_2245,N_2082);
or U3470 (N_3470,N_2466,N_1447);
nor U3471 (N_3471,N_2276,N_1721);
or U3472 (N_3472,N_2313,N_1876);
and U3473 (N_3473,N_1523,N_1386);
xnor U3474 (N_3474,N_2314,N_1958);
and U3475 (N_3475,N_1886,N_1678);
nand U3476 (N_3476,N_1812,N_1949);
and U3477 (N_3477,N_1848,N_1566);
xor U3478 (N_3478,N_2367,N_2454);
or U3479 (N_3479,N_1457,N_2240);
xnor U3480 (N_3480,N_2371,N_1715);
and U3481 (N_3481,N_1423,N_1822);
nand U3482 (N_3482,N_2413,N_1616);
nand U3483 (N_3483,N_2185,N_1266);
nand U3484 (N_3484,N_1360,N_1293);
xnor U3485 (N_3485,N_1937,N_2147);
or U3486 (N_3486,N_1983,N_2453);
and U3487 (N_3487,N_1317,N_1789);
and U3488 (N_3488,N_1271,N_1527);
nor U3489 (N_3489,N_1947,N_1602);
or U3490 (N_3490,N_1558,N_1751);
and U3491 (N_3491,N_1461,N_2405);
and U3492 (N_3492,N_2058,N_2236);
or U3493 (N_3493,N_2119,N_1665);
nand U3494 (N_3494,N_1738,N_1520);
nor U3495 (N_3495,N_1974,N_1497);
nor U3496 (N_3496,N_1752,N_1608);
nand U3497 (N_3497,N_1884,N_1486);
xnor U3498 (N_3498,N_1862,N_2075);
or U3499 (N_3499,N_2339,N_2192);
nand U3500 (N_3500,N_1601,N_2352);
xnor U3501 (N_3501,N_1718,N_1724);
and U3502 (N_3502,N_2235,N_2425);
and U3503 (N_3503,N_1813,N_1362);
and U3504 (N_3504,N_2385,N_1746);
xnor U3505 (N_3505,N_2391,N_2256);
or U3506 (N_3506,N_2100,N_1972);
or U3507 (N_3507,N_1770,N_1449);
nand U3508 (N_3508,N_1962,N_1973);
or U3509 (N_3509,N_2241,N_2160);
and U3510 (N_3510,N_1959,N_2395);
and U3511 (N_3511,N_1548,N_2174);
and U3512 (N_3512,N_1947,N_2186);
nor U3513 (N_3513,N_1591,N_1693);
and U3514 (N_3514,N_1988,N_2098);
xnor U3515 (N_3515,N_1947,N_2014);
nor U3516 (N_3516,N_2499,N_1800);
nor U3517 (N_3517,N_1705,N_1645);
nand U3518 (N_3518,N_2038,N_2096);
or U3519 (N_3519,N_1985,N_2137);
nor U3520 (N_3520,N_1661,N_2282);
xnor U3521 (N_3521,N_2184,N_1665);
and U3522 (N_3522,N_1390,N_2388);
nand U3523 (N_3523,N_1711,N_1493);
and U3524 (N_3524,N_1765,N_2369);
xnor U3525 (N_3525,N_2290,N_1352);
or U3526 (N_3526,N_2025,N_1767);
or U3527 (N_3527,N_1543,N_1683);
or U3528 (N_3528,N_1308,N_1436);
and U3529 (N_3529,N_2276,N_1290);
xnor U3530 (N_3530,N_1723,N_1394);
and U3531 (N_3531,N_1362,N_2174);
or U3532 (N_3532,N_1443,N_2095);
nand U3533 (N_3533,N_1367,N_1420);
nor U3534 (N_3534,N_2159,N_1842);
xnor U3535 (N_3535,N_1564,N_1395);
or U3536 (N_3536,N_2170,N_1686);
or U3537 (N_3537,N_1286,N_1906);
nand U3538 (N_3538,N_2072,N_2155);
nor U3539 (N_3539,N_1465,N_1513);
xnor U3540 (N_3540,N_1934,N_1724);
nor U3541 (N_3541,N_2046,N_1446);
or U3542 (N_3542,N_1856,N_1340);
and U3543 (N_3543,N_2000,N_2094);
or U3544 (N_3544,N_1762,N_1628);
xor U3545 (N_3545,N_2063,N_2482);
nand U3546 (N_3546,N_1530,N_1276);
nor U3547 (N_3547,N_1485,N_1283);
xnor U3548 (N_3548,N_1865,N_2254);
nor U3549 (N_3549,N_2244,N_1824);
xnor U3550 (N_3550,N_2492,N_1774);
or U3551 (N_3551,N_2406,N_2082);
or U3552 (N_3552,N_1329,N_2456);
and U3553 (N_3553,N_2335,N_2337);
and U3554 (N_3554,N_1600,N_1754);
nand U3555 (N_3555,N_1467,N_2013);
nor U3556 (N_3556,N_1339,N_1524);
and U3557 (N_3557,N_1346,N_2385);
and U3558 (N_3558,N_2027,N_1324);
xor U3559 (N_3559,N_1969,N_2346);
and U3560 (N_3560,N_1795,N_2001);
and U3561 (N_3561,N_1713,N_2080);
or U3562 (N_3562,N_1994,N_2201);
xnor U3563 (N_3563,N_1358,N_2134);
nor U3564 (N_3564,N_1717,N_1344);
nor U3565 (N_3565,N_2279,N_1879);
and U3566 (N_3566,N_1435,N_2014);
or U3567 (N_3567,N_1901,N_1517);
nand U3568 (N_3568,N_1512,N_1621);
xnor U3569 (N_3569,N_2274,N_1396);
nand U3570 (N_3570,N_2038,N_2232);
or U3571 (N_3571,N_2033,N_1982);
and U3572 (N_3572,N_2393,N_1471);
and U3573 (N_3573,N_2364,N_2316);
xnor U3574 (N_3574,N_1596,N_1645);
nor U3575 (N_3575,N_1498,N_2428);
xnor U3576 (N_3576,N_1394,N_1580);
or U3577 (N_3577,N_2244,N_1597);
xnor U3578 (N_3578,N_1654,N_2051);
nand U3579 (N_3579,N_1925,N_1702);
or U3580 (N_3580,N_1359,N_2125);
xor U3581 (N_3581,N_1601,N_1688);
nor U3582 (N_3582,N_1508,N_2019);
xor U3583 (N_3583,N_2062,N_1718);
and U3584 (N_3584,N_2346,N_1634);
nand U3585 (N_3585,N_1977,N_1943);
nor U3586 (N_3586,N_1904,N_1533);
nor U3587 (N_3587,N_2368,N_1959);
and U3588 (N_3588,N_1470,N_1926);
xnor U3589 (N_3589,N_1673,N_1489);
nand U3590 (N_3590,N_2049,N_2073);
and U3591 (N_3591,N_1755,N_1578);
nand U3592 (N_3592,N_2078,N_1570);
nor U3593 (N_3593,N_1335,N_2398);
nor U3594 (N_3594,N_2382,N_2185);
and U3595 (N_3595,N_1784,N_2169);
or U3596 (N_3596,N_1347,N_2082);
xnor U3597 (N_3597,N_1356,N_2251);
and U3598 (N_3598,N_2008,N_2229);
nor U3599 (N_3599,N_2155,N_1946);
nor U3600 (N_3600,N_2314,N_2015);
and U3601 (N_3601,N_2412,N_1810);
nand U3602 (N_3602,N_1953,N_1372);
nor U3603 (N_3603,N_2212,N_2463);
xor U3604 (N_3604,N_2073,N_1377);
and U3605 (N_3605,N_2478,N_2025);
and U3606 (N_3606,N_2139,N_2480);
and U3607 (N_3607,N_2336,N_2459);
xor U3608 (N_3608,N_2162,N_1581);
nand U3609 (N_3609,N_1274,N_1726);
nand U3610 (N_3610,N_2007,N_1658);
xor U3611 (N_3611,N_2297,N_1589);
nor U3612 (N_3612,N_1669,N_2098);
xor U3613 (N_3613,N_2252,N_1439);
nand U3614 (N_3614,N_2183,N_1379);
and U3615 (N_3615,N_1974,N_2440);
and U3616 (N_3616,N_1261,N_1423);
nand U3617 (N_3617,N_2275,N_1986);
nand U3618 (N_3618,N_2199,N_1325);
and U3619 (N_3619,N_1714,N_1346);
nor U3620 (N_3620,N_2071,N_1371);
xor U3621 (N_3621,N_1697,N_1575);
xor U3622 (N_3622,N_1937,N_1393);
nand U3623 (N_3623,N_2090,N_1814);
and U3624 (N_3624,N_1858,N_2156);
or U3625 (N_3625,N_2403,N_1673);
nor U3626 (N_3626,N_1386,N_1562);
and U3627 (N_3627,N_2481,N_2431);
xnor U3628 (N_3628,N_2188,N_1975);
nand U3629 (N_3629,N_2418,N_1917);
or U3630 (N_3630,N_2039,N_2086);
and U3631 (N_3631,N_1486,N_1384);
xnor U3632 (N_3632,N_1800,N_2417);
and U3633 (N_3633,N_2321,N_2226);
or U3634 (N_3634,N_1727,N_2476);
nand U3635 (N_3635,N_2412,N_1405);
and U3636 (N_3636,N_1555,N_2221);
and U3637 (N_3637,N_1454,N_2123);
nand U3638 (N_3638,N_1446,N_1791);
nand U3639 (N_3639,N_1882,N_1830);
nor U3640 (N_3640,N_1433,N_1377);
and U3641 (N_3641,N_1856,N_1589);
nand U3642 (N_3642,N_1409,N_2254);
nand U3643 (N_3643,N_1722,N_1290);
nand U3644 (N_3644,N_1711,N_1635);
nand U3645 (N_3645,N_2313,N_1950);
and U3646 (N_3646,N_2255,N_2388);
or U3647 (N_3647,N_2161,N_2027);
or U3648 (N_3648,N_2110,N_1600);
nor U3649 (N_3649,N_2154,N_2017);
nor U3650 (N_3650,N_1985,N_1279);
nand U3651 (N_3651,N_2000,N_2010);
or U3652 (N_3652,N_1617,N_2129);
or U3653 (N_3653,N_1666,N_1746);
nor U3654 (N_3654,N_1976,N_2398);
or U3655 (N_3655,N_2030,N_2344);
or U3656 (N_3656,N_1612,N_1718);
nand U3657 (N_3657,N_1547,N_2208);
nand U3658 (N_3658,N_2188,N_2225);
nand U3659 (N_3659,N_1366,N_2193);
nand U3660 (N_3660,N_2233,N_1724);
and U3661 (N_3661,N_1380,N_1549);
or U3662 (N_3662,N_2006,N_1923);
nor U3663 (N_3663,N_1565,N_1467);
and U3664 (N_3664,N_2127,N_2050);
and U3665 (N_3665,N_1913,N_2317);
and U3666 (N_3666,N_2452,N_1582);
and U3667 (N_3667,N_1434,N_1291);
nand U3668 (N_3668,N_1253,N_1320);
or U3669 (N_3669,N_1346,N_2444);
or U3670 (N_3670,N_2496,N_2057);
nand U3671 (N_3671,N_1785,N_1583);
nor U3672 (N_3672,N_1349,N_1606);
nand U3673 (N_3673,N_2063,N_2093);
nand U3674 (N_3674,N_1745,N_1327);
and U3675 (N_3675,N_1511,N_1568);
nand U3676 (N_3676,N_1297,N_1820);
xnor U3677 (N_3677,N_2258,N_1907);
xnor U3678 (N_3678,N_2200,N_1350);
and U3679 (N_3679,N_1727,N_2186);
xnor U3680 (N_3680,N_2217,N_2240);
nor U3681 (N_3681,N_1712,N_2184);
and U3682 (N_3682,N_1681,N_1745);
xnor U3683 (N_3683,N_1652,N_2187);
and U3684 (N_3684,N_2152,N_1796);
and U3685 (N_3685,N_2102,N_2432);
xnor U3686 (N_3686,N_1349,N_1497);
xor U3687 (N_3687,N_1519,N_2052);
xor U3688 (N_3688,N_2490,N_1712);
and U3689 (N_3689,N_2499,N_2447);
and U3690 (N_3690,N_1631,N_1942);
xnor U3691 (N_3691,N_1510,N_2389);
nand U3692 (N_3692,N_2072,N_2191);
nand U3693 (N_3693,N_1510,N_2075);
nand U3694 (N_3694,N_1347,N_2164);
nor U3695 (N_3695,N_2231,N_2345);
or U3696 (N_3696,N_2213,N_1919);
and U3697 (N_3697,N_1943,N_1907);
nand U3698 (N_3698,N_2077,N_2188);
xnor U3699 (N_3699,N_2448,N_1555);
nand U3700 (N_3700,N_2128,N_2438);
nand U3701 (N_3701,N_2062,N_2017);
or U3702 (N_3702,N_1520,N_1638);
xor U3703 (N_3703,N_2316,N_1374);
nor U3704 (N_3704,N_2266,N_1544);
or U3705 (N_3705,N_1364,N_1555);
nor U3706 (N_3706,N_2484,N_2201);
and U3707 (N_3707,N_2079,N_2438);
nor U3708 (N_3708,N_1310,N_2447);
and U3709 (N_3709,N_1459,N_2438);
xnor U3710 (N_3710,N_1998,N_1588);
and U3711 (N_3711,N_2371,N_1908);
nor U3712 (N_3712,N_2046,N_2031);
or U3713 (N_3713,N_2467,N_1590);
xor U3714 (N_3714,N_2273,N_2236);
and U3715 (N_3715,N_1801,N_1606);
and U3716 (N_3716,N_1694,N_2348);
and U3717 (N_3717,N_1803,N_2436);
or U3718 (N_3718,N_2393,N_1946);
nor U3719 (N_3719,N_1708,N_1558);
and U3720 (N_3720,N_2024,N_1523);
nand U3721 (N_3721,N_1642,N_1768);
or U3722 (N_3722,N_2268,N_1878);
and U3723 (N_3723,N_1665,N_1318);
xnor U3724 (N_3724,N_1987,N_1714);
nand U3725 (N_3725,N_1279,N_1882);
nand U3726 (N_3726,N_2255,N_1576);
nand U3727 (N_3727,N_1740,N_1690);
or U3728 (N_3728,N_2299,N_1806);
or U3729 (N_3729,N_1926,N_1526);
nor U3730 (N_3730,N_1965,N_2250);
xnor U3731 (N_3731,N_1690,N_1333);
nand U3732 (N_3732,N_2498,N_1381);
xor U3733 (N_3733,N_1778,N_1745);
xor U3734 (N_3734,N_2389,N_2154);
nand U3735 (N_3735,N_2290,N_2270);
or U3736 (N_3736,N_2228,N_1310);
nand U3737 (N_3737,N_1777,N_1973);
xor U3738 (N_3738,N_2384,N_2398);
xnor U3739 (N_3739,N_1401,N_1356);
xnor U3740 (N_3740,N_2463,N_1690);
and U3741 (N_3741,N_1286,N_1940);
or U3742 (N_3742,N_2404,N_1528);
and U3743 (N_3743,N_1976,N_1575);
and U3744 (N_3744,N_1265,N_1417);
nor U3745 (N_3745,N_1426,N_1589);
nand U3746 (N_3746,N_1371,N_1667);
and U3747 (N_3747,N_2462,N_1438);
nor U3748 (N_3748,N_1352,N_2147);
and U3749 (N_3749,N_1977,N_1886);
xor U3750 (N_3750,N_2913,N_3033);
and U3751 (N_3751,N_3267,N_3490);
or U3752 (N_3752,N_3320,N_3656);
nor U3753 (N_3753,N_3429,N_2517);
xnor U3754 (N_3754,N_2682,N_3297);
or U3755 (N_3755,N_3091,N_2527);
or U3756 (N_3756,N_2824,N_2816);
nand U3757 (N_3757,N_2658,N_3343);
nand U3758 (N_3758,N_2942,N_2989);
nor U3759 (N_3759,N_3349,N_3118);
xnor U3760 (N_3760,N_3261,N_2822);
nand U3761 (N_3761,N_3417,N_3218);
and U3762 (N_3762,N_3010,N_3306);
nand U3763 (N_3763,N_2814,N_2876);
xor U3764 (N_3764,N_3679,N_3152);
nand U3765 (N_3765,N_3649,N_3743);
nor U3766 (N_3766,N_3541,N_2736);
nor U3767 (N_3767,N_3073,N_2661);
nor U3768 (N_3768,N_3702,N_3722);
xor U3769 (N_3769,N_2568,N_2811);
nor U3770 (N_3770,N_3068,N_3256);
xnor U3771 (N_3771,N_2983,N_3381);
and U3772 (N_3772,N_2589,N_3403);
xnor U3773 (N_3773,N_3504,N_3575);
nand U3774 (N_3774,N_2614,N_3131);
or U3775 (N_3775,N_2677,N_3627);
and U3776 (N_3776,N_3479,N_2696);
and U3777 (N_3777,N_3112,N_2738);
or U3778 (N_3778,N_3132,N_2698);
nor U3779 (N_3779,N_3147,N_3527);
xnor U3780 (N_3780,N_3317,N_3470);
nand U3781 (N_3781,N_2821,N_2979);
nor U3782 (N_3782,N_2735,N_2866);
xor U3783 (N_3783,N_3310,N_3720);
nand U3784 (N_3784,N_3681,N_2687);
and U3785 (N_3785,N_2536,N_2785);
xor U3786 (N_3786,N_3712,N_3356);
and U3787 (N_3787,N_2671,N_2935);
nor U3788 (N_3788,N_3055,N_2774);
and U3789 (N_3789,N_3345,N_2744);
nand U3790 (N_3790,N_3071,N_3225);
and U3791 (N_3791,N_3264,N_2553);
or U3792 (N_3792,N_2549,N_3038);
or U3793 (N_3793,N_2692,N_2723);
and U3794 (N_3794,N_3259,N_2753);
and U3795 (N_3795,N_2654,N_3483);
nor U3796 (N_3796,N_3704,N_3005);
xnor U3797 (N_3797,N_3083,N_2513);
or U3798 (N_3798,N_3206,N_3555);
xnor U3799 (N_3799,N_2604,N_3051);
or U3800 (N_3800,N_2707,N_3011);
or U3801 (N_3801,N_2665,N_3420);
and U3802 (N_3802,N_3528,N_3523);
nand U3803 (N_3803,N_2904,N_2647);
nand U3804 (N_3804,N_3154,N_3582);
nor U3805 (N_3805,N_3579,N_2885);
nor U3806 (N_3806,N_3397,N_3244);
or U3807 (N_3807,N_2962,N_2512);
or U3808 (N_3808,N_2590,N_3458);
nand U3809 (N_3809,N_3623,N_2588);
nor U3810 (N_3810,N_2628,N_3733);
nor U3811 (N_3811,N_3373,N_3738);
nor U3812 (N_3812,N_2778,N_3561);
or U3813 (N_3813,N_3725,N_3090);
nor U3814 (N_3814,N_2612,N_3336);
nor U3815 (N_3815,N_3107,N_3439);
or U3816 (N_3816,N_3181,N_2930);
nand U3817 (N_3817,N_3583,N_2873);
or U3818 (N_3818,N_3276,N_3000);
and U3819 (N_3819,N_2722,N_3248);
or U3820 (N_3820,N_3468,N_3441);
nand U3821 (N_3821,N_2789,N_2515);
nor U3822 (N_3822,N_3353,N_3632);
nand U3823 (N_3823,N_2842,N_3238);
nor U3824 (N_3824,N_2781,N_2804);
nand U3825 (N_3825,N_2859,N_2543);
or U3826 (N_3826,N_3066,N_3654);
and U3827 (N_3827,N_2884,N_2847);
and U3828 (N_3828,N_3390,N_2598);
xor U3829 (N_3829,N_2636,N_3697);
and U3830 (N_3830,N_3499,N_2971);
and U3831 (N_3831,N_3492,N_2887);
nor U3832 (N_3832,N_2525,N_3331);
and U3833 (N_3833,N_2668,N_3495);
nand U3834 (N_3834,N_2681,N_3172);
and U3835 (N_3835,N_3675,N_2911);
nand U3836 (N_3836,N_3642,N_3683);
xnor U3837 (N_3837,N_2910,N_3707);
nor U3838 (N_3838,N_3569,N_2531);
and U3839 (N_3839,N_2666,N_2902);
nand U3840 (N_3840,N_3393,N_2796);
or U3841 (N_3841,N_3173,N_3482);
nor U3842 (N_3842,N_3544,N_2786);
or U3843 (N_3843,N_3277,N_3467);
nor U3844 (N_3844,N_2906,N_3494);
and U3845 (N_3845,N_3551,N_3060);
or U3846 (N_3846,N_2769,N_3574);
and U3847 (N_3847,N_3601,N_3568);
and U3848 (N_3848,N_3175,N_2932);
nor U3849 (N_3849,N_3588,N_3489);
xor U3850 (N_3850,N_2702,N_3700);
nor U3851 (N_3851,N_3059,N_2745);
and U3852 (N_3852,N_3315,N_3339);
nand U3853 (N_3853,N_2924,N_3240);
xnor U3854 (N_3854,N_3521,N_3084);
nor U3855 (N_3855,N_3602,N_3460);
nand U3856 (N_3856,N_3703,N_2909);
nand U3857 (N_3857,N_3556,N_2990);
xnor U3858 (N_3858,N_3043,N_2936);
and U3859 (N_3859,N_2922,N_3137);
xor U3860 (N_3860,N_2664,N_3485);
nand U3861 (N_3861,N_3730,N_3678);
nor U3862 (N_3862,N_3616,N_2505);
nor U3863 (N_3863,N_3028,N_2503);
xnor U3864 (N_3864,N_3061,N_3701);
xnor U3865 (N_3865,N_2894,N_3493);
and U3866 (N_3866,N_2504,N_3526);
xnor U3867 (N_3867,N_2943,N_2896);
and U3868 (N_3868,N_3635,N_2556);
or U3869 (N_3869,N_3198,N_2779);
nor U3870 (N_3870,N_3130,N_2939);
nor U3871 (N_3871,N_2584,N_3324);
or U3872 (N_3872,N_2891,N_3149);
xnor U3873 (N_3873,N_3472,N_3138);
xor U3874 (N_3874,N_2831,N_2624);
xnor U3875 (N_3875,N_3204,N_2637);
or U3876 (N_3876,N_3682,N_3186);
nor U3877 (N_3877,N_2791,N_3419);
or U3878 (N_3878,N_3525,N_3507);
nand U3879 (N_3879,N_3039,N_3653);
and U3880 (N_3880,N_3257,N_2923);
or U3881 (N_3881,N_2729,N_2975);
xnor U3882 (N_3882,N_3471,N_3572);
or U3883 (N_3883,N_2730,N_2806);
or U3884 (N_3884,N_3481,N_3219);
xor U3885 (N_3885,N_3295,N_3271);
nand U3886 (N_3886,N_2965,N_3311);
nand U3887 (N_3887,N_3533,N_3550);
and U3888 (N_3888,N_3562,N_2558);
or U3889 (N_3889,N_2620,N_2949);
xor U3890 (N_3890,N_3387,N_3369);
nor U3891 (N_3891,N_2581,N_3136);
or U3892 (N_3892,N_3727,N_2925);
nor U3893 (N_3893,N_2907,N_3056);
xnor U3894 (N_3894,N_3411,N_3203);
or U3895 (N_3895,N_3126,N_2711);
or U3896 (N_3896,N_2599,N_2714);
and U3897 (N_3897,N_3386,N_2602);
nor U3898 (N_3898,N_3148,N_3615);
nand U3899 (N_3899,N_2748,N_2691);
or U3900 (N_3900,N_3690,N_2921);
or U3901 (N_3901,N_3652,N_3625);
nand U3902 (N_3902,N_2900,N_3414);
and U3903 (N_3903,N_3170,N_3183);
and U3904 (N_3904,N_2838,N_3057);
and U3905 (N_3905,N_2863,N_3634);
or U3906 (N_3906,N_3480,N_3564);
and U3907 (N_3907,N_3484,N_2659);
or U3908 (N_3908,N_3451,N_3536);
nor U3909 (N_3909,N_3191,N_3402);
nor U3910 (N_3910,N_2856,N_2807);
xor U3911 (N_3911,N_3037,N_2693);
and U3912 (N_3912,N_3721,N_3698);
and U3913 (N_3913,N_3178,N_3629);
nand U3914 (N_3914,N_2746,N_3158);
nor U3915 (N_3915,N_3109,N_3252);
xnor U3916 (N_3916,N_2537,N_3025);
xor U3917 (N_3917,N_3724,N_3580);
nor U3918 (N_3918,N_2716,N_3278);
nand U3919 (N_3919,N_3294,N_3367);
nand U3920 (N_3920,N_2782,N_3245);
or U3921 (N_3921,N_3094,N_3344);
xnor U3922 (N_3922,N_3554,N_2643);
or U3923 (N_3923,N_2882,N_3024);
nand U3924 (N_3924,N_3391,N_3065);
nor U3925 (N_3925,N_3321,N_3049);
or U3926 (N_3926,N_3229,N_3141);
and U3927 (N_3927,N_2669,N_3101);
nor U3928 (N_3928,N_3664,N_2713);
nor U3929 (N_3929,N_3736,N_2552);
nor U3930 (N_3930,N_2572,N_3217);
nand U3931 (N_3931,N_2964,N_2697);
nand U3932 (N_3932,N_3041,N_2890);
xor U3933 (N_3933,N_2733,N_3437);
nand U3934 (N_3934,N_2802,N_3513);
or U3935 (N_3935,N_2564,N_3202);
xnor U3936 (N_3936,N_2893,N_2960);
xnor U3937 (N_3937,N_3416,N_3630);
nand U3938 (N_3938,N_3425,N_2644);
and U3939 (N_3939,N_2954,N_3571);
nand U3940 (N_3940,N_3230,N_2724);
xor U3941 (N_3941,N_2656,N_3508);
nor U3942 (N_3942,N_3027,N_3226);
xnor U3943 (N_3943,N_3124,N_3274);
nor U3944 (N_3944,N_2818,N_2749);
xor U3945 (N_3945,N_3286,N_2800);
xor U3946 (N_3946,N_2974,N_2805);
xnor U3947 (N_3947,N_3079,N_3749);
nor U3948 (N_3948,N_2538,N_2817);
nor U3949 (N_3949,N_3577,N_2867);
nor U3950 (N_3950,N_2550,N_3099);
or U3951 (N_3951,N_2596,N_3398);
nand U3952 (N_3952,N_2747,N_3449);
or U3953 (N_3953,N_3434,N_2988);
and U3954 (N_3954,N_3201,N_3475);
nand U3955 (N_3955,N_3503,N_3742);
and U3956 (N_3956,N_3436,N_3168);
xnor U3957 (N_3957,N_3077,N_2917);
nor U3958 (N_3958,N_3631,N_3641);
nor U3959 (N_3959,N_3044,N_2653);
nand U3960 (N_3960,N_3313,N_3714);
and U3961 (N_3961,N_3740,N_3680);
and U3962 (N_3962,N_3666,N_2507);
nor U3963 (N_3963,N_3422,N_3358);
xnor U3964 (N_3964,N_3308,N_3007);
nand U3965 (N_3965,N_2751,N_2928);
or U3966 (N_3966,N_3705,N_3624);
or U3967 (N_3967,N_2732,N_2768);
nor U3968 (N_3968,N_3734,N_2919);
nor U3969 (N_3969,N_3455,N_3171);
or U3970 (N_3970,N_3184,N_2511);
or U3971 (N_3971,N_2554,N_3281);
xnor U3972 (N_3972,N_2667,N_2845);
nand U3973 (N_3973,N_2872,N_3578);
xnor U3974 (N_3974,N_3323,N_2575);
and U3975 (N_3975,N_2903,N_2871);
and U3976 (N_3976,N_3549,N_2577);
nand U3977 (N_3977,N_2870,N_2686);
nand U3978 (N_3978,N_3535,N_2993);
xor U3979 (N_3979,N_3164,N_3200);
or U3980 (N_3980,N_2840,N_3511);
nand U3981 (N_3981,N_3696,N_3280);
and U3982 (N_3982,N_2999,N_2648);
nand U3983 (N_3983,N_3223,N_3553);
xor U3984 (N_3984,N_3473,N_3161);
and U3985 (N_3985,N_3426,N_2679);
nand U3986 (N_3986,N_3302,N_2623);
or U3987 (N_3987,N_2819,N_3019);
nor U3988 (N_3988,N_2798,N_3305);
and U3989 (N_3989,N_3097,N_2597);
and U3990 (N_3990,N_2897,N_3266);
nand U3991 (N_3991,N_3212,N_2908);
or U3992 (N_3992,N_2984,N_3529);
xnor U3993 (N_3993,N_3500,N_2670);
and U3994 (N_3994,N_3466,N_3585);
xor U3995 (N_3995,N_3092,N_2547);
or U3996 (N_3996,N_3524,N_3594);
nand U3997 (N_3997,N_3328,N_2613);
xnor U3998 (N_3998,N_3260,N_3663);
nor U3999 (N_3999,N_2569,N_3192);
or U4000 (N_4000,N_3213,N_3231);
or U4001 (N_4001,N_2756,N_3089);
or U4002 (N_4002,N_3383,N_2823);
and U4003 (N_4003,N_3012,N_3341);
and U4004 (N_4004,N_3163,N_3384);
xor U4005 (N_4005,N_3478,N_3224);
or U4006 (N_4006,N_2795,N_2708);
or U4007 (N_4007,N_2948,N_2851);
or U4008 (N_4008,N_3412,N_2961);
and U4009 (N_4009,N_3016,N_3453);
or U4010 (N_4010,N_2833,N_2721);
xnor U4011 (N_4011,N_3346,N_2642);
nor U4012 (N_4012,N_3116,N_3177);
and U4013 (N_4013,N_3318,N_2632);
and U4014 (N_4014,N_3014,N_3273);
or U4015 (N_4015,N_3423,N_2898);
xnor U4016 (N_4016,N_2991,N_2740);
nor U4017 (N_4017,N_2663,N_3459);
nor U4018 (N_4018,N_2530,N_2675);
nand U4019 (N_4019,N_3214,N_3618);
xnor U4020 (N_4020,N_3023,N_2826);
nor U4021 (N_4021,N_3581,N_3247);
or U4022 (N_4022,N_3253,N_2973);
or U4023 (N_4023,N_2947,N_3570);
xor U4024 (N_4024,N_3462,N_3543);
nand U4025 (N_4025,N_3102,N_3539);
xor U4026 (N_4026,N_3001,N_3607);
nand U4027 (N_4027,N_3193,N_3319);
nand U4028 (N_4028,N_2699,N_3665);
nor U4029 (N_4029,N_2758,N_2690);
nor U4030 (N_4030,N_3352,N_2874);
and U4031 (N_4031,N_3316,N_3254);
or U4032 (N_4032,N_3669,N_2743);
nor U4033 (N_4033,N_2627,N_2830);
and U4034 (N_4034,N_3537,N_3235);
nor U4035 (N_4035,N_3687,N_3715);
xnor U4036 (N_4036,N_3400,N_2715);
xnor U4037 (N_4037,N_2757,N_2883);
nand U4038 (N_4038,N_3337,N_3379);
and U4039 (N_4039,N_2764,N_3729);
and U4040 (N_4040,N_2912,N_2680);
xnor U4041 (N_4041,N_3165,N_2944);
xor U4042 (N_4042,N_2646,N_3643);
and U4043 (N_4043,N_3100,N_2762);
and U4044 (N_4044,N_2520,N_2809);
nor U4045 (N_4045,N_3408,N_2559);
and U4046 (N_4046,N_2931,N_3667);
nor U4047 (N_4047,N_3452,N_3135);
or U4048 (N_4048,N_3444,N_3140);
nand U4049 (N_4049,N_3628,N_3128);
xnor U4050 (N_4050,N_3435,N_3519);
xnor U4051 (N_4051,N_3354,N_3620);
nor U4052 (N_4052,N_2546,N_3211);
nand U4053 (N_4053,N_3693,N_3166);
or U4054 (N_4054,N_2524,N_2563);
nand U4055 (N_4055,N_3127,N_3143);
and U4056 (N_4056,N_2742,N_2560);
and U4057 (N_4057,N_2638,N_3695);
and U4058 (N_4058,N_2618,N_2765);
or U4059 (N_4059,N_3427,N_2880);
nor U4060 (N_4060,N_2548,N_3366);
nand U4061 (N_4061,N_3283,N_3232);
and U4062 (N_4062,N_3476,N_3325);
nor U4063 (N_4063,N_3189,N_2850);
nand U4064 (N_4064,N_3176,N_2683);
or U4065 (N_4065,N_2771,N_3456);
and U4066 (N_4066,N_3668,N_2706);
and U4067 (N_4067,N_3610,N_3545);
and U4068 (N_4068,N_3002,N_2980);
and U4069 (N_4069,N_2593,N_3021);
and U4070 (N_4070,N_3560,N_2797);
and U4071 (N_4071,N_2532,N_2727);
or U4072 (N_4072,N_3598,N_3103);
nand U4073 (N_4073,N_3591,N_3399);
nor U4074 (N_4074,N_3361,N_2739);
nor U4075 (N_4075,N_3246,N_3409);
xnor U4076 (N_4076,N_2545,N_2500);
nor U4077 (N_4077,N_3241,N_2508);
nand U4078 (N_4078,N_3626,N_2578);
nand U4079 (N_4079,N_2834,N_3650);
and U4080 (N_4080,N_3413,N_2995);
nand U4081 (N_4081,N_3491,N_2986);
xor U4082 (N_4082,N_3078,N_3015);
or U4083 (N_4083,N_2875,N_3329);
and U4084 (N_4084,N_3685,N_2889);
nor U4085 (N_4085,N_2676,N_3122);
nand U4086 (N_4086,N_3454,N_2997);
nor U4087 (N_4087,N_3717,N_3671);
xnor U4088 (N_4088,N_2619,N_3314);
and U4089 (N_4089,N_3081,N_2854);
and U4090 (N_4090,N_3121,N_2516);
or U4091 (N_4091,N_3639,N_3080);
nand U4092 (N_4092,N_2792,N_3157);
and U4093 (N_4093,N_3732,N_3646);
or U4094 (N_4094,N_3442,N_3162);
or U4095 (N_4095,N_2934,N_3054);
or U4096 (N_4096,N_2752,N_3405);
and U4097 (N_4097,N_3129,N_3350);
nor U4098 (N_4098,N_2719,N_3009);
and U4099 (N_4099,N_2678,N_3389);
or U4100 (N_4100,N_3293,N_3522);
or U4101 (N_4101,N_3558,N_3735);
xnor U4102 (N_4102,N_3067,N_3250);
xor U4103 (N_4103,N_3401,N_3603);
or U4104 (N_4104,N_2703,N_2565);
nor U4105 (N_4105,N_2937,N_3637);
nand U4106 (N_4106,N_3307,N_2825);
or U4107 (N_4107,N_3622,N_2591);
nand U4108 (N_4108,N_3388,N_3430);
nor U4109 (N_4109,N_3377,N_2726);
nor U4110 (N_4110,N_2855,N_3446);
and U4111 (N_4111,N_3301,N_3120);
and U4112 (N_4112,N_3392,N_3082);
nand U4113 (N_4113,N_2535,N_3676);
and U4114 (N_4114,N_3069,N_2561);
nor U4115 (N_4115,N_3565,N_3220);
nor U4116 (N_4116,N_3505,N_3029);
nor U4117 (N_4117,N_2881,N_3364);
xnor U4118 (N_4118,N_2640,N_3205);
and U4119 (N_4119,N_3547,N_3394);
nor U4120 (N_4120,N_3605,N_2794);
nor U4121 (N_4121,N_3110,N_3370);
or U4122 (N_4122,N_3125,N_3180);
nor U4123 (N_4123,N_3375,N_2555);
or U4124 (N_4124,N_3359,N_2501);
or U4125 (N_4125,N_2860,N_2868);
xor U4126 (N_4126,N_3123,N_2985);
nor U4127 (N_4127,N_3531,N_3284);
and U4128 (N_4128,N_3406,N_2601);
nand U4129 (N_4129,N_2837,N_3368);
xnor U4130 (N_4130,N_2694,N_3300);
xor U4131 (N_4131,N_3593,N_2629);
nor U4132 (N_4132,N_3443,N_2586);
nand U4133 (N_4133,N_2521,N_2631);
and U4134 (N_4134,N_3040,N_2731);
nand U4135 (N_4135,N_3322,N_2585);
nand U4136 (N_4136,N_2841,N_3279);
and U4137 (N_4137,N_3469,N_2953);
nand U4138 (N_4138,N_3621,N_2607);
xnor U4139 (N_4139,N_3728,N_3167);
nand U4140 (N_4140,N_2626,N_3106);
and U4141 (N_4141,N_3087,N_3008);
nand U4142 (N_4142,N_3378,N_3418);
or U4143 (N_4143,N_3196,N_3590);
xnor U4144 (N_4144,N_3619,N_3584);
or U4145 (N_4145,N_3255,N_2976);
or U4146 (N_4146,N_3215,N_2580);
and U4147 (N_4147,N_3382,N_3333);
or U4148 (N_4148,N_3496,N_3360);
or U4149 (N_4149,N_2633,N_2760);
and U4150 (N_4150,N_2522,N_3233);
or U4151 (N_4151,N_3239,N_3372);
or U4152 (N_4152,N_2570,N_3612);
and U4153 (N_4153,N_2672,N_2788);
and U4154 (N_4154,N_3731,N_2829);
and U4155 (N_4155,N_2750,N_3699);
and U4156 (N_4156,N_2968,N_2869);
xor U4157 (N_4157,N_2835,N_3509);
nand U4158 (N_4158,N_2886,N_2918);
nor U4159 (N_4159,N_2709,N_2542);
nor U4160 (N_4160,N_2783,N_3465);
nor U4161 (N_4161,N_2566,N_3312);
or U4162 (N_4162,N_2509,N_2801);
and U4163 (N_4163,N_2609,N_3433);
or U4164 (N_4164,N_3516,N_2526);
nand U4165 (N_4165,N_2622,N_2583);
nand U4166 (N_4166,N_3672,N_2810);
xor U4167 (N_4167,N_2978,N_3488);
or U4168 (N_4168,N_3748,N_3188);
or U4169 (N_4169,N_3546,N_2777);
and U4170 (N_4170,N_3611,N_3088);
nand U4171 (N_4171,N_3557,N_3114);
or U4172 (N_4172,N_3146,N_3365);
xor U4173 (N_4173,N_2787,N_3348);
and U4174 (N_4174,N_3265,N_3216);
nor U4175 (N_4175,N_2684,N_2674);
xnor U4176 (N_4176,N_3415,N_3046);
and U4177 (N_4177,N_2587,N_3661);
nor U4178 (N_4178,N_3221,N_2877);
xor U4179 (N_4179,N_2784,N_2926);
xnor U4180 (N_4180,N_3708,N_3096);
nor U4181 (N_4181,N_3063,N_3119);
or U4182 (N_4182,N_3692,N_2963);
and U4183 (N_4183,N_2813,N_3022);
or U4184 (N_4184,N_3694,N_3563);
or U4185 (N_4185,N_2861,N_2528);
or U4186 (N_4186,N_3351,N_3440);
nand U4187 (N_4187,N_3062,N_2630);
nand U4188 (N_4188,N_3645,N_3638);
nor U4189 (N_4189,N_3520,N_3395);
nor U4190 (N_4190,N_3438,N_3013);
nor U4191 (N_4191,N_3142,N_3272);
xor U4192 (N_4192,N_3604,N_3269);
and U4193 (N_4193,N_2717,N_3552);
and U4194 (N_4194,N_3113,N_2895);
and U4195 (N_4195,N_2506,N_2582);
nand U4196 (N_4196,N_2518,N_2815);
and U4197 (N_4197,N_2970,N_3338);
xor U4198 (N_4198,N_3709,N_3017);
nor U4199 (N_4199,N_2862,N_3020);
and U4200 (N_4200,N_3463,N_2579);
or U4201 (N_4201,N_3237,N_2767);
and U4202 (N_4202,N_3340,N_3291);
and U4203 (N_4203,N_3609,N_3518);
nor U4204 (N_4204,N_2892,N_2650);
nand U4205 (N_4205,N_3153,N_2969);
or U4206 (N_4206,N_2852,N_2849);
or U4207 (N_4207,N_3182,N_2865);
or U4208 (N_4208,N_3498,N_2879);
nand U4209 (N_4209,N_3108,N_3159);
and U4210 (N_4210,N_2941,N_3380);
or U4211 (N_4211,N_3744,N_3534);
nor U4212 (N_4212,N_2808,N_3457);
nand U4213 (N_4213,N_2625,N_2832);
nor U4214 (N_4214,N_2915,N_3673);
xnor U4215 (N_4215,N_2574,N_3195);
or U4216 (N_4216,N_2639,N_3035);
nor U4217 (N_4217,N_3289,N_3711);
xnor U4218 (N_4218,N_2950,N_3600);
xnor U4219 (N_4219,N_3573,N_3407);
xor U4220 (N_4220,N_2951,N_3053);
nor U4221 (N_4221,N_3243,N_3385);
xnor U4222 (N_4222,N_3648,N_3139);
xor U4223 (N_4223,N_3236,N_3258);
and U4224 (N_4224,N_2755,N_3086);
xor U4225 (N_4225,N_3737,N_3477);
and U4226 (N_4226,N_3270,N_2966);
nor U4227 (N_4227,N_3160,N_3093);
and U4228 (N_4228,N_2899,N_2780);
nor U4229 (N_4229,N_3559,N_3228);
and U4230 (N_4230,N_3633,N_3227);
xnor U4231 (N_4231,N_3145,N_3532);
xnor U4232 (N_4232,N_2701,N_2945);
nor U4233 (N_4233,N_3155,N_2938);
and U4234 (N_4234,N_2534,N_3501);
nor U4235 (N_4235,N_2621,N_2615);
nand U4236 (N_4236,N_3309,N_3031);
and U4237 (N_4237,N_2864,N_3647);
xor U4238 (N_4238,N_2967,N_3515);
xor U4239 (N_4239,N_3596,N_3156);
nand U4240 (N_4240,N_3670,N_3614);
xor U4241 (N_4241,N_3357,N_3150);
nand U4242 (N_4242,N_3303,N_3045);
xor U4243 (N_4243,N_3739,N_2734);
and U4244 (N_4244,N_2929,N_3330);
nand U4245 (N_4245,N_3288,N_3719);
xnor U4246 (N_4246,N_3464,N_2634);
or U4247 (N_4247,N_3432,N_2858);
and U4248 (N_4248,N_3599,N_3662);
nor U4249 (N_4249,N_2957,N_3404);
and U4250 (N_4250,N_3474,N_3296);
nor U4251 (N_4251,N_3197,N_3445);
or U4252 (N_4252,N_2741,N_3677);
xnor U4253 (N_4253,N_2611,N_3117);
nor U4254 (N_4254,N_3234,N_3174);
or U4255 (N_4255,N_3595,N_3208);
xor U4256 (N_4256,N_3502,N_3251);
or U4257 (N_4257,N_2617,N_2523);
and U4258 (N_4258,N_2952,N_3074);
and U4259 (N_4259,N_2776,N_3263);
nand U4260 (N_4260,N_3047,N_3487);
nand U4261 (N_4261,N_3510,N_3034);
nor U4262 (N_4262,N_2651,N_2994);
or U4263 (N_4263,N_2649,N_3542);
nand U4264 (N_4264,N_2914,N_3587);
nor U4265 (N_4265,N_2972,N_3608);
and U4266 (N_4266,N_3371,N_2737);
or U4267 (N_4267,N_3589,N_2901);
nor U4268 (N_4268,N_2959,N_2660);
nand U4269 (N_4269,N_2657,N_3032);
and U4270 (N_4270,N_3282,N_2595);
and U4271 (N_4271,N_2977,N_2514);
nand U4272 (N_4272,N_2608,N_3396);
nor U4273 (N_4273,N_3072,N_2704);
xor U4274 (N_4274,N_3644,N_3710);
and U4275 (N_4275,N_3249,N_3058);
xor U4276 (N_4276,N_2759,N_2853);
xnor U4277 (N_4277,N_2754,N_3660);
or U4278 (N_4278,N_3741,N_3085);
and U4279 (N_4279,N_3242,N_3207);
or U4280 (N_4280,N_2793,N_3374);
and U4281 (N_4281,N_2645,N_2539);
xor U4282 (N_4282,N_2848,N_3651);
and U4283 (N_4283,N_2946,N_2533);
or U4284 (N_4284,N_3190,N_2635);
nand U4285 (N_4285,N_2888,N_2562);
nor U4286 (N_4286,N_3144,N_3355);
or U4287 (N_4287,N_2955,N_2700);
xnor U4288 (N_4288,N_3640,N_2673);
xor U4289 (N_4289,N_2606,N_3030);
nor U4290 (N_4290,N_2710,N_3421);
or U4291 (N_4291,N_3098,N_3548);
nand U4292 (N_4292,N_3655,N_3111);
or U4293 (N_4293,N_3428,N_3179);
or U4294 (N_4294,N_3538,N_3448);
xor U4295 (N_4295,N_3567,N_3424);
nand U4296 (N_4296,N_2958,N_3362);
or U4297 (N_4297,N_3745,N_3342);
xnor U4298 (N_4298,N_3376,N_3530);
xnor U4299 (N_4299,N_3746,N_3209);
nor U4300 (N_4300,N_3684,N_3723);
nand U4301 (N_4301,N_3410,N_3688);
or U4302 (N_4302,N_3275,N_3115);
nand U4303 (N_4303,N_3747,N_2510);
and U4304 (N_4304,N_3185,N_2655);
and U4305 (N_4305,N_2662,N_2770);
nand U4306 (N_4306,N_2529,N_3050);
xor U4307 (N_4307,N_2772,N_2905);
nand U4308 (N_4308,N_2576,N_2933);
xor U4309 (N_4309,N_2616,N_3210);
xnor U4310 (N_4310,N_2844,N_2685);
nor U4311 (N_4311,N_3566,N_2519);
or U4312 (N_4312,N_2705,N_3299);
xor U4313 (N_4313,N_3613,N_3706);
or U4314 (N_4314,N_3486,N_2766);
xor U4315 (N_4315,N_3268,N_3586);
xor U4316 (N_4316,N_3018,N_2541);
nor U4317 (N_4317,N_3689,N_2920);
or U4318 (N_4318,N_2610,N_2956);
nand U4319 (N_4319,N_3076,N_2718);
or U4320 (N_4320,N_3095,N_3105);
xor U4321 (N_4321,N_3070,N_3327);
nand U4322 (N_4322,N_2987,N_3134);
xor U4323 (N_4323,N_3517,N_3512);
nor U4324 (N_4324,N_3674,N_3004);
or U4325 (N_4325,N_2551,N_3716);
nand U4326 (N_4326,N_3592,N_3718);
xor U4327 (N_4327,N_3576,N_3334);
and U4328 (N_4328,N_3659,N_3506);
and U4329 (N_4329,N_2544,N_2828);
nand U4330 (N_4330,N_3461,N_2998);
and U4331 (N_4331,N_2773,N_3048);
xnor U4332 (N_4332,N_3657,N_2592);
xor U4333 (N_4333,N_2763,N_3431);
and U4334 (N_4334,N_3658,N_3597);
xnor U4335 (N_4335,N_3363,N_2843);
nand U4336 (N_4336,N_3287,N_2688);
nand U4337 (N_4337,N_2839,N_3447);
xnor U4338 (N_4338,N_3133,N_3540);
nand U4339 (N_4339,N_3052,N_2605);
and U4340 (N_4340,N_3169,N_3026);
or U4341 (N_4341,N_2799,N_3686);
or U4342 (N_4342,N_2652,N_2712);
xnor U4343 (N_4343,N_3042,N_3151);
nor U4344 (N_4344,N_3347,N_3262);
nand U4345 (N_4345,N_2836,N_2725);
and U4346 (N_4346,N_2695,N_2982);
xnor U4347 (N_4347,N_2927,N_3326);
xnor U4348 (N_4348,N_3003,N_2720);
xor U4349 (N_4349,N_2812,N_2803);
nand U4350 (N_4350,N_3726,N_3497);
and U4351 (N_4351,N_3713,N_2981);
xor U4352 (N_4352,N_2600,N_2573);
xor U4353 (N_4353,N_3304,N_2594);
nor U4354 (N_4354,N_2761,N_3104);
and U4355 (N_4355,N_2603,N_3199);
and U4356 (N_4356,N_2820,N_3036);
xor U4357 (N_4357,N_3187,N_2775);
and U4358 (N_4358,N_3617,N_2728);
nor U4359 (N_4359,N_3292,N_2916);
nor U4360 (N_4360,N_3514,N_2502);
nor U4361 (N_4361,N_3075,N_3335);
and U4362 (N_4362,N_2827,N_2996);
nor U4363 (N_4363,N_3064,N_2846);
or U4364 (N_4364,N_2567,N_2992);
nor U4365 (N_4365,N_2857,N_2641);
nand U4366 (N_4366,N_2878,N_3290);
xnor U4367 (N_4367,N_2940,N_3006);
nor U4368 (N_4368,N_3450,N_3298);
and U4369 (N_4369,N_3285,N_2540);
nand U4370 (N_4370,N_3222,N_2557);
nor U4371 (N_4371,N_3691,N_3636);
xor U4372 (N_4372,N_2571,N_2689);
nand U4373 (N_4373,N_3606,N_3194);
nor U4374 (N_4374,N_3332,N_2790);
nor U4375 (N_4375,N_3474,N_3147);
nor U4376 (N_4376,N_3669,N_2953);
xor U4377 (N_4377,N_2937,N_2502);
and U4378 (N_4378,N_3456,N_3211);
nor U4379 (N_4379,N_3114,N_3403);
xor U4380 (N_4380,N_3318,N_2508);
nand U4381 (N_4381,N_3282,N_3735);
nand U4382 (N_4382,N_3131,N_3080);
nor U4383 (N_4383,N_3307,N_2918);
and U4384 (N_4384,N_2584,N_2641);
nor U4385 (N_4385,N_3574,N_3340);
or U4386 (N_4386,N_3740,N_2699);
and U4387 (N_4387,N_2920,N_3571);
and U4388 (N_4388,N_2884,N_2828);
xor U4389 (N_4389,N_3602,N_3713);
and U4390 (N_4390,N_2944,N_3405);
and U4391 (N_4391,N_3203,N_3186);
or U4392 (N_4392,N_3715,N_3326);
nand U4393 (N_4393,N_2522,N_3436);
and U4394 (N_4394,N_3332,N_3484);
nand U4395 (N_4395,N_3114,N_3293);
xor U4396 (N_4396,N_3118,N_2986);
nor U4397 (N_4397,N_3039,N_2550);
or U4398 (N_4398,N_3399,N_2910);
and U4399 (N_4399,N_3639,N_2572);
nand U4400 (N_4400,N_3036,N_3133);
nand U4401 (N_4401,N_3109,N_3449);
or U4402 (N_4402,N_3494,N_2930);
nand U4403 (N_4403,N_3253,N_3507);
nor U4404 (N_4404,N_3284,N_3401);
nand U4405 (N_4405,N_2521,N_2879);
xnor U4406 (N_4406,N_2542,N_2994);
nor U4407 (N_4407,N_3509,N_3251);
or U4408 (N_4408,N_3583,N_2944);
xnor U4409 (N_4409,N_2780,N_2972);
or U4410 (N_4410,N_3210,N_3578);
nor U4411 (N_4411,N_3703,N_3140);
xor U4412 (N_4412,N_3403,N_3187);
and U4413 (N_4413,N_3065,N_3687);
or U4414 (N_4414,N_2698,N_3183);
or U4415 (N_4415,N_3231,N_2991);
nand U4416 (N_4416,N_3274,N_3332);
xnor U4417 (N_4417,N_3386,N_3394);
or U4418 (N_4418,N_2956,N_3559);
or U4419 (N_4419,N_3101,N_3450);
and U4420 (N_4420,N_3238,N_3443);
nand U4421 (N_4421,N_2787,N_3568);
xor U4422 (N_4422,N_3178,N_2533);
xor U4423 (N_4423,N_3030,N_3187);
and U4424 (N_4424,N_2527,N_3249);
and U4425 (N_4425,N_3404,N_3192);
xor U4426 (N_4426,N_3268,N_3455);
xnor U4427 (N_4427,N_3058,N_3166);
xor U4428 (N_4428,N_2651,N_2922);
xor U4429 (N_4429,N_2548,N_3316);
or U4430 (N_4430,N_2509,N_2643);
or U4431 (N_4431,N_3246,N_3715);
and U4432 (N_4432,N_3385,N_3278);
xor U4433 (N_4433,N_2546,N_2595);
or U4434 (N_4434,N_2791,N_3073);
and U4435 (N_4435,N_3534,N_2746);
nor U4436 (N_4436,N_2518,N_3468);
nor U4437 (N_4437,N_3271,N_3283);
and U4438 (N_4438,N_3533,N_3021);
nand U4439 (N_4439,N_2927,N_3176);
nand U4440 (N_4440,N_2833,N_2674);
and U4441 (N_4441,N_2645,N_3491);
and U4442 (N_4442,N_3710,N_3334);
nand U4443 (N_4443,N_3381,N_2571);
or U4444 (N_4444,N_3705,N_2848);
nor U4445 (N_4445,N_3367,N_2842);
nand U4446 (N_4446,N_3338,N_3085);
or U4447 (N_4447,N_3126,N_3084);
nand U4448 (N_4448,N_2941,N_3640);
or U4449 (N_4449,N_2829,N_3082);
or U4450 (N_4450,N_2567,N_2509);
and U4451 (N_4451,N_3072,N_3407);
or U4452 (N_4452,N_2683,N_2500);
nor U4453 (N_4453,N_2956,N_2550);
or U4454 (N_4454,N_2786,N_2500);
xor U4455 (N_4455,N_2633,N_3423);
nand U4456 (N_4456,N_2620,N_3199);
nand U4457 (N_4457,N_3052,N_3395);
nand U4458 (N_4458,N_3205,N_2703);
xor U4459 (N_4459,N_2715,N_3251);
xor U4460 (N_4460,N_3095,N_3594);
nor U4461 (N_4461,N_2866,N_3491);
or U4462 (N_4462,N_3474,N_3675);
and U4463 (N_4463,N_3701,N_2693);
or U4464 (N_4464,N_2892,N_2710);
or U4465 (N_4465,N_3105,N_3382);
nor U4466 (N_4466,N_2594,N_3727);
and U4467 (N_4467,N_3023,N_3321);
or U4468 (N_4468,N_2749,N_2947);
nor U4469 (N_4469,N_3475,N_3410);
nor U4470 (N_4470,N_3734,N_3193);
nor U4471 (N_4471,N_3681,N_2876);
nand U4472 (N_4472,N_3126,N_3083);
and U4473 (N_4473,N_3486,N_3720);
nor U4474 (N_4474,N_2912,N_3247);
nor U4475 (N_4475,N_3297,N_3074);
nor U4476 (N_4476,N_3370,N_3459);
nor U4477 (N_4477,N_2623,N_3374);
or U4478 (N_4478,N_3441,N_2619);
nand U4479 (N_4479,N_3067,N_2779);
nor U4480 (N_4480,N_3675,N_2617);
xor U4481 (N_4481,N_3298,N_3459);
and U4482 (N_4482,N_3217,N_3229);
or U4483 (N_4483,N_2787,N_3345);
xnor U4484 (N_4484,N_2732,N_2889);
or U4485 (N_4485,N_3625,N_2556);
nand U4486 (N_4486,N_3408,N_3074);
or U4487 (N_4487,N_2597,N_3746);
and U4488 (N_4488,N_3558,N_3147);
nor U4489 (N_4489,N_2787,N_2670);
nand U4490 (N_4490,N_3183,N_2560);
or U4491 (N_4491,N_3077,N_2914);
xnor U4492 (N_4492,N_3633,N_3285);
and U4493 (N_4493,N_2989,N_3084);
or U4494 (N_4494,N_3262,N_3088);
and U4495 (N_4495,N_3211,N_2753);
and U4496 (N_4496,N_2609,N_2937);
nand U4497 (N_4497,N_3549,N_3175);
nand U4498 (N_4498,N_3215,N_3680);
xor U4499 (N_4499,N_3667,N_3428);
xnor U4500 (N_4500,N_3663,N_3551);
or U4501 (N_4501,N_3337,N_3714);
or U4502 (N_4502,N_2543,N_2742);
nand U4503 (N_4503,N_3069,N_2752);
and U4504 (N_4504,N_3402,N_2695);
and U4505 (N_4505,N_3571,N_3464);
or U4506 (N_4506,N_2504,N_3051);
and U4507 (N_4507,N_2735,N_3248);
or U4508 (N_4508,N_2581,N_3450);
nand U4509 (N_4509,N_3263,N_3450);
xnor U4510 (N_4510,N_2913,N_3389);
and U4511 (N_4511,N_3419,N_2591);
nand U4512 (N_4512,N_2715,N_3268);
or U4513 (N_4513,N_3469,N_3647);
or U4514 (N_4514,N_2893,N_3729);
and U4515 (N_4515,N_2610,N_3028);
nand U4516 (N_4516,N_3203,N_2853);
nor U4517 (N_4517,N_2907,N_2688);
nand U4518 (N_4518,N_2553,N_3031);
and U4519 (N_4519,N_3111,N_2700);
nand U4520 (N_4520,N_3004,N_2729);
nor U4521 (N_4521,N_2769,N_2588);
nor U4522 (N_4522,N_2773,N_2536);
and U4523 (N_4523,N_2737,N_3589);
and U4524 (N_4524,N_3556,N_3442);
nor U4525 (N_4525,N_2747,N_3385);
and U4526 (N_4526,N_2682,N_3032);
and U4527 (N_4527,N_3056,N_3547);
xnor U4528 (N_4528,N_3254,N_3182);
or U4529 (N_4529,N_2660,N_3697);
nand U4530 (N_4530,N_3638,N_2657);
nor U4531 (N_4531,N_3488,N_3544);
xnor U4532 (N_4532,N_3037,N_3079);
or U4533 (N_4533,N_3722,N_3320);
nand U4534 (N_4534,N_3565,N_3515);
and U4535 (N_4535,N_3081,N_3094);
or U4536 (N_4536,N_2610,N_3230);
nor U4537 (N_4537,N_2863,N_2829);
and U4538 (N_4538,N_3486,N_3610);
xor U4539 (N_4539,N_3332,N_2767);
xor U4540 (N_4540,N_3205,N_3627);
xnor U4541 (N_4541,N_3488,N_3119);
nand U4542 (N_4542,N_3468,N_2677);
nor U4543 (N_4543,N_3647,N_3165);
and U4544 (N_4544,N_2529,N_3403);
nand U4545 (N_4545,N_2705,N_3575);
nor U4546 (N_4546,N_2895,N_3024);
or U4547 (N_4547,N_2721,N_2889);
nor U4548 (N_4548,N_3458,N_3255);
nor U4549 (N_4549,N_2637,N_3339);
or U4550 (N_4550,N_3221,N_2693);
or U4551 (N_4551,N_2693,N_2912);
or U4552 (N_4552,N_3694,N_2793);
or U4553 (N_4553,N_3185,N_3124);
nor U4554 (N_4554,N_3304,N_3240);
or U4555 (N_4555,N_3732,N_3461);
and U4556 (N_4556,N_2552,N_3050);
nand U4557 (N_4557,N_2512,N_3011);
nand U4558 (N_4558,N_2706,N_2598);
nand U4559 (N_4559,N_3739,N_3746);
xnor U4560 (N_4560,N_3605,N_3347);
nand U4561 (N_4561,N_3237,N_2962);
xnor U4562 (N_4562,N_3539,N_3540);
nor U4563 (N_4563,N_3594,N_2914);
nor U4564 (N_4564,N_3655,N_2993);
or U4565 (N_4565,N_2818,N_2877);
nor U4566 (N_4566,N_3034,N_3582);
xor U4567 (N_4567,N_3280,N_2954);
or U4568 (N_4568,N_3217,N_2934);
nor U4569 (N_4569,N_3532,N_2501);
nor U4570 (N_4570,N_3294,N_3379);
or U4571 (N_4571,N_3480,N_3301);
or U4572 (N_4572,N_3634,N_3010);
nor U4573 (N_4573,N_3252,N_2790);
and U4574 (N_4574,N_2924,N_2938);
xnor U4575 (N_4575,N_2881,N_2726);
or U4576 (N_4576,N_3503,N_3458);
nor U4577 (N_4577,N_3737,N_3553);
or U4578 (N_4578,N_2586,N_3196);
or U4579 (N_4579,N_2798,N_3131);
xnor U4580 (N_4580,N_3340,N_3195);
nor U4581 (N_4581,N_2787,N_2834);
xor U4582 (N_4582,N_3394,N_3076);
xnor U4583 (N_4583,N_3658,N_2701);
or U4584 (N_4584,N_3016,N_2543);
nand U4585 (N_4585,N_3000,N_3220);
or U4586 (N_4586,N_2532,N_3292);
nor U4587 (N_4587,N_3096,N_3207);
and U4588 (N_4588,N_3376,N_3018);
nand U4589 (N_4589,N_3445,N_2644);
and U4590 (N_4590,N_2775,N_3253);
or U4591 (N_4591,N_3408,N_3545);
or U4592 (N_4592,N_3458,N_2760);
nor U4593 (N_4593,N_3191,N_3188);
and U4594 (N_4594,N_2545,N_2622);
nor U4595 (N_4595,N_3537,N_3673);
xnor U4596 (N_4596,N_3235,N_3485);
nor U4597 (N_4597,N_3418,N_3503);
nand U4598 (N_4598,N_3689,N_2593);
nor U4599 (N_4599,N_3700,N_2605);
nor U4600 (N_4600,N_2664,N_2771);
nand U4601 (N_4601,N_3692,N_2961);
nand U4602 (N_4602,N_3538,N_2868);
or U4603 (N_4603,N_3635,N_3030);
or U4604 (N_4604,N_3372,N_3120);
or U4605 (N_4605,N_3553,N_2787);
nand U4606 (N_4606,N_3277,N_3476);
nor U4607 (N_4607,N_2593,N_3598);
or U4608 (N_4608,N_3435,N_2718);
or U4609 (N_4609,N_3632,N_2813);
nor U4610 (N_4610,N_2504,N_2966);
and U4611 (N_4611,N_3737,N_2502);
nor U4612 (N_4612,N_3546,N_3609);
nand U4613 (N_4613,N_3397,N_2539);
nor U4614 (N_4614,N_2630,N_3041);
or U4615 (N_4615,N_3117,N_2647);
xnor U4616 (N_4616,N_3411,N_2852);
nand U4617 (N_4617,N_3320,N_3224);
or U4618 (N_4618,N_3690,N_2552);
nor U4619 (N_4619,N_2567,N_3480);
or U4620 (N_4620,N_2974,N_3416);
xnor U4621 (N_4621,N_3386,N_2685);
nand U4622 (N_4622,N_3624,N_2850);
xnor U4623 (N_4623,N_2828,N_2930);
nor U4624 (N_4624,N_2819,N_3442);
xnor U4625 (N_4625,N_3531,N_3050);
nor U4626 (N_4626,N_2537,N_2896);
and U4627 (N_4627,N_2901,N_3623);
or U4628 (N_4628,N_3325,N_3357);
and U4629 (N_4629,N_2768,N_3269);
or U4630 (N_4630,N_2607,N_3303);
xor U4631 (N_4631,N_2941,N_2649);
and U4632 (N_4632,N_3194,N_3660);
nor U4633 (N_4633,N_2535,N_2542);
or U4634 (N_4634,N_2828,N_2733);
and U4635 (N_4635,N_3518,N_3483);
or U4636 (N_4636,N_3199,N_2611);
xnor U4637 (N_4637,N_2971,N_3123);
or U4638 (N_4638,N_2658,N_3012);
xor U4639 (N_4639,N_3259,N_2658);
or U4640 (N_4640,N_3146,N_2797);
xnor U4641 (N_4641,N_3021,N_3563);
and U4642 (N_4642,N_3172,N_3539);
or U4643 (N_4643,N_3454,N_3615);
nand U4644 (N_4644,N_2691,N_2655);
xor U4645 (N_4645,N_3684,N_2565);
nor U4646 (N_4646,N_3730,N_2716);
xnor U4647 (N_4647,N_3256,N_3740);
nand U4648 (N_4648,N_2618,N_2803);
or U4649 (N_4649,N_2526,N_2912);
or U4650 (N_4650,N_2840,N_3411);
or U4651 (N_4651,N_3413,N_2501);
or U4652 (N_4652,N_2885,N_2913);
and U4653 (N_4653,N_3186,N_3118);
or U4654 (N_4654,N_3180,N_3375);
xnor U4655 (N_4655,N_2860,N_3115);
nand U4656 (N_4656,N_2974,N_3444);
xor U4657 (N_4657,N_2600,N_3693);
nor U4658 (N_4658,N_2740,N_2967);
nor U4659 (N_4659,N_3000,N_3560);
nor U4660 (N_4660,N_2694,N_2511);
nand U4661 (N_4661,N_3101,N_3462);
or U4662 (N_4662,N_3332,N_2558);
or U4663 (N_4663,N_3063,N_2772);
xor U4664 (N_4664,N_2737,N_2783);
xor U4665 (N_4665,N_2598,N_2522);
nor U4666 (N_4666,N_3241,N_2884);
and U4667 (N_4667,N_3068,N_2892);
nor U4668 (N_4668,N_2915,N_3531);
or U4669 (N_4669,N_3367,N_3049);
xor U4670 (N_4670,N_2528,N_3385);
nor U4671 (N_4671,N_2962,N_3266);
xnor U4672 (N_4672,N_3034,N_3406);
nand U4673 (N_4673,N_3553,N_3727);
and U4674 (N_4674,N_2865,N_2637);
nor U4675 (N_4675,N_3032,N_2783);
nor U4676 (N_4676,N_3698,N_3460);
xnor U4677 (N_4677,N_2765,N_3424);
and U4678 (N_4678,N_3538,N_2748);
and U4679 (N_4679,N_2754,N_3026);
nand U4680 (N_4680,N_3518,N_2525);
and U4681 (N_4681,N_3097,N_3738);
nand U4682 (N_4682,N_3233,N_3694);
nor U4683 (N_4683,N_3019,N_2778);
nand U4684 (N_4684,N_3354,N_3336);
nor U4685 (N_4685,N_3304,N_2826);
nand U4686 (N_4686,N_3314,N_2900);
and U4687 (N_4687,N_3153,N_2507);
and U4688 (N_4688,N_2716,N_3118);
xnor U4689 (N_4689,N_3578,N_3160);
and U4690 (N_4690,N_2817,N_2819);
xor U4691 (N_4691,N_2926,N_3344);
or U4692 (N_4692,N_3011,N_3352);
nor U4693 (N_4693,N_3408,N_2922);
nand U4694 (N_4694,N_2778,N_3365);
xnor U4695 (N_4695,N_2968,N_3059);
or U4696 (N_4696,N_2689,N_3630);
nand U4697 (N_4697,N_3499,N_3549);
nand U4698 (N_4698,N_3632,N_3208);
xnor U4699 (N_4699,N_2646,N_2812);
and U4700 (N_4700,N_3469,N_2883);
nor U4701 (N_4701,N_3304,N_3026);
nand U4702 (N_4702,N_3234,N_3707);
and U4703 (N_4703,N_2737,N_2571);
nand U4704 (N_4704,N_3705,N_3496);
or U4705 (N_4705,N_3714,N_3571);
and U4706 (N_4706,N_2542,N_3343);
nand U4707 (N_4707,N_3006,N_2987);
or U4708 (N_4708,N_3387,N_2904);
and U4709 (N_4709,N_2735,N_3686);
nand U4710 (N_4710,N_3431,N_3156);
xor U4711 (N_4711,N_3681,N_2922);
nand U4712 (N_4712,N_3661,N_3254);
nor U4713 (N_4713,N_2893,N_3268);
xor U4714 (N_4714,N_2917,N_3434);
nor U4715 (N_4715,N_2897,N_3270);
nand U4716 (N_4716,N_2724,N_3737);
and U4717 (N_4717,N_3057,N_3178);
or U4718 (N_4718,N_2778,N_3369);
or U4719 (N_4719,N_3501,N_3196);
or U4720 (N_4720,N_2676,N_3658);
or U4721 (N_4721,N_2733,N_3492);
or U4722 (N_4722,N_3352,N_3354);
or U4723 (N_4723,N_3089,N_3055);
nor U4724 (N_4724,N_3419,N_3708);
and U4725 (N_4725,N_3682,N_3717);
or U4726 (N_4726,N_3173,N_3144);
or U4727 (N_4727,N_2777,N_3624);
and U4728 (N_4728,N_3537,N_3332);
and U4729 (N_4729,N_2707,N_2521);
xnor U4730 (N_4730,N_3622,N_3625);
xnor U4731 (N_4731,N_3273,N_3199);
nand U4732 (N_4732,N_3147,N_3035);
nand U4733 (N_4733,N_3108,N_3323);
nand U4734 (N_4734,N_3685,N_2580);
and U4735 (N_4735,N_3006,N_2800);
nor U4736 (N_4736,N_3371,N_3376);
nor U4737 (N_4737,N_3109,N_2808);
xnor U4738 (N_4738,N_3621,N_3514);
nor U4739 (N_4739,N_2590,N_3675);
or U4740 (N_4740,N_3435,N_3487);
nand U4741 (N_4741,N_3633,N_3599);
nand U4742 (N_4742,N_2852,N_3525);
nor U4743 (N_4743,N_2865,N_3407);
or U4744 (N_4744,N_3081,N_3280);
and U4745 (N_4745,N_3349,N_3560);
and U4746 (N_4746,N_3024,N_3122);
nor U4747 (N_4747,N_2911,N_3234);
nor U4748 (N_4748,N_3516,N_3439);
nand U4749 (N_4749,N_3528,N_2910);
nand U4750 (N_4750,N_2631,N_2805);
nor U4751 (N_4751,N_3261,N_3567);
and U4752 (N_4752,N_2985,N_3620);
nand U4753 (N_4753,N_3333,N_3523);
and U4754 (N_4754,N_3329,N_3026);
nand U4755 (N_4755,N_3375,N_2842);
and U4756 (N_4756,N_3197,N_2511);
nor U4757 (N_4757,N_3080,N_3596);
xnor U4758 (N_4758,N_2766,N_3733);
or U4759 (N_4759,N_2656,N_2572);
and U4760 (N_4760,N_3425,N_3195);
nand U4761 (N_4761,N_2845,N_3312);
nor U4762 (N_4762,N_3435,N_2548);
or U4763 (N_4763,N_2882,N_2818);
nand U4764 (N_4764,N_3742,N_2778);
nor U4765 (N_4765,N_2847,N_3528);
and U4766 (N_4766,N_2800,N_3517);
nor U4767 (N_4767,N_3513,N_2798);
nor U4768 (N_4768,N_2855,N_3390);
and U4769 (N_4769,N_3676,N_3004);
or U4770 (N_4770,N_3185,N_2917);
nor U4771 (N_4771,N_3534,N_2679);
or U4772 (N_4772,N_3364,N_3133);
xor U4773 (N_4773,N_3083,N_3601);
nand U4774 (N_4774,N_3605,N_2545);
and U4775 (N_4775,N_3474,N_3588);
nand U4776 (N_4776,N_3744,N_3220);
xor U4777 (N_4777,N_2707,N_3026);
xor U4778 (N_4778,N_2991,N_2957);
nand U4779 (N_4779,N_2691,N_2624);
nand U4780 (N_4780,N_3131,N_3493);
and U4781 (N_4781,N_3736,N_3387);
and U4782 (N_4782,N_3070,N_2820);
nor U4783 (N_4783,N_3254,N_3603);
nand U4784 (N_4784,N_2970,N_3656);
and U4785 (N_4785,N_2915,N_3605);
nor U4786 (N_4786,N_3460,N_3370);
and U4787 (N_4787,N_2934,N_2802);
nand U4788 (N_4788,N_3258,N_3261);
nand U4789 (N_4789,N_3590,N_3167);
and U4790 (N_4790,N_3115,N_3336);
and U4791 (N_4791,N_3541,N_3397);
nand U4792 (N_4792,N_3431,N_3021);
xnor U4793 (N_4793,N_3435,N_3020);
nor U4794 (N_4794,N_3642,N_2707);
and U4795 (N_4795,N_3604,N_3579);
or U4796 (N_4796,N_2870,N_3085);
xnor U4797 (N_4797,N_3167,N_3653);
nand U4798 (N_4798,N_3599,N_3597);
and U4799 (N_4799,N_2837,N_3016);
nand U4800 (N_4800,N_3298,N_3086);
nand U4801 (N_4801,N_3668,N_3176);
or U4802 (N_4802,N_2777,N_3435);
nand U4803 (N_4803,N_3107,N_3244);
xor U4804 (N_4804,N_3484,N_3159);
and U4805 (N_4805,N_2822,N_3422);
and U4806 (N_4806,N_3668,N_2973);
or U4807 (N_4807,N_3094,N_3254);
and U4808 (N_4808,N_3441,N_3036);
nor U4809 (N_4809,N_2504,N_3353);
and U4810 (N_4810,N_3246,N_2971);
nand U4811 (N_4811,N_2914,N_3240);
nand U4812 (N_4812,N_3595,N_3081);
xnor U4813 (N_4813,N_2892,N_3604);
nand U4814 (N_4814,N_2597,N_2637);
and U4815 (N_4815,N_2573,N_2839);
and U4816 (N_4816,N_3291,N_2528);
nor U4817 (N_4817,N_3014,N_3196);
nand U4818 (N_4818,N_3237,N_2615);
xnor U4819 (N_4819,N_2974,N_2679);
nand U4820 (N_4820,N_2831,N_3235);
nor U4821 (N_4821,N_3284,N_3070);
xnor U4822 (N_4822,N_3629,N_3504);
nor U4823 (N_4823,N_3479,N_2658);
xnor U4824 (N_4824,N_3058,N_3101);
and U4825 (N_4825,N_3084,N_3017);
nor U4826 (N_4826,N_2703,N_2506);
xnor U4827 (N_4827,N_3644,N_3486);
nor U4828 (N_4828,N_3596,N_3573);
or U4829 (N_4829,N_2667,N_3195);
nand U4830 (N_4830,N_2529,N_3463);
or U4831 (N_4831,N_3060,N_3435);
nand U4832 (N_4832,N_2995,N_3361);
xor U4833 (N_4833,N_2939,N_2846);
and U4834 (N_4834,N_2964,N_2698);
nor U4835 (N_4835,N_3104,N_3091);
nor U4836 (N_4836,N_3308,N_3414);
and U4837 (N_4837,N_2600,N_3221);
and U4838 (N_4838,N_3393,N_3700);
nand U4839 (N_4839,N_2535,N_3042);
xor U4840 (N_4840,N_2725,N_2814);
nand U4841 (N_4841,N_3187,N_3659);
xnor U4842 (N_4842,N_2735,N_3739);
or U4843 (N_4843,N_3011,N_3179);
nor U4844 (N_4844,N_2875,N_3307);
and U4845 (N_4845,N_3291,N_2893);
nor U4846 (N_4846,N_3484,N_2791);
nand U4847 (N_4847,N_3484,N_3210);
and U4848 (N_4848,N_3209,N_3486);
and U4849 (N_4849,N_3257,N_3239);
xor U4850 (N_4850,N_3225,N_2673);
nand U4851 (N_4851,N_3166,N_3600);
and U4852 (N_4852,N_3739,N_2787);
xnor U4853 (N_4853,N_2636,N_2683);
nor U4854 (N_4854,N_3711,N_2576);
xor U4855 (N_4855,N_3623,N_2975);
nor U4856 (N_4856,N_3417,N_3575);
nand U4857 (N_4857,N_2982,N_3399);
or U4858 (N_4858,N_3221,N_3531);
or U4859 (N_4859,N_2548,N_3223);
or U4860 (N_4860,N_2714,N_2733);
or U4861 (N_4861,N_3348,N_2503);
or U4862 (N_4862,N_3291,N_3052);
or U4863 (N_4863,N_2786,N_3505);
nand U4864 (N_4864,N_2967,N_2580);
or U4865 (N_4865,N_2895,N_3532);
or U4866 (N_4866,N_3427,N_3632);
xnor U4867 (N_4867,N_2538,N_3597);
nor U4868 (N_4868,N_3080,N_3620);
nor U4869 (N_4869,N_3173,N_3601);
and U4870 (N_4870,N_3740,N_3534);
nor U4871 (N_4871,N_2928,N_3284);
and U4872 (N_4872,N_2868,N_3521);
nor U4873 (N_4873,N_3177,N_2650);
or U4874 (N_4874,N_3017,N_2797);
xor U4875 (N_4875,N_3484,N_3215);
or U4876 (N_4876,N_3210,N_3169);
and U4877 (N_4877,N_3256,N_3710);
xor U4878 (N_4878,N_2655,N_2551);
nor U4879 (N_4879,N_2556,N_3073);
nor U4880 (N_4880,N_2515,N_3456);
nand U4881 (N_4881,N_3590,N_3704);
xnor U4882 (N_4882,N_3566,N_2663);
and U4883 (N_4883,N_3280,N_2556);
or U4884 (N_4884,N_3664,N_2857);
nor U4885 (N_4885,N_3539,N_3721);
or U4886 (N_4886,N_2845,N_2660);
nand U4887 (N_4887,N_2820,N_3174);
nor U4888 (N_4888,N_3529,N_3270);
and U4889 (N_4889,N_2561,N_3687);
nor U4890 (N_4890,N_2574,N_3009);
or U4891 (N_4891,N_2525,N_2615);
nor U4892 (N_4892,N_2614,N_3521);
and U4893 (N_4893,N_3629,N_2917);
and U4894 (N_4894,N_2795,N_3709);
and U4895 (N_4895,N_2611,N_2676);
nor U4896 (N_4896,N_3061,N_3363);
and U4897 (N_4897,N_3434,N_3548);
xor U4898 (N_4898,N_2565,N_3332);
nand U4899 (N_4899,N_2871,N_3709);
or U4900 (N_4900,N_3214,N_2636);
or U4901 (N_4901,N_3579,N_3042);
nor U4902 (N_4902,N_3342,N_3628);
nand U4903 (N_4903,N_2903,N_3308);
or U4904 (N_4904,N_3236,N_3647);
nand U4905 (N_4905,N_3241,N_3708);
and U4906 (N_4906,N_2822,N_2685);
or U4907 (N_4907,N_3301,N_3572);
xnor U4908 (N_4908,N_3183,N_2675);
xor U4909 (N_4909,N_3272,N_2981);
or U4910 (N_4910,N_3604,N_3407);
and U4911 (N_4911,N_3374,N_3076);
or U4912 (N_4912,N_3046,N_3160);
nor U4913 (N_4913,N_3385,N_3037);
and U4914 (N_4914,N_3049,N_2827);
nand U4915 (N_4915,N_2951,N_2869);
and U4916 (N_4916,N_3401,N_3269);
and U4917 (N_4917,N_3391,N_2934);
nor U4918 (N_4918,N_3739,N_2773);
nand U4919 (N_4919,N_2784,N_3180);
xnor U4920 (N_4920,N_3693,N_2533);
or U4921 (N_4921,N_3234,N_2663);
and U4922 (N_4922,N_3608,N_3507);
nor U4923 (N_4923,N_2556,N_2933);
or U4924 (N_4924,N_2995,N_3119);
nand U4925 (N_4925,N_3441,N_2747);
nand U4926 (N_4926,N_2926,N_3364);
nor U4927 (N_4927,N_2931,N_2790);
or U4928 (N_4928,N_3190,N_3218);
xor U4929 (N_4929,N_2784,N_3731);
or U4930 (N_4930,N_3370,N_2892);
and U4931 (N_4931,N_3281,N_3013);
and U4932 (N_4932,N_3320,N_3535);
nor U4933 (N_4933,N_3006,N_3318);
nor U4934 (N_4934,N_3702,N_2818);
or U4935 (N_4935,N_3197,N_3357);
xor U4936 (N_4936,N_2727,N_3034);
and U4937 (N_4937,N_2615,N_3092);
nor U4938 (N_4938,N_2721,N_3257);
or U4939 (N_4939,N_3516,N_3076);
nor U4940 (N_4940,N_2742,N_2735);
and U4941 (N_4941,N_2554,N_3688);
nand U4942 (N_4942,N_3720,N_3684);
and U4943 (N_4943,N_3071,N_2839);
nor U4944 (N_4944,N_2913,N_3743);
or U4945 (N_4945,N_2519,N_2581);
or U4946 (N_4946,N_2718,N_3027);
or U4947 (N_4947,N_2565,N_2935);
and U4948 (N_4948,N_2789,N_3735);
nand U4949 (N_4949,N_3142,N_2987);
nand U4950 (N_4950,N_2948,N_2927);
nand U4951 (N_4951,N_3717,N_2519);
xnor U4952 (N_4952,N_3389,N_2808);
and U4953 (N_4953,N_3109,N_3121);
nor U4954 (N_4954,N_3699,N_3153);
xnor U4955 (N_4955,N_3575,N_3499);
nor U4956 (N_4956,N_3512,N_2643);
xor U4957 (N_4957,N_3530,N_2764);
or U4958 (N_4958,N_2548,N_2883);
xor U4959 (N_4959,N_2721,N_2634);
and U4960 (N_4960,N_2846,N_2678);
and U4961 (N_4961,N_2545,N_3446);
and U4962 (N_4962,N_3432,N_3295);
xnor U4963 (N_4963,N_3273,N_3691);
xnor U4964 (N_4964,N_3735,N_3145);
and U4965 (N_4965,N_2599,N_3339);
nor U4966 (N_4966,N_2860,N_3326);
nor U4967 (N_4967,N_3203,N_2768);
xor U4968 (N_4968,N_3556,N_2822);
and U4969 (N_4969,N_3477,N_3121);
or U4970 (N_4970,N_3013,N_2654);
nor U4971 (N_4971,N_3588,N_3129);
nor U4972 (N_4972,N_3536,N_3544);
nor U4973 (N_4973,N_3565,N_2684);
xnor U4974 (N_4974,N_3398,N_3543);
or U4975 (N_4975,N_3077,N_3704);
nand U4976 (N_4976,N_2893,N_2684);
xor U4977 (N_4977,N_2987,N_2665);
nand U4978 (N_4978,N_2541,N_3488);
xor U4979 (N_4979,N_3568,N_3706);
and U4980 (N_4980,N_3262,N_3727);
nand U4981 (N_4981,N_3676,N_3709);
nand U4982 (N_4982,N_3615,N_2769);
or U4983 (N_4983,N_2792,N_2747);
nand U4984 (N_4984,N_3401,N_3108);
nor U4985 (N_4985,N_2652,N_3404);
or U4986 (N_4986,N_3650,N_2806);
and U4987 (N_4987,N_3489,N_3658);
and U4988 (N_4988,N_3049,N_3386);
nor U4989 (N_4989,N_2552,N_2932);
nor U4990 (N_4990,N_3052,N_2686);
nand U4991 (N_4991,N_3366,N_3482);
or U4992 (N_4992,N_2723,N_3360);
nor U4993 (N_4993,N_3663,N_2791);
and U4994 (N_4994,N_3403,N_3590);
nand U4995 (N_4995,N_2945,N_2975);
xor U4996 (N_4996,N_3164,N_2690);
nor U4997 (N_4997,N_2559,N_2578);
nor U4998 (N_4998,N_2971,N_3120);
nor U4999 (N_4999,N_2584,N_3380);
nand U5000 (N_5000,N_4842,N_4156);
and U5001 (N_5001,N_4005,N_4825);
or U5002 (N_5002,N_3948,N_4903);
xnor U5003 (N_5003,N_4907,N_4951);
nor U5004 (N_5004,N_4760,N_4937);
and U5005 (N_5005,N_3924,N_4984);
xnor U5006 (N_5006,N_4302,N_4378);
or U5007 (N_5007,N_4839,N_4433);
nand U5008 (N_5008,N_4772,N_4536);
xnor U5009 (N_5009,N_4203,N_4813);
or U5010 (N_5010,N_4904,N_4961);
xor U5011 (N_5011,N_4475,N_4797);
nor U5012 (N_5012,N_4333,N_4351);
or U5013 (N_5013,N_4212,N_4502);
xnor U5014 (N_5014,N_4809,N_3910);
or U5015 (N_5015,N_4720,N_4017);
xor U5016 (N_5016,N_4528,N_4257);
nand U5017 (N_5017,N_4589,N_4299);
or U5018 (N_5018,N_3997,N_4316);
and U5019 (N_5019,N_4624,N_4294);
and U5020 (N_5020,N_4328,N_3994);
nand U5021 (N_5021,N_4312,N_4640);
and U5022 (N_5022,N_4140,N_4301);
nor U5023 (N_5023,N_3951,N_4417);
nand U5024 (N_5024,N_4777,N_3939);
nand U5025 (N_5025,N_4222,N_3870);
or U5026 (N_5026,N_4991,N_4785);
xnor U5027 (N_5027,N_4229,N_4437);
and U5028 (N_5028,N_4694,N_4572);
or U5029 (N_5029,N_4002,N_4943);
nor U5030 (N_5030,N_4710,N_4290);
and U5031 (N_5031,N_4373,N_4996);
and U5032 (N_5032,N_4662,N_4132);
xnor U5033 (N_5033,N_4912,N_3900);
xor U5034 (N_5034,N_4462,N_3841);
nand U5035 (N_5035,N_4269,N_4288);
or U5036 (N_5036,N_4563,N_4449);
nor U5037 (N_5037,N_4634,N_3821);
xnor U5038 (N_5038,N_4165,N_4040);
nand U5039 (N_5039,N_3979,N_3960);
nor U5040 (N_5040,N_4385,N_4239);
xnor U5041 (N_5041,N_3932,N_3944);
or U5042 (N_5042,N_4551,N_3856);
and U5043 (N_5043,N_4675,N_4224);
nor U5044 (N_5044,N_4711,N_4761);
or U5045 (N_5045,N_4603,N_4958);
and U5046 (N_5046,N_4013,N_4554);
and U5047 (N_5047,N_4338,N_4076);
xnor U5048 (N_5048,N_4493,N_4500);
and U5049 (N_5049,N_4564,N_3757);
nor U5050 (N_5050,N_4047,N_4235);
xnor U5051 (N_5051,N_4345,N_4916);
nand U5052 (N_5052,N_3969,N_4773);
nand U5053 (N_5053,N_4356,N_4410);
nand U5054 (N_5054,N_4108,N_4771);
nor U5055 (N_5055,N_4431,N_4159);
nor U5056 (N_5056,N_4866,N_4453);
or U5057 (N_5057,N_4786,N_4778);
and U5058 (N_5058,N_4104,N_4174);
and U5059 (N_5059,N_4464,N_4518);
xor U5060 (N_5060,N_4230,N_3965);
or U5061 (N_5061,N_4249,N_4890);
or U5062 (N_5062,N_4262,N_4731);
nand U5063 (N_5063,N_4689,N_4205);
nand U5064 (N_5064,N_4506,N_3785);
or U5065 (N_5065,N_3797,N_4256);
nand U5066 (N_5066,N_4261,N_4881);
nand U5067 (N_5067,N_4079,N_4178);
xor U5068 (N_5068,N_4319,N_3780);
nand U5069 (N_5069,N_3966,N_4549);
nor U5070 (N_5070,N_4401,N_3838);
nor U5071 (N_5071,N_3847,N_4614);
or U5072 (N_5072,N_4359,N_3971);
and U5073 (N_5073,N_4346,N_4483);
nor U5074 (N_5074,N_3929,N_4821);
nand U5075 (N_5075,N_3992,N_4255);
or U5076 (N_5076,N_4678,N_4807);
nand U5077 (N_5077,N_4781,N_4587);
and U5078 (N_5078,N_4664,N_4730);
or U5079 (N_5079,N_4643,N_4657);
nor U5080 (N_5080,N_3904,N_4562);
and U5081 (N_5081,N_4695,N_3831);
nor U5082 (N_5082,N_4962,N_4399);
xnor U5083 (N_5083,N_3915,N_4238);
nor U5084 (N_5084,N_4905,N_4154);
and U5085 (N_5085,N_4339,N_4194);
xor U5086 (N_5086,N_4295,N_4582);
or U5087 (N_5087,N_4846,N_4700);
xnor U5088 (N_5088,N_4116,N_4281);
and U5089 (N_5089,N_4292,N_4347);
nand U5090 (N_5090,N_4107,N_4880);
xnor U5091 (N_5091,N_4902,N_4086);
nor U5092 (N_5092,N_4136,N_4567);
xnor U5093 (N_5093,N_3921,N_4062);
xnor U5094 (N_5094,N_4161,N_4418);
nand U5095 (N_5095,N_4069,N_4800);
and U5096 (N_5096,N_4535,N_4382);
xor U5097 (N_5097,N_4066,N_3760);
nor U5098 (N_5098,N_3919,N_4114);
and U5099 (N_5099,N_4636,N_3923);
or U5100 (N_5100,N_3998,N_4323);
xor U5101 (N_5101,N_4539,N_4298);
nor U5102 (N_5102,N_4628,N_4920);
xor U5103 (N_5103,N_3893,N_4349);
and U5104 (N_5104,N_4598,N_3896);
xor U5105 (N_5105,N_4514,N_4758);
xnor U5106 (N_5106,N_4612,N_4503);
nor U5107 (N_5107,N_4621,N_3816);
nand U5108 (N_5108,N_4172,N_4847);
xnor U5109 (N_5109,N_4213,N_4888);
or U5110 (N_5110,N_3917,N_4420);
xor U5111 (N_5111,N_4123,N_4663);
nand U5112 (N_5112,N_4801,N_4548);
nand U5113 (N_5113,N_4595,N_4867);
nor U5114 (N_5114,N_4602,N_3782);
and U5115 (N_5115,N_4220,N_4364);
xnor U5116 (N_5116,N_3809,N_4638);
xnor U5117 (N_5117,N_4613,N_4189);
nor U5118 (N_5118,N_4181,N_4976);
nand U5119 (N_5119,N_4780,N_4811);
or U5120 (N_5120,N_4309,N_4436);
nor U5121 (N_5121,N_3943,N_4791);
and U5122 (N_5122,N_4163,N_4210);
or U5123 (N_5123,N_4980,N_4085);
nand U5124 (N_5124,N_3793,N_4990);
and U5125 (N_5125,N_4956,N_4673);
xnor U5126 (N_5126,N_4273,N_4470);
nor U5127 (N_5127,N_4241,N_4573);
nor U5128 (N_5128,N_4246,N_4885);
and U5129 (N_5129,N_4303,N_4666);
and U5130 (N_5130,N_4153,N_4358);
xnor U5131 (N_5131,N_4134,N_4726);
or U5132 (N_5132,N_4889,N_4147);
nor U5133 (N_5133,N_4537,N_4152);
xnor U5134 (N_5134,N_4626,N_4987);
xnor U5135 (N_5135,N_4073,N_3898);
nand U5136 (N_5136,N_4392,N_4995);
xor U5137 (N_5137,N_4327,N_4524);
or U5138 (N_5138,N_4361,N_3788);
nand U5139 (N_5139,N_4688,N_4275);
nor U5140 (N_5140,N_3887,N_4074);
and U5141 (N_5141,N_3810,N_4899);
nand U5142 (N_5142,N_3762,N_4856);
and U5143 (N_5143,N_4714,N_3974);
or U5144 (N_5144,N_4830,N_3753);
xnor U5145 (N_5145,N_4250,N_4787);
xnor U5146 (N_5146,N_3907,N_4950);
xor U5147 (N_5147,N_3769,N_3895);
or U5148 (N_5148,N_4057,N_4928);
and U5149 (N_5149,N_4739,N_4986);
xnor U5150 (N_5150,N_3854,N_4642);
and U5151 (N_5151,N_4735,N_4698);
nand U5152 (N_5152,N_4233,N_4372);
or U5153 (N_5153,N_4315,N_3763);
and U5154 (N_5154,N_4498,N_4578);
nor U5155 (N_5155,N_4287,N_4585);
or U5156 (N_5156,N_4941,N_3863);
nor U5157 (N_5157,N_3899,N_3869);
or U5158 (N_5158,N_4512,N_3937);
nor U5159 (N_5159,N_4182,N_4862);
or U5160 (N_5160,N_4874,N_4533);
xor U5161 (N_5161,N_4455,N_3891);
or U5162 (N_5162,N_4148,N_4124);
xor U5163 (N_5163,N_3912,N_4765);
xor U5164 (N_5164,N_4102,N_4266);
xnor U5165 (N_5165,N_4044,N_4425);
and U5166 (N_5166,N_4505,N_4769);
and U5167 (N_5167,N_3975,N_4305);
nor U5168 (N_5168,N_4690,N_4329);
xor U5169 (N_5169,N_4532,N_4314);
xor U5170 (N_5170,N_4805,N_4369);
xnor U5171 (N_5171,N_4764,N_3791);
and U5172 (N_5172,N_4463,N_4218);
or U5173 (N_5173,N_4403,N_4137);
nor U5174 (N_5174,N_4712,N_3866);
and U5175 (N_5175,N_4878,N_4783);
nor U5176 (N_5176,N_4041,N_4348);
nor U5177 (N_5177,N_4759,N_3968);
nor U5178 (N_5178,N_4820,N_3949);
nand U5179 (N_5179,N_4908,N_3787);
and U5180 (N_5180,N_3830,N_4571);
nand U5181 (N_5181,N_4402,N_4946);
nand U5182 (N_5182,N_4016,N_4831);
xnor U5183 (N_5183,N_4576,N_4383);
and U5184 (N_5184,N_4293,N_4701);
nor U5185 (N_5185,N_4193,N_4665);
nor U5186 (N_5186,N_4547,N_4183);
nand U5187 (N_5187,N_4419,N_4118);
nand U5188 (N_5188,N_4499,N_4604);
or U5189 (N_5189,N_4893,N_4196);
nor U5190 (N_5190,N_4489,N_4515);
nor U5191 (N_5191,N_4670,N_3964);
xnor U5192 (N_5192,N_4708,N_4414);
or U5193 (N_5193,N_3872,N_3967);
xnor U5194 (N_5194,N_3982,N_4009);
or U5195 (N_5195,N_3973,N_4597);
xnor U5196 (N_5196,N_4151,N_4072);
nor U5197 (N_5197,N_4226,N_3824);
xor U5198 (N_5198,N_4119,N_3773);
and U5199 (N_5199,N_4993,N_4396);
xor U5200 (N_5200,N_3882,N_4855);
nand U5201 (N_5201,N_4448,N_3772);
nand U5202 (N_5202,N_4947,N_4814);
and U5203 (N_5203,N_3999,N_4767);
or U5204 (N_5204,N_3796,N_3852);
and U5205 (N_5205,N_4812,N_4077);
nand U5206 (N_5206,N_4723,N_4858);
or U5207 (N_5207,N_4185,N_4482);
nor U5208 (N_5208,N_4051,N_4426);
nand U5209 (N_5209,N_4468,N_4265);
nand U5210 (N_5210,N_4342,N_3859);
or U5211 (N_5211,N_4798,N_4929);
or U5212 (N_5212,N_4353,N_4952);
nor U5213 (N_5213,N_4741,N_4616);
nand U5214 (N_5214,N_3873,N_4087);
xnor U5215 (N_5215,N_4822,N_4629);
nor U5216 (N_5216,N_4432,N_4439);
nand U5217 (N_5217,N_4718,N_4924);
xnor U5218 (N_5218,N_4596,N_4452);
nand U5219 (N_5219,N_3795,N_4003);
nor U5220 (N_5220,N_3800,N_4763);
or U5221 (N_5221,N_4627,N_3835);
and U5222 (N_5222,N_4917,N_4456);
nand U5223 (N_5223,N_4094,N_4721);
xor U5224 (N_5224,N_4579,N_4744);
xor U5225 (N_5225,N_4569,N_4216);
xnor U5226 (N_5226,N_4451,N_4538);
nor U5227 (N_5227,N_4560,N_3799);
or U5228 (N_5228,N_3851,N_4803);
nand U5229 (N_5229,N_4474,N_4651);
xor U5230 (N_5230,N_4860,N_4715);
xor U5231 (N_5231,N_4817,N_4367);
or U5232 (N_5232,N_4509,N_4750);
nand U5233 (N_5233,N_4975,N_4208);
xor U5234 (N_5234,N_4092,N_4245);
nor U5235 (N_5235,N_4001,N_3826);
and U5236 (N_5236,N_4555,N_4832);
or U5237 (N_5237,N_3892,N_4055);
and U5238 (N_5238,N_4519,N_4479);
and U5239 (N_5239,N_3993,N_4306);
xnor U5240 (N_5240,N_4891,N_4697);
nor U5241 (N_5241,N_4829,N_4411);
nand U5242 (N_5242,N_4160,N_3876);
nor U5243 (N_5243,N_4511,N_4901);
and U5244 (N_5244,N_4240,N_4979);
nor U5245 (N_5245,N_4459,N_4054);
xnor U5246 (N_5246,N_4490,N_4125);
nand U5247 (N_5247,N_4209,N_3933);
and U5248 (N_5248,N_4552,N_4836);
nand U5249 (N_5249,N_4387,N_4093);
nor U5250 (N_5250,N_4989,N_4611);
xnor U5251 (N_5251,N_4206,N_4960);
xnor U5252 (N_5252,N_4162,N_3767);
nor U5253 (N_5253,N_3931,N_4157);
xnor U5254 (N_5254,N_4258,N_4486);
nor U5255 (N_5255,N_4244,N_4816);
xnor U5256 (N_5256,N_4601,N_3885);
nand U5257 (N_5257,N_4752,N_4215);
nor U5258 (N_5258,N_4313,N_4211);
xnor U5259 (N_5259,N_4794,N_4408);
or U5260 (N_5260,N_4592,N_4869);
or U5261 (N_5261,N_3776,N_3991);
or U5262 (N_5262,N_4568,N_4248);
xnor U5263 (N_5263,N_4179,N_3811);
xor U5264 (N_5264,N_4913,N_4749);
nor U5265 (N_5265,N_4610,N_3930);
nor U5266 (N_5266,N_4757,N_4296);
nor U5267 (N_5267,N_4412,N_4792);
nor U5268 (N_5268,N_3976,N_4930);
and U5269 (N_5269,N_3777,N_4068);
nor U5270 (N_5270,N_4450,N_4932);
and U5271 (N_5271,N_3823,N_4007);
nand U5272 (N_5272,N_4308,N_4440);
or U5273 (N_5273,N_4877,N_3812);
or U5274 (N_5274,N_4268,N_4438);
xnor U5275 (N_5275,N_4404,N_4921);
or U5276 (N_5276,N_4070,N_4082);
and U5277 (N_5277,N_4546,N_4191);
and U5278 (N_5278,N_4755,N_4310);
xnor U5279 (N_5279,N_4897,N_4078);
or U5280 (N_5280,N_4472,N_4398);
nand U5281 (N_5281,N_3759,N_4925);
and U5282 (N_5282,N_3750,N_4898);
nand U5283 (N_5283,N_4659,N_4553);
xor U5284 (N_5284,N_4034,N_4982);
and U5285 (N_5285,N_4588,N_3985);
and U5286 (N_5286,N_3954,N_4168);
nand U5287 (N_5287,N_4127,N_4672);
xnor U5288 (N_5288,N_4445,N_4335);
and U5289 (N_5289,N_4045,N_3828);
xnor U5290 (N_5290,N_4321,N_4059);
or U5291 (N_5291,N_4198,N_4635);
nor U5292 (N_5292,N_4868,N_4705);
nand U5293 (N_5293,N_4032,N_4377);
or U5294 (N_5294,N_4594,N_3756);
nor U5295 (N_5295,N_4743,N_4325);
xor U5296 (N_5296,N_4722,N_4819);
xor U5297 (N_5297,N_4593,N_3978);
nor U5298 (N_5298,N_3990,N_4103);
and U5299 (N_5299,N_4969,N_4128);
or U5300 (N_5300,N_3765,N_4095);
nor U5301 (N_5301,N_4927,N_3857);
and U5302 (N_5302,N_4391,N_4828);
nor U5303 (N_5303,N_4331,N_3947);
xnor U5304 (N_5304,N_4677,N_3807);
and U5305 (N_5305,N_4326,N_3906);
xnor U5306 (N_5306,N_3911,N_4130);
and U5307 (N_5307,N_4894,N_4607);
and U5308 (N_5308,N_4175,N_4379);
xnor U5309 (N_5309,N_3958,N_4609);
nor U5310 (N_5310,N_3996,N_4716);
nor U5311 (N_5311,N_4135,N_3995);
or U5312 (N_5312,N_3981,N_3842);
nor U5313 (N_5313,N_4854,N_3903);
nor U5314 (N_5314,N_4129,N_4618);
xnor U5315 (N_5315,N_4530,N_3935);
xor U5316 (N_5316,N_3956,N_3774);
xnor U5317 (N_5317,N_3813,N_4071);
or U5318 (N_5318,N_4740,N_4354);
nor U5319 (N_5319,N_4802,N_4606);
or U5320 (N_5320,N_3846,N_4967);
nand U5321 (N_5321,N_4038,N_4466);
or U5322 (N_5322,N_4138,N_4696);
or U5323 (N_5323,N_4823,N_3789);
xnor U5324 (N_5324,N_3945,N_3865);
and U5325 (N_5325,N_4409,N_3920);
or U5326 (N_5326,N_4766,N_4075);
or U5327 (N_5327,N_4746,N_4232);
xnor U5328 (N_5328,N_4337,N_3881);
nor U5329 (N_5329,N_4388,N_4729);
nand U5330 (N_5330,N_3934,N_4341);
and U5331 (N_5331,N_4442,N_3875);
or U5332 (N_5332,N_4652,N_4944);
nor U5333 (N_5333,N_4285,N_3980);
xor U5334 (N_5334,N_4632,N_4622);
xnor U5335 (N_5335,N_3905,N_3808);
xnor U5336 (N_5336,N_4520,N_4260);
or U5337 (N_5337,N_4375,N_3853);
nor U5338 (N_5338,N_4838,N_4141);
xor U5339 (N_5339,N_3784,N_3849);
nand U5340 (N_5340,N_4926,N_4365);
nand U5341 (N_5341,N_4340,N_4747);
nand U5342 (N_5342,N_4030,N_4671);
xnor U5343 (N_5343,N_3794,N_3890);
or U5344 (N_5344,N_4692,N_4434);
nor U5345 (N_5345,N_4155,N_4166);
or U5346 (N_5346,N_4574,N_4906);
nor U5347 (N_5347,N_4983,N_4397);
nand U5348 (N_5348,N_4895,N_3833);
or U5349 (N_5349,N_4501,N_3805);
and U5350 (N_5350,N_4097,N_4406);
nor U5351 (N_5351,N_4279,N_4035);
nor U5352 (N_5352,N_4717,N_4237);
xor U5353 (N_5353,N_4217,N_4080);
and U5354 (N_5354,N_4413,N_4173);
and U5355 (N_5355,N_4922,N_4355);
and U5356 (N_5356,N_4117,N_4508);
nand U5357 (N_5357,N_3860,N_4150);
and U5358 (N_5358,N_3926,N_4542);
or U5359 (N_5359,N_4557,N_3972);
or U5360 (N_5360,N_4940,N_3977);
or U5361 (N_5361,N_4732,N_4344);
or U5362 (N_5362,N_3755,N_4586);
xnor U5363 (N_5363,N_4972,N_4892);
xnor U5364 (N_5364,N_4158,N_4971);
or U5365 (N_5365,N_3804,N_4872);
nor U5366 (N_5366,N_4177,N_4541);
and U5367 (N_5367,N_4201,N_4186);
nand U5368 (N_5368,N_4565,N_3751);
xnor U5369 (N_5369,N_4703,N_4471);
nor U5370 (N_5370,N_4476,N_4029);
xnor U5371 (N_5371,N_4371,N_3874);
xnor U5372 (N_5372,N_4407,N_4048);
and U5373 (N_5373,N_4039,N_4142);
xor U5374 (N_5374,N_4775,N_4488);
xnor U5375 (N_5375,N_4790,N_4283);
nor U5376 (N_5376,N_4865,N_4204);
xnor U5377 (N_5377,N_3959,N_3902);
and U5378 (N_5378,N_4352,N_4648);
and U5379 (N_5379,N_3983,N_4014);
nand U5380 (N_5380,N_4247,N_3850);
nor U5381 (N_5381,N_4254,N_4376);
nand U5382 (N_5382,N_4133,N_4728);
xor U5383 (N_5383,N_3832,N_4599);
nor U5384 (N_5384,N_4522,N_4873);
nand U5385 (N_5385,N_4774,N_4768);
nand U5386 (N_5386,N_3840,N_4112);
or U5387 (N_5387,N_4496,N_4687);
or U5388 (N_5388,N_3908,N_3825);
nor U5389 (N_5389,N_4473,N_4144);
xnor U5390 (N_5390,N_4707,N_4581);
and U5391 (N_5391,N_4973,N_4046);
xor U5392 (N_5392,N_4540,N_3962);
xor U5393 (N_5393,N_4953,N_4970);
nand U5394 (N_5394,N_3819,N_4487);
nor U5395 (N_5395,N_4655,N_4997);
nand U5396 (N_5396,N_3839,N_4200);
xnor U5397 (N_5397,N_3986,N_4264);
xor U5398 (N_5398,N_4639,N_4422);
nor U5399 (N_5399,N_4837,N_3758);
or U5400 (N_5400,N_4111,N_3889);
nand U5401 (N_5401,N_4458,N_4004);
xor U5402 (N_5402,N_4966,N_4745);
nand U5403 (N_5403,N_3942,N_4024);
or U5404 (N_5404,N_4988,N_4526);
nor U5405 (N_5405,N_4608,N_4948);
and U5406 (N_5406,N_4336,N_4693);
or U5407 (N_5407,N_4738,N_4042);
or U5408 (N_5408,N_4242,N_3761);
nor U5409 (N_5409,N_4400,N_4497);
or U5410 (N_5410,N_4390,N_3922);
nor U5411 (N_5411,N_4274,N_4938);
nand U5412 (N_5412,N_4291,N_3775);
or U5413 (N_5413,N_4019,N_3927);
xnor U5414 (N_5414,N_4699,N_3768);
xnor U5415 (N_5415,N_4060,N_4637);
nor U5416 (N_5416,N_4793,N_4380);
nand U5417 (N_5417,N_4277,N_4911);
nor U5418 (N_5418,N_4423,N_4334);
and U5419 (N_5419,N_4859,N_4619);
nor U5420 (N_5420,N_4089,N_4806);
or U5421 (N_5421,N_4214,N_3855);
nand U5422 (N_5422,N_4110,N_4685);
xnor U5423 (N_5423,N_4478,N_4507);
or U5424 (N_5424,N_4919,N_4650);
and U5425 (N_5425,N_4441,N_4504);
or U5426 (N_5426,N_3770,N_4884);
nor U5427 (N_5427,N_4307,N_4968);
nand U5428 (N_5428,N_3878,N_4827);
nand U5429 (N_5429,N_3883,N_4799);
xor U5430 (N_5430,N_4228,N_4756);
and U5431 (N_5431,N_3901,N_4343);
xnor U5432 (N_5432,N_4605,N_4864);
nor U5433 (N_5433,N_4416,N_4225);
and U5434 (N_5434,N_4556,N_4949);
nand U5435 (N_5435,N_4955,N_4709);
nor U5436 (N_5436,N_4580,N_4320);
xnor U5437 (N_5437,N_4282,N_4570);
and U5438 (N_5438,N_4465,N_4770);
xnor U5439 (N_5439,N_4143,N_3848);
nor U5440 (N_5440,N_4415,N_4188);
xnor U5441 (N_5441,N_4053,N_4681);
nor U5442 (N_5442,N_3963,N_4513);
or U5443 (N_5443,N_4366,N_4914);
and U5444 (N_5444,N_4534,N_4485);
or U5445 (N_5445,N_4600,N_3928);
and U5446 (N_5446,N_4481,N_4886);
nor U5447 (N_5447,N_4959,N_4835);
nand U5448 (N_5448,N_3867,N_4167);
and U5449 (N_5449,N_4495,N_3864);
or U5450 (N_5450,N_4936,N_4028);
nor U5451 (N_5451,N_4405,N_3888);
or U5452 (N_5452,N_3834,N_4527);
nor U5453 (N_5453,N_4945,N_4317);
nand U5454 (N_5454,N_4063,N_4427);
xor U5455 (N_5455,N_4357,N_4272);
and U5456 (N_5456,N_4789,N_3837);
nand U5457 (N_5457,N_4558,N_4667);
nand U5458 (N_5458,N_4942,N_3814);
xor U5459 (N_5459,N_4724,N_3766);
and U5460 (N_5460,N_4680,N_4682);
xor U5461 (N_5461,N_4559,N_3916);
xnor U5462 (N_5462,N_4978,N_4683);
and U5463 (N_5463,N_4644,N_3806);
and U5464 (N_5464,N_3792,N_4737);
nand U5465 (N_5465,N_4067,N_4202);
nor U5466 (N_5466,N_3946,N_4126);
xnor U5467 (N_5467,N_4840,N_4516);
nand U5468 (N_5468,N_4957,N_4645);
and U5469 (N_5469,N_4311,N_4430);
or U5470 (N_5470,N_4517,N_4289);
and U5471 (N_5471,N_3802,N_4469);
or U5472 (N_5472,N_3925,N_4023);
and U5473 (N_5473,N_4615,N_3941);
and U5474 (N_5474,N_4088,N_4467);
or U5475 (N_5475,N_4259,N_4727);
nand U5476 (N_5476,N_4583,N_4460);
nand U5477 (N_5477,N_4871,N_4050);
or U5478 (N_5478,N_4020,N_4243);
and U5479 (N_5479,N_4139,N_4849);
or U5480 (N_5480,N_4625,N_4751);
nor U5481 (N_5481,N_4036,N_4852);
and U5482 (N_5482,N_4098,N_4368);
and U5483 (N_5483,N_4857,N_4706);
nor U5484 (N_5484,N_4918,N_4815);
xor U5485 (N_5485,N_4454,N_4954);
xnor U5486 (N_5486,N_4389,N_4617);
xor U5487 (N_5487,N_4974,N_4253);
and U5488 (N_5488,N_4545,N_4525);
nand U5489 (N_5489,N_4845,N_4018);
nand U5490 (N_5490,N_3771,N_4641);
nor U5491 (N_5491,N_4101,N_4896);
and U5492 (N_5492,N_4330,N_3940);
and U5493 (N_5493,N_4804,N_3779);
nand U5494 (N_5494,N_4934,N_4236);
nand U5495 (N_5495,N_4736,N_4145);
and U5496 (N_5496,N_4171,N_4457);
nand U5497 (N_5497,N_3820,N_4011);
and U5498 (N_5498,N_4360,N_3952);
nor U5499 (N_5499,N_4684,N_3897);
nor U5500 (N_5500,N_4267,N_4844);
and U5501 (N_5501,N_4850,N_4350);
xor U5502 (N_5502,N_4853,N_4049);
or U5503 (N_5503,N_4106,N_4480);
nand U5504 (N_5504,N_4964,N_4221);
nand U5505 (N_5505,N_4491,N_4753);
nor U5506 (N_5506,N_4297,N_3836);
and U5507 (N_5507,N_4170,N_4748);
xor U5508 (N_5508,N_3886,N_4362);
or U5509 (N_5509,N_3909,N_4674);
xor U5510 (N_5510,N_3987,N_4381);
nand U5511 (N_5511,N_4105,N_4660);
xor U5512 (N_5512,N_4661,N_4649);
xor U5513 (N_5513,N_4719,N_4164);
or U5514 (N_5514,N_4795,N_4374);
and U5515 (N_5515,N_4000,N_3845);
and U5516 (N_5516,N_4447,N_4190);
and U5517 (N_5517,N_4861,N_4529);
and U5518 (N_5518,N_4271,N_3798);
or U5519 (N_5519,N_4192,N_4064);
nor U5520 (N_5520,N_4833,N_4015);
nand U5521 (N_5521,N_4676,N_4494);
or U5522 (N_5522,N_4394,N_3790);
nor U5523 (N_5523,N_4318,N_3871);
nand U5524 (N_5524,N_4061,N_3880);
and U5525 (N_5525,N_3781,N_4931);
nand U5526 (N_5526,N_3877,N_4824);
xnor U5527 (N_5527,N_4591,N_4848);
xor U5528 (N_5528,N_4056,N_4841);
nand U5529 (N_5529,N_4779,N_4115);
xnor U5530 (N_5530,N_3822,N_4006);
and U5531 (N_5531,N_4742,N_3957);
nand U5532 (N_5532,N_4733,N_3817);
nor U5533 (N_5533,N_4923,N_3914);
nor U5534 (N_5534,N_3970,N_4304);
nand U5535 (N_5535,N_4584,N_4590);
xor U5536 (N_5536,N_3858,N_4395);
or U5537 (N_5537,N_3803,N_4882);
nand U5538 (N_5538,N_4184,N_4484);
xor U5539 (N_5539,N_4630,N_4084);
xor U5540 (N_5540,N_3988,N_4322);
nor U5541 (N_5541,N_3862,N_4421);
and U5542 (N_5542,N_4083,N_4669);
nand U5543 (N_5543,N_3989,N_4754);
nand U5544 (N_5544,N_4096,N_4843);
or U5545 (N_5545,N_4531,N_4025);
or U5546 (N_5546,N_4909,N_4252);
xor U5547 (N_5547,N_4052,N_4713);
nor U5548 (N_5548,N_4900,N_4021);
and U5549 (N_5549,N_4550,N_4037);
nor U5550 (N_5550,N_4725,N_4444);
nor U5551 (N_5551,N_3754,N_4492);
nand U5552 (N_5552,N_4324,N_3936);
and U5553 (N_5553,N_4782,N_4027);
or U5554 (N_5554,N_4818,N_4656);
or U5555 (N_5555,N_3843,N_4734);
xnor U5556 (N_5556,N_4620,N_4278);
xor U5557 (N_5557,N_3818,N_4300);
xor U5558 (N_5558,N_4965,N_4543);
and U5559 (N_5559,N_4653,N_4424);
and U5560 (N_5560,N_4477,N_4933);
or U5561 (N_5561,N_4704,N_4384);
xor U5562 (N_5562,N_4131,N_4031);
xor U5563 (N_5563,N_4658,N_4981);
and U5564 (N_5564,N_4654,N_4363);
nor U5565 (N_5565,N_4043,N_3764);
and U5566 (N_5566,N_3879,N_4234);
or U5567 (N_5567,N_4523,N_4810);
or U5568 (N_5568,N_4702,N_4910);
and U5569 (N_5569,N_4879,N_4691);
xor U5570 (N_5570,N_3786,N_4090);
xnor U5571 (N_5571,N_4149,N_4646);
and U5572 (N_5572,N_4270,N_4808);
nor U5573 (N_5573,N_3938,N_4561);
or U5574 (N_5574,N_3783,N_4826);
or U5575 (N_5575,N_4994,N_4109);
or U5576 (N_5576,N_4686,N_4939);
nand U5577 (N_5577,N_4197,N_4461);
and U5578 (N_5578,N_3801,N_4146);
or U5579 (N_5579,N_4010,N_4985);
and U5580 (N_5580,N_3894,N_4386);
or U5581 (N_5581,N_3918,N_4446);
nor U5582 (N_5582,N_4963,N_4577);
and U5583 (N_5583,N_4195,N_4679);
and U5584 (N_5584,N_4834,N_4863);
or U5585 (N_5585,N_4370,N_4207);
nand U5586 (N_5586,N_3955,N_4219);
xnor U5587 (N_5587,N_4199,N_3961);
nand U5588 (N_5588,N_3844,N_3778);
nand U5589 (N_5589,N_4113,N_4876);
and U5590 (N_5590,N_4544,N_4796);
and U5591 (N_5591,N_4875,N_4633);
or U5592 (N_5592,N_4393,N_4058);
xnor U5593 (N_5593,N_4915,N_4223);
xor U5594 (N_5594,N_4231,N_4120);
nor U5595 (N_5595,N_3913,N_3752);
nor U5596 (N_5596,N_3884,N_4977);
and U5597 (N_5597,N_4566,N_4121);
or U5598 (N_5598,N_4180,N_4081);
and U5599 (N_5599,N_4091,N_4870);
nand U5600 (N_5600,N_4251,N_4762);
xor U5601 (N_5601,N_4647,N_4999);
and U5602 (N_5602,N_4263,N_4033);
xnor U5603 (N_5603,N_3829,N_4443);
nor U5604 (N_5604,N_4099,N_4286);
nor U5605 (N_5605,N_4883,N_4776);
nand U5606 (N_5606,N_3984,N_4276);
xnor U5607 (N_5607,N_4187,N_4575);
nor U5608 (N_5608,N_4280,N_4429);
and U5609 (N_5609,N_4851,N_3868);
nor U5610 (N_5610,N_3827,N_3815);
and U5611 (N_5611,N_4122,N_4026);
xnor U5612 (N_5612,N_3953,N_4935);
xor U5613 (N_5613,N_4998,N_4428);
and U5614 (N_5614,N_4784,N_4631);
and U5615 (N_5615,N_3861,N_4065);
and U5616 (N_5616,N_4284,N_4012);
nor U5617 (N_5617,N_4992,N_4668);
xnor U5618 (N_5618,N_4008,N_4887);
xor U5619 (N_5619,N_3950,N_4435);
nand U5620 (N_5620,N_4510,N_4788);
nor U5621 (N_5621,N_4521,N_4100);
nor U5622 (N_5622,N_4022,N_4623);
or U5623 (N_5623,N_4332,N_4227);
or U5624 (N_5624,N_4176,N_4169);
nor U5625 (N_5625,N_4912,N_4927);
nand U5626 (N_5626,N_4161,N_4337);
nor U5627 (N_5627,N_4949,N_4607);
xor U5628 (N_5628,N_4553,N_4531);
and U5629 (N_5629,N_4546,N_4157);
nand U5630 (N_5630,N_4206,N_4089);
xnor U5631 (N_5631,N_4747,N_4644);
nand U5632 (N_5632,N_3753,N_3782);
nor U5633 (N_5633,N_4512,N_4731);
nor U5634 (N_5634,N_4630,N_4952);
and U5635 (N_5635,N_4921,N_4426);
xor U5636 (N_5636,N_4820,N_4023);
nor U5637 (N_5637,N_4883,N_4131);
or U5638 (N_5638,N_4964,N_4880);
nand U5639 (N_5639,N_4077,N_4630);
and U5640 (N_5640,N_3819,N_4320);
nand U5641 (N_5641,N_4763,N_4793);
nand U5642 (N_5642,N_4873,N_4634);
xnor U5643 (N_5643,N_4615,N_3794);
nor U5644 (N_5644,N_4768,N_3773);
xor U5645 (N_5645,N_4857,N_4340);
nand U5646 (N_5646,N_4409,N_4094);
and U5647 (N_5647,N_4589,N_4612);
and U5648 (N_5648,N_4471,N_4031);
nor U5649 (N_5649,N_3795,N_4573);
xnor U5650 (N_5650,N_4650,N_4283);
or U5651 (N_5651,N_4064,N_4448);
xnor U5652 (N_5652,N_4398,N_4180);
xor U5653 (N_5653,N_3757,N_3790);
and U5654 (N_5654,N_4577,N_3815);
or U5655 (N_5655,N_3839,N_4154);
xor U5656 (N_5656,N_3859,N_4743);
and U5657 (N_5657,N_4690,N_4055);
or U5658 (N_5658,N_4157,N_4642);
or U5659 (N_5659,N_3956,N_4951);
or U5660 (N_5660,N_4174,N_4195);
xor U5661 (N_5661,N_4008,N_4883);
nor U5662 (N_5662,N_4651,N_4118);
and U5663 (N_5663,N_4192,N_3942);
xor U5664 (N_5664,N_4311,N_4579);
nor U5665 (N_5665,N_4581,N_4443);
or U5666 (N_5666,N_4576,N_4253);
nor U5667 (N_5667,N_4942,N_4919);
or U5668 (N_5668,N_4012,N_4721);
xnor U5669 (N_5669,N_3758,N_3887);
xnor U5670 (N_5670,N_4297,N_4506);
and U5671 (N_5671,N_4097,N_4330);
nor U5672 (N_5672,N_4379,N_4691);
and U5673 (N_5673,N_4731,N_4689);
or U5674 (N_5674,N_3752,N_4589);
nor U5675 (N_5675,N_4408,N_4927);
or U5676 (N_5676,N_4816,N_4588);
xor U5677 (N_5677,N_4067,N_4293);
nor U5678 (N_5678,N_4696,N_4091);
or U5679 (N_5679,N_4739,N_3759);
nor U5680 (N_5680,N_4542,N_4900);
or U5681 (N_5681,N_3832,N_4984);
or U5682 (N_5682,N_4427,N_4841);
and U5683 (N_5683,N_4439,N_4031);
nand U5684 (N_5684,N_4950,N_4492);
and U5685 (N_5685,N_4452,N_4211);
and U5686 (N_5686,N_4133,N_4175);
nand U5687 (N_5687,N_4327,N_3897);
nor U5688 (N_5688,N_4251,N_4037);
xnor U5689 (N_5689,N_4400,N_4525);
nor U5690 (N_5690,N_4688,N_4225);
nor U5691 (N_5691,N_4297,N_4899);
xor U5692 (N_5692,N_4521,N_4829);
nand U5693 (N_5693,N_3886,N_4060);
or U5694 (N_5694,N_4261,N_4429);
nand U5695 (N_5695,N_4565,N_4474);
and U5696 (N_5696,N_4486,N_4976);
nand U5697 (N_5697,N_3964,N_4343);
or U5698 (N_5698,N_4304,N_4651);
xor U5699 (N_5699,N_4937,N_4110);
and U5700 (N_5700,N_4986,N_4115);
and U5701 (N_5701,N_3854,N_4553);
xor U5702 (N_5702,N_4158,N_4443);
nor U5703 (N_5703,N_4341,N_4817);
and U5704 (N_5704,N_4259,N_4251);
and U5705 (N_5705,N_4154,N_4443);
nand U5706 (N_5706,N_4414,N_4584);
nand U5707 (N_5707,N_3780,N_4553);
nor U5708 (N_5708,N_3751,N_4913);
nor U5709 (N_5709,N_4622,N_4141);
nand U5710 (N_5710,N_3973,N_4070);
xor U5711 (N_5711,N_4047,N_4035);
xnor U5712 (N_5712,N_4354,N_4716);
and U5713 (N_5713,N_4647,N_3762);
nand U5714 (N_5714,N_4779,N_4638);
nor U5715 (N_5715,N_4335,N_4492);
or U5716 (N_5716,N_4037,N_4291);
and U5717 (N_5717,N_4737,N_4261);
nor U5718 (N_5718,N_4248,N_4265);
and U5719 (N_5719,N_4754,N_3947);
nand U5720 (N_5720,N_3827,N_4439);
nand U5721 (N_5721,N_4253,N_4656);
and U5722 (N_5722,N_4533,N_4733);
and U5723 (N_5723,N_3752,N_4962);
nor U5724 (N_5724,N_4091,N_4129);
xor U5725 (N_5725,N_4011,N_4930);
nand U5726 (N_5726,N_4809,N_4475);
nand U5727 (N_5727,N_4343,N_3894);
and U5728 (N_5728,N_4272,N_4325);
and U5729 (N_5729,N_3944,N_4211);
or U5730 (N_5730,N_4801,N_4662);
nor U5731 (N_5731,N_4230,N_4394);
nand U5732 (N_5732,N_4768,N_4675);
or U5733 (N_5733,N_4024,N_4199);
and U5734 (N_5734,N_4319,N_4757);
nand U5735 (N_5735,N_3972,N_4459);
nor U5736 (N_5736,N_4071,N_4716);
and U5737 (N_5737,N_4942,N_4990);
xor U5738 (N_5738,N_4359,N_4366);
and U5739 (N_5739,N_4558,N_3770);
nor U5740 (N_5740,N_3993,N_4264);
and U5741 (N_5741,N_4135,N_4049);
nor U5742 (N_5742,N_3959,N_4990);
nor U5743 (N_5743,N_3839,N_4708);
nand U5744 (N_5744,N_4097,N_4554);
xnor U5745 (N_5745,N_4333,N_4629);
nand U5746 (N_5746,N_4054,N_4991);
nand U5747 (N_5747,N_4835,N_4193);
nand U5748 (N_5748,N_4645,N_4924);
and U5749 (N_5749,N_3881,N_4499);
and U5750 (N_5750,N_4201,N_4173);
xnor U5751 (N_5751,N_4203,N_4652);
nor U5752 (N_5752,N_3829,N_4488);
nor U5753 (N_5753,N_4400,N_4987);
nand U5754 (N_5754,N_4827,N_4433);
xor U5755 (N_5755,N_4545,N_4629);
and U5756 (N_5756,N_4220,N_4458);
xor U5757 (N_5757,N_4446,N_4420);
or U5758 (N_5758,N_3894,N_4340);
nand U5759 (N_5759,N_4174,N_4473);
nor U5760 (N_5760,N_4489,N_4181);
xor U5761 (N_5761,N_4026,N_4003);
nor U5762 (N_5762,N_4293,N_4182);
xor U5763 (N_5763,N_4548,N_4923);
nand U5764 (N_5764,N_3812,N_4106);
nand U5765 (N_5765,N_4208,N_4227);
nand U5766 (N_5766,N_4305,N_4605);
xnor U5767 (N_5767,N_4824,N_4985);
nor U5768 (N_5768,N_3905,N_4678);
and U5769 (N_5769,N_4420,N_4786);
or U5770 (N_5770,N_4538,N_4249);
nor U5771 (N_5771,N_4445,N_4508);
and U5772 (N_5772,N_4024,N_4093);
nor U5773 (N_5773,N_4654,N_3774);
nand U5774 (N_5774,N_4083,N_4832);
nand U5775 (N_5775,N_4394,N_4350);
nand U5776 (N_5776,N_4429,N_4986);
and U5777 (N_5777,N_4711,N_4385);
or U5778 (N_5778,N_4439,N_4484);
and U5779 (N_5779,N_4209,N_4454);
or U5780 (N_5780,N_4293,N_4454);
nand U5781 (N_5781,N_4458,N_4093);
nor U5782 (N_5782,N_3846,N_3828);
nor U5783 (N_5783,N_4556,N_3783);
or U5784 (N_5784,N_3849,N_4832);
nor U5785 (N_5785,N_4178,N_3806);
xnor U5786 (N_5786,N_4115,N_4551);
nand U5787 (N_5787,N_4831,N_4169);
nor U5788 (N_5788,N_4767,N_4918);
xnor U5789 (N_5789,N_3985,N_3802);
and U5790 (N_5790,N_4477,N_3766);
xor U5791 (N_5791,N_3880,N_4196);
xnor U5792 (N_5792,N_4272,N_4647);
and U5793 (N_5793,N_4989,N_3759);
and U5794 (N_5794,N_3909,N_3928);
and U5795 (N_5795,N_4034,N_4459);
nand U5796 (N_5796,N_4899,N_3786);
or U5797 (N_5797,N_4984,N_4837);
nand U5798 (N_5798,N_4036,N_4161);
xor U5799 (N_5799,N_4711,N_4489);
nand U5800 (N_5800,N_4707,N_3945);
or U5801 (N_5801,N_4854,N_4855);
or U5802 (N_5802,N_3968,N_4863);
and U5803 (N_5803,N_4238,N_3964);
xnor U5804 (N_5804,N_4733,N_4017);
xnor U5805 (N_5805,N_4495,N_4354);
or U5806 (N_5806,N_4934,N_4983);
or U5807 (N_5807,N_3938,N_4112);
nor U5808 (N_5808,N_4616,N_3825);
nor U5809 (N_5809,N_4827,N_4643);
xor U5810 (N_5810,N_4211,N_3828);
or U5811 (N_5811,N_4514,N_4367);
xor U5812 (N_5812,N_3941,N_4101);
xor U5813 (N_5813,N_4219,N_4414);
or U5814 (N_5814,N_4649,N_4371);
xor U5815 (N_5815,N_4996,N_4386);
or U5816 (N_5816,N_4534,N_3906);
nor U5817 (N_5817,N_4691,N_4684);
and U5818 (N_5818,N_4466,N_4368);
or U5819 (N_5819,N_4499,N_4715);
nor U5820 (N_5820,N_4956,N_3780);
or U5821 (N_5821,N_4229,N_3901);
nand U5822 (N_5822,N_4683,N_4202);
and U5823 (N_5823,N_4700,N_3771);
nor U5824 (N_5824,N_4410,N_4919);
nor U5825 (N_5825,N_4980,N_4613);
or U5826 (N_5826,N_4635,N_4831);
nand U5827 (N_5827,N_4806,N_4018);
xor U5828 (N_5828,N_4275,N_4570);
xnor U5829 (N_5829,N_4657,N_4434);
nand U5830 (N_5830,N_4659,N_3912);
or U5831 (N_5831,N_4697,N_4209);
or U5832 (N_5832,N_4665,N_4880);
nor U5833 (N_5833,N_3893,N_3937);
nor U5834 (N_5834,N_4236,N_4704);
nand U5835 (N_5835,N_4354,N_4985);
and U5836 (N_5836,N_4721,N_4789);
or U5837 (N_5837,N_4764,N_4904);
and U5838 (N_5838,N_4778,N_4379);
and U5839 (N_5839,N_3922,N_4232);
or U5840 (N_5840,N_4300,N_3929);
nor U5841 (N_5841,N_4231,N_4823);
xnor U5842 (N_5842,N_4590,N_4866);
xor U5843 (N_5843,N_4737,N_4340);
xnor U5844 (N_5844,N_4411,N_4054);
nor U5845 (N_5845,N_4285,N_4715);
nor U5846 (N_5846,N_4007,N_4829);
nor U5847 (N_5847,N_4564,N_3929);
or U5848 (N_5848,N_4571,N_4149);
nor U5849 (N_5849,N_4957,N_4625);
xor U5850 (N_5850,N_4010,N_4608);
xor U5851 (N_5851,N_4948,N_3963);
xnor U5852 (N_5852,N_4901,N_3911);
nand U5853 (N_5853,N_4319,N_4253);
nand U5854 (N_5854,N_4575,N_4538);
and U5855 (N_5855,N_4817,N_4553);
and U5856 (N_5856,N_4560,N_4733);
nand U5857 (N_5857,N_3941,N_4651);
nand U5858 (N_5858,N_3819,N_4029);
nand U5859 (N_5859,N_3930,N_4529);
nor U5860 (N_5860,N_4967,N_4778);
nand U5861 (N_5861,N_4331,N_3841);
or U5862 (N_5862,N_4122,N_4411);
nand U5863 (N_5863,N_4983,N_4726);
nand U5864 (N_5864,N_4764,N_3970);
or U5865 (N_5865,N_3916,N_4642);
nand U5866 (N_5866,N_4043,N_4004);
xnor U5867 (N_5867,N_4814,N_3819);
xnor U5868 (N_5868,N_3793,N_4976);
nor U5869 (N_5869,N_4694,N_4880);
xor U5870 (N_5870,N_3868,N_3951);
xnor U5871 (N_5871,N_4847,N_4423);
and U5872 (N_5872,N_3805,N_4041);
xor U5873 (N_5873,N_3791,N_3939);
nor U5874 (N_5874,N_4129,N_4262);
and U5875 (N_5875,N_4302,N_4606);
or U5876 (N_5876,N_4738,N_3816);
and U5877 (N_5877,N_4481,N_3990);
and U5878 (N_5878,N_4210,N_4455);
and U5879 (N_5879,N_4839,N_4785);
xor U5880 (N_5880,N_4990,N_3806);
nand U5881 (N_5881,N_4061,N_4190);
xnor U5882 (N_5882,N_3827,N_4326);
or U5883 (N_5883,N_4759,N_4117);
xor U5884 (N_5884,N_4060,N_3814);
nor U5885 (N_5885,N_3750,N_4882);
xnor U5886 (N_5886,N_4041,N_4219);
xnor U5887 (N_5887,N_4537,N_4959);
or U5888 (N_5888,N_4938,N_4466);
nor U5889 (N_5889,N_4552,N_4716);
xor U5890 (N_5890,N_4076,N_4111);
xnor U5891 (N_5891,N_4274,N_3935);
xor U5892 (N_5892,N_4949,N_4816);
xor U5893 (N_5893,N_4039,N_4448);
xnor U5894 (N_5894,N_4226,N_4673);
and U5895 (N_5895,N_4078,N_3834);
xor U5896 (N_5896,N_4193,N_4020);
nor U5897 (N_5897,N_4065,N_4021);
xor U5898 (N_5898,N_3789,N_3953);
or U5899 (N_5899,N_4627,N_3978);
or U5900 (N_5900,N_4857,N_4855);
nand U5901 (N_5901,N_4072,N_4135);
nand U5902 (N_5902,N_4166,N_4267);
xor U5903 (N_5903,N_4181,N_4591);
nand U5904 (N_5904,N_4144,N_3855);
and U5905 (N_5905,N_4705,N_4627);
xor U5906 (N_5906,N_3822,N_4882);
and U5907 (N_5907,N_4226,N_4234);
xor U5908 (N_5908,N_4072,N_4556);
and U5909 (N_5909,N_4383,N_4828);
nor U5910 (N_5910,N_3772,N_4991);
nand U5911 (N_5911,N_3887,N_4686);
nor U5912 (N_5912,N_3979,N_4127);
and U5913 (N_5913,N_4378,N_3817);
nand U5914 (N_5914,N_4326,N_4379);
nand U5915 (N_5915,N_4195,N_4212);
xor U5916 (N_5916,N_4674,N_4210);
and U5917 (N_5917,N_4105,N_4338);
nand U5918 (N_5918,N_4205,N_4139);
nand U5919 (N_5919,N_4886,N_4063);
nor U5920 (N_5920,N_4743,N_4906);
and U5921 (N_5921,N_4116,N_3889);
nand U5922 (N_5922,N_4976,N_4078);
or U5923 (N_5923,N_4288,N_4646);
nand U5924 (N_5924,N_4726,N_4222);
xor U5925 (N_5925,N_4078,N_4076);
or U5926 (N_5926,N_4740,N_4140);
or U5927 (N_5927,N_4400,N_4237);
nor U5928 (N_5928,N_3912,N_3962);
and U5929 (N_5929,N_4292,N_4577);
nor U5930 (N_5930,N_4395,N_3844);
or U5931 (N_5931,N_4615,N_4908);
xnor U5932 (N_5932,N_4331,N_3800);
or U5933 (N_5933,N_4092,N_4776);
and U5934 (N_5934,N_3904,N_4944);
nand U5935 (N_5935,N_4317,N_4669);
and U5936 (N_5936,N_3811,N_4398);
and U5937 (N_5937,N_4471,N_4208);
nand U5938 (N_5938,N_4860,N_4145);
or U5939 (N_5939,N_3893,N_3795);
and U5940 (N_5940,N_4839,N_4954);
nand U5941 (N_5941,N_4017,N_4569);
and U5942 (N_5942,N_4472,N_4250);
or U5943 (N_5943,N_4141,N_4365);
nor U5944 (N_5944,N_4292,N_4473);
xnor U5945 (N_5945,N_4450,N_4089);
nand U5946 (N_5946,N_4879,N_4765);
nor U5947 (N_5947,N_3839,N_3868);
and U5948 (N_5948,N_4488,N_3869);
or U5949 (N_5949,N_4650,N_4359);
nor U5950 (N_5950,N_4355,N_4165);
and U5951 (N_5951,N_4696,N_4429);
xnor U5952 (N_5952,N_4528,N_4026);
nand U5953 (N_5953,N_4825,N_3894);
nor U5954 (N_5954,N_4392,N_4809);
nor U5955 (N_5955,N_4950,N_4252);
or U5956 (N_5956,N_3854,N_3816);
nand U5957 (N_5957,N_4777,N_4744);
xor U5958 (N_5958,N_4686,N_3972);
or U5959 (N_5959,N_4460,N_4027);
nor U5960 (N_5960,N_4487,N_4499);
xnor U5961 (N_5961,N_3882,N_3915);
and U5962 (N_5962,N_4997,N_4912);
nand U5963 (N_5963,N_4208,N_4521);
nor U5964 (N_5964,N_4687,N_4744);
and U5965 (N_5965,N_4596,N_4024);
and U5966 (N_5966,N_4546,N_4325);
xnor U5967 (N_5967,N_4921,N_4499);
xor U5968 (N_5968,N_3903,N_3965);
or U5969 (N_5969,N_4122,N_4258);
xor U5970 (N_5970,N_4808,N_4456);
nand U5971 (N_5971,N_4902,N_4233);
nand U5972 (N_5972,N_3959,N_4770);
or U5973 (N_5973,N_3956,N_3835);
and U5974 (N_5974,N_3974,N_4296);
xnor U5975 (N_5975,N_3903,N_4399);
or U5976 (N_5976,N_4488,N_3991);
and U5977 (N_5977,N_4318,N_3870);
nand U5978 (N_5978,N_4729,N_4503);
xor U5979 (N_5979,N_4051,N_4617);
and U5980 (N_5980,N_4733,N_4307);
nor U5981 (N_5981,N_4304,N_3939);
or U5982 (N_5982,N_3820,N_4085);
xor U5983 (N_5983,N_3848,N_3923);
or U5984 (N_5984,N_4094,N_3902);
or U5985 (N_5985,N_3935,N_4317);
or U5986 (N_5986,N_3786,N_4018);
and U5987 (N_5987,N_4392,N_4572);
nor U5988 (N_5988,N_3894,N_4852);
or U5989 (N_5989,N_4137,N_3795);
xor U5990 (N_5990,N_4955,N_4244);
nand U5991 (N_5991,N_3803,N_4201);
and U5992 (N_5992,N_4500,N_4542);
and U5993 (N_5993,N_4162,N_4935);
nand U5994 (N_5994,N_3868,N_4590);
nor U5995 (N_5995,N_4612,N_4286);
or U5996 (N_5996,N_3888,N_4284);
or U5997 (N_5997,N_4173,N_4750);
nand U5998 (N_5998,N_3836,N_4917);
and U5999 (N_5999,N_4675,N_4247);
xnor U6000 (N_6000,N_4130,N_4741);
nand U6001 (N_6001,N_3832,N_4379);
or U6002 (N_6002,N_4901,N_3845);
and U6003 (N_6003,N_4820,N_4435);
xor U6004 (N_6004,N_4154,N_4121);
and U6005 (N_6005,N_4808,N_4103);
nor U6006 (N_6006,N_4584,N_4921);
and U6007 (N_6007,N_4049,N_4080);
nor U6008 (N_6008,N_4878,N_4555);
nor U6009 (N_6009,N_4069,N_4444);
nor U6010 (N_6010,N_4447,N_4158);
xor U6011 (N_6011,N_4961,N_4277);
and U6012 (N_6012,N_4444,N_3898);
nor U6013 (N_6013,N_4568,N_4382);
xnor U6014 (N_6014,N_4963,N_4415);
nand U6015 (N_6015,N_4631,N_4714);
nor U6016 (N_6016,N_4343,N_3798);
or U6017 (N_6017,N_4927,N_4939);
and U6018 (N_6018,N_4897,N_3776);
xnor U6019 (N_6019,N_4631,N_4447);
nor U6020 (N_6020,N_4201,N_4634);
nand U6021 (N_6021,N_4592,N_4310);
and U6022 (N_6022,N_4307,N_3795);
or U6023 (N_6023,N_4696,N_4130);
and U6024 (N_6024,N_4150,N_4029);
and U6025 (N_6025,N_4831,N_4291);
or U6026 (N_6026,N_4869,N_4766);
and U6027 (N_6027,N_4192,N_3778);
nand U6028 (N_6028,N_4544,N_3848);
nor U6029 (N_6029,N_4190,N_4126);
nand U6030 (N_6030,N_4761,N_3893);
nand U6031 (N_6031,N_4864,N_3969);
and U6032 (N_6032,N_4960,N_3961);
and U6033 (N_6033,N_3884,N_4586);
and U6034 (N_6034,N_4544,N_3788);
or U6035 (N_6035,N_3838,N_3934);
and U6036 (N_6036,N_4676,N_4777);
xor U6037 (N_6037,N_4171,N_3755);
or U6038 (N_6038,N_4745,N_4319);
nand U6039 (N_6039,N_3829,N_4770);
xnor U6040 (N_6040,N_4393,N_4347);
nor U6041 (N_6041,N_3808,N_4669);
and U6042 (N_6042,N_4069,N_4936);
nor U6043 (N_6043,N_4782,N_4080);
nand U6044 (N_6044,N_4562,N_4892);
nand U6045 (N_6045,N_4563,N_4479);
or U6046 (N_6046,N_4299,N_4698);
and U6047 (N_6047,N_4928,N_4641);
or U6048 (N_6048,N_4225,N_4119);
nand U6049 (N_6049,N_4451,N_4147);
or U6050 (N_6050,N_4017,N_4428);
nand U6051 (N_6051,N_4848,N_4298);
xnor U6052 (N_6052,N_3923,N_3966);
nand U6053 (N_6053,N_4536,N_4473);
or U6054 (N_6054,N_3948,N_4345);
and U6055 (N_6055,N_3957,N_3906);
nand U6056 (N_6056,N_4422,N_4885);
xnor U6057 (N_6057,N_4530,N_4783);
nor U6058 (N_6058,N_4149,N_3778);
nand U6059 (N_6059,N_4444,N_4639);
and U6060 (N_6060,N_4519,N_4635);
and U6061 (N_6061,N_4613,N_4397);
and U6062 (N_6062,N_4758,N_3761);
nand U6063 (N_6063,N_4972,N_4002);
or U6064 (N_6064,N_4585,N_4184);
nand U6065 (N_6065,N_3753,N_3907);
xnor U6066 (N_6066,N_3780,N_4784);
xnor U6067 (N_6067,N_4415,N_4340);
or U6068 (N_6068,N_3919,N_3957);
nor U6069 (N_6069,N_4379,N_4101);
xor U6070 (N_6070,N_4045,N_4552);
or U6071 (N_6071,N_4862,N_3818);
nand U6072 (N_6072,N_4423,N_3983);
and U6073 (N_6073,N_4691,N_4317);
xnor U6074 (N_6074,N_3963,N_4619);
xor U6075 (N_6075,N_4385,N_4945);
and U6076 (N_6076,N_4403,N_4129);
nand U6077 (N_6077,N_4730,N_4833);
xnor U6078 (N_6078,N_3828,N_3941);
xnor U6079 (N_6079,N_3938,N_4194);
nand U6080 (N_6080,N_4245,N_4753);
nand U6081 (N_6081,N_4922,N_4598);
or U6082 (N_6082,N_4038,N_4732);
and U6083 (N_6083,N_4605,N_4722);
or U6084 (N_6084,N_4292,N_4772);
xnor U6085 (N_6085,N_4780,N_3912);
nand U6086 (N_6086,N_4256,N_4298);
nor U6087 (N_6087,N_4479,N_4537);
and U6088 (N_6088,N_4342,N_3848);
and U6089 (N_6089,N_4566,N_4411);
nor U6090 (N_6090,N_3909,N_4719);
or U6091 (N_6091,N_3941,N_4622);
and U6092 (N_6092,N_4837,N_4909);
xnor U6093 (N_6093,N_3925,N_4922);
and U6094 (N_6094,N_4418,N_4237);
and U6095 (N_6095,N_4134,N_4609);
xor U6096 (N_6096,N_4465,N_4773);
and U6097 (N_6097,N_3788,N_4106);
and U6098 (N_6098,N_4269,N_4005);
and U6099 (N_6099,N_4181,N_3973);
xnor U6100 (N_6100,N_4590,N_4089);
and U6101 (N_6101,N_3905,N_4132);
and U6102 (N_6102,N_4480,N_4595);
xnor U6103 (N_6103,N_4705,N_4369);
xor U6104 (N_6104,N_4269,N_4421);
nand U6105 (N_6105,N_3763,N_4866);
nor U6106 (N_6106,N_3916,N_4251);
nor U6107 (N_6107,N_3782,N_4056);
xor U6108 (N_6108,N_4176,N_4318);
nand U6109 (N_6109,N_4505,N_3905);
or U6110 (N_6110,N_4257,N_4190);
nor U6111 (N_6111,N_4019,N_4072);
and U6112 (N_6112,N_4719,N_4387);
xnor U6113 (N_6113,N_4979,N_4664);
nand U6114 (N_6114,N_4759,N_4104);
nor U6115 (N_6115,N_4299,N_4312);
or U6116 (N_6116,N_4274,N_4056);
and U6117 (N_6117,N_4996,N_4753);
and U6118 (N_6118,N_4644,N_4328);
nand U6119 (N_6119,N_4667,N_4821);
nand U6120 (N_6120,N_4138,N_4993);
or U6121 (N_6121,N_4986,N_4344);
nor U6122 (N_6122,N_4990,N_4265);
nor U6123 (N_6123,N_3898,N_4595);
xnor U6124 (N_6124,N_4286,N_4336);
nand U6125 (N_6125,N_4096,N_4401);
nand U6126 (N_6126,N_3776,N_3907);
or U6127 (N_6127,N_3877,N_4539);
xor U6128 (N_6128,N_4893,N_4346);
and U6129 (N_6129,N_4387,N_4074);
nor U6130 (N_6130,N_4481,N_4684);
nor U6131 (N_6131,N_4203,N_4149);
nand U6132 (N_6132,N_4563,N_4370);
or U6133 (N_6133,N_4660,N_4766);
xor U6134 (N_6134,N_3812,N_4228);
and U6135 (N_6135,N_4760,N_4482);
nor U6136 (N_6136,N_4850,N_4430);
nor U6137 (N_6137,N_4401,N_4792);
xor U6138 (N_6138,N_4212,N_4306);
xnor U6139 (N_6139,N_4801,N_4333);
or U6140 (N_6140,N_4094,N_4421);
or U6141 (N_6141,N_3820,N_3752);
or U6142 (N_6142,N_4894,N_4649);
nand U6143 (N_6143,N_4723,N_4170);
nor U6144 (N_6144,N_4103,N_4444);
nand U6145 (N_6145,N_4083,N_4357);
nand U6146 (N_6146,N_3959,N_4928);
xor U6147 (N_6147,N_4302,N_4463);
xnor U6148 (N_6148,N_4038,N_4975);
xnor U6149 (N_6149,N_4110,N_4735);
and U6150 (N_6150,N_4882,N_3896);
or U6151 (N_6151,N_4326,N_4874);
and U6152 (N_6152,N_4987,N_4162);
nor U6153 (N_6153,N_4199,N_4116);
xnor U6154 (N_6154,N_4053,N_4847);
xnor U6155 (N_6155,N_4482,N_4936);
and U6156 (N_6156,N_4395,N_4051);
nand U6157 (N_6157,N_4859,N_4776);
nor U6158 (N_6158,N_4864,N_4936);
or U6159 (N_6159,N_3873,N_4750);
or U6160 (N_6160,N_4912,N_4858);
nand U6161 (N_6161,N_4552,N_4984);
or U6162 (N_6162,N_3875,N_4903);
nor U6163 (N_6163,N_3801,N_4120);
xor U6164 (N_6164,N_4111,N_3752);
xnor U6165 (N_6165,N_4038,N_4012);
nor U6166 (N_6166,N_4989,N_4000);
and U6167 (N_6167,N_3976,N_4948);
or U6168 (N_6168,N_4664,N_4578);
and U6169 (N_6169,N_3940,N_4185);
or U6170 (N_6170,N_4367,N_4394);
nand U6171 (N_6171,N_4635,N_4018);
nand U6172 (N_6172,N_4005,N_4308);
and U6173 (N_6173,N_4090,N_4626);
nand U6174 (N_6174,N_4638,N_4637);
nor U6175 (N_6175,N_3979,N_4210);
xnor U6176 (N_6176,N_4833,N_4108);
nor U6177 (N_6177,N_4785,N_3930);
nor U6178 (N_6178,N_4595,N_3962);
xor U6179 (N_6179,N_4604,N_4712);
nor U6180 (N_6180,N_4686,N_4497);
nand U6181 (N_6181,N_4925,N_3952);
or U6182 (N_6182,N_3956,N_3926);
and U6183 (N_6183,N_4575,N_4012);
and U6184 (N_6184,N_4157,N_4821);
and U6185 (N_6185,N_4899,N_4536);
or U6186 (N_6186,N_4225,N_4822);
nor U6187 (N_6187,N_4043,N_4104);
nand U6188 (N_6188,N_3862,N_4198);
xnor U6189 (N_6189,N_4664,N_4496);
and U6190 (N_6190,N_3836,N_3917);
or U6191 (N_6191,N_4940,N_4366);
and U6192 (N_6192,N_4419,N_3923);
nor U6193 (N_6193,N_4021,N_4959);
nand U6194 (N_6194,N_4524,N_4032);
nand U6195 (N_6195,N_4851,N_4517);
or U6196 (N_6196,N_3751,N_4536);
nor U6197 (N_6197,N_4142,N_4782);
xnor U6198 (N_6198,N_4841,N_4458);
nor U6199 (N_6199,N_4697,N_4841);
nor U6200 (N_6200,N_3814,N_4756);
or U6201 (N_6201,N_3991,N_4247);
nand U6202 (N_6202,N_3853,N_3848);
nand U6203 (N_6203,N_4486,N_4387);
or U6204 (N_6204,N_4104,N_4042);
or U6205 (N_6205,N_4256,N_4344);
nor U6206 (N_6206,N_4381,N_4396);
xnor U6207 (N_6207,N_4184,N_4089);
xor U6208 (N_6208,N_4668,N_4344);
and U6209 (N_6209,N_4198,N_3917);
and U6210 (N_6210,N_4477,N_4674);
nand U6211 (N_6211,N_4640,N_4332);
and U6212 (N_6212,N_4615,N_4071);
xnor U6213 (N_6213,N_3921,N_4824);
or U6214 (N_6214,N_4894,N_4537);
xor U6215 (N_6215,N_4349,N_4422);
nand U6216 (N_6216,N_3908,N_4779);
or U6217 (N_6217,N_3961,N_4443);
nand U6218 (N_6218,N_4102,N_3997);
and U6219 (N_6219,N_3869,N_4173);
xnor U6220 (N_6220,N_4940,N_4893);
nand U6221 (N_6221,N_4826,N_4239);
nor U6222 (N_6222,N_3846,N_4694);
nand U6223 (N_6223,N_4223,N_4837);
and U6224 (N_6224,N_4634,N_4849);
nor U6225 (N_6225,N_3978,N_4532);
xnor U6226 (N_6226,N_4793,N_4728);
nor U6227 (N_6227,N_3963,N_4724);
nand U6228 (N_6228,N_4884,N_4250);
xor U6229 (N_6229,N_4422,N_3919);
nand U6230 (N_6230,N_4260,N_3858);
xnor U6231 (N_6231,N_4929,N_4139);
nor U6232 (N_6232,N_4837,N_4763);
or U6233 (N_6233,N_4323,N_4443);
nand U6234 (N_6234,N_4148,N_4530);
nor U6235 (N_6235,N_4697,N_4583);
and U6236 (N_6236,N_4581,N_3835);
nor U6237 (N_6237,N_4020,N_4583);
or U6238 (N_6238,N_4988,N_4345);
nand U6239 (N_6239,N_4215,N_4724);
and U6240 (N_6240,N_3775,N_4312);
xnor U6241 (N_6241,N_4042,N_4651);
xor U6242 (N_6242,N_3887,N_4517);
nor U6243 (N_6243,N_4878,N_4506);
xor U6244 (N_6244,N_4387,N_3755);
and U6245 (N_6245,N_4848,N_4069);
xnor U6246 (N_6246,N_4953,N_4298);
or U6247 (N_6247,N_4883,N_3822);
nor U6248 (N_6248,N_4940,N_4476);
xnor U6249 (N_6249,N_4796,N_3903);
and U6250 (N_6250,N_5774,N_5014);
xor U6251 (N_6251,N_5161,N_5435);
nand U6252 (N_6252,N_5610,N_5583);
or U6253 (N_6253,N_5265,N_5682);
and U6254 (N_6254,N_5166,N_5157);
xnor U6255 (N_6255,N_5366,N_5137);
nand U6256 (N_6256,N_5750,N_6033);
or U6257 (N_6257,N_5864,N_5874);
nor U6258 (N_6258,N_5333,N_5293);
nand U6259 (N_6259,N_6089,N_5647);
xnor U6260 (N_6260,N_5499,N_5162);
xor U6261 (N_6261,N_5724,N_5302);
and U6262 (N_6262,N_5716,N_5117);
nand U6263 (N_6263,N_5245,N_5894);
or U6264 (N_6264,N_5773,N_5702);
nand U6265 (N_6265,N_5381,N_5490);
or U6266 (N_6266,N_5730,N_6172);
xnor U6267 (N_6267,N_5028,N_5115);
nand U6268 (N_6268,N_5072,N_5844);
and U6269 (N_6269,N_5050,N_6083);
xnor U6270 (N_6270,N_5421,N_5980);
nor U6271 (N_6271,N_6065,N_5908);
nor U6272 (N_6272,N_6047,N_6192);
nand U6273 (N_6273,N_5862,N_5810);
nand U6274 (N_6274,N_5815,N_6231);
or U6275 (N_6275,N_5272,N_5714);
nor U6276 (N_6276,N_5651,N_6141);
nand U6277 (N_6277,N_6096,N_5200);
xor U6278 (N_6278,N_5653,N_5939);
xnor U6279 (N_6279,N_5589,N_5005);
and U6280 (N_6280,N_5854,N_6003);
xor U6281 (N_6281,N_5936,N_5349);
xor U6282 (N_6282,N_5229,N_5711);
xnor U6283 (N_6283,N_5378,N_5213);
nor U6284 (N_6284,N_5769,N_5994);
or U6285 (N_6285,N_5822,N_5422);
and U6286 (N_6286,N_5607,N_5158);
and U6287 (N_6287,N_5738,N_5767);
and U6288 (N_6288,N_5344,N_5972);
and U6289 (N_6289,N_5118,N_5690);
nor U6290 (N_6290,N_5664,N_5827);
nand U6291 (N_6291,N_6148,N_6064);
nand U6292 (N_6292,N_5561,N_6098);
nand U6293 (N_6293,N_5903,N_5974);
nor U6294 (N_6294,N_5726,N_5276);
nor U6295 (N_6295,N_5102,N_5342);
nand U6296 (N_6296,N_5065,N_5728);
xor U6297 (N_6297,N_6113,N_5725);
nand U6298 (N_6298,N_6163,N_5802);
xnor U6299 (N_6299,N_6228,N_6165);
nand U6300 (N_6300,N_5996,N_5643);
or U6301 (N_6301,N_5965,N_5734);
nand U6302 (N_6302,N_5476,N_5929);
xnor U6303 (N_6303,N_6120,N_5485);
and U6304 (N_6304,N_5839,N_5443);
nand U6305 (N_6305,N_5469,N_5517);
or U6306 (N_6306,N_5202,N_5587);
or U6307 (N_6307,N_5759,N_5480);
nor U6308 (N_6308,N_5203,N_5018);
xnor U6309 (N_6309,N_6205,N_5294);
nand U6310 (N_6310,N_5247,N_6219);
nor U6311 (N_6311,N_5787,N_5695);
nand U6312 (N_6312,N_5244,N_5508);
xnor U6313 (N_6313,N_6152,N_5308);
nand U6314 (N_6314,N_6224,N_5393);
and U6315 (N_6315,N_5627,N_5883);
xor U6316 (N_6316,N_5592,N_5012);
or U6317 (N_6317,N_5145,N_5900);
nor U6318 (N_6318,N_5870,N_5323);
nand U6319 (N_6319,N_5257,N_5122);
and U6320 (N_6320,N_5928,N_5792);
xor U6321 (N_6321,N_5681,N_5328);
and U6322 (N_6322,N_5588,N_5925);
xnor U6323 (N_6323,N_5842,N_5009);
and U6324 (N_6324,N_6051,N_5614);
xor U6325 (N_6325,N_5116,N_5068);
nand U6326 (N_6326,N_6230,N_6106);
nor U6327 (N_6327,N_5321,N_5875);
or U6328 (N_6328,N_5631,N_5367);
and U6329 (N_6329,N_5295,N_6057);
xor U6330 (N_6330,N_5857,N_5804);
and U6331 (N_6331,N_5484,N_5825);
xnor U6332 (N_6332,N_5374,N_5222);
xor U6333 (N_6333,N_5687,N_5548);
nor U6334 (N_6334,N_5677,N_5935);
and U6335 (N_6335,N_5261,N_5639);
xor U6336 (N_6336,N_5940,N_5088);
nand U6337 (N_6337,N_5676,N_5955);
xor U6338 (N_6338,N_5616,N_5943);
or U6339 (N_6339,N_6093,N_5135);
or U6340 (N_6340,N_5348,N_5579);
xnor U6341 (N_6341,N_5309,N_5895);
xnor U6342 (N_6342,N_5569,N_5466);
nor U6343 (N_6343,N_6121,N_6158);
nor U6344 (N_6344,N_5345,N_5199);
or U6345 (N_6345,N_5004,N_5432);
nand U6346 (N_6346,N_5729,N_5733);
and U6347 (N_6347,N_5034,N_5696);
nand U6348 (N_6348,N_5154,N_5277);
and U6349 (N_6349,N_5745,N_6218);
xnor U6350 (N_6350,N_5584,N_5255);
nand U6351 (N_6351,N_6056,N_6118);
nand U6352 (N_6352,N_5658,N_6114);
xor U6353 (N_6353,N_5095,N_5542);
or U6354 (N_6354,N_5789,N_5577);
xnor U6355 (N_6355,N_5826,N_5160);
xor U6356 (N_6356,N_5352,N_5701);
xor U6357 (N_6357,N_6050,N_5392);
nor U6358 (N_6358,N_6168,N_5156);
or U6359 (N_6359,N_6081,N_5568);
nand U6360 (N_6360,N_5927,N_5578);
xor U6361 (N_6361,N_5477,N_6097);
or U6362 (N_6362,N_6073,N_5471);
nor U6363 (N_6363,N_6142,N_5281);
or U6364 (N_6364,N_5315,N_5192);
nor U6365 (N_6365,N_5661,N_5560);
and U6366 (N_6366,N_5020,N_5510);
nand U6367 (N_6367,N_5977,N_5678);
nand U6368 (N_6368,N_5470,N_5475);
nand U6369 (N_6369,N_6014,N_5762);
nand U6370 (N_6370,N_6227,N_5455);
xor U6371 (N_6371,N_5305,N_5566);
or U6372 (N_6372,N_5452,N_5000);
xnor U6373 (N_6373,N_5371,N_6061);
nor U6374 (N_6374,N_5872,N_5986);
or U6375 (N_6375,N_5002,N_5772);
or U6376 (N_6376,N_5386,N_5163);
and U6377 (N_6377,N_6013,N_5140);
nand U6378 (N_6378,N_5880,N_5298);
or U6379 (N_6379,N_6104,N_5620);
xnor U6380 (N_6380,N_6167,N_5128);
or U6381 (N_6381,N_5076,N_6030);
nand U6382 (N_6382,N_6229,N_5217);
or U6383 (N_6383,N_5586,N_5081);
xor U6384 (N_6384,N_5524,N_5377);
nand U6385 (N_6385,N_5752,N_6049);
nor U6386 (N_6386,N_5554,N_5411);
or U6387 (N_6387,N_6105,N_6072);
or U6388 (N_6388,N_5101,N_5087);
and U6389 (N_6389,N_5181,N_5211);
xor U6390 (N_6390,N_5189,N_6087);
or U6391 (N_6391,N_5246,N_5093);
and U6392 (N_6392,N_5365,N_6000);
xor U6393 (N_6393,N_5650,N_6235);
xnor U6394 (N_6394,N_5462,N_5106);
nor U6395 (N_6395,N_5628,N_5278);
nand U6396 (N_6396,N_5159,N_5420);
nand U6397 (N_6397,N_5855,N_6066);
or U6398 (N_6398,N_5543,N_6078);
xor U6399 (N_6399,N_5464,N_5694);
nor U6400 (N_6400,N_5040,N_5585);
nand U6401 (N_6401,N_5882,N_5399);
nor U6402 (N_6402,N_5888,N_5791);
or U6403 (N_6403,N_5805,N_5867);
nand U6404 (N_6404,N_6074,N_6201);
and U6405 (N_6405,N_5722,N_5416);
nor U6406 (N_6406,N_6191,N_5948);
or U6407 (N_6407,N_6226,N_5394);
and U6408 (N_6408,N_6108,N_5871);
and U6409 (N_6409,N_5617,N_5788);
nor U6410 (N_6410,N_5066,N_6238);
nand U6411 (N_6411,N_6067,N_5251);
and U6412 (N_6412,N_5672,N_5183);
and U6413 (N_6413,N_5613,N_5231);
nand U6414 (N_6414,N_5152,N_5454);
nor U6415 (N_6415,N_5131,N_5039);
and U6416 (N_6416,N_5515,N_5434);
or U6417 (N_6417,N_5803,N_5536);
nand U6418 (N_6418,N_5336,N_5016);
xor U6419 (N_6419,N_5307,N_5129);
nor U6420 (N_6420,N_5912,N_6237);
and U6421 (N_6421,N_5615,N_6214);
and U6422 (N_6422,N_5141,N_5313);
or U6423 (N_6423,N_6159,N_5194);
and U6424 (N_6424,N_5838,N_5148);
nor U6425 (N_6425,N_6086,N_6063);
nor U6426 (N_6426,N_6101,N_5492);
nand U6427 (N_6427,N_6135,N_5498);
xnor U6428 (N_6428,N_5937,N_6052);
nand U6429 (N_6429,N_6025,N_6156);
nand U6430 (N_6430,N_5460,N_6054);
nand U6431 (N_6431,N_5735,N_5384);
or U6432 (N_6432,N_5057,N_5124);
nand U6433 (N_6433,N_5654,N_5758);
nand U6434 (N_6434,N_5011,N_6139);
nand U6435 (N_6435,N_5896,N_5234);
and U6436 (N_6436,N_5144,N_6005);
or U6437 (N_6437,N_5784,N_6055);
and U6438 (N_6438,N_6207,N_5709);
nand U6439 (N_6439,N_5723,N_5852);
or U6440 (N_6440,N_5227,N_6138);
nand U6441 (N_6441,N_5840,N_6040);
nand U6442 (N_6442,N_5080,N_5109);
or U6443 (N_6443,N_6107,N_5567);
nand U6444 (N_6444,N_5742,N_6177);
nand U6445 (N_6445,N_5970,N_5429);
nand U6446 (N_6446,N_5132,N_5755);
nor U6447 (N_6447,N_5120,N_5624);
and U6448 (N_6448,N_5973,N_5021);
or U6449 (N_6449,N_5893,N_5680);
and U6450 (N_6450,N_5982,N_6234);
and U6451 (N_6451,N_5509,N_5916);
nor U6452 (N_6452,N_5611,N_5388);
nand U6453 (N_6453,N_5179,N_5488);
nor U6454 (N_6454,N_5898,N_5878);
and U6455 (N_6455,N_5059,N_5642);
xor U6456 (N_6456,N_5901,N_6085);
xor U6457 (N_6457,N_5847,N_5280);
and U6458 (N_6458,N_5530,N_6016);
and U6459 (N_6459,N_6164,N_5529);
nor U6460 (N_6460,N_5914,N_5559);
or U6461 (N_6461,N_5877,N_6195);
nor U6462 (N_6462,N_6112,N_6143);
or U6463 (N_6463,N_5235,N_5666);
nand U6464 (N_6464,N_5551,N_6193);
nor U6465 (N_6465,N_5727,N_6242);
nor U6466 (N_6466,N_5541,N_5030);
nor U6467 (N_6467,N_6161,N_5649);
or U6468 (N_6468,N_5155,N_5688);
nor U6469 (N_6469,N_5770,N_6088);
nand U6470 (N_6470,N_6090,N_5941);
nand U6471 (N_6471,N_5299,N_6128);
xor U6472 (N_6472,N_6092,N_6182);
nand U6473 (N_6473,N_6111,N_5022);
nor U6474 (N_6474,N_6004,N_5634);
or U6475 (N_6475,N_5552,N_6011);
nand U6476 (N_6476,N_5410,N_5191);
nor U6477 (N_6477,N_5397,N_5290);
nand U6478 (N_6478,N_5926,N_5453);
or U6479 (N_6479,N_5494,N_5591);
nor U6480 (N_6480,N_5673,N_5351);
and U6481 (N_6481,N_5123,N_5845);
or U6482 (N_6482,N_6058,N_5683);
xor U6483 (N_6483,N_5099,N_5419);
nor U6484 (N_6484,N_6185,N_5286);
nor U6485 (N_6485,N_5899,N_5346);
nor U6486 (N_6486,N_5172,N_6035);
nand U6487 (N_6487,N_5902,N_5232);
xnor U6488 (N_6488,N_5330,N_5461);
nor U6489 (N_6489,N_5049,N_5019);
and U6490 (N_6490,N_5915,N_5482);
or U6491 (N_6491,N_5786,N_6213);
or U6492 (N_6492,N_6175,N_5186);
nor U6493 (N_6493,N_6077,N_5423);
xor U6494 (N_6494,N_5090,N_5623);
and U6495 (N_6495,N_5881,N_5104);
nand U6496 (N_6496,N_6184,N_5311);
nand U6497 (N_6497,N_5026,N_5856);
xor U6498 (N_6498,N_6070,N_5473);
nor U6499 (N_6499,N_5267,N_5350);
nand U6500 (N_6500,N_6020,N_5291);
and U6501 (N_6501,N_5641,N_6069);
nand U6502 (N_6502,N_5771,N_5987);
xor U6503 (N_6503,N_5873,N_5303);
nor U6504 (N_6504,N_6146,N_5017);
and U6505 (N_6505,N_5830,N_5151);
nor U6506 (N_6506,N_6059,N_5989);
and U6507 (N_6507,N_5175,N_5932);
or U6508 (N_6508,N_5174,N_5547);
xor U6509 (N_6509,N_6117,N_6129);
nor U6510 (N_6510,N_6102,N_5775);
nor U6511 (N_6511,N_6075,N_5886);
nor U6512 (N_6512,N_5999,N_5525);
or U6513 (N_6513,N_5168,N_5817);
xnor U6514 (N_6514,N_5983,N_6041);
and U6515 (N_6515,N_5138,N_5660);
nor U6516 (N_6516,N_5210,N_5979);
or U6517 (N_6517,N_5513,N_6140);
nor U6518 (N_6518,N_6209,N_6157);
xnor U6519 (N_6519,N_5923,N_5981);
nor U6520 (N_6520,N_5663,N_5415);
nand U6521 (N_6521,N_5630,N_5086);
and U6522 (N_6522,N_5966,N_6217);
and U6523 (N_6523,N_6126,N_5753);
nand U6524 (N_6524,N_5165,N_5256);
xnor U6525 (N_6525,N_5546,N_5736);
and U6526 (N_6526,N_6053,N_5783);
or U6527 (N_6527,N_5100,N_6180);
nor U6528 (N_6528,N_5865,N_5142);
xnor U6529 (N_6529,N_5938,N_6239);
or U6530 (N_6530,N_5204,N_5749);
or U6531 (N_6531,N_5853,N_6045);
and U6532 (N_6532,N_5438,N_5190);
and U6533 (N_6533,N_5967,N_5555);
or U6534 (N_6534,N_5780,N_5287);
nor U6535 (N_6535,N_5077,N_5357);
xnor U6536 (N_6536,N_5035,N_5218);
or U6537 (N_6537,N_5337,N_5369);
nor U6538 (N_6538,N_5674,N_6008);
nor U6539 (N_6539,N_5465,N_5570);
nand U6540 (N_6540,N_5814,N_5376);
and U6541 (N_6541,N_5604,N_5075);
or U6542 (N_6542,N_5139,N_5959);
or U6543 (N_6543,N_5505,N_5644);
nor U6544 (N_6544,N_5402,N_5706);
or U6545 (N_6545,N_5924,N_5317);
or U6546 (N_6546,N_6243,N_5684);
xnor U6547 (N_6547,N_5236,N_5091);
nand U6548 (N_6548,N_5380,N_5521);
xor U6549 (N_6549,N_5952,N_5364);
and U6550 (N_6550,N_5708,N_5667);
xnor U6551 (N_6551,N_5233,N_6189);
and U6552 (N_6552,N_5990,N_5041);
xnor U6553 (N_6553,N_5212,N_6154);
nor U6554 (N_6554,N_5445,N_5562);
and U6555 (N_6555,N_5799,N_5282);
xnor U6556 (N_6556,N_5069,N_5608);
and U6557 (N_6557,N_5169,N_5637);
or U6558 (N_6558,N_5887,N_5060);
or U6559 (N_6559,N_5851,N_5909);
nand U6560 (N_6560,N_6194,N_5114);
nor U6561 (N_6561,N_5489,N_5431);
and U6562 (N_6562,N_6095,N_5503);
nand U6563 (N_6563,N_5031,N_5747);
or U6564 (N_6564,N_5539,N_5668);
or U6565 (N_6565,N_5763,N_5514);
and U6566 (N_6566,N_5963,N_6130);
or U6567 (N_6567,N_5008,N_5013);
xor U6568 (N_6568,N_5910,N_5646);
nor U6569 (N_6569,N_5809,N_5495);
xor U6570 (N_6570,N_5359,N_5876);
nor U6571 (N_6571,N_5836,N_5905);
nand U6572 (N_6572,N_5575,N_5697);
nor U6573 (N_6573,N_5250,N_5931);
xor U6574 (N_6574,N_5969,N_5713);
nand U6575 (N_6575,N_5430,N_5754);
xnor U6576 (N_6576,N_5954,N_5861);
xnor U6577 (N_6577,N_5576,N_5127);
xor U6578 (N_6578,N_5563,N_5180);
xnor U6579 (N_6579,N_5626,N_5051);
xnor U6580 (N_6580,N_5632,N_5582);
xnor U6581 (N_6581,N_5300,N_5372);
and U6582 (N_6582,N_6171,N_6208);
nor U6583 (N_6583,N_5597,N_5382);
xnor U6584 (N_6584,N_5848,N_5717);
or U6585 (N_6585,N_5340,N_5698);
nand U6586 (N_6586,N_5528,N_5596);
and U6587 (N_6587,N_5474,N_5042);
xor U6588 (N_6588,N_6080,N_6115);
nor U6589 (N_6589,N_5712,N_5648);
and U6590 (N_6590,N_5593,N_5662);
nor U6591 (N_6591,N_5441,N_5831);
and U6592 (N_6592,N_6188,N_6124);
nor U6593 (N_6593,N_6187,N_6244);
xor U6594 (N_6594,N_5292,N_5073);
xnor U6595 (N_6595,N_5507,N_5496);
xnor U6596 (N_6596,N_5125,N_6007);
and U6597 (N_6597,N_5868,N_5849);
nand U6598 (N_6598,N_5437,N_5418);
nand U6599 (N_6599,N_5944,N_5025);
nand U6600 (N_6600,N_5595,N_5686);
or U6601 (N_6601,N_5133,N_5571);
nor U6602 (N_6602,N_5297,N_5500);
and U6603 (N_6603,N_5829,N_5010);
xor U6604 (N_6604,N_6215,N_5198);
nand U6605 (N_6605,N_5052,N_6166);
nor U6606 (N_6606,N_5493,N_5519);
xor U6607 (N_6607,N_5756,N_5007);
or U6608 (N_6608,N_5718,N_5779);
nand U6609 (N_6609,N_5329,N_5835);
nand U6610 (N_6610,N_5195,N_5964);
xor U6611 (N_6611,N_5228,N_5258);
xnor U6612 (N_6612,N_5064,N_5679);
and U6613 (N_6613,N_6220,N_6169);
xnor U6614 (N_6614,N_5998,N_5121);
nor U6615 (N_6615,N_6018,N_6178);
nand U6616 (N_6616,N_5268,N_5549);
or U6617 (N_6617,N_5240,N_5621);
and U6618 (N_6618,N_5837,N_5130);
and U6619 (N_6619,N_5483,N_5220);
and U6620 (N_6620,N_5691,N_5373);
nor U6621 (N_6621,N_5045,N_5890);
xor U6622 (N_6622,N_5564,N_6137);
and U6623 (N_6623,N_5044,N_5573);
or U6624 (N_6624,N_5523,N_5375);
nor U6625 (N_6625,N_5995,N_5670);
or U6626 (N_6626,N_5097,N_5618);
and U6627 (N_6627,N_5834,N_6186);
nor U6628 (N_6628,N_5544,N_5176);
nor U6629 (N_6629,N_6046,N_5859);
nor U6630 (N_6630,N_5098,N_5215);
and U6631 (N_6631,N_5993,N_5408);
nor U6632 (N_6632,N_5574,N_5846);
and U6633 (N_6633,N_5304,N_5143);
nand U6634 (N_6634,N_5417,N_5720);
nor U6635 (N_6635,N_5396,N_5946);
or U6636 (N_6636,N_5598,N_5807);
or U6637 (N_6637,N_5395,N_5055);
or U6638 (N_6638,N_5556,N_5656);
and U6639 (N_6639,N_5391,N_5710);
and U6640 (N_6640,N_6149,N_6136);
xor U6641 (N_6641,N_5322,N_6198);
xnor U6642 (N_6642,N_5401,N_5732);
or U6643 (N_6643,N_5289,N_5897);
xnor U6644 (N_6644,N_5645,N_5652);
and U6645 (N_6645,N_5638,N_5640);
xor U6646 (N_6646,N_6245,N_6038);
or U6647 (N_6647,N_5033,N_5223);
xor U6648 (N_6648,N_5793,N_5197);
xor U6649 (N_6649,N_5491,N_6196);
nand U6650 (N_6650,N_6131,N_5283);
and U6651 (N_6651,N_5226,N_5334);
nor U6652 (N_6652,N_6071,N_5037);
nand U6653 (N_6653,N_5119,N_5406);
or U6654 (N_6654,N_5083,N_6134);
or U6655 (N_6655,N_5209,N_5933);
nor U6656 (N_6656,N_5361,N_5450);
xnor U6657 (N_6657,N_5458,N_5860);
or U6658 (N_6658,N_5146,N_5599);
xor U6659 (N_6659,N_5306,N_5126);
nand U6660 (N_6660,N_5383,N_6155);
nor U6661 (N_6661,N_5777,N_6091);
nand U6662 (N_6662,N_5600,N_6019);
and U6663 (N_6663,N_5748,N_5545);
and U6664 (N_6664,N_5043,N_6028);
nor U6665 (N_6665,N_6153,N_5619);
or U6666 (N_6666,N_6110,N_5355);
nand U6667 (N_6667,N_6012,N_5572);
or U6668 (N_6668,N_5414,N_5858);
nor U6669 (N_6669,N_5047,N_5107);
or U6670 (N_6670,N_5794,N_5015);
and U6671 (N_6671,N_5920,N_5238);
and U6672 (N_6672,N_5061,N_6002);
or U6673 (N_6673,N_6026,N_6246);
and U6674 (N_6674,N_5533,N_5719);
xnor U6675 (N_6675,N_5207,N_5451);
nand U6676 (N_6676,N_5188,N_5746);
nand U6677 (N_6677,N_6109,N_6162);
and U6678 (N_6678,N_5796,N_6127);
xnor U6679 (N_6679,N_5693,N_6133);
nand U6680 (N_6680,N_5085,N_5806);
xor U6681 (N_6681,N_5006,N_5526);
or U6682 (N_6682,N_6029,N_5721);
xor U6683 (N_6683,N_5692,N_5550);
nor U6684 (N_6684,N_5820,N_5655);
and U6685 (N_6685,N_5707,N_5379);
nor U6686 (N_6686,N_5024,N_5553);
nand U6687 (N_6687,N_6151,N_5961);
xor U6688 (N_6688,N_5284,N_5766);
xor U6689 (N_6689,N_5518,N_5606);
and U6690 (N_6690,N_5316,N_5906);
xor U6691 (N_6691,N_5478,N_6001);
xnor U6692 (N_6692,N_5703,N_6204);
and U6693 (N_6693,N_5092,N_5270);
or U6694 (N_6694,N_5992,N_5400);
and U6695 (N_6695,N_5689,N_5456);
or U6696 (N_6696,N_6084,N_5739);
and U6697 (N_6697,N_6147,N_5744);
xor U6698 (N_6698,N_5918,N_5003);
or U6699 (N_6699,N_5581,N_5447);
or U6700 (N_6700,N_5063,N_5070);
xnor U6701 (N_6701,N_5960,N_5765);
nand U6702 (N_6702,N_5962,N_6099);
nand U6703 (N_6703,N_5459,N_5193);
and U6704 (N_6704,N_5531,N_5808);
or U6705 (N_6705,N_5412,N_5889);
and U6706 (N_6706,N_6039,N_5913);
xor U6707 (N_6707,N_5413,N_5958);
nand U6708 (N_6708,N_5254,N_5259);
and U6709 (N_6709,N_5971,N_5850);
and U6710 (N_6710,N_5237,N_6024);
and U6711 (N_6711,N_6181,N_5343);
and U6712 (N_6712,N_6247,N_5260);
or U6713 (N_6713,N_5326,N_5285);
xnor U6714 (N_6714,N_5335,N_5404);
or U6715 (N_6715,N_5502,N_6068);
nor U6716 (N_6716,N_5824,N_5046);
nand U6717 (N_6717,N_6015,N_5327);
and U6718 (N_6718,N_5084,N_6043);
or U6719 (N_6719,N_5731,N_5038);
or U6720 (N_6720,N_5332,N_5934);
xor U6721 (N_6721,N_6037,N_6027);
or U6722 (N_6722,N_5310,N_6241);
or U6723 (N_6723,N_5105,N_6223);
xnor U6724 (N_6724,N_5398,N_5813);
and U6725 (N_6725,N_5978,N_5387);
xnor U6726 (N_6726,N_5150,N_5094);
nor U6727 (N_6727,N_5705,N_5699);
nor U6728 (N_6728,N_5479,N_5472);
nor U6729 (N_6729,N_5764,N_5884);
nand U6730 (N_6730,N_5975,N_5532);
nand U6731 (N_6731,N_5950,N_5512);
nor U6732 (N_6732,N_5319,N_5869);
or U6733 (N_6733,N_5785,N_5605);
xnor U6734 (N_6734,N_5216,N_6119);
and U6735 (N_6735,N_5953,N_5230);
nor U6736 (N_6736,N_5288,N_5023);
nor U6737 (N_6737,N_5205,N_5390);
xnor U6738 (N_6738,N_5685,N_5439);
nor U6739 (N_6739,N_5601,N_5782);
nand U6740 (N_6740,N_5801,N_5405);
xnor U6741 (N_6741,N_5173,N_6210);
or U6742 (N_6742,N_5968,N_5629);
and U6743 (N_6743,N_5446,N_6232);
nor U6744 (N_6744,N_5241,N_5919);
nor U6745 (N_6745,N_5985,N_5248);
nand U6746 (N_6746,N_5448,N_5930);
or U6747 (N_6747,N_5922,N_5761);
and U6748 (N_6748,N_6225,N_5239);
or U6749 (N_6749,N_5704,N_5273);
xor U6750 (N_6750,N_5740,N_6199);
xor U6751 (N_6751,N_5428,N_5800);
or U6752 (N_6752,N_5540,N_5436);
xor U6753 (N_6753,N_5486,N_5219);
nor U6754 (N_6754,N_5296,N_5949);
nand U6755 (N_6755,N_5997,N_6125);
or U6756 (N_6756,N_5904,N_5062);
or U6757 (N_6757,N_5768,N_5885);
xnor U6758 (N_6758,N_6183,N_5942);
and U6759 (N_6759,N_5565,N_5403);
and U6760 (N_6760,N_5389,N_5185);
nor U6761 (N_6761,N_6031,N_5225);
nand U6762 (N_6762,N_5468,N_5467);
nor U6763 (N_6763,N_6170,N_5338);
nor U6764 (N_6764,N_5504,N_5027);
nand U6765 (N_6765,N_5622,N_5187);
or U6766 (N_6766,N_5036,N_5609);
or U6767 (N_6767,N_5032,N_5635);
and U6768 (N_6768,N_5368,N_5602);
nand U6769 (N_6769,N_5590,N_6202);
nand U6770 (N_6770,N_6173,N_6079);
and U6771 (N_6771,N_5951,N_5659);
or U6772 (N_6772,N_5358,N_6021);
or U6773 (N_6773,N_6212,N_5096);
nand U6774 (N_6774,N_5798,N_5527);
xnor U6775 (N_6775,N_5449,N_5339);
nand U6776 (N_6776,N_5177,N_5108);
nor U6777 (N_6777,N_5790,N_6094);
xor U6778 (N_6778,N_5892,N_5275);
and U6779 (N_6779,N_5497,N_5751);
nand U6780 (N_6780,N_5113,N_5487);
or U6781 (N_6781,N_5669,N_5249);
and U6782 (N_6782,N_5612,N_5074);
nor U6783 (N_6783,N_5048,N_5818);
xnor U6784 (N_6784,N_5426,N_6179);
xnor U6785 (N_6785,N_5221,N_5506);
and U6786 (N_6786,N_5269,N_5812);
and U6787 (N_6787,N_5153,N_5353);
and U6788 (N_6788,N_5440,N_5843);
nor U6789 (N_6789,N_5424,N_5262);
or U6790 (N_6790,N_5301,N_5457);
nor U6791 (N_6791,N_5314,N_5743);
nor U6792 (N_6792,N_5347,N_5700);
nand U6793 (N_6793,N_5945,N_5665);
or U6794 (N_6794,N_5866,N_5201);
and U6795 (N_6795,N_5331,N_5224);
nor U6796 (N_6796,N_6150,N_6044);
and U6797 (N_6797,N_6076,N_5167);
nand U6798 (N_6798,N_5657,N_5511);
and U6799 (N_6799,N_5832,N_5208);
xor U6800 (N_6800,N_5111,N_5427);
xor U6801 (N_6801,N_6082,N_5538);
nor U6802 (N_6802,N_6022,N_5911);
or U6803 (N_6803,N_6062,N_5433);
xnor U6804 (N_6804,N_5947,N_5671);
xor U6805 (N_6805,N_5891,N_6197);
or U6806 (N_6806,N_5580,N_5921);
xnor U6807 (N_6807,N_6132,N_6203);
nor U6808 (N_6808,N_6221,N_6211);
or U6809 (N_6809,N_5325,N_5136);
nand U6810 (N_6810,N_5558,N_5534);
nor U6811 (N_6811,N_6144,N_5795);
and U6812 (N_6812,N_5320,N_5833);
nor U6813 (N_6813,N_6048,N_5907);
nor U6814 (N_6814,N_5078,N_6042);
xnor U6815 (N_6815,N_5385,N_5957);
nand U6816 (N_6816,N_5196,N_5603);
and U6817 (N_6817,N_5737,N_5149);
nand U6818 (N_6818,N_5147,N_5263);
nand U6819 (N_6819,N_6116,N_5134);
and U6820 (N_6820,N_6206,N_6176);
nand U6821 (N_6821,N_6006,N_5797);
nor U6822 (N_6822,N_6174,N_5991);
or U6823 (N_6823,N_5407,N_5242);
xnor U6824 (N_6824,N_5819,N_6103);
nor U6825 (N_6825,N_5520,N_6123);
or U6826 (N_6826,N_6100,N_5082);
nor U6827 (N_6827,N_5984,N_5089);
nand U6828 (N_6828,N_5001,N_5409);
and U6829 (N_6829,N_5988,N_5781);
or U6830 (N_6830,N_6249,N_5370);
xnor U6831 (N_6831,N_5253,N_5760);
nor U6832 (N_6832,N_5164,N_5633);
and U6833 (N_6833,N_5252,N_5776);
xor U6834 (N_6834,N_6222,N_5442);
nand U6835 (N_6835,N_5079,N_5279);
nor U6836 (N_6836,N_6060,N_5171);
and U6837 (N_6837,N_5594,N_5841);
nand U6838 (N_6838,N_5112,N_5206);
xnor U6839 (N_6839,N_5053,N_5741);
xnor U6840 (N_6840,N_6032,N_5274);
xor U6841 (N_6841,N_6145,N_6010);
or U6842 (N_6842,N_6248,N_5318);
and U6843 (N_6843,N_6233,N_5463);
and U6844 (N_6844,N_5715,N_5360);
nand U6845 (N_6845,N_5056,N_5956);
xnor U6846 (N_6846,N_5029,N_5058);
nand U6847 (N_6847,N_5271,N_5675);
or U6848 (N_6848,N_6160,N_5481);
nor U6849 (N_6849,N_5535,N_5324);
or U6850 (N_6850,N_5184,N_5243);
xor U6851 (N_6851,N_6017,N_6036);
and U6852 (N_6852,N_5341,N_5110);
xnor U6853 (N_6853,N_5823,N_6034);
or U6854 (N_6854,N_6240,N_6190);
and U6855 (N_6855,N_5356,N_6200);
xor U6856 (N_6856,N_5363,N_5067);
xnor U6857 (N_6857,N_5170,N_5182);
nand U6858 (N_6858,N_5811,N_6236);
or U6859 (N_6859,N_5425,N_5757);
nand U6860 (N_6860,N_5214,N_5557);
nor U6861 (N_6861,N_5071,N_6216);
or U6862 (N_6862,N_5625,N_5054);
and U6863 (N_6863,N_6023,N_5312);
xor U6864 (N_6864,N_5354,N_5636);
or U6865 (N_6865,N_5178,N_5444);
nand U6866 (N_6866,N_5537,N_5103);
nand U6867 (N_6867,N_5816,N_5264);
nor U6868 (N_6868,N_5828,N_5879);
nand U6869 (N_6869,N_5516,N_5501);
nand U6870 (N_6870,N_5917,N_5976);
nand U6871 (N_6871,N_5362,N_5266);
and U6872 (N_6872,N_5778,N_5821);
nor U6873 (N_6873,N_5522,N_5863);
and U6874 (N_6874,N_6122,N_6009);
xor U6875 (N_6875,N_6097,N_5592);
or U6876 (N_6876,N_5938,N_6002);
or U6877 (N_6877,N_6188,N_5777);
nand U6878 (N_6878,N_5485,N_6157);
nand U6879 (N_6879,N_6060,N_6032);
and U6880 (N_6880,N_5732,N_5821);
or U6881 (N_6881,N_5604,N_5765);
xor U6882 (N_6882,N_5204,N_5377);
xor U6883 (N_6883,N_5584,N_5119);
or U6884 (N_6884,N_6122,N_5301);
nor U6885 (N_6885,N_5454,N_6040);
and U6886 (N_6886,N_6227,N_5184);
xor U6887 (N_6887,N_5950,N_5836);
and U6888 (N_6888,N_6231,N_6145);
or U6889 (N_6889,N_6031,N_6048);
and U6890 (N_6890,N_5682,N_5710);
nor U6891 (N_6891,N_5433,N_5103);
or U6892 (N_6892,N_5573,N_6215);
and U6893 (N_6893,N_5681,N_5035);
nor U6894 (N_6894,N_6117,N_5074);
nand U6895 (N_6895,N_5396,N_5750);
and U6896 (N_6896,N_5556,N_5680);
nand U6897 (N_6897,N_5670,N_5475);
nand U6898 (N_6898,N_5879,N_5636);
xor U6899 (N_6899,N_5349,N_5212);
or U6900 (N_6900,N_5004,N_5167);
or U6901 (N_6901,N_5989,N_5747);
or U6902 (N_6902,N_6169,N_6243);
nand U6903 (N_6903,N_5948,N_5311);
nand U6904 (N_6904,N_5703,N_5570);
xor U6905 (N_6905,N_5727,N_5792);
nor U6906 (N_6906,N_5031,N_5096);
and U6907 (N_6907,N_5125,N_5515);
and U6908 (N_6908,N_5157,N_6169);
nand U6909 (N_6909,N_5143,N_5820);
nor U6910 (N_6910,N_5274,N_5748);
nand U6911 (N_6911,N_6074,N_5314);
nand U6912 (N_6912,N_5567,N_5558);
xor U6913 (N_6913,N_6222,N_5544);
and U6914 (N_6914,N_5091,N_5753);
nand U6915 (N_6915,N_5544,N_5255);
and U6916 (N_6916,N_6011,N_6151);
xnor U6917 (N_6917,N_5085,N_5498);
or U6918 (N_6918,N_6165,N_5709);
xor U6919 (N_6919,N_6023,N_5977);
nand U6920 (N_6920,N_5038,N_6190);
or U6921 (N_6921,N_5426,N_5967);
or U6922 (N_6922,N_5987,N_5576);
nand U6923 (N_6923,N_6001,N_5928);
nand U6924 (N_6924,N_5025,N_5332);
and U6925 (N_6925,N_5665,N_5203);
xnor U6926 (N_6926,N_5119,N_5508);
xnor U6927 (N_6927,N_6081,N_6008);
and U6928 (N_6928,N_5387,N_6155);
nand U6929 (N_6929,N_5717,N_5611);
or U6930 (N_6930,N_5938,N_5167);
and U6931 (N_6931,N_5548,N_5726);
xnor U6932 (N_6932,N_5127,N_5561);
or U6933 (N_6933,N_5069,N_5649);
and U6934 (N_6934,N_5515,N_5815);
and U6935 (N_6935,N_5311,N_5835);
xnor U6936 (N_6936,N_5272,N_5994);
or U6937 (N_6937,N_5710,N_5650);
nand U6938 (N_6938,N_5269,N_6195);
or U6939 (N_6939,N_5526,N_5678);
xor U6940 (N_6940,N_5326,N_5551);
nor U6941 (N_6941,N_5369,N_6172);
and U6942 (N_6942,N_5074,N_6019);
nand U6943 (N_6943,N_5691,N_6005);
or U6944 (N_6944,N_5105,N_6088);
nand U6945 (N_6945,N_5290,N_5537);
and U6946 (N_6946,N_5577,N_6170);
and U6947 (N_6947,N_6226,N_6023);
and U6948 (N_6948,N_5510,N_6197);
or U6949 (N_6949,N_5043,N_5946);
nor U6950 (N_6950,N_5295,N_5464);
or U6951 (N_6951,N_5490,N_6058);
nor U6952 (N_6952,N_5360,N_5833);
xor U6953 (N_6953,N_5973,N_6092);
xnor U6954 (N_6954,N_5811,N_5702);
xor U6955 (N_6955,N_6201,N_5261);
or U6956 (N_6956,N_6238,N_5808);
nand U6957 (N_6957,N_5798,N_5601);
and U6958 (N_6958,N_5407,N_5071);
xor U6959 (N_6959,N_5700,N_5315);
and U6960 (N_6960,N_5078,N_5761);
and U6961 (N_6961,N_5326,N_5412);
nor U6962 (N_6962,N_5233,N_6245);
or U6963 (N_6963,N_6169,N_5028);
nor U6964 (N_6964,N_5117,N_5802);
xnor U6965 (N_6965,N_5542,N_5605);
nor U6966 (N_6966,N_5435,N_5767);
and U6967 (N_6967,N_5303,N_6240);
or U6968 (N_6968,N_5672,N_5378);
nand U6969 (N_6969,N_5841,N_5186);
or U6970 (N_6970,N_5155,N_6053);
and U6971 (N_6971,N_5350,N_5487);
nor U6972 (N_6972,N_5909,N_5411);
and U6973 (N_6973,N_5007,N_5291);
and U6974 (N_6974,N_5694,N_5789);
nor U6975 (N_6975,N_5419,N_6128);
or U6976 (N_6976,N_5461,N_6001);
or U6977 (N_6977,N_5669,N_5202);
nor U6978 (N_6978,N_5134,N_5817);
nand U6979 (N_6979,N_6006,N_6234);
nand U6980 (N_6980,N_5753,N_5256);
nand U6981 (N_6981,N_5986,N_5459);
and U6982 (N_6982,N_5357,N_5408);
or U6983 (N_6983,N_5922,N_6084);
and U6984 (N_6984,N_5360,N_5951);
and U6985 (N_6985,N_6155,N_6149);
xor U6986 (N_6986,N_5721,N_5013);
nor U6987 (N_6987,N_5729,N_5139);
xnor U6988 (N_6988,N_5559,N_5660);
nor U6989 (N_6989,N_5988,N_5109);
nand U6990 (N_6990,N_5538,N_5324);
or U6991 (N_6991,N_5220,N_5975);
nor U6992 (N_6992,N_5030,N_5935);
xnor U6993 (N_6993,N_6232,N_5831);
xor U6994 (N_6994,N_5382,N_6075);
or U6995 (N_6995,N_5486,N_5643);
and U6996 (N_6996,N_5667,N_6017);
nand U6997 (N_6997,N_5356,N_5495);
nor U6998 (N_6998,N_5930,N_5497);
xnor U6999 (N_6999,N_5931,N_5401);
nor U7000 (N_7000,N_5034,N_5308);
nand U7001 (N_7001,N_5370,N_5725);
or U7002 (N_7002,N_5423,N_5220);
xor U7003 (N_7003,N_5856,N_5409);
nand U7004 (N_7004,N_5853,N_5505);
xor U7005 (N_7005,N_5211,N_5304);
xnor U7006 (N_7006,N_5012,N_5713);
xnor U7007 (N_7007,N_5139,N_5153);
or U7008 (N_7008,N_5747,N_5395);
or U7009 (N_7009,N_6083,N_5892);
nor U7010 (N_7010,N_5157,N_5767);
xnor U7011 (N_7011,N_5399,N_5121);
nand U7012 (N_7012,N_5149,N_5296);
xnor U7013 (N_7013,N_6038,N_6082);
and U7014 (N_7014,N_5521,N_5100);
nor U7015 (N_7015,N_5362,N_5017);
or U7016 (N_7016,N_5968,N_5904);
or U7017 (N_7017,N_6092,N_5777);
nor U7018 (N_7018,N_5498,N_5909);
nor U7019 (N_7019,N_5646,N_6059);
or U7020 (N_7020,N_6028,N_5323);
and U7021 (N_7021,N_5247,N_5003);
nand U7022 (N_7022,N_5267,N_6138);
xor U7023 (N_7023,N_5110,N_5642);
and U7024 (N_7024,N_6129,N_5140);
xor U7025 (N_7025,N_5819,N_5215);
xnor U7026 (N_7026,N_5281,N_5622);
nand U7027 (N_7027,N_6186,N_5421);
or U7028 (N_7028,N_5377,N_5296);
and U7029 (N_7029,N_5620,N_6235);
and U7030 (N_7030,N_5869,N_5701);
xnor U7031 (N_7031,N_5690,N_6217);
nand U7032 (N_7032,N_5038,N_5605);
and U7033 (N_7033,N_5333,N_5899);
nor U7034 (N_7034,N_6127,N_5984);
nand U7035 (N_7035,N_5647,N_6197);
nand U7036 (N_7036,N_5805,N_5747);
and U7037 (N_7037,N_5556,N_5636);
and U7038 (N_7038,N_5205,N_5570);
nand U7039 (N_7039,N_5824,N_5457);
and U7040 (N_7040,N_6104,N_5434);
nor U7041 (N_7041,N_5079,N_6059);
xnor U7042 (N_7042,N_5970,N_6046);
nor U7043 (N_7043,N_5690,N_5180);
xor U7044 (N_7044,N_5197,N_6115);
nand U7045 (N_7045,N_5378,N_5261);
xnor U7046 (N_7046,N_5724,N_6121);
xor U7047 (N_7047,N_5576,N_5117);
nor U7048 (N_7048,N_6076,N_5555);
or U7049 (N_7049,N_5770,N_5147);
xnor U7050 (N_7050,N_6044,N_5800);
nor U7051 (N_7051,N_5247,N_5495);
nand U7052 (N_7052,N_5280,N_5622);
nor U7053 (N_7053,N_5050,N_5808);
and U7054 (N_7054,N_5114,N_5942);
nand U7055 (N_7055,N_6144,N_5859);
and U7056 (N_7056,N_5315,N_5596);
nor U7057 (N_7057,N_5884,N_5816);
nand U7058 (N_7058,N_6215,N_5546);
or U7059 (N_7059,N_5763,N_6100);
and U7060 (N_7060,N_5267,N_5700);
nand U7061 (N_7061,N_5518,N_5269);
and U7062 (N_7062,N_5292,N_5373);
nor U7063 (N_7063,N_5285,N_5459);
nor U7064 (N_7064,N_5268,N_5352);
or U7065 (N_7065,N_5748,N_6054);
or U7066 (N_7066,N_5813,N_6011);
nand U7067 (N_7067,N_5858,N_5131);
nor U7068 (N_7068,N_6038,N_5838);
nand U7069 (N_7069,N_5898,N_5927);
and U7070 (N_7070,N_5873,N_5555);
xnor U7071 (N_7071,N_5687,N_5304);
nand U7072 (N_7072,N_5958,N_5145);
and U7073 (N_7073,N_6127,N_5673);
or U7074 (N_7074,N_5366,N_5959);
or U7075 (N_7075,N_5575,N_5920);
or U7076 (N_7076,N_5721,N_5903);
and U7077 (N_7077,N_5915,N_6071);
nand U7078 (N_7078,N_5191,N_5190);
nor U7079 (N_7079,N_5267,N_5454);
nor U7080 (N_7080,N_5047,N_5925);
or U7081 (N_7081,N_5845,N_5776);
and U7082 (N_7082,N_5263,N_6205);
or U7083 (N_7083,N_5434,N_6030);
nand U7084 (N_7084,N_5062,N_5898);
and U7085 (N_7085,N_5999,N_5768);
nor U7086 (N_7086,N_5864,N_5593);
nor U7087 (N_7087,N_5563,N_5490);
or U7088 (N_7088,N_5069,N_5702);
xor U7089 (N_7089,N_6060,N_5375);
or U7090 (N_7090,N_5154,N_6174);
nand U7091 (N_7091,N_5407,N_6114);
xor U7092 (N_7092,N_6103,N_5226);
nor U7093 (N_7093,N_5673,N_5018);
and U7094 (N_7094,N_5065,N_6065);
and U7095 (N_7095,N_5174,N_6079);
nand U7096 (N_7096,N_5636,N_5003);
or U7097 (N_7097,N_5996,N_5312);
nand U7098 (N_7098,N_5368,N_5687);
and U7099 (N_7099,N_6146,N_5598);
nor U7100 (N_7100,N_5495,N_5198);
nand U7101 (N_7101,N_5432,N_5503);
nand U7102 (N_7102,N_6097,N_5515);
nor U7103 (N_7103,N_5083,N_5143);
and U7104 (N_7104,N_6117,N_6038);
nor U7105 (N_7105,N_5857,N_5956);
nor U7106 (N_7106,N_5973,N_6039);
nand U7107 (N_7107,N_5308,N_5046);
nor U7108 (N_7108,N_5530,N_6091);
or U7109 (N_7109,N_6000,N_5602);
nand U7110 (N_7110,N_5993,N_5979);
or U7111 (N_7111,N_6073,N_5439);
xor U7112 (N_7112,N_5107,N_5500);
and U7113 (N_7113,N_5654,N_5235);
nor U7114 (N_7114,N_6007,N_6070);
or U7115 (N_7115,N_5083,N_5780);
xor U7116 (N_7116,N_5836,N_6101);
and U7117 (N_7117,N_5897,N_5760);
or U7118 (N_7118,N_5223,N_5559);
nand U7119 (N_7119,N_5779,N_5413);
and U7120 (N_7120,N_6245,N_5430);
or U7121 (N_7121,N_6034,N_5868);
nand U7122 (N_7122,N_5608,N_5743);
and U7123 (N_7123,N_5746,N_5113);
nor U7124 (N_7124,N_5084,N_5622);
nor U7125 (N_7125,N_5435,N_5898);
nor U7126 (N_7126,N_5034,N_5640);
or U7127 (N_7127,N_5758,N_6058);
xnor U7128 (N_7128,N_5606,N_5031);
xor U7129 (N_7129,N_6121,N_5125);
xor U7130 (N_7130,N_5187,N_5718);
nand U7131 (N_7131,N_5640,N_5301);
and U7132 (N_7132,N_5479,N_5534);
or U7133 (N_7133,N_5429,N_5692);
or U7134 (N_7134,N_6118,N_5485);
xor U7135 (N_7135,N_6180,N_5392);
and U7136 (N_7136,N_5177,N_5794);
nand U7137 (N_7137,N_5279,N_5645);
nor U7138 (N_7138,N_6115,N_5674);
or U7139 (N_7139,N_5660,N_5632);
and U7140 (N_7140,N_5957,N_5334);
nand U7141 (N_7141,N_5835,N_5870);
or U7142 (N_7142,N_5041,N_6201);
nor U7143 (N_7143,N_5217,N_6132);
or U7144 (N_7144,N_5566,N_5593);
xor U7145 (N_7145,N_5703,N_5718);
and U7146 (N_7146,N_5317,N_5095);
or U7147 (N_7147,N_5294,N_6024);
xnor U7148 (N_7148,N_5490,N_6110);
xor U7149 (N_7149,N_5343,N_6150);
nand U7150 (N_7150,N_5274,N_5070);
nand U7151 (N_7151,N_5293,N_6201);
xor U7152 (N_7152,N_5581,N_5272);
and U7153 (N_7153,N_6132,N_5590);
nor U7154 (N_7154,N_5520,N_5543);
xor U7155 (N_7155,N_5955,N_5735);
or U7156 (N_7156,N_6076,N_5211);
and U7157 (N_7157,N_5111,N_5886);
xnor U7158 (N_7158,N_5293,N_5365);
or U7159 (N_7159,N_5417,N_5813);
xnor U7160 (N_7160,N_5374,N_5641);
and U7161 (N_7161,N_5866,N_5868);
xor U7162 (N_7162,N_5028,N_5476);
nand U7163 (N_7163,N_5405,N_5516);
nand U7164 (N_7164,N_5159,N_5118);
xor U7165 (N_7165,N_6209,N_6167);
nand U7166 (N_7166,N_5751,N_5469);
nand U7167 (N_7167,N_6030,N_5854);
or U7168 (N_7168,N_5609,N_5680);
nand U7169 (N_7169,N_5898,N_5388);
or U7170 (N_7170,N_5766,N_5219);
or U7171 (N_7171,N_5688,N_6077);
or U7172 (N_7172,N_5877,N_6139);
or U7173 (N_7173,N_5195,N_6145);
xnor U7174 (N_7174,N_5262,N_5808);
nand U7175 (N_7175,N_5449,N_5383);
nand U7176 (N_7176,N_5129,N_5621);
nand U7177 (N_7177,N_5261,N_5287);
xnor U7178 (N_7178,N_6095,N_5491);
or U7179 (N_7179,N_5920,N_5122);
or U7180 (N_7180,N_5731,N_5221);
and U7181 (N_7181,N_6034,N_6058);
xnor U7182 (N_7182,N_5356,N_5917);
nand U7183 (N_7183,N_5677,N_5396);
or U7184 (N_7184,N_5702,N_6191);
nor U7185 (N_7185,N_5073,N_5003);
and U7186 (N_7186,N_5030,N_5446);
and U7187 (N_7187,N_5074,N_5281);
nand U7188 (N_7188,N_5212,N_5161);
or U7189 (N_7189,N_6124,N_5981);
and U7190 (N_7190,N_5841,N_5790);
nand U7191 (N_7191,N_5176,N_5813);
and U7192 (N_7192,N_5850,N_5467);
nand U7193 (N_7193,N_5296,N_5139);
nor U7194 (N_7194,N_5818,N_5586);
nor U7195 (N_7195,N_5770,N_5425);
and U7196 (N_7196,N_5670,N_6192);
xnor U7197 (N_7197,N_5477,N_6017);
and U7198 (N_7198,N_6096,N_5836);
or U7199 (N_7199,N_5233,N_5363);
nor U7200 (N_7200,N_5737,N_5575);
nor U7201 (N_7201,N_6218,N_5722);
and U7202 (N_7202,N_6211,N_5733);
or U7203 (N_7203,N_5537,N_5792);
nor U7204 (N_7204,N_6062,N_5787);
and U7205 (N_7205,N_5950,N_5688);
or U7206 (N_7206,N_5507,N_5056);
nand U7207 (N_7207,N_5978,N_5208);
or U7208 (N_7208,N_6081,N_6206);
or U7209 (N_7209,N_5684,N_5460);
xnor U7210 (N_7210,N_5846,N_5948);
nor U7211 (N_7211,N_5768,N_5172);
xnor U7212 (N_7212,N_6142,N_5957);
xor U7213 (N_7213,N_5996,N_5833);
xor U7214 (N_7214,N_5580,N_6112);
or U7215 (N_7215,N_6098,N_5281);
or U7216 (N_7216,N_6231,N_6217);
or U7217 (N_7217,N_5646,N_5527);
or U7218 (N_7218,N_5176,N_5276);
nor U7219 (N_7219,N_6029,N_6192);
xnor U7220 (N_7220,N_5758,N_6214);
and U7221 (N_7221,N_5940,N_5767);
and U7222 (N_7222,N_5102,N_5643);
nor U7223 (N_7223,N_6046,N_6128);
nand U7224 (N_7224,N_6223,N_6043);
xnor U7225 (N_7225,N_5229,N_5694);
nand U7226 (N_7226,N_6200,N_5648);
xor U7227 (N_7227,N_5418,N_5855);
or U7228 (N_7228,N_5880,N_5782);
and U7229 (N_7229,N_5679,N_5800);
xnor U7230 (N_7230,N_5799,N_5935);
nand U7231 (N_7231,N_5253,N_5121);
nor U7232 (N_7232,N_5890,N_5135);
xor U7233 (N_7233,N_6141,N_6049);
xnor U7234 (N_7234,N_5558,N_6071);
or U7235 (N_7235,N_5159,N_5212);
xor U7236 (N_7236,N_5254,N_5178);
and U7237 (N_7237,N_5479,N_5542);
nor U7238 (N_7238,N_5190,N_6244);
nor U7239 (N_7239,N_6136,N_5730);
nor U7240 (N_7240,N_5213,N_5783);
xnor U7241 (N_7241,N_5326,N_6048);
or U7242 (N_7242,N_5757,N_6026);
xor U7243 (N_7243,N_5299,N_5834);
nand U7244 (N_7244,N_6024,N_5541);
and U7245 (N_7245,N_5182,N_5534);
or U7246 (N_7246,N_5867,N_5205);
and U7247 (N_7247,N_5758,N_5227);
nand U7248 (N_7248,N_5733,N_5623);
or U7249 (N_7249,N_5857,N_5486);
nand U7250 (N_7250,N_6225,N_5752);
nand U7251 (N_7251,N_5302,N_5295);
or U7252 (N_7252,N_5103,N_5929);
xnor U7253 (N_7253,N_5084,N_5513);
nand U7254 (N_7254,N_6160,N_5018);
nand U7255 (N_7255,N_5879,N_6235);
nand U7256 (N_7256,N_6239,N_5469);
and U7257 (N_7257,N_6015,N_5794);
nand U7258 (N_7258,N_5056,N_5875);
and U7259 (N_7259,N_6209,N_5442);
nand U7260 (N_7260,N_5857,N_5784);
nand U7261 (N_7261,N_5325,N_6071);
nor U7262 (N_7262,N_5933,N_5626);
and U7263 (N_7263,N_6181,N_5494);
and U7264 (N_7264,N_6186,N_5268);
nor U7265 (N_7265,N_5137,N_5503);
and U7266 (N_7266,N_5507,N_5858);
or U7267 (N_7267,N_5143,N_5426);
and U7268 (N_7268,N_6100,N_5980);
or U7269 (N_7269,N_5796,N_5355);
nor U7270 (N_7270,N_6076,N_5907);
or U7271 (N_7271,N_5328,N_6079);
and U7272 (N_7272,N_5179,N_6175);
and U7273 (N_7273,N_5086,N_6119);
xnor U7274 (N_7274,N_5120,N_5409);
nor U7275 (N_7275,N_5330,N_5071);
or U7276 (N_7276,N_6082,N_5505);
nand U7277 (N_7277,N_5492,N_5388);
nor U7278 (N_7278,N_6246,N_5637);
nor U7279 (N_7279,N_5445,N_5298);
or U7280 (N_7280,N_5419,N_5388);
xnor U7281 (N_7281,N_5467,N_5772);
nand U7282 (N_7282,N_6035,N_5873);
or U7283 (N_7283,N_5358,N_5505);
xnor U7284 (N_7284,N_5964,N_5604);
or U7285 (N_7285,N_6015,N_5609);
xnor U7286 (N_7286,N_5334,N_6128);
xnor U7287 (N_7287,N_6065,N_5110);
xnor U7288 (N_7288,N_5182,N_5578);
nor U7289 (N_7289,N_5271,N_5934);
nor U7290 (N_7290,N_5924,N_6086);
or U7291 (N_7291,N_5746,N_5882);
xor U7292 (N_7292,N_5631,N_6047);
nor U7293 (N_7293,N_5086,N_5804);
xnor U7294 (N_7294,N_5693,N_5187);
or U7295 (N_7295,N_6197,N_5201);
nand U7296 (N_7296,N_5464,N_5895);
nor U7297 (N_7297,N_5609,N_5398);
or U7298 (N_7298,N_6085,N_5372);
nand U7299 (N_7299,N_5907,N_5750);
xor U7300 (N_7300,N_5421,N_5865);
xor U7301 (N_7301,N_6244,N_6051);
xnor U7302 (N_7302,N_5499,N_5008);
nand U7303 (N_7303,N_6013,N_5583);
nand U7304 (N_7304,N_5631,N_6086);
nor U7305 (N_7305,N_5428,N_5300);
nor U7306 (N_7306,N_6103,N_5852);
or U7307 (N_7307,N_6051,N_5140);
or U7308 (N_7308,N_5463,N_5112);
xnor U7309 (N_7309,N_5026,N_5229);
and U7310 (N_7310,N_5273,N_5747);
nand U7311 (N_7311,N_5624,N_5170);
nor U7312 (N_7312,N_5425,N_5136);
xnor U7313 (N_7313,N_5401,N_5740);
or U7314 (N_7314,N_6032,N_6074);
xnor U7315 (N_7315,N_5535,N_5899);
nor U7316 (N_7316,N_5811,N_5475);
xnor U7317 (N_7317,N_5726,N_5720);
or U7318 (N_7318,N_6189,N_5508);
nand U7319 (N_7319,N_5974,N_5268);
xor U7320 (N_7320,N_5710,N_5933);
or U7321 (N_7321,N_5953,N_5232);
xnor U7322 (N_7322,N_5244,N_5156);
xnor U7323 (N_7323,N_5325,N_6038);
or U7324 (N_7324,N_5767,N_5839);
and U7325 (N_7325,N_5108,N_5050);
nand U7326 (N_7326,N_5050,N_5900);
and U7327 (N_7327,N_5326,N_5698);
xnor U7328 (N_7328,N_5161,N_5488);
or U7329 (N_7329,N_5929,N_6008);
and U7330 (N_7330,N_6192,N_5941);
or U7331 (N_7331,N_6054,N_5299);
nor U7332 (N_7332,N_5033,N_5384);
or U7333 (N_7333,N_5420,N_5715);
xnor U7334 (N_7334,N_5868,N_6029);
nor U7335 (N_7335,N_6120,N_5086);
and U7336 (N_7336,N_5788,N_5690);
nand U7337 (N_7337,N_5412,N_5288);
or U7338 (N_7338,N_6164,N_5656);
or U7339 (N_7339,N_5889,N_5875);
or U7340 (N_7340,N_6236,N_5220);
nand U7341 (N_7341,N_5590,N_6018);
xor U7342 (N_7342,N_6008,N_5124);
or U7343 (N_7343,N_6016,N_5483);
nor U7344 (N_7344,N_5174,N_5471);
and U7345 (N_7345,N_5161,N_5554);
nor U7346 (N_7346,N_6165,N_5852);
and U7347 (N_7347,N_5708,N_5693);
nor U7348 (N_7348,N_5803,N_5567);
or U7349 (N_7349,N_5697,N_5688);
or U7350 (N_7350,N_5616,N_5452);
nand U7351 (N_7351,N_5178,N_5310);
or U7352 (N_7352,N_5443,N_5860);
or U7353 (N_7353,N_6154,N_6098);
or U7354 (N_7354,N_6191,N_5087);
nand U7355 (N_7355,N_5499,N_5984);
and U7356 (N_7356,N_5284,N_5471);
or U7357 (N_7357,N_6234,N_5277);
xnor U7358 (N_7358,N_5838,N_5591);
and U7359 (N_7359,N_5626,N_5321);
or U7360 (N_7360,N_5180,N_5560);
and U7361 (N_7361,N_5736,N_5471);
or U7362 (N_7362,N_5552,N_5701);
and U7363 (N_7363,N_5571,N_5838);
nand U7364 (N_7364,N_5370,N_6002);
nor U7365 (N_7365,N_6167,N_5946);
or U7366 (N_7366,N_5658,N_5619);
and U7367 (N_7367,N_5311,N_5738);
nand U7368 (N_7368,N_5247,N_5374);
nand U7369 (N_7369,N_6067,N_5936);
nor U7370 (N_7370,N_5697,N_5064);
and U7371 (N_7371,N_5414,N_5260);
nor U7372 (N_7372,N_5269,N_5953);
nand U7373 (N_7373,N_5178,N_6201);
and U7374 (N_7374,N_5386,N_5339);
nand U7375 (N_7375,N_5120,N_5718);
and U7376 (N_7376,N_5843,N_5501);
or U7377 (N_7377,N_5798,N_5075);
xnor U7378 (N_7378,N_6097,N_5957);
or U7379 (N_7379,N_6041,N_5986);
nor U7380 (N_7380,N_5972,N_5607);
nand U7381 (N_7381,N_5192,N_5169);
or U7382 (N_7382,N_5682,N_5258);
xor U7383 (N_7383,N_5802,N_5798);
or U7384 (N_7384,N_5288,N_5015);
xor U7385 (N_7385,N_5364,N_5010);
xnor U7386 (N_7386,N_5150,N_5838);
nor U7387 (N_7387,N_5515,N_5012);
nand U7388 (N_7388,N_5082,N_5406);
and U7389 (N_7389,N_6044,N_5418);
nand U7390 (N_7390,N_5294,N_5065);
nand U7391 (N_7391,N_6143,N_6132);
nand U7392 (N_7392,N_5814,N_5898);
and U7393 (N_7393,N_5563,N_5136);
xor U7394 (N_7394,N_5107,N_6176);
and U7395 (N_7395,N_5370,N_5277);
xor U7396 (N_7396,N_5482,N_5389);
nand U7397 (N_7397,N_5440,N_5500);
nor U7398 (N_7398,N_5085,N_5535);
nor U7399 (N_7399,N_6200,N_6093);
nor U7400 (N_7400,N_5691,N_6097);
xor U7401 (N_7401,N_5779,N_6180);
nor U7402 (N_7402,N_5965,N_5195);
nand U7403 (N_7403,N_5333,N_6168);
xnor U7404 (N_7404,N_5139,N_5888);
and U7405 (N_7405,N_5842,N_5408);
or U7406 (N_7406,N_5976,N_5430);
xnor U7407 (N_7407,N_5060,N_5033);
and U7408 (N_7408,N_5029,N_5107);
and U7409 (N_7409,N_5308,N_5740);
or U7410 (N_7410,N_5539,N_5315);
xnor U7411 (N_7411,N_5737,N_5447);
and U7412 (N_7412,N_6031,N_5320);
nor U7413 (N_7413,N_5595,N_5211);
and U7414 (N_7414,N_5690,N_5113);
or U7415 (N_7415,N_5472,N_6241);
or U7416 (N_7416,N_5763,N_5379);
xor U7417 (N_7417,N_5797,N_5759);
nand U7418 (N_7418,N_6139,N_6220);
nor U7419 (N_7419,N_5705,N_5462);
xnor U7420 (N_7420,N_6185,N_5952);
and U7421 (N_7421,N_5137,N_5641);
nand U7422 (N_7422,N_5353,N_5603);
and U7423 (N_7423,N_5330,N_6009);
nor U7424 (N_7424,N_5307,N_5860);
and U7425 (N_7425,N_5476,N_5151);
nor U7426 (N_7426,N_5115,N_5195);
nand U7427 (N_7427,N_5073,N_6246);
nor U7428 (N_7428,N_5860,N_5028);
xor U7429 (N_7429,N_5525,N_6001);
nor U7430 (N_7430,N_6086,N_6126);
or U7431 (N_7431,N_5887,N_5488);
xor U7432 (N_7432,N_5931,N_5010);
and U7433 (N_7433,N_5645,N_5633);
or U7434 (N_7434,N_5817,N_5751);
nand U7435 (N_7435,N_5562,N_6008);
xnor U7436 (N_7436,N_5176,N_5966);
nand U7437 (N_7437,N_6155,N_5221);
nand U7438 (N_7438,N_5475,N_5321);
nand U7439 (N_7439,N_6178,N_5914);
and U7440 (N_7440,N_5462,N_5662);
xor U7441 (N_7441,N_5077,N_5168);
and U7442 (N_7442,N_5267,N_5443);
xor U7443 (N_7443,N_5593,N_5921);
nor U7444 (N_7444,N_5229,N_5669);
nor U7445 (N_7445,N_6022,N_5976);
nand U7446 (N_7446,N_6041,N_5564);
and U7447 (N_7447,N_5413,N_5954);
nand U7448 (N_7448,N_6101,N_5640);
xor U7449 (N_7449,N_5279,N_5334);
or U7450 (N_7450,N_5175,N_5976);
or U7451 (N_7451,N_5880,N_6099);
nand U7452 (N_7452,N_5675,N_5769);
or U7453 (N_7453,N_6037,N_6020);
or U7454 (N_7454,N_5384,N_5995);
or U7455 (N_7455,N_6207,N_5508);
xor U7456 (N_7456,N_5966,N_5006);
nor U7457 (N_7457,N_5516,N_6058);
nor U7458 (N_7458,N_5859,N_5362);
xor U7459 (N_7459,N_5144,N_5833);
nand U7460 (N_7460,N_5310,N_5858);
and U7461 (N_7461,N_6116,N_6106);
and U7462 (N_7462,N_5040,N_5756);
xor U7463 (N_7463,N_5310,N_5615);
or U7464 (N_7464,N_6134,N_5176);
xnor U7465 (N_7465,N_5875,N_5807);
or U7466 (N_7466,N_5004,N_5803);
xor U7467 (N_7467,N_5472,N_5875);
or U7468 (N_7468,N_5541,N_5312);
and U7469 (N_7469,N_5674,N_5052);
nand U7470 (N_7470,N_5457,N_6170);
and U7471 (N_7471,N_5523,N_6230);
nor U7472 (N_7472,N_5533,N_5702);
nand U7473 (N_7473,N_5476,N_5383);
nor U7474 (N_7474,N_6035,N_5419);
or U7475 (N_7475,N_5047,N_5214);
nand U7476 (N_7476,N_6220,N_5614);
nand U7477 (N_7477,N_5278,N_5695);
xnor U7478 (N_7478,N_5730,N_5738);
xor U7479 (N_7479,N_5048,N_5918);
nand U7480 (N_7480,N_5245,N_6086);
xor U7481 (N_7481,N_5116,N_5159);
or U7482 (N_7482,N_5701,N_6189);
nor U7483 (N_7483,N_5076,N_5159);
nand U7484 (N_7484,N_5562,N_6109);
or U7485 (N_7485,N_5709,N_5550);
xor U7486 (N_7486,N_6020,N_6017);
and U7487 (N_7487,N_5530,N_5633);
nor U7488 (N_7488,N_5831,N_5513);
or U7489 (N_7489,N_6006,N_6163);
nand U7490 (N_7490,N_5560,N_5287);
or U7491 (N_7491,N_5419,N_5755);
nand U7492 (N_7492,N_5779,N_6021);
nor U7493 (N_7493,N_6147,N_5147);
or U7494 (N_7494,N_5635,N_5138);
nand U7495 (N_7495,N_5638,N_5878);
nor U7496 (N_7496,N_6174,N_5683);
and U7497 (N_7497,N_5696,N_5451);
nor U7498 (N_7498,N_5867,N_5690);
nor U7499 (N_7499,N_6024,N_5587);
nor U7500 (N_7500,N_7145,N_6486);
nand U7501 (N_7501,N_7417,N_7029);
or U7502 (N_7502,N_6583,N_7066);
or U7503 (N_7503,N_7074,N_7445);
and U7504 (N_7504,N_7405,N_6342);
xnor U7505 (N_7505,N_6551,N_6271);
or U7506 (N_7506,N_7050,N_7456);
xor U7507 (N_7507,N_6339,N_7449);
xnor U7508 (N_7508,N_6933,N_7304);
xnor U7509 (N_7509,N_6924,N_7305);
and U7510 (N_7510,N_7493,N_6672);
or U7511 (N_7511,N_6347,N_7184);
nand U7512 (N_7512,N_6594,N_7046);
nand U7513 (N_7513,N_7147,N_7261);
or U7514 (N_7514,N_6430,N_6791);
nand U7515 (N_7515,N_6429,N_6773);
nand U7516 (N_7516,N_6563,N_7220);
nor U7517 (N_7517,N_7152,N_6362);
xnor U7518 (N_7518,N_7331,N_7133);
xnor U7519 (N_7519,N_6971,N_6310);
nor U7520 (N_7520,N_6836,N_7019);
nor U7521 (N_7521,N_7059,N_6759);
or U7522 (N_7522,N_7093,N_6397);
nand U7523 (N_7523,N_6734,N_6522);
nor U7524 (N_7524,N_7287,N_6875);
nand U7525 (N_7525,N_7497,N_6585);
nand U7526 (N_7526,N_7276,N_6580);
and U7527 (N_7527,N_6958,N_7150);
or U7528 (N_7528,N_6846,N_6291);
nor U7529 (N_7529,N_6802,N_7372);
xor U7530 (N_7530,N_6957,N_7266);
or U7531 (N_7531,N_6649,N_6476);
nand U7532 (N_7532,N_6653,N_6976);
nand U7533 (N_7533,N_7325,N_6929);
or U7534 (N_7534,N_6609,N_6380);
nor U7535 (N_7535,N_7139,N_6900);
nor U7536 (N_7536,N_6326,N_6645);
nand U7537 (N_7537,N_6296,N_6788);
and U7538 (N_7538,N_6545,N_6889);
and U7539 (N_7539,N_7337,N_6252);
xor U7540 (N_7540,N_6543,N_7165);
and U7541 (N_7541,N_7267,N_7045);
and U7542 (N_7542,N_7191,N_7199);
or U7543 (N_7543,N_6518,N_6826);
nand U7544 (N_7544,N_7010,N_6473);
nor U7545 (N_7545,N_6573,N_6972);
or U7546 (N_7546,N_6620,N_7211);
nor U7547 (N_7547,N_6469,N_6870);
and U7548 (N_7548,N_6956,N_7469);
or U7549 (N_7549,N_6819,N_6657);
or U7550 (N_7550,N_7175,N_6570);
nand U7551 (N_7551,N_6992,N_7312);
and U7552 (N_7552,N_6696,N_7213);
and U7553 (N_7553,N_6415,N_6599);
xor U7554 (N_7554,N_6552,N_7064);
or U7555 (N_7555,N_6771,N_6315);
xor U7556 (N_7556,N_6717,N_6452);
nand U7557 (N_7557,N_6996,N_6745);
nor U7558 (N_7558,N_7376,N_6388);
or U7559 (N_7559,N_7039,N_6716);
nand U7560 (N_7560,N_6743,N_7072);
and U7561 (N_7561,N_6521,N_7016);
and U7562 (N_7562,N_6989,N_7244);
xnor U7563 (N_7563,N_6411,N_6911);
xor U7564 (N_7564,N_6309,N_6517);
or U7565 (N_7565,N_7056,N_7086);
nor U7566 (N_7566,N_6595,N_6891);
and U7567 (N_7567,N_7227,N_6634);
nor U7568 (N_7568,N_7311,N_6384);
and U7569 (N_7569,N_7142,N_7431);
nor U7570 (N_7570,N_7434,N_7430);
nor U7571 (N_7571,N_7128,N_7189);
and U7572 (N_7572,N_6779,N_6981);
nor U7573 (N_7573,N_7108,N_6554);
nand U7574 (N_7574,N_7452,N_6530);
xor U7575 (N_7575,N_7342,N_6343);
xor U7576 (N_7576,N_7300,N_6789);
nand U7577 (N_7577,N_7371,N_6269);
and U7578 (N_7578,N_6673,N_6772);
nand U7579 (N_7579,N_7296,N_7023);
or U7580 (N_7580,N_6753,N_7071);
nor U7581 (N_7581,N_7200,N_6508);
nand U7582 (N_7582,N_6709,N_6295);
and U7583 (N_7583,N_7381,N_6810);
or U7584 (N_7584,N_6421,N_6394);
nor U7585 (N_7585,N_6426,N_7454);
nand U7586 (N_7586,N_7030,N_6665);
xnor U7587 (N_7587,N_6861,N_6444);
nand U7588 (N_7588,N_7359,N_7309);
and U7589 (N_7589,N_6302,N_6336);
or U7590 (N_7590,N_7140,N_6379);
xnor U7591 (N_7591,N_6481,N_6671);
nand U7592 (N_7592,N_6766,N_7339);
or U7593 (N_7593,N_6726,N_6623);
or U7594 (N_7594,N_6281,N_7104);
nand U7595 (N_7595,N_7384,N_6507);
nor U7596 (N_7596,N_6414,N_7396);
nand U7597 (N_7597,N_7186,N_7317);
or U7598 (N_7598,N_6286,N_6393);
nand U7599 (N_7599,N_6450,N_7228);
nor U7600 (N_7600,N_6525,N_6806);
nor U7601 (N_7601,N_7097,N_6764);
nand U7602 (N_7602,N_7410,N_7033);
nor U7603 (N_7603,N_7051,N_6539);
or U7604 (N_7604,N_6356,N_6962);
and U7605 (N_7605,N_7096,N_6798);
xor U7606 (N_7606,N_7102,N_6495);
xnor U7607 (N_7607,N_6966,N_6320);
or U7608 (N_7608,N_6297,N_7391);
nand U7609 (N_7609,N_7185,N_7256);
xnor U7610 (N_7610,N_7241,N_7457);
and U7611 (N_7611,N_6496,N_6256);
nand U7612 (N_7612,N_7187,N_7323);
xor U7613 (N_7613,N_6809,N_6733);
xor U7614 (N_7614,N_6279,N_7301);
and U7615 (N_7615,N_7048,N_7057);
nor U7616 (N_7616,N_7069,N_6589);
nand U7617 (N_7617,N_6678,N_6558);
nand U7618 (N_7618,N_6600,N_7164);
nor U7619 (N_7619,N_6923,N_7310);
nor U7620 (N_7620,N_6794,N_7327);
or U7621 (N_7621,N_6333,N_6542);
nand U7622 (N_7622,N_6330,N_7487);
nand U7623 (N_7623,N_6782,N_6267);
xnor U7624 (N_7624,N_7407,N_7237);
nor U7625 (N_7625,N_6401,N_6964);
and U7626 (N_7626,N_6317,N_7049);
or U7627 (N_7627,N_7306,N_6830);
nand U7628 (N_7628,N_6675,N_7040);
xnor U7629 (N_7629,N_7465,N_6986);
xor U7630 (N_7630,N_6728,N_7078);
nor U7631 (N_7631,N_6775,N_6626);
and U7632 (N_7632,N_7247,N_6820);
xnor U7633 (N_7633,N_7460,N_7031);
and U7634 (N_7634,N_6953,N_7148);
and U7635 (N_7635,N_6456,N_7113);
or U7636 (N_7636,N_7014,N_7362);
or U7637 (N_7637,N_6372,N_6579);
nand U7638 (N_7638,N_6660,N_6284);
and U7639 (N_7639,N_6998,N_6916);
xor U7640 (N_7640,N_7171,N_6399);
and U7641 (N_7641,N_6859,N_6905);
xor U7642 (N_7642,N_7011,N_6804);
xor U7643 (N_7643,N_7238,N_6799);
nor U7644 (N_7644,N_6708,N_6698);
nor U7645 (N_7645,N_7271,N_7091);
or U7646 (N_7646,N_6361,N_6639);
xor U7647 (N_7647,N_6987,N_6959);
nor U7648 (N_7648,N_6529,N_7061);
xnor U7649 (N_7649,N_7421,N_7308);
and U7650 (N_7650,N_6607,N_6559);
and U7651 (N_7651,N_6458,N_7277);
nand U7652 (N_7652,N_6534,N_6305);
xor U7653 (N_7653,N_6723,N_6867);
xnor U7654 (N_7654,N_6774,N_6949);
or U7655 (N_7655,N_6781,N_7089);
nand U7656 (N_7656,N_7183,N_7122);
nor U7657 (N_7657,N_6541,N_7321);
or U7658 (N_7658,N_7005,N_6922);
xor U7659 (N_7659,N_6566,N_7341);
nand U7660 (N_7660,N_7024,N_7136);
xnor U7661 (N_7661,N_7118,N_6390);
and U7662 (N_7662,N_6635,N_7135);
xnor U7663 (N_7663,N_7115,N_6434);
xor U7664 (N_7664,N_6903,N_6669);
and U7665 (N_7665,N_7324,N_7217);
nor U7666 (N_7666,N_6686,N_6640);
nand U7667 (N_7667,N_6571,N_6879);
and U7668 (N_7668,N_6676,N_6970);
or U7669 (N_7669,N_6428,N_6370);
nand U7670 (N_7670,N_7218,N_7223);
or U7671 (N_7671,N_6294,N_6658);
nand U7672 (N_7672,N_6457,N_6837);
nand U7673 (N_7673,N_7022,N_7436);
nor U7674 (N_7674,N_7340,N_6690);
nand U7675 (N_7675,N_6502,N_6777);
xnor U7676 (N_7676,N_7475,N_7486);
nand U7677 (N_7677,N_6868,N_6722);
nand U7678 (N_7678,N_7007,N_7060);
xnor U7679 (N_7679,N_6387,N_6615);
or U7680 (N_7680,N_6472,N_7208);
xnor U7681 (N_7681,N_7485,N_6259);
xor U7682 (N_7682,N_6590,N_6625);
nand U7683 (N_7683,N_7044,N_6453);
nand U7684 (N_7684,N_6679,N_7418);
xnor U7685 (N_7685,N_7000,N_7105);
nand U7686 (N_7686,N_7178,N_7169);
and U7687 (N_7687,N_6459,N_6366);
nand U7688 (N_7688,N_6516,N_6492);
xnor U7689 (N_7689,N_6610,N_7110);
nand U7690 (N_7690,N_7215,N_7119);
xnor U7691 (N_7691,N_7289,N_6519);
nor U7692 (N_7692,N_6264,N_7193);
xnor U7693 (N_7693,N_6618,N_7077);
xor U7694 (N_7694,N_6700,N_7082);
or U7695 (N_7695,N_6955,N_6331);
nor U7696 (N_7696,N_7219,N_6592);
xnor U7697 (N_7697,N_6883,N_6694);
nor U7698 (N_7698,N_6852,N_6278);
or U7699 (N_7699,N_6392,N_6967);
nor U7700 (N_7700,N_7155,N_6944);
nand U7701 (N_7701,N_7131,N_7320);
nand U7702 (N_7702,N_6562,N_6300);
and U7703 (N_7703,N_6853,N_6695);
or U7704 (N_7704,N_6290,N_7288);
nand U7705 (N_7705,N_7390,N_6482);
xnor U7706 (N_7706,N_6783,N_6963);
nor U7707 (N_7707,N_7146,N_7173);
nor U7708 (N_7708,N_6556,N_6602);
nor U7709 (N_7709,N_6285,N_6800);
nand U7710 (N_7710,N_6896,N_6822);
or U7711 (N_7711,N_6767,N_7043);
xnor U7712 (N_7712,N_7166,N_6593);
nor U7713 (N_7713,N_6914,N_6376);
or U7714 (N_7714,N_6869,N_7402);
and U7715 (N_7715,N_6423,N_6437);
and U7716 (N_7716,N_6641,N_7470);
or U7717 (N_7717,N_6681,N_7283);
xnor U7718 (N_7718,N_6648,N_6514);
nor U7719 (N_7719,N_7443,N_6650);
nand U7720 (N_7720,N_7207,N_6877);
xnor U7721 (N_7721,N_6608,N_6311);
xor U7722 (N_7722,N_7176,N_7103);
xnor U7723 (N_7723,N_7035,N_6805);
nor U7724 (N_7724,N_6997,N_7290);
or U7725 (N_7725,N_7466,N_7388);
nor U7726 (N_7726,N_6991,N_7013);
or U7727 (N_7727,N_6646,N_7361);
nand U7728 (N_7728,N_6715,N_7326);
or U7729 (N_7729,N_6913,N_6439);
xnor U7730 (N_7730,N_7037,N_6280);
or U7731 (N_7731,N_6402,N_6849);
xnor U7732 (N_7732,N_6856,N_7251);
and U7733 (N_7733,N_6329,N_7157);
and U7734 (N_7734,N_7481,N_7280);
nand U7735 (N_7735,N_6301,N_7409);
nand U7736 (N_7736,N_7406,N_6843);
and U7737 (N_7737,N_7448,N_7275);
and U7738 (N_7738,N_6817,N_7236);
and U7739 (N_7739,N_7492,N_6501);
nand U7740 (N_7740,N_7479,N_6371);
xor U7741 (N_7741,N_6776,N_7412);
nor U7742 (N_7742,N_6282,N_7441);
nor U7743 (N_7743,N_6364,N_7243);
or U7744 (N_7744,N_7116,N_6928);
and U7745 (N_7745,N_6289,N_7248);
nor U7746 (N_7746,N_6627,N_6619);
and U7747 (N_7747,N_7447,N_6358);
xor U7748 (N_7748,N_7464,N_6898);
xnor U7749 (N_7749,N_6863,N_6498);
and U7750 (N_7750,N_7130,N_7225);
or U7751 (N_7751,N_7413,N_6744);
nand U7752 (N_7752,N_6666,N_6360);
nor U7753 (N_7753,N_6761,N_6951);
nor U7754 (N_7754,N_6835,N_7281);
nor U7755 (N_7755,N_6250,N_6613);
and U7756 (N_7756,N_6749,N_7451);
or U7757 (N_7757,N_7254,N_6720);
xnor U7758 (N_7758,N_7374,N_6467);
nand U7759 (N_7759,N_7137,N_6617);
and U7760 (N_7760,N_6885,N_7313);
or U7761 (N_7761,N_6793,N_6742);
nor U7762 (N_7762,N_6550,N_7279);
nor U7763 (N_7763,N_7174,N_6582);
or U7764 (N_7764,N_6438,N_7222);
or U7765 (N_7765,N_6480,N_7483);
or U7766 (N_7766,N_7335,N_6474);
or U7767 (N_7767,N_6866,N_6383);
xnor U7768 (N_7768,N_6265,N_7076);
and U7769 (N_7769,N_7012,N_7075);
nor U7770 (N_7770,N_6655,N_6834);
and U7771 (N_7771,N_6939,N_6892);
and U7772 (N_7772,N_6418,N_7387);
or U7773 (N_7773,N_7099,N_6621);
or U7774 (N_7774,N_6258,N_7003);
xor U7775 (N_7775,N_6765,N_6780);
nand U7776 (N_7776,N_7168,N_7004);
nand U7777 (N_7777,N_7363,N_6973);
nand U7778 (N_7778,N_6847,N_7239);
or U7779 (N_7779,N_6328,N_6803);
and U7780 (N_7780,N_6841,N_7274);
nor U7781 (N_7781,N_6901,N_7295);
nor U7782 (N_7782,N_6605,N_6493);
nor U7783 (N_7783,N_6864,N_6569);
nand U7784 (N_7784,N_7322,N_6851);
xor U7785 (N_7785,N_7260,N_6948);
nor U7786 (N_7786,N_6353,N_7214);
nand U7787 (N_7787,N_6536,N_7408);
nor U7788 (N_7788,N_7299,N_7425);
nor U7789 (N_7789,N_6833,N_6292);
or U7790 (N_7790,N_7333,N_7401);
nor U7791 (N_7791,N_7380,N_6752);
nand U7792 (N_7792,N_7230,N_6979);
and U7793 (N_7793,N_7411,N_7158);
or U7794 (N_7794,N_6389,N_7126);
or U7795 (N_7795,N_6446,N_6825);
xnor U7796 (N_7796,N_6829,N_7382);
or U7797 (N_7797,N_7491,N_6855);
xor U7798 (N_7798,N_7088,N_7375);
nand U7799 (N_7799,N_7291,N_7224);
nor U7800 (N_7800,N_6818,N_6832);
xor U7801 (N_7801,N_7458,N_6478);
or U7802 (N_7802,N_7083,N_7161);
and U7803 (N_7803,N_6980,N_6306);
nor U7804 (N_7804,N_6455,N_6369);
and U7805 (N_7805,N_6906,N_6577);
nand U7806 (N_7806,N_6701,N_6950);
nand U7807 (N_7807,N_7009,N_6413);
nand U7808 (N_7808,N_6425,N_7293);
nor U7809 (N_7809,N_7265,N_6448);
nand U7810 (N_7810,N_7285,N_6268);
and U7811 (N_7811,N_7478,N_6642);
nand U7812 (N_7812,N_6785,N_6858);
or U7813 (N_7813,N_7018,N_6688);
nand U7814 (N_7814,N_6930,N_6591);
or U7815 (N_7815,N_6643,N_6882);
xnor U7816 (N_7816,N_6266,N_6537);
and U7817 (N_7817,N_7393,N_6812);
nor U7818 (N_7818,N_7025,N_6895);
and U7819 (N_7819,N_6344,N_6598);
nand U7820 (N_7820,N_7006,N_7399);
nand U7821 (N_7821,N_6821,N_7038);
nor U7822 (N_7822,N_7453,N_7353);
xnor U7823 (N_7823,N_7355,N_6560);
xor U7824 (N_7824,N_6942,N_6433);
and U7825 (N_7825,N_6318,N_7428);
or U7826 (N_7826,N_6540,N_6662);
nand U7827 (N_7827,N_6523,N_6790);
nand U7828 (N_7828,N_7416,N_6897);
nand U7829 (N_7829,N_6629,N_6367);
or U7830 (N_7830,N_6597,N_6739);
and U7831 (N_7831,N_6547,N_7336);
and U7832 (N_7832,N_6403,N_7414);
or U7833 (N_7833,N_7160,N_6628);
nand U7834 (N_7834,N_6887,N_7002);
xnor U7835 (N_7835,N_7494,N_6422);
nand U7836 (N_7836,N_7346,N_7444);
and U7837 (N_7837,N_6878,N_6638);
nor U7838 (N_7838,N_7196,N_6324);
and U7839 (N_7839,N_7070,N_6873);
and U7840 (N_7840,N_7201,N_6750);
or U7841 (N_7841,N_6365,N_6985);
nor U7842 (N_7842,N_7149,N_7028);
and U7843 (N_7843,N_6952,N_6746);
nand U7844 (N_7844,N_6736,N_7440);
or U7845 (N_7845,N_6406,N_6975);
nor U7846 (N_7846,N_6575,N_6490);
nand U7847 (N_7847,N_6483,N_7182);
or U7848 (N_7848,N_6664,N_7472);
nor U7849 (N_7849,N_7482,N_6854);
nand U7850 (N_7850,N_7188,N_7107);
or U7851 (N_7851,N_6603,N_6352);
nand U7852 (N_7852,N_6647,N_7092);
nand U7853 (N_7853,N_7047,N_6661);
nand U7854 (N_7854,N_6355,N_6299);
and U7855 (N_7855,N_7360,N_7053);
nor U7856 (N_7856,N_7085,N_7204);
and U7857 (N_7857,N_7463,N_6886);
and U7858 (N_7858,N_6340,N_6656);
or U7859 (N_7859,N_6893,N_7245);
nand U7860 (N_7860,N_7419,N_6824);
nor U7861 (N_7861,N_6308,N_6586);
nor U7862 (N_7862,N_6533,N_6811);
or U7863 (N_7863,N_7383,N_7427);
xnor U7864 (N_7864,N_7143,N_7206);
xnor U7865 (N_7865,N_6351,N_7034);
xor U7866 (N_7866,N_7490,N_7259);
and U7867 (N_7867,N_6298,N_6935);
xor U7868 (N_7868,N_7471,N_6756);
or U7869 (N_7869,N_6348,N_7163);
or U7870 (N_7870,N_6815,N_6845);
xor U7871 (N_7871,N_7153,N_6663);
or U7872 (N_7872,N_7499,N_6479);
and U7873 (N_7873,N_6477,N_6270);
nand U7874 (N_7874,N_6451,N_6505);
and U7875 (N_7875,N_6961,N_6405);
nand U7876 (N_7876,N_6748,N_6398);
nor U7877 (N_7877,N_6601,N_7109);
or U7878 (N_7878,N_7235,N_7282);
nand U7879 (N_7879,N_6578,N_6506);
nor U7880 (N_7880,N_7209,N_7216);
xor U7881 (N_7881,N_7358,N_6727);
xnor U7882 (N_7882,N_6630,N_7151);
nand U7883 (N_7883,N_6564,N_7098);
xnor U7884 (N_7884,N_6524,N_6374);
nor U7885 (N_7885,N_7226,N_6947);
and U7886 (N_7886,N_6915,N_6707);
nor U7887 (N_7887,N_6614,N_6888);
nor U7888 (N_7888,N_6945,N_6710);
xnor U7889 (N_7889,N_6978,N_7258);
and U7890 (N_7890,N_6338,N_7292);
nor U7891 (N_7891,N_7015,N_6460);
nand U7892 (N_7892,N_7055,N_6632);
and U7893 (N_7893,N_7041,N_7087);
xnor U7894 (N_7894,N_6527,N_7307);
xnor U7895 (N_7895,N_6346,N_6463);
or U7896 (N_7896,N_6999,N_6737);
or U7897 (N_7897,N_6327,N_7008);
or U7898 (N_7898,N_6731,N_7488);
nand U7899 (N_7899,N_6936,N_6968);
and U7900 (N_7900,N_6862,N_6431);
or U7901 (N_7901,N_6497,N_6969);
nor U7902 (N_7902,N_7170,N_6488);
nand U7903 (N_7903,N_7262,N_7272);
or U7904 (N_7904,N_7273,N_7350);
and U7905 (N_7905,N_7474,N_6321);
and U7906 (N_7906,N_7446,N_7231);
or U7907 (N_7907,N_6555,N_6874);
xor U7908 (N_7908,N_6499,N_6485);
nor U7909 (N_7909,N_6946,N_7141);
and U7910 (N_7910,N_6357,N_6907);
nor U7911 (N_7911,N_6740,N_6509);
xor U7912 (N_7912,N_7080,N_7202);
xor U7913 (N_7913,N_7192,N_6561);
or U7914 (N_7914,N_6816,N_6526);
nand U7915 (N_7915,N_6407,N_6706);
and U7916 (N_7916,N_6738,N_7386);
and U7917 (N_7917,N_6719,N_6932);
xor U7918 (N_7918,N_6680,N_7229);
nand U7919 (N_7919,N_6751,N_6904);
and U7920 (N_7920,N_6844,N_7318);
nand U7921 (N_7921,N_6319,N_6382);
or U7922 (N_7922,N_6303,N_7400);
nor U7923 (N_7923,N_7462,N_7233);
nand U7924 (N_7924,N_7084,N_7450);
nor U7925 (N_7925,N_7398,N_7255);
and U7926 (N_7926,N_7438,N_7062);
xnor U7927 (N_7927,N_7194,N_6674);
xnor U7928 (N_7928,N_6400,N_7348);
nand U7929 (N_7929,N_6910,N_6977);
xor U7930 (N_7930,N_7268,N_6409);
xor U7931 (N_7931,N_6631,N_7422);
nor U7932 (N_7932,N_7101,N_6471);
xor U7933 (N_7933,N_7468,N_7354);
and U7934 (N_7934,N_6940,N_6462);
nand U7935 (N_7935,N_7352,N_6465);
nor U7936 (N_7936,N_6682,N_6274);
or U7937 (N_7937,N_7052,N_6865);
nand U7938 (N_7938,N_6652,N_6386);
xor U7939 (N_7939,N_6993,N_7332);
or U7940 (N_7940,N_7042,N_7370);
nor U7941 (N_7941,N_7439,N_6699);
or U7942 (N_7942,N_6718,N_7257);
and U7943 (N_7943,N_7121,N_6890);
xor U7944 (N_7944,N_6807,N_7392);
or U7945 (N_7945,N_7032,N_6612);
or U7946 (N_7946,N_6735,N_7058);
nor U7947 (N_7947,N_6795,N_6293);
nand U7948 (N_7948,N_7286,N_6454);
or U7949 (N_7949,N_6633,N_6500);
xor U7950 (N_7950,N_7394,N_6334);
xor U7951 (N_7951,N_7111,N_7476);
nand U7952 (N_7952,N_7036,N_6712);
nor U7953 (N_7953,N_6503,N_6729);
nand U7954 (N_7954,N_6762,N_6416);
nand U7955 (N_7955,N_7242,N_7349);
xnor U7956 (N_7956,N_7377,N_6322);
nor U7957 (N_7957,N_7095,N_6741);
nand U7958 (N_7958,N_6670,N_7156);
nor U7959 (N_7959,N_7437,N_7426);
or U7960 (N_7960,N_6732,N_6754);
and U7961 (N_7961,N_7298,N_7297);
and U7962 (N_7962,N_7269,N_7278);
and U7963 (N_7963,N_7403,N_7343);
and U7964 (N_7964,N_6801,N_7351);
nand U7965 (N_7965,N_6567,N_6814);
and U7966 (N_7966,N_6312,N_7210);
nor U7967 (N_7967,N_7435,N_6683);
or U7968 (N_7968,N_7344,N_6823);
xor U7969 (N_7969,N_6881,N_6902);
nand U7970 (N_7970,N_6994,N_6797);
or U7971 (N_7971,N_7079,N_7144);
and U7972 (N_7972,N_6468,N_7179);
or U7973 (N_7973,N_6515,N_6813);
nor U7974 (N_7974,N_6842,N_7369);
or U7975 (N_7975,N_6848,N_6395);
or U7976 (N_7976,N_6934,N_6404);
and U7977 (N_7977,N_6850,N_6624);
xnor U7978 (N_7978,N_6899,N_6553);
xor U7979 (N_7979,N_7270,N_6876);
xnor U7980 (N_7980,N_7132,N_6549);
nand U7981 (N_7981,N_6304,N_6769);
and U7982 (N_7982,N_6778,N_6325);
nor U7983 (N_7983,N_7180,N_6511);
xor U7984 (N_7984,N_6787,N_6381);
or U7985 (N_7985,N_6828,N_6919);
or U7986 (N_7986,N_6721,N_7316);
nor U7987 (N_7987,N_6894,N_6510);
nand U7988 (N_7988,N_6927,N_6960);
xor U7989 (N_7989,N_6713,N_7489);
xnor U7990 (N_7990,N_6359,N_6449);
nor U7991 (N_7991,N_6637,N_7404);
and U7992 (N_7992,N_6341,N_7159);
and U7993 (N_7993,N_7433,N_6984);
and U7994 (N_7994,N_6918,N_6692);
and U7995 (N_7995,N_6435,N_7424);
nor U7996 (N_7996,N_7415,N_6260);
xor U7997 (N_7997,N_7100,N_7389);
nor U7998 (N_7998,N_7420,N_6704);
and U7999 (N_7999,N_7345,N_6314);
nor U8000 (N_8000,N_6941,N_7094);
nor U8001 (N_8001,N_7197,N_6644);
nor U8002 (N_8002,N_6368,N_6484);
nor U8003 (N_8003,N_7246,N_7467);
nand U8004 (N_8004,N_7026,N_6757);
and U8005 (N_8005,N_7114,N_6349);
xnor U8006 (N_8006,N_6768,N_7252);
xor U8007 (N_8007,N_7240,N_6255);
nand U8008 (N_8008,N_6363,N_6931);
nor U8009 (N_8009,N_6375,N_6307);
or U8010 (N_8010,N_7017,N_6654);
or U8011 (N_8011,N_6831,N_6565);
nand U8012 (N_8012,N_6354,N_6316);
nand U8013 (N_8013,N_6687,N_7081);
nand U8014 (N_8014,N_6827,N_6667);
nand U8015 (N_8015,N_7330,N_6464);
nand U8016 (N_8016,N_7162,N_6588);
nand U8017 (N_8017,N_7063,N_6489);
nor U8018 (N_8018,N_7120,N_7395);
nor U8019 (N_8019,N_6396,N_6587);
nand U8020 (N_8020,N_7459,N_7021);
or U8021 (N_8021,N_6677,N_6335);
or U8022 (N_8022,N_6920,N_6763);
nor U8023 (N_8023,N_7379,N_7498);
or U8024 (N_8024,N_7328,N_6568);
nor U8025 (N_8025,N_6880,N_6792);
and U8026 (N_8026,N_7429,N_7397);
xnor U8027 (N_8027,N_7367,N_7368);
and U8028 (N_8028,N_7315,N_6703);
xnor U8029 (N_8029,N_6491,N_6995);
xor U8030 (N_8030,N_6659,N_6840);
and U8031 (N_8031,N_6276,N_7203);
xnor U8032 (N_8032,N_7181,N_6668);
or U8033 (N_8033,N_7067,N_7154);
xor U8034 (N_8034,N_6412,N_6584);
xnor U8035 (N_8035,N_6373,N_6513);
xnor U8036 (N_8036,N_6871,N_7378);
nor U8037 (N_8037,N_7338,N_6636);
nand U8038 (N_8038,N_7294,N_6436);
xor U8039 (N_8039,N_7167,N_6417);
xnor U8040 (N_8040,N_7117,N_7106);
nand U8041 (N_8041,N_7123,N_6747);
nand U8042 (N_8042,N_6912,N_7496);
and U8043 (N_8043,N_7190,N_7129);
nand U8044 (N_8044,N_7027,N_7090);
or U8045 (N_8045,N_6261,N_7329);
and U8046 (N_8046,N_6538,N_6684);
nand U8047 (N_8047,N_6937,N_6808);
nor U8048 (N_8048,N_6974,N_6611);
xor U8049 (N_8049,N_6725,N_6755);
nand U8050 (N_8050,N_6693,N_6410);
or U8051 (N_8051,N_6925,N_6254);
and U8052 (N_8052,N_6535,N_7373);
nand U8053 (N_8053,N_7134,N_7232);
nand U8054 (N_8054,N_6908,N_6424);
xnor U8055 (N_8055,N_6487,N_6954);
xor U8056 (N_8056,N_6758,N_7484);
and U8057 (N_8057,N_6943,N_6572);
or U8058 (N_8058,N_7172,N_7001);
xnor U8059 (N_8059,N_6714,N_6872);
xor U8060 (N_8060,N_6420,N_7249);
nor U8061 (N_8061,N_6504,N_6917);
nand U8062 (N_8062,N_7205,N_7480);
nand U8063 (N_8063,N_6251,N_6427);
nand U8064 (N_8064,N_6702,N_7138);
nand U8065 (N_8065,N_6983,N_6857);
and U8066 (N_8066,N_6273,N_6576);
or U8067 (N_8067,N_6786,N_6691);
nor U8068 (N_8068,N_7253,N_6884);
nand U8069 (N_8069,N_6283,N_7365);
xor U8070 (N_8070,N_6253,N_7356);
xor U8071 (N_8071,N_6685,N_7127);
or U8072 (N_8072,N_7221,N_6606);
or U8073 (N_8073,N_6622,N_7357);
xnor U8074 (N_8074,N_6377,N_6730);
nand U8075 (N_8075,N_7263,N_6548);
and U8076 (N_8076,N_6604,N_6796);
nor U8077 (N_8077,N_7264,N_6965);
nor U8078 (N_8078,N_7495,N_6461);
nand U8079 (N_8079,N_6345,N_7302);
nor U8080 (N_8080,N_6475,N_7432);
or U8081 (N_8081,N_6288,N_6350);
nand U8082 (N_8082,N_6990,N_7212);
nand U8083 (N_8083,N_6926,N_7125);
and U8084 (N_8084,N_6378,N_6440);
nand U8085 (N_8085,N_6544,N_7124);
nor U8086 (N_8086,N_6546,N_6512);
and U8087 (N_8087,N_7068,N_6470);
nor U8088 (N_8088,N_6557,N_6445);
and U8089 (N_8089,N_6528,N_7473);
or U8090 (N_8090,N_6262,N_7334);
or U8091 (N_8091,N_7250,N_6323);
xnor U8092 (N_8092,N_7477,N_7364);
nor U8093 (N_8093,N_6443,N_6494);
nor U8094 (N_8094,N_6581,N_6313);
or U8095 (N_8095,N_6596,N_6760);
nand U8096 (N_8096,N_6466,N_6574);
and U8097 (N_8097,N_7314,N_7054);
and U8098 (N_8098,N_7442,N_6337);
or U8099 (N_8099,N_7195,N_6921);
or U8100 (N_8100,N_6784,N_7198);
or U8101 (N_8101,N_6711,N_7112);
nand U8102 (N_8102,N_6432,N_7347);
nand U8103 (N_8103,N_7020,N_6705);
or U8104 (N_8104,N_6616,N_6839);
nor U8105 (N_8105,N_6408,N_6531);
nor U8106 (N_8106,N_6938,N_7423);
nor U8107 (N_8107,N_6332,N_6275);
or U8108 (N_8108,N_6272,N_6770);
nand U8109 (N_8109,N_7073,N_6447);
or U8110 (N_8110,N_6287,N_7284);
and U8111 (N_8111,N_6724,N_6697);
or U8112 (N_8112,N_6277,N_6860);
nand U8113 (N_8113,N_6982,N_6988);
and U8114 (N_8114,N_6532,N_6385);
and U8115 (N_8115,N_7234,N_7455);
nor U8116 (N_8116,N_6520,N_6391);
nand U8117 (N_8117,N_6689,N_7177);
xnor U8118 (N_8118,N_6441,N_6651);
nand U8119 (N_8119,N_6257,N_6442);
nand U8120 (N_8120,N_7303,N_7385);
nor U8121 (N_8121,N_7461,N_6909);
or U8122 (N_8122,N_7065,N_7366);
or U8123 (N_8123,N_6263,N_6838);
nand U8124 (N_8124,N_6419,N_7319);
xnor U8125 (N_8125,N_6499,N_7238);
nand U8126 (N_8126,N_6808,N_6923);
nand U8127 (N_8127,N_6410,N_7077);
nor U8128 (N_8128,N_6734,N_6356);
or U8129 (N_8129,N_6324,N_7189);
nand U8130 (N_8130,N_7209,N_6906);
xnor U8131 (N_8131,N_6354,N_7384);
or U8132 (N_8132,N_7050,N_6717);
or U8133 (N_8133,N_7395,N_7461);
or U8134 (N_8134,N_6497,N_6797);
and U8135 (N_8135,N_7413,N_7309);
nand U8136 (N_8136,N_6756,N_6560);
nor U8137 (N_8137,N_6918,N_6322);
or U8138 (N_8138,N_7075,N_6564);
nor U8139 (N_8139,N_6647,N_6861);
and U8140 (N_8140,N_6281,N_6524);
and U8141 (N_8141,N_7345,N_6458);
xnor U8142 (N_8142,N_7319,N_6473);
and U8143 (N_8143,N_6811,N_7362);
nor U8144 (N_8144,N_6520,N_7098);
or U8145 (N_8145,N_6565,N_6800);
xor U8146 (N_8146,N_6271,N_6379);
xor U8147 (N_8147,N_7176,N_7055);
xnor U8148 (N_8148,N_6297,N_7499);
nor U8149 (N_8149,N_6856,N_6764);
and U8150 (N_8150,N_6476,N_7393);
or U8151 (N_8151,N_6992,N_7402);
nand U8152 (N_8152,N_6899,N_7396);
nor U8153 (N_8153,N_7218,N_6443);
and U8154 (N_8154,N_6619,N_6917);
xor U8155 (N_8155,N_7136,N_6683);
nand U8156 (N_8156,N_6747,N_6306);
nand U8157 (N_8157,N_6524,N_7439);
nand U8158 (N_8158,N_6770,N_7023);
or U8159 (N_8159,N_6312,N_6663);
nor U8160 (N_8160,N_6948,N_6602);
xor U8161 (N_8161,N_7082,N_6484);
or U8162 (N_8162,N_6253,N_7368);
and U8163 (N_8163,N_6590,N_7388);
nand U8164 (N_8164,N_7206,N_6737);
nor U8165 (N_8165,N_7387,N_6633);
nor U8166 (N_8166,N_6581,N_6827);
and U8167 (N_8167,N_6824,N_6741);
or U8168 (N_8168,N_6937,N_7191);
or U8169 (N_8169,N_7483,N_7357);
nand U8170 (N_8170,N_6293,N_6768);
nand U8171 (N_8171,N_7165,N_7258);
or U8172 (N_8172,N_6570,N_6933);
or U8173 (N_8173,N_6266,N_6385);
nand U8174 (N_8174,N_7128,N_6597);
xor U8175 (N_8175,N_6338,N_7038);
xnor U8176 (N_8176,N_6773,N_6978);
or U8177 (N_8177,N_6891,N_6551);
nor U8178 (N_8178,N_6835,N_6435);
and U8179 (N_8179,N_7297,N_6866);
xnor U8180 (N_8180,N_6803,N_7333);
nand U8181 (N_8181,N_7279,N_6284);
nand U8182 (N_8182,N_7257,N_7065);
and U8183 (N_8183,N_6612,N_6962);
xor U8184 (N_8184,N_6935,N_7208);
xnor U8185 (N_8185,N_7321,N_7038);
nor U8186 (N_8186,N_6453,N_6866);
xor U8187 (N_8187,N_6936,N_6966);
or U8188 (N_8188,N_6657,N_7471);
and U8189 (N_8189,N_6901,N_6773);
nor U8190 (N_8190,N_7239,N_6572);
and U8191 (N_8191,N_6250,N_6529);
and U8192 (N_8192,N_6496,N_6820);
or U8193 (N_8193,N_7341,N_6426);
or U8194 (N_8194,N_7315,N_6564);
xnor U8195 (N_8195,N_7046,N_7020);
and U8196 (N_8196,N_6812,N_7351);
or U8197 (N_8197,N_6572,N_6933);
xor U8198 (N_8198,N_7482,N_6443);
and U8199 (N_8199,N_6740,N_7079);
or U8200 (N_8200,N_7088,N_6392);
or U8201 (N_8201,N_6535,N_7400);
xnor U8202 (N_8202,N_7067,N_7498);
nand U8203 (N_8203,N_7227,N_7118);
nand U8204 (N_8204,N_7367,N_7107);
nand U8205 (N_8205,N_6307,N_6911);
and U8206 (N_8206,N_7244,N_7042);
xor U8207 (N_8207,N_7241,N_7243);
nor U8208 (N_8208,N_6363,N_6849);
or U8209 (N_8209,N_6633,N_7128);
and U8210 (N_8210,N_7391,N_6861);
or U8211 (N_8211,N_6586,N_7475);
nand U8212 (N_8212,N_6382,N_6267);
nand U8213 (N_8213,N_6464,N_6397);
nor U8214 (N_8214,N_6830,N_6392);
nor U8215 (N_8215,N_7104,N_6309);
or U8216 (N_8216,N_7454,N_6796);
nor U8217 (N_8217,N_6413,N_7436);
xnor U8218 (N_8218,N_6886,N_6450);
nand U8219 (N_8219,N_7139,N_6281);
and U8220 (N_8220,N_7357,N_6883);
or U8221 (N_8221,N_6657,N_6469);
nor U8222 (N_8222,N_6435,N_6560);
and U8223 (N_8223,N_6257,N_7088);
or U8224 (N_8224,N_6597,N_7041);
or U8225 (N_8225,N_6662,N_6306);
nor U8226 (N_8226,N_6874,N_7338);
xnor U8227 (N_8227,N_7103,N_7081);
nor U8228 (N_8228,N_6582,N_7408);
xor U8229 (N_8229,N_6269,N_6679);
xnor U8230 (N_8230,N_6565,N_7303);
nor U8231 (N_8231,N_6361,N_6635);
xor U8232 (N_8232,N_7030,N_6727);
xor U8233 (N_8233,N_6272,N_7090);
nand U8234 (N_8234,N_6684,N_6381);
xor U8235 (N_8235,N_6791,N_6695);
nand U8236 (N_8236,N_6927,N_6867);
xnor U8237 (N_8237,N_7398,N_7464);
xnor U8238 (N_8238,N_6721,N_7117);
and U8239 (N_8239,N_6455,N_6265);
nor U8240 (N_8240,N_7162,N_6482);
and U8241 (N_8241,N_6514,N_6874);
xnor U8242 (N_8242,N_7194,N_6990);
xnor U8243 (N_8243,N_6762,N_6710);
or U8244 (N_8244,N_6847,N_6960);
nand U8245 (N_8245,N_7477,N_6683);
nor U8246 (N_8246,N_6382,N_6837);
nand U8247 (N_8247,N_6557,N_6834);
and U8248 (N_8248,N_6756,N_6860);
nand U8249 (N_8249,N_6998,N_6485);
nor U8250 (N_8250,N_7082,N_7460);
nand U8251 (N_8251,N_6513,N_7122);
nor U8252 (N_8252,N_6565,N_7482);
nand U8253 (N_8253,N_6456,N_7237);
and U8254 (N_8254,N_6448,N_7021);
xnor U8255 (N_8255,N_6310,N_6744);
xor U8256 (N_8256,N_7097,N_7380);
nand U8257 (N_8257,N_7318,N_6524);
and U8258 (N_8258,N_6271,N_6267);
xor U8259 (N_8259,N_6555,N_7205);
xor U8260 (N_8260,N_6326,N_6363);
nor U8261 (N_8261,N_6636,N_7199);
nand U8262 (N_8262,N_7247,N_6714);
nand U8263 (N_8263,N_6838,N_6827);
nor U8264 (N_8264,N_7345,N_7422);
xnor U8265 (N_8265,N_6404,N_6330);
nor U8266 (N_8266,N_6283,N_6291);
xnor U8267 (N_8267,N_6473,N_6485);
nand U8268 (N_8268,N_6685,N_7056);
xor U8269 (N_8269,N_6538,N_6670);
nand U8270 (N_8270,N_7065,N_6540);
or U8271 (N_8271,N_6365,N_7318);
nor U8272 (N_8272,N_6319,N_7343);
xor U8273 (N_8273,N_7016,N_6904);
or U8274 (N_8274,N_6730,N_7006);
xnor U8275 (N_8275,N_7281,N_6520);
and U8276 (N_8276,N_6997,N_6265);
or U8277 (N_8277,N_6545,N_7231);
nor U8278 (N_8278,N_6916,N_6991);
nor U8279 (N_8279,N_7364,N_7025);
nor U8280 (N_8280,N_6527,N_6476);
nand U8281 (N_8281,N_6588,N_6802);
nand U8282 (N_8282,N_6859,N_7390);
nand U8283 (N_8283,N_6593,N_7320);
nand U8284 (N_8284,N_7205,N_6548);
nand U8285 (N_8285,N_6331,N_7080);
xnor U8286 (N_8286,N_7108,N_6956);
and U8287 (N_8287,N_6557,N_6982);
nand U8288 (N_8288,N_6304,N_6334);
nor U8289 (N_8289,N_6810,N_7358);
and U8290 (N_8290,N_6823,N_6325);
xnor U8291 (N_8291,N_6485,N_6451);
nor U8292 (N_8292,N_6354,N_6835);
or U8293 (N_8293,N_6392,N_7069);
xnor U8294 (N_8294,N_7499,N_7400);
nand U8295 (N_8295,N_7440,N_7387);
and U8296 (N_8296,N_7196,N_6446);
and U8297 (N_8297,N_6616,N_7398);
and U8298 (N_8298,N_6613,N_6971);
or U8299 (N_8299,N_7399,N_7459);
and U8300 (N_8300,N_6421,N_6708);
or U8301 (N_8301,N_6922,N_6606);
nand U8302 (N_8302,N_6827,N_6320);
and U8303 (N_8303,N_6290,N_6414);
nor U8304 (N_8304,N_6845,N_7212);
xor U8305 (N_8305,N_7465,N_6505);
nor U8306 (N_8306,N_7089,N_6466);
nor U8307 (N_8307,N_6489,N_7347);
nor U8308 (N_8308,N_7163,N_6907);
xor U8309 (N_8309,N_6468,N_7304);
nand U8310 (N_8310,N_7434,N_6693);
and U8311 (N_8311,N_6644,N_7276);
and U8312 (N_8312,N_6884,N_6588);
and U8313 (N_8313,N_6393,N_6918);
and U8314 (N_8314,N_6764,N_6506);
or U8315 (N_8315,N_6444,N_6437);
nand U8316 (N_8316,N_7309,N_7439);
or U8317 (N_8317,N_7338,N_6680);
nor U8318 (N_8318,N_7362,N_6961);
or U8319 (N_8319,N_6618,N_7046);
nor U8320 (N_8320,N_6297,N_6692);
and U8321 (N_8321,N_6921,N_7227);
and U8322 (N_8322,N_7177,N_6356);
xnor U8323 (N_8323,N_7144,N_7446);
or U8324 (N_8324,N_6457,N_6382);
nor U8325 (N_8325,N_7230,N_6255);
xnor U8326 (N_8326,N_7148,N_7347);
nand U8327 (N_8327,N_6549,N_6485);
and U8328 (N_8328,N_7351,N_6950);
or U8329 (N_8329,N_6964,N_6867);
or U8330 (N_8330,N_6610,N_6951);
xnor U8331 (N_8331,N_7415,N_6932);
and U8332 (N_8332,N_6629,N_6368);
nand U8333 (N_8333,N_6436,N_7139);
xor U8334 (N_8334,N_6716,N_6342);
and U8335 (N_8335,N_6901,N_7237);
nand U8336 (N_8336,N_7020,N_7097);
and U8337 (N_8337,N_7180,N_6607);
nor U8338 (N_8338,N_6278,N_7011);
xor U8339 (N_8339,N_6419,N_7373);
or U8340 (N_8340,N_7383,N_6472);
nor U8341 (N_8341,N_7270,N_7437);
nand U8342 (N_8342,N_6920,N_6391);
xnor U8343 (N_8343,N_6325,N_7069);
xnor U8344 (N_8344,N_6639,N_7464);
xnor U8345 (N_8345,N_7381,N_7476);
and U8346 (N_8346,N_6528,N_6705);
nand U8347 (N_8347,N_6339,N_6750);
nor U8348 (N_8348,N_6481,N_6354);
or U8349 (N_8349,N_6280,N_7228);
or U8350 (N_8350,N_6256,N_6475);
nand U8351 (N_8351,N_7287,N_6667);
xnor U8352 (N_8352,N_7325,N_6917);
or U8353 (N_8353,N_7180,N_6314);
nor U8354 (N_8354,N_6589,N_6508);
xor U8355 (N_8355,N_6273,N_6833);
xor U8356 (N_8356,N_6312,N_6965);
nor U8357 (N_8357,N_7248,N_6515);
xor U8358 (N_8358,N_7016,N_6310);
or U8359 (N_8359,N_7499,N_7047);
xor U8360 (N_8360,N_6379,N_7459);
and U8361 (N_8361,N_7139,N_6936);
nor U8362 (N_8362,N_6685,N_7284);
nor U8363 (N_8363,N_7029,N_6312);
or U8364 (N_8364,N_7261,N_7331);
and U8365 (N_8365,N_6545,N_6968);
xor U8366 (N_8366,N_6852,N_7176);
nand U8367 (N_8367,N_7061,N_6659);
nand U8368 (N_8368,N_7294,N_6882);
and U8369 (N_8369,N_7123,N_7092);
nand U8370 (N_8370,N_7397,N_7244);
and U8371 (N_8371,N_6864,N_7040);
nand U8372 (N_8372,N_7113,N_6506);
nor U8373 (N_8373,N_7226,N_6581);
or U8374 (N_8374,N_7258,N_7348);
xor U8375 (N_8375,N_7093,N_6317);
or U8376 (N_8376,N_6446,N_7308);
nor U8377 (N_8377,N_6498,N_6611);
nor U8378 (N_8378,N_6982,N_6688);
xor U8379 (N_8379,N_7284,N_6402);
nand U8380 (N_8380,N_7304,N_6982);
or U8381 (N_8381,N_6829,N_6755);
or U8382 (N_8382,N_6661,N_6462);
and U8383 (N_8383,N_6963,N_6521);
xor U8384 (N_8384,N_7269,N_6859);
and U8385 (N_8385,N_7354,N_6355);
and U8386 (N_8386,N_6580,N_6404);
nor U8387 (N_8387,N_7313,N_6540);
nand U8388 (N_8388,N_7182,N_7249);
nand U8389 (N_8389,N_6488,N_7207);
nand U8390 (N_8390,N_6643,N_6779);
nor U8391 (N_8391,N_7256,N_6572);
xnor U8392 (N_8392,N_7071,N_6960);
nor U8393 (N_8393,N_6949,N_6735);
nand U8394 (N_8394,N_6874,N_6764);
nor U8395 (N_8395,N_6656,N_6487);
nand U8396 (N_8396,N_6776,N_6356);
nand U8397 (N_8397,N_6488,N_7480);
xor U8398 (N_8398,N_7367,N_7294);
xnor U8399 (N_8399,N_6312,N_7349);
and U8400 (N_8400,N_6419,N_6968);
nand U8401 (N_8401,N_7113,N_7424);
xor U8402 (N_8402,N_7393,N_7377);
and U8403 (N_8403,N_7222,N_6591);
xnor U8404 (N_8404,N_6348,N_6583);
xnor U8405 (N_8405,N_7300,N_7223);
or U8406 (N_8406,N_7093,N_6698);
or U8407 (N_8407,N_6272,N_6408);
nor U8408 (N_8408,N_6378,N_6517);
xnor U8409 (N_8409,N_6869,N_6544);
and U8410 (N_8410,N_6308,N_6657);
xnor U8411 (N_8411,N_6681,N_7056);
and U8412 (N_8412,N_6678,N_6583);
and U8413 (N_8413,N_7034,N_7334);
or U8414 (N_8414,N_6897,N_6278);
or U8415 (N_8415,N_6902,N_7011);
nand U8416 (N_8416,N_6874,N_7153);
and U8417 (N_8417,N_7093,N_7032);
and U8418 (N_8418,N_6848,N_7374);
xor U8419 (N_8419,N_7305,N_7230);
and U8420 (N_8420,N_7244,N_6348);
nand U8421 (N_8421,N_6796,N_7491);
or U8422 (N_8422,N_7301,N_6320);
or U8423 (N_8423,N_6940,N_6718);
or U8424 (N_8424,N_7150,N_6288);
or U8425 (N_8425,N_7308,N_6319);
and U8426 (N_8426,N_6860,N_6515);
and U8427 (N_8427,N_7185,N_6748);
nor U8428 (N_8428,N_7074,N_7465);
nand U8429 (N_8429,N_6442,N_7433);
nor U8430 (N_8430,N_7023,N_7223);
xor U8431 (N_8431,N_7053,N_7056);
and U8432 (N_8432,N_6636,N_6475);
nand U8433 (N_8433,N_6534,N_6752);
or U8434 (N_8434,N_7118,N_7273);
and U8435 (N_8435,N_7291,N_6560);
or U8436 (N_8436,N_6699,N_6731);
xor U8437 (N_8437,N_7485,N_7372);
xnor U8438 (N_8438,N_6433,N_6834);
and U8439 (N_8439,N_6536,N_6783);
nor U8440 (N_8440,N_6312,N_7092);
nor U8441 (N_8441,N_6946,N_6844);
nand U8442 (N_8442,N_7211,N_6680);
nor U8443 (N_8443,N_6886,N_7186);
nand U8444 (N_8444,N_7051,N_7286);
nor U8445 (N_8445,N_7010,N_6497);
or U8446 (N_8446,N_6915,N_6684);
nand U8447 (N_8447,N_6607,N_7284);
or U8448 (N_8448,N_6369,N_6308);
or U8449 (N_8449,N_6585,N_7379);
and U8450 (N_8450,N_6393,N_6982);
and U8451 (N_8451,N_6920,N_6930);
nor U8452 (N_8452,N_6724,N_7159);
nand U8453 (N_8453,N_6667,N_6578);
and U8454 (N_8454,N_7034,N_6369);
nand U8455 (N_8455,N_6911,N_6299);
nand U8456 (N_8456,N_6641,N_6257);
xnor U8457 (N_8457,N_7230,N_6330);
and U8458 (N_8458,N_7234,N_6976);
or U8459 (N_8459,N_6775,N_7213);
nor U8460 (N_8460,N_6675,N_7213);
nor U8461 (N_8461,N_6337,N_6687);
or U8462 (N_8462,N_7403,N_6354);
nand U8463 (N_8463,N_7411,N_7111);
nor U8464 (N_8464,N_6456,N_7435);
and U8465 (N_8465,N_7161,N_6250);
and U8466 (N_8466,N_7167,N_6489);
and U8467 (N_8467,N_6861,N_7015);
nor U8468 (N_8468,N_7444,N_6464);
and U8469 (N_8469,N_7192,N_7062);
nor U8470 (N_8470,N_6616,N_6902);
nand U8471 (N_8471,N_6980,N_6431);
nor U8472 (N_8472,N_6727,N_7106);
nand U8473 (N_8473,N_6461,N_6959);
xnor U8474 (N_8474,N_6685,N_6665);
or U8475 (N_8475,N_6572,N_7029);
xnor U8476 (N_8476,N_6846,N_7148);
or U8477 (N_8477,N_6301,N_7356);
and U8478 (N_8478,N_6270,N_7270);
and U8479 (N_8479,N_6595,N_6967);
xor U8480 (N_8480,N_7132,N_6974);
nand U8481 (N_8481,N_6641,N_7109);
and U8482 (N_8482,N_6459,N_6472);
and U8483 (N_8483,N_7146,N_7274);
or U8484 (N_8484,N_7068,N_6752);
or U8485 (N_8485,N_7235,N_6295);
nand U8486 (N_8486,N_6520,N_7308);
nand U8487 (N_8487,N_7395,N_7053);
and U8488 (N_8488,N_7495,N_6893);
xnor U8489 (N_8489,N_6344,N_7246);
nand U8490 (N_8490,N_6967,N_6454);
nor U8491 (N_8491,N_6937,N_6612);
nand U8492 (N_8492,N_7087,N_6796);
or U8493 (N_8493,N_6642,N_7226);
and U8494 (N_8494,N_6877,N_6696);
and U8495 (N_8495,N_6344,N_7361);
or U8496 (N_8496,N_6717,N_7394);
nor U8497 (N_8497,N_6316,N_6481);
nand U8498 (N_8498,N_6648,N_6372);
nand U8499 (N_8499,N_7187,N_7336);
nor U8500 (N_8500,N_6250,N_6740);
and U8501 (N_8501,N_6884,N_7036);
nand U8502 (N_8502,N_6310,N_7119);
and U8503 (N_8503,N_6331,N_6799);
and U8504 (N_8504,N_6939,N_7345);
nor U8505 (N_8505,N_7172,N_6734);
or U8506 (N_8506,N_6264,N_6490);
nand U8507 (N_8507,N_6928,N_6978);
or U8508 (N_8508,N_6630,N_6984);
nor U8509 (N_8509,N_7210,N_6618);
nor U8510 (N_8510,N_7458,N_7381);
and U8511 (N_8511,N_6693,N_6657);
nand U8512 (N_8512,N_6263,N_6580);
and U8513 (N_8513,N_7407,N_7039);
nand U8514 (N_8514,N_6272,N_6799);
and U8515 (N_8515,N_6391,N_6957);
xnor U8516 (N_8516,N_6762,N_7418);
xnor U8517 (N_8517,N_6833,N_7384);
and U8518 (N_8518,N_7056,N_7129);
and U8519 (N_8519,N_6633,N_7099);
or U8520 (N_8520,N_7408,N_6883);
nor U8521 (N_8521,N_6725,N_6599);
xnor U8522 (N_8522,N_7165,N_7175);
and U8523 (N_8523,N_6705,N_7485);
nand U8524 (N_8524,N_6280,N_7466);
nor U8525 (N_8525,N_7448,N_6618);
and U8526 (N_8526,N_7212,N_7216);
xnor U8527 (N_8527,N_7109,N_7232);
xor U8528 (N_8528,N_7399,N_7069);
or U8529 (N_8529,N_6375,N_6627);
xor U8530 (N_8530,N_6447,N_6861);
nor U8531 (N_8531,N_7077,N_6911);
xnor U8532 (N_8532,N_6611,N_7250);
nand U8533 (N_8533,N_6563,N_7247);
nand U8534 (N_8534,N_6536,N_6846);
or U8535 (N_8535,N_6727,N_6521);
nand U8536 (N_8536,N_7121,N_6710);
xnor U8537 (N_8537,N_7182,N_6830);
or U8538 (N_8538,N_6737,N_7153);
xor U8539 (N_8539,N_6823,N_7052);
nor U8540 (N_8540,N_6770,N_7033);
and U8541 (N_8541,N_6690,N_6862);
nor U8542 (N_8542,N_6398,N_6504);
nand U8543 (N_8543,N_6964,N_6558);
nand U8544 (N_8544,N_6363,N_7351);
or U8545 (N_8545,N_6431,N_7164);
or U8546 (N_8546,N_7238,N_6875);
xor U8547 (N_8547,N_7162,N_6645);
or U8548 (N_8548,N_7499,N_7381);
or U8549 (N_8549,N_6421,N_7206);
or U8550 (N_8550,N_6434,N_6312);
and U8551 (N_8551,N_6851,N_6876);
nand U8552 (N_8552,N_6673,N_6830);
nand U8553 (N_8553,N_7183,N_7043);
nand U8554 (N_8554,N_6516,N_7251);
xnor U8555 (N_8555,N_6931,N_6980);
nand U8556 (N_8556,N_7419,N_7132);
and U8557 (N_8557,N_6705,N_6296);
xor U8558 (N_8558,N_7009,N_6876);
nand U8559 (N_8559,N_6252,N_6505);
nand U8560 (N_8560,N_7111,N_6780);
and U8561 (N_8561,N_6694,N_6493);
xor U8562 (N_8562,N_6788,N_6987);
nand U8563 (N_8563,N_6265,N_6980);
and U8564 (N_8564,N_7341,N_7127);
or U8565 (N_8565,N_6461,N_7244);
nand U8566 (N_8566,N_6510,N_7034);
nand U8567 (N_8567,N_6346,N_6310);
xnor U8568 (N_8568,N_6827,N_7003);
xor U8569 (N_8569,N_7251,N_7127);
and U8570 (N_8570,N_6728,N_6600);
nor U8571 (N_8571,N_7072,N_6338);
xnor U8572 (N_8572,N_6883,N_7267);
or U8573 (N_8573,N_7298,N_6338);
or U8574 (N_8574,N_6403,N_7256);
xor U8575 (N_8575,N_7367,N_6259);
nand U8576 (N_8576,N_7407,N_6445);
nand U8577 (N_8577,N_7359,N_6816);
and U8578 (N_8578,N_7487,N_6846);
xor U8579 (N_8579,N_6821,N_6618);
xor U8580 (N_8580,N_6609,N_6730);
and U8581 (N_8581,N_6327,N_7319);
nand U8582 (N_8582,N_7160,N_7153);
and U8583 (N_8583,N_6963,N_7347);
nor U8584 (N_8584,N_7241,N_6998);
or U8585 (N_8585,N_6580,N_7061);
xor U8586 (N_8586,N_6906,N_6763);
xor U8587 (N_8587,N_6840,N_7139);
or U8588 (N_8588,N_6750,N_6573);
and U8589 (N_8589,N_6516,N_6868);
and U8590 (N_8590,N_6408,N_6637);
nor U8591 (N_8591,N_7460,N_6831);
nand U8592 (N_8592,N_6492,N_7234);
and U8593 (N_8593,N_6779,N_6352);
nor U8594 (N_8594,N_7464,N_7321);
nor U8595 (N_8595,N_6323,N_6331);
xor U8596 (N_8596,N_7456,N_6458);
xor U8597 (N_8597,N_7235,N_7089);
nand U8598 (N_8598,N_6303,N_7494);
or U8599 (N_8599,N_6482,N_7276);
and U8600 (N_8600,N_6566,N_6269);
or U8601 (N_8601,N_6993,N_6933);
and U8602 (N_8602,N_6660,N_7436);
or U8603 (N_8603,N_7493,N_6719);
nand U8604 (N_8604,N_7224,N_7319);
nor U8605 (N_8605,N_6504,N_6848);
or U8606 (N_8606,N_7258,N_6277);
nor U8607 (N_8607,N_7155,N_7371);
nor U8608 (N_8608,N_6840,N_7181);
xnor U8609 (N_8609,N_6296,N_6443);
or U8610 (N_8610,N_7493,N_6737);
xor U8611 (N_8611,N_7323,N_6341);
nand U8612 (N_8612,N_6558,N_6895);
or U8613 (N_8613,N_6543,N_7498);
nand U8614 (N_8614,N_6308,N_6594);
xnor U8615 (N_8615,N_6507,N_7255);
or U8616 (N_8616,N_6855,N_6703);
nand U8617 (N_8617,N_7306,N_7157);
or U8618 (N_8618,N_7320,N_7050);
or U8619 (N_8619,N_6292,N_6257);
nor U8620 (N_8620,N_6541,N_6255);
and U8621 (N_8621,N_7122,N_6512);
xnor U8622 (N_8622,N_7485,N_6747);
nand U8623 (N_8623,N_6635,N_6349);
and U8624 (N_8624,N_6724,N_7349);
nand U8625 (N_8625,N_7292,N_6343);
nor U8626 (N_8626,N_7377,N_6757);
nor U8627 (N_8627,N_6954,N_7441);
and U8628 (N_8628,N_6364,N_6387);
nand U8629 (N_8629,N_7340,N_6643);
xor U8630 (N_8630,N_6691,N_7196);
and U8631 (N_8631,N_6656,N_6914);
or U8632 (N_8632,N_6731,N_6622);
or U8633 (N_8633,N_6609,N_6735);
or U8634 (N_8634,N_7017,N_7374);
nand U8635 (N_8635,N_7477,N_6608);
xnor U8636 (N_8636,N_6316,N_6742);
nor U8637 (N_8637,N_7244,N_6846);
nand U8638 (N_8638,N_6649,N_7241);
nand U8639 (N_8639,N_6907,N_6999);
xor U8640 (N_8640,N_6978,N_6270);
nor U8641 (N_8641,N_7391,N_6446);
and U8642 (N_8642,N_6359,N_7408);
and U8643 (N_8643,N_6900,N_7315);
or U8644 (N_8644,N_7347,N_6604);
xnor U8645 (N_8645,N_7418,N_7458);
and U8646 (N_8646,N_7378,N_6669);
and U8647 (N_8647,N_7179,N_6809);
nand U8648 (N_8648,N_7311,N_6767);
or U8649 (N_8649,N_7121,N_7073);
or U8650 (N_8650,N_6514,N_6766);
nor U8651 (N_8651,N_6444,N_7143);
nor U8652 (N_8652,N_6912,N_6511);
xnor U8653 (N_8653,N_7366,N_6897);
xnor U8654 (N_8654,N_6282,N_6767);
or U8655 (N_8655,N_6407,N_6957);
nand U8656 (N_8656,N_7321,N_6655);
and U8657 (N_8657,N_6545,N_6326);
and U8658 (N_8658,N_7201,N_7170);
and U8659 (N_8659,N_7383,N_7135);
nor U8660 (N_8660,N_6820,N_6793);
xor U8661 (N_8661,N_7029,N_6844);
nand U8662 (N_8662,N_6307,N_7187);
nor U8663 (N_8663,N_6528,N_7068);
and U8664 (N_8664,N_6790,N_6642);
or U8665 (N_8665,N_6296,N_6691);
nand U8666 (N_8666,N_7352,N_7276);
or U8667 (N_8667,N_6962,N_6770);
xor U8668 (N_8668,N_7391,N_6621);
xor U8669 (N_8669,N_7440,N_6641);
and U8670 (N_8670,N_6289,N_6483);
nand U8671 (N_8671,N_7219,N_7109);
or U8672 (N_8672,N_6591,N_6999);
nor U8673 (N_8673,N_7331,N_6427);
xnor U8674 (N_8674,N_6973,N_6999);
xor U8675 (N_8675,N_6355,N_7391);
or U8676 (N_8676,N_6903,N_7092);
and U8677 (N_8677,N_6367,N_7161);
and U8678 (N_8678,N_6818,N_6892);
nor U8679 (N_8679,N_7395,N_6892);
nand U8680 (N_8680,N_7197,N_6302);
xor U8681 (N_8681,N_6812,N_7386);
nor U8682 (N_8682,N_6585,N_7378);
and U8683 (N_8683,N_7348,N_6265);
xor U8684 (N_8684,N_7294,N_6983);
nor U8685 (N_8685,N_7288,N_7056);
xor U8686 (N_8686,N_7024,N_6552);
xor U8687 (N_8687,N_7290,N_6992);
xor U8688 (N_8688,N_6386,N_6479);
or U8689 (N_8689,N_7270,N_6710);
nand U8690 (N_8690,N_6712,N_7193);
nand U8691 (N_8691,N_6808,N_7203);
nor U8692 (N_8692,N_7044,N_6862);
or U8693 (N_8693,N_6643,N_7224);
nand U8694 (N_8694,N_6275,N_7299);
and U8695 (N_8695,N_6694,N_7357);
and U8696 (N_8696,N_6725,N_6825);
and U8697 (N_8697,N_7155,N_6409);
and U8698 (N_8698,N_6370,N_7220);
and U8699 (N_8699,N_6916,N_6958);
and U8700 (N_8700,N_6336,N_6419);
nor U8701 (N_8701,N_7284,N_6986);
nor U8702 (N_8702,N_6716,N_7123);
and U8703 (N_8703,N_7450,N_6787);
nand U8704 (N_8704,N_7100,N_6958);
or U8705 (N_8705,N_6999,N_7336);
nand U8706 (N_8706,N_6296,N_7223);
and U8707 (N_8707,N_6839,N_6954);
nand U8708 (N_8708,N_6893,N_7097);
and U8709 (N_8709,N_7157,N_7404);
or U8710 (N_8710,N_7219,N_6907);
nand U8711 (N_8711,N_7379,N_6313);
xor U8712 (N_8712,N_7041,N_6678);
or U8713 (N_8713,N_6677,N_6406);
or U8714 (N_8714,N_7294,N_7299);
or U8715 (N_8715,N_6885,N_7275);
or U8716 (N_8716,N_6907,N_6901);
or U8717 (N_8717,N_6968,N_7026);
xnor U8718 (N_8718,N_6985,N_6696);
nor U8719 (N_8719,N_6459,N_7259);
nand U8720 (N_8720,N_7084,N_6980);
nand U8721 (N_8721,N_6544,N_6966);
nand U8722 (N_8722,N_7180,N_6689);
xnor U8723 (N_8723,N_7479,N_6266);
and U8724 (N_8724,N_7061,N_6878);
xor U8725 (N_8725,N_6623,N_6382);
xnor U8726 (N_8726,N_7298,N_7014);
nand U8727 (N_8727,N_7348,N_7442);
nand U8728 (N_8728,N_7203,N_6977);
or U8729 (N_8729,N_6906,N_6603);
or U8730 (N_8730,N_6482,N_6273);
nand U8731 (N_8731,N_6577,N_7017);
xnor U8732 (N_8732,N_7202,N_6920);
nand U8733 (N_8733,N_6649,N_7095);
nand U8734 (N_8734,N_7456,N_7132);
xor U8735 (N_8735,N_6948,N_6920);
xor U8736 (N_8736,N_7411,N_7125);
or U8737 (N_8737,N_6629,N_7089);
nand U8738 (N_8738,N_6536,N_6541);
nand U8739 (N_8739,N_6425,N_6901);
nor U8740 (N_8740,N_6583,N_7058);
nor U8741 (N_8741,N_7258,N_6595);
and U8742 (N_8742,N_6399,N_7378);
nor U8743 (N_8743,N_6334,N_6546);
nor U8744 (N_8744,N_6944,N_6539);
nand U8745 (N_8745,N_6696,N_6259);
and U8746 (N_8746,N_7239,N_7462);
nand U8747 (N_8747,N_6396,N_7420);
or U8748 (N_8748,N_6679,N_7336);
xnor U8749 (N_8749,N_6521,N_6702);
and U8750 (N_8750,N_8719,N_8384);
and U8751 (N_8751,N_8121,N_7940);
nand U8752 (N_8752,N_8674,N_8311);
xor U8753 (N_8753,N_8471,N_7696);
nand U8754 (N_8754,N_8458,N_8456);
nor U8755 (N_8755,N_8481,N_8747);
nor U8756 (N_8756,N_7870,N_7664);
and U8757 (N_8757,N_7902,N_7653);
nor U8758 (N_8758,N_7500,N_8109);
xnor U8759 (N_8759,N_7869,N_8163);
and U8760 (N_8760,N_8137,N_7674);
nand U8761 (N_8761,N_7603,N_8687);
xnor U8762 (N_8762,N_7876,N_8556);
xnor U8763 (N_8763,N_8020,N_7969);
xor U8764 (N_8764,N_8124,N_7544);
nor U8765 (N_8765,N_7518,N_8247);
xnor U8766 (N_8766,N_8675,N_8062);
or U8767 (N_8767,N_8573,N_7974);
xnor U8768 (N_8768,N_7889,N_8451);
nand U8769 (N_8769,N_7853,N_8141);
nand U8770 (N_8770,N_8161,N_7545);
or U8771 (N_8771,N_8391,N_7846);
nor U8772 (N_8772,N_7875,N_8206);
and U8773 (N_8773,N_8363,N_7935);
nor U8774 (N_8774,N_7807,N_7893);
and U8775 (N_8775,N_7560,N_8192);
nand U8776 (N_8776,N_7933,N_7977);
or U8777 (N_8777,N_7826,N_7612);
nor U8778 (N_8778,N_8144,N_8092);
and U8779 (N_8779,N_7712,N_7700);
nor U8780 (N_8780,N_7804,N_8531);
nand U8781 (N_8781,N_8592,N_8389);
nor U8782 (N_8782,N_8193,N_7947);
and U8783 (N_8783,N_7963,N_7620);
and U8784 (N_8784,N_7583,N_8671);
xor U8785 (N_8785,N_8469,N_8076);
or U8786 (N_8786,N_8231,N_7618);
xor U8787 (N_8787,N_8105,N_8640);
nand U8788 (N_8788,N_8194,N_7514);
and U8789 (N_8789,N_8511,N_7646);
xor U8790 (N_8790,N_8225,N_7801);
nor U8791 (N_8791,N_8061,N_8660);
or U8792 (N_8792,N_7625,N_8632);
nor U8793 (N_8793,N_8348,N_8122);
nor U8794 (N_8794,N_7591,N_8084);
xnor U8795 (N_8795,N_8078,N_7719);
xnor U8796 (N_8796,N_8744,N_8568);
nand U8797 (N_8797,N_8284,N_8228);
or U8798 (N_8798,N_8606,N_7636);
nand U8799 (N_8799,N_8641,N_7578);
and U8800 (N_8800,N_8642,N_8296);
or U8801 (N_8801,N_7989,N_8443);
or U8802 (N_8802,N_8631,N_8026);
nand U8803 (N_8803,N_8306,N_8737);
xnor U8804 (N_8804,N_7951,N_8167);
and U8805 (N_8805,N_8169,N_8683);
nand U8806 (N_8806,N_7557,N_7827);
xnor U8807 (N_8807,N_8003,N_7526);
nor U8808 (N_8808,N_7914,N_7967);
and U8809 (N_8809,N_7856,N_7930);
nand U8810 (N_8810,N_7589,N_8682);
or U8811 (N_8811,N_8620,N_7608);
nand U8812 (N_8812,N_8037,N_8523);
nor U8813 (N_8813,N_8290,N_7550);
and U8814 (N_8814,N_8328,N_7692);
nand U8815 (N_8815,N_7873,N_8442);
nor U8816 (N_8816,N_8318,N_8224);
nor U8817 (N_8817,N_7723,N_8381);
and U8818 (N_8818,N_8221,N_7927);
nor U8819 (N_8819,N_7568,N_7602);
nor U8820 (N_8820,N_8411,N_8291);
nand U8821 (N_8821,N_8212,N_7971);
and U8822 (N_8822,N_8689,N_8204);
nor U8823 (N_8823,N_8602,N_8482);
nor U8824 (N_8824,N_7781,N_8582);
or U8825 (N_8825,N_7616,N_7736);
or U8826 (N_8826,N_8370,N_8255);
nor U8827 (N_8827,N_7507,N_7813);
nand U8828 (N_8828,N_7740,N_8388);
or U8829 (N_8829,N_7837,N_7996);
nand U8830 (N_8830,N_8303,N_7660);
nand U8831 (N_8831,N_7650,N_8168);
nor U8832 (N_8832,N_8201,N_7798);
and U8833 (N_8833,N_8509,N_7998);
nor U8834 (N_8834,N_7665,N_7655);
or U8835 (N_8835,N_8659,N_7934);
or U8836 (N_8836,N_8483,N_8400);
nor U8837 (N_8837,N_8251,N_7732);
nor U8838 (N_8838,N_8651,N_8664);
and U8839 (N_8839,N_8114,N_8677);
xnor U8840 (N_8840,N_8293,N_7982);
or U8841 (N_8841,N_8358,N_8190);
nor U8842 (N_8842,N_7685,N_7566);
xnor U8843 (N_8843,N_8505,N_7872);
xor U8844 (N_8844,N_8089,N_8151);
nor U8845 (N_8845,N_8007,N_8101);
or U8846 (N_8846,N_7884,N_8472);
nor U8847 (N_8847,N_7906,N_7919);
and U8848 (N_8848,N_8177,N_8213);
and U8849 (N_8849,N_8629,N_8010);
nand U8850 (N_8850,N_8365,N_8490);
or U8851 (N_8851,N_7605,N_7727);
xnor U8852 (N_8852,N_8520,N_7690);
xnor U8853 (N_8853,N_8262,N_8267);
nand U8854 (N_8854,N_8305,N_7531);
and U8855 (N_8855,N_8579,N_8713);
nand U8856 (N_8856,N_7792,N_7763);
or U8857 (N_8857,N_7905,N_8253);
nor U8858 (N_8858,N_7777,N_8325);
xor U8859 (N_8859,N_8567,N_7888);
and U8860 (N_8860,N_7921,N_8434);
nand U8861 (N_8861,N_8200,N_8743);
xor U8862 (N_8862,N_8383,N_8650);
nor U8863 (N_8863,N_8009,N_7858);
and U8864 (N_8864,N_7667,N_8716);
and U8865 (N_8865,N_7673,N_7656);
nor U8866 (N_8866,N_7842,N_7759);
xor U8867 (N_8867,N_7599,N_8367);
and U8868 (N_8868,N_7613,N_8741);
nor U8869 (N_8869,N_7783,N_8210);
nor U8870 (N_8870,N_7534,N_8615);
nor U8871 (N_8871,N_8613,N_8197);
and U8872 (N_8872,N_7627,N_8135);
or U8873 (N_8873,N_8745,N_8202);
or U8874 (N_8874,N_7725,N_7894);
or U8875 (N_8875,N_7693,N_8227);
or U8876 (N_8876,N_8050,N_8676);
and U8877 (N_8877,N_8599,N_7623);
and U8878 (N_8878,N_8188,N_7698);
or U8879 (N_8879,N_7574,N_7867);
or U8880 (N_8880,N_8006,N_7991);
or U8881 (N_8881,N_8712,N_8102);
or U8882 (N_8882,N_8685,N_8045);
nor U8883 (N_8883,N_8015,N_7900);
nand U8884 (N_8884,N_7746,N_8056);
nor U8885 (N_8885,N_8023,N_8618);
or U8886 (N_8886,N_8260,N_8211);
xor U8887 (N_8887,N_8080,N_8628);
xor U8888 (N_8888,N_8277,N_8692);
or U8889 (N_8889,N_7766,N_8178);
nand U8890 (N_8890,N_8332,N_8610);
nand U8891 (N_8891,N_7672,N_8216);
xnor U8892 (N_8892,N_8131,N_8595);
nand U8893 (N_8893,N_8425,N_8438);
and U8894 (N_8894,N_7502,N_8081);
nor U8895 (N_8895,N_7942,N_7536);
xor U8896 (N_8896,N_7587,N_8258);
nand U8897 (N_8897,N_7735,N_8316);
nor U8898 (N_8898,N_7786,N_8150);
nor U8899 (N_8899,N_8396,N_8115);
nand U8900 (N_8900,N_8681,N_8055);
nand U8901 (N_8901,N_8274,N_8230);
xor U8902 (N_8902,N_7720,N_8662);
xor U8903 (N_8903,N_8619,N_8229);
nor U8904 (N_8904,N_7953,N_8140);
nand U8905 (N_8905,N_7887,N_8729);
and U8906 (N_8906,N_8341,N_8678);
nor U8907 (N_8907,N_8517,N_8624);
or U8908 (N_8908,N_7615,N_7908);
nor U8909 (N_8909,N_8427,N_8696);
nand U8910 (N_8910,N_7999,N_7810);
and U8911 (N_8911,N_8627,N_8565);
or U8912 (N_8912,N_7993,N_8295);
xnor U8913 (N_8913,N_8580,N_8380);
and U8914 (N_8914,N_7530,N_8239);
and U8915 (N_8915,N_7768,N_8571);
xnor U8916 (N_8916,N_8362,N_7678);
nand U8917 (N_8917,N_8466,N_7808);
xnor U8918 (N_8918,N_8715,N_8343);
or U8919 (N_8919,N_7744,N_8594);
nor U8920 (N_8920,N_7885,N_8421);
xor U8921 (N_8921,N_7979,N_8724);
nand U8922 (N_8922,N_7776,N_8695);
and U8923 (N_8923,N_8346,N_8215);
or U8924 (N_8924,N_7515,N_8209);
and U8925 (N_8925,N_7997,N_8237);
nand U8926 (N_8926,N_7686,N_8461);
xnor U8927 (N_8927,N_8138,N_7699);
and U8928 (N_8928,N_8680,N_8699);
xor U8929 (N_8929,N_7710,N_8576);
nand U8930 (N_8930,N_8444,N_8272);
xnor U8931 (N_8931,N_8090,N_8263);
nand U8932 (N_8932,N_7772,N_8235);
and U8933 (N_8933,N_8002,N_8653);
or U8934 (N_8934,N_7958,N_8726);
nand U8935 (N_8935,N_8666,N_8082);
xnor U8936 (N_8936,N_8068,N_8589);
nand U8937 (N_8937,N_8693,N_8570);
and U8938 (N_8938,N_7717,N_8537);
or U8939 (N_8939,N_7572,N_7955);
or U8940 (N_8940,N_7980,N_8175);
nand U8941 (N_8941,N_7961,N_8176);
nand U8942 (N_8942,N_7950,N_7702);
xor U8943 (N_8943,N_7898,N_8526);
or U8944 (N_8944,N_8249,N_8017);
xnor U8945 (N_8945,N_7848,N_8551);
or U8946 (N_8946,N_7806,N_8364);
and U8947 (N_8947,N_8491,N_8220);
nor U8948 (N_8948,N_7600,N_7718);
nand U8949 (N_8949,N_8746,N_8448);
xnor U8950 (N_8950,N_7839,N_7595);
and U8951 (N_8951,N_8463,N_8000);
xor U8952 (N_8952,N_8285,N_8283);
nor U8953 (N_8953,N_8304,N_8563);
nor U8954 (N_8954,N_7542,N_7880);
or U8955 (N_8955,N_7541,N_8475);
and U8956 (N_8956,N_8673,N_8402);
nand U8957 (N_8957,N_8372,N_7948);
xor U8958 (N_8958,N_7941,N_8652);
nor U8959 (N_8959,N_7936,N_7903);
nor U8960 (N_8960,N_8334,N_8607);
or U8961 (N_8961,N_8538,N_7923);
nand U8962 (N_8962,N_8587,N_7931);
xor U8963 (N_8963,N_8377,N_8725);
or U8964 (N_8964,N_8073,N_7715);
nor U8965 (N_8965,N_8091,N_7863);
nand U8966 (N_8966,N_7701,N_8585);
and U8967 (N_8967,N_8162,N_7745);
nand U8968 (N_8968,N_8052,N_7661);
xnor U8969 (N_8969,N_8093,N_8172);
or U8970 (N_8970,N_8345,N_8241);
nor U8971 (N_8971,N_8173,N_8368);
or U8972 (N_8972,N_7859,N_8035);
xnor U8973 (N_8973,N_8495,N_7762);
and U8974 (N_8974,N_8621,N_8711);
or U8975 (N_8975,N_7992,N_8540);
or U8976 (N_8976,N_8516,N_7754);
or U8977 (N_8977,N_7657,N_7543);
or U8978 (N_8978,N_8539,N_8654);
and U8979 (N_8979,N_7524,N_8180);
and U8980 (N_8980,N_8616,N_7928);
xor U8981 (N_8981,N_8441,N_7562);
nand U8982 (N_8982,N_8271,N_8536);
nor U8983 (N_8983,N_7904,N_8067);
xnor U8984 (N_8984,N_7555,N_8468);
or U8985 (N_8985,N_7552,N_8426);
nor U8986 (N_8986,N_8488,N_8494);
nor U8987 (N_8987,N_8104,N_8480);
nor U8988 (N_8988,N_8191,N_7622);
and U8989 (N_8989,N_7610,N_8123);
xnor U8990 (N_8990,N_7585,N_7681);
and U8991 (N_8991,N_8515,N_7790);
nand U8992 (N_8992,N_7682,N_8484);
nand U8993 (N_8993,N_8694,N_8722);
nand U8994 (N_8994,N_8170,N_7851);
xor U8995 (N_8995,N_7504,N_8710);
and U8996 (N_8996,N_7789,N_8099);
and U8997 (N_8997,N_8548,N_8658);
or U8998 (N_8998,N_8256,N_7516);
xor U8999 (N_8999,N_8740,N_7509);
and U9000 (N_9000,N_7779,N_8530);
nor U9001 (N_9001,N_7816,N_8057);
and U9002 (N_9002,N_8510,N_7617);
nor U9003 (N_9003,N_8485,N_8219);
xor U9004 (N_9004,N_8038,N_8085);
or U9005 (N_9005,N_8299,N_7771);
nand U9006 (N_9006,N_7932,N_7774);
or U9007 (N_9007,N_8074,N_7817);
or U9008 (N_9008,N_8129,N_7539);
nand U9009 (N_9009,N_8184,N_7797);
nor U9010 (N_9010,N_8111,N_8354);
nor U9011 (N_9011,N_8455,N_8004);
and U9012 (N_9012,N_8408,N_8054);
or U9013 (N_9013,N_7695,N_8029);
or U9014 (N_9014,N_8612,N_8070);
or U9015 (N_9015,N_8700,N_7820);
and U9016 (N_9016,N_8244,N_7604);
or U9017 (N_9017,N_8250,N_8043);
nor U9018 (N_9018,N_8697,N_7831);
nand U9019 (N_9019,N_8561,N_8376);
and U9020 (N_9020,N_8012,N_8493);
xnor U9021 (N_9021,N_8502,N_8339);
or U9022 (N_9022,N_8022,N_8656);
xor U9023 (N_9023,N_8242,N_8183);
and U9024 (N_9024,N_8721,N_7582);
xnor U9025 (N_9025,N_8717,N_8665);
and U9026 (N_9026,N_8347,N_7822);
xnor U9027 (N_9027,N_7973,N_8519);
nand U9028 (N_9028,N_8406,N_8139);
and U9029 (N_9029,N_7684,N_7590);
or U9030 (N_9030,N_8185,N_8727);
nor U9031 (N_9031,N_7828,N_8326);
or U9032 (N_9032,N_8590,N_7739);
or U9033 (N_9033,N_8330,N_7588);
or U9034 (N_9034,N_8546,N_8452);
xor U9035 (N_9035,N_8103,N_8223);
and U9036 (N_9036,N_8748,N_7501);
xnor U9037 (N_9037,N_7952,N_8684);
xor U9038 (N_9038,N_8532,N_8428);
or U9039 (N_9039,N_7824,N_7576);
xor U9040 (N_9040,N_7891,N_8401);
and U9041 (N_9041,N_7659,N_8269);
nand U9042 (N_9042,N_8147,N_7624);
nor U9043 (N_9043,N_8668,N_8087);
and U9044 (N_9044,N_8142,N_8447);
nand U9045 (N_9045,N_7749,N_7528);
xor U9046 (N_9046,N_7563,N_8307);
or U9047 (N_9047,N_8550,N_8155);
and U9048 (N_9048,N_8403,N_8031);
nor U9049 (N_9049,N_7883,N_8672);
and U9050 (N_9050,N_7675,N_8337);
nor U9051 (N_9051,N_8478,N_8507);
nor U9052 (N_9052,N_8557,N_7634);
and U9053 (N_9053,N_8222,N_8643);
or U9054 (N_9054,N_8707,N_7983);
xnor U9055 (N_9055,N_8243,N_8270);
and U9056 (N_9056,N_8107,N_8355);
xnor U9057 (N_9057,N_7546,N_8518);
xor U9058 (N_9058,N_7943,N_7737);
nor U9059 (N_9059,N_8547,N_7957);
and U9060 (N_9060,N_7733,N_8634);
xor U9061 (N_9061,N_7742,N_8701);
xnor U9062 (N_9062,N_7954,N_8351);
nor U9063 (N_9063,N_8436,N_8691);
xor U9064 (N_9064,N_8025,N_7743);
nor U9065 (N_9065,N_8094,N_8259);
and U9066 (N_9066,N_8597,N_7811);
or U9067 (N_9067,N_8011,N_8153);
or U9068 (N_9068,N_7795,N_8075);
nand U9069 (N_9069,N_7975,N_8657);
nand U9070 (N_9070,N_7529,N_8578);
nand U9071 (N_9071,N_8527,N_8553);
and U9072 (N_9072,N_8498,N_8288);
xnor U9073 (N_9073,N_7532,N_7879);
nor U9074 (N_9074,N_7775,N_7800);
xnor U9075 (N_9075,N_7548,N_7554);
xnor U9076 (N_9076,N_8460,N_8280);
xor U9077 (N_9077,N_7823,N_7965);
and U9078 (N_9078,N_8001,N_8186);
xnor U9079 (N_9079,N_7713,N_8110);
xor U9080 (N_9080,N_8117,N_8287);
or U9081 (N_9081,N_7791,N_7629);
xnor U9082 (N_9082,N_8027,N_7860);
and U9083 (N_9083,N_7758,N_7938);
nor U9084 (N_9084,N_8489,N_7632);
and U9085 (N_9085,N_8649,N_8601);
xnor U9086 (N_9086,N_8419,N_8036);
and U9087 (N_9087,N_8116,N_7614);
nor U9088 (N_9088,N_8508,N_7812);
xnor U9089 (N_9089,N_8112,N_7918);
xor U9090 (N_9090,N_7939,N_7986);
nor U9091 (N_9091,N_8042,N_7878);
nand U9092 (N_9092,N_8541,N_7586);
and U9093 (N_9093,N_7910,N_8008);
xnor U9094 (N_9094,N_8095,N_8562);
and U9095 (N_9095,N_7988,N_8203);
xor U9096 (N_9096,N_8106,N_8399);
or U9097 (N_9097,N_7508,N_7577);
or U9098 (N_9098,N_7925,N_7607);
xnor U9099 (N_9099,N_8583,N_7521);
and U9100 (N_9100,N_8321,N_7920);
or U9101 (N_9101,N_7756,N_8449);
nand U9102 (N_9102,N_7628,N_8706);
and U9103 (N_9103,N_8181,N_8476);
nand U9104 (N_9104,N_8723,N_7929);
nor U9105 (N_9105,N_8273,N_7547);
nor U9106 (N_9106,N_8331,N_7729);
xor U9107 (N_9107,N_7784,N_7706);
nand U9108 (N_9108,N_7892,N_8395);
nor U9109 (N_9109,N_8072,N_7639);
or U9110 (N_9110,N_8039,N_8047);
and U9111 (N_9111,N_8282,N_7597);
xnor U9112 (N_9112,N_7609,N_7778);
xnor U9113 (N_9113,N_8063,N_8335);
or U9114 (N_9114,N_8734,N_8430);
and U9115 (N_9115,N_7581,N_7649);
nand U9116 (N_9116,N_7598,N_8432);
xnor U9117 (N_9117,N_8360,N_7734);
nand U9118 (N_9118,N_8603,N_7909);
or U9119 (N_9119,N_8257,N_7654);
nand U9120 (N_9120,N_7567,N_7716);
and U9121 (N_9121,N_7881,N_8459);
nor U9122 (N_9122,N_7707,N_8324);
nor U9123 (N_9123,N_8098,N_8513);
or U9124 (N_9124,N_7575,N_8608);
nand U9125 (N_9125,N_8559,N_8386);
xor U9126 (N_9126,N_8148,N_7704);
and U9127 (N_9127,N_8301,N_8083);
xor U9128 (N_9128,N_8423,N_8187);
and U9129 (N_9129,N_8166,N_8266);
nor U9130 (N_9130,N_8604,N_8118);
nand U9131 (N_9131,N_7840,N_7945);
nor U9132 (N_9132,N_8378,N_7663);
or U9133 (N_9133,N_8416,N_7606);
nor U9134 (N_9134,N_7630,N_7794);
and U9135 (N_9135,N_7726,N_7922);
xor U9136 (N_9136,N_8234,N_8647);
xnor U9137 (N_9137,N_8446,N_8265);
nand U9138 (N_9138,N_7592,N_8030);
nand U9139 (N_9139,N_8728,N_7959);
or U9140 (N_9140,N_8644,N_7631);
or U9141 (N_9141,N_7512,N_8623);
xor U9142 (N_9142,N_8645,N_8544);
nor U9143 (N_9143,N_8160,N_8207);
or U9144 (N_9144,N_7551,N_7506);
nor U9145 (N_9145,N_7689,N_8302);
nand U9146 (N_9146,N_8633,N_8069);
nor U9147 (N_9147,N_8132,N_8096);
nand U9148 (N_9148,N_7694,N_8445);
or U9149 (N_9149,N_8394,N_8584);
nand U9150 (N_9150,N_8313,N_7917);
and U9151 (N_9151,N_7666,N_8382);
nand U9152 (N_9152,N_8312,N_8731);
xnor U9153 (N_9153,N_8670,N_8390);
xor U9154 (N_9154,N_8504,N_8245);
and U9155 (N_9155,N_8214,N_7565);
nor U9156 (N_9156,N_7679,N_8357);
nand U9157 (N_9157,N_7890,N_7912);
nor U9158 (N_9158,N_8314,N_8698);
nor U9159 (N_9159,N_8322,N_8246);
and U9160 (N_9160,N_7976,N_7815);
xnor U9161 (N_9161,N_8286,N_8393);
or U9162 (N_9162,N_8046,N_8600);
xnor U9163 (N_9163,N_7573,N_7829);
xnor U9164 (N_9164,N_7833,N_8232);
xnor U9165 (N_9165,N_8108,N_8412);
nor U9166 (N_9166,N_7787,N_7561);
or U9167 (N_9167,N_7946,N_8709);
xor U9168 (N_9168,N_8614,N_7966);
or U9169 (N_9169,N_7844,N_7852);
nand U9170 (N_9170,N_8514,N_8338);
and U9171 (N_9171,N_8268,N_8136);
nor U9172 (N_9172,N_7559,N_8577);
xor U9173 (N_9173,N_7564,N_8336);
xnor U9174 (N_9174,N_7751,N_8189);
or U9175 (N_9175,N_7821,N_8611);
nor U9176 (N_9176,N_7949,N_8450);
and U9177 (N_9177,N_7937,N_8159);
or U9178 (N_9178,N_8617,N_7793);
nand U9179 (N_9179,N_7594,N_7895);
nor U9180 (N_9180,N_7871,N_7956);
nand U9181 (N_9181,N_8344,N_7533);
or U9182 (N_9182,N_7611,N_7832);
or U9183 (N_9183,N_8024,N_7962);
xnor U9184 (N_9184,N_8409,N_8487);
nor U9185 (N_9185,N_8352,N_8405);
nand U9186 (N_9186,N_7651,N_8703);
nor U9187 (N_9187,N_8356,N_8066);
and U9188 (N_9188,N_8240,N_8646);
nand U9189 (N_9189,N_7981,N_8199);
xor U9190 (N_9190,N_7676,N_8733);
or U9191 (N_9191,N_8424,N_8238);
or U9192 (N_9192,N_8431,N_8048);
xnor U9193 (N_9193,N_7984,N_7721);
xor U9194 (N_9194,N_8555,N_7834);
nand U9195 (N_9195,N_8467,N_8414);
xnor U9196 (N_9196,N_8586,N_8679);
or U9197 (N_9197,N_8264,N_8500);
nor U9198 (N_9198,N_7558,N_8317);
xor U9199 (N_9199,N_8625,N_8560);
or U9200 (N_9200,N_8182,N_7540);
or U9201 (N_9201,N_8143,N_8044);
nor U9202 (N_9202,N_7596,N_8146);
nand U9203 (N_9203,N_8077,N_7711);
and U9204 (N_9204,N_7964,N_8040);
or U9205 (N_9205,N_8392,N_8113);
and U9206 (N_9206,N_7841,N_8196);
and U9207 (N_9207,N_8648,N_8439);
and U9208 (N_9208,N_7671,N_8718);
and U9209 (N_9209,N_7714,N_8327);
nor U9210 (N_9210,N_8667,N_8126);
xor U9211 (N_9211,N_8477,N_8473);
or U9212 (N_9212,N_8535,N_8499);
xnor U9213 (N_9213,N_7513,N_8366);
xor U9214 (N_9214,N_7978,N_8252);
nand U9215 (N_9215,N_8254,N_7697);
and U9216 (N_9216,N_8034,N_8521);
or U9217 (N_9217,N_8542,N_8097);
nand U9218 (N_9218,N_7520,N_8492);
or U9219 (N_9219,N_7802,N_8417);
xor U9220 (N_9220,N_7511,N_7722);
or U9221 (N_9221,N_8569,N_7911);
xnor U9222 (N_9222,N_7724,N_8635);
xor U9223 (N_9223,N_8622,N_7537);
or U9224 (N_9224,N_8564,N_8379);
or U9225 (N_9225,N_8742,N_8418);
or U9226 (N_9226,N_8217,N_8353);
xnor U9227 (N_9227,N_8152,N_7854);
nand U9228 (N_9228,N_7645,N_8738);
and U9229 (N_9229,N_7640,N_8720);
xor U9230 (N_9230,N_8410,N_7799);
xnor U9231 (N_9231,N_8315,N_7527);
nand U9232 (N_9232,N_8134,N_8065);
xor U9233 (N_9233,N_7845,N_8574);
and U9234 (N_9234,N_7926,N_8059);
or U9235 (N_9235,N_7882,N_7579);
nand U9236 (N_9236,N_8749,N_8522);
or U9237 (N_9237,N_8323,N_8486);
nand U9238 (N_9238,N_8373,N_7505);
nand U9239 (N_9239,N_8236,N_8437);
and U9240 (N_9240,N_7658,N_8133);
or U9241 (N_9241,N_8735,N_7990);
xnor U9242 (N_9242,N_8702,N_7519);
nor U9243 (N_9243,N_8413,N_7730);
or U9244 (N_9244,N_8596,N_7788);
or U9245 (N_9245,N_7868,N_8119);
and U9246 (N_9246,N_8233,N_8591);
nor U9247 (N_9247,N_7897,N_8598);
and U9248 (N_9248,N_7994,N_8310);
nand U9249 (N_9249,N_8429,N_8479);
xor U9250 (N_9250,N_7752,N_7662);
xnor U9251 (N_9251,N_8686,N_8032);
nor U9252 (N_9252,N_7857,N_8533);
or U9253 (N_9253,N_7843,N_8736);
xnor U9254 (N_9254,N_7862,N_7647);
nor U9255 (N_9255,N_8435,N_8350);
nand U9256 (N_9256,N_7677,N_8088);
xnor U9257 (N_9257,N_8407,N_8014);
nor U9258 (N_9258,N_8558,N_7773);
nand U9259 (N_9259,N_8397,N_7782);
or U9260 (N_9260,N_8198,N_8609);
or U9261 (N_9261,N_8289,N_8566);
xor U9262 (N_9262,N_7861,N_8525);
nor U9263 (N_9263,N_7750,N_7865);
and U9264 (N_9264,N_7916,N_8154);
nor U9265 (N_9265,N_7760,N_7522);
nand U9266 (N_9266,N_8297,N_8058);
nor U9267 (N_9267,N_7648,N_7741);
or U9268 (N_9268,N_8605,N_8704);
or U9269 (N_9269,N_8506,N_8018);
xor U9270 (N_9270,N_7819,N_8454);
nand U9271 (N_9271,N_7510,N_7738);
nor U9272 (N_9272,N_8549,N_8422);
nand U9273 (N_9273,N_7641,N_8545);
or U9274 (N_9274,N_7601,N_7761);
xnor U9275 (N_9275,N_8349,N_8309);
xor U9276 (N_9276,N_8300,N_7644);
nand U9277 (N_9277,N_7944,N_8528);
nor U9278 (N_9278,N_8404,N_7825);
or U9279 (N_9279,N_7642,N_8501);
or U9280 (N_9280,N_7866,N_7830);
and U9281 (N_9281,N_8638,N_8661);
nand U9282 (N_9282,N_7549,N_7764);
xor U9283 (N_9283,N_7755,N_7652);
nor U9284 (N_9284,N_8636,N_8626);
or U9285 (N_9285,N_8021,N_7847);
xnor U9286 (N_9286,N_8060,N_7593);
and U9287 (N_9287,N_8512,N_7874);
and U9288 (N_9288,N_7643,N_7691);
or U9289 (N_9289,N_8275,N_8385);
xnor U9290 (N_9290,N_8453,N_8016);
or U9291 (N_9291,N_8639,N_8375);
or U9292 (N_9292,N_7995,N_8149);
nand U9293 (N_9293,N_8171,N_8019);
nor U9294 (N_9294,N_8524,N_8276);
xor U9295 (N_9295,N_7809,N_8329);
nand U9296 (N_9296,N_8292,N_8028);
or U9297 (N_9297,N_7855,N_7683);
nor U9298 (N_9298,N_7780,N_7688);
or U9299 (N_9299,N_8165,N_8732);
nor U9300 (N_9300,N_8218,N_7748);
or U9301 (N_9301,N_8226,N_7769);
nand U9302 (N_9302,N_8474,N_7523);
or U9303 (N_9303,N_8398,N_8100);
nand U9304 (N_9304,N_7638,N_8127);
nor U9305 (N_9305,N_8496,N_8158);
nand U9306 (N_9306,N_7747,N_8041);
or U9307 (N_9307,N_8433,N_8572);
xor U9308 (N_9308,N_7818,N_8071);
xnor U9309 (N_9309,N_7626,N_7517);
nor U9310 (N_9310,N_8125,N_8261);
or U9311 (N_9311,N_8308,N_7886);
nor U9312 (N_9312,N_8457,N_7987);
xor U9313 (N_9313,N_7571,N_8359);
nor U9314 (N_9314,N_8369,N_7814);
and U9315 (N_9315,N_8298,N_8157);
xor U9316 (N_9316,N_8714,N_8630);
xor U9317 (N_9317,N_7569,N_7896);
xnor U9318 (N_9318,N_7584,N_8462);
xnor U9319 (N_9319,N_7803,N_8208);
and U9320 (N_9320,N_7924,N_7753);
nand U9321 (N_9321,N_7680,N_7570);
and U9322 (N_9322,N_7836,N_7796);
nor U9323 (N_9323,N_7669,N_7728);
and U9324 (N_9324,N_8464,N_7970);
nor U9325 (N_9325,N_8588,N_8415);
nand U9326 (N_9326,N_8145,N_8465);
or U9327 (N_9327,N_7687,N_7907);
or U9328 (N_9328,N_8248,N_8279);
xor U9329 (N_9329,N_8739,N_8005);
or U9330 (N_9330,N_8333,N_8195);
xnor U9331 (N_9331,N_8340,N_7535);
xor U9332 (N_9332,N_8470,N_8663);
xnor U9333 (N_9333,N_8534,N_8705);
or U9334 (N_9334,N_7635,N_8440);
nor U9335 (N_9335,N_8387,N_8320);
xor U9336 (N_9336,N_7705,N_7633);
and U9337 (N_9337,N_7985,N_7785);
or U9338 (N_9338,N_8708,N_8503);
nand U9339 (N_9339,N_8174,N_8688);
nand U9340 (N_9340,N_7580,N_7968);
or U9341 (N_9341,N_8064,N_7849);
nor U9342 (N_9342,N_8593,N_8205);
nand U9343 (N_9343,N_8371,N_7538);
xnor U9344 (N_9344,N_8164,N_8575);
xor U9345 (N_9345,N_7850,N_8669);
nor U9346 (N_9346,N_8554,N_8342);
nor U9347 (N_9347,N_7709,N_8179);
or U9348 (N_9348,N_7668,N_8294);
xor U9349 (N_9349,N_8051,N_7838);
or U9350 (N_9350,N_8053,N_7670);
xor U9351 (N_9351,N_7899,N_7703);
nor U9352 (N_9352,N_8581,N_8637);
nor U9353 (N_9353,N_7901,N_8361);
nand U9354 (N_9354,N_8049,N_7805);
nand U9355 (N_9355,N_7913,N_7972);
nand U9356 (N_9356,N_8497,N_7765);
xor U9357 (N_9357,N_7757,N_7731);
nor U9358 (N_9358,N_7770,N_7525);
nor U9359 (N_9359,N_7767,N_7619);
xor U9360 (N_9360,N_7503,N_8130);
xor U9361 (N_9361,N_8543,N_8156);
and U9362 (N_9362,N_8529,N_8374);
and U9363 (N_9363,N_8278,N_8120);
nand U9364 (N_9364,N_8079,N_7556);
xor U9365 (N_9365,N_8552,N_8281);
and U9366 (N_9366,N_8319,N_7864);
xor U9367 (N_9367,N_8033,N_8655);
and U9368 (N_9368,N_7637,N_8086);
and U9369 (N_9369,N_7553,N_8128);
nor U9370 (N_9370,N_7835,N_8013);
nand U9371 (N_9371,N_8690,N_7877);
nor U9372 (N_9372,N_8420,N_7708);
and U9373 (N_9373,N_7621,N_7915);
nand U9374 (N_9374,N_7960,N_8730);
xor U9375 (N_9375,N_8066,N_7907);
or U9376 (N_9376,N_8101,N_8619);
nor U9377 (N_9377,N_8438,N_8318);
or U9378 (N_9378,N_8445,N_8147);
nand U9379 (N_9379,N_8586,N_8264);
or U9380 (N_9380,N_8269,N_7848);
or U9381 (N_9381,N_8372,N_7513);
nor U9382 (N_9382,N_7829,N_7869);
nand U9383 (N_9383,N_7921,N_8508);
xor U9384 (N_9384,N_7574,N_8286);
and U9385 (N_9385,N_7785,N_8090);
nor U9386 (N_9386,N_7564,N_7865);
or U9387 (N_9387,N_8704,N_8691);
nand U9388 (N_9388,N_8561,N_8672);
nand U9389 (N_9389,N_8326,N_8524);
xor U9390 (N_9390,N_7770,N_8617);
and U9391 (N_9391,N_7901,N_8695);
xnor U9392 (N_9392,N_7941,N_8302);
and U9393 (N_9393,N_8367,N_8717);
xor U9394 (N_9394,N_8731,N_8443);
xor U9395 (N_9395,N_8682,N_8731);
or U9396 (N_9396,N_7522,N_8595);
nand U9397 (N_9397,N_8533,N_7655);
or U9398 (N_9398,N_7882,N_8647);
nor U9399 (N_9399,N_7703,N_8273);
xnor U9400 (N_9400,N_8600,N_8240);
nor U9401 (N_9401,N_8512,N_8245);
and U9402 (N_9402,N_7552,N_8358);
or U9403 (N_9403,N_8326,N_8414);
and U9404 (N_9404,N_8375,N_8016);
or U9405 (N_9405,N_8645,N_7608);
xnor U9406 (N_9406,N_8545,N_7612);
nand U9407 (N_9407,N_8430,N_8149);
xnor U9408 (N_9408,N_8621,N_7566);
nand U9409 (N_9409,N_7777,N_8515);
nor U9410 (N_9410,N_8421,N_8364);
nand U9411 (N_9411,N_8698,N_8700);
nand U9412 (N_9412,N_8323,N_8707);
nand U9413 (N_9413,N_7505,N_8111);
or U9414 (N_9414,N_7983,N_7755);
or U9415 (N_9415,N_8385,N_7730);
xnor U9416 (N_9416,N_8401,N_8491);
and U9417 (N_9417,N_7755,N_8547);
xor U9418 (N_9418,N_8287,N_8014);
or U9419 (N_9419,N_7592,N_8213);
xnor U9420 (N_9420,N_8296,N_8324);
and U9421 (N_9421,N_7825,N_7729);
and U9422 (N_9422,N_8683,N_7937);
nor U9423 (N_9423,N_7981,N_8107);
or U9424 (N_9424,N_8668,N_7975);
nand U9425 (N_9425,N_7925,N_8245);
nor U9426 (N_9426,N_8427,N_7679);
nor U9427 (N_9427,N_7705,N_8540);
and U9428 (N_9428,N_8430,N_7519);
and U9429 (N_9429,N_8288,N_8236);
or U9430 (N_9430,N_8084,N_7833);
nand U9431 (N_9431,N_7966,N_8136);
nand U9432 (N_9432,N_8473,N_7943);
and U9433 (N_9433,N_7655,N_8045);
or U9434 (N_9434,N_8726,N_7880);
nand U9435 (N_9435,N_8725,N_8164);
nand U9436 (N_9436,N_8504,N_7601);
xnor U9437 (N_9437,N_8235,N_7591);
nor U9438 (N_9438,N_7714,N_8302);
nor U9439 (N_9439,N_8482,N_7587);
xor U9440 (N_9440,N_8727,N_8028);
xnor U9441 (N_9441,N_8550,N_8129);
xor U9442 (N_9442,N_8299,N_8723);
xor U9443 (N_9443,N_7565,N_8220);
nand U9444 (N_9444,N_8728,N_8416);
nor U9445 (N_9445,N_8626,N_8099);
nor U9446 (N_9446,N_8099,N_7812);
nor U9447 (N_9447,N_7904,N_8617);
and U9448 (N_9448,N_7863,N_8534);
nor U9449 (N_9449,N_8279,N_7679);
nor U9450 (N_9450,N_7801,N_8345);
and U9451 (N_9451,N_8682,N_8124);
xor U9452 (N_9452,N_7862,N_8301);
xnor U9453 (N_9453,N_7755,N_8434);
nor U9454 (N_9454,N_7982,N_7837);
xnor U9455 (N_9455,N_8348,N_8603);
xor U9456 (N_9456,N_8432,N_8445);
nor U9457 (N_9457,N_8372,N_8537);
nor U9458 (N_9458,N_8555,N_8332);
and U9459 (N_9459,N_8524,N_7885);
nor U9460 (N_9460,N_8490,N_8742);
and U9461 (N_9461,N_8197,N_7553);
or U9462 (N_9462,N_8489,N_8529);
or U9463 (N_9463,N_8212,N_8049);
nor U9464 (N_9464,N_8563,N_8065);
nor U9465 (N_9465,N_8444,N_8343);
nor U9466 (N_9466,N_7549,N_7617);
or U9467 (N_9467,N_8292,N_7644);
nor U9468 (N_9468,N_8098,N_7709);
nor U9469 (N_9469,N_8678,N_8725);
or U9470 (N_9470,N_8104,N_8232);
and U9471 (N_9471,N_8447,N_8450);
xor U9472 (N_9472,N_8034,N_8299);
nor U9473 (N_9473,N_8128,N_8739);
nor U9474 (N_9474,N_8577,N_8417);
or U9475 (N_9475,N_7879,N_8113);
xor U9476 (N_9476,N_8367,N_7697);
or U9477 (N_9477,N_8144,N_8354);
xor U9478 (N_9478,N_8455,N_8507);
nor U9479 (N_9479,N_8459,N_7823);
nand U9480 (N_9480,N_8465,N_8300);
and U9481 (N_9481,N_8243,N_8199);
xnor U9482 (N_9482,N_8549,N_7932);
nor U9483 (N_9483,N_8363,N_8336);
nand U9484 (N_9484,N_8697,N_8236);
nor U9485 (N_9485,N_8566,N_8689);
xnor U9486 (N_9486,N_8450,N_7913);
or U9487 (N_9487,N_8106,N_8498);
nand U9488 (N_9488,N_8185,N_7583);
nand U9489 (N_9489,N_8107,N_7559);
nor U9490 (N_9490,N_8174,N_7539);
or U9491 (N_9491,N_7961,N_8322);
nor U9492 (N_9492,N_8364,N_7771);
xnor U9493 (N_9493,N_7981,N_8304);
or U9494 (N_9494,N_7501,N_7754);
nand U9495 (N_9495,N_8056,N_8730);
or U9496 (N_9496,N_8733,N_7716);
or U9497 (N_9497,N_8591,N_8373);
or U9498 (N_9498,N_8565,N_7819);
or U9499 (N_9499,N_8093,N_7553);
or U9500 (N_9500,N_8650,N_8272);
and U9501 (N_9501,N_7835,N_8380);
nor U9502 (N_9502,N_8007,N_8004);
nand U9503 (N_9503,N_8001,N_8704);
xor U9504 (N_9504,N_8233,N_7714);
xnor U9505 (N_9505,N_8635,N_7747);
and U9506 (N_9506,N_8672,N_7523);
or U9507 (N_9507,N_8079,N_7867);
or U9508 (N_9508,N_8490,N_8272);
and U9509 (N_9509,N_8543,N_7533);
xnor U9510 (N_9510,N_7576,N_8665);
nor U9511 (N_9511,N_8451,N_7791);
or U9512 (N_9512,N_8387,N_8280);
nor U9513 (N_9513,N_8385,N_8261);
xnor U9514 (N_9514,N_8285,N_8231);
and U9515 (N_9515,N_7695,N_7765);
nor U9516 (N_9516,N_8172,N_7708);
xnor U9517 (N_9517,N_8384,N_7598);
or U9518 (N_9518,N_8520,N_8357);
or U9519 (N_9519,N_8374,N_8144);
or U9520 (N_9520,N_8708,N_8474);
nor U9521 (N_9521,N_8597,N_7914);
nor U9522 (N_9522,N_8359,N_8072);
or U9523 (N_9523,N_7999,N_8545);
xor U9524 (N_9524,N_8290,N_7549);
nand U9525 (N_9525,N_8384,N_8208);
nor U9526 (N_9526,N_8047,N_8037);
nand U9527 (N_9527,N_7795,N_8293);
or U9528 (N_9528,N_7865,N_7951);
or U9529 (N_9529,N_8613,N_8693);
or U9530 (N_9530,N_8250,N_8141);
nor U9531 (N_9531,N_8095,N_8404);
nand U9532 (N_9532,N_7638,N_8154);
xnor U9533 (N_9533,N_8201,N_8295);
or U9534 (N_9534,N_8282,N_8194);
or U9535 (N_9535,N_8313,N_8065);
or U9536 (N_9536,N_8143,N_8553);
xor U9537 (N_9537,N_8045,N_8645);
and U9538 (N_9538,N_8045,N_8743);
and U9539 (N_9539,N_7949,N_8175);
and U9540 (N_9540,N_7877,N_7809);
nand U9541 (N_9541,N_8250,N_8210);
and U9542 (N_9542,N_7900,N_7545);
or U9543 (N_9543,N_7521,N_8354);
or U9544 (N_9544,N_7903,N_7802);
or U9545 (N_9545,N_8372,N_8188);
or U9546 (N_9546,N_7866,N_8364);
or U9547 (N_9547,N_8601,N_7740);
nand U9548 (N_9548,N_8023,N_7671);
and U9549 (N_9549,N_8347,N_7676);
xor U9550 (N_9550,N_7804,N_8310);
or U9551 (N_9551,N_8407,N_7856);
nand U9552 (N_9552,N_7756,N_8331);
nand U9553 (N_9553,N_8616,N_7671);
nor U9554 (N_9554,N_7649,N_8454);
and U9555 (N_9555,N_8236,N_7630);
nand U9556 (N_9556,N_8519,N_8253);
nor U9557 (N_9557,N_8749,N_8031);
nor U9558 (N_9558,N_8455,N_8203);
nand U9559 (N_9559,N_7643,N_8045);
nor U9560 (N_9560,N_7782,N_7655);
or U9561 (N_9561,N_8745,N_8588);
nor U9562 (N_9562,N_7989,N_8706);
nand U9563 (N_9563,N_7923,N_8090);
nand U9564 (N_9564,N_8429,N_7839);
nor U9565 (N_9565,N_8551,N_7717);
and U9566 (N_9566,N_7781,N_7719);
or U9567 (N_9567,N_8581,N_8159);
nor U9568 (N_9568,N_8350,N_8377);
xnor U9569 (N_9569,N_7946,N_8453);
xnor U9570 (N_9570,N_8306,N_7967);
nor U9571 (N_9571,N_7758,N_8424);
or U9572 (N_9572,N_8159,N_7893);
nor U9573 (N_9573,N_8054,N_8150);
xnor U9574 (N_9574,N_8587,N_8495);
and U9575 (N_9575,N_8616,N_8037);
or U9576 (N_9576,N_8416,N_7696);
or U9577 (N_9577,N_7763,N_7942);
and U9578 (N_9578,N_8070,N_8401);
and U9579 (N_9579,N_7549,N_8357);
and U9580 (N_9580,N_8591,N_8158);
nand U9581 (N_9581,N_8344,N_8451);
or U9582 (N_9582,N_8705,N_7945);
or U9583 (N_9583,N_8060,N_7644);
and U9584 (N_9584,N_7754,N_7667);
xor U9585 (N_9585,N_8338,N_8449);
and U9586 (N_9586,N_7873,N_7907);
nor U9587 (N_9587,N_7600,N_7570);
and U9588 (N_9588,N_8343,N_8313);
and U9589 (N_9589,N_7544,N_7629);
or U9590 (N_9590,N_7967,N_7549);
or U9591 (N_9591,N_7810,N_8316);
nor U9592 (N_9592,N_8026,N_8721);
nand U9593 (N_9593,N_8519,N_7802);
nor U9594 (N_9594,N_7585,N_8335);
or U9595 (N_9595,N_7739,N_7652);
or U9596 (N_9596,N_7903,N_8427);
or U9597 (N_9597,N_8501,N_8496);
xor U9598 (N_9598,N_7668,N_7724);
and U9599 (N_9599,N_7865,N_8521);
and U9600 (N_9600,N_8727,N_8174);
nand U9601 (N_9601,N_8251,N_8384);
or U9602 (N_9602,N_8533,N_8440);
or U9603 (N_9603,N_7984,N_8113);
nand U9604 (N_9604,N_8573,N_7856);
and U9605 (N_9605,N_7615,N_8596);
xnor U9606 (N_9606,N_8720,N_8595);
or U9607 (N_9607,N_8043,N_7774);
and U9608 (N_9608,N_7515,N_8253);
and U9609 (N_9609,N_8691,N_7747);
nor U9610 (N_9610,N_8355,N_7647);
xnor U9611 (N_9611,N_8226,N_8670);
xor U9612 (N_9612,N_7807,N_7729);
xor U9613 (N_9613,N_8024,N_7744);
or U9614 (N_9614,N_8447,N_8059);
xor U9615 (N_9615,N_7757,N_8158);
xor U9616 (N_9616,N_8557,N_8737);
nand U9617 (N_9617,N_7820,N_8675);
or U9618 (N_9618,N_7513,N_7523);
and U9619 (N_9619,N_8725,N_8378);
nand U9620 (N_9620,N_8396,N_8435);
or U9621 (N_9621,N_8472,N_8432);
xnor U9622 (N_9622,N_7587,N_8597);
nand U9623 (N_9623,N_8255,N_8171);
xor U9624 (N_9624,N_8694,N_8283);
nand U9625 (N_9625,N_8719,N_8351);
nor U9626 (N_9626,N_8162,N_8021);
nand U9627 (N_9627,N_8624,N_7527);
nor U9628 (N_9628,N_8023,N_8521);
nand U9629 (N_9629,N_8504,N_8725);
and U9630 (N_9630,N_7816,N_7880);
xor U9631 (N_9631,N_8420,N_7931);
xnor U9632 (N_9632,N_8534,N_8202);
xor U9633 (N_9633,N_7975,N_7887);
nand U9634 (N_9634,N_8718,N_7836);
xor U9635 (N_9635,N_8476,N_7624);
nor U9636 (N_9636,N_8552,N_7574);
and U9637 (N_9637,N_8419,N_8564);
and U9638 (N_9638,N_8427,N_8562);
xor U9639 (N_9639,N_8585,N_8540);
nor U9640 (N_9640,N_8049,N_8675);
or U9641 (N_9641,N_7743,N_8545);
nand U9642 (N_9642,N_8017,N_8737);
nand U9643 (N_9643,N_8614,N_7515);
xnor U9644 (N_9644,N_7923,N_8474);
nor U9645 (N_9645,N_7889,N_7818);
or U9646 (N_9646,N_7888,N_7761);
nand U9647 (N_9647,N_7802,N_8744);
xor U9648 (N_9648,N_8038,N_8417);
xnor U9649 (N_9649,N_8633,N_7858);
nor U9650 (N_9650,N_8013,N_8483);
nor U9651 (N_9651,N_7585,N_8064);
and U9652 (N_9652,N_8498,N_8298);
and U9653 (N_9653,N_8651,N_8064);
nand U9654 (N_9654,N_7770,N_7592);
xnor U9655 (N_9655,N_8073,N_7576);
nand U9656 (N_9656,N_8259,N_8511);
or U9657 (N_9657,N_8334,N_7723);
xnor U9658 (N_9658,N_8662,N_7834);
or U9659 (N_9659,N_7819,N_8312);
nor U9660 (N_9660,N_7665,N_8575);
and U9661 (N_9661,N_7699,N_7850);
nand U9662 (N_9662,N_7604,N_7833);
nand U9663 (N_9663,N_7648,N_7515);
xnor U9664 (N_9664,N_7940,N_7669);
and U9665 (N_9665,N_8424,N_8151);
and U9666 (N_9666,N_8045,N_7616);
xor U9667 (N_9667,N_8013,N_8711);
nor U9668 (N_9668,N_7666,N_7661);
nor U9669 (N_9669,N_7807,N_8621);
and U9670 (N_9670,N_7552,N_8341);
xnor U9671 (N_9671,N_8384,N_8371);
and U9672 (N_9672,N_8530,N_7989);
or U9673 (N_9673,N_8599,N_7807);
or U9674 (N_9674,N_8233,N_8526);
or U9675 (N_9675,N_7600,N_8563);
or U9676 (N_9676,N_7699,N_8526);
xnor U9677 (N_9677,N_8443,N_8092);
nand U9678 (N_9678,N_8073,N_8723);
or U9679 (N_9679,N_8616,N_8440);
nand U9680 (N_9680,N_8697,N_8259);
and U9681 (N_9681,N_8693,N_8705);
nand U9682 (N_9682,N_8205,N_8333);
or U9683 (N_9683,N_8277,N_8391);
xor U9684 (N_9684,N_8733,N_7868);
nor U9685 (N_9685,N_8661,N_8645);
xor U9686 (N_9686,N_8155,N_8421);
nor U9687 (N_9687,N_7775,N_7958);
nor U9688 (N_9688,N_7874,N_8019);
xnor U9689 (N_9689,N_7895,N_8017);
nor U9690 (N_9690,N_7765,N_7912);
nand U9691 (N_9691,N_8557,N_8337);
nor U9692 (N_9692,N_8698,N_7845);
nor U9693 (N_9693,N_8576,N_8219);
nand U9694 (N_9694,N_8638,N_8378);
xor U9695 (N_9695,N_8404,N_8042);
or U9696 (N_9696,N_7552,N_7695);
or U9697 (N_9697,N_8103,N_8119);
nand U9698 (N_9698,N_8628,N_8508);
nor U9699 (N_9699,N_8717,N_8119);
nor U9700 (N_9700,N_8035,N_8516);
or U9701 (N_9701,N_7843,N_7618);
and U9702 (N_9702,N_7548,N_7629);
nor U9703 (N_9703,N_8197,N_7708);
xor U9704 (N_9704,N_7604,N_7948);
xnor U9705 (N_9705,N_7926,N_8314);
xnor U9706 (N_9706,N_8081,N_8719);
and U9707 (N_9707,N_7537,N_7566);
nor U9708 (N_9708,N_8051,N_8072);
xor U9709 (N_9709,N_7641,N_8482);
nand U9710 (N_9710,N_8085,N_7717);
nand U9711 (N_9711,N_8701,N_8493);
nand U9712 (N_9712,N_8549,N_7733);
or U9713 (N_9713,N_8312,N_7694);
and U9714 (N_9714,N_8476,N_8504);
and U9715 (N_9715,N_8422,N_8041);
or U9716 (N_9716,N_8208,N_8232);
nand U9717 (N_9717,N_8580,N_8480);
nor U9718 (N_9718,N_7784,N_8416);
nor U9719 (N_9719,N_8254,N_7789);
and U9720 (N_9720,N_8104,N_7669);
xnor U9721 (N_9721,N_7774,N_7841);
xor U9722 (N_9722,N_8447,N_8199);
or U9723 (N_9723,N_7615,N_8093);
and U9724 (N_9724,N_8001,N_8742);
nor U9725 (N_9725,N_7869,N_8051);
or U9726 (N_9726,N_7839,N_8096);
nor U9727 (N_9727,N_8418,N_8544);
and U9728 (N_9728,N_8664,N_7919);
nor U9729 (N_9729,N_8428,N_7629);
nand U9730 (N_9730,N_7766,N_8639);
or U9731 (N_9731,N_7761,N_8112);
nor U9732 (N_9732,N_8200,N_8466);
or U9733 (N_9733,N_7588,N_8395);
and U9734 (N_9734,N_8476,N_7516);
and U9735 (N_9735,N_7721,N_7559);
xor U9736 (N_9736,N_8351,N_7849);
nor U9737 (N_9737,N_8697,N_8057);
or U9738 (N_9738,N_8302,N_8151);
xnor U9739 (N_9739,N_8223,N_8746);
and U9740 (N_9740,N_7919,N_8733);
nor U9741 (N_9741,N_8621,N_8053);
and U9742 (N_9742,N_8023,N_8022);
or U9743 (N_9743,N_8470,N_7896);
and U9744 (N_9744,N_7944,N_7817);
and U9745 (N_9745,N_8479,N_8114);
and U9746 (N_9746,N_7959,N_8053);
or U9747 (N_9747,N_8476,N_8300);
nand U9748 (N_9748,N_8050,N_8580);
xnor U9749 (N_9749,N_8627,N_8087);
nor U9750 (N_9750,N_8376,N_7575);
nor U9751 (N_9751,N_7909,N_8706);
nor U9752 (N_9752,N_8445,N_8458);
nor U9753 (N_9753,N_8683,N_8444);
or U9754 (N_9754,N_7713,N_8216);
nand U9755 (N_9755,N_8340,N_8708);
or U9756 (N_9756,N_8360,N_7572);
nand U9757 (N_9757,N_7767,N_7510);
nand U9758 (N_9758,N_7866,N_8672);
nor U9759 (N_9759,N_7585,N_8546);
xnor U9760 (N_9760,N_8732,N_7804);
nor U9761 (N_9761,N_7560,N_8297);
or U9762 (N_9762,N_7870,N_7945);
nand U9763 (N_9763,N_8063,N_7553);
xnor U9764 (N_9764,N_7525,N_8217);
xnor U9765 (N_9765,N_8341,N_7987);
and U9766 (N_9766,N_8029,N_7557);
xnor U9767 (N_9767,N_8748,N_7956);
xor U9768 (N_9768,N_7861,N_8015);
xnor U9769 (N_9769,N_8448,N_8059);
nand U9770 (N_9770,N_8402,N_8121);
nor U9771 (N_9771,N_8325,N_7893);
or U9772 (N_9772,N_8416,N_8200);
nand U9773 (N_9773,N_7515,N_8437);
or U9774 (N_9774,N_8139,N_7868);
nor U9775 (N_9775,N_7891,N_7949);
nand U9776 (N_9776,N_8345,N_8031);
xnor U9777 (N_9777,N_7908,N_8626);
or U9778 (N_9778,N_8350,N_7920);
and U9779 (N_9779,N_8733,N_8683);
nand U9780 (N_9780,N_7969,N_7563);
xor U9781 (N_9781,N_7975,N_8364);
or U9782 (N_9782,N_7569,N_8499);
nand U9783 (N_9783,N_8354,N_8192);
nand U9784 (N_9784,N_8330,N_7975);
xnor U9785 (N_9785,N_7778,N_7505);
or U9786 (N_9786,N_7798,N_7725);
xor U9787 (N_9787,N_8000,N_8524);
and U9788 (N_9788,N_8680,N_8169);
xor U9789 (N_9789,N_8409,N_7660);
xnor U9790 (N_9790,N_8715,N_8283);
or U9791 (N_9791,N_8000,N_7939);
nand U9792 (N_9792,N_8628,N_8477);
nand U9793 (N_9793,N_8250,N_8603);
nor U9794 (N_9794,N_8394,N_7781);
or U9795 (N_9795,N_7618,N_8385);
xnor U9796 (N_9796,N_8367,N_7735);
or U9797 (N_9797,N_7769,N_7917);
or U9798 (N_9798,N_7994,N_7660);
nand U9799 (N_9799,N_8445,N_8468);
xnor U9800 (N_9800,N_8333,N_7689);
or U9801 (N_9801,N_7854,N_7844);
or U9802 (N_9802,N_8371,N_7613);
or U9803 (N_9803,N_8263,N_8692);
or U9804 (N_9804,N_8483,N_7698);
nor U9805 (N_9805,N_7583,N_7915);
nand U9806 (N_9806,N_7509,N_8241);
and U9807 (N_9807,N_8229,N_8184);
nor U9808 (N_9808,N_7811,N_7710);
nand U9809 (N_9809,N_7848,N_7619);
or U9810 (N_9810,N_8355,N_7976);
nor U9811 (N_9811,N_7589,N_7601);
nand U9812 (N_9812,N_7741,N_7588);
or U9813 (N_9813,N_7540,N_7586);
nor U9814 (N_9814,N_8164,N_8549);
nand U9815 (N_9815,N_8005,N_8167);
and U9816 (N_9816,N_8556,N_8043);
and U9817 (N_9817,N_7666,N_8446);
and U9818 (N_9818,N_8281,N_8345);
xor U9819 (N_9819,N_8411,N_8696);
or U9820 (N_9820,N_8551,N_8213);
nand U9821 (N_9821,N_7766,N_7677);
nand U9822 (N_9822,N_8306,N_8044);
nor U9823 (N_9823,N_8085,N_7589);
and U9824 (N_9824,N_8470,N_8570);
nand U9825 (N_9825,N_7562,N_7795);
nor U9826 (N_9826,N_8423,N_7621);
nand U9827 (N_9827,N_7806,N_8478);
or U9828 (N_9828,N_8121,N_7863);
nor U9829 (N_9829,N_7879,N_8727);
and U9830 (N_9830,N_8170,N_8443);
xor U9831 (N_9831,N_7997,N_7633);
nor U9832 (N_9832,N_8017,N_8234);
xor U9833 (N_9833,N_7786,N_7739);
nor U9834 (N_9834,N_7608,N_8365);
nor U9835 (N_9835,N_8226,N_8496);
nor U9836 (N_9836,N_8060,N_8603);
nand U9837 (N_9837,N_7637,N_7639);
nor U9838 (N_9838,N_8246,N_7994);
or U9839 (N_9839,N_8202,N_7653);
nand U9840 (N_9840,N_8414,N_7839);
xnor U9841 (N_9841,N_8103,N_7518);
nand U9842 (N_9842,N_7829,N_8363);
nor U9843 (N_9843,N_8028,N_7998);
xnor U9844 (N_9844,N_8660,N_8725);
or U9845 (N_9845,N_8209,N_8190);
nor U9846 (N_9846,N_8724,N_8344);
and U9847 (N_9847,N_7881,N_8075);
xor U9848 (N_9848,N_7580,N_8091);
xnor U9849 (N_9849,N_7880,N_8022);
nor U9850 (N_9850,N_8266,N_8197);
nand U9851 (N_9851,N_7777,N_8629);
xnor U9852 (N_9852,N_8360,N_7810);
nor U9853 (N_9853,N_7656,N_7530);
nand U9854 (N_9854,N_7523,N_7581);
and U9855 (N_9855,N_7650,N_7952);
nor U9856 (N_9856,N_8661,N_7783);
and U9857 (N_9857,N_7613,N_7623);
or U9858 (N_9858,N_8318,N_7972);
xor U9859 (N_9859,N_7939,N_8122);
or U9860 (N_9860,N_8494,N_8011);
xor U9861 (N_9861,N_8371,N_8742);
nor U9862 (N_9862,N_8046,N_7838);
nand U9863 (N_9863,N_8447,N_7711);
nor U9864 (N_9864,N_8693,N_8418);
nor U9865 (N_9865,N_8330,N_8456);
xor U9866 (N_9866,N_8638,N_8243);
or U9867 (N_9867,N_8150,N_8730);
and U9868 (N_9868,N_7970,N_8258);
xnor U9869 (N_9869,N_8659,N_7637);
or U9870 (N_9870,N_7735,N_8138);
or U9871 (N_9871,N_7835,N_8719);
xnor U9872 (N_9872,N_8497,N_8041);
nor U9873 (N_9873,N_7582,N_7516);
or U9874 (N_9874,N_7701,N_8139);
xor U9875 (N_9875,N_8077,N_7688);
and U9876 (N_9876,N_7803,N_8323);
and U9877 (N_9877,N_7816,N_7656);
or U9878 (N_9878,N_8519,N_7862);
and U9879 (N_9879,N_8683,N_8057);
and U9880 (N_9880,N_8511,N_8104);
nand U9881 (N_9881,N_8432,N_8423);
xnor U9882 (N_9882,N_8641,N_8395);
or U9883 (N_9883,N_7996,N_7867);
nor U9884 (N_9884,N_8672,N_8571);
or U9885 (N_9885,N_7888,N_8223);
or U9886 (N_9886,N_8275,N_8717);
nand U9887 (N_9887,N_8075,N_7956);
or U9888 (N_9888,N_8199,N_8422);
nand U9889 (N_9889,N_8089,N_7913);
xnor U9890 (N_9890,N_8671,N_8155);
or U9891 (N_9891,N_8520,N_7986);
and U9892 (N_9892,N_8351,N_8070);
or U9893 (N_9893,N_8464,N_8620);
nand U9894 (N_9894,N_8193,N_8630);
nor U9895 (N_9895,N_8527,N_8747);
and U9896 (N_9896,N_8161,N_8700);
or U9897 (N_9897,N_7765,N_8094);
and U9898 (N_9898,N_8207,N_7751);
nor U9899 (N_9899,N_7821,N_8533);
xor U9900 (N_9900,N_7934,N_7657);
or U9901 (N_9901,N_8345,N_7780);
and U9902 (N_9902,N_8028,N_8725);
and U9903 (N_9903,N_8062,N_7712);
or U9904 (N_9904,N_7664,N_7990);
nor U9905 (N_9905,N_7787,N_7936);
and U9906 (N_9906,N_8392,N_8553);
or U9907 (N_9907,N_8611,N_8093);
nor U9908 (N_9908,N_7521,N_8171);
nor U9909 (N_9909,N_7527,N_8581);
nor U9910 (N_9910,N_8112,N_7588);
and U9911 (N_9911,N_7513,N_8030);
xnor U9912 (N_9912,N_8098,N_8339);
nand U9913 (N_9913,N_8744,N_7741);
nand U9914 (N_9914,N_8369,N_7522);
nand U9915 (N_9915,N_8012,N_7762);
or U9916 (N_9916,N_8338,N_8614);
nor U9917 (N_9917,N_7673,N_8647);
xor U9918 (N_9918,N_8087,N_8548);
xor U9919 (N_9919,N_8058,N_7512);
or U9920 (N_9920,N_8342,N_8598);
xnor U9921 (N_9921,N_8636,N_7945);
and U9922 (N_9922,N_8130,N_7622);
nor U9923 (N_9923,N_8000,N_7715);
and U9924 (N_9924,N_8298,N_8441);
and U9925 (N_9925,N_7685,N_8199);
and U9926 (N_9926,N_8149,N_8199);
and U9927 (N_9927,N_8686,N_7788);
xor U9928 (N_9928,N_7564,N_8429);
and U9929 (N_9929,N_7710,N_7663);
nand U9930 (N_9930,N_7572,N_8525);
or U9931 (N_9931,N_8282,N_7607);
xnor U9932 (N_9932,N_8481,N_7974);
nor U9933 (N_9933,N_7505,N_8116);
and U9934 (N_9934,N_8390,N_8080);
xor U9935 (N_9935,N_8278,N_7866);
nor U9936 (N_9936,N_8077,N_8013);
and U9937 (N_9937,N_7655,N_7540);
and U9938 (N_9938,N_8294,N_7655);
nor U9939 (N_9939,N_7577,N_7840);
nand U9940 (N_9940,N_8700,N_8321);
nand U9941 (N_9941,N_8511,N_8717);
nand U9942 (N_9942,N_8038,N_7513);
or U9943 (N_9943,N_8142,N_8534);
xnor U9944 (N_9944,N_8571,N_8385);
nor U9945 (N_9945,N_7662,N_7961);
xnor U9946 (N_9946,N_7577,N_7986);
nand U9947 (N_9947,N_8432,N_7814);
nor U9948 (N_9948,N_8011,N_8637);
xor U9949 (N_9949,N_7521,N_8318);
nor U9950 (N_9950,N_8128,N_7582);
nand U9951 (N_9951,N_7963,N_7742);
or U9952 (N_9952,N_7954,N_7994);
or U9953 (N_9953,N_8265,N_7955);
nand U9954 (N_9954,N_7738,N_7707);
or U9955 (N_9955,N_7791,N_8664);
xnor U9956 (N_9956,N_7900,N_8217);
or U9957 (N_9957,N_7614,N_7822);
nand U9958 (N_9958,N_8031,N_8458);
xor U9959 (N_9959,N_8058,N_8069);
xor U9960 (N_9960,N_7972,N_8696);
nor U9961 (N_9961,N_7541,N_7547);
nor U9962 (N_9962,N_7707,N_8604);
xnor U9963 (N_9963,N_7898,N_8681);
xor U9964 (N_9964,N_7504,N_7507);
and U9965 (N_9965,N_8617,N_8704);
or U9966 (N_9966,N_8536,N_7667);
nand U9967 (N_9967,N_7968,N_8410);
nand U9968 (N_9968,N_8270,N_7608);
xor U9969 (N_9969,N_8046,N_8312);
xor U9970 (N_9970,N_7802,N_7672);
and U9971 (N_9971,N_7927,N_8099);
and U9972 (N_9972,N_7692,N_7839);
or U9973 (N_9973,N_8522,N_8084);
or U9974 (N_9974,N_8627,N_8444);
nand U9975 (N_9975,N_7631,N_7618);
nor U9976 (N_9976,N_8362,N_8363);
nor U9977 (N_9977,N_7880,N_7567);
xor U9978 (N_9978,N_8536,N_7871);
and U9979 (N_9979,N_8123,N_8164);
nor U9980 (N_9980,N_8189,N_8487);
nor U9981 (N_9981,N_8254,N_8242);
and U9982 (N_9982,N_7635,N_7745);
and U9983 (N_9983,N_8194,N_8039);
or U9984 (N_9984,N_7621,N_8408);
nand U9985 (N_9985,N_8571,N_7803);
xor U9986 (N_9986,N_8180,N_8498);
and U9987 (N_9987,N_7513,N_8020);
nor U9988 (N_9988,N_8319,N_8523);
nor U9989 (N_9989,N_7959,N_7853);
nand U9990 (N_9990,N_8070,N_7672);
xnor U9991 (N_9991,N_8550,N_8396);
nand U9992 (N_9992,N_8318,N_7528);
nand U9993 (N_9993,N_7612,N_8303);
xor U9994 (N_9994,N_8391,N_8215);
xnor U9995 (N_9995,N_7709,N_8269);
or U9996 (N_9996,N_8447,N_7886);
nor U9997 (N_9997,N_8089,N_8048);
nand U9998 (N_9998,N_8584,N_8351);
and U9999 (N_9999,N_8067,N_8450);
or U10000 (N_10000,N_9816,N_9122);
or U10001 (N_10001,N_9817,N_9377);
or U10002 (N_10002,N_9514,N_9685);
xnor U10003 (N_10003,N_9914,N_8805);
nor U10004 (N_10004,N_9114,N_9938);
nor U10005 (N_10005,N_9020,N_9118);
or U10006 (N_10006,N_9992,N_9522);
nand U10007 (N_10007,N_9135,N_9392);
nor U10008 (N_10008,N_9418,N_9765);
xor U10009 (N_10009,N_8912,N_8878);
xnor U10010 (N_10010,N_9443,N_9417);
xor U10011 (N_10011,N_9773,N_9137);
and U10012 (N_10012,N_9464,N_9103);
xor U10013 (N_10013,N_9111,N_9515);
xor U10014 (N_10014,N_9769,N_9278);
xnor U10015 (N_10015,N_9946,N_9391);
or U10016 (N_10016,N_9008,N_9825);
xnor U10017 (N_10017,N_9529,N_9584);
nor U10018 (N_10018,N_9566,N_9186);
xor U10019 (N_10019,N_9979,N_9876);
nand U10020 (N_10020,N_9797,N_9722);
or U10021 (N_10021,N_9751,N_9962);
nand U10022 (N_10022,N_9253,N_9244);
nor U10023 (N_10023,N_9156,N_9819);
nand U10024 (N_10024,N_8993,N_9198);
nand U10025 (N_10025,N_8972,N_9766);
or U10026 (N_10026,N_8864,N_8853);
and U10027 (N_10027,N_9617,N_9881);
or U10028 (N_10028,N_9396,N_8832);
xor U10029 (N_10029,N_9826,N_9295);
nand U10030 (N_10030,N_9098,N_8957);
xor U10031 (N_10031,N_9601,N_9900);
nor U10032 (N_10032,N_9034,N_8986);
nand U10033 (N_10033,N_8758,N_9344);
and U10034 (N_10034,N_8874,N_9864);
nand U10035 (N_10035,N_9126,N_9412);
nor U10036 (N_10036,N_9154,N_9559);
or U10037 (N_10037,N_9018,N_9021);
or U10038 (N_10038,N_9099,N_9645);
nand U10039 (N_10039,N_9586,N_9809);
and U10040 (N_10040,N_9376,N_8838);
or U10041 (N_10041,N_9243,N_8934);
nor U10042 (N_10042,N_9657,N_9503);
nor U10043 (N_10043,N_9678,N_9739);
nor U10044 (N_10044,N_9644,N_9889);
xnor U10045 (N_10045,N_9505,N_9270);
xnor U10046 (N_10046,N_8975,N_8795);
nand U10047 (N_10047,N_9594,N_9507);
nand U10048 (N_10048,N_9692,N_8911);
nor U10049 (N_10049,N_9955,N_9671);
or U10050 (N_10050,N_9228,N_9022);
and U10051 (N_10051,N_9466,N_8898);
and U10052 (N_10052,N_9052,N_9128);
xor U10053 (N_10053,N_9906,N_9481);
and U10054 (N_10054,N_9235,N_9368);
nor U10055 (N_10055,N_9339,N_8850);
and U10056 (N_10056,N_9375,N_9066);
nor U10057 (N_10057,N_8796,N_9266);
nor U10058 (N_10058,N_9095,N_8858);
and U10059 (N_10059,N_8777,N_9291);
xnor U10060 (N_10060,N_9465,N_9901);
or U10061 (N_10061,N_9595,N_9567);
or U10062 (N_10062,N_9406,N_9690);
nand U10063 (N_10063,N_9132,N_9611);
and U10064 (N_10064,N_8762,N_9632);
nor U10065 (N_10065,N_9129,N_8941);
xor U10066 (N_10066,N_9172,N_9106);
and U10067 (N_10067,N_9297,N_9776);
and U10068 (N_10068,N_9059,N_9957);
nand U10069 (N_10069,N_9770,N_9155);
and U10070 (N_10070,N_9312,N_9153);
nor U10071 (N_10071,N_8990,N_9738);
or U10072 (N_10072,N_9423,N_9063);
nand U10073 (N_10073,N_9878,N_8906);
nor U10074 (N_10074,N_9164,N_9110);
xor U10075 (N_10075,N_9163,N_9145);
xor U10076 (N_10076,N_8959,N_9745);
and U10077 (N_10077,N_9089,N_9355);
xor U10078 (N_10078,N_9585,N_8797);
or U10079 (N_10079,N_8902,N_9292);
or U10080 (N_10080,N_9072,N_8918);
xor U10081 (N_10081,N_9785,N_8835);
or U10082 (N_10082,N_8824,N_9065);
and U10083 (N_10083,N_9887,N_8991);
nor U10084 (N_10084,N_9252,N_9053);
xor U10085 (N_10085,N_9650,N_9613);
and U10086 (N_10086,N_9393,N_9610);
or U10087 (N_10087,N_9929,N_9786);
nand U10088 (N_10088,N_9943,N_9997);
xnor U10089 (N_10089,N_9225,N_9659);
and U10090 (N_10090,N_9171,N_9985);
and U10091 (N_10091,N_9910,N_9778);
nand U10092 (N_10092,N_8813,N_9397);
xnor U10093 (N_10093,N_9638,N_9415);
or U10094 (N_10094,N_9905,N_8879);
and U10095 (N_10095,N_8794,N_9345);
or U10096 (N_10096,N_9779,N_9774);
xnor U10097 (N_10097,N_9702,N_9044);
and U10098 (N_10098,N_9074,N_9994);
xnor U10099 (N_10099,N_9170,N_8877);
nand U10100 (N_10100,N_8892,N_8760);
or U10101 (N_10101,N_9724,N_9036);
xnor U10102 (N_10102,N_9472,N_9798);
and U10103 (N_10103,N_9913,N_9402);
nor U10104 (N_10104,N_9795,N_9080);
xnor U10105 (N_10105,N_9307,N_9136);
nor U10106 (N_10106,N_9551,N_9082);
nor U10107 (N_10107,N_8816,N_9879);
xnor U10108 (N_10108,N_8871,N_9840);
nand U10109 (N_10109,N_9682,N_9708);
and U10110 (N_10110,N_9248,N_9374);
xnor U10111 (N_10111,N_9272,N_9880);
xor U10112 (N_10112,N_9734,N_9832);
nand U10113 (N_10113,N_9823,N_9207);
or U10114 (N_10114,N_9311,N_9577);
nor U10115 (N_10115,N_9200,N_9653);
nor U10116 (N_10116,N_9771,N_9408);
nand U10117 (N_10117,N_8793,N_9075);
xor U10118 (N_10118,N_9356,N_8982);
nor U10119 (N_10119,N_9231,N_9602);
or U10120 (N_10120,N_9629,N_8828);
or U10121 (N_10121,N_9818,N_9283);
or U10122 (N_10122,N_9805,N_9214);
and U10123 (N_10123,N_8854,N_9705);
or U10124 (N_10124,N_9820,N_8951);
nand U10125 (N_10125,N_8889,N_9325);
and U10126 (N_10126,N_9860,N_9768);
or U10127 (N_10127,N_9326,N_9509);
and U10128 (N_10128,N_8984,N_9492);
xnor U10129 (N_10129,N_9750,N_9721);
nor U10130 (N_10130,N_9409,N_8910);
nor U10131 (N_10131,N_8946,N_9056);
xnor U10132 (N_10132,N_9564,N_8868);
nand U10133 (N_10133,N_9043,N_9570);
xor U10134 (N_10134,N_9027,N_9616);
and U10135 (N_10135,N_9411,N_8861);
or U10136 (N_10136,N_9201,N_8862);
and U10137 (N_10137,N_9933,N_8926);
nor U10138 (N_10138,N_9015,N_8952);
nand U10139 (N_10139,N_9333,N_9342);
or U10140 (N_10140,N_9512,N_9152);
nor U10141 (N_10141,N_9789,N_8856);
nor U10142 (N_10142,N_8843,N_9861);
nand U10143 (N_10143,N_9309,N_9358);
or U10144 (N_10144,N_9193,N_9643);
and U10145 (N_10145,N_9019,N_9160);
and U10146 (N_10146,N_8846,N_9433);
and U10147 (N_10147,N_9723,N_9640);
xor U10148 (N_10148,N_9633,N_9069);
and U10149 (N_10149,N_9932,N_9289);
or U10150 (N_10150,N_9926,N_9536);
and U10151 (N_10151,N_9016,N_8851);
or U10152 (N_10152,N_9084,N_9205);
xor U10153 (N_10153,N_9531,N_8833);
or U10154 (N_10154,N_9220,N_9500);
or U10155 (N_10155,N_9064,N_8875);
nor U10156 (N_10156,N_8936,N_9234);
or U10157 (N_10157,N_9484,N_9268);
and U10158 (N_10158,N_9664,N_8948);
xnor U10159 (N_10159,N_8921,N_9236);
nor U10160 (N_10160,N_9331,N_9183);
nand U10161 (N_10161,N_9538,N_8823);
xor U10162 (N_10162,N_9324,N_9005);
or U10163 (N_10163,N_9456,N_9212);
and U10164 (N_10164,N_9561,N_8989);
and U10165 (N_10165,N_9542,N_8869);
nand U10166 (N_10166,N_9867,N_9006);
and U10167 (N_10167,N_9775,N_9660);
nand U10168 (N_10168,N_9603,N_9918);
nor U10169 (N_10169,N_9865,N_9323);
or U10170 (N_10170,N_8790,N_8779);
and U10171 (N_10171,N_9141,N_8988);
nor U10172 (N_10172,N_9665,N_9092);
nand U10173 (N_10173,N_9907,N_9873);
or U10174 (N_10174,N_9953,N_9897);
or U10175 (N_10175,N_9589,N_9026);
nor U10176 (N_10176,N_8840,N_8970);
and U10177 (N_10177,N_9945,N_9274);
or U10178 (N_10178,N_8755,N_9387);
nor U10179 (N_10179,N_8787,N_9639);
nor U10180 (N_10180,N_9508,N_8827);
nor U10181 (N_10181,N_9810,N_9661);
and U10182 (N_10182,N_9454,N_9086);
and U10183 (N_10183,N_9647,N_9803);
xor U10184 (N_10184,N_9506,N_9223);
and U10185 (N_10185,N_8776,N_9458);
nor U10186 (N_10186,N_9176,N_9662);
nor U10187 (N_10187,N_9337,N_9516);
nor U10188 (N_10188,N_9365,N_9714);
and U10189 (N_10189,N_9988,N_9648);
and U10190 (N_10190,N_9029,N_9697);
nor U10191 (N_10191,N_9711,N_9502);
or U10192 (N_10192,N_8927,N_9002);
or U10193 (N_10193,N_9038,N_9814);
nand U10194 (N_10194,N_9909,N_9035);
and U10195 (N_10195,N_9378,N_9104);
or U10196 (N_10196,N_9039,N_9666);
and U10197 (N_10197,N_9058,N_8935);
xnor U10198 (N_10198,N_9047,N_9130);
nand U10199 (N_10199,N_9424,N_9085);
and U10200 (N_10200,N_8981,N_8891);
or U10201 (N_10201,N_9032,N_9960);
nand U10202 (N_10202,N_8973,N_8907);
and U10203 (N_10203,N_9582,N_9190);
nand U10204 (N_10204,N_9302,N_9485);
nor U10205 (N_10205,N_8860,N_9476);
nor U10206 (N_10206,N_9802,N_9419);
nor U10207 (N_10207,N_9158,N_9781);
nor U10208 (N_10208,N_9833,N_9656);
nand U10209 (N_10209,N_8817,N_9849);
nand U10210 (N_10210,N_9294,N_8826);
xor U10211 (N_10211,N_9247,N_9313);
and U10212 (N_10212,N_9090,N_9389);
xnor U10213 (N_10213,N_9438,N_9699);
nand U10214 (N_10214,N_8999,N_9563);
nor U10215 (N_10215,N_9608,N_9287);
nand U10216 (N_10216,N_9232,N_9532);
and U10217 (N_10217,N_9706,N_9893);
nand U10218 (N_10218,N_9490,N_9218);
nand U10219 (N_10219,N_9894,N_9037);
and U10220 (N_10220,N_9627,N_9348);
nand U10221 (N_10221,N_8782,N_9859);
xnor U10222 (N_10222,N_9870,N_9413);
xnor U10223 (N_10223,N_9761,N_9187);
or U10224 (N_10224,N_9545,N_8844);
nand U10225 (N_10225,N_9354,N_8766);
and U10226 (N_10226,N_9868,N_9742);
and U10227 (N_10227,N_9477,N_9442);
nand U10228 (N_10228,N_8998,N_8802);
and U10229 (N_10229,N_9794,N_9612);
nor U10230 (N_10230,N_9139,N_8945);
nor U10231 (N_10231,N_9550,N_9320);
or U10232 (N_10232,N_9952,N_9680);
nor U10233 (N_10233,N_9581,N_9941);
nand U10234 (N_10234,N_9917,N_9405);
xor U10235 (N_10235,N_9281,N_9314);
nor U10236 (N_10236,N_9524,N_9931);
xnor U10237 (N_10237,N_9134,N_8808);
nand U10238 (N_10238,N_9336,N_9959);
nor U10239 (N_10239,N_9679,N_8820);
nor U10240 (N_10240,N_9970,N_9166);
nor U10241 (N_10241,N_9296,N_9984);
xor U10242 (N_10242,N_9731,N_8914);
nor U10243 (N_10243,N_8801,N_9630);
or U10244 (N_10244,N_9669,N_8958);
and U10245 (N_10245,N_9259,N_9804);
or U10246 (N_10246,N_9410,N_8809);
xnor U10247 (N_10247,N_9380,N_9950);
or U10248 (N_10248,N_9691,N_9730);
or U10249 (N_10249,N_9591,N_9912);
or U10250 (N_10250,N_9927,N_9045);
or U10251 (N_10251,N_9548,N_9684);
nand U10252 (N_10252,N_9222,N_9604);
nor U10253 (N_10253,N_9807,N_9256);
or U10254 (N_10254,N_9535,N_9670);
nor U10255 (N_10255,N_9767,N_9758);
nand U10256 (N_10256,N_8822,N_9527);
and U10257 (N_10257,N_9240,N_9319);
nor U10258 (N_10258,N_9523,N_9199);
or U10259 (N_10259,N_9254,N_8847);
nor U10260 (N_10260,N_8894,N_8916);
xor U10261 (N_10261,N_9364,N_9401);
nand U10262 (N_10262,N_9973,N_9216);
xor U10263 (N_10263,N_9431,N_9658);
and U10264 (N_10264,N_9206,N_9108);
nand U10265 (N_10265,N_9347,N_8899);
or U10266 (N_10266,N_9173,N_9701);
xor U10267 (N_10267,N_8873,N_9123);
and U10268 (N_10268,N_9133,N_9150);
and U10269 (N_10269,N_9635,N_8919);
or U10270 (N_10270,N_9367,N_9293);
nor U10271 (N_10271,N_9203,N_9196);
or U10272 (N_10272,N_8947,N_8929);
and U10273 (N_10273,N_8992,N_9161);
or U10274 (N_10274,N_8956,N_8922);
xnor U10275 (N_10275,N_9185,N_9017);
and U10276 (N_10276,N_9855,N_9882);
nor U10277 (N_10277,N_9383,N_9366);
nor U10278 (N_10278,N_9245,N_9330);
nand U10279 (N_10279,N_9470,N_9899);
nor U10280 (N_10280,N_9578,N_9471);
nor U10281 (N_10281,N_9167,N_9197);
and U10282 (N_10282,N_9087,N_9384);
nand U10283 (N_10283,N_9068,N_9300);
xor U10284 (N_10284,N_9195,N_9261);
nor U10285 (N_10285,N_8821,N_8799);
nor U10286 (N_10286,N_8750,N_9273);
nor U10287 (N_10287,N_9863,N_9360);
and U10288 (N_10288,N_8996,N_9636);
and U10289 (N_10289,N_9760,N_9696);
nand U10290 (N_10290,N_8841,N_9838);
nand U10291 (N_10291,N_9713,N_8839);
and U10292 (N_10292,N_9262,N_9530);
or U10293 (N_10293,N_9057,N_8849);
and U10294 (N_10294,N_9131,N_8870);
or U10295 (N_10295,N_9381,N_9028);
nor U10296 (N_10296,N_8950,N_9501);
or U10297 (N_10297,N_9127,N_9568);
nor U10298 (N_10298,N_9519,N_8814);
nor U10299 (N_10299,N_9965,N_9012);
nand U10300 (N_10300,N_9625,N_9491);
xor U10301 (N_10301,N_9862,N_9306);
or U10302 (N_10302,N_9482,N_9301);
nor U10303 (N_10303,N_9493,N_9263);
xor U10304 (N_10304,N_8834,N_9971);
or U10305 (N_10305,N_9553,N_9908);
nor U10306 (N_10306,N_9168,N_9483);
nor U10307 (N_10307,N_9400,N_8818);
nor U10308 (N_10308,N_9569,N_9974);
or U10309 (N_10309,N_9457,N_8836);
xor U10310 (N_10310,N_9762,N_9451);
or U10311 (N_10311,N_9772,N_9871);
or U10312 (N_10312,N_9023,N_9782);
nor U10313 (N_10313,N_9736,N_8830);
or U10314 (N_10314,N_8983,N_8882);
xnor U10315 (N_10315,N_9606,N_9054);
and U10316 (N_10316,N_9432,N_9487);
nor U10317 (N_10317,N_9041,N_9416);
xnor U10318 (N_10318,N_9159,N_8798);
nand U10319 (N_10319,N_9049,N_9618);
nand U10320 (N_10320,N_9688,N_9208);
or U10321 (N_10321,N_9732,N_9479);
nor U10322 (N_10322,N_8944,N_9703);
or U10323 (N_10323,N_9600,N_9162);
and U10324 (N_10324,N_9654,N_9846);
and U10325 (N_10325,N_8803,N_9352);
nor U10326 (N_10326,N_9452,N_9073);
nor U10327 (N_10327,N_8893,N_9982);
or U10328 (N_10328,N_9681,N_8763);
or U10329 (N_10329,N_9321,N_9753);
or U10330 (N_10330,N_9042,N_9242);
xnor U10331 (N_10331,N_9362,N_9717);
xnor U10332 (N_10332,N_9728,N_9940);
nor U10333 (N_10333,N_8812,N_9229);
xor U10334 (N_10334,N_9290,N_9450);
and U10335 (N_10335,N_9888,N_8938);
and U10336 (N_10336,N_8961,N_9983);
and U10337 (N_10337,N_9398,N_9828);
and U10338 (N_10338,N_9842,N_9791);
xnor U10339 (N_10339,N_9841,N_9796);
xnor U10340 (N_10340,N_9105,N_9284);
nor U10341 (N_10341,N_9898,N_9689);
and U10342 (N_10342,N_8757,N_9441);
nor U10343 (N_10343,N_9009,N_9449);
xor U10344 (N_10344,N_9546,N_9373);
and U10345 (N_10345,N_9874,N_8829);
xor U10346 (N_10346,N_9783,N_9904);
or U10347 (N_10347,N_9718,N_9372);
nor U10348 (N_10348,N_9265,N_9989);
and U10349 (N_10349,N_9621,N_8971);
or U10350 (N_10350,N_9537,N_9831);
nand U10351 (N_10351,N_9539,N_8789);
nor U10352 (N_10352,N_9202,N_9921);
xor U10353 (N_10353,N_9672,N_9544);
or U10354 (N_10354,N_9866,N_9540);
xnor U10355 (N_10355,N_9445,N_9003);
or U10356 (N_10356,N_8977,N_9067);
or U10357 (N_10357,N_9453,N_9673);
and U10358 (N_10358,N_9676,N_9649);
nand U10359 (N_10359,N_8881,N_8885);
nand U10360 (N_10360,N_8754,N_9322);
nand U10361 (N_10361,N_9478,N_9497);
and U10362 (N_10362,N_9520,N_8859);
nand U10363 (N_10363,N_9191,N_9007);
xor U10364 (N_10364,N_8940,N_9759);
and U10365 (N_10365,N_9115,N_9787);
nor U10366 (N_10366,N_9050,N_8774);
nor U10367 (N_10367,N_9716,N_9857);
and U10368 (N_10368,N_9720,N_9175);
nand U10369 (N_10369,N_8985,N_9936);
nor U10370 (N_10370,N_9693,N_9010);
nand U10371 (N_10371,N_9250,N_9780);
xor U10372 (N_10372,N_9436,N_9174);
nor U10373 (N_10373,N_9588,N_9430);
xor U10374 (N_10374,N_9428,N_9046);
xnor U10375 (N_10375,N_9459,N_8764);
and U10376 (N_10376,N_9213,N_9386);
or U10377 (N_10377,N_8756,N_9226);
and U10378 (N_10378,N_9844,N_9737);
or U10379 (N_10379,N_9615,N_9088);
nand U10380 (N_10380,N_9641,N_9024);
nand U10381 (N_10381,N_8807,N_8968);
nor U10382 (N_10382,N_9598,N_8752);
nor U10383 (N_10383,N_9363,N_9964);
or U10384 (N_10384,N_9217,N_8932);
or U10385 (N_10385,N_9286,N_9461);
or U10386 (N_10386,N_9157,N_9475);
nand U10387 (N_10387,N_9267,N_9510);
nor U10388 (N_10388,N_9390,N_8930);
xor U10389 (N_10389,N_9729,N_8953);
xor U10390 (N_10390,N_9260,N_9277);
nand U10391 (N_10391,N_9683,N_9148);
xnor U10392 (N_10392,N_9623,N_8905);
nand U10393 (N_10393,N_9496,N_9467);
or U10394 (N_10394,N_8837,N_9435);
or U10395 (N_10395,N_9219,N_9583);
and U10396 (N_10396,N_9102,N_9719);
and U10397 (N_10397,N_8886,N_8772);
nand U10398 (N_10398,N_9258,N_9958);
xnor U10399 (N_10399,N_9975,N_9460);
xnor U10400 (N_10400,N_8960,N_8939);
xnor U10401 (N_10401,N_9562,N_9837);
nor U10402 (N_10402,N_9555,N_9712);
xor U10403 (N_10403,N_9756,N_9239);
xnor U10404 (N_10404,N_9579,N_9427);
xnor U10405 (N_10405,N_8759,N_9305);
or U10406 (N_10406,N_9070,N_9829);
nand U10407 (N_10407,N_9434,N_9609);
or U10408 (N_10408,N_9246,N_9593);
xnor U10409 (N_10409,N_9238,N_8887);
nor U10410 (N_10410,N_9061,N_8933);
or U10411 (N_10411,N_9571,N_8791);
and U10412 (N_10412,N_8848,N_9151);
and U10413 (N_10413,N_9093,N_9851);
and U10414 (N_10414,N_9192,N_9533);
nor U10415 (N_10415,N_9303,N_9149);
nand U10416 (N_10416,N_8866,N_8872);
or U10417 (N_10417,N_9715,N_9329);
or U10418 (N_10418,N_9969,N_9308);
nand U10419 (N_10419,N_9597,N_8857);
and U10420 (N_10420,N_9437,N_8753);
nor U10421 (N_10421,N_8903,N_9637);
or U10422 (N_10422,N_8995,N_9013);
nor U10423 (N_10423,N_9793,N_9463);
nand U10424 (N_10424,N_9668,N_9839);
xnor U10425 (N_10425,N_9651,N_9967);
nor U10426 (N_10426,N_9079,N_9474);
xnor U10427 (N_10427,N_9369,N_9554);
xnor U10428 (N_10428,N_9513,N_9001);
or U10429 (N_10429,N_9448,N_8969);
nand U10430 (N_10430,N_9182,N_9343);
or U10431 (N_10431,N_9394,N_9875);
or U10432 (N_10432,N_9573,N_8867);
nor U10433 (N_10433,N_9221,N_9920);
nand U10434 (N_10434,N_9987,N_9556);
nor U10435 (N_10435,N_9947,N_9371);
and U10436 (N_10436,N_9830,N_9891);
xnor U10437 (N_10437,N_9580,N_9704);
nor U10438 (N_10438,N_9279,N_9446);
or U10439 (N_10439,N_9511,N_9499);
or U10440 (N_10440,N_9966,N_9993);
nand U10441 (N_10441,N_9119,N_8997);
or U10442 (N_10442,N_8884,N_9370);
and U10443 (N_10443,N_9425,N_9599);
nor U10444 (N_10444,N_9178,N_9264);
and U10445 (N_10445,N_9241,N_9469);
nand U10446 (N_10446,N_9977,N_9572);
xnor U10447 (N_10447,N_8786,N_9557);
nor U10448 (N_10448,N_9144,N_8931);
or U10449 (N_10449,N_9414,N_9146);
and U10450 (N_10450,N_8783,N_8785);
nand U10451 (N_10451,N_8962,N_9784);
nand U10452 (N_10452,N_9327,N_9674);
and U10453 (N_10453,N_8980,N_9961);
nand U10454 (N_10454,N_9619,N_9318);
nor U10455 (N_10455,N_9925,N_9000);
nor U10456 (N_10456,N_9147,N_9030);
or U10457 (N_10457,N_8778,N_9317);
nand U10458 (N_10458,N_9815,N_9025);
xnor U10459 (N_10459,N_8876,N_9298);
xor U10460 (N_10460,N_9518,N_9922);
and U10461 (N_10461,N_9605,N_9255);
nor U10462 (N_10462,N_9097,N_8966);
xnor U10463 (N_10463,N_9112,N_9338);
nor U10464 (N_10464,N_8880,N_9916);
xor U10465 (N_10465,N_9655,N_9942);
xnor U10466 (N_10466,N_9930,N_9121);
or U10467 (N_10467,N_9677,N_8978);
and U10468 (N_10468,N_9934,N_8920);
nand U10469 (N_10469,N_8771,N_9488);
or U10470 (N_10470,N_8942,N_9299);
nor U10471 (N_10471,N_9468,N_9835);
nor U10472 (N_10472,N_9328,N_8804);
xnor U10473 (N_10473,N_9040,N_9634);
or U10474 (N_10474,N_9801,N_9346);
nor U10475 (N_10475,N_9349,N_8806);
nand U10476 (N_10476,N_9116,N_8917);
and U10477 (N_10477,N_9525,N_9340);
nand U10478 (N_10478,N_9473,N_9560);
or U10479 (N_10479,N_9790,N_9071);
nor U10480 (N_10480,N_9822,N_9140);
nand U10481 (N_10481,N_8965,N_9062);
xor U10482 (N_10482,N_9420,N_9237);
nor U10483 (N_10483,N_9051,N_9725);
and U10484 (N_10484,N_9972,N_8896);
nand U10485 (N_10485,N_9854,N_9179);
nor U10486 (N_10486,N_8811,N_8937);
and U10487 (N_10487,N_9494,N_9495);
xnor U10488 (N_10488,N_8987,N_9078);
nand U10489 (N_10489,N_9120,N_9727);
nand U10490 (N_10490,N_8788,N_9209);
nor U10491 (N_10491,N_8761,N_9091);
and U10492 (N_10492,N_9885,N_9504);
and U10493 (N_10493,N_8773,N_8775);
nor U10494 (N_10494,N_9575,N_9915);
or U10495 (N_10495,N_9902,N_9251);
or U10496 (N_10496,N_8904,N_9033);
and U10497 (N_10497,N_9361,N_9903);
xnor U10498 (N_10498,N_8909,N_9543);
nand U10499 (N_10499,N_8943,N_9836);
and U10500 (N_10500,N_9565,N_9194);
nand U10501 (N_10501,N_8770,N_8792);
xnor U10502 (N_10502,N_9357,N_9698);
nand U10503 (N_10503,N_9924,N_9403);
nor U10504 (N_10504,N_9271,N_9694);
xor U10505 (N_10505,N_9892,N_9048);
nand U10506 (N_10506,N_9498,N_9843);
or U10507 (N_10507,N_8800,N_9895);
and U10508 (N_10508,N_9777,N_9877);
nand U10509 (N_10509,N_8897,N_9998);
nor U10510 (N_10510,N_9276,N_9596);
nand U10511 (N_10511,N_9549,N_9142);
and U10512 (N_10512,N_9848,N_8784);
xor U10513 (N_10513,N_9620,N_9275);
nand U10514 (N_10514,N_9031,N_8767);
xor U10515 (N_10515,N_9060,N_9847);
xor U10516 (N_10516,N_9890,N_9856);
nand U10517 (N_10517,N_9227,N_9757);
and U10518 (N_10518,N_9455,N_9353);
xor U10519 (N_10519,N_9304,N_9334);
and U10520 (N_10520,N_8819,N_9911);
and U10521 (N_10521,N_9076,N_9257);
and U10522 (N_10522,N_8976,N_9686);
xnor U10523 (N_10523,N_9886,N_9919);
nor U10524 (N_10524,N_8925,N_9351);
nand U10525 (N_10525,N_9944,N_9138);
xnor U10526 (N_10526,N_9749,N_9980);
nor U10527 (N_10527,N_9675,N_9752);
xor U10528 (N_10528,N_9552,N_9986);
and U10529 (N_10529,N_9990,N_9642);
nand U10530 (N_10530,N_9489,N_9746);
or U10531 (N_10531,N_9101,N_9928);
nand U10532 (N_10532,N_9935,N_9687);
nand U10533 (N_10533,N_9646,N_9821);
nor U10534 (N_10534,N_9741,N_9624);
nor U10535 (N_10535,N_9956,N_9124);
nor U10536 (N_10536,N_8883,N_9249);
nand U10537 (N_10537,N_8954,N_9592);
and U10538 (N_10538,N_9447,N_9444);
nand U10539 (N_10539,N_9341,N_8895);
or U10540 (N_10540,N_8855,N_9695);
nand U10541 (N_10541,N_9014,N_9827);
xnor U10542 (N_10542,N_9981,N_9845);
nor U10543 (N_10543,N_9735,N_9335);
xnor U10544 (N_10544,N_9521,N_9100);
xor U10545 (N_10545,N_9954,N_8963);
and U10546 (N_10546,N_9663,N_9350);
and U10547 (N_10547,N_9763,N_9165);
or U10548 (N_10548,N_9824,N_8845);
nor U10549 (N_10549,N_9884,N_8890);
xor U10550 (N_10550,N_9747,N_9896);
and U10551 (N_10551,N_9385,N_9733);
nand U10552 (N_10552,N_8924,N_9421);
and U10553 (N_10553,N_9652,N_9404);
nand U10554 (N_10554,N_9576,N_9230);
and U10555 (N_10555,N_9107,N_8974);
or U10556 (N_10556,N_9177,N_9744);
nand U10557 (N_10557,N_8831,N_8979);
xor U10558 (N_10558,N_9285,N_9590);
xor U10559 (N_10559,N_9883,N_9462);
or U10560 (N_10560,N_9799,N_9188);
nand U10561 (N_10561,N_9631,N_9233);
nor U10562 (N_10562,N_9976,N_9316);
nor U10563 (N_10563,N_8964,N_8923);
nor U10564 (N_10564,N_9211,N_9109);
and U10565 (N_10565,N_9743,N_9978);
xnor U10566 (N_10566,N_9991,N_9923);
or U10567 (N_10567,N_9528,N_9755);
nand U10568 (N_10568,N_9614,N_9858);
nor U10569 (N_10569,N_9143,N_9748);
nor U10570 (N_10570,N_9407,N_8810);
or U10571 (N_10571,N_9184,N_9288);
nor U10572 (N_10572,N_9709,N_8865);
nor U10573 (N_10573,N_9181,N_9440);
xnor U10574 (N_10574,N_9332,N_9754);
xor U10575 (N_10575,N_9834,N_8825);
nor U10576 (N_10576,N_8955,N_9426);
nand U10577 (N_10577,N_9740,N_9282);
nand U10578 (N_10578,N_9169,N_9077);
nor U10579 (N_10579,N_9710,N_9853);
or U10580 (N_10580,N_8900,N_8751);
xnor U10581 (N_10581,N_9558,N_9949);
or U10582 (N_10582,N_9204,N_9083);
nor U10583 (N_10583,N_8842,N_8768);
and U10584 (N_10584,N_9094,N_9996);
nor U10585 (N_10585,N_9269,N_9395);
or U10586 (N_10586,N_9937,N_9869);
nand U10587 (N_10587,N_9399,N_9948);
or U10588 (N_10588,N_9574,N_9999);
or U10589 (N_10589,N_8888,N_9382);
nor U10590 (N_10590,N_8863,N_8928);
xnor U10591 (N_10591,N_9180,N_9526);
nand U10592 (N_10592,N_9004,N_8769);
or U10593 (N_10593,N_8781,N_9280);
and U10594 (N_10594,N_8908,N_9315);
nand U10595 (N_10595,N_9125,N_9963);
xnor U10596 (N_10596,N_9011,N_9359);
nand U10597 (N_10597,N_8915,N_9517);
or U10598 (N_10598,N_9726,N_9429);
nor U10599 (N_10599,N_9310,N_9486);
or U10600 (N_10600,N_9872,N_9995);
nand U10601 (N_10601,N_9788,N_9764);
or U10602 (N_10602,N_9813,N_9534);
nand U10603 (N_10603,N_9096,N_9850);
xnor U10604 (N_10604,N_9667,N_8815);
xor U10605 (N_10605,N_9628,N_9806);
or U10606 (N_10606,N_8994,N_9215);
nand U10607 (N_10607,N_9388,N_9480);
nand U10608 (N_10608,N_9811,N_9968);
nor U10609 (N_10609,N_9607,N_8967);
nor U10610 (N_10610,N_9189,N_8852);
and U10611 (N_10611,N_9081,N_8765);
or U10612 (N_10612,N_9700,N_9210);
or U10613 (N_10613,N_9055,N_9224);
nand U10614 (N_10614,N_8780,N_9422);
nor U10615 (N_10615,N_8901,N_9439);
and U10616 (N_10616,N_9113,N_8913);
or U10617 (N_10617,N_9812,N_9626);
nand U10618 (N_10618,N_9117,N_9939);
or U10619 (N_10619,N_9800,N_9951);
nand U10620 (N_10620,N_9379,N_9547);
nand U10621 (N_10621,N_9808,N_8949);
nand U10622 (N_10622,N_9587,N_9622);
and U10623 (N_10623,N_9707,N_9852);
or U10624 (N_10624,N_9792,N_9541);
xor U10625 (N_10625,N_9360,N_9919);
nor U10626 (N_10626,N_9842,N_9016);
xor U10627 (N_10627,N_9497,N_9500);
nand U10628 (N_10628,N_9485,N_9895);
nor U10629 (N_10629,N_9806,N_9928);
and U10630 (N_10630,N_8885,N_8948);
nand U10631 (N_10631,N_9338,N_9204);
or U10632 (N_10632,N_9450,N_9590);
nor U10633 (N_10633,N_9332,N_9736);
and U10634 (N_10634,N_9257,N_8943);
nor U10635 (N_10635,N_9440,N_9263);
xor U10636 (N_10636,N_9325,N_9176);
and U10637 (N_10637,N_9437,N_9071);
xor U10638 (N_10638,N_8904,N_8886);
xor U10639 (N_10639,N_9714,N_9977);
or U10640 (N_10640,N_9376,N_9410);
nor U10641 (N_10641,N_9865,N_8768);
and U10642 (N_10642,N_8884,N_9955);
nand U10643 (N_10643,N_9175,N_8872);
or U10644 (N_10644,N_9722,N_9307);
or U10645 (N_10645,N_9457,N_9321);
or U10646 (N_10646,N_8902,N_8943);
nand U10647 (N_10647,N_9461,N_9954);
nand U10648 (N_10648,N_8754,N_9062);
and U10649 (N_10649,N_8850,N_9240);
nand U10650 (N_10650,N_9684,N_9865);
nand U10651 (N_10651,N_9290,N_9309);
xor U10652 (N_10652,N_9477,N_9403);
nor U10653 (N_10653,N_9413,N_9685);
xnor U10654 (N_10654,N_8890,N_8909);
and U10655 (N_10655,N_8991,N_8841);
or U10656 (N_10656,N_9174,N_9753);
nor U10657 (N_10657,N_9944,N_9255);
nor U10658 (N_10658,N_9504,N_9472);
xor U10659 (N_10659,N_9753,N_9201);
nand U10660 (N_10660,N_9584,N_9504);
nand U10661 (N_10661,N_9672,N_9265);
xnor U10662 (N_10662,N_9097,N_9709);
xor U10663 (N_10663,N_9502,N_9029);
nor U10664 (N_10664,N_9243,N_9681);
and U10665 (N_10665,N_9870,N_8846);
or U10666 (N_10666,N_9626,N_9078);
and U10667 (N_10667,N_9479,N_9348);
nor U10668 (N_10668,N_9070,N_9210);
xnor U10669 (N_10669,N_8991,N_9855);
or U10670 (N_10670,N_9005,N_9810);
nand U10671 (N_10671,N_9373,N_9593);
or U10672 (N_10672,N_9068,N_9134);
and U10673 (N_10673,N_9789,N_9704);
and U10674 (N_10674,N_8828,N_9731);
nor U10675 (N_10675,N_9841,N_9229);
xnor U10676 (N_10676,N_9967,N_9442);
nand U10677 (N_10677,N_9014,N_9077);
or U10678 (N_10678,N_9028,N_9087);
xor U10679 (N_10679,N_9848,N_9284);
nand U10680 (N_10680,N_8779,N_9765);
or U10681 (N_10681,N_8943,N_9913);
and U10682 (N_10682,N_9403,N_9038);
or U10683 (N_10683,N_8824,N_9156);
nand U10684 (N_10684,N_9360,N_9986);
nand U10685 (N_10685,N_9451,N_9606);
xor U10686 (N_10686,N_8860,N_8767);
or U10687 (N_10687,N_9275,N_8882);
xnor U10688 (N_10688,N_8763,N_9995);
nand U10689 (N_10689,N_9493,N_9912);
nor U10690 (N_10690,N_9604,N_8820);
or U10691 (N_10691,N_8846,N_9263);
xnor U10692 (N_10692,N_8788,N_9085);
nor U10693 (N_10693,N_9564,N_9649);
xor U10694 (N_10694,N_9655,N_8939);
nand U10695 (N_10695,N_9458,N_9461);
xnor U10696 (N_10696,N_9614,N_9667);
nand U10697 (N_10697,N_9760,N_8848);
nand U10698 (N_10698,N_9179,N_8803);
nor U10699 (N_10699,N_9064,N_9476);
nor U10700 (N_10700,N_9407,N_9983);
nor U10701 (N_10701,N_8889,N_9167);
nor U10702 (N_10702,N_8810,N_8984);
nor U10703 (N_10703,N_9836,N_9058);
nor U10704 (N_10704,N_9104,N_8850);
nand U10705 (N_10705,N_9937,N_9850);
nor U10706 (N_10706,N_9740,N_9763);
nand U10707 (N_10707,N_9580,N_9963);
and U10708 (N_10708,N_9095,N_9084);
and U10709 (N_10709,N_9645,N_8758);
and U10710 (N_10710,N_9395,N_8786);
and U10711 (N_10711,N_9694,N_9026);
and U10712 (N_10712,N_9265,N_9828);
xor U10713 (N_10713,N_9382,N_9283);
or U10714 (N_10714,N_8945,N_9003);
nor U10715 (N_10715,N_9015,N_8934);
and U10716 (N_10716,N_9247,N_9746);
and U10717 (N_10717,N_9217,N_9423);
nand U10718 (N_10718,N_9270,N_9844);
or U10719 (N_10719,N_8832,N_8956);
and U10720 (N_10720,N_9861,N_9827);
nand U10721 (N_10721,N_9071,N_9652);
nand U10722 (N_10722,N_9273,N_8985);
xor U10723 (N_10723,N_8924,N_9426);
xnor U10724 (N_10724,N_9178,N_8779);
nand U10725 (N_10725,N_9443,N_9483);
nor U10726 (N_10726,N_9456,N_9955);
nor U10727 (N_10727,N_9428,N_9663);
or U10728 (N_10728,N_9201,N_9714);
or U10729 (N_10729,N_9894,N_9054);
or U10730 (N_10730,N_9876,N_9140);
or U10731 (N_10731,N_9995,N_9071);
or U10732 (N_10732,N_9234,N_8877);
and U10733 (N_10733,N_9327,N_9528);
xor U10734 (N_10734,N_9850,N_9792);
nor U10735 (N_10735,N_9563,N_9469);
xnor U10736 (N_10736,N_9239,N_8774);
or U10737 (N_10737,N_9055,N_9923);
nand U10738 (N_10738,N_9176,N_9608);
or U10739 (N_10739,N_8768,N_9757);
xor U10740 (N_10740,N_9508,N_8878);
nor U10741 (N_10741,N_9800,N_8820);
nor U10742 (N_10742,N_8823,N_9692);
xor U10743 (N_10743,N_8874,N_8897);
nand U10744 (N_10744,N_9486,N_9524);
nand U10745 (N_10745,N_9699,N_9709);
and U10746 (N_10746,N_9079,N_9102);
and U10747 (N_10747,N_9721,N_9588);
and U10748 (N_10748,N_9465,N_9752);
nand U10749 (N_10749,N_9994,N_9693);
and U10750 (N_10750,N_9715,N_9164);
nor U10751 (N_10751,N_9415,N_9978);
xnor U10752 (N_10752,N_9655,N_9097);
or U10753 (N_10753,N_9557,N_8964);
nand U10754 (N_10754,N_9849,N_9113);
or U10755 (N_10755,N_9543,N_9528);
and U10756 (N_10756,N_9024,N_9978);
or U10757 (N_10757,N_9124,N_9816);
and U10758 (N_10758,N_9195,N_9677);
and U10759 (N_10759,N_9050,N_9714);
xnor U10760 (N_10760,N_8757,N_9237);
nand U10761 (N_10761,N_9699,N_9527);
and U10762 (N_10762,N_9013,N_9422);
and U10763 (N_10763,N_9522,N_9851);
xnor U10764 (N_10764,N_9123,N_9761);
nor U10765 (N_10765,N_8795,N_9578);
or U10766 (N_10766,N_8755,N_8963);
nor U10767 (N_10767,N_9242,N_9761);
nand U10768 (N_10768,N_9762,N_9348);
xor U10769 (N_10769,N_9917,N_9339);
or U10770 (N_10770,N_9080,N_9504);
nor U10771 (N_10771,N_9744,N_8826);
nor U10772 (N_10772,N_9023,N_9792);
nor U10773 (N_10773,N_9188,N_9555);
nand U10774 (N_10774,N_9753,N_9157);
nor U10775 (N_10775,N_9490,N_9926);
or U10776 (N_10776,N_9109,N_8800);
and U10777 (N_10777,N_9202,N_9019);
xnor U10778 (N_10778,N_9937,N_9423);
or U10779 (N_10779,N_9629,N_9005);
nand U10780 (N_10780,N_9148,N_8890);
and U10781 (N_10781,N_9964,N_9225);
or U10782 (N_10782,N_9041,N_9347);
xnor U10783 (N_10783,N_9268,N_8759);
or U10784 (N_10784,N_9637,N_9207);
nor U10785 (N_10785,N_8982,N_9429);
and U10786 (N_10786,N_8827,N_9582);
nand U10787 (N_10787,N_9371,N_9497);
or U10788 (N_10788,N_9056,N_9842);
nand U10789 (N_10789,N_9601,N_9600);
and U10790 (N_10790,N_9026,N_9251);
and U10791 (N_10791,N_9703,N_9449);
nand U10792 (N_10792,N_9072,N_9615);
or U10793 (N_10793,N_9611,N_9421);
nor U10794 (N_10794,N_9581,N_9702);
or U10795 (N_10795,N_9485,N_8933);
and U10796 (N_10796,N_9640,N_8997);
xnor U10797 (N_10797,N_9203,N_9235);
and U10798 (N_10798,N_9508,N_9427);
nor U10799 (N_10799,N_8818,N_9247);
xnor U10800 (N_10800,N_8785,N_9342);
xor U10801 (N_10801,N_8858,N_8847);
or U10802 (N_10802,N_9470,N_9775);
or U10803 (N_10803,N_9353,N_9498);
or U10804 (N_10804,N_9051,N_9749);
and U10805 (N_10805,N_9470,N_9360);
and U10806 (N_10806,N_9621,N_9785);
and U10807 (N_10807,N_9348,N_9270);
nor U10808 (N_10808,N_9572,N_9096);
xor U10809 (N_10809,N_9455,N_9475);
xor U10810 (N_10810,N_8780,N_8918);
and U10811 (N_10811,N_9123,N_8996);
nor U10812 (N_10812,N_8897,N_9375);
or U10813 (N_10813,N_9702,N_9112);
and U10814 (N_10814,N_9946,N_9240);
nor U10815 (N_10815,N_9078,N_9674);
xnor U10816 (N_10816,N_9228,N_9083);
or U10817 (N_10817,N_9099,N_9891);
nand U10818 (N_10818,N_9233,N_9822);
nand U10819 (N_10819,N_9225,N_8761);
or U10820 (N_10820,N_9895,N_9847);
nand U10821 (N_10821,N_9495,N_9552);
or U10822 (N_10822,N_9055,N_9443);
or U10823 (N_10823,N_9478,N_9577);
and U10824 (N_10824,N_9144,N_8940);
nand U10825 (N_10825,N_9928,N_9102);
xnor U10826 (N_10826,N_9754,N_8880);
nand U10827 (N_10827,N_9298,N_9717);
nor U10828 (N_10828,N_9072,N_9768);
nor U10829 (N_10829,N_9923,N_9061);
or U10830 (N_10830,N_9759,N_8928);
xor U10831 (N_10831,N_8950,N_8855);
or U10832 (N_10832,N_9446,N_9044);
or U10833 (N_10833,N_8919,N_9207);
xnor U10834 (N_10834,N_8949,N_9013);
nor U10835 (N_10835,N_9748,N_9154);
xor U10836 (N_10836,N_9056,N_9441);
nor U10837 (N_10837,N_9568,N_9132);
or U10838 (N_10838,N_9793,N_9169);
or U10839 (N_10839,N_8988,N_9545);
nand U10840 (N_10840,N_9107,N_9351);
and U10841 (N_10841,N_9112,N_8845);
or U10842 (N_10842,N_9819,N_9328);
and U10843 (N_10843,N_8794,N_9325);
and U10844 (N_10844,N_8786,N_9037);
nand U10845 (N_10845,N_8781,N_9664);
and U10846 (N_10846,N_8769,N_8874);
nand U10847 (N_10847,N_9599,N_9517);
nand U10848 (N_10848,N_9623,N_9603);
or U10849 (N_10849,N_9152,N_9099);
xnor U10850 (N_10850,N_9758,N_9860);
and U10851 (N_10851,N_9162,N_9752);
nor U10852 (N_10852,N_9828,N_9526);
nand U10853 (N_10853,N_9432,N_9447);
nor U10854 (N_10854,N_9446,N_9693);
or U10855 (N_10855,N_9112,N_9211);
xor U10856 (N_10856,N_9685,N_9149);
xnor U10857 (N_10857,N_8847,N_9669);
or U10858 (N_10858,N_8918,N_9115);
or U10859 (N_10859,N_9157,N_9352);
nand U10860 (N_10860,N_9465,N_9822);
xor U10861 (N_10861,N_9352,N_9396);
or U10862 (N_10862,N_9923,N_9001);
nor U10863 (N_10863,N_9024,N_9739);
and U10864 (N_10864,N_9191,N_9977);
xor U10865 (N_10865,N_9090,N_9101);
nand U10866 (N_10866,N_8992,N_9862);
xnor U10867 (N_10867,N_8995,N_9744);
xnor U10868 (N_10868,N_9793,N_9687);
xnor U10869 (N_10869,N_9774,N_9255);
nand U10870 (N_10870,N_9121,N_9706);
nor U10871 (N_10871,N_8850,N_9844);
xnor U10872 (N_10872,N_9046,N_9316);
or U10873 (N_10873,N_9287,N_9066);
nand U10874 (N_10874,N_9194,N_8939);
and U10875 (N_10875,N_9135,N_9989);
and U10876 (N_10876,N_9976,N_8988);
nor U10877 (N_10877,N_9527,N_9099);
and U10878 (N_10878,N_9267,N_9729);
nand U10879 (N_10879,N_9072,N_8967);
xor U10880 (N_10880,N_9323,N_9097);
and U10881 (N_10881,N_8837,N_9521);
or U10882 (N_10882,N_9678,N_9947);
or U10883 (N_10883,N_9651,N_9064);
nand U10884 (N_10884,N_9051,N_8935);
xnor U10885 (N_10885,N_8820,N_9892);
xnor U10886 (N_10886,N_8789,N_9412);
and U10887 (N_10887,N_9446,N_8859);
xnor U10888 (N_10888,N_9057,N_9515);
and U10889 (N_10889,N_8928,N_9736);
and U10890 (N_10890,N_8963,N_8791);
nor U10891 (N_10891,N_9424,N_9984);
or U10892 (N_10892,N_9024,N_9487);
nor U10893 (N_10893,N_8927,N_9037);
and U10894 (N_10894,N_8943,N_9470);
xor U10895 (N_10895,N_9892,N_9600);
and U10896 (N_10896,N_9159,N_9261);
nand U10897 (N_10897,N_9689,N_9799);
nand U10898 (N_10898,N_9013,N_9152);
nor U10899 (N_10899,N_9553,N_9055);
or U10900 (N_10900,N_9167,N_9523);
and U10901 (N_10901,N_9259,N_9305);
nand U10902 (N_10902,N_9847,N_9574);
or U10903 (N_10903,N_9702,N_9115);
nand U10904 (N_10904,N_9242,N_9924);
or U10905 (N_10905,N_9896,N_9695);
and U10906 (N_10906,N_9563,N_9896);
or U10907 (N_10907,N_9411,N_9341);
xor U10908 (N_10908,N_9087,N_9601);
nand U10909 (N_10909,N_9084,N_9580);
nor U10910 (N_10910,N_8757,N_9260);
or U10911 (N_10911,N_9270,N_9121);
and U10912 (N_10912,N_8979,N_9375);
nand U10913 (N_10913,N_9722,N_9530);
nand U10914 (N_10914,N_9974,N_8906);
xor U10915 (N_10915,N_9197,N_9616);
nand U10916 (N_10916,N_9911,N_8920);
xnor U10917 (N_10917,N_9535,N_9017);
and U10918 (N_10918,N_9026,N_9525);
and U10919 (N_10919,N_9464,N_9131);
and U10920 (N_10920,N_9276,N_9305);
and U10921 (N_10921,N_9027,N_9257);
xnor U10922 (N_10922,N_9733,N_8961);
and U10923 (N_10923,N_9512,N_9122);
nand U10924 (N_10924,N_8772,N_9989);
and U10925 (N_10925,N_8833,N_8857);
xnor U10926 (N_10926,N_9220,N_8972);
and U10927 (N_10927,N_9616,N_9560);
nor U10928 (N_10928,N_9108,N_9442);
nor U10929 (N_10929,N_9402,N_9646);
and U10930 (N_10930,N_9341,N_9332);
nor U10931 (N_10931,N_9479,N_9812);
or U10932 (N_10932,N_9889,N_9267);
or U10933 (N_10933,N_9219,N_9057);
xor U10934 (N_10934,N_9392,N_9826);
or U10935 (N_10935,N_8889,N_9218);
xnor U10936 (N_10936,N_9627,N_9332);
nor U10937 (N_10937,N_9836,N_9095);
or U10938 (N_10938,N_9221,N_9327);
nand U10939 (N_10939,N_9184,N_9803);
nor U10940 (N_10940,N_9367,N_9540);
or U10941 (N_10941,N_9428,N_9489);
and U10942 (N_10942,N_9072,N_9306);
and U10943 (N_10943,N_8820,N_9978);
or U10944 (N_10944,N_9762,N_8865);
xnor U10945 (N_10945,N_9323,N_8957);
and U10946 (N_10946,N_9976,N_9396);
nor U10947 (N_10947,N_9402,N_9353);
and U10948 (N_10948,N_9020,N_9878);
nor U10949 (N_10949,N_9939,N_8997);
or U10950 (N_10950,N_8808,N_8757);
nand U10951 (N_10951,N_9436,N_8861);
nand U10952 (N_10952,N_8855,N_9878);
or U10953 (N_10953,N_9913,N_9669);
xor U10954 (N_10954,N_9796,N_9728);
or U10955 (N_10955,N_9446,N_9729);
nor U10956 (N_10956,N_9379,N_9095);
nor U10957 (N_10957,N_9374,N_8976);
or U10958 (N_10958,N_9458,N_9342);
or U10959 (N_10959,N_8971,N_9546);
and U10960 (N_10960,N_9288,N_9633);
nor U10961 (N_10961,N_9134,N_9858);
and U10962 (N_10962,N_8970,N_9667);
nor U10963 (N_10963,N_9269,N_9731);
nor U10964 (N_10964,N_8990,N_9764);
nand U10965 (N_10965,N_8803,N_9821);
and U10966 (N_10966,N_9680,N_9320);
and U10967 (N_10967,N_9632,N_9194);
nand U10968 (N_10968,N_9827,N_9126);
xnor U10969 (N_10969,N_9158,N_9309);
nand U10970 (N_10970,N_9042,N_9108);
nor U10971 (N_10971,N_8906,N_8894);
and U10972 (N_10972,N_9126,N_8851);
and U10973 (N_10973,N_9601,N_9211);
and U10974 (N_10974,N_9482,N_9169);
nand U10975 (N_10975,N_9475,N_9539);
xnor U10976 (N_10976,N_9245,N_9240);
or U10977 (N_10977,N_8975,N_9084);
nor U10978 (N_10978,N_8879,N_9296);
and U10979 (N_10979,N_9529,N_9431);
nor U10980 (N_10980,N_9380,N_8966);
xnor U10981 (N_10981,N_9312,N_9209);
nor U10982 (N_10982,N_9672,N_8890);
xnor U10983 (N_10983,N_9136,N_9033);
or U10984 (N_10984,N_9980,N_9998);
xor U10985 (N_10985,N_9898,N_8836);
or U10986 (N_10986,N_9429,N_8779);
xnor U10987 (N_10987,N_8916,N_9937);
and U10988 (N_10988,N_8909,N_9202);
nand U10989 (N_10989,N_9190,N_9235);
and U10990 (N_10990,N_9265,N_8872);
xnor U10991 (N_10991,N_9177,N_9600);
nand U10992 (N_10992,N_9863,N_9638);
nor U10993 (N_10993,N_9601,N_9270);
and U10994 (N_10994,N_8877,N_9292);
or U10995 (N_10995,N_9231,N_9208);
xnor U10996 (N_10996,N_9674,N_9091);
xor U10997 (N_10997,N_9858,N_9800);
and U10998 (N_10998,N_9622,N_9294);
xor U10999 (N_10999,N_9007,N_8881);
nor U11000 (N_11000,N_9336,N_9853);
and U11001 (N_11001,N_8773,N_9434);
xnor U11002 (N_11002,N_8967,N_9706);
xnor U11003 (N_11003,N_9993,N_9134);
nand U11004 (N_11004,N_8933,N_9474);
nor U11005 (N_11005,N_9830,N_9988);
nor U11006 (N_11006,N_8773,N_9376);
or U11007 (N_11007,N_8877,N_9161);
nor U11008 (N_11008,N_8871,N_9491);
nor U11009 (N_11009,N_9658,N_8926);
xnor U11010 (N_11010,N_9849,N_9678);
and U11011 (N_11011,N_9381,N_8814);
xor U11012 (N_11012,N_9051,N_9112);
nand U11013 (N_11013,N_9407,N_8764);
nand U11014 (N_11014,N_9016,N_8850);
or U11015 (N_11015,N_9291,N_9901);
and U11016 (N_11016,N_9278,N_9220);
or U11017 (N_11017,N_9608,N_8859);
xnor U11018 (N_11018,N_9721,N_9473);
nor U11019 (N_11019,N_9727,N_8928);
nor U11020 (N_11020,N_9550,N_9799);
or U11021 (N_11021,N_9551,N_8904);
nand U11022 (N_11022,N_9602,N_9084);
nand U11023 (N_11023,N_9469,N_9398);
xnor U11024 (N_11024,N_9070,N_9321);
or U11025 (N_11025,N_8866,N_9158);
nand U11026 (N_11026,N_9281,N_9476);
and U11027 (N_11027,N_9266,N_8779);
xnor U11028 (N_11028,N_9899,N_9453);
or U11029 (N_11029,N_9621,N_8826);
nand U11030 (N_11030,N_9149,N_8843);
and U11031 (N_11031,N_9398,N_9748);
and U11032 (N_11032,N_9562,N_9507);
nand U11033 (N_11033,N_9546,N_9046);
or U11034 (N_11034,N_8958,N_9154);
nand U11035 (N_11035,N_9737,N_9422);
xnor U11036 (N_11036,N_9839,N_9457);
xnor U11037 (N_11037,N_8938,N_9296);
or U11038 (N_11038,N_9388,N_9212);
xor U11039 (N_11039,N_8886,N_9308);
and U11040 (N_11040,N_9488,N_9852);
xnor U11041 (N_11041,N_9372,N_9917);
nor U11042 (N_11042,N_9455,N_9759);
nor U11043 (N_11043,N_9843,N_9329);
nand U11044 (N_11044,N_8909,N_9264);
and U11045 (N_11045,N_9289,N_9453);
and U11046 (N_11046,N_8800,N_9349);
xnor U11047 (N_11047,N_9674,N_9337);
or U11048 (N_11048,N_9766,N_9197);
nor U11049 (N_11049,N_8862,N_9331);
or U11050 (N_11050,N_8954,N_9322);
and U11051 (N_11051,N_9027,N_8755);
and U11052 (N_11052,N_9368,N_9593);
xor U11053 (N_11053,N_8865,N_9883);
xor U11054 (N_11054,N_9054,N_9591);
and U11055 (N_11055,N_9114,N_9446);
or U11056 (N_11056,N_9046,N_9664);
or U11057 (N_11057,N_9709,N_9954);
and U11058 (N_11058,N_8921,N_9012);
xnor U11059 (N_11059,N_8960,N_9121);
or U11060 (N_11060,N_9047,N_9692);
or U11061 (N_11061,N_9520,N_8953);
and U11062 (N_11062,N_9266,N_8842);
or U11063 (N_11063,N_9907,N_9918);
and U11064 (N_11064,N_9870,N_9083);
or U11065 (N_11065,N_9203,N_9086);
nor U11066 (N_11066,N_9663,N_9665);
xor U11067 (N_11067,N_8915,N_8828);
xor U11068 (N_11068,N_9257,N_9187);
xor U11069 (N_11069,N_9091,N_9828);
nor U11070 (N_11070,N_9672,N_8853);
nor U11071 (N_11071,N_9732,N_9067);
and U11072 (N_11072,N_8826,N_8757);
and U11073 (N_11073,N_9624,N_9996);
and U11074 (N_11074,N_9799,N_9924);
nor U11075 (N_11075,N_9501,N_9270);
nand U11076 (N_11076,N_9600,N_9296);
or U11077 (N_11077,N_9274,N_9907);
xor U11078 (N_11078,N_9392,N_9534);
nor U11079 (N_11079,N_8933,N_9008);
and U11080 (N_11080,N_9898,N_9002);
xnor U11081 (N_11081,N_9552,N_8927);
nor U11082 (N_11082,N_9263,N_9625);
xnor U11083 (N_11083,N_9617,N_9734);
nor U11084 (N_11084,N_9607,N_9495);
or U11085 (N_11085,N_8772,N_9416);
xnor U11086 (N_11086,N_9974,N_9793);
or U11087 (N_11087,N_9988,N_9372);
nand U11088 (N_11088,N_9347,N_8840);
nand U11089 (N_11089,N_9148,N_9850);
nand U11090 (N_11090,N_9300,N_9465);
xnor U11091 (N_11091,N_9721,N_9624);
nor U11092 (N_11092,N_9376,N_9732);
xnor U11093 (N_11093,N_9913,N_9547);
xor U11094 (N_11094,N_8828,N_9053);
xnor U11095 (N_11095,N_9171,N_9778);
nand U11096 (N_11096,N_8935,N_9703);
or U11097 (N_11097,N_9372,N_9668);
or U11098 (N_11098,N_9688,N_9820);
nor U11099 (N_11099,N_9027,N_9986);
nor U11100 (N_11100,N_9738,N_9172);
nor U11101 (N_11101,N_9532,N_9738);
and U11102 (N_11102,N_9949,N_9229);
nor U11103 (N_11103,N_8867,N_9953);
nand U11104 (N_11104,N_9939,N_9382);
and U11105 (N_11105,N_9302,N_8872);
or U11106 (N_11106,N_9928,N_9168);
or U11107 (N_11107,N_9963,N_9834);
and U11108 (N_11108,N_9588,N_9055);
or U11109 (N_11109,N_9557,N_9215);
or U11110 (N_11110,N_9686,N_9023);
nor U11111 (N_11111,N_9919,N_9323);
or U11112 (N_11112,N_9509,N_9555);
or U11113 (N_11113,N_8771,N_8917);
nor U11114 (N_11114,N_8915,N_8993);
or U11115 (N_11115,N_9423,N_9070);
nand U11116 (N_11116,N_9813,N_9369);
and U11117 (N_11117,N_9623,N_9663);
nand U11118 (N_11118,N_9076,N_9848);
xnor U11119 (N_11119,N_9081,N_8843);
or U11120 (N_11120,N_9325,N_9416);
or U11121 (N_11121,N_8857,N_9134);
nand U11122 (N_11122,N_9750,N_9014);
xor U11123 (N_11123,N_9686,N_8822);
or U11124 (N_11124,N_9228,N_9765);
xnor U11125 (N_11125,N_9558,N_9951);
xnor U11126 (N_11126,N_9595,N_8982);
nor U11127 (N_11127,N_9463,N_9049);
nand U11128 (N_11128,N_9552,N_9865);
xnor U11129 (N_11129,N_8833,N_9123);
nand U11130 (N_11130,N_9001,N_8775);
and U11131 (N_11131,N_8928,N_9886);
or U11132 (N_11132,N_9291,N_8822);
nand U11133 (N_11133,N_9119,N_9472);
or U11134 (N_11134,N_9834,N_9572);
xor U11135 (N_11135,N_9271,N_9301);
or U11136 (N_11136,N_9026,N_9955);
xor U11137 (N_11137,N_9713,N_9566);
xnor U11138 (N_11138,N_9737,N_9901);
nand U11139 (N_11139,N_9357,N_9976);
nor U11140 (N_11140,N_9637,N_9099);
xor U11141 (N_11141,N_9086,N_8975);
xor U11142 (N_11142,N_9957,N_9794);
xor U11143 (N_11143,N_9204,N_9730);
xnor U11144 (N_11144,N_9469,N_9286);
xnor U11145 (N_11145,N_9455,N_9936);
nor U11146 (N_11146,N_9590,N_9317);
and U11147 (N_11147,N_9382,N_9544);
or U11148 (N_11148,N_8995,N_9668);
and U11149 (N_11149,N_8787,N_9739);
or U11150 (N_11150,N_9221,N_9143);
and U11151 (N_11151,N_9308,N_9119);
nor U11152 (N_11152,N_9341,N_9212);
and U11153 (N_11153,N_8954,N_9448);
xnor U11154 (N_11154,N_8913,N_9575);
nand U11155 (N_11155,N_9880,N_9796);
or U11156 (N_11156,N_8998,N_9288);
xnor U11157 (N_11157,N_9512,N_8788);
or U11158 (N_11158,N_8762,N_9555);
or U11159 (N_11159,N_9827,N_9854);
xor U11160 (N_11160,N_9241,N_9417);
xnor U11161 (N_11161,N_9199,N_9756);
xor U11162 (N_11162,N_9038,N_9940);
nor U11163 (N_11163,N_9056,N_9562);
or U11164 (N_11164,N_9855,N_9229);
nand U11165 (N_11165,N_9703,N_9212);
xor U11166 (N_11166,N_9027,N_9788);
and U11167 (N_11167,N_9863,N_9268);
or U11168 (N_11168,N_9030,N_9989);
xnor U11169 (N_11169,N_9788,N_9272);
xnor U11170 (N_11170,N_9641,N_9585);
xnor U11171 (N_11171,N_9195,N_8800);
and U11172 (N_11172,N_9690,N_9092);
and U11173 (N_11173,N_9587,N_9600);
and U11174 (N_11174,N_8752,N_9342);
nor U11175 (N_11175,N_9093,N_9927);
xnor U11176 (N_11176,N_9560,N_9941);
or U11177 (N_11177,N_9709,N_9932);
or U11178 (N_11178,N_9935,N_9496);
nor U11179 (N_11179,N_9910,N_9428);
and U11180 (N_11180,N_9833,N_8921);
nor U11181 (N_11181,N_9885,N_9958);
and U11182 (N_11182,N_8825,N_9767);
and U11183 (N_11183,N_9572,N_8898);
or U11184 (N_11184,N_9651,N_9166);
xnor U11185 (N_11185,N_9945,N_9312);
nor U11186 (N_11186,N_9780,N_9178);
xnor U11187 (N_11187,N_9992,N_9533);
and U11188 (N_11188,N_9017,N_9619);
xor U11189 (N_11189,N_9946,N_9412);
nor U11190 (N_11190,N_9193,N_9299);
xnor U11191 (N_11191,N_9344,N_9768);
xor U11192 (N_11192,N_9682,N_9559);
nand U11193 (N_11193,N_9995,N_9402);
xnor U11194 (N_11194,N_9575,N_9131);
nor U11195 (N_11195,N_8888,N_9105);
nand U11196 (N_11196,N_9247,N_9922);
nor U11197 (N_11197,N_9408,N_9766);
nor U11198 (N_11198,N_8828,N_8950);
and U11199 (N_11199,N_9741,N_9261);
xnor U11200 (N_11200,N_9571,N_8845);
and U11201 (N_11201,N_9754,N_9109);
nor U11202 (N_11202,N_9253,N_9490);
or U11203 (N_11203,N_8985,N_8965);
and U11204 (N_11204,N_9356,N_9249);
nand U11205 (N_11205,N_9523,N_9737);
nor U11206 (N_11206,N_9288,N_9940);
xnor U11207 (N_11207,N_9069,N_9967);
and U11208 (N_11208,N_9113,N_8929);
and U11209 (N_11209,N_9095,N_8754);
and U11210 (N_11210,N_9312,N_9634);
or U11211 (N_11211,N_9421,N_9949);
nor U11212 (N_11212,N_9574,N_9610);
nor U11213 (N_11213,N_9171,N_9863);
xnor U11214 (N_11214,N_9175,N_9029);
nand U11215 (N_11215,N_8920,N_8976);
nor U11216 (N_11216,N_9033,N_9836);
or U11217 (N_11217,N_9788,N_9235);
or U11218 (N_11218,N_9292,N_8784);
or U11219 (N_11219,N_9861,N_9804);
xnor U11220 (N_11220,N_8876,N_9267);
and U11221 (N_11221,N_9198,N_9916);
nand U11222 (N_11222,N_9761,N_9277);
or U11223 (N_11223,N_9023,N_9728);
xor U11224 (N_11224,N_8807,N_9589);
xor U11225 (N_11225,N_9702,N_9760);
nand U11226 (N_11226,N_9572,N_9810);
and U11227 (N_11227,N_9958,N_9466);
nand U11228 (N_11228,N_9849,N_9357);
nor U11229 (N_11229,N_9808,N_9264);
nor U11230 (N_11230,N_9614,N_9523);
nor U11231 (N_11231,N_8869,N_9810);
and U11232 (N_11232,N_9525,N_9231);
nor U11233 (N_11233,N_9789,N_8954);
nand U11234 (N_11234,N_9184,N_9768);
or U11235 (N_11235,N_9894,N_9491);
xor U11236 (N_11236,N_8958,N_9979);
xnor U11237 (N_11237,N_9756,N_9333);
and U11238 (N_11238,N_9889,N_9843);
nor U11239 (N_11239,N_9640,N_9933);
or U11240 (N_11240,N_9057,N_8930);
nand U11241 (N_11241,N_9016,N_9023);
xnor U11242 (N_11242,N_9816,N_9566);
xnor U11243 (N_11243,N_9216,N_9560);
or U11244 (N_11244,N_9924,N_9969);
nand U11245 (N_11245,N_9923,N_9930);
xnor U11246 (N_11246,N_9326,N_8999);
xor U11247 (N_11247,N_9665,N_9914);
xnor U11248 (N_11248,N_9429,N_9047);
and U11249 (N_11249,N_9301,N_8807);
nor U11250 (N_11250,N_10241,N_10084);
and U11251 (N_11251,N_10096,N_10928);
xor U11252 (N_11252,N_10612,N_11177);
and U11253 (N_11253,N_10193,N_10757);
nand U11254 (N_11254,N_10208,N_10499);
nand U11255 (N_11255,N_10798,N_10466);
or U11256 (N_11256,N_10300,N_10401);
nor U11257 (N_11257,N_10664,N_10232);
nand U11258 (N_11258,N_10908,N_10873);
or U11259 (N_11259,N_10441,N_10089);
nand U11260 (N_11260,N_11025,N_11202);
and U11261 (N_11261,N_11149,N_10942);
nand U11262 (N_11262,N_10633,N_10091);
xnor U11263 (N_11263,N_10440,N_10897);
nand U11264 (N_11264,N_10352,N_10429);
xor U11265 (N_11265,N_10880,N_10251);
nor U11266 (N_11266,N_10181,N_10587);
xor U11267 (N_11267,N_11018,N_10981);
or U11268 (N_11268,N_10222,N_10107);
and U11269 (N_11269,N_10801,N_10565);
and U11270 (N_11270,N_10226,N_10504);
xnor U11271 (N_11271,N_10087,N_10487);
nor U11272 (N_11272,N_10535,N_11020);
xnor U11273 (N_11273,N_10468,N_11185);
and U11274 (N_11274,N_10436,N_10849);
nor U11275 (N_11275,N_10263,N_10304);
nand U11276 (N_11276,N_10442,N_10407);
xnor U11277 (N_11277,N_10695,N_11138);
or U11278 (N_11278,N_11012,N_10256);
and U11279 (N_11279,N_10116,N_10771);
xor U11280 (N_11280,N_10839,N_11193);
xor U11281 (N_11281,N_10496,N_10000);
nand U11282 (N_11282,N_11087,N_11118);
or U11283 (N_11283,N_10493,N_10976);
or U11284 (N_11284,N_10891,N_11186);
xor U11285 (N_11285,N_10437,N_10604);
nor U11286 (N_11286,N_11192,N_11155);
xnor U11287 (N_11287,N_11044,N_10481);
nand U11288 (N_11288,N_11211,N_11077);
nor U11289 (N_11289,N_10531,N_10592);
nand U11290 (N_11290,N_11230,N_10172);
and U11291 (N_11291,N_11246,N_10915);
xnor U11292 (N_11292,N_10058,N_10563);
xnor U11293 (N_11293,N_11204,N_10174);
nand U11294 (N_11294,N_10934,N_10858);
and U11295 (N_11295,N_10713,N_10862);
or U11296 (N_11296,N_10344,N_10660);
or U11297 (N_11297,N_10259,N_10417);
and U11298 (N_11298,N_10744,N_10685);
or U11299 (N_11299,N_10818,N_11059);
and U11300 (N_11300,N_11161,N_10649);
and U11301 (N_11301,N_10912,N_10902);
and U11302 (N_11302,N_10761,N_10180);
nor U11303 (N_11303,N_10541,N_10234);
xnor U11304 (N_11304,N_10213,N_11124);
xor U11305 (N_11305,N_10638,N_10829);
nor U11306 (N_11306,N_10736,N_10384);
nor U11307 (N_11307,N_10475,N_11234);
nor U11308 (N_11308,N_10673,N_10528);
nor U11309 (N_11309,N_11136,N_10192);
nor U11310 (N_11310,N_10701,N_10783);
xor U11311 (N_11311,N_11047,N_10999);
nor U11312 (N_11312,N_10539,N_10828);
nand U11313 (N_11313,N_10388,N_10435);
xor U11314 (N_11314,N_11003,N_10517);
and U11315 (N_11315,N_11141,N_10859);
or U11316 (N_11316,N_10372,N_10663);
xor U11317 (N_11317,N_10167,N_10467);
or U11318 (N_11318,N_11001,N_11152);
and U11319 (N_11319,N_10892,N_10692);
or U11320 (N_11320,N_10038,N_10671);
nor U11321 (N_11321,N_10670,N_11144);
or U11322 (N_11322,N_10317,N_10510);
and U11323 (N_11323,N_10291,N_10484);
and U11324 (N_11324,N_10595,N_10963);
or U11325 (N_11325,N_10720,N_10139);
nor U11326 (N_11326,N_10187,N_10398);
nor U11327 (N_11327,N_11052,N_10060);
or U11328 (N_11328,N_10746,N_11080);
or U11329 (N_11329,N_10723,N_10681);
xor U11330 (N_11330,N_10877,N_10586);
and U11331 (N_11331,N_10396,N_10944);
or U11332 (N_11332,N_10933,N_10762);
xnor U11333 (N_11333,N_10556,N_10279);
nor U11334 (N_11334,N_10888,N_10056);
or U11335 (N_11335,N_10792,N_10733);
nor U11336 (N_11336,N_10766,N_10257);
or U11337 (N_11337,N_10355,N_10110);
or U11338 (N_11338,N_10814,N_10628);
or U11339 (N_11339,N_10566,N_10969);
nor U11340 (N_11340,N_10412,N_10486);
and U11341 (N_11341,N_10893,N_10753);
and U11342 (N_11342,N_10986,N_11169);
nand U11343 (N_11343,N_10315,N_10739);
nor U11344 (N_11344,N_11109,N_10408);
nand U11345 (N_11345,N_10146,N_10325);
nand U11346 (N_11346,N_10579,N_11183);
nor U11347 (N_11347,N_11135,N_10306);
and U11348 (N_11348,N_10597,N_10201);
xnor U11349 (N_11349,N_10299,N_10223);
and U11350 (N_11350,N_10458,N_10190);
and U11351 (N_11351,N_10086,N_10006);
and U11352 (N_11352,N_10572,N_10918);
nor U11353 (N_11353,N_10947,N_10104);
xor U11354 (N_11354,N_11039,N_10361);
nor U11355 (N_11355,N_10972,N_10735);
and U11356 (N_11356,N_10952,N_11134);
nor U11357 (N_11357,N_10549,N_10785);
and U11358 (N_11358,N_10769,N_10029);
xor U11359 (N_11359,N_10802,N_10793);
and U11360 (N_11360,N_10422,N_10666);
and U11361 (N_11361,N_10092,N_10101);
nor U11362 (N_11362,N_10163,N_10812);
or U11363 (N_11363,N_10327,N_10932);
nor U11364 (N_11364,N_10634,N_10654);
xor U11365 (N_11365,N_10980,N_10030);
nor U11366 (N_11366,N_10079,N_10069);
xor U11367 (N_11367,N_10901,N_11235);
nor U11368 (N_11368,N_10109,N_10474);
xnor U11369 (N_11369,N_10519,N_11239);
xor U11370 (N_11370,N_11198,N_11166);
xor U11371 (N_11371,N_10584,N_10909);
nor U11372 (N_11372,N_10018,N_11164);
xor U11373 (N_11373,N_10874,N_10276);
nand U11374 (N_11374,N_10249,N_10825);
and U11375 (N_11375,N_10805,N_10293);
nor U11376 (N_11376,N_11036,N_11181);
nor U11377 (N_11377,N_10062,N_10377);
xnor U11378 (N_11378,N_11244,N_10882);
xnor U11379 (N_11379,N_10009,N_10042);
or U11380 (N_11380,N_10378,N_10130);
nor U11381 (N_11381,N_10289,N_10227);
or U11382 (N_11382,N_10358,N_11098);
nand U11383 (N_11383,N_10143,N_10215);
xor U11384 (N_11384,N_10323,N_10285);
xor U11385 (N_11385,N_10710,N_10497);
nor U11386 (N_11386,N_10609,N_10832);
and U11387 (N_11387,N_10400,N_10658);
or U11388 (N_11388,N_11088,N_10644);
or U11389 (N_11389,N_11129,N_10640);
xor U11390 (N_11390,N_10748,N_10477);
xnor U11391 (N_11391,N_10051,N_11053);
and U11392 (N_11392,N_10948,N_10480);
nand U11393 (N_11393,N_10583,N_11043);
xor U11394 (N_11394,N_10900,N_10758);
and U11395 (N_11395,N_11106,N_10406);
xor U11396 (N_11396,N_10575,N_10749);
xnor U11397 (N_11397,N_10320,N_10191);
nand U11398 (N_11398,N_10262,N_10790);
nand U11399 (N_11399,N_10730,N_10610);
nor U11400 (N_11400,N_10068,N_11223);
nor U11401 (N_11401,N_11127,N_11048);
or U11402 (N_11402,N_10033,N_11123);
nand U11403 (N_11403,N_10444,N_10558);
nand U11404 (N_11404,N_11160,N_10830);
xnor U11405 (N_11405,N_10864,N_10596);
and U11406 (N_11406,N_11242,N_11222);
or U11407 (N_11407,N_10472,N_10155);
xor U11408 (N_11408,N_10703,N_10287);
and U11409 (N_11409,N_10426,N_10799);
or U11410 (N_11410,N_10534,N_10652);
xnor U11411 (N_11411,N_11147,N_10581);
or U11412 (N_11412,N_10278,N_10984);
xor U11413 (N_11413,N_10153,N_10374);
and U11414 (N_11414,N_10211,N_10935);
nor U11415 (N_11415,N_10837,N_11099);
nand U11416 (N_11416,N_10445,N_10979);
and U11417 (N_11417,N_10356,N_10577);
xnor U11418 (N_11418,N_10381,N_10571);
and U11419 (N_11419,N_11221,N_10376);
and U11420 (N_11420,N_11030,N_10602);
nand U11421 (N_11421,N_10423,N_11095);
xor U11422 (N_11422,N_10359,N_11035);
nand U11423 (N_11423,N_11125,N_11197);
nor U11424 (N_11424,N_10696,N_11157);
or U11425 (N_11425,N_11076,N_10831);
or U11426 (N_11426,N_10275,N_11074);
xnor U11427 (N_11427,N_11031,N_10686);
xor U11428 (N_11428,N_11007,N_10639);
nand U11429 (N_11429,N_10419,N_10144);
nor U11430 (N_11430,N_10931,N_10889);
xnor U11431 (N_11431,N_10264,N_11010);
xnor U11432 (N_11432,N_10760,N_10387);
or U11433 (N_11433,N_10844,N_11100);
nand U11434 (N_11434,N_10258,N_10751);
nor U11435 (N_11435,N_10464,N_11201);
nand U11436 (N_11436,N_10626,N_10250);
nor U11437 (N_11437,N_10283,N_10495);
nand U11438 (N_11438,N_11180,N_10509);
nor U11439 (N_11439,N_10796,N_10034);
nand U11440 (N_11440,N_10741,N_10854);
nor U11441 (N_11441,N_10951,N_10724);
and U11442 (N_11442,N_10763,N_10850);
and U11443 (N_11443,N_10290,N_10852);
and U11444 (N_11444,N_11014,N_10272);
or U11445 (N_11445,N_10483,N_10759);
nor U11446 (N_11446,N_10819,N_10917);
and U11447 (N_11447,N_10871,N_11112);
or U11448 (N_11448,N_11119,N_11082);
and U11449 (N_11449,N_10151,N_10808);
or U11450 (N_11450,N_10675,N_10329);
nand U11451 (N_11451,N_10603,N_11050);
or U11452 (N_11452,N_10843,N_10453);
xnor U11453 (N_11453,N_10059,N_10813);
or U11454 (N_11454,N_11062,N_10625);
and U11455 (N_11455,N_11196,N_10856);
and U11456 (N_11456,N_10156,N_10840);
and U11457 (N_11457,N_10364,N_10745);
nand U11458 (N_11458,N_10238,N_10938);
or U11459 (N_11459,N_11115,N_10732);
xnor U11460 (N_11460,N_11200,N_10053);
nand U11461 (N_11461,N_10463,N_10836);
nor U11462 (N_11462,N_10807,N_11143);
nand U11463 (N_11463,N_10775,N_11203);
or U11464 (N_11464,N_11154,N_10946);
nand U11465 (N_11465,N_10788,N_11175);
nor U11466 (N_11466,N_10131,N_10017);
and U11467 (N_11467,N_11116,N_10135);
nor U11468 (N_11468,N_10786,N_10270);
nand U11469 (N_11469,N_10594,N_11219);
xor U11470 (N_11470,N_10339,N_10218);
nor U11471 (N_11471,N_10321,N_10055);
nand U11472 (N_11472,N_10608,N_11008);
and U11473 (N_11473,N_10574,N_10505);
or U11474 (N_11474,N_10898,N_10080);
or U11475 (N_11475,N_10557,N_10379);
nor U11476 (N_11476,N_10997,N_10550);
and U11477 (N_11477,N_10421,N_10225);
nor U11478 (N_11478,N_10899,N_10476);
xnor U11479 (N_11479,N_10182,N_10943);
or U11480 (N_11480,N_11206,N_10386);
and U11481 (N_11481,N_10318,N_10026);
xnor U11482 (N_11482,N_10036,N_10173);
xor U11483 (N_11483,N_10473,N_10134);
and U11484 (N_11484,N_10129,N_11148);
nand U11485 (N_11485,N_10373,N_11041);
nand U11486 (N_11486,N_10067,N_10369);
or U11487 (N_11487,N_11170,N_10044);
xnor U11488 (N_11488,N_10605,N_11055);
nor U11489 (N_11489,N_10567,N_10185);
nand U11490 (N_11490,N_10688,N_11113);
or U11491 (N_11491,N_10288,N_10332);
or U11492 (N_11492,N_10842,N_10545);
nand U11493 (N_11493,N_10661,N_10085);
and U11494 (N_11494,N_10623,N_10168);
nand U11495 (N_11495,N_11225,N_11209);
xnor U11496 (N_11496,N_11199,N_10806);
nand U11497 (N_11497,N_10368,N_10590);
nor U11498 (N_11498,N_11060,N_11248);
or U11499 (N_11499,N_10301,N_11179);
or U11500 (N_11500,N_10667,N_10341);
xnor U11501 (N_11501,N_10731,N_10770);
nor U11502 (N_11502,N_10618,N_10169);
and U11503 (N_11503,N_10237,N_10452);
nor U11504 (N_11504,N_10553,N_10456);
and U11505 (N_11505,N_10929,N_10491);
and U11506 (N_11506,N_10455,N_11061);
xor U11507 (N_11507,N_10274,N_11006);
or U11508 (N_11508,N_10221,N_10552);
nor U11509 (N_11509,N_10811,N_10012);
nor U11510 (N_11510,N_10410,N_11187);
and U11511 (N_11511,N_10296,N_11151);
nor U11512 (N_11512,N_11069,N_10525);
or U11513 (N_11513,N_11224,N_11058);
and U11514 (N_11514,N_10375,N_10971);
xor U11515 (N_11515,N_10261,N_10527);
and U11516 (N_11516,N_10013,N_10048);
xor U11517 (N_11517,N_10451,N_11086);
nor U11518 (N_11518,N_10702,N_11146);
or U11519 (N_11519,N_10657,N_10869);
xor U11520 (N_11520,N_10564,N_10360);
or U11521 (N_11521,N_10157,N_10896);
or U11522 (N_11522,N_10125,N_10175);
xnor U11523 (N_11523,N_11184,N_10668);
and U11524 (N_11524,N_10551,N_10975);
or U11525 (N_11525,N_10342,N_10209);
or U11526 (N_11526,N_10106,N_10651);
xor U11527 (N_11527,N_10548,N_10680);
xnor U11528 (N_11528,N_10367,N_10511);
nand U11529 (N_11529,N_10070,N_10432);
xnor U11530 (N_11530,N_10292,N_10127);
nor U11531 (N_11531,N_10028,N_10524);
nor U11532 (N_11532,N_11017,N_10032);
or U11533 (N_11533,N_10016,N_10921);
nand U11534 (N_11534,N_10507,N_10057);
or U11535 (N_11535,N_11212,N_11101);
xor U11536 (N_11536,N_11172,N_10500);
xor U11537 (N_11537,N_10489,N_10962);
xor U11538 (N_11538,N_10365,N_10239);
xor U11539 (N_11539,N_11153,N_10073);
or U11540 (N_11540,N_10188,N_10336);
or U11541 (N_11541,N_10202,N_10041);
or U11542 (N_11542,N_10987,N_11238);
nand U11543 (N_11543,N_10968,N_10004);
and U11544 (N_11544,N_11140,N_10331);
nor U11545 (N_11545,N_10810,N_11033);
or U11546 (N_11546,N_10046,N_11178);
and U11547 (N_11547,N_10789,N_11057);
nor U11548 (N_11548,N_10189,N_10719);
and U11549 (N_11549,N_10704,N_11207);
nand U11550 (N_11550,N_10648,N_10210);
nand U11551 (N_11551,N_10878,N_10447);
nand U11552 (N_11552,N_10161,N_11091);
nand U11553 (N_11553,N_10308,N_10415);
nor U11554 (N_11554,N_10521,N_10820);
and U11555 (N_11555,N_11173,N_10413);
or U11556 (N_11556,N_10978,N_10983);
or U11557 (N_11557,N_10956,N_10311);
nand U11558 (N_11558,N_10449,N_10752);
nor U11559 (N_11559,N_10727,N_10093);
xnor U11560 (N_11560,N_10284,N_10111);
nand U11561 (N_11561,N_10217,N_10309);
nand U11562 (N_11562,N_11015,N_11188);
nor U11563 (N_11563,N_10076,N_10351);
or U11564 (N_11564,N_10536,N_10243);
xor U11565 (N_11565,N_10996,N_10868);
xnor U11566 (N_11566,N_10676,N_10606);
nand U11567 (N_11567,N_10848,N_11073);
xnor U11568 (N_11568,N_11215,N_10522);
xor U11569 (N_11569,N_10298,N_10782);
and U11570 (N_11570,N_10949,N_11210);
or U11571 (N_11571,N_10199,N_11167);
nor U11572 (N_11572,N_10443,N_10098);
xor U11573 (N_11573,N_10402,N_10506);
nor U11574 (N_11574,N_10324,N_11027);
nor U11575 (N_11575,N_11105,N_10371);
nand U11576 (N_11576,N_11108,N_11132);
xor U11577 (N_11577,N_10824,N_10863);
nand U11578 (N_11578,N_10991,N_10177);
and U11579 (N_11579,N_10973,N_10136);
or U11580 (N_11580,N_10303,N_10020);
and U11581 (N_11581,N_11065,N_11032);
nand U11582 (N_11582,N_10273,N_10112);
xor U11583 (N_11583,N_10872,N_11046);
xnor U11584 (N_11584,N_10128,N_10392);
nand U11585 (N_11585,N_10043,N_10039);
and U11586 (N_11586,N_10122,N_10431);
or U11587 (N_11587,N_10940,N_11159);
nand U11588 (N_11588,N_10726,N_10071);
xnor U11589 (N_11589,N_10390,N_10974);
nand U11590 (N_11590,N_10490,N_10265);
nor U11591 (N_11591,N_10659,N_11038);
xor U11592 (N_11592,N_11195,N_10001);
and U11593 (N_11593,N_10767,N_10765);
or U11594 (N_11594,N_10152,N_10939);
xnor U11595 (N_11595,N_10936,N_10523);
and U11596 (N_11596,N_11208,N_11023);
or U11597 (N_11597,N_10773,N_10526);
nor U11598 (N_11598,N_10920,N_10229);
xor U11599 (N_11599,N_10682,N_10047);
nand U11600 (N_11600,N_10121,N_10513);
xor U11601 (N_11601,N_11162,N_10988);
xnor U11602 (N_11602,N_10886,N_10160);
nor U11603 (N_11603,N_10340,N_10236);
or U11604 (N_11604,N_10772,N_10691);
or U11605 (N_11605,N_11121,N_11227);
xor U11606 (N_11606,N_10008,N_10835);
xnor U11607 (N_11607,N_10197,N_11231);
xnor U11608 (N_11608,N_10865,N_10138);
or U11609 (N_11609,N_10147,N_10591);
nor U11610 (N_11610,N_10573,N_11243);
xor U11611 (N_11611,N_10077,N_10543);
or U11612 (N_11612,N_10240,N_10314);
nand U11613 (N_11613,N_10794,N_11075);
and U11614 (N_11614,N_11176,N_10363);
xor U11615 (N_11615,N_10580,N_10970);
xor U11616 (N_11616,N_10914,N_10598);
and U11617 (N_11617,N_10647,N_11037);
and U11618 (N_11618,N_11114,N_10740);
nand U11619 (N_11619,N_11220,N_10281);
and U11620 (N_11620,N_10994,N_10471);
xor U11621 (N_11621,N_11205,N_10697);
xor U11622 (N_11622,N_10957,N_10665);
xor U11623 (N_11623,N_11110,N_11103);
nand U11624 (N_11624,N_11079,N_10890);
nand U11625 (N_11625,N_10601,N_10065);
nand U11626 (N_11626,N_11232,N_10853);
xor U11627 (N_11627,N_10540,N_10738);
or U11628 (N_11628,N_10699,N_10833);
xor U11629 (N_11629,N_10637,N_10313);
nor U11630 (N_11630,N_10672,N_10502);
or U11631 (N_11631,N_10460,N_11016);
xnor U11632 (N_11632,N_10319,N_10613);
nor U11633 (N_11633,N_10022,N_10958);
and U11634 (N_11634,N_10170,N_11247);
nor U11635 (N_11635,N_10630,N_10282);
xnor U11636 (N_11636,N_10679,N_11150);
nand U11637 (N_11637,N_11042,N_10636);
nand U11638 (N_11638,N_10108,N_10774);
nor U11639 (N_11639,N_10887,N_10930);
and U11640 (N_11640,N_10870,N_11011);
nor U11641 (N_11641,N_10570,N_10684);
nor U11642 (N_11642,N_10937,N_10641);
xor U11643 (N_11643,N_10516,N_10409);
nand U11644 (N_11644,N_10049,N_10158);
xor U11645 (N_11645,N_10926,N_10267);
or U11646 (N_11646,N_10478,N_11171);
nand U11647 (N_11647,N_10438,N_10924);
or U11648 (N_11648,N_10544,N_10002);
and U11649 (N_11649,N_10411,N_10955);
nand U11650 (N_11650,N_10063,N_11051);
and U11651 (N_11651,N_10380,N_10066);
xnor U11652 (N_11652,N_11090,N_10714);
nand U11653 (N_11653,N_11245,N_10297);
nand U11654 (N_11654,N_10224,N_10354);
or U11655 (N_11655,N_10366,N_10800);
xnor U11656 (N_11656,N_10459,N_10183);
or U11657 (N_11657,N_10120,N_10847);
nor U11658 (N_11658,N_10922,N_10866);
nor U11659 (N_11659,N_10252,N_11104);
or U11660 (N_11660,N_10503,N_11156);
nand U11661 (N_11661,N_10050,N_11093);
nand U11662 (N_11662,N_10150,N_11189);
nor U11663 (N_11663,N_10635,N_10919);
and U11664 (N_11664,N_11249,N_11111);
or U11665 (N_11665,N_10662,N_10074);
or U11666 (N_11666,N_10142,N_11094);
xnor U11667 (N_11667,N_10742,N_10599);
or U11668 (N_11668,N_10576,N_10725);
xor U11669 (N_11669,N_11218,N_11045);
xor U11670 (N_11670,N_10328,N_10821);
or U11671 (N_11671,N_11102,N_10383);
or U11672 (N_11672,N_10778,N_10841);
and U11673 (N_11673,N_11064,N_11190);
xnor U11674 (N_11674,N_10014,N_10561);
xnor U11675 (N_11675,N_10619,N_10405);
and U11676 (N_11676,N_11165,N_10011);
xor U11677 (N_11677,N_11107,N_10809);
nand U11678 (N_11678,N_10655,N_10622);
nor U11679 (N_11679,N_10428,N_10953);
and U11680 (N_11680,N_10734,N_11028);
xnor U11681 (N_11681,N_10656,N_10706);
and U11682 (N_11682,N_10391,N_10764);
xnor U11683 (N_11683,N_10728,N_11026);
and U11684 (N_11684,N_10488,N_10966);
nand U11685 (N_11685,N_11226,N_10322);
or U11686 (N_11686,N_10399,N_10345);
or U11687 (N_11687,N_10537,N_10271);
xor U11688 (N_11688,N_10233,N_10216);
xor U11689 (N_11689,N_10479,N_10950);
or U11690 (N_11690,N_11096,N_10616);
nand U11691 (N_11691,N_10439,N_10582);
nand U11692 (N_11692,N_10708,N_10141);
xor U11693 (N_11693,N_10834,N_10268);
xnor U11694 (N_11694,N_10119,N_10925);
xnor U11695 (N_11695,N_10588,N_10876);
and U11696 (N_11696,N_10905,N_10709);
xor U11697 (N_11697,N_10054,N_10389);
nand U11698 (N_11698,N_10114,N_10492);
and U11699 (N_11699,N_10260,N_10993);
nand U11700 (N_11700,N_10040,N_10784);
xnor U11701 (N_11701,N_10838,N_10214);
or U11702 (N_11702,N_11097,N_10425);
and U11703 (N_11703,N_10916,N_11145);
nor U11704 (N_11704,N_10307,N_10154);
and U11705 (N_11705,N_10515,N_10027);
and U11706 (N_11706,N_11214,N_10791);
and U11707 (N_11707,N_11126,N_10338);
xor U11708 (N_11708,N_10310,N_10985);
or U11709 (N_11709,N_10397,N_10021);
or U11710 (N_11710,N_10712,N_10508);
nand U11711 (N_11711,N_10721,N_10910);
xnor U11712 (N_11712,N_11019,N_11128);
xnor U11713 (N_11713,N_10906,N_10090);
xnor U11714 (N_11714,N_10514,N_10642);
xor U11715 (N_11715,N_10061,N_10795);
nand U11716 (N_11716,N_10815,N_10382);
xor U11717 (N_11717,N_10879,N_10266);
xnor U11718 (N_11718,N_11002,N_10248);
nor U11719 (N_11719,N_10927,N_10099);
nand U11720 (N_11720,N_10904,N_10617);
or U11721 (N_11721,N_11217,N_10857);
nor U11722 (N_11722,N_11131,N_10532);
or U11723 (N_11723,N_10007,N_11067);
nor U11724 (N_11724,N_10694,N_10242);
nand U11725 (N_11725,N_10015,N_10228);
xor U11726 (N_11726,N_10755,N_10600);
nor U11727 (N_11727,N_10420,N_10149);
xor U11728 (N_11728,N_11241,N_11191);
and U11729 (N_11729,N_10578,N_10530);
xnor U11730 (N_11730,N_10964,N_10822);
nor U11731 (N_11731,N_11092,N_10195);
nor U11732 (N_11732,N_10780,N_10498);
or U11733 (N_11733,N_10117,N_10416);
and U11734 (N_11734,N_10031,N_10094);
nand U11735 (N_11735,N_11004,N_10088);
xnor U11736 (N_11736,N_10255,N_10959);
nor U11737 (N_11737,N_10559,N_10620);
and U11738 (N_11738,N_10393,N_10343);
nand U11739 (N_11739,N_10961,N_10333);
xnor U11740 (N_11740,N_10294,N_10967);
or U11741 (N_11741,N_11009,N_10203);
nand U11742 (N_11742,N_10023,N_11029);
or U11743 (N_11743,N_10097,N_10204);
nor U11744 (N_11744,N_11120,N_11085);
nand U11745 (N_11745,N_10145,N_10518);
nor U11746 (N_11746,N_10219,N_10632);
or U11747 (N_11747,N_10166,N_10722);
xor U11748 (N_11748,N_10019,N_10176);
nand U11749 (N_11749,N_10072,N_11078);
and U11750 (N_11750,N_10454,N_10277);
or U11751 (N_11751,N_10280,N_10171);
or U11752 (N_11752,N_10716,N_11024);
nand U11753 (N_11753,N_10082,N_10103);
xnor U11754 (N_11754,N_10433,N_11142);
nand U11755 (N_11755,N_10430,N_10747);
nor U11756 (N_11756,N_10178,N_10253);
nand U11757 (N_11757,N_11034,N_10105);
and U11758 (N_11758,N_10132,N_10235);
or U11759 (N_11759,N_10353,N_10164);
nor U11760 (N_11760,N_10945,N_11063);
nor U11761 (N_11761,N_11182,N_10207);
nand U11762 (N_11762,N_10348,N_10200);
or U11763 (N_11763,N_10124,N_10003);
nor U11764 (N_11764,N_11158,N_10729);
xor U11765 (N_11765,N_10385,N_11083);
or U11766 (N_11766,N_10115,N_10700);
nor U11767 (N_11767,N_10705,N_10078);
and U11768 (N_11768,N_10562,N_10689);
or U11769 (N_11769,N_11229,N_10650);
xnor U11770 (N_11770,N_10881,N_10855);
nor U11771 (N_11771,N_10403,N_10718);
and U11772 (N_11772,N_10081,N_10424);
nand U11773 (N_11773,N_10555,N_10005);
or U11774 (N_11774,N_10037,N_10826);
and U11775 (N_11775,N_10095,N_11117);
nand U11776 (N_11776,N_10624,N_10394);
xor U11777 (N_11777,N_10941,N_10269);
nand U11778 (N_11778,N_11194,N_10469);
nand U11779 (N_11779,N_10295,N_10494);
xor U11780 (N_11780,N_10646,N_10585);
or U11781 (N_11781,N_10512,N_10247);
nand U11782 (N_11782,N_10024,N_11068);
nand U11783 (N_11783,N_11013,N_10804);
xnor U11784 (N_11784,N_10627,N_10075);
or U11785 (N_11785,N_10230,N_10614);
xnor U11786 (N_11786,N_10052,N_10643);
and U11787 (N_11787,N_10992,N_10414);
xnor U11788 (N_11788,N_10347,N_10885);
and U11789 (N_11789,N_11139,N_10687);
nand U11790 (N_11790,N_11054,N_11133);
nand U11791 (N_11791,N_10462,N_10350);
and U11792 (N_11792,N_10349,N_10448);
nand U11793 (N_11793,N_11228,N_10913);
xor U11794 (N_11794,N_11066,N_11072);
and U11795 (N_11795,N_10960,N_10894);
and U11796 (N_11796,N_10861,N_10186);
xor U11797 (N_11797,N_11040,N_11084);
nand U11798 (N_11798,N_10827,N_10148);
xnor U11799 (N_11799,N_10998,N_10777);
or U11800 (N_11800,N_10669,N_11240);
nor U11801 (N_11801,N_10743,N_10977);
or U11802 (N_11802,N_10045,N_10754);
and U11803 (N_11803,N_10823,N_10907);
xnor U11804 (N_11804,N_10254,N_10589);
xor U11805 (N_11805,N_10485,N_10446);
nand U11806 (N_11806,N_10846,N_10165);
and U11807 (N_11807,N_10787,N_10212);
xnor U11808 (N_11808,N_10334,N_10547);
and U11809 (N_11809,N_10860,N_11070);
nor U11810 (N_11810,N_10162,N_10717);
or U11811 (N_11811,N_10715,N_10615);
xnor U11812 (N_11812,N_10965,N_10010);
or U11813 (N_11813,N_10737,N_10501);
xor U11814 (N_11814,N_10246,N_10677);
and U11815 (N_11815,N_10100,N_10370);
xnor U11816 (N_11816,N_10690,N_11213);
nand U11817 (N_11817,N_10404,N_11216);
and U11818 (N_11818,N_10126,N_11071);
and U11819 (N_11819,N_10707,N_10337);
or U11820 (N_11820,N_10911,N_10330);
xor U11821 (N_11821,N_10803,N_10995);
xnor U11822 (N_11822,N_10923,N_10568);
and U11823 (N_11823,N_10990,N_10231);
nor U11824 (N_11824,N_10653,N_11237);
or U11825 (N_11825,N_10427,N_10845);
or U11826 (N_11826,N_10123,N_10118);
nor U11827 (N_11827,N_11174,N_11022);
nor U11828 (N_11828,N_10883,N_10554);
nand U11829 (N_11829,N_10159,N_11049);
nor U11830 (N_11830,N_10851,N_10631);
or U11831 (N_11831,N_10245,N_10779);
xor U11832 (N_11832,N_10621,N_10546);
and U11833 (N_11833,N_11021,N_10206);
or U11834 (N_11834,N_10674,N_11000);
nand U11835 (N_11835,N_10645,N_10244);
nor U11836 (N_11836,N_10542,N_10982);
nor U11837 (N_11837,N_10133,N_10768);
xnor U11838 (N_11838,N_10205,N_10750);
xnor U11839 (N_11839,N_10179,N_10693);
nor U11840 (N_11840,N_10989,N_10357);
or U11841 (N_11841,N_10312,N_11130);
and U11842 (N_11842,N_11089,N_10302);
nor U11843 (N_11843,N_10346,N_10470);
xor U11844 (N_11844,N_10678,N_10607);
or U11845 (N_11845,N_10533,N_10220);
and U11846 (N_11846,N_11056,N_10629);
nor U11847 (N_11847,N_10064,N_10875);
xnor U11848 (N_11848,N_10529,N_10611);
or U11849 (N_11849,N_10781,N_10035);
xnor U11850 (N_11850,N_10198,N_10395);
or U11851 (N_11851,N_10593,N_11137);
nand U11852 (N_11852,N_10194,N_10316);
nand U11853 (N_11853,N_10113,N_10461);
nor U11854 (N_11854,N_10326,N_10698);
nand U11855 (N_11855,N_10569,N_11081);
or U11856 (N_11856,N_10335,N_10137);
or U11857 (N_11857,N_11005,N_11163);
and U11858 (N_11858,N_10895,N_10196);
or U11859 (N_11859,N_10184,N_10817);
nand U11860 (N_11860,N_10286,N_10140);
or U11861 (N_11861,N_10520,N_11122);
and U11862 (N_11862,N_10797,N_11168);
and U11863 (N_11863,N_10305,N_11236);
xor U11864 (N_11864,N_10954,N_10884);
nand U11865 (N_11865,N_10362,N_10102);
nor U11866 (N_11866,N_10457,N_10776);
nor U11867 (N_11867,N_10816,N_10083);
nand U11868 (N_11868,N_10482,N_10465);
or U11869 (N_11869,N_10025,N_10711);
nand U11870 (N_11870,N_11233,N_10560);
xnor U11871 (N_11871,N_10450,N_10903);
nor U11872 (N_11872,N_10867,N_10538);
and U11873 (N_11873,N_10418,N_10434);
nor U11874 (N_11874,N_10756,N_10683);
nor U11875 (N_11875,N_10469,N_10575);
xor U11876 (N_11876,N_10169,N_11181);
nor U11877 (N_11877,N_10827,N_11219);
and U11878 (N_11878,N_11111,N_10254);
xnor U11879 (N_11879,N_10291,N_10714);
nand U11880 (N_11880,N_10626,N_10129);
or U11881 (N_11881,N_10867,N_10360);
or U11882 (N_11882,N_10326,N_10661);
nand U11883 (N_11883,N_10580,N_10386);
nor U11884 (N_11884,N_10898,N_11060);
nand U11885 (N_11885,N_10110,N_10672);
or U11886 (N_11886,N_10657,N_10876);
xor U11887 (N_11887,N_10515,N_10173);
xnor U11888 (N_11888,N_10704,N_10060);
and U11889 (N_11889,N_11017,N_10582);
nor U11890 (N_11890,N_10596,N_11145);
nand U11891 (N_11891,N_11017,N_10920);
nor U11892 (N_11892,N_10645,N_10722);
nor U11893 (N_11893,N_10483,N_10778);
nand U11894 (N_11894,N_10322,N_10346);
or U11895 (N_11895,N_10282,N_10300);
xnor U11896 (N_11896,N_10072,N_10619);
and U11897 (N_11897,N_10209,N_10689);
xnor U11898 (N_11898,N_10145,N_10871);
nor U11899 (N_11899,N_10926,N_10910);
nor U11900 (N_11900,N_10350,N_11124);
xor U11901 (N_11901,N_10086,N_10004);
nor U11902 (N_11902,N_10578,N_10843);
or U11903 (N_11903,N_10052,N_10202);
and U11904 (N_11904,N_11074,N_10175);
and U11905 (N_11905,N_11016,N_10068);
and U11906 (N_11906,N_10119,N_10890);
xnor U11907 (N_11907,N_10418,N_11103);
nor U11908 (N_11908,N_10153,N_10369);
xor U11909 (N_11909,N_11231,N_10053);
xnor U11910 (N_11910,N_10090,N_10766);
or U11911 (N_11911,N_10343,N_10318);
and U11912 (N_11912,N_10039,N_10253);
nand U11913 (N_11913,N_11218,N_10616);
nand U11914 (N_11914,N_10805,N_10485);
nand U11915 (N_11915,N_10701,N_10929);
nand U11916 (N_11916,N_11199,N_11177);
nand U11917 (N_11917,N_11242,N_10978);
or U11918 (N_11918,N_10016,N_10547);
or U11919 (N_11919,N_10375,N_11016);
nor U11920 (N_11920,N_10105,N_10138);
xnor U11921 (N_11921,N_10173,N_10644);
xnor U11922 (N_11922,N_11191,N_10900);
nor U11923 (N_11923,N_11219,N_10430);
nand U11924 (N_11924,N_10713,N_10499);
xnor U11925 (N_11925,N_10453,N_10401);
xor U11926 (N_11926,N_10347,N_10549);
and U11927 (N_11927,N_10786,N_11048);
nor U11928 (N_11928,N_10726,N_10123);
nor U11929 (N_11929,N_11074,N_10363);
nand U11930 (N_11930,N_10464,N_10588);
or U11931 (N_11931,N_10713,N_11204);
or U11932 (N_11932,N_10675,N_10844);
and U11933 (N_11933,N_10137,N_10063);
and U11934 (N_11934,N_10898,N_10715);
nor U11935 (N_11935,N_10483,N_10368);
or U11936 (N_11936,N_11132,N_10823);
nand U11937 (N_11937,N_10213,N_10549);
nor U11938 (N_11938,N_10749,N_10373);
and U11939 (N_11939,N_10632,N_11114);
or U11940 (N_11940,N_10108,N_10235);
nand U11941 (N_11941,N_10828,N_10541);
and U11942 (N_11942,N_10931,N_10936);
nor U11943 (N_11943,N_10664,N_10242);
nor U11944 (N_11944,N_10850,N_10539);
nor U11945 (N_11945,N_10626,N_10711);
xnor U11946 (N_11946,N_10970,N_10958);
nand U11947 (N_11947,N_10278,N_10424);
nand U11948 (N_11948,N_10502,N_10375);
nor U11949 (N_11949,N_11227,N_10884);
xnor U11950 (N_11950,N_10851,N_10638);
or U11951 (N_11951,N_11017,N_10679);
and U11952 (N_11952,N_10764,N_11129);
nor U11953 (N_11953,N_11072,N_10562);
xnor U11954 (N_11954,N_10632,N_10466);
xor U11955 (N_11955,N_10180,N_10152);
nand U11956 (N_11956,N_10530,N_10331);
nand U11957 (N_11957,N_10041,N_11039);
or U11958 (N_11958,N_10804,N_10632);
nand U11959 (N_11959,N_10558,N_11248);
xor U11960 (N_11960,N_10135,N_10175);
nor U11961 (N_11961,N_11078,N_10913);
and U11962 (N_11962,N_10959,N_10324);
xnor U11963 (N_11963,N_10666,N_11026);
and U11964 (N_11964,N_10921,N_10398);
and U11965 (N_11965,N_10064,N_10334);
nand U11966 (N_11966,N_10689,N_10044);
nand U11967 (N_11967,N_10845,N_10915);
nand U11968 (N_11968,N_10101,N_10175);
nand U11969 (N_11969,N_11180,N_10525);
or U11970 (N_11970,N_10518,N_10148);
nor U11971 (N_11971,N_10782,N_10775);
nor U11972 (N_11972,N_10749,N_10107);
xnor U11973 (N_11973,N_10088,N_10410);
nor U11974 (N_11974,N_10187,N_10077);
nor U11975 (N_11975,N_10431,N_10913);
xnor U11976 (N_11976,N_11244,N_10367);
nor U11977 (N_11977,N_10873,N_10077);
and U11978 (N_11978,N_11229,N_11019);
nor U11979 (N_11979,N_10233,N_11088);
or U11980 (N_11980,N_10767,N_11073);
or U11981 (N_11981,N_10010,N_10093);
xnor U11982 (N_11982,N_11144,N_10082);
xor U11983 (N_11983,N_10619,N_11146);
or U11984 (N_11984,N_11133,N_10707);
nor U11985 (N_11985,N_10987,N_10720);
or U11986 (N_11986,N_10256,N_10468);
xnor U11987 (N_11987,N_11245,N_10688);
nor U11988 (N_11988,N_10621,N_10056);
nor U11989 (N_11989,N_11124,N_10247);
xnor U11990 (N_11990,N_10159,N_10819);
xor U11991 (N_11991,N_10765,N_11073);
and U11992 (N_11992,N_10640,N_10602);
and U11993 (N_11993,N_11113,N_11138);
and U11994 (N_11994,N_10871,N_10573);
nor U11995 (N_11995,N_10181,N_10159);
xor U11996 (N_11996,N_10228,N_11093);
nor U11997 (N_11997,N_11101,N_10609);
xor U11998 (N_11998,N_11192,N_11103);
and U11999 (N_11999,N_11236,N_10408);
or U12000 (N_12000,N_10369,N_10499);
or U12001 (N_12001,N_10197,N_10151);
nand U12002 (N_12002,N_10147,N_10019);
and U12003 (N_12003,N_10988,N_10106);
nor U12004 (N_12004,N_10307,N_10497);
nor U12005 (N_12005,N_11107,N_10864);
xor U12006 (N_12006,N_10292,N_10858);
and U12007 (N_12007,N_10454,N_10086);
nor U12008 (N_12008,N_10737,N_10308);
nand U12009 (N_12009,N_10511,N_10557);
and U12010 (N_12010,N_10649,N_10217);
or U12011 (N_12011,N_10604,N_10047);
and U12012 (N_12012,N_10370,N_10267);
and U12013 (N_12013,N_10158,N_10997);
or U12014 (N_12014,N_11047,N_10363);
xor U12015 (N_12015,N_10036,N_10122);
or U12016 (N_12016,N_10337,N_11037);
and U12017 (N_12017,N_10134,N_10215);
or U12018 (N_12018,N_11075,N_10073);
nor U12019 (N_12019,N_10286,N_10744);
nand U12020 (N_12020,N_10477,N_10196);
or U12021 (N_12021,N_10195,N_10937);
and U12022 (N_12022,N_10970,N_10099);
xor U12023 (N_12023,N_10205,N_11174);
xnor U12024 (N_12024,N_11208,N_10395);
and U12025 (N_12025,N_11083,N_11146);
nor U12026 (N_12026,N_11187,N_10361);
nor U12027 (N_12027,N_10648,N_11083);
nor U12028 (N_12028,N_10792,N_10440);
nor U12029 (N_12029,N_10593,N_10667);
nand U12030 (N_12030,N_10704,N_10712);
xor U12031 (N_12031,N_10824,N_10241);
nand U12032 (N_12032,N_10384,N_10780);
xor U12033 (N_12033,N_11158,N_11071);
and U12034 (N_12034,N_10693,N_10985);
xor U12035 (N_12035,N_10879,N_10604);
nor U12036 (N_12036,N_10338,N_11193);
and U12037 (N_12037,N_10250,N_10162);
nor U12038 (N_12038,N_10860,N_10548);
and U12039 (N_12039,N_10629,N_10904);
nand U12040 (N_12040,N_10851,N_11157);
xnor U12041 (N_12041,N_10596,N_10964);
xor U12042 (N_12042,N_10628,N_10397);
xnor U12043 (N_12043,N_11141,N_10816);
nor U12044 (N_12044,N_10736,N_10441);
and U12045 (N_12045,N_10878,N_11119);
or U12046 (N_12046,N_10125,N_10168);
or U12047 (N_12047,N_11162,N_10080);
or U12048 (N_12048,N_10784,N_10324);
xnor U12049 (N_12049,N_10710,N_10342);
xor U12050 (N_12050,N_10171,N_10644);
xor U12051 (N_12051,N_10297,N_10270);
nor U12052 (N_12052,N_10078,N_10207);
or U12053 (N_12053,N_10709,N_10676);
xnor U12054 (N_12054,N_11186,N_10775);
xnor U12055 (N_12055,N_11075,N_10950);
nor U12056 (N_12056,N_10825,N_10181);
nand U12057 (N_12057,N_10305,N_11096);
and U12058 (N_12058,N_10741,N_10817);
or U12059 (N_12059,N_10461,N_10988);
xor U12060 (N_12060,N_11038,N_10560);
nand U12061 (N_12061,N_10470,N_10530);
or U12062 (N_12062,N_10604,N_11146);
nand U12063 (N_12063,N_11182,N_10038);
or U12064 (N_12064,N_11199,N_10892);
and U12065 (N_12065,N_10346,N_10338);
nand U12066 (N_12066,N_11004,N_11134);
or U12067 (N_12067,N_11101,N_11002);
nand U12068 (N_12068,N_11094,N_10307);
xnor U12069 (N_12069,N_10304,N_11239);
and U12070 (N_12070,N_10352,N_10094);
xor U12071 (N_12071,N_10761,N_10105);
or U12072 (N_12072,N_10921,N_11222);
or U12073 (N_12073,N_10015,N_11217);
or U12074 (N_12074,N_10182,N_10704);
xor U12075 (N_12075,N_10905,N_10648);
xor U12076 (N_12076,N_10442,N_10026);
nor U12077 (N_12077,N_10238,N_10175);
or U12078 (N_12078,N_10622,N_10595);
and U12079 (N_12079,N_10451,N_10905);
nor U12080 (N_12080,N_10609,N_10389);
nor U12081 (N_12081,N_11143,N_11131);
xor U12082 (N_12082,N_10873,N_10379);
xnor U12083 (N_12083,N_10766,N_10184);
and U12084 (N_12084,N_10130,N_10268);
xnor U12085 (N_12085,N_10441,N_10414);
xnor U12086 (N_12086,N_10264,N_10206);
nor U12087 (N_12087,N_10280,N_10405);
or U12088 (N_12088,N_10452,N_10733);
nor U12089 (N_12089,N_10172,N_10701);
nor U12090 (N_12090,N_11172,N_10983);
or U12091 (N_12091,N_11003,N_11216);
nor U12092 (N_12092,N_10170,N_11227);
and U12093 (N_12093,N_10660,N_10778);
nand U12094 (N_12094,N_10644,N_11030);
and U12095 (N_12095,N_10909,N_10564);
or U12096 (N_12096,N_10422,N_10310);
xnor U12097 (N_12097,N_10227,N_10185);
or U12098 (N_12098,N_10492,N_10242);
or U12099 (N_12099,N_10926,N_10174);
and U12100 (N_12100,N_10624,N_11029);
xor U12101 (N_12101,N_10266,N_10366);
xnor U12102 (N_12102,N_10665,N_10620);
nand U12103 (N_12103,N_10845,N_10064);
or U12104 (N_12104,N_10932,N_10200);
nor U12105 (N_12105,N_10384,N_10877);
nand U12106 (N_12106,N_10328,N_10908);
nand U12107 (N_12107,N_10806,N_11237);
nand U12108 (N_12108,N_10268,N_10966);
nor U12109 (N_12109,N_10749,N_10883);
nor U12110 (N_12110,N_10906,N_10460);
nand U12111 (N_12111,N_10227,N_10238);
and U12112 (N_12112,N_10581,N_10297);
and U12113 (N_12113,N_10762,N_11037);
or U12114 (N_12114,N_10769,N_11244);
xnor U12115 (N_12115,N_10210,N_10309);
or U12116 (N_12116,N_10553,N_10649);
or U12117 (N_12117,N_11031,N_10454);
xnor U12118 (N_12118,N_10370,N_10372);
nor U12119 (N_12119,N_10142,N_10212);
nor U12120 (N_12120,N_11093,N_10910);
nor U12121 (N_12121,N_11120,N_10512);
nor U12122 (N_12122,N_10690,N_10702);
xor U12123 (N_12123,N_10439,N_10037);
xnor U12124 (N_12124,N_10220,N_11189);
and U12125 (N_12125,N_10316,N_10780);
xnor U12126 (N_12126,N_10773,N_10486);
nand U12127 (N_12127,N_10505,N_11177);
xor U12128 (N_12128,N_11160,N_10810);
nor U12129 (N_12129,N_11140,N_10851);
or U12130 (N_12130,N_10426,N_10463);
and U12131 (N_12131,N_10752,N_10378);
and U12132 (N_12132,N_10990,N_10619);
and U12133 (N_12133,N_11034,N_10223);
nand U12134 (N_12134,N_10276,N_11105);
or U12135 (N_12135,N_10767,N_11230);
nand U12136 (N_12136,N_10161,N_11070);
nor U12137 (N_12137,N_10395,N_10782);
and U12138 (N_12138,N_10750,N_10929);
nand U12139 (N_12139,N_10795,N_11197);
xnor U12140 (N_12140,N_10526,N_11172);
nand U12141 (N_12141,N_10557,N_10960);
nor U12142 (N_12142,N_11204,N_10003);
or U12143 (N_12143,N_11048,N_11120);
or U12144 (N_12144,N_10787,N_10401);
or U12145 (N_12145,N_10139,N_10271);
xor U12146 (N_12146,N_10730,N_10142);
nand U12147 (N_12147,N_10939,N_11184);
nor U12148 (N_12148,N_11134,N_10161);
xor U12149 (N_12149,N_10970,N_10192);
xor U12150 (N_12150,N_10692,N_10097);
and U12151 (N_12151,N_10827,N_10230);
nand U12152 (N_12152,N_10645,N_10686);
and U12153 (N_12153,N_10115,N_10867);
nand U12154 (N_12154,N_10488,N_10909);
and U12155 (N_12155,N_10880,N_10153);
nor U12156 (N_12156,N_10825,N_10980);
nor U12157 (N_12157,N_11111,N_11218);
nand U12158 (N_12158,N_10520,N_10846);
or U12159 (N_12159,N_10683,N_10271);
nand U12160 (N_12160,N_11134,N_10028);
nor U12161 (N_12161,N_10851,N_10266);
or U12162 (N_12162,N_10929,N_10311);
xor U12163 (N_12163,N_10733,N_11180);
or U12164 (N_12164,N_10690,N_10784);
nand U12165 (N_12165,N_11133,N_10823);
or U12166 (N_12166,N_10895,N_11060);
nor U12167 (N_12167,N_10361,N_10245);
and U12168 (N_12168,N_10412,N_10044);
xnor U12169 (N_12169,N_11175,N_10131);
nand U12170 (N_12170,N_10202,N_10751);
or U12171 (N_12171,N_10131,N_10856);
and U12172 (N_12172,N_10007,N_10986);
nand U12173 (N_12173,N_10832,N_10051);
nand U12174 (N_12174,N_10115,N_10987);
and U12175 (N_12175,N_10563,N_10183);
nor U12176 (N_12176,N_10737,N_10602);
and U12177 (N_12177,N_10840,N_10824);
or U12178 (N_12178,N_10401,N_10980);
nor U12179 (N_12179,N_10984,N_10397);
and U12180 (N_12180,N_10812,N_10750);
nor U12181 (N_12181,N_11052,N_10746);
or U12182 (N_12182,N_11101,N_10449);
nor U12183 (N_12183,N_10777,N_11065);
or U12184 (N_12184,N_11244,N_10678);
nand U12185 (N_12185,N_10703,N_10733);
and U12186 (N_12186,N_10570,N_10326);
nor U12187 (N_12187,N_10363,N_10229);
and U12188 (N_12188,N_10687,N_10893);
and U12189 (N_12189,N_10302,N_10993);
and U12190 (N_12190,N_10847,N_10711);
nor U12191 (N_12191,N_11247,N_11148);
or U12192 (N_12192,N_10306,N_10209);
nand U12193 (N_12193,N_10111,N_10779);
xnor U12194 (N_12194,N_10331,N_10309);
nand U12195 (N_12195,N_10435,N_11047);
and U12196 (N_12196,N_10455,N_10833);
xor U12197 (N_12197,N_10666,N_10928);
xor U12198 (N_12198,N_10795,N_10168);
xor U12199 (N_12199,N_10661,N_10553);
nand U12200 (N_12200,N_10537,N_10050);
and U12201 (N_12201,N_10151,N_10559);
xor U12202 (N_12202,N_10982,N_10408);
and U12203 (N_12203,N_10238,N_10505);
and U12204 (N_12204,N_10446,N_10558);
and U12205 (N_12205,N_11034,N_10177);
nor U12206 (N_12206,N_10925,N_11047);
or U12207 (N_12207,N_10441,N_10371);
or U12208 (N_12208,N_10890,N_10316);
or U12209 (N_12209,N_10171,N_10875);
nor U12210 (N_12210,N_10652,N_10785);
nand U12211 (N_12211,N_10130,N_10655);
or U12212 (N_12212,N_11088,N_10599);
nor U12213 (N_12213,N_10104,N_11099);
xor U12214 (N_12214,N_10613,N_11143);
xor U12215 (N_12215,N_10605,N_11245);
and U12216 (N_12216,N_10807,N_10799);
nand U12217 (N_12217,N_11239,N_10759);
nor U12218 (N_12218,N_10336,N_10127);
or U12219 (N_12219,N_10965,N_10835);
and U12220 (N_12220,N_10636,N_11139);
and U12221 (N_12221,N_10523,N_10135);
or U12222 (N_12222,N_10168,N_11227);
nor U12223 (N_12223,N_10757,N_11106);
xor U12224 (N_12224,N_10425,N_11016);
or U12225 (N_12225,N_10173,N_10467);
nor U12226 (N_12226,N_10300,N_10653);
nand U12227 (N_12227,N_10885,N_10226);
xnor U12228 (N_12228,N_10931,N_10768);
nand U12229 (N_12229,N_10431,N_10079);
and U12230 (N_12230,N_10858,N_10595);
and U12231 (N_12231,N_10370,N_10813);
or U12232 (N_12232,N_10628,N_10586);
and U12233 (N_12233,N_10825,N_10040);
nand U12234 (N_12234,N_10276,N_10408);
or U12235 (N_12235,N_10555,N_10734);
or U12236 (N_12236,N_10182,N_10849);
or U12237 (N_12237,N_10416,N_10131);
nand U12238 (N_12238,N_10986,N_10253);
and U12239 (N_12239,N_10534,N_10325);
nand U12240 (N_12240,N_10310,N_10963);
and U12241 (N_12241,N_11214,N_10349);
nand U12242 (N_12242,N_10647,N_10017);
or U12243 (N_12243,N_10078,N_11218);
and U12244 (N_12244,N_10409,N_10889);
nor U12245 (N_12245,N_11161,N_10165);
nor U12246 (N_12246,N_11090,N_11113);
nand U12247 (N_12247,N_10037,N_10228);
xor U12248 (N_12248,N_10338,N_11033);
nand U12249 (N_12249,N_11201,N_11223);
xor U12250 (N_12250,N_10384,N_10464);
and U12251 (N_12251,N_10460,N_10937);
nor U12252 (N_12252,N_11130,N_10929);
nand U12253 (N_12253,N_10315,N_10316);
nand U12254 (N_12254,N_10757,N_10538);
xnor U12255 (N_12255,N_10556,N_10204);
nor U12256 (N_12256,N_10012,N_10481);
or U12257 (N_12257,N_10943,N_11235);
nand U12258 (N_12258,N_10584,N_11078);
nor U12259 (N_12259,N_10304,N_10985);
nand U12260 (N_12260,N_10974,N_11043);
xor U12261 (N_12261,N_10274,N_10289);
or U12262 (N_12262,N_10031,N_11035);
and U12263 (N_12263,N_10248,N_10139);
and U12264 (N_12264,N_10764,N_10146);
nand U12265 (N_12265,N_10277,N_10297);
nor U12266 (N_12266,N_11188,N_11206);
xor U12267 (N_12267,N_11232,N_10012);
or U12268 (N_12268,N_10319,N_10338);
or U12269 (N_12269,N_10187,N_10049);
nand U12270 (N_12270,N_10323,N_10811);
nand U12271 (N_12271,N_10000,N_10712);
or U12272 (N_12272,N_10272,N_10089);
nand U12273 (N_12273,N_10775,N_10140);
nor U12274 (N_12274,N_10138,N_10171);
xor U12275 (N_12275,N_10453,N_10820);
xnor U12276 (N_12276,N_11053,N_10912);
nor U12277 (N_12277,N_10602,N_11185);
nor U12278 (N_12278,N_10232,N_10483);
or U12279 (N_12279,N_10817,N_10050);
xnor U12280 (N_12280,N_10721,N_10792);
and U12281 (N_12281,N_10171,N_10433);
nor U12282 (N_12282,N_10013,N_10096);
and U12283 (N_12283,N_10760,N_10931);
and U12284 (N_12284,N_10823,N_11098);
and U12285 (N_12285,N_10790,N_11083);
or U12286 (N_12286,N_10978,N_10789);
nor U12287 (N_12287,N_10818,N_10313);
and U12288 (N_12288,N_10784,N_10310);
xor U12289 (N_12289,N_11210,N_11008);
nor U12290 (N_12290,N_10154,N_11061);
xor U12291 (N_12291,N_10883,N_10489);
or U12292 (N_12292,N_10452,N_10264);
or U12293 (N_12293,N_10685,N_10428);
nand U12294 (N_12294,N_10460,N_10903);
xnor U12295 (N_12295,N_10593,N_10944);
nor U12296 (N_12296,N_10435,N_11044);
nand U12297 (N_12297,N_10672,N_10707);
or U12298 (N_12298,N_10280,N_10536);
nor U12299 (N_12299,N_11005,N_11107);
nor U12300 (N_12300,N_10582,N_11136);
or U12301 (N_12301,N_10817,N_11233);
and U12302 (N_12302,N_10235,N_10036);
xnor U12303 (N_12303,N_10922,N_10030);
xnor U12304 (N_12304,N_11097,N_10822);
nand U12305 (N_12305,N_10652,N_10746);
nand U12306 (N_12306,N_10270,N_10849);
nand U12307 (N_12307,N_10792,N_10232);
or U12308 (N_12308,N_10172,N_10242);
or U12309 (N_12309,N_10057,N_11170);
and U12310 (N_12310,N_10421,N_10909);
xnor U12311 (N_12311,N_10263,N_11194);
nand U12312 (N_12312,N_11213,N_10320);
nor U12313 (N_12313,N_10264,N_11247);
nand U12314 (N_12314,N_10115,N_11188);
nand U12315 (N_12315,N_11039,N_10562);
xor U12316 (N_12316,N_11095,N_10794);
and U12317 (N_12317,N_10866,N_10200);
xnor U12318 (N_12318,N_10369,N_10155);
nand U12319 (N_12319,N_10473,N_11089);
or U12320 (N_12320,N_10001,N_10385);
nand U12321 (N_12321,N_11037,N_10241);
and U12322 (N_12322,N_10048,N_10247);
or U12323 (N_12323,N_10782,N_11096);
xnor U12324 (N_12324,N_10581,N_10093);
and U12325 (N_12325,N_11236,N_11219);
xnor U12326 (N_12326,N_10938,N_10812);
xnor U12327 (N_12327,N_10763,N_10766);
and U12328 (N_12328,N_11117,N_10458);
or U12329 (N_12329,N_10998,N_11109);
nand U12330 (N_12330,N_11197,N_10549);
or U12331 (N_12331,N_10887,N_11152);
nand U12332 (N_12332,N_11130,N_11142);
or U12333 (N_12333,N_10402,N_10167);
or U12334 (N_12334,N_10080,N_11221);
nand U12335 (N_12335,N_10989,N_10040);
nand U12336 (N_12336,N_10337,N_11081);
or U12337 (N_12337,N_10963,N_10486);
or U12338 (N_12338,N_11213,N_10798);
nor U12339 (N_12339,N_10785,N_10725);
nand U12340 (N_12340,N_11079,N_10449);
or U12341 (N_12341,N_10937,N_10504);
xnor U12342 (N_12342,N_10228,N_10104);
and U12343 (N_12343,N_10417,N_10221);
nand U12344 (N_12344,N_10006,N_10483);
and U12345 (N_12345,N_11237,N_10719);
or U12346 (N_12346,N_11054,N_10218);
nand U12347 (N_12347,N_10695,N_10709);
nand U12348 (N_12348,N_11127,N_10613);
and U12349 (N_12349,N_11016,N_10247);
and U12350 (N_12350,N_11120,N_10793);
or U12351 (N_12351,N_10992,N_10563);
xor U12352 (N_12352,N_10924,N_10422);
xnor U12353 (N_12353,N_11171,N_10903);
and U12354 (N_12354,N_11101,N_10789);
or U12355 (N_12355,N_11186,N_10107);
nand U12356 (N_12356,N_10526,N_11247);
or U12357 (N_12357,N_11103,N_10657);
xor U12358 (N_12358,N_10652,N_11086);
or U12359 (N_12359,N_10833,N_10430);
xnor U12360 (N_12360,N_10595,N_10915);
nor U12361 (N_12361,N_10142,N_11021);
nor U12362 (N_12362,N_10601,N_11156);
nand U12363 (N_12363,N_10063,N_10823);
xor U12364 (N_12364,N_10015,N_10650);
nor U12365 (N_12365,N_10402,N_10065);
xnor U12366 (N_12366,N_11195,N_10594);
nor U12367 (N_12367,N_10358,N_10278);
and U12368 (N_12368,N_10552,N_10377);
nor U12369 (N_12369,N_11175,N_10911);
nor U12370 (N_12370,N_10811,N_10891);
and U12371 (N_12371,N_10189,N_10572);
and U12372 (N_12372,N_10202,N_10604);
and U12373 (N_12373,N_10221,N_10484);
and U12374 (N_12374,N_10004,N_10712);
or U12375 (N_12375,N_10525,N_10881);
xor U12376 (N_12376,N_11008,N_10330);
nand U12377 (N_12377,N_10609,N_10758);
nand U12378 (N_12378,N_10537,N_10462);
nor U12379 (N_12379,N_11203,N_10023);
and U12380 (N_12380,N_11102,N_11238);
nor U12381 (N_12381,N_10088,N_11230);
xnor U12382 (N_12382,N_10453,N_10591);
or U12383 (N_12383,N_10468,N_10744);
nor U12384 (N_12384,N_10829,N_10187);
xnor U12385 (N_12385,N_10560,N_10678);
nand U12386 (N_12386,N_10998,N_11187);
nand U12387 (N_12387,N_10338,N_11162);
or U12388 (N_12388,N_10423,N_11170);
and U12389 (N_12389,N_10957,N_10928);
nor U12390 (N_12390,N_10305,N_11013);
nand U12391 (N_12391,N_10461,N_10433);
nor U12392 (N_12392,N_11240,N_11212);
and U12393 (N_12393,N_10127,N_11008);
or U12394 (N_12394,N_10301,N_10782);
or U12395 (N_12395,N_10475,N_11045);
xor U12396 (N_12396,N_10407,N_10014);
xnor U12397 (N_12397,N_10692,N_10647);
xor U12398 (N_12398,N_10760,N_10620);
nand U12399 (N_12399,N_11199,N_11174);
and U12400 (N_12400,N_10959,N_10195);
nand U12401 (N_12401,N_10719,N_10134);
or U12402 (N_12402,N_10867,N_10133);
nor U12403 (N_12403,N_10306,N_10454);
xor U12404 (N_12404,N_10428,N_10184);
xnor U12405 (N_12405,N_10405,N_11230);
and U12406 (N_12406,N_10014,N_10866);
or U12407 (N_12407,N_10045,N_11217);
or U12408 (N_12408,N_10231,N_11187);
and U12409 (N_12409,N_10440,N_10232);
and U12410 (N_12410,N_11235,N_11116);
xor U12411 (N_12411,N_10059,N_10716);
nor U12412 (N_12412,N_10628,N_10233);
xnor U12413 (N_12413,N_10874,N_10768);
nand U12414 (N_12414,N_10012,N_11197);
nand U12415 (N_12415,N_11215,N_10952);
nand U12416 (N_12416,N_10879,N_10005);
nand U12417 (N_12417,N_10229,N_10469);
and U12418 (N_12418,N_10835,N_11057);
nand U12419 (N_12419,N_10280,N_10915);
nand U12420 (N_12420,N_10588,N_10338);
or U12421 (N_12421,N_10739,N_11004);
xor U12422 (N_12422,N_10730,N_10264);
nand U12423 (N_12423,N_10961,N_10593);
nor U12424 (N_12424,N_10993,N_11215);
or U12425 (N_12425,N_10826,N_10678);
nor U12426 (N_12426,N_11142,N_10545);
and U12427 (N_12427,N_10189,N_11224);
and U12428 (N_12428,N_11206,N_10124);
and U12429 (N_12429,N_10150,N_10531);
nor U12430 (N_12430,N_10069,N_10868);
nand U12431 (N_12431,N_10258,N_11238);
nor U12432 (N_12432,N_10731,N_11203);
or U12433 (N_12433,N_10727,N_10319);
nor U12434 (N_12434,N_10595,N_11021);
or U12435 (N_12435,N_10235,N_10592);
nor U12436 (N_12436,N_10979,N_11056);
nand U12437 (N_12437,N_10582,N_10923);
nand U12438 (N_12438,N_10927,N_10129);
nand U12439 (N_12439,N_10860,N_10646);
or U12440 (N_12440,N_10972,N_10329);
nor U12441 (N_12441,N_10144,N_10074);
nor U12442 (N_12442,N_10759,N_10336);
nor U12443 (N_12443,N_10832,N_11167);
or U12444 (N_12444,N_10114,N_10858);
or U12445 (N_12445,N_10951,N_10968);
nand U12446 (N_12446,N_10625,N_10891);
xnor U12447 (N_12447,N_10460,N_10711);
and U12448 (N_12448,N_10197,N_10036);
and U12449 (N_12449,N_11219,N_10107);
nand U12450 (N_12450,N_10608,N_10423);
or U12451 (N_12451,N_10318,N_11094);
nor U12452 (N_12452,N_10548,N_10102);
nor U12453 (N_12453,N_10712,N_10317);
xnor U12454 (N_12454,N_11211,N_11001);
nor U12455 (N_12455,N_11248,N_11216);
xor U12456 (N_12456,N_10947,N_10811);
or U12457 (N_12457,N_10101,N_10347);
xnor U12458 (N_12458,N_11142,N_11012);
or U12459 (N_12459,N_10966,N_10659);
nand U12460 (N_12460,N_10842,N_10880);
or U12461 (N_12461,N_10358,N_10440);
and U12462 (N_12462,N_10956,N_10116);
and U12463 (N_12463,N_10392,N_10617);
nand U12464 (N_12464,N_10549,N_11246);
xor U12465 (N_12465,N_10939,N_10106);
or U12466 (N_12466,N_10580,N_10592);
nor U12467 (N_12467,N_11239,N_11088);
nor U12468 (N_12468,N_11109,N_10835);
and U12469 (N_12469,N_11170,N_11151);
xnor U12470 (N_12470,N_10695,N_10518);
xor U12471 (N_12471,N_10696,N_10960);
or U12472 (N_12472,N_10487,N_11113);
xor U12473 (N_12473,N_10801,N_10247);
nand U12474 (N_12474,N_10610,N_10004);
and U12475 (N_12475,N_11149,N_10547);
and U12476 (N_12476,N_10146,N_10096);
nand U12477 (N_12477,N_11054,N_11212);
or U12478 (N_12478,N_11061,N_10907);
and U12479 (N_12479,N_10774,N_10829);
xor U12480 (N_12480,N_11243,N_10776);
xor U12481 (N_12481,N_10313,N_10894);
nand U12482 (N_12482,N_10315,N_10177);
nand U12483 (N_12483,N_10054,N_10408);
nand U12484 (N_12484,N_11137,N_10582);
and U12485 (N_12485,N_11029,N_11164);
or U12486 (N_12486,N_10227,N_10746);
and U12487 (N_12487,N_10913,N_11062);
nand U12488 (N_12488,N_10476,N_10450);
nor U12489 (N_12489,N_10874,N_10608);
nand U12490 (N_12490,N_10068,N_10211);
or U12491 (N_12491,N_11121,N_10998);
and U12492 (N_12492,N_11097,N_10675);
nor U12493 (N_12493,N_10711,N_10218);
xor U12494 (N_12494,N_10162,N_11152);
or U12495 (N_12495,N_10249,N_10224);
nor U12496 (N_12496,N_11055,N_10203);
or U12497 (N_12497,N_10426,N_10717);
nor U12498 (N_12498,N_10237,N_10415);
and U12499 (N_12499,N_11171,N_11140);
nand U12500 (N_12500,N_12334,N_11875);
xnor U12501 (N_12501,N_12030,N_11587);
and U12502 (N_12502,N_12226,N_11990);
and U12503 (N_12503,N_11674,N_11568);
nor U12504 (N_12504,N_11931,N_11452);
and U12505 (N_12505,N_11838,N_12212);
nor U12506 (N_12506,N_12323,N_11262);
and U12507 (N_12507,N_11324,N_11684);
nand U12508 (N_12508,N_12231,N_12169);
nor U12509 (N_12509,N_12408,N_11398);
nor U12510 (N_12510,N_11626,N_12383);
nand U12511 (N_12511,N_11852,N_11708);
or U12512 (N_12512,N_11279,N_11645);
nand U12513 (N_12513,N_11910,N_11333);
nor U12514 (N_12514,N_12019,N_11507);
nand U12515 (N_12515,N_12402,N_11636);
xnor U12516 (N_12516,N_11331,N_11999);
nor U12517 (N_12517,N_12477,N_11476);
nor U12518 (N_12518,N_12213,N_11969);
xor U12519 (N_12519,N_11478,N_11375);
nand U12520 (N_12520,N_12374,N_11276);
or U12521 (N_12521,N_11939,N_12349);
and U12522 (N_12522,N_11797,N_11935);
xor U12523 (N_12523,N_11892,N_12494);
nor U12524 (N_12524,N_12443,N_12411);
or U12525 (N_12525,N_11702,N_11434);
nor U12526 (N_12526,N_12435,N_11715);
or U12527 (N_12527,N_12307,N_12051);
or U12528 (N_12528,N_11914,N_11421);
xnor U12529 (N_12529,N_11401,N_12220);
xnor U12530 (N_12530,N_12309,N_11533);
nor U12531 (N_12531,N_11686,N_12109);
nor U12532 (N_12532,N_12321,N_11778);
xnor U12533 (N_12533,N_11815,N_12485);
xor U12534 (N_12534,N_11373,N_11558);
xor U12535 (N_12535,N_12209,N_11773);
nand U12536 (N_12536,N_11295,N_11376);
xnor U12537 (N_12537,N_11657,N_12407);
xnor U12538 (N_12538,N_12018,N_11497);
or U12539 (N_12539,N_12430,N_11997);
and U12540 (N_12540,N_11275,N_11573);
and U12541 (N_12541,N_11588,N_11747);
nand U12542 (N_12542,N_11802,N_11406);
nand U12543 (N_12543,N_11785,N_12341);
nor U12544 (N_12544,N_11775,N_12160);
or U12545 (N_12545,N_11627,N_11765);
or U12546 (N_12546,N_11368,N_11466);
xnor U12547 (N_12547,N_12172,N_11728);
and U12548 (N_12548,N_11795,N_11515);
nand U12549 (N_12549,N_11799,N_11800);
nor U12550 (N_12550,N_11296,N_11944);
or U12551 (N_12551,N_12211,N_12175);
nor U12552 (N_12552,N_12085,N_12029);
nor U12553 (N_12553,N_12056,N_11283);
and U12554 (N_12554,N_12215,N_11846);
and U12555 (N_12555,N_12201,N_11536);
or U12556 (N_12556,N_11635,N_11766);
and U12557 (N_12557,N_12222,N_11679);
nand U12558 (N_12558,N_11571,N_11693);
and U12559 (N_12559,N_12134,N_11943);
nor U12560 (N_12560,N_11856,N_11726);
nor U12561 (N_12561,N_12141,N_12096);
nor U12562 (N_12562,N_11362,N_12204);
or U12563 (N_12563,N_11941,N_11574);
nand U12564 (N_12564,N_11263,N_11567);
nand U12565 (N_12565,N_11489,N_12199);
nor U12566 (N_12566,N_12296,N_12177);
xnor U12567 (N_12567,N_11970,N_11600);
and U12568 (N_12568,N_11719,N_12126);
or U12569 (N_12569,N_11818,N_11869);
or U12570 (N_12570,N_12099,N_12406);
nor U12571 (N_12571,N_11413,N_12198);
xor U12572 (N_12572,N_12456,N_11641);
nor U12573 (N_12573,N_11624,N_12033);
and U12574 (N_12574,N_11353,N_11481);
and U12575 (N_12575,N_12373,N_12100);
nand U12576 (N_12576,N_11357,N_12291);
or U12577 (N_12577,N_11953,N_12398);
and U12578 (N_12578,N_11666,N_11658);
nand U12579 (N_12579,N_11864,N_11435);
or U12580 (N_12580,N_12252,N_11267);
xor U12581 (N_12581,N_11720,N_11438);
and U12582 (N_12582,N_11891,N_11330);
nor U12583 (N_12583,N_11902,N_12132);
nor U12584 (N_12584,N_12083,N_11467);
or U12585 (N_12585,N_12144,N_11447);
or U12586 (N_12586,N_12433,N_11655);
nor U12587 (N_12587,N_11252,N_11359);
nand U12588 (N_12588,N_11286,N_11819);
and U12589 (N_12589,N_12289,N_12377);
xnor U12590 (N_12590,N_11534,N_12354);
nand U12591 (N_12591,N_12326,N_11549);
xor U12592 (N_12592,N_11502,N_12042);
or U12593 (N_12593,N_11973,N_12125);
nor U12594 (N_12594,N_11312,N_12228);
nor U12595 (N_12595,N_11493,N_11423);
nand U12596 (N_12596,N_11964,N_12118);
nand U12597 (N_12597,N_12437,N_11451);
xor U12598 (N_12598,N_12483,N_12188);
or U12599 (N_12599,N_12223,N_11590);
xnor U12600 (N_12600,N_11461,N_11881);
or U12601 (N_12601,N_12255,N_11586);
or U12602 (N_12602,N_11299,N_11794);
nand U12603 (N_12603,N_11683,N_12330);
or U12604 (N_12604,N_11724,N_11991);
nor U12605 (N_12605,N_11979,N_11448);
and U12606 (N_12606,N_12470,N_12282);
nand U12607 (N_12607,N_12122,N_12185);
and U12608 (N_12608,N_11705,N_12396);
nand U12609 (N_12609,N_12283,N_11430);
nand U12610 (N_12610,N_12343,N_11374);
nand U12611 (N_12611,N_12195,N_12284);
and U12612 (N_12612,N_12459,N_11858);
xnor U12613 (N_12613,N_11524,N_11789);
nand U12614 (N_12614,N_12305,N_12129);
nor U12615 (N_12615,N_12389,N_11397);
and U12616 (N_12616,N_12062,N_11685);
nor U12617 (N_12617,N_12465,N_11909);
or U12618 (N_12618,N_11922,N_11475);
xnor U12619 (N_12619,N_12165,N_11872);
and U12620 (N_12620,N_11425,N_12439);
and U12621 (N_12621,N_12166,N_12445);
xor U12622 (N_12622,N_11446,N_11455);
nor U12623 (N_12623,N_12131,N_12194);
or U12624 (N_12624,N_11700,N_11848);
and U12625 (N_12625,N_12397,N_12332);
nor U12626 (N_12626,N_11623,N_11537);
or U12627 (N_12627,N_11343,N_12176);
or U12628 (N_12628,N_12329,N_12210);
and U12629 (N_12629,N_11517,N_12164);
or U12630 (N_12630,N_12196,N_11965);
nor U12631 (N_12631,N_11668,N_11394);
nand U12632 (N_12632,N_12191,N_12487);
nand U12633 (N_12633,N_12192,N_11598);
nor U12634 (N_12634,N_12367,N_12225);
or U12635 (N_12635,N_11584,N_12026);
nor U12636 (N_12636,N_12163,N_12257);
nand U12637 (N_12637,N_11740,N_11566);
nand U12638 (N_12638,N_11580,N_11621);
xnor U12639 (N_12639,N_11436,N_11727);
nand U12640 (N_12640,N_11561,N_11923);
xor U12641 (N_12641,N_11649,N_11912);
xnor U12642 (N_12642,N_12253,N_12145);
xor U12643 (N_12643,N_11801,N_12286);
xor U12644 (N_12644,N_12107,N_12205);
xor U12645 (N_12645,N_12092,N_11605);
or U12646 (N_12646,N_11487,N_12369);
or U12647 (N_12647,N_11601,N_12313);
nand U12648 (N_12648,N_11273,N_12234);
nand U12649 (N_12649,N_12281,N_11433);
or U12650 (N_12650,N_11297,N_11745);
nor U12651 (N_12651,N_12386,N_12152);
nand U12652 (N_12652,N_12073,N_11615);
nand U12653 (N_12653,N_11774,N_11871);
and U12654 (N_12654,N_12306,N_11490);
or U12655 (N_12655,N_12379,N_11913);
xnor U12656 (N_12656,N_11464,N_12499);
xnor U12657 (N_12657,N_11553,N_11281);
nor U12658 (N_12658,N_11529,N_11689);
and U12659 (N_12659,N_11651,N_11335);
xor U12660 (N_12660,N_12111,N_11748);
or U12661 (N_12661,N_12009,N_11697);
or U12662 (N_12662,N_11604,N_12393);
and U12663 (N_12663,N_12048,N_11753);
and U12664 (N_12664,N_12346,N_12424);
nand U12665 (N_12665,N_11501,N_11250);
xnor U12666 (N_12666,N_11602,N_12221);
and U12667 (N_12667,N_11504,N_11760);
xor U12668 (N_12668,N_11739,N_11508);
nor U12669 (N_12669,N_12387,N_11255);
and U12670 (N_12670,N_12075,N_11995);
nand U12671 (N_12671,N_12475,N_11396);
nor U12672 (N_12672,N_11405,N_12368);
or U12673 (N_12673,N_11264,N_11827);
nor U12674 (N_12674,N_11652,N_11477);
xnor U12675 (N_12675,N_12143,N_11890);
nand U12676 (N_12676,N_11659,N_11366);
nor U12677 (N_12677,N_11293,N_12431);
nor U12678 (N_12678,N_12298,N_12245);
xor U12679 (N_12679,N_12034,N_12136);
xor U12680 (N_12680,N_11538,N_12130);
or U12681 (N_12681,N_11422,N_11387);
nor U12682 (N_12682,N_12300,N_12401);
and U12683 (N_12683,N_12361,N_11850);
nor U12684 (N_12684,N_11690,N_11593);
or U12685 (N_12685,N_11514,N_11480);
and U12686 (N_12686,N_11418,N_11551);
xor U12687 (N_12687,N_12327,N_11642);
nor U12688 (N_12688,N_11783,N_11288);
nand U12689 (N_12689,N_12405,N_11866);
or U12690 (N_12690,N_12376,N_12032);
and U12691 (N_12691,N_11344,N_11400);
or U12692 (N_12692,N_11287,N_12458);
and U12693 (N_12693,N_11861,N_12295);
and U12694 (N_12694,N_11810,N_12279);
or U12695 (N_12695,N_11661,N_12348);
and U12696 (N_12696,N_11518,N_12390);
nand U12697 (N_12697,N_11429,N_11579);
nand U12698 (N_12698,N_12123,N_12310);
and U12699 (N_12699,N_12496,N_12412);
and U12700 (N_12700,N_12473,N_11831);
or U12701 (N_12701,N_12214,N_12498);
xor U12702 (N_12702,N_11860,N_11749);
or U12703 (N_12703,N_12187,N_11730);
or U12704 (N_12704,N_11959,N_11614);
or U12705 (N_12705,N_11793,N_11301);
nand U12706 (N_12706,N_12243,N_11315);
and U12707 (N_12707,N_11687,N_12106);
or U12708 (N_12708,N_12474,N_12331);
or U12709 (N_12709,N_11611,N_12432);
or U12710 (N_12710,N_11417,N_11257);
xnor U12711 (N_12711,N_11884,N_12380);
xnor U12712 (N_12712,N_12482,N_12442);
or U12713 (N_12713,N_11329,N_11901);
nand U12714 (N_12714,N_12035,N_11332);
and U12715 (N_12715,N_12087,N_12014);
nand U12716 (N_12716,N_12128,N_12202);
or U12717 (N_12717,N_12149,N_12248);
or U12718 (N_12718,N_11613,N_11812);
and U12719 (N_12719,N_11826,N_12124);
or U12720 (N_12720,N_11814,N_11951);
or U12721 (N_12721,N_11302,N_11867);
or U12722 (N_12722,N_11894,N_11998);
and U12723 (N_12723,N_11414,N_11703);
nand U12724 (N_12724,N_11261,N_12311);
or U12725 (N_12725,N_12001,N_12059);
nand U12726 (N_12726,N_12469,N_11936);
nand U12727 (N_12727,N_11419,N_12338);
and U12728 (N_12728,N_11805,N_11532);
nor U12729 (N_12729,N_12325,N_12312);
nand U12730 (N_12730,N_12449,N_11522);
or U12731 (N_12731,N_11628,N_11842);
nand U12732 (N_12732,N_11948,N_11771);
nor U12733 (N_12733,N_11495,N_11638);
or U12734 (N_12734,N_12044,N_12491);
nor U12735 (N_12735,N_12319,N_11907);
or U12736 (N_12736,N_12121,N_12015);
or U12737 (N_12737,N_11407,N_11284);
nand U12738 (N_12738,N_11844,N_12242);
or U12739 (N_12739,N_12471,N_11701);
nor U12740 (N_12740,N_11439,N_12171);
xor U12741 (N_12741,N_11355,N_12237);
nand U12742 (N_12742,N_11443,N_12448);
and U12743 (N_12743,N_12249,N_11639);
and U12744 (N_12744,N_12489,N_11325);
nand U12745 (N_12745,N_12247,N_11980);
and U12746 (N_12746,N_11699,N_11757);
or U12747 (N_12747,N_11971,N_11554);
and U12748 (N_12748,N_12084,N_11606);
xor U12749 (N_12749,N_12318,N_11963);
nand U12750 (N_12750,N_12478,N_12037);
nor U12751 (N_12751,N_11498,N_12434);
nor U12752 (N_12752,N_11806,N_12404);
xor U12753 (N_12753,N_12182,N_12425);
nand U12754 (N_12754,N_12022,N_11555);
nor U12755 (N_12755,N_12046,N_11752);
or U12756 (N_12756,N_11460,N_11472);
nor U12757 (N_12757,N_12352,N_11632);
xor U12758 (N_12758,N_11918,N_11637);
or U12759 (N_12759,N_11839,N_11383);
or U12760 (N_12760,N_12161,N_11986);
nand U12761 (N_12761,N_12285,N_11395);
or U12762 (N_12762,N_11449,N_11432);
nand U12763 (N_12763,N_11424,N_11440);
nand U12764 (N_12764,N_11525,N_12197);
nor U12765 (N_12765,N_11928,N_11854);
nor U12766 (N_12766,N_12292,N_12098);
xnor U12767 (N_12767,N_11847,N_11706);
nor U12768 (N_12768,N_12208,N_11294);
or U12769 (N_12769,N_12277,N_11259);
nor U12770 (N_12770,N_12039,N_12230);
nor U12771 (N_12771,N_11988,N_12333);
nor U12772 (N_12772,N_12244,N_11987);
xnor U12773 (N_12773,N_12495,N_11880);
nand U12774 (N_12774,N_11303,N_12480);
and U12775 (N_12775,N_12154,N_11653);
or U12776 (N_12776,N_12464,N_11692);
nand U12777 (N_12777,N_12133,N_12429);
xor U12778 (N_12778,N_11305,N_11565);
and U12779 (N_12779,N_11318,N_11560);
nor U12780 (N_12780,N_11754,N_12103);
and U12781 (N_12781,N_11798,N_11589);
xnor U12782 (N_12782,N_12440,N_12423);
or U12783 (N_12783,N_11863,N_11254);
nor U12784 (N_12784,N_11306,N_11688);
nand U12785 (N_12785,N_12254,N_11469);
xnor U12786 (N_12786,N_11711,N_12421);
nand U12787 (N_12787,N_11932,N_12320);
xnor U12788 (N_12788,N_12382,N_12274);
or U12789 (N_12789,N_11340,N_12267);
nand U12790 (N_12790,N_11895,N_12224);
xnor U12791 (N_12791,N_11535,N_11924);
nand U12792 (N_12792,N_11807,N_11746);
nand U12793 (N_12793,N_11742,N_12078);
nor U12794 (N_12794,N_11879,N_11870);
nand U12795 (N_12795,N_11888,N_12476);
or U12796 (N_12796,N_11712,N_12114);
and U12797 (N_12797,N_11542,N_11736);
xor U12798 (N_12798,N_11270,N_12216);
xnor U12799 (N_12799,N_12219,N_12358);
xor U12800 (N_12800,N_12259,N_11269);
and U12801 (N_12801,N_11350,N_11713);
and U12802 (N_12802,N_11966,N_12265);
nor U12803 (N_12803,N_12345,N_11280);
nand U12804 (N_12804,N_12120,N_12273);
nand U12805 (N_12805,N_12488,N_12385);
or U12806 (N_12806,N_11337,N_12372);
and U12807 (N_12807,N_11483,N_11426);
nand U12808 (N_12808,N_12146,N_11955);
nor U12809 (N_12809,N_11519,N_11485);
and U12810 (N_12810,N_12142,N_11358);
and U12811 (N_12811,N_11817,N_12180);
nor U12812 (N_12812,N_11564,N_11972);
xnor U12813 (N_12813,N_12066,N_11572);
and U12814 (N_12814,N_11882,N_11360);
nor U12815 (N_12815,N_12184,N_11528);
or U12816 (N_12816,N_11516,N_11442);
xor U12817 (N_12817,N_12317,N_12436);
nor U12818 (N_12818,N_12147,N_12293);
xor U12819 (N_12819,N_11716,N_12416);
xor U12820 (N_12820,N_11550,N_11876);
nor U12821 (N_12821,N_12189,N_12117);
xor U12822 (N_12822,N_11769,N_11386);
nand U12823 (N_12823,N_11342,N_11889);
xnor U12824 (N_12824,N_11512,N_12155);
xor U12825 (N_12825,N_11364,N_11834);
nand U12826 (N_12826,N_11629,N_11622);
nor U12827 (N_12827,N_11384,N_11796);
xor U12828 (N_12828,N_11725,N_11729);
xnor U12829 (N_12829,N_12240,N_11505);
xnor U12830 (N_12830,N_11906,N_11527);
nor U12831 (N_12831,N_12262,N_12183);
nand U12832 (N_12832,N_11857,N_12316);
xnor U12833 (N_12833,N_12441,N_11723);
xnor U12834 (N_12834,N_11570,N_11268);
and U12835 (N_12835,N_11908,N_11833);
xor U12836 (N_12836,N_11462,N_11513);
nand U12837 (N_12837,N_11595,N_12270);
or U12838 (N_12838,N_11791,N_12472);
nand U12839 (N_12839,N_11321,N_11996);
xnor U12840 (N_12840,N_11695,N_11897);
xnor U12841 (N_12841,N_11777,N_11569);
xor U12842 (N_12842,N_11619,N_11751);
and U12843 (N_12843,N_11272,N_11921);
nand U12844 (N_12844,N_11367,N_11552);
or U12845 (N_12845,N_12094,N_12112);
nand U12846 (N_12846,N_12454,N_11258);
nor U12847 (N_12847,N_11934,N_11671);
nor U12848 (N_12848,N_11597,N_11468);
or U12849 (N_12849,N_12236,N_11738);
xor U12850 (N_12850,N_11691,N_11544);
nor U12851 (N_12851,N_12467,N_11582);
nor U12852 (N_12852,N_11886,N_11563);
nand U12853 (N_12853,N_11670,N_11278);
xor U12854 (N_12854,N_11954,N_11285);
xnor U12855 (N_12855,N_11823,N_11946);
or U12856 (N_12856,N_12359,N_12012);
and U12857 (N_12857,N_11486,N_11585);
or U12858 (N_12858,N_12027,N_11506);
xor U12859 (N_12859,N_12162,N_12303);
and U12860 (N_12860,N_11616,N_11511);
nand U12861 (N_12861,N_12079,N_12008);
or U12862 (N_12862,N_11764,N_11577);
xnor U12863 (N_12863,N_12088,N_12428);
nand U12864 (N_12864,N_12113,N_12074);
nor U12865 (N_12865,N_11694,N_11371);
or U12866 (N_12866,N_12297,N_12420);
or U12867 (N_12867,N_11804,N_11381);
or U12868 (N_12868,N_12468,N_11415);
and U12869 (N_12869,N_12399,N_12006);
nor U12870 (N_12870,N_11457,N_11410);
nor U12871 (N_12871,N_11408,N_11993);
nand U12872 (N_12872,N_11859,N_11427);
or U12873 (N_12873,N_11441,N_12378);
nand U12874 (N_12874,N_11416,N_11596);
nor U12875 (N_12875,N_12031,N_11351);
or U12876 (N_12876,N_12233,N_11898);
or U12877 (N_12877,N_11458,N_11821);
nand U12878 (N_12878,N_12238,N_11737);
and U12879 (N_12879,N_11710,N_11920);
xnor U12880 (N_12880,N_11562,N_11664);
nand U12881 (N_12881,N_11917,N_11938);
nor U12882 (N_12882,N_12347,N_12025);
nor U12883 (N_12883,N_12115,N_12021);
xor U12884 (N_12884,N_12381,N_12452);
nor U12885 (N_12885,N_11669,N_11307);
xnor U12886 (N_12886,N_11646,N_12045);
and U12887 (N_12887,N_12064,N_11835);
xor U12888 (N_12888,N_12350,N_11952);
xnor U12889 (N_12889,N_11885,N_12360);
nand U12890 (N_12890,N_11811,N_11378);
nand U12891 (N_12891,N_12336,N_11482);
xnor U12892 (N_12892,N_11780,N_12076);
xor U12893 (N_12893,N_12328,N_11992);
and U12894 (N_12894,N_11456,N_12186);
and U12895 (N_12895,N_12040,N_11790);
nand U12896 (N_12896,N_12461,N_11349);
and U12897 (N_12897,N_11548,N_12093);
nand U12898 (N_12898,N_12446,N_12190);
nor U12899 (N_12899,N_12353,N_11837);
xor U12900 (N_12900,N_11832,N_12426);
nor U12901 (N_12901,N_11559,N_11784);
nor U12902 (N_12902,N_11316,N_11968);
nand U12903 (N_12903,N_12068,N_12258);
nand U12904 (N_12904,N_12451,N_12174);
and U12905 (N_12905,N_11650,N_12067);
or U12906 (N_12906,N_12097,N_11828);
xnor U12907 (N_12907,N_12486,N_11663);
nor U12908 (N_12908,N_11412,N_11292);
or U12909 (N_12909,N_11682,N_11454);
xor U12910 (N_12910,N_12250,N_11896);
xor U12911 (N_12911,N_11370,N_12235);
nor U12912 (N_12912,N_12391,N_12139);
nor U12913 (N_12913,N_12036,N_11768);
nor U12914 (N_12914,N_12127,N_11759);
xnor U12915 (N_12915,N_11782,N_12049);
nor U12916 (N_12916,N_11665,N_11274);
or U12917 (N_12917,N_12153,N_12357);
or U12918 (N_12918,N_12304,N_11741);
xor U12919 (N_12919,N_11289,N_11260);
and U12920 (N_12920,N_12414,N_12447);
nor U12921 (N_12921,N_12264,N_11925);
nor U12922 (N_12922,N_11709,N_12041);
xnor U12923 (N_12923,N_11949,N_11392);
and U12924 (N_12924,N_12028,N_11776);
or U12925 (N_12925,N_11251,N_11531);
xnor U12926 (N_12926,N_11680,N_12444);
and U12927 (N_12927,N_11758,N_11873);
nor U12928 (N_12928,N_11905,N_11471);
and U12929 (N_12929,N_12371,N_11445);
nor U12930 (N_12930,N_11609,N_12324);
xnor U12931 (N_12931,N_12070,N_11750);
xnor U12932 (N_12932,N_11372,N_11958);
nor U12933 (N_12933,N_12339,N_11382);
nor U12934 (N_12934,N_12102,N_11271);
xor U12935 (N_12935,N_12410,N_11520);
nor U12936 (N_12936,N_11494,N_11822);
or U12937 (N_12937,N_11983,N_11961);
or U12938 (N_12938,N_12355,N_12150);
and U12939 (N_12939,N_12272,N_11678);
nand U12940 (N_12940,N_12043,N_11530);
or U12941 (N_12941,N_11523,N_11291);
nor U12942 (N_12942,N_12460,N_11770);
xor U12943 (N_12943,N_11403,N_12137);
or U12944 (N_12944,N_11761,N_11660);
nand U12945 (N_12945,N_11735,N_12256);
and U12946 (N_12946,N_11911,N_12010);
and U12947 (N_12947,N_11904,N_11836);
nor U12948 (N_12948,N_12290,N_12417);
and U12949 (N_12949,N_11625,N_11803);
or U12950 (N_12950,N_12229,N_12322);
or U12951 (N_12951,N_11865,N_12344);
nand U12952 (N_12952,N_11341,N_12151);
and U12953 (N_12953,N_12002,N_11385);
xnor U12954 (N_12954,N_11957,N_12157);
and U12955 (N_12955,N_11633,N_12455);
nand U12956 (N_12956,N_11521,N_11594);
nor U12957 (N_12957,N_11479,N_11300);
or U12958 (N_12958,N_11320,N_12217);
and U12959 (N_12959,N_12302,N_12119);
xnor U12960 (N_12960,N_11265,N_12024);
xor U12961 (N_12961,N_11672,N_12466);
nor U12962 (N_12962,N_11323,N_12438);
or U12963 (N_12963,N_11450,N_12206);
nor U12964 (N_12964,N_11608,N_11640);
nor U12965 (N_12965,N_11266,N_11734);
nor U12966 (N_12966,N_12138,N_11820);
or U12967 (N_12967,N_11339,N_12400);
and U12968 (N_12968,N_11930,N_11813);
or U12969 (N_12969,N_12462,N_12308);
xor U12970 (N_12970,N_12158,N_12101);
or U12971 (N_12971,N_12016,N_11610);
and U12972 (N_12972,N_12271,N_12193);
or U12973 (N_12973,N_12057,N_11298);
nor U12974 (N_12974,N_11313,N_11974);
and U12975 (N_12975,N_12203,N_11714);
and U12976 (N_12976,N_11919,N_12314);
nand U12977 (N_12977,N_12268,N_12362);
and U12978 (N_12978,N_12492,N_12072);
and U12979 (N_12979,N_11363,N_11576);
xor U12980 (N_12980,N_12261,N_11676);
or U12981 (N_12981,N_11841,N_12065);
xnor U12982 (N_12982,N_11772,N_11862);
or U12983 (N_12983,N_11781,N_11463);
nor U12984 (N_12984,N_11704,N_12061);
nor U12985 (N_12985,N_11786,N_12450);
xnor U12986 (N_12986,N_12419,N_11978);
or U12987 (N_12987,N_11756,N_11453);
or U12988 (N_12988,N_12071,N_11592);
xor U12989 (N_12989,N_11960,N_11314);
nor U12990 (N_12990,N_11940,N_11620);
xnor U12991 (N_12991,N_12178,N_12409);
or U12992 (N_12992,N_12490,N_12058);
or U12993 (N_12993,N_12418,N_12457);
or U12994 (N_12994,N_11887,N_11634);
and U12995 (N_12995,N_11399,N_12038);
xor U12996 (N_12996,N_12052,N_12013);
or U12997 (N_12997,N_12497,N_12340);
or U12998 (N_12998,N_11903,N_12395);
xor U12999 (N_12999,N_11962,N_11369);
xnor U13000 (N_13000,N_12005,N_11420);
and U13001 (N_13001,N_12269,N_12080);
nor U13002 (N_13002,N_11868,N_11809);
and U13003 (N_13003,N_12337,N_11336);
nor U13004 (N_13004,N_11644,N_11825);
nor U13005 (N_13005,N_11982,N_11763);
and U13006 (N_13006,N_12463,N_11681);
and U13007 (N_13007,N_11732,N_11603);
and U13008 (N_13008,N_11843,N_11977);
and U13009 (N_13009,N_11607,N_11411);
or U13010 (N_13010,N_11792,N_11916);
xnor U13011 (N_13011,N_11308,N_11322);
nand U13012 (N_13012,N_11779,N_11929);
xnor U13013 (N_13013,N_12181,N_11354);
nor U13014 (N_13014,N_11851,N_11981);
and U13015 (N_13015,N_11317,N_12365);
nor U13016 (N_13016,N_12140,N_11540);
nor U13017 (N_13017,N_11282,N_12091);
and U13018 (N_13018,N_11583,N_12110);
and U13019 (N_13019,N_11365,N_11618);
xor U13020 (N_13020,N_11346,N_12227);
xor U13021 (N_13021,N_12493,N_11877);
xor U13022 (N_13022,N_11762,N_12413);
nor U13023 (N_13023,N_12294,N_11677);
nor U13024 (N_13024,N_11824,N_12108);
nor U13025 (N_13025,N_11488,N_11547);
xnor U13026 (N_13026,N_11830,N_11277);
or U13027 (N_13027,N_11492,N_12388);
nand U13028 (N_13028,N_11389,N_12116);
or U13029 (N_13029,N_11256,N_11667);
xor U13030 (N_13030,N_11431,N_11444);
nor U13031 (N_13031,N_12260,N_11361);
or U13032 (N_13032,N_11428,N_11722);
nand U13033 (N_13033,N_11578,N_11356);
nand U13034 (N_13034,N_12023,N_12342);
xnor U13035 (N_13035,N_12050,N_11840);
and U13036 (N_13036,N_12280,N_12167);
or U13037 (N_13037,N_12105,N_11380);
and U13038 (N_13038,N_11883,N_11473);
and U13039 (N_13039,N_11575,N_11643);
and U13040 (N_13040,N_11617,N_12453);
or U13041 (N_13041,N_12299,N_12422);
xnor U13042 (N_13042,N_12179,N_11484);
xor U13043 (N_13043,N_12288,N_11327);
xor U13044 (N_13044,N_12351,N_11304);
nor U13045 (N_13045,N_11377,N_12366);
or U13046 (N_13046,N_11874,N_11721);
and U13047 (N_13047,N_11345,N_12484);
nand U13048 (N_13048,N_11338,N_12148);
nand U13049 (N_13049,N_12135,N_11581);
xnor U13050 (N_13050,N_11767,N_12081);
nor U13051 (N_13051,N_12363,N_12156);
xor U13052 (N_13052,N_11927,N_12207);
or U13053 (N_13053,N_11612,N_12055);
xor U13054 (N_13054,N_11947,N_12017);
nand U13055 (N_13055,N_12375,N_11718);
and U13056 (N_13056,N_12000,N_11326);
xnor U13057 (N_13057,N_12275,N_11733);
xor U13058 (N_13058,N_12315,N_11989);
xor U13059 (N_13059,N_12403,N_12415);
nand U13060 (N_13060,N_11755,N_11557);
nor U13061 (N_13061,N_11539,N_11352);
xnor U13062 (N_13062,N_11591,N_11743);
xnor U13063 (N_13063,N_12007,N_11474);
and U13064 (N_13064,N_11845,N_12276);
nand U13065 (N_13065,N_11500,N_11290);
or U13066 (N_13066,N_11465,N_12095);
xor U13067 (N_13067,N_11391,N_12266);
and U13068 (N_13068,N_11526,N_11648);
xnor U13069 (N_13069,N_11503,N_12356);
nand U13070 (N_13070,N_11975,N_11253);
nor U13071 (N_13071,N_12479,N_12232);
or U13072 (N_13072,N_11808,N_11731);
nor U13073 (N_13073,N_12020,N_11409);
xnor U13074 (N_13074,N_12069,N_11545);
nor U13075 (N_13075,N_11599,N_12104);
nor U13076 (N_13076,N_12263,N_11950);
nand U13077 (N_13077,N_11390,N_11404);
nand U13078 (N_13078,N_11900,N_11662);
nand U13079 (N_13079,N_11788,N_12241);
or U13080 (N_13080,N_12370,N_11976);
xor U13081 (N_13081,N_11556,N_12086);
nor U13082 (N_13082,N_12287,N_12251);
nor U13083 (N_13083,N_11673,N_12077);
or U13084 (N_13084,N_11348,N_11319);
or U13085 (N_13085,N_11459,N_11379);
nand U13086 (N_13086,N_12384,N_12301);
or U13087 (N_13087,N_12170,N_11347);
and U13088 (N_13088,N_12053,N_12218);
and U13089 (N_13089,N_12392,N_12246);
or U13090 (N_13090,N_11543,N_12063);
xnor U13091 (N_13091,N_11631,N_11491);
or U13092 (N_13092,N_12090,N_12394);
nand U13093 (N_13093,N_11334,N_11942);
nand U13094 (N_13094,N_11945,N_11933);
or U13095 (N_13095,N_11698,N_11496);
nand U13096 (N_13096,N_11967,N_12082);
or U13097 (N_13097,N_11328,N_12335);
and U13098 (N_13098,N_11899,N_11311);
xnor U13099 (N_13099,N_11402,N_11829);
and U13100 (N_13100,N_11656,N_12060);
and U13101 (N_13101,N_12278,N_11388);
nor U13102 (N_13102,N_12054,N_11654);
and U13103 (N_13103,N_11470,N_11787);
or U13104 (N_13104,N_12173,N_11855);
nor U13105 (N_13105,N_11509,N_12011);
xnor U13106 (N_13106,N_12481,N_11546);
or U13107 (N_13107,N_11717,N_12089);
nand U13108 (N_13108,N_11984,N_11309);
xor U13109 (N_13109,N_11310,N_12159);
nor U13110 (N_13110,N_12004,N_11878);
xnor U13111 (N_13111,N_11696,N_11437);
nor U13112 (N_13112,N_11816,N_11510);
nor U13113 (N_13113,N_11744,N_11675);
xnor U13114 (N_13114,N_11393,N_12003);
nor U13115 (N_13115,N_11541,N_12427);
nor U13116 (N_13116,N_11994,N_11893);
or U13117 (N_13117,N_11853,N_11937);
xor U13118 (N_13118,N_11849,N_11630);
nor U13119 (N_13119,N_11956,N_12239);
nand U13120 (N_13120,N_11985,N_12364);
and U13121 (N_13121,N_12047,N_11915);
nand U13122 (N_13122,N_12168,N_11499);
or U13123 (N_13123,N_12200,N_11647);
or U13124 (N_13124,N_11926,N_11707);
or U13125 (N_13125,N_12016,N_11619);
xnor U13126 (N_13126,N_11419,N_11441);
nor U13127 (N_13127,N_11407,N_11500);
nand U13128 (N_13128,N_12279,N_12281);
or U13129 (N_13129,N_11951,N_12306);
xnor U13130 (N_13130,N_11801,N_11407);
or U13131 (N_13131,N_11712,N_11658);
or U13132 (N_13132,N_11479,N_11506);
nor U13133 (N_13133,N_11304,N_11888);
or U13134 (N_13134,N_11546,N_12060);
and U13135 (N_13135,N_11675,N_11473);
nand U13136 (N_13136,N_12418,N_12254);
nand U13137 (N_13137,N_12337,N_11429);
and U13138 (N_13138,N_11762,N_11250);
and U13139 (N_13139,N_11826,N_11545);
and U13140 (N_13140,N_11325,N_12468);
or U13141 (N_13141,N_11793,N_11693);
nand U13142 (N_13142,N_12473,N_12442);
nor U13143 (N_13143,N_11944,N_11994);
nor U13144 (N_13144,N_12402,N_11535);
and U13145 (N_13145,N_11494,N_12493);
xor U13146 (N_13146,N_11346,N_11739);
nor U13147 (N_13147,N_11676,N_11916);
and U13148 (N_13148,N_12287,N_12246);
xnor U13149 (N_13149,N_12137,N_12482);
and U13150 (N_13150,N_11442,N_11881);
and U13151 (N_13151,N_11856,N_12092);
or U13152 (N_13152,N_11877,N_11724);
xor U13153 (N_13153,N_11668,N_11951);
xnor U13154 (N_13154,N_12016,N_11605);
nor U13155 (N_13155,N_12359,N_12047);
nor U13156 (N_13156,N_11259,N_12060);
and U13157 (N_13157,N_12287,N_11905);
xnor U13158 (N_13158,N_12096,N_12341);
and U13159 (N_13159,N_11689,N_12146);
or U13160 (N_13160,N_11558,N_11905);
nor U13161 (N_13161,N_11882,N_12348);
nand U13162 (N_13162,N_11897,N_11504);
and U13163 (N_13163,N_11465,N_11441);
nor U13164 (N_13164,N_12103,N_12437);
xor U13165 (N_13165,N_11391,N_11263);
nand U13166 (N_13166,N_12014,N_11635);
xor U13167 (N_13167,N_12303,N_12347);
and U13168 (N_13168,N_12160,N_12086);
and U13169 (N_13169,N_11720,N_11790);
xnor U13170 (N_13170,N_11695,N_11563);
or U13171 (N_13171,N_11977,N_11635);
nand U13172 (N_13172,N_11699,N_11301);
xnor U13173 (N_13173,N_12358,N_11443);
or U13174 (N_13174,N_12084,N_11339);
and U13175 (N_13175,N_12461,N_11632);
or U13176 (N_13176,N_11522,N_12363);
or U13177 (N_13177,N_11762,N_11823);
or U13178 (N_13178,N_12031,N_11627);
xnor U13179 (N_13179,N_11931,N_11298);
xnor U13180 (N_13180,N_11575,N_11533);
and U13181 (N_13181,N_12279,N_12423);
or U13182 (N_13182,N_11538,N_12079);
nand U13183 (N_13183,N_12307,N_12182);
xor U13184 (N_13184,N_12276,N_11326);
nor U13185 (N_13185,N_11562,N_11444);
nor U13186 (N_13186,N_11379,N_12239);
nor U13187 (N_13187,N_11992,N_12152);
or U13188 (N_13188,N_11539,N_12087);
and U13189 (N_13189,N_11716,N_11574);
nor U13190 (N_13190,N_12458,N_11824);
nand U13191 (N_13191,N_12303,N_12065);
xor U13192 (N_13192,N_12019,N_12079);
nor U13193 (N_13193,N_11800,N_12327);
nor U13194 (N_13194,N_11817,N_11371);
nand U13195 (N_13195,N_12151,N_12471);
xor U13196 (N_13196,N_11849,N_12376);
and U13197 (N_13197,N_11437,N_11717);
xor U13198 (N_13198,N_11838,N_11954);
nor U13199 (N_13199,N_11650,N_11614);
and U13200 (N_13200,N_12256,N_11450);
xnor U13201 (N_13201,N_11288,N_11417);
and U13202 (N_13202,N_12300,N_12350);
and U13203 (N_13203,N_11726,N_12076);
xnor U13204 (N_13204,N_11436,N_12343);
xnor U13205 (N_13205,N_11929,N_12176);
xnor U13206 (N_13206,N_12213,N_11582);
or U13207 (N_13207,N_12457,N_11278);
xnor U13208 (N_13208,N_12339,N_11683);
and U13209 (N_13209,N_11619,N_12490);
nor U13210 (N_13210,N_11761,N_11839);
and U13211 (N_13211,N_11687,N_11423);
xor U13212 (N_13212,N_11533,N_11898);
xnor U13213 (N_13213,N_11698,N_11260);
nor U13214 (N_13214,N_12405,N_12122);
nand U13215 (N_13215,N_11736,N_11252);
xor U13216 (N_13216,N_11953,N_11392);
nor U13217 (N_13217,N_12200,N_11754);
nor U13218 (N_13218,N_11963,N_12467);
nor U13219 (N_13219,N_12146,N_11428);
nor U13220 (N_13220,N_12256,N_12167);
xnor U13221 (N_13221,N_12099,N_11660);
nand U13222 (N_13222,N_11468,N_12153);
and U13223 (N_13223,N_11327,N_12042);
xnor U13224 (N_13224,N_11620,N_11340);
and U13225 (N_13225,N_12183,N_12263);
nor U13226 (N_13226,N_11581,N_11800);
and U13227 (N_13227,N_12078,N_11349);
and U13228 (N_13228,N_12483,N_12080);
xnor U13229 (N_13229,N_11692,N_12412);
and U13230 (N_13230,N_11544,N_12464);
or U13231 (N_13231,N_11378,N_12049);
or U13232 (N_13232,N_11510,N_11772);
or U13233 (N_13233,N_11258,N_11778);
and U13234 (N_13234,N_11363,N_12222);
xnor U13235 (N_13235,N_12484,N_11658);
and U13236 (N_13236,N_12445,N_11393);
or U13237 (N_13237,N_11951,N_12262);
xor U13238 (N_13238,N_11295,N_11763);
xor U13239 (N_13239,N_11656,N_12007);
and U13240 (N_13240,N_11525,N_12177);
and U13241 (N_13241,N_11942,N_11382);
and U13242 (N_13242,N_12281,N_11833);
and U13243 (N_13243,N_12024,N_12128);
xnor U13244 (N_13244,N_12365,N_12400);
nand U13245 (N_13245,N_12354,N_11546);
or U13246 (N_13246,N_12407,N_11824);
or U13247 (N_13247,N_11808,N_11807);
xnor U13248 (N_13248,N_12329,N_11666);
nand U13249 (N_13249,N_11351,N_12280);
and U13250 (N_13250,N_12481,N_11985);
nor U13251 (N_13251,N_11808,N_11604);
nand U13252 (N_13252,N_12260,N_11785);
nand U13253 (N_13253,N_11380,N_11337);
and U13254 (N_13254,N_11768,N_11476);
xnor U13255 (N_13255,N_12199,N_11352);
and U13256 (N_13256,N_12224,N_12362);
and U13257 (N_13257,N_12087,N_11988);
and U13258 (N_13258,N_12189,N_12149);
and U13259 (N_13259,N_11692,N_12068);
nand U13260 (N_13260,N_11336,N_11405);
nor U13261 (N_13261,N_11401,N_11490);
nand U13262 (N_13262,N_12418,N_11522);
xnor U13263 (N_13263,N_12476,N_11787);
xnor U13264 (N_13264,N_12299,N_12262);
xnor U13265 (N_13265,N_11391,N_11280);
nor U13266 (N_13266,N_12102,N_12033);
xor U13267 (N_13267,N_12131,N_12005);
xor U13268 (N_13268,N_11675,N_11490);
nor U13269 (N_13269,N_11985,N_12243);
nor U13270 (N_13270,N_12322,N_11939);
nor U13271 (N_13271,N_12359,N_11694);
or U13272 (N_13272,N_11977,N_11736);
nor U13273 (N_13273,N_12093,N_11621);
nand U13274 (N_13274,N_12176,N_12222);
nand U13275 (N_13275,N_11966,N_12194);
or U13276 (N_13276,N_11931,N_11370);
or U13277 (N_13277,N_12484,N_11588);
xor U13278 (N_13278,N_11405,N_11986);
and U13279 (N_13279,N_11672,N_12276);
nand U13280 (N_13280,N_11550,N_11948);
nor U13281 (N_13281,N_12019,N_11687);
xnor U13282 (N_13282,N_12321,N_12342);
nor U13283 (N_13283,N_11879,N_12065);
nor U13284 (N_13284,N_12393,N_11260);
and U13285 (N_13285,N_11367,N_12267);
and U13286 (N_13286,N_12437,N_11650);
xor U13287 (N_13287,N_12303,N_11493);
or U13288 (N_13288,N_11864,N_11866);
xnor U13289 (N_13289,N_11424,N_12332);
and U13290 (N_13290,N_12380,N_11489);
nand U13291 (N_13291,N_12391,N_11328);
or U13292 (N_13292,N_12014,N_11741);
and U13293 (N_13293,N_12004,N_12450);
or U13294 (N_13294,N_11532,N_12385);
or U13295 (N_13295,N_12056,N_11716);
nand U13296 (N_13296,N_12197,N_11322);
and U13297 (N_13297,N_12136,N_11321);
or U13298 (N_13298,N_11996,N_11526);
xnor U13299 (N_13299,N_12269,N_11477);
nor U13300 (N_13300,N_11683,N_11651);
and U13301 (N_13301,N_11466,N_12000);
nand U13302 (N_13302,N_11309,N_12248);
xor U13303 (N_13303,N_11781,N_12125);
nor U13304 (N_13304,N_11845,N_11473);
and U13305 (N_13305,N_11905,N_12058);
nor U13306 (N_13306,N_11819,N_11315);
nand U13307 (N_13307,N_11801,N_11572);
xor U13308 (N_13308,N_12117,N_12197);
nand U13309 (N_13309,N_12117,N_11302);
or U13310 (N_13310,N_11921,N_12462);
or U13311 (N_13311,N_12224,N_12283);
xor U13312 (N_13312,N_12404,N_11392);
nand U13313 (N_13313,N_11254,N_11542);
nor U13314 (N_13314,N_11810,N_12313);
nor U13315 (N_13315,N_11796,N_12279);
xor U13316 (N_13316,N_12421,N_11926);
xor U13317 (N_13317,N_12298,N_12465);
xor U13318 (N_13318,N_11873,N_11331);
or U13319 (N_13319,N_11424,N_12039);
and U13320 (N_13320,N_11947,N_11441);
and U13321 (N_13321,N_11635,N_11601);
nand U13322 (N_13322,N_11671,N_12424);
nor U13323 (N_13323,N_11834,N_11921);
xnor U13324 (N_13324,N_12092,N_11608);
or U13325 (N_13325,N_11382,N_11784);
and U13326 (N_13326,N_11702,N_11656);
nand U13327 (N_13327,N_11819,N_11996);
xnor U13328 (N_13328,N_11963,N_12164);
and U13329 (N_13329,N_11671,N_12002);
and U13330 (N_13330,N_12215,N_11427);
and U13331 (N_13331,N_12469,N_11289);
xor U13332 (N_13332,N_12309,N_12317);
nand U13333 (N_13333,N_12433,N_11704);
xor U13334 (N_13334,N_11685,N_12100);
or U13335 (N_13335,N_11324,N_11473);
nor U13336 (N_13336,N_11534,N_11683);
or U13337 (N_13337,N_11546,N_12325);
nor U13338 (N_13338,N_12077,N_11661);
or U13339 (N_13339,N_11548,N_12452);
or U13340 (N_13340,N_11984,N_12266);
or U13341 (N_13341,N_12023,N_12179);
nand U13342 (N_13342,N_11927,N_12107);
and U13343 (N_13343,N_12064,N_11766);
and U13344 (N_13344,N_11448,N_12178);
xor U13345 (N_13345,N_11522,N_12045);
xnor U13346 (N_13346,N_11897,N_12397);
or U13347 (N_13347,N_12499,N_11729);
nand U13348 (N_13348,N_12281,N_12066);
and U13349 (N_13349,N_12139,N_12041);
or U13350 (N_13350,N_12399,N_12306);
xor U13351 (N_13351,N_11637,N_12328);
nor U13352 (N_13352,N_11300,N_12070);
and U13353 (N_13353,N_11846,N_11333);
or U13354 (N_13354,N_12362,N_12370);
and U13355 (N_13355,N_11811,N_12463);
and U13356 (N_13356,N_11633,N_12374);
nand U13357 (N_13357,N_12289,N_12027);
xor U13358 (N_13358,N_11848,N_11967);
and U13359 (N_13359,N_12048,N_12226);
or U13360 (N_13360,N_11840,N_11731);
and U13361 (N_13361,N_12240,N_11322);
and U13362 (N_13362,N_12198,N_12283);
nand U13363 (N_13363,N_11748,N_11415);
nor U13364 (N_13364,N_12056,N_11743);
or U13365 (N_13365,N_11661,N_11611);
nand U13366 (N_13366,N_12156,N_12016);
nand U13367 (N_13367,N_11723,N_12001);
or U13368 (N_13368,N_12046,N_11989);
or U13369 (N_13369,N_11661,N_11311);
and U13370 (N_13370,N_12485,N_12462);
or U13371 (N_13371,N_11989,N_12194);
or U13372 (N_13372,N_11556,N_11463);
nand U13373 (N_13373,N_11750,N_11553);
and U13374 (N_13374,N_11573,N_11931);
and U13375 (N_13375,N_11362,N_11763);
nand U13376 (N_13376,N_11583,N_11324);
or U13377 (N_13377,N_11712,N_11259);
or U13378 (N_13378,N_12151,N_11633);
or U13379 (N_13379,N_12143,N_12489);
nand U13380 (N_13380,N_12148,N_11287);
nand U13381 (N_13381,N_12133,N_11583);
xnor U13382 (N_13382,N_12400,N_12118);
nand U13383 (N_13383,N_11272,N_11654);
xor U13384 (N_13384,N_11264,N_12115);
or U13385 (N_13385,N_11390,N_12152);
or U13386 (N_13386,N_12139,N_11901);
or U13387 (N_13387,N_11768,N_11533);
and U13388 (N_13388,N_12371,N_12415);
nor U13389 (N_13389,N_11413,N_11593);
nor U13390 (N_13390,N_12421,N_11826);
and U13391 (N_13391,N_11488,N_12146);
nor U13392 (N_13392,N_12103,N_12252);
nor U13393 (N_13393,N_12059,N_11286);
xnor U13394 (N_13394,N_11490,N_11448);
nand U13395 (N_13395,N_11640,N_11578);
and U13396 (N_13396,N_11659,N_12448);
or U13397 (N_13397,N_12132,N_11854);
or U13398 (N_13398,N_11456,N_11510);
or U13399 (N_13399,N_12146,N_11792);
and U13400 (N_13400,N_12011,N_12481);
or U13401 (N_13401,N_12149,N_11974);
or U13402 (N_13402,N_12077,N_11690);
nor U13403 (N_13403,N_12132,N_12233);
xnor U13404 (N_13404,N_12378,N_11577);
nor U13405 (N_13405,N_12400,N_11518);
nor U13406 (N_13406,N_11361,N_11499);
or U13407 (N_13407,N_11601,N_12110);
xnor U13408 (N_13408,N_12243,N_11846);
nor U13409 (N_13409,N_11761,N_11752);
xnor U13410 (N_13410,N_12428,N_11943);
xor U13411 (N_13411,N_11443,N_12171);
and U13412 (N_13412,N_12302,N_11804);
and U13413 (N_13413,N_11433,N_11509);
and U13414 (N_13414,N_11447,N_11588);
nand U13415 (N_13415,N_12084,N_11896);
and U13416 (N_13416,N_11748,N_12141);
and U13417 (N_13417,N_11851,N_11451);
nand U13418 (N_13418,N_11725,N_11387);
and U13419 (N_13419,N_12404,N_11927);
or U13420 (N_13420,N_12413,N_12120);
or U13421 (N_13421,N_11932,N_11439);
nor U13422 (N_13422,N_12453,N_12078);
nand U13423 (N_13423,N_12499,N_11452);
or U13424 (N_13424,N_11594,N_11342);
nand U13425 (N_13425,N_11514,N_11568);
and U13426 (N_13426,N_11296,N_11682);
and U13427 (N_13427,N_11645,N_11995);
nand U13428 (N_13428,N_11690,N_12373);
or U13429 (N_13429,N_11820,N_12274);
or U13430 (N_13430,N_11302,N_11265);
or U13431 (N_13431,N_11585,N_12480);
and U13432 (N_13432,N_12366,N_12338);
and U13433 (N_13433,N_11280,N_12087);
nor U13434 (N_13434,N_12117,N_11256);
and U13435 (N_13435,N_12086,N_12194);
xor U13436 (N_13436,N_11692,N_12045);
and U13437 (N_13437,N_11385,N_12106);
or U13438 (N_13438,N_12110,N_11642);
nor U13439 (N_13439,N_11894,N_11962);
nor U13440 (N_13440,N_12468,N_11740);
or U13441 (N_13441,N_12442,N_11692);
nand U13442 (N_13442,N_11300,N_11588);
and U13443 (N_13443,N_11460,N_11988);
and U13444 (N_13444,N_11842,N_12491);
nand U13445 (N_13445,N_12310,N_12206);
or U13446 (N_13446,N_12141,N_12107);
or U13447 (N_13447,N_12031,N_11623);
nand U13448 (N_13448,N_11342,N_11486);
nor U13449 (N_13449,N_12439,N_12248);
nor U13450 (N_13450,N_11567,N_11640);
or U13451 (N_13451,N_12438,N_11569);
xnor U13452 (N_13452,N_11449,N_11332);
nand U13453 (N_13453,N_11799,N_11439);
nor U13454 (N_13454,N_11812,N_12306);
and U13455 (N_13455,N_11681,N_12460);
nand U13456 (N_13456,N_11414,N_11647);
and U13457 (N_13457,N_11857,N_11440);
xor U13458 (N_13458,N_12382,N_11416);
xnor U13459 (N_13459,N_12277,N_11587);
nand U13460 (N_13460,N_11286,N_12013);
and U13461 (N_13461,N_11359,N_11597);
and U13462 (N_13462,N_11295,N_11258);
or U13463 (N_13463,N_12077,N_12430);
nand U13464 (N_13464,N_12286,N_12486);
and U13465 (N_13465,N_11485,N_11569);
xor U13466 (N_13466,N_11711,N_12469);
nor U13467 (N_13467,N_11961,N_11444);
and U13468 (N_13468,N_12202,N_11380);
or U13469 (N_13469,N_12336,N_12008);
xnor U13470 (N_13470,N_11730,N_11312);
xor U13471 (N_13471,N_12372,N_11259);
nand U13472 (N_13472,N_12117,N_11575);
xnor U13473 (N_13473,N_12193,N_12316);
or U13474 (N_13474,N_12157,N_11686);
nor U13475 (N_13475,N_12150,N_12031);
or U13476 (N_13476,N_11879,N_12454);
and U13477 (N_13477,N_11976,N_11700);
and U13478 (N_13478,N_12046,N_11688);
and U13479 (N_13479,N_11469,N_11913);
or U13480 (N_13480,N_12038,N_11531);
xor U13481 (N_13481,N_11916,N_11685);
nor U13482 (N_13482,N_11322,N_12217);
xor U13483 (N_13483,N_11325,N_11746);
or U13484 (N_13484,N_11846,N_11679);
nor U13485 (N_13485,N_11778,N_11418);
and U13486 (N_13486,N_11715,N_11487);
nor U13487 (N_13487,N_11980,N_12173);
or U13488 (N_13488,N_11825,N_11926);
nor U13489 (N_13489,N_11736,N_12458);
and U13490 (N_13490,N_11409,N_12173);
or U13491 (N_13491,N_12449,N_12030);
and U13492 (N_13492,N_12197,N_12057);
and U13493 (N_13493,N_11611,N_11935);
nand U13494 (N_13494,N_12444,N_11855);
nand U13495 (N_13495,N_11280,N_11889);
xnor U13496 (N_13496,N_11660,N_12017);
nor U13497 (N_13497,N_12195,N_12280);
nand U13498 (N_13498,N_12187,N_12248);
xnor U13499 (N_13499,N_12386,N_11799);
nand U13500 (N_13500,N_11736,N_12032);
or U13501 (N_13501,N_12260,N_12144);
xnor U13502 (N_13502,N_11380,N_11481);
xnor U13503 (N_13503,N_11820,N_12466);
or U13504 (N_13504,N_11766,N_11372);
and U13505 (N_13505,N_11817,N_11476);
nor U13506 (N_13506,N_12337,N_11455);
xnor U13507 (N_13507,N_11286,N_12143);
or U13508 (N_13508,N_11306,N_11877);
nor U13509 (N_13509,N_12309,N_11627);
and U13510 (N_13510,N_12237,N_11459);
nand U13511 (N_13511,N_11496,N_11611);
or U13512 (N_13512,N_11276,N_11814);
nand U13513 (N_13513,N_11434,N_12388);
nand U13514 (N_13514,N_11733,N_11942);
and U13515 (N_13515,N_12028,N_11326);
nand U13516 (N_13516,N_12419,N_12489);
and U13517 (N_13517,N_12396,N_11537);
and U13518 (N_13518,N_11598,N_12386);
xor U13519 (N_13519,N_11808,N_11929);
nor U13520 (N_13520,N_11398,N_11412);
xor U13521 (N_13521,N_11544,N_11555);
and U13522 (N_13522,N_11863,N_11527);
nor U13523 (N_13523,N_12070,N_12312);
xor U13524 (N_13524,N_12449,N_12348);
or U13525 (N_13525,N_11967,N_12450);
nand U13526 (N_13526,N_12299,N_12015);
nand U13527 (N_13527,N_11554,N_11610);
or U13528 (N_13528,N_11279,N_11679);
xor U13529 (N_13529,N_12022,N_11345);
nor U13530 (N_13530,N_12152,N_11502);
nand U13531 (N_13531,N_11791,N_11927);
nor U13532 (N_13532,N_12399,N_12249);
xnor U13533 (N_13533,N_12270,N_11524);
and U13534 (N_13534,N_12487,N_11486);
or U13535 (N_13535,N_11856,N_11913);
and U13536 (N_13536,N_12416,N_11771);
or U13537 (N_13537,N_11366,N_12031);
and U13538 (N_13538,N_11712,N_12058);
or U13539 (N_13539,N_12465,N_11948);
nand U13540 (N_13540,N_11436,N_11893);
xnor U13541 (N_13541,N_12346,N_11681);
nand U13542 (N_13542,N_11843,N_11706);
nor U13543 (N_13543,N_11560,N_11552);
xor U13544 (N_13544,N_11449,N_12061);
nor U13545 (N_13545,N_11652,N_11595);
nand U13546 (N_13546,N_11809,N_11556);
nor U13547 (N_13547,N_11378,N_12148);
xor U13548 (N_13548,N_11753,N_11939);
nor U13549 (N_13549,N_11797,N_11833);
nand U13550 (N_13550,N_12227,N_12493);
nor U13551 (N_13551,N_12153,N_11745);
or U13552 (N_13552,N_11705,N_12206);
or U13553 (N_13553,N_11865,N_11382);
nor U13554 (N_13554,N_12218,N_12485);
or U13555 (N_13555,N_11750,N_12142);
nor U13556 (N_13556,N_11618,N_11279);
xor U13557 (N_13557,N_12013,N_12453);
nand U13558 (N_13558,N_11560,N_12126);
nor U13559 (N_13559,N_11631,N_12476);
nand U13560 (N_13560,N_11936,N_11676);
or U13561 (N_13561,N_11337,N_11339);
and U13562 (N_13562,N_11460,N_11841);
xor U13563 (N_13563,N_11769,N_12089);
and U13564 (N_13564,N_12298,N_11503);
nand U13565 (N_13565,N_12240,N_12262);
nor U13566 (N_13566,N_11436,N_12390);
and U13567 (N_13567,N_12125,N_12298);
nand U13568 (N_13568,N_11373,N_11498);
nand U13569 (N_13569,N_11735,N_11610);
and U13570 (N_13570,N_11445,N_11911);
nor U13571 (N_13571,N_11726,N_11342);
nor U13572 (N_13572,N_12456,N_12232);
or U13573 (N_13573,N_11272,N_12461);
and U13574 (N_13574,N_11618,N_12468);
xor U13575 (N_13575,N_11814,N_12467);
nand U13576 (N_13576,N_11483,N_11528);
nand U13577 (N_13577,N_12420,N_11909);
nor U13578 (N_13578,N_12466,N_11595);
or U13579 (N_13579,N_11826,N_12269);
and U13580 (N_13580,N_12354,N_11355);
nor U13581 (N_13581,N_11510,N_11904);
xnor U13582 (N_13582,N_12474,N_12204);
xnor U13583 (N_13583,N_11459,N_12327);
and U13584 (N_13584,N_11319,N_11838);
and U13585 (N_13585,N_11983,N_11954);
nor U13586 (N_13586,N_11999,N_12446);
nor U13587 (N_13587,N_12115,N_11918);
nor U13588 (N_13588,N_11943,N_11963);
or U13589 (N_13589,N_11489,N_12362);
nand U13590 (N_13590,N_11439,N_12257);
and U13591 (N_13591,N_12074,N_12177);
nor U13592 (N_13592,N_12163,N_11907);
xor U13593 (N_13593,N_12398,N_11890);
nor U13594 (N_13594,N_11971,N_11644);
xnor U13595 (N_13595,N_11836,N_11458);
or U13596 (N_13596,N_11782,N_12480);
nand U13597 (N_13597,N_11845,N_11697);
nand U13598 (N_13598,N_12200,N_12334);
nand U13599 (N_13599,N_12338,N_11728);
nor U13600 (N_13600,N_12305,N_11704);
or U13601 (N_13601,N_11410,N_11906);
nand U13602 (N_13602,N_12272,N_11904);
nor U13603 (N_13603,N_11397,N_11943);
and U13604 (N_13604,N_12306,N_11409);
xnor U13605 (N_13605,N_11824,N_12479);
xnor U13606 (N_13606,N_11612,N_11488);
xnor U13607 (N_13607,N_11602,N_11825);
or U13608 (N_13608,N_12306,N_12003);
or U13609 (N_13609,N_11416,N_11670);
xor U13610 (N_13610,N_11498,N_12145);
xnor U13611 (N_13611,N_11894,N_11840);
xnor U13612 (N_13612,N_11711,N_11892);
nand U13613 (N_13613,N_12043,N_11592);
or U13614 (N_13614,N_11868,N_11311);
or U13615 (N_13615,N_11731,N_11967);
xnor U13616 (N_13616,N_12396,N_11846);
xnor U13617 (N_13617,N_11618,N_11903);
nor U13618 (N_13618,N_11914,N_12168);
and U13619 (N_13619,N_11936,N_11967);
xnor U13620 (N_13620,N_12279,N_12321);
and U13621 (N_13621,N_11574,N_11874);
nor U13622 (N_13622,N_11738,N_11572);
nor U13623 (N_13623,N_11535,N_11984);
nor U13624 (N_13624,N_11804,N_11449);
and U13625 (N_13625,N_12410,N_12169);
nor U13626 (N_13626,N_11278,N_11319);
and U13627 (N_13627,N_12390,N_12328);
or U13628 (N_13628,N_11570,N_11644);
nand U13629 (N_13629,N_11798,N_11556);
or U13630 (N_13630,N_12018,N_11271);
and U13631 (N_13631,N_11882,N_11595);
and U13632 (N_13632,N_11454,N_11613);
and U13633 (N_13633,N_11542,N_12070);
and U13634 (N_13634,N_11993,N_11802);
or U13635 (N_13635,N_11744,N_12323);
or U13636 (N_13636,N_11878,N_11869);
nand U13637 (N_13637,N_11884,N_12196);
xor U13638 (N_13638,N_12052,N_11345);
nor U13639 (N_13639,N_12451,N_12051);
or U13640 (N_13640,N_12218,N_11633);
nand U13641 (N_13641,N_11382,N_11391);
and U13642 (N_13642,N_11857,N_11808);
nand U13643 (N_13643,N_11914,N_12194);
nor U13644 (N_13644,N_12240,N_11581);
and U13645 (N_13645,N_11566,N_12065);
nand U13646 (N_13646,N_11435,N_11531);
xnor U13647 (N_13647,N_11874,N_11671);
nand U13648 (N_13648,N_11915,N_12459);
xnor U13649 (N_13649,N_11753,N_11309);
xnor U13650 (N_13650,N_11589,N_12303);
and U13651 (N_13651,N_11485,N_11436);
or U13652 (N_13652,N_11336,N_11438);
xnor U13653 (N_13653,N_11918,N_11509);
or U13654 (N_13654,N_12123,N_12111);
nand U13655 (N_13655,N_11510,N_11761);
and U13656 (N_13656,N_11983,N_12364);
and U13657 (N_13657,N_12154,N_11828);
nand U13658 (N_13658,N_11471,N_11926);
nand U13659 (N_13659,N_12479,N_12452);
or U13660 (N_13660,N_11893,N_11395);
nor U13661 (N_13661,N_11717,N_12480);
and U13662 (N_13662,N_11323,N_11396);
xor U13663 (N_13663,N_11456,N_11526);
and U13664 (N_13664,N_11340,N_12050);
xor U13665 (N_13665,N_12118,N_11907);
xor U13666 (N_13666,N_11341,N_12410);
or U13667 (N_13667,N_11927,N_11274);
xnor U13668 (N_13668,N_12431,N_12116);
xnor U13669 (N_13669,N_11723,N_12334);
nor U13670 (N_13670,N_12116,N_11927);
nor U13671 (N_13671,N_12470,N_11931);
or U13672 (N_13672,N_11750,N_11960);
or U13673 (N_13673,N_11404,N_12013);
nand U13674 (N_13674,N_12172,N_12166);
nor U13675 (N_13675,N_11399,N_11578);
or U13676 (N_13676,N_12149,N_12148);
nor U13677 (N_13677,N_11495,N_12257);
and U13678 (N_13678,N_11251,N_11266);
xnor U13679 (N_13679,N_11976,N_12379);
and U13680 (N_13680,N_12133,N_11504);
nor U13681 (N_13681,N_11772,N_11385);
xnor U13682 (N_13682,N_12340,N_11838);
or U13683 (N_13683,N_12436,N_11589);
and U13684 (N_13684,N_12352,N_11904);
xnor U13685 (N_13685,N_11381,N_11936);
or U13686 (N_13686,N_12288,N_11904);
nand U13687 (N_13687,N_11771,N_11853);
and U13688 (N_13688,N_11335,N_12333);
or U13689 (N_13689,N_11992,N_11331);
nor U13690 (N_13690,N_12384,N_11717);
nor U13691 (N_13691,N_11656,N_11265);
and U13692 (N_13692,N_11360,N_12077);
nor U13693 (N_13693,N_12095,N_11909);
xor U13694 (N_13694,N_11478,N_11929);
nor U13695 (N_13695,N_11722,N_11277);
xor U13696 (N_13696,N_12103,N_12070);
xnor U13697 (N_13697,N_11808,N_12435);
or U13698 (N_13698,N_11296,N_12153);
nand U13699 (N_13699,N_12153,N_12413);
or U13700 (N_13700,N_11850,N_11341);
xor U13701 (N_13701,N_12359,N_11427);
and U13702 (N_13702,N_12293,N_12367);
nand U13703 (N_13703,N_11691,N_11435);
nand U13704 (N_13704,N_12395,N_12033);
nand U13705 (N_13705,N_11258,N_11688);
or U13706 (N_13706,N_11386,N_11902);
nor U13707 (N_13707,N_11657,N_11661);
and U13708 (N_13708,N_11729,N_11826);
and U13709 (N_13709,N_11960,N_12492);
nand U13710 (N_13710,N_11499,N_11416);
nand U13711 (N_13711,N_11648,N_11915);
nor U13712 (N_13712,N_11435,N_12172);
or U13713 (N_13713,N_12025,N_12239);
or U13714 (N_13714,N_11866,N_11332);
or U13715 (N_13715,N_12282,N_12489);
nor U13716 (N_13716,N_12036,N_12395);
nand U13717 (N_13717,N_12268,N_11698);
xor U13718 (N_13718,N_12038,N_11980);
and U13719 (N_13719,N_11603,N_12080);
or U13720 (N_13720,N_11553,N_12107);
nor U13721 (N_13721,N_11772,N_11764);
nand U13722 (N_13722,N_11572,N_11632);
or U13723 (N_13723,N_11534,N_11941);
or U13724 (N_13724,N_12321,N_12099);
nor U13725 (N_13725,N_11384,N_11845);
xnor U13726 (N_13726,N_12329,N_11333);
xor U13727 (N_13727,N_12187,N_11573);
xnor U13728 (N_13728,N_11951,N_11626);
and U13729 (N_13729,N_12436,N_12453);
xnor U13730 (N_13730,N_12203,N_11780);
nor U13731 (N_13731,N_11612,N_11720);
nand U13732 (N_13732,N_11272,N_11918);
nor U13733 (N_13733,N_11420,N_12277);
nor U13734 (N_13734,N_11623,N_12275);
and U13735 (N_13735,N_11284,N_11926);
and U13736 (N_13736,N_11815,N_12093);
xor U13737 (N_13737,N_12261,N_12410);
and U13738 (N_13738,N_11349,N_11945);
nand U13739 (N_13739,N_12129,N_11337);
xnor U13740 (N_13740,N_11284,N_11814);
and U13741 (N_13741,N_12350,N_12295);
and U13742 (N_13742,N_11890,N_11704);
xnor U13743 (N_13743,N_11352,N_12487);
xnor U13744 (N_13744,N_11812,N_11831);
and U13745 (N_13745,N_12285,N_12253);
nand U13746 (N_13746,N_11542,N_12215);
or U13747 (N_13747,N_11435,N_11670);
nand U13748 (N_13748,N_11761,N_12200);
nor U13749 (N_13749,N_11818,N_11830);
nor U13750 (N_13750,N_13480,N_13150);
nand U13751 (N_13751,N_12641,N_13092);
nor U13752 (N_13752,N_12747,N_12524);
xor U13753 (N_13753,N_13327,N_13069);
or U13754 (N_13754,N_12781,N_13559);
and U13755 (N_13755,N_12975,N_12752);
xnor U13756 (N_13756,N_13739,N_13414);
xor U13757 (N_13757,N_13408,N_12736);
nand U13758 (N_13758,N_13481,N_12871);
and U13759 (N_13759,N_12814,N_13280);
xnor U13760 (N_13760,N_13415,N_13261);
nand U13761 (N_13761,N_12527,N_13484);
nor U13762 (N_13762,N_12670,N_12938);
or U13763 (N_13763,N_12679,N_13273);
xor U13764 (N_13764,N_13310,N_13749);
and U13765 (N_13765,N_13291,N_12651);
and U13766 (N_13766,N_12865,N_13726);
nor U13767 (N_13767,N_13445,N_12601);
nand U13768 (N_13768,N_13448,N_12775);
or U13769 (N_13769,N_12545,N_12903);
nor U13770 (N_13770,N_13269,N_13602);
xor U13771 (N_13771,N_13257,N_13248);
xnor U13772 (N_13772,N_13373,N_13376);
or U13773 (N_13773,N_13122,N_13637);
xnor U13774 (N_13774,N_12897,N_13178);
or U13775 (N_13775,N_13260,N_12984);
nor U13776 (N_13776,N_12932,N_12896);
nor U13777 (N_13777,N_13404,N_13125);
and U13778 (N_13778,N_13411,N_12990);
or U13779 (N_13779,N_13106,N_13645);
xor U13780 (N_13780,N_13317,N_13627);
and U13781 (N_13781,N_13501,N_13543);
nor U13782 (N_13782,N_12861,N_13278);
and U13783 (N_13783,N_12754,N_13004);
nor U13784 (N_13784,N_13532,N_12999);
nor U13785 (N_13785,N_13616,N_12866);
xnor U13786 (N_13786,N_12538,N_12839);
xor U13787 (N_13787,N_13675,N_12771);
xnor U13788 (N_13788,N_12878,N_13155);
or U13789 (N_13789,N_13416,N_12940);
nor U13790 (N_13790,N_12912,N_13427);
and U13791 (N_13791,N_12962,N_13297);
xnor U13792 (N_13792,N_13697,N_12684);
nor U13793 (N_13793,N_13518,N_13563);
or U13794 (N_13794,N_13277,N_12535);
nor U13795 (N_13795,N_13080,N_12623);
nand U13796 (N_13796,N_12842,N_12743);
nand U13797 (N_13797,N_12612,N_12846);
nor U13798 (N_13798,N_12525,N_13172);
and U13799 (N_13799,N_13499,N_12572);
nor U13800 (N_13800,N_13186,N_13288);
and U13801 (N_13801,N_13465,N_12630);
nor U13802 (N_13802,N_13275,N_13372);
xor U13803 (N_13803,N_12915,N_12616);
or U13804 (N_13804,N_12909,N_12762);
or U13805 (N_13805,N_13202,N_12926);
xnor U13806 (N_13806,N_12646,N_13265);
and U13807 (N_13807,N_12832,N_13086);
nand U13808 (N_13808,N_13459,N_13457);
nor U13809 (N_13809,N_13059,N_13422);
nor U13810 (N_13810,N_12834,N_13599);
and U13811 (N_13811,N_12959,N_12508);
nor U13812 (N_13812,N_12617,N_13068);
or U13813 (N_13813,N_13633,N_12738);
nor U13814 (N_13814,N_12979,N_13730);
nor U13815 (N_13815,N_12943,N_12677);
and U13816 (N_13816,N_12996,N_12750);
nand U13817 (N_13817,N_12674,N_13177);
xnor U13818 (N_13818,N_12580,N_12873);
or U13819 (N_13819,N_13581,N_13453);
or U13820 (N_13820,N_12886,N_13201);
xor U13821 (N_13821,N_12544,N_13168);
nor U13822 (N_13822,N_13723,N_13712);
nor U13823 (N_13823,N_13205,N_13469);
and U13824 (N_13824,N_13213,N_12960);
nand U13825 (N_13825,N_12589,N_13597);
nand U13826 (N_13826,N_13511,N_12526);
nand U13827 (N_13827,N_13164,N_12767);
xor U13828 (N_13828,N_13671,N_13340);
and U13829 (N_13829,N_12642,N_13737);
or U13830 (N_13830,N_13311,N_13742);
nor U13831 (N_13831,N_13724,N_12579);
or U13832 (N_13832,N_12735,N_13699);
xnor U13833 (N_13833,N_13466,N_13182);
or U13834 (N_13834,N_13160,N_12520);
and U13835 (N_13835,N_13234,N_13077);
nand U13836 (N_13836,N_13668,N_13074);
nand U13837 (N_13837,N_13121,N_13019);
nand U13838 (N_13838,N_12607,N_12902);
and U13839 (N_13839,N_12536,N_12561);
and U13840 (N_13840,N_12796,N_12764);
nor U13841 (N_13841,N_13323,N_13304);
nand U13842 (N_13842,N_12934,N_13272);
nand U13843 (N_13843,N_13512,N_13577);
nand U13844 (N_13844,N_13392,N_13196);
xnor U13845 (N_13845,N_13203,N_13630);
xnor U13846 (N_13846,N_13126,N_13556);
nor U13847 (N_13847,N_13364,N_13617);
and U13848 (N_13848,N_13173,N_13589);
nand U13849 (N_13849,N_13190,N_13085);
and U13850 (N_13850,N_13555,N_13104);
and U13851 (N_13851,N_13072,N_12574);
xnor U13852 (N_13852,N_12737,N_13655);
xor U13853 (N_13853,N_13442,N_12806);
xnor U13854 (N_13854,N_12748,N_13250);
and U13855 (N_13855,N_12863,N_13028);
xnor U13856 (N_13856,N_13434,N_13333);
or U13857 (N_13857,N_13266,N_13526);
nor U13858 (N_13858,N_13088,N_13281);
and U13859 (N_13859,N_13672,N_13657);
and U13860 (N_13860,N_13316,N_13390);
and U13861 (N_13861,N_12898,N_12790);
nand U13862 (N_13862,N_12560,N_12672);
and U13863 (N_13863,N_13684,N_12680);
and U13864 (N_13864,N_13594,N_13676);
nand U13865 (N_13865,N_12598,N_12779);
nor U13866 (N_13866,N_12744,N_13174);
nor U13867 (N_13867,N_13537,N_13334);
nor U13868 (N_13868,N_13216,N_13718);
xor U13869 (N_13869,N_13460,N_12826);
xnor U13870 (N_13870,N_13076,N_12660);
and U13871 (N_13871,N_12787,N_12840);
nor U13872 (N_13872,N_13063,N_12780);
or U13873 (N_13873,N_12565,N_13393);
or U13874 (N_13874,N_12869,N_12968);
and U13875 (N_13875,N_13554,N_13079);
nor U13876 (N_13876,N_13176,N_12974);
xnor U13877 (N_13877,N_12682,N_13038);
nor U13878 (N_13878,N_13349,N_13625);
and U13879 (N_13879,N_13394,N_12945);
xnor U13880 (N_13880,N_13410,N_12751);
or U13881 (N_13881,N_12914,N_12969);
nor U13882 (N_13882,N_13535,N_13097);
nor U13883 (N_13883,N_13037,N_13574);
or U13884 (N_13884,N_12860,N_12503);
xor U13885 (N_13885,N_12913,N_13325);
nor U13886 (N_13886,N_12952,N_12676);
xor U13887 (N_13887,N_13436,N_13221);
xnor U13888 (N_13888,N_13228,N_13474);
and U13889 (N_13889,N_12788,N_13306);
nand U13890 (N_13890,N_13057,N_12944);
nor U13891 (N_13891,N_13508,N_13600);
xnor U13892 (N_13892,N_12592,N_13530);
xor U13893 (N_13893,N_12685,N_13748);
nand U13894 (N_13894,N_12655,N_12883);
xnor U13895 (N_13895,N_12740,N_13175);
and U13896 (N_13896,N_13268,N_13167);
and U13897 (N_13897,N_13588,N_12824);
or U13898 (N_13898,N_13437,N_12856);
or U13899 (N_13899,N_12608,N_13255);
xnor U13900 (N_13900,N_13400,N_12681);
nor U13901 (N_13901,N_13103,N_13447);
xnor U13902 (N_13902,N_12563,N_12529);
xor U13903 (N_13903,N_12541,N_13362);
nor U13904 (N_13904,N_13720,N_12852);
or U13905 (N_13905,N_13188,N_13496);
and U13906 (N_13906,N_12837,N_12718);
nand U13907 (N_13907,N_13507,N_12605);
and U13908 (N_13908,N_13421,N_12755);
or U13909 (N_13909,N_13223,N_12858);
or U13910 (N_13910,N_12813,N_13674);
nand U13911 (N_13911,N_13598,N_12537);
or U13912 (N_13912,N_13326,N_13579);
and U13913 (N_13913,N_13263,N_12573);
xor U13914 (N_13914,N_13145,N_12910);
and U13915 (N_13915,N_12784,N_13099);
xor U13916 (N_13916,N_13307,N_12964);
or U13917 (N_13917,N_13612,N_12675);
nand U13918 (N_13918,N_12803,N_13711);
nand U13919 (N_13919,N_13383,N_12987);
xor U13920 (N_13920,N_12916,N_12733);
and U13921 (N_13921,N_13568,N_12922);
and U13922 (N_13922,N_12937,N_13045);
nor U13923 (N_13923,N_12864,N_13536);
or U13924 (N_13924,N_12827,N_12844);
xnor U13925 (N_13925,N_13519,N_12719);
nand U13926 (N_13926,N_12804,N_13485);
nor U13927 (N_13927,N_13418,N_13386);
or U13928 (N_13928,N_13267,N_13032);
or U13929 (N_13929,N_13331,N_13198);
and U13930 (N_13930,N_13565,N_12627);
xor U13931 (N_13931,N_12568,N_13653);
or U13932 (N_13932,N_13670,N_13603);
nor U13933 (N_13933,N_12638,N_13271);
nand U13934 (N_13934,N_12625,N_13232);
xor U13935 (N_13935,N_12518,N_13450);
and U13936 (N_13936,N_12724,N_13135);
xor U13937 (N_13937,N_13521,N_13678);
xnor U13938 (N_13938,N_13548,N_13580);
nand U13939 (N_13939,N_12941,N_13082);
and U13940 (N_13940,N_13506,N_12694);
xor U13941 (N_13941,N_12571,N_12559);
or U13942 (N_13942,N_13371,N_13694);
nor U13943 (N_13943,N_12895,N_13254);
and U13944 (N_13944,N_13707,N_13609);
nand U13945 (N_13945,N_13227,N_12976);
nand U13946 (N_13946,N_13596,N_13571);
xor U13947 (N_13947,N_13479,N_13025);
nand U13948 (N_13948,N_13241,N_13001);
or U13949 (N_13949,N_12648,N_13181);
nand U13950 (N_13950,N_12758,N_13187);
and U13951 (N_13951,N_12849,N_13132);
nor U13952 (N_13952,N_12956,N_13000);
nor U13953 (N_13953,N_13443,N_13628);
or U13954 (N_13954,N_13247,N_13608);
or U13955 (N_13955,N_12859,N_13704);
and U13956 (N_13956,N_12519,N_13370);
xor U13957 (N_13957,N_12765,N_13401);
or U13958 (N_13958,N_12785,N_13626);
nand U13959 (N_13959,N_13215,N_13397);
xor U13960 (N_13960,N_13593,N_12506);
nor U13961 (N_13961,N_13540,N_13528);
xor U13962 (N_13962,N_13446,N_13710);
xor U13963 (N_13963,N_13464,N_13298);
and U13964 (N_13964,N_12829,N_13014);
and U13965 (N_13965,N_13222,N_12889);
or U13966 (N_13966,N_13570,N_13683);
nor U13967 (N_13967,N_13243,N_13312);
nor U13968 (N_13968,N_13350,N_13191);
nand U13969 (N_13969,N_12633,N_13677);
xor U13970 (N_13970,N_12695,N_13360);
xnor U13971 (N_13971,N_13039,N_13515);
or U13972 (N_13972,N_13302,N_12721);
nor U13973 (N_13973,N_12973,N_12853);
and U13974 (N_13974,N_13100,N_12776);
xor U13975 (N_13975,N_13572,N_13412);
nand U13976 (N_13976,N_13052,N_12635);
and U13977 (N_13977,N_13315,N_12933);
xor U13978 (N_13978,N_13128,N_13592);
nor U13979 (N_13979,N_12663,N_12961);
or U13980 (N_13980,N_12661,N_12576);
or U13981 (N_13981,N_13368,N_13488);
nor U13982 (N_13982,N_13139,N_12986);
and U13983 (N_13983,N_13017,N_13495);
nand U13984 (N_13984,N_13680,N_12575);
and U13985 (N_13985,N_12647,N_12801);
xnor U13986 (N_13986,N_13026,N_13081);
or U13987 (N_13987,N_13041,N_13043);
and U13988 (N_13988,N_12591,N_12577);
and U13989 (N_13989,N_13286,N_13516);
nor U13990 (N_13990,N_12557,N_12930);
nand U13991 (N_13991,N_12821,N_13300);
or U13992 (N_13992,N_13044,N_12516);
xor U13993 (N_13993,N_12786,N_12845);
or U13994 (N_13994,N_12900,N_13116);
nor U13995 (N_13995,N_12805,N_13236);
nor U13996 (N_13996,N_13557,N_12777);
xor U13997 (N_13997,N_12502,N_12951);
and U13998 (N_13998,N_13523,N_13138);
nor U13999 (N_13999,N_12954,N_13705);
or U14000 (N_14000,N_13652,N_12875);
or U14001 (N_14001,N_13635,N_13006);
or U14002 (N_14002,N_13287,N_13649);
and U14003 (N_14003,N_13134,N_12728);
nand U14004 (N_14004,N_13567,N_13681);
xnor U14005 (N_14005,N_13429,N_13691);
or U14006 (N_14006,N_13153,N_13229);
or U14007 (N_14007,N_13478,N_12809);
xor U14008 (N_14008,N_12700,N_13522);
nand U14009 (N_14009,N_12683,N_13432);
and U14010 (N_14010,N_13098,N_12504);
nor U14011 (N_14011,N_12687,N_12901);
nand U14012 (N_14012,N_12794,N_13391);
xnor U14013 (N_14013,N_13170,N_13115);
or U14014 (N_14014,N_12795,N_13462);
xnor U14015 (N_14015,N_12971,N_13365);
nor U14016 (N_14016,N_12978,N_12688);
nand U14017 (N_14017,N_13729,N_13458);
nor U14018 (N_14018,N_13470,N_12997);
or U14019 (N_14019,N_13345,N_13366);
nor U14020 (N_14020,N_13669,N_12550);
and U14021 (N_14021,N_13529,N_12998);
nand U14022 (N_14022,N_13091,N_12739);
xnor U14023 (N_14023,N_13127,N_13015);
or U14024 (N_14024,N_13613,N_12972);
nor U14025 (N_14025,N_13010,N_13621);
nand U14026 (N_14026,N_12985,N_13225);
and U14027 (N_14027,N_13406,N_12907);
and U14028 (N_14028,N_13611,N_13018);
xor U14029 (N_14029,N_12967,N_12982);
xor U14030 (N_14030,N_13431,N_13193);
nor U14031 (N_14031,N_13320,N_12578);
nand U14032 (N_14032,N_13276,N_13113);
or U14033 (N_14033,N_13258,N_13740);
nand U14034 (N_14034,N_13237,N_12634);
or U14035 (N_14035,N_13643,N_13533);
or U14036 (N_14036,N_13053,N_13040);
or U14037 (N_14037,N_13264,N_13639);
and U14038 (N_14038,N_13096,N_12699);
xnor U14039 (N_14039,N_12888,N_12993);
and U14040 (N_14040,N_13746,N_13207);
nor U14041 (N_14041,N_12947,N_12551);
and U14042 (N_14042,N_13089,N_13405);
nor U14043 (N_14043,N_13008,N_12818);
and U14044 (N_14044,N_12935,N_12816);
nand U14045 (N_14045,N_13623,N_13509);
and U14046 (N_14046,N_12667,N_13463);
nor U14047 (N_14047,N_12703,N_12594);
and U14048 (N_14048,N_12673,N_13148);
xnor U14049 (N_14049,N_12949,N_13294);
or U14050 (N_14050,N_13124,N_13409);
xor U14051 (N_14051,N_12970,N_13741);
nor U14052 (N_14052,N_12929,N_12802);
or U14053 (N_14053,N_12723,N_13654);
or U14054 (N_14054,N_12911,N_13144);
xnor U14055 (N_14055,N_13256,N_13706);
and U14056 (N_14056,N_13354,N_13693);
nand U14057 (N_14057,N_12882,N_12644);
or U14058 (N_14058,N_12570,N_12531);
nor U14059 (N_14059,N_13467,N_13289);
nor U14060 (N_14060,N_13606,N_13541);
nand U14061 (N_14061,N_12981,N_13424);
nor U14062 (N_14062,N_12862,N_13192);
and U14063 (N_14063,N_12712,N_13631);
xnor U14064 (N_14064,N_13083,N_13619);
or U14065 (N_14065,N_13332,N_13067);
nand U14066 (N_14066,N_13292,N_13547);
nand U14067 (N_14067,N_13717,N_13377);
nor U14068 (N_14068,N_12581,N_13149);
or U14069 (N_14069,N_13378,N_13342);
and U14070 (N_14070,N_12534,N_12988);
and U14071 (N_14071,N_13582,N_12953);
and U14072 (N_14072,N_13435,N_13615);
nor U14073 (N_14073,N_13283,N_12727);
nor U14074 (N_14074,N_13585,N_12950);
xnor U14075 (N_14075,N_12822,N_12815);
nand U14076 (N_14076,N_13455,N_12783);
xor U14077 (N_14077,N_13388,N_12880);
and U14078 (N_14078,N_12606,N_13514);
nand U14079 (N_14079,N_12710,N_13456);
nor U14080 (N_14080,N_12992,N_13259);
nor U14081 (N_14081,N_13583,N_12893);
nor U14082 (N_14082,N_12587,N_13157);
and U14083 (N_14083,N_12847,N_13199);
nor U14084 (N_14084,N_13295,N_13238);
or U14085 (N_14085,N_12881,N_13071);
xor U14086 (N_14086,N_12991,N_12686);
nor U14087 (N_14087,N_13344,N_13195);
and U14088 (N_14088,N_12678,N_12593);
or U14089 (N_14089,N_12600,N_12774);
nor U14090 (N_14090,N_12624,N_13698);
or U14091 (N_14091,N_12705,N_13438);
or U14092 (N_14092,N_12766,N_12753);
and U14093 (N_14093,N_12749,N_13539);
xnor U14094 (N_14094,N_12514,N_12836);
nor U14095 (N_14095,N_13209,N_13189);
xor U14096 (N_14096,N_12904,N_13648);
and U14097 (N_14097,N_12620,N_13420);
nor U14098 (N_14098,N_13387,N_13527);
or U14099 (N_14099,N_12921,N_12556);
xnor U14100 (N_14100,N_13566,N_13065);
nor U14101 (N_14101,N_13550,N_12717);
and U14102 (N_14102,N_12989,N_12807);
or U14103 (N_14103,N_12597,N_13584);
nand U14104 (N_14104,N_12917,N_12511);
xor U14105 (N_14105,N_13517,N_13733);
or U14106 (N_14106,N_13564,N_13058);
nand U14107 (N_14107,N_13702,N_12547);
and U14108 (N_14108,N_13636,N_13673);
or U14109 (N_14109,N_13647,N_13073);
or U14110 (N_14110,N_13715,N_13313);
and U14111 (N_14111,N_13218,N_13348);
and U14112 (N_14112,N_13658,N_13735);
nor U14113 (N_14113,N_13747,N_13503);
or U14114 (N_14114,N_12817,N_13449);
nand U14115 (N_14115,N_12994,N_12931);
and U14116 (N_14116,N_13451,N_13558);
or U14117 (N_14117,N_12808,N_13646);
or U14118 (N_14118,N_13664,N_13047);
or U14119 (N_14119,N_12626,N_13070);
or U14120 (N_14120,N_12746,N_13208);
xor U14121 (N_14121,N_13549,N_13504);
nand U14122 (N_14122,N_12637,N_12509);
and U14123 (N_14123,N_13473,N_12905);
xor U14124 (N_14124,N_13355,N_13102);
nor U14125 (N_14125,N_12632,N_13211);
and U14126 (N_14126,N_12761,N_12825);
and U14127 (N_14127,N_13308,N_13033);
xnor U14128 (N_14128,N_13171,N_12868);
or U14129 (N_14129,N_13477,N_13016);
xnor U14130 (N_14130,N_13604,N_12763);
nand U14131 (N_14131,N_13486,N_13475);
nor U14132 (N_14132,N_12564,N_12923);
nor U14133 (N_14133,N_13212,N_13687);
nand U14134 (N_14134,N_13651,N_13398);
and U14135 (N_14135,N_13007,N_13367);
nand U14136 (N_14136,N_13358,N_13251);
and U14137 (N_14137,N_13725,N_13112);
and U14138 (N_14138,N_13339,N_13337);
nor U14139 (N_14139,N_13641,N_13736);
nor U14140 (N_14140,N_13296,N_12500);
or U14141 (N_14141,N_13607,N_12588);
or U14142 (N_14142,N_13353,N_12855);
or U14143 (N_14143,N_13700,N_13142);
xnor U14144 (N_14144,N_13494,N_12957);
nand U14145 (N_14145,N_12874,N_12697);
nor U14146 (N_14146,N_13380,N_13719);
or U14147 (N_14147,N_13575,N_12963);
or U14148 (N_14148,N_12867,N_13396);
xnor U14149 (N_14149,N_13246,N_12918);
and U14150 (N_14150,N_13361,N_13601);
xor U14151 (N_14151,N_13184,N_12879);
nor U14152 (N_14152,N_13546,N_13105);
xnor U14153 (N_14153,N_13491,N_12621);
and U14154 (N_14154,N_12730,N_13389);
xnor U14155 (N_14155,N_13385,N_13659);
and U14156 (N_14156,N_12942,N_12958);
or U14157 (N_14157,N_13011,N_13140);
nor U14158 (N_14158,N_12562,N_12995);
or U14159 (N_14159,N_13665,N_13513);
nor U14160 (N_14160,N_12769,N_13423);
nor U14161 (N_14161,N_12702,N_13305);
xor U14162 (N_14162,N_12831,N_12797);
or U14163 (N_14163,N_13062,N_13728);
nor U14164 (N_14164,N_13194,N_13183);
or U14165 (N_14165,N_13703,N_12851);
and U14166 (N_14166,N_13217,N_12828);
and U14167 (N_14167,N_13440,N_13510);
and U14168 (N_14168,N_13562,N_13489);
and U14169 (N_14169,N_13716,N_12657);
xor U14170 (N_14170,N_13525,N_12558);
and U14171 (N_14171,N_12654,N_12890);
and U14172 (N_14172,N_13330,N_13210);
nand U14173 (N_14173,N_12515,N_12857);
nor U14174 (N_14174,N_12894,N_13690);
nor U14175 (N_14175,N_13204,N_12778);
xnor U14176 (N_14176,N_13030,N_13303);
xor U14177 (N_14177,N_13375,N_12732);
nor U14178 (N_14178,N_13586,N_12798);
nand U14179 (N_14179,N_13663,N_12887);
nand U14180 (N_14180,N_12810,N_13338);
or U14181 (N_14181,N_12666,N_13472);
nand U14182 (N_14182,N_12722,N_12946);
nor U14183 (N_14183,N_12936,N_13319);
xnor U14184 (N_14184,N_13162,N_12792);
or U14185 (N_14185,N_13009,N_12920);
nor U14186 (N_14186,N_13642,N_12583);
and U14187 (N_14187,N_12522,N_13587);
xnor U14188 (N_14188,N_13341,N_12799);
nor U14189 (N_14189,N_13111,N_12716);
or U14190 (N_14190,N_12709,N_12823);
or U14191 (N_14191,N_13156,N_13552);
nor U14192 (N_14192,N_12629,N_12908);
or U14193 (N_14193,N_13235,N_13335);
xor U14194 (N_14194,N_13087,N_13561);
and U14195 (N_14195,N_13290,N_13284);
and U14196 (N_14196,N_12980,N_13682);
xor U14197 (N_14197,N_13721,N_12553);
nand U14198 (N_14198,N_13137,N_13656);
and U14199 (N_14199,N_13545,N_13428);
nor U14200 (N_14200,N_13231,N_13200);
nand U14201 (N_14201,N_13629,N_13049);
nand U14202 (N_14202,N_12800,N_13224);
or U14203 (N_14203,N_13356,N_12604);
nor U14204 (N_14204,N_12793,N_13230);
nor U14205 (N_14205,N_13696,N_13042);
nor U14206 (N_14206,N_12734,N_13012);
or U14207 (N_14207,N_13708,N_13542);
xor U14208 (N_14208,N_13108,N_13471);
or U14209 (N_14209,N_13056,N_12772);
and U14210 (N_14210,N_13036,N_13638);
nor U14211 (N_14211,N_13695,N_13169);
nand U14212 (N_14212,N_13064,N_13051);
xnor U14213 (N_14213,N_13027,N_12668);
xor U14214 (N_14214,N_13163,N_13066);
and U14215 (N_14215,N_13093,N_13403);
nand U14216 (N_14216,N_13461,N_13329);
nor U14217 (N_14217,N_13560,N_13743);
xnor U14218 (N_14218,N_13352,N_12528);
and U14219 (N_14219,N_13090,N_13321);
nor U14220 (N_14220,N_13133,N_12569);
and U14221 (N_14221,N_13576,N_13569);
and U14222 (N_14222,N_12701,N_13035);
xnor U14223 (N_14223,N_13732,N_13023);
nor U14224 (N_14224,N_13245,N_12843);
nor U14225 (N_14225,N_12854,N_13114);
and U14226 (N_14226,N_12540,N_12512);
or U14227 (N_14227,N_13328,N_12848);
and U14228 (N_14228,N_12885,N_12628);
and U14229 (N_14229,N_12725,N_13322);
or U14230 (N_14230,N_13206,N_13220);
or U14231 (N_14231,N_13662,N_13402);
and U14232 (N_14232,N_12939,N_12870);
nor U14233 (N_14233,N_13279,N_13553);
nand U14234 (N_14234,N_13242,N_13034);
or U14235 (N_14235,N_12707,N_13357);
nor U14236 (N_14236,N_13524,N_13487);
nor U14237 (N_14237,N_13381,N_13021);
and U14238 (N_14238,N_12554,N_12636);
and U14239 (N_14239,N_13551,N_13640);
xor U14240 (N_14240,N_13159,N_12532);
nand U14241 (N_14241,N_12596,N_13590);
nand U14242 (N_14242,N_13413,N_13476);
nand U14243 (N_14243,N_12517,N_12530);
nor U14244 (N_14244,N_12838,N_13614);
or U14245 (N_14245,N_13013,N_12745);
or U14246 (N_14246,N_13055,N_13226);
or U14247 (N_14247,N_13731,N_13622);
xor U14248 (N_14248,N_12653,N_12631);
xor U14249 (N_14249,N_13544,N_13734);
nor U14250 (N_14250,N_12698,N_13502);
xnor U14251 (N_14251,N_12613,N_13084);
or U14252 (N_14252,N_13197,N_12513);
and U14253 (N_14253,N_13426,N_13395);
xnor U14254 (N_14254,N_12590,N_12773);
nand U14255 (N_14255,N_13407,N_12671);
nor U14256 (N_14256,N_12708,N_13129);
xnor U14257 (N_14257,N_13118,N_12689);
nand U14258 (N_14258,N_13002,N_12542);
xor U14259 (N_14259,N_12665,N_12830);
or U14260 (N_14260,N_13417,N_13482);
nand U14261 (N_14261,N_12523,N_13003);
nand U14262 (N_14262,N_12820,N_12603);
xnor U14263 (N_14263,N_13152,N_13433);
nor U14264 (N_14264,N_12891,N_13618);
or U14265 (N_14265,N_12555,N_12884);
and U14266 (N_14266,N_12706,N_13078);
nor U14267 (N_14267,N_12760,N_12731);
nor U14268 (N_14268,N_13620,N_13685);
or U14269 (N_14269,N_13050,N_13031);
xnor U14270 (N_14270,N_12811,N_13179);
and U14271 (N_14271,N_12906,N_13439);
nor U14272 (N_14272,N_13109,N_12584);
and U14273 (N_14273,N_13101,N_13701);
nor U14274 (N_14274,N_13165,N_13666);
or U14275 (N_14275,N_12876,N_13692);
or U14276 (N_14276,N_12696,N_12715);
nor U14277 (N_14277,N_13146,N_13573);
or U14278 (N_14278,N_12595,N_12789);
or U14279 (N_14279,N_13382,N_13722);
or U14280 (N_14280,N_13343,N_13713);
or U14281 (N_14281,N_12919,N_13219);
xor U14282 (N_14282,N_12741,N_12928);
or U14283 (N_14283,N_12693,N_12567);
nor U14284 (N_14284,N_12649,N_13595);
and U14285 (N_14285,N_12872,N_12622);
and U14286 (N_14286,N_12877,N_13147);
xnor U14287 (N_14287,N_12768,N_12614);
nor U14288 (N_14288,N_12602,N_13301);
and U14289 (N_14289,N_13632,N_12599);
nor U14290 (N_14290,N_13046,N_13660);
nand U14291 (N_14291,N_13253,N_12925);
and U14292 (N_14292,N_12507,N_13154);
nor U14293 (N_14293,N_13425,N_13500);
nand U14294 (N_14294,N_13324,N_13531);
or U14295 (N_14295,N_13240,N_13120);
or U14296 (N_14296,N_12501,N_13095);
or U14297 (N_14297,N_13060,N_13029);
or U14298 (N_14298,N_13444,N_12692);
xor U14299 (N_14299,N_13110,N_12726);
nor U14300 (N_14300,N_13346,N_13634);
nor U14301 (N_14301,N_13374,N_13610);
or U14302 (N_14302,N_12609,N_13161);
nor U14303 (N_14303,N_12582,N_12610);
nand U14304 (N_14304,N_13244,N_13538);
nor U14305 (N_14305,N_12662,N_13369);
or U14306 (N_14306,N_13262,N_12643);
nor U14307 (N_14307,N_13490,N_12835);
nor U14308 (N_14308,N_12658,N_12756);
nor U14309 (N_14309,N_13347,N_13644);
xnor U14310 (N_14310,N_13468,N_13314);
or U14311 (N_14311,N_12983,N_13185);
nor U14312 (N_14312,N_13744,N_13123);
nor U14313 (N_14313,N_13454,N_12782);
xnor U14314 (N_14314,N_13578,N_12704);
and U14315 (N_14315,N_12585,N_13107);
or U14316 (N_14316,N_12714,N_13667);
and U14317 (N_14317,N_12656,N_13309);
and U14318 (N_14318,N_13299,N_13094);
and U14319 (N_14319,N_12720,N_13498);
nand U14320 (N_14320,N_13119,N_12690);
and U14321 (N_14321,N_12645,N_12729);
nor U14322 (N_14322,N_13022,N_12640);
nor U14323 (N_14323,N_12618,N_12948);
and U14324 (N_14324,N_13214,N_13650);
nor U14325 (N_14325,N_12543,N_13430);
or U14326 (N_14326,N_12691,N_12850);
nand U14327 (N_14327,N_13624,N_13714);
nand U14328 (N_14328,N_13151,N_13180);
or U14329 (N_14329,N_13399,N_13452);
xnor U14330 (N_14330,N_13061,N_13351);
nor U14331 (N_14331,N_13709,N_12819);
nor U14332 (N_14332,N_13727,N_13605);
or U14333 (N_14333,N_13075,N_13282);
and U14334 (N_14334,N_12924,N_12552);
nor U14335 (N_14335,N_12791,N_12770);
xor U14336 (N_14336,N_13143,N_13233);
xor U14337 (N_14337,N_13131,N_12742);
nor U14338 (N_14338,N_12619,N_12611);
nor U14339 (N_14339,N_12892,N_13005);
xor U14340 (N_14340,N_13661,N_13441);
or U14341 (N_14341,N_13136,N_13520);
and U14342 (N_14342,N_13492,N_13270);
xnor U14343 (N_14343,N_12546,N_13493);
nor U14344 (N_14344,N_12899,N_13591);
nor U14345 (N_14345,N_13679,N_12650);
xnor U14346 (N_14346,N_13274,N_12505);
xnor U14347 (N_14347,N_12510,N_13054);
nor U14348 (N_14348,N_13249,N_13285);
xnor U14349 (N_14349,N_12639,N_13048);
nand U14350 (N_14350,N_12841,N_13130);
nand U14351 (N_14351,N_12833,N_13166);
nand U14352 (N_14352,N_12533,N_12757);
nand U14353 (N_14353,N_12713,N_13239);
and U14354 (N_14354,N_13252,N_13419);
and U14355 (N_14355,N_12966,N_13686);
and U14356 (N_14356,N_12759,N_12566);
xor U14357 (N_14357,N_13483,N_13020);
xnor U14358 (N_14358,N_13379,N_13141);
xnor U14359 (N_14359,N_12548,N_13293);
or U14360 (N_14360,N_12539,N_13384);
or U14361 (N_14361,N_12549,N_12659);
xnor U14362 (N_14362,N_12521,N_13497);
nand U14363 (N_14363,N_13359,N_13688);
or U14364 (N_14364,N_12965,N_12615);
or U14365 (N_14365,N_12711,N_12955);
nand U14366 (N_14366,N_13689,N_13158);
and U14367 (N_14367,N_13336,N_12652);
and U14368 (N_14368,N_13117,N_12927);
or U14369 (N_14369,N_12669,N_12664);
and U14370 (N_14370,N_13534,N_13505);
xor U14371 (N_14371,N_12977,N_13363);
and U14372 (N_14372,N_13318,N_12812);
nand U14373 (N_14373,N_13745,N_13738);
or U14374 (N_14374,N_12586,N_13024);
xnor U14375 (N_14375,N_13296,N_13374);
or U14376 (N_14376,N_13110,N_13618);
or U14377 (N_14377,N_13351,N_12955);
or U14378 (N_14378,N_13249,N_12990);
and U14379 (N_14379,N_13006,N_13163);
nand U14380 (N_14380,N_12622,N_12992);
nand U14381 (N_14381,N_12823,N_12572);
and U14382 (N_14382,N_13585,N_13471);
and U14383 (N_14383,N_13368,N_13167);
or U14384 (N_14384,N_13036,N_12651);
or U14385 (N_14385,N_12884,N_12630);
nor U14386 (N_14386,N_12996,N_13079);
nand U14387 (N_14387,N_12919,N_13346);
nor U14388 (N_14388,N_12539,N_13168);
and U14389 (N_14389,N_12834,N_12901);
and U14390 (N_14390,N_12558,N_13712);
nand U14391 (N_14391,N_12725,N_13471);
and U14392 (N_14392,N_12824,N_12516);
xor U14393 (N_14393,N_13201,N_13546);
xnor U14394 (N_14394,N_13105,N_13351);
or U14395 (N_14395,N_13730,N_13030);
xor U14396 (N_14396,N_13548,N_13570);
nand U14397 (N_14397,N_12834,N_13423);
nand U14398 (N_14398,N_13068,N_13392);
xnor U14399 (N_14399,N_13405,N_12710);
or U14400 (N_14400,N_13600,N_13040);
or U14401 (N_14401,N_12773,N_13141);
and U14402 (N_14402,N_13275,N_13050);
nand U14403 (N_14403,N_13441,N_12558);
nor U14404 (N_14404,N_13071,N_13486);
xnor U14405 (N_14405,N_13407,N_12765);
nand U14406 (N_14406,N_12892,N_13533);
nand U14407 (N_14407,N_12765,N_12867);
and U14408 (N_14408,N_12859,N_12828);
nor U14409 (N_14409,N_13335,N_13377);
and U14410 (N_14410,N_13383,N_12538);
xor U14411 (N_14411,N_12660,N_13204);
and U14412 (N_14412,N_13522,N_13293);
and U14413 (N_14413,N_13228,N_13255);
xor U14414 (N_14414,N_13276,N_13528);
xnor U14415 (N_14415,N_13236,N_12860);
nor U14416 (N_14416,N_13635,N_13626);
nand U14417 (N_14417,N_12893,N_13236);
xnor U14418 (N_14418,N_13068,N_12732);
or U14419 (N_14419,N_13090,N_12854);
xor U14420 (N_14420,N_12971,N_12750);
or U14421 (N_14421,N_13669,N_12885);
nand U14422 (N_14422,N_13367,N_12785);
or U14423 (N_14423,N_12618,N_12752);
nor U14424 (N_14424,N_13015,N_12524);
nor U14425 (N_14425,N_13294,N_12688);
and U14426 (N_14426,N_12845,N_13616);
nand U14427 (N_14427,N_13154,N_13641);
xor U14428 (N_14428,N_13577,N_13134);
nand U14429 (N_14429,N_13375,N_12767);
and U14430 (N_14430,N_12830,N_13746);
and U14431 (N_14431,N_13358,N_13467);
and U14432 (N_14432,N_12923,N_13190);
nand U14433 (N_14433,N_13736,N_13538);
and U14434 (N_14434,N_13179,N_13567);
or U14435 (N_14435,N_12838,N_12925);
or U14436 (N_14436,N_13166,N_13448);
nand U14437 (N_14437,N_13023,N_12709);
and U14438 (N_14438,N_13449,N_12659);
nand U14439 (N_14439,N_12887,N_13232);
and U14440 (N_14440,N_13457,N_13682);
nor U14441 (N_14441,N_13205,N_12700);
and U14442 (N_14442,N_13179,N_13085);
nor U14443 (N_14443,N_13179,N_12547);
xnor U14444 (N_14444,N_13538,N_12549);
xor U14445 (N_14445,N_13510,N_13449);
nand U14446 (N_14446,N_13140,N_13644);
nor U14447 (N_14447,N_13193,N_12577);
and U14448 (N_14448,N_13474,N_12777);
or U14449 (N_14449,N_12611,N_12833);
and U14450 (N_14450,N_12650,N_13731);
and U14451 (N_14451,N_13432,N_13707);
and U14452 (N_14452,N_12813,N_13214);
xor U14453 (N_14453,N_12873,N_12827);
nor U14454 (N_14454,N_13574,N_12624);
nor U14455 (N_14455,N_13655,N_12868);
xor U14456 (N_14456,N_13643,N_13311);
nand U14457 (N_14457,N_12511,N_13398);
nand U14458 (N_14458,N_12553,N_12700);
and U14459 (N_14459,N_12798,N_13005);
nor U14460 (N_14460,N_13405,N_12529);
nand U14461 (N_14461,N_13051,N_13617);
nand U14462 (N_14462,N_12961,N_13015);
and U14463 (N_14463,N_13498,N_13165);
and U14464 (N_14464,N_12903,N_13072);
nor U14465 (N_14465,N_13448,N_13343);
nor U14466 (N_14466,N_12893,N_13379);
nor U14467 (N_14467,N_12732,N_13427);
xnor U14468 (N_14468,N_12672,N_12828);
nor U14469 (N_14469,N_12722,N_13339);
nand U14470 (N_14470,N_13076,N_12518);
or U14471 (N_14471,N_13443,N_13171);
nand U14472 (N_14472,N_12898,N_13359);
nor U14473 (N_14473,N_12723,N_13154);
nand U14474 (N_14474,N_13029,N_13686);
and U14475 (N_14475,N_13234,N_12641);
or U14476 (N_14476,N_13190,N_12674);
nor U14477 (N_14477,N_13730,N_12835);
nand U14478 (N_14478,N_12963,N_13188);
xor U14479 (N_14479,N_12562,N_13192);
xor U14480 (N_14480,N_12922,N_13587);
xnor U14481 (N_14481,N_13485,N_12819);
nor U14482 (N_14482,N_13360,N_13594);
nand U14483 (N_14483,N_12537,N_12617);
or U14484 (N_14484,N_13426,N_12756);
xor U14485 (N_14485,N_13687,N_13718);
xnor U14486 (N_14486,N_13309,N_12556);
and U14487 (N_14487,N_12641,N_13509);
nand U14488 (N_14488,N_13124,N_13054);
xor U14489 (N_14489,N_12722,N_13473);
nor U14490 (N_14490,N_12659,N_12526);
or U14491 (N_14491,N_13336,N_12630);
or U14492 (N_14492,N_12947,N_13253);
xnor U14493 (N_14493,N_12770,N_13059);
or U14494 (N_14494,N_13692,N_13353);
or U14495 (N_14495,N_13062,N_13060);
nand U14496 (N_14496,N_12774,N_13291);
or U14497 (N_14497,N_12681,N_13349);
or U14498 (N_14498,N_12694,N_13079);
and U14499 (N_14499,N_13542,N_13570);
xnor U14500 (N_14500,N_13391,N_13118);
nor U14501 (N_14501,N_13692,N_13446);
or U14502 (N_14502,N_13721,N_13138);
xnor U14503 (N_14503,N_13342,N_12727);
nor U14504 (N_14504,N_12879,N_12655);
and U14505 (N_14505,N_13064,N_13459);
nor U14506 (N_14506,N_13223,N_13672);
nor U14507 (N_14507,N_13570,N_13529);
nor U14508 (N_14508,N_12867,N_12883);
nor U14509 (N_14509,N_12871,N_13082);
xnor U14510 (N_14510,N_13468,N_12655);
or U14511 (N_14511,N_13657,N_12597);
nand U14512 (N_14512,N_12820,N_12673);
xor U14513 (N_14513,N_12982,N_13248);
nand U14514 (N_14514,N_12583,N_12848);
nor U14515 (N_14515,N_12817,N_12738);
xor U14516 (N_14516,N_13089,N_13302);
nor U14517 (N_14517,N_13585,N_13172);
nor U14518 (N_14518,N_13641,N_12639);
and U14519 (N_14519,N_13449,N_12666);
and U14520 (N_14520,N_12842,N_12977);
xnor U14521 (N_14521,N_12728,N_13274);
xnor U14522 (N_14522,N_13188,N_12810);
nand U14523 (N_14523,N_13070,N_13324);
nor U14524 (N_14524,N_12672,N_12510);
nand U14525 (N_14525,N_12554,N_13127);
nand U14526 (N_14526,N_13462,N_12888);
nand U14527 (N_14527,N_13379,N_12657);
nand U14528 (N_14528,N_12946,N_13051);
xor U14529 (N_14529,N_13361,N_13426);
or U14530 (N_14530,N_13091,N_13472);
and U14531 (N_14531,N_13433,N_13096);
nor U14532 (N_14532,N_13295,N_13378);
and U14533 (N_14533,N_13626,N_13262);
xor U14534 (N_14534,N_13350,N_13666);
nor U14535 (N_14535,N_12524,N_12756);
and U14536 (N_14536,N_13303,N_13087);
xnor U14537 (N_14537,N_13592,N_13239);
and U14538 (N_14538,N_13222,N_13173);
nor U14539 (N_14539,N_13125,N_13425);
or U14540 (N_14540,N_13185,N_13146);
nor U14541 (N_14541,N_12559,N_13357);
xnor U14542 (N_14542,N_12627,N_12662);
nand U14543 (N_14543,N_12952,N_13088);
nor U14544 (N_14544,N_13487,N_13106);
or U14545 (N_14545,N_12812,N_13425);
nor U14546 (N_14546,N_12519,N_13040);
and U14547 (N_14547,N_12796,N_12918);
and U14548 (N_14548,N_12801,N_13434);
xor U14549 (N_14549,N_12862,N_13131);
or U14550 (N_14550,N_13135,N_12911);
and U14551 (N_14551,N_13672,N_12591);
nor U14552 (N_14552,N_12977,N_12820);
or U14553 (N_14553,N_13667,N_12992);
xnor U14554 (N_14554,N_13661,N_12861);
and U14555 (N_14555,N_13311,N_12502);
or U14556 (N_14556,N_13168,N_12582);
nor U14557 (N_14557,N_13710,N_13070);
xor U14558 (N_14558,N_12871,N_13596);
and U14559 (N_14559,N_12881,N_13748);
nand U14560 (N_14560,N_13004,N_13713);
and U14561 (N_14561,N_13504,N_13192);
nor U14562 (N_14562,N_13544,N_13376);
nor U14563 (N_14563,N_13724,N_13091);
and U14564 (N_14564,N_13503,N_13390);
and U14565 (N_14565,N_13347,N_12944);
nand U14566 (N_14566,N_12694,N_13686);
nand U14567 (N_14567,N_13586,N_13120);
xor U14568 (N_14568,N_13219,N_13416);
xnor U14569 (N_14569,N_12536,N_12830);
nand U14570 (N_14570,N_13064,N_12965);
nor U14571 (N_14571,N_12956,N_12729);
nor U14572 (N_14572,N_13499,N_13364);
nand U14573 (N_14573,N_12855,N_12723);
nand U14574 (N_14574,N_13236,N_13417);
or U14575 (N_14575,N_12684,N_13008);
and U14576 (N_14576,N_13263,N_13280);
nor U14577 (N_14577,N_13383,N_13284);
xor U14578 (N_14578,N_12512,N_13663);
or U14579 (N_14579,N_12789,N_12863);
nor U14580 (N_14580,N_13578,N_13187);
xor U14581 (N_14581,N_12687,N_13197);
nand U14582 (N_14582,N_12879,N_12799);
or U14583 (N_14583,N_13526,N_12583);
xnor U14584 (N_14584,N_12946,N_13133);
nand U14585 (N_14585,N_12883,N_13389);
nand U14586 (N_14586,N_12570,N_13462);
or U14587 (N_14587,N_12934,N_13154);
nand U14588 (N_14588,N_13108,N_13033);
and U14589 (N_14589,N_13190,N_13686);
and U14590 (N_14590,N_13631,N_13545);
and U14591 (N_14591,N_13584,N_13025);
nor U14592 (N_14592,N_13369,N_12563);
nand U14593 (N_14593,N_12806,N_13464);
nand U14594 (N_14594,N_12901,N_13142);
nor U14595 (N_14595,N_12679,N_13131);
and U14596 (N_14596,N_13300,N_12525);
xor U14597 (N_14597,N_12563,N_12995);
nand U14598 (N_14598,N_13101,N_13613);
nand U14599 (N_14599,N_13540,N_12792);
nand U14600 (N_14600,N_12876,N_12867);
and U14601 (N_14601,N_13381,N_13611);
nand U14602 (N_14602,N_13080,N_13097);
or U14603 (N_14603,N_12603,N_12691);
nor U14604 (N_14604,N_13025,N_13586);
or U14605 (N_14605,N_13566,N_13205);
xnor U14606 (N_14606,N_12751,N_12875);
nor U14607 (N_14607,N_13158,N_13429);
xnor U14608 (N_14608,N_13224,N_13562);
or U14609 (N_14609,N_13701,N_13605);
xor U14610 (N_14610,N_13203,N_12818);
xor U14611 (N_14611,N_13207,N_13340);
and U14612 (N_14612,N_12518,N_13135);
nand U14613 (N_14613,N_13658,N_12676);
and U14614 (N_14614,N_13154,N_13376);
and U14615 (N_14615,N_13009,N_13062);
nand U14616 (N_14616,N_12533,N_12651);
nor U14617 (N_14617,N_12970,N_13557);
or U14618 (N_14618,N_12666,N_13723);
xnor U14619 (N_14619,N_12944,N_13016);
nand U14620 (N_14620,N_13216,N_12710);
and U14621 (N_14621,N_13187,N_12552);
and U14622 (N_14622,N_12599,N_13253);
and U14623 (N_14623,N_13340,N_13076);
and U14624 (N_14624,N_13370,N_12864);
nor U14625 (N_14625,N_13186,N_12694);
and U14626 (N_14626,N_13252,N_12781);
nor U14627 (N_14627,N_13485,N_13415);
and U14628 (N_14628,N_12519,N_13497);
and U14629 (N_14629,N_13255,N_13613);
and U14630 (N_14630,N_12855,N_12654);
or U14631 (N_14631,N_13262,N_12708);
nand U14632 (N_14632,N_13694,N_12867);
or U14633 (N_14633,N_13632,N_12812);
nor U14634 (N_14634,N_12880,N_13499);
xnor U14635 (N_14635,N_12770,N_13561);
xor U14636 (N_14636,N_13387,N_13226);
and U14637 (N_14637,N_13588,N_13294);
or U14638 (N_14638,N_13495,N_13022);
and U14639 (N_14639,N_12954,N_13505);
and U14640 (N_14640,N_13177,N_12536);
or U14641 (N_14641,N_13744,N_13503);
nor U14642 (N_14642,N_13559,N_12653);
xor U14643 (N_14643,N_13071,N_12820);
or U14644 (N_14644,N_13631,N_12535);
and U14645 (N_14645,N_13730,N_13013);
xor U14646 (N_14646,N_12652,N_13375);
nand U14647 (N_14647,N_13522,N_12653);
and U14648 (N_14648,N_13265,N_12787);
nor U14649 (N_14649,N_13107,N_12973);
xnor U14650 (N_14650,N_13084,N_13601);
and U14651 (N_14651,N_12836,N_13021);
and U14652 (N_14652,N_13147,N_13491);
or U14653 (N_14653,N_13631,N_13358);
and U14654 (N_14654,N_13123,N_13682);
or U14655 (N_14655,N_12739,N_13431);
or U14656 (N_14656,N_13702,N_13196);
or U14657 (N_14657,N_12674,N_12584);
xnor U14658 (N_14658,N_12843,N_13663);
nor U14659 (N_14659,N_13282,N_12511);
nor U14660 (N_14660,N_13094,N_13535);
nor U14661 (N_14661,N_12736,N_13179);
or U14662 (N_14662,N_13601,N_13258);
nor U14663 (N_14663,N_13266,N_13560);
or U14664 (N_14664,N_12941,N_13488);
or U14665 (N_14665,N_13402,N_12891);
or U14666 (N_14666,N_12868,N_12684);
nor U14667 (N_14667,N_13457,N_12641);
or U14668 (N_14668,N_12861,N_12683);
nand U14669 (N_14669,N_12961,N_13195);
nand U14670 (N_14670,N_13262,N_13512);
nor U14671 (N_14671,N_12715,N_13571);
nor U14672 (N_14672,N_12953,N_13554);
nor U14673 (N_14673,N_13003,N_13579);
or U14674 (N_14674,N_12752,N_12985);
xnor U14675 (N_14675,N_13687,N_13171);
or U14676 (N_14676,N_13183,N_13149);
nor U14677 (N_14677,N_13731,N_13300);
and U14678 (N_14678,N_12556,N_13111);
xor U14679 (N_14679,N_12525,N_13627);
and U14680 (N_14680,N_12768,N_12751);
or U14681 (N_14681,N_13602,N_13613);
and U14682 (N_14682,N_12562,N_13410);
or U14683 (N_14683,N_12942,N_13290);
or U14684 (N_14684,N_12733,N_13233);
nand U14685 (N_14685,N_13534,N_13287);
or U14686 (N_14686,N_12515,N_12538);
and U14687 (N_14687,N_12868,N_12580);
nand U14688 (N_14688,N_12715,N_12694);
nor U14689 (N_14689,N_12952,N_13123);
and U14690 (N_14690,N_13507,N_12939);
nand U14691 (N_14691,N_13180,N_13647);
and U14692 (N_14692,N_12944,N_13327);
or U14693 (N_14693,N_12682,N_13601);
xnor U14694 (N_14694,N_13602,N_12519);
nand U14695 (N_14695,N_13488,N_12964);
xor U14696 (N_14696,N_13508,N_13395);
nand U14697 (N_14697,N_12500,N_12974);
nor U14698 (N_14698,N_13485,N_12754);
nand U14699 (N_14699,N_12980,N_13442);
nand U14700 (N_14700,N_13016,N_13687);
nor U14701 (N_14701,N_13663,N_12993);
and U14702 (N_14702,N_12514,N_13617);
or U14703 (N_14703,N_12984,N_12744);
and U14704 (N_14704,N_12744,N_12558);
or U14705 (N_14705,N_13462,N_13584);
nand U14706 (N_14706,N_12556,N_13340);
nor U14707 (N_14707,N_13424,N_13549);
nor U14708 (N_14708,N_12667,N_12622);
nor U14709 (N_14709,N_13459,N_13196);
and U14710 (N_14710,N_12853,N_13178);
nand U14711 (N_14711,N_13425,N_12791);
nand U14712 (N_14712,N_13002,N_13738);
xor U14713 (N_14713,N_13114,N_13508);
and U14714 (N_14714,N_13615,N_12933);
nor U14715 (N_14715,N_13578,N_13355);
and U14716 (N_14716,N_13051,N_12560);
xnor U14717 (N_14717,N_12799,N_13155);
and U14718 (N_14718,N_13438,N_13290);
and U14719 (N_14719,N_13641,N_12784);
nor U14720 (N_14720,N_12945,N_13243);
nand U14721 (N_14721,N_12992,N_13112);
nand U14722 (N_14722,N_13247,N_12993);
and U14723 (N_14723,N_12720,N_13524);
nand U14724 (N_14724,N_13625,N_12887);
nor U14725 (N_14725,N_13513,N_13486);
or U14726 (N_14726,N_13082,N_13459);
and U14727 (N_14727,N_12623,N_12834);
or U14728 (N_14728,N_13485,N_12916);
or U14729 (N_14729,N_12754,N_12749);
xor U14730 (N_14730,N_13084,N_13730);
xor U14731 (N_14731,N_13084,N_13612);
nand U14732 (N_14732,N_13170,N_13623);
or U14733 (N_14733,N_12995,N_12801);
or U14734 (N_14734,N_12940,N_12822);
and U14735 (N_14735,N_12895,N_13449);
nand U14736 (N_14736,N_13511,N_13108);
nor U14737 (N_14737,N_13216,N_12705);
xnor U14738 (N_14738,N_13434,N_13548);
and U14739 (N_14739,N_13015,N_13525);
or U14740 (N_14740,N_13175,N_13067);
and U14741 (N_14741,N_12821,N_12870);
xnor U14742 (N_14742,N_12862,N_13311);
nor U14743 (N_14743,N_13599,N_12646);
nand U14744 (N_14744,N_13605,N_13459);
and U14745 (N_14745,N_13581,N_13412);
nor U14746 (N_14746,N_13106,N_13352);
xor U14747 (N_14747,N_13059,N_13586);
xnor U14748 (N_14748,N_13180,N_12545);
and U14749 (N_14749,N_13114,N_12758);
or U14750 (N_14750,N_13505,N_12589);
nor U14751 (N_14751,N_12966,N_12969);
nor U14752 (N_14752,N_12541,N_12790);
or U14753 (N_14753,N_13615,N_13194);
and U14754 (N_14754,N_13529,N_12907);
xor U14755 (N_14755,N_13525,N_13424);
nand U14756 (N_14756,N_13551,N_12584);
or U14757 (N_14757,N_12565,N_12567);
or U14758 (N_14758,N_13558,N_12599);
nand U14759 (N_14759,N_12722,N_12546);
xnor U14760 (N_14760,N_12786,N_13127);
nor U14761 (N_14761,N_12669,N_13215);
nand U14762 (N_14762,N_13018,N_12826);
nand U14763 (N_14763,N_13327,N_12943);
nand U14764 (N_14764,N_13029,N_13718);
nor U14765 (N_14765,N_12733,N_12694);
xor U14766 (N_14766,N_13566,N_13263);
and U14767 (N_14767,N_12766,N_12882);
and U14768 (N_14768,N_12804,N_13391);
nor U14769 (N_14769,N_12932,N_13429);
or U14770 (N_14770,N_12933,N_13232);
or U14771 (N_14771,N_13140,N_12690);
or U14772 (N_14772,N_12989,N_12902);
nand U14773 (N_14773,N_13186,N_12986);
xnor U14774 (N_14774,N_12561,N_12815);
nand U14775 (N_14775,N_13351,N_12608);
or U14776 (N_14776,N_13511,N_12692);
nor U14777 (N_14777,N_13255,N_13618);
or U14778 (N_14778,N_13401,N_12838);
nand U14779 (N_14779,N_12587,N_12937);
nor U14780 (N_14780,N_13045,N_13068);
xnor U14781 (N_14781,N_12715,N_12597);
and U14782 (N_14782,N_12835,N_13139);
nand U14783 (N_14783,N_13486,N_12893);
xnor U14784 (N_14784,N_13261,N_13454);
xnor U14785 (N_14785,N_12566,N_13577);
and U14786 (N_14786,N_13014,N_13692);
or U14787 (N_14787,N_12814,N_12804);
and U14788 (N_14788,N_13283,N_12704);
or U14789 (N_14789,N_13414,N_12961);
xnor U14790 (N_14790,N_13122,N_13492);
xor U14791 (N_14791,N_13533,N_13096);
xnor U14792 (N_14792,N_13318,N_12593);
nand U14793 (N_14793,N_12922,N_13492);
nor U14794 (N_14794,N_12745,N_13173);
or U14795 (N_14795,N_12853,N_13468);
and U14796 (N_14796,N_13321,N_13449);
or U14797 (N_14797,N_13607,N_12538);
xor U14798 (N_14798,N_13105,N_12603);
and U14799 (N_14799,N_13118,N_13226);
xor U14800 (N_14800,N_12797,N_12983);
nand U14801 (N_14801,N_12956,N_13435);
and U14802 (N_14802,N_12699,N_12626);
nand U14803 (N_14803,N_12808,N_13260);
and U14804 (N_14804,N_13715,N_13563);
nand U14805 (N_14805,N_12977,N_13397);
or U14806 (N_14806,N_13392,N_13393);
nand U14807 (N_14807,N_13390,N_12509);
nand U14808 (N_14808,N_13035,N_13183);
xor U14809 (N_14809,N_13546,N_12656);
nand U14810 (N_14810,N_12903,N_12668);
and U14811 (N_14811,N_12810,N_13225);
nor U14812 (N_14812,N_12955,N_13337);
xnor U14813 (N_14813,N_13263,N_13498);
nor U14814 (N_14814,N_13545,N_12626);
nand U14815 (N_14815,N_13451,N_12505);
nor U14816 (N_14816,N_13214,N_12664);
or U14817 (N_14817,N_13327,N_12868);
or U14818 (N_14818,N_13578,N_12530);
nand U14819 (N_14819,N_13196,N_12646);
and U14820 (N_14820,N_13456,N_12859);
xnor U14821 (N_14821,N_13581,N_12574);
nand U14822 (N_14822,N_13476,N_13688);
or U14823 (N_14823,N_13149,N_13302);
xor U14824 (N_14824,N_13191,N_12657);
or U14825 (N_14825,N_13577,N_13036);
nor U14826 (N_14826,N_13425,N_12538);
nand U14827 (N_14827,N_13582,N_13201);
or U14828 (N_14828,N_12581,N_13410);
and U14829 (N_14829,N_13377,N_13509);
and U14830 (N_14830,N_12781,N_12615);
and U14831 (N_14831,N_13389,N_13443);
nor U14832 (N_14832,N_13226,N_13506);
nand U14833 (N_14833,N_13136,N_12821);
xor U14834 (N_14834,N_12577,N_13445);
nand U14835 (N_14835,N_13683,N_13440);
and U14836 (N_14836,N_13060,N_13625);
nor U14837 (N_14837,N_12965,N_13355);
nand U14838 (N_14838,N_13145,N_12935);
xnor U14839 (N_14839,N_13125,N_13030);
nand U14840 (N_14840,N_13328,N_13563);
nor U14841 (N_14841,N_12795,N_13622);
and U14842 (N_14842,N_13368,N_13377);
nand U14843 (N_14843,N_13694,N_12971);
nand U14844 (N_14844,N_13248,N_12767);
and U14845 (N_14845,N_13277,N_13649);
and U14846 (N_14846,N_13586,N_13676);
nand U14847 (N_14847,N_13188,N_12691);
and U14848 (N_14848,N_12964,N_13473);
nand U14849 (N_14849,N_13628,N_13668);
nor U14850 (N_14850,N_12811,N_12612);
or U14851 (N_14851,N_13086,N_13180);
xor U14852 (N_14852,N_13411,N_13185);
nand U14853 (N_14853,N_13605,N_12671);
nand U14854 (N_14854,N_13300,N_13502);
nor U14855 (N_14855,N_13181,N_12913);
nor U14856 (N_14856,N_13719,N_12949);
and U14857 (N_14857,N_12806,N_13086);
and U14858 (N_14858,N_13675,N_12583);
and U14859 (N_14859,N_12597,N_13173);
or U14860 (N_14860,N_12641,N_13307);
nand U14861 (N_14861,N_13385,N_13021);
nor U14862 (N_14862,N_12596,N_13602);
xor U14863 (N_14863,N_13194,N_12713);
xnor U14864 (N_14864,N_12653,N_13297);
nand U14865 (N_14865,N_13265,N_12699);
or U14866 (N_14866,N_12538,N_13414);
xnor U14867 (N_14867,N_12986,N_12770);
nand U14868 (N_14868,N_13187,N_13099);
xor U14869 (N_14869,N_13727,N_13221);
nor U14870 (N_14870,N_13415,N_13749);
xnor U14871 (N_14871,N_12530,N_12724);
or U14872 (N_14872,N_13143,N_13126);
nand U14873 (N_14873,N_13338,N_13420);
xor U14874 (N_14874,N_12538,N_12957);
nor U14875 (N_14875,N_13499,N_13695);
xnor U14876 (N_14876,N_12974,N_13254);
nand U14877 (N_14877,N_13738,N_13439);
and U14878 (N_14878,N_12762,N_12522);
or U14879 (N_14879,N_13597,N_13728);
nor U14880 (N_14880,N_12666,N_13167);
nor U14881 (N_14881,N_12845,N_13452);
xor U14882 (N_14882,N_12874,N_13318);
or U14883 (N_14883,N_13661,N_13618);
nand U14884 (N_14884,N_13542,N_13180);
and U14885 (N_14885,N_13108,N_13313);
and U14886 (N_14886,N_13244,N_13594);
and U14887 (N_14887,N_13667,N_12794);
nand U14888 (N_14888,N_12931,N_12997);
xor U14889 (N_14889,N_13178,N_12998);
xnor U14890 (N_14890,N_12538,N_13408);
nand U14891 (N_14891,N_13642,N_13563);
and U14892 (N_14892,N_13208,N_12543);
and U14893 (N_14893,N_13738,N_13300);
nor U14894 (N_14894,N_13598,N_12812);
xnor U14895 (N_14895,N_12685,N_13276);
and U14896 (N_14896,N_12612,N_13347);
and U14897 (N_14897,N_12823,N_13548);
nand U14898 (N_14898,N_12739,N_13025);
xnor U14899 (N_14899,N_12681,N_12829);
nand U14900 (N_14900,N_12823,N_13016);
nor U14901 (N_14901,N_13437,N_13200);
and U14902 (N_14902,N_13268,N_13554);
nand U14903 (N_14903,N_13687,N_13360);
xor U14904 (N_14904,N_12943,N_12998);
nand U14905 (N_14905,N_13368,N_13231);
nor U14906 (N_14906,N_12742,N_13529);
or U14907 (N_14907,N_13512,N_13146);
and U14908 (N_14908,N_13621,N_12848);
and U14909 (N_14909,N_13630,N_13647);
xnor U14910 (N_14910,N_12673,N_12637);
or U14911 (N_14911,N_13692,N_12853);
nor U14912 (N_14912,N_13381,N_12708);
and U14913 (N_14913,N_13290,N_13089);
xnor U14914 (N_14914,N_12639,N_13118);
and U14915 (N_14915,N_12951,N_13589);
nand U14916 (N_14916,N_12651,N_12692);
and U14917 (N_14917,N_13297,N_13518);
xor U14918 (N_14918,N_12612,N_13482);
or U14919 (N_14919,N_13410,N_12697);
nand U14920 (N_14920,N_13162,N_13709);
nand U14921 (N_14921,N_13302,N_13156);
xnor U14922 (N_14922,N_12943,N_12847);
and U14923 (N_14923,N_13047,N_12827);
and U14924 (N_14924,N_13551,N_13497);
xnor U14925 (N_14925,N_13010,N_13604);
and U14926 (N_14926,N_13503,N_13138);
or U14927 (N_14927,N_12853,N_13460);
nor U14928 (N_14928,N_12840,N_12666);
and U14929 (N_14929,N_12848,N_13062);
xor U14930 (N_14930,N_12781,N_13021);
or U14931 (N_14931,N_12754,N_13218);
nor U14932 (N_14932,N_13480,N_12649);
nand U14933 (N_14933,N_13559,N_13153);
nor U14934 (N_14934,N_12920,N_12753);
nor U14935 (N_14935,N_13165,N_13386);
or U14936 (N_14936,N_13721,N_13158);
or U14937 (N_14937,N_12561,N_12556);
nor U14938 (N_14938,N_13554,N_12986);
xnor U14939 (N_14939,N_12517,N_13279);
nor U14940 (N_14940,N_13229,N_13387);
or U14941 (N_14941,N_13672,N_12880);
and U14942 (N_14942,N_12667,N_13193);
or U14943 (N_14943,N_13480,N_12782);
nor U14944 (N_14944,N_13124,N_13178);
nor U14945 (N_14945,N_12809,N_12619);
and U14946 (N_14946,N_13247,N_13492);
and U14947 (N_14947,N_13087,N_12964);
nand U14948 (N_14948,N_13247,N_12987);
xnor U14949 (N_14949,N_12932,N_13747);
nor U14950 (N_14950,N_13179,N_13392);
or U14951 (N_14951,N_12963,N_13624);
or U14952 (N_14952,N_12823,N_13107);
nor U14953 (N_14953,N_12543,N_13721);
xor U14954 (N_14954,N_12543,N_12942);
nor U14955 (N_14955,N_12704,N_12515);
or U14956 (N_14956,N_13117,N_13037);
or U14957 (N_14957,N_13591,N_13598);
nor U14958 (N_14958,N_12770,N_13227);
and U14959 (N_14959,N_13008,N_13562);
and U14960 (N_14960,N_13740,N_13486);
nor U14961 (N_14961,N_13344,N_12831);
nand U14962 (N_14962,N_13350,N_13510);
and U14963 (N_14963,N_12694,N_12820);
and U14964 (N_14964,N_13030,N_13060);
nor U14965 (N_14965,N_12786,N_13590);
and U14966 (N_14966,N_13157,N_13321);
nand U14967 (N_14967,N_12760,N_13429);
nand U14968 (N_14968,N_12527,N_12831);
or U14969 (N_14969,N_13066,N_12762);
nor U14970 (N_14970,N_13178,N_12822);
xor U14971 (N_14971,N_12543,N_13247);
nand U14972 (N_14972,N_13678,N_13005);
nand U14973 (N_14973,N_13489,N_12638);
and U14974 (N_14974,N_12640,N_13607);
and U14975 (N_14975,N_12622,N_13259);
or U14976 (N_14976,N_13700,N_13005);
and U14977 (N_14977,N_13691,N_12578);
xnor U14978 (N_14978,N_12810,N_13343);
or U14979 (N_14979,N_13446,N_12704);
nor U14980 (N_14980,N_13345,N_12542);
and U14981 (N_14981,N_13649,N_13666);
or U14982 (N_14982,N_13429,N_13391);
nand U14983 (N_14983,N_13563,N_13365);
xor U14984 (N_14984,N_13215,N_12729);
and U14985 (N_14985,N_13094,N_13003);
nor U14986 (N_14986,N_12530,N_13104);
or U14987 (N_14987,N_12665,N_12867);
and U14988 (N_14988,N_13145,N_12867);
or U14989 (N_14989,N_13092,N_13316);
or U14990 (N_14990,N_12584,N_13118);
and U14991 (N_14991,N_12744,N_13711);
nor U14992 (N_14992,N_12661,N_13386);
and U14993 (N_14993,N_13384,N_13273);
and U14994 (N_14994,N_13167,N_13489);
nor U14995 (N_14995,N_13337,N_13445);
and U14996 (N_14996,N_12635,N_13089);
xnor U14997 (N_14997,N_13406,N_12993);
xor U14998 (N_14998,N_13542,N_12997);
nand U14999 (N_14999,N_13608,N_13462);
nand U15000 (N_15000,N_14377,N_14130);
nand U15001 (N_15001,N_14892,N_13801);
or U15002 (N_15002,N_13880,N_13773);
and U15003 (N_15003,N_14072,N_14161);
xor U15004 (N_15004,N_14766,N_14959);
nor U15005 (N_15005,N_14156,N_14250);
nand U15006 (N_15006,N_14327,N_14822);
and U15007 (N_15007,N_14466,N_14227);
and U15008 (N_15008,N_14106,N_14011);
and U15009 (N_15009,N_14095,N_14748);
or U15010 (N_15010,N_14331,N_14303);
or U15011 (N_15011,N_14527,N_13938);
and U15012 (N_15012,N_14253,N_13785);
nand U15013 (N_15013,N_14512,N_14643);
nand U15014 (N_15014,N_14413,N_13949);
and U15015 (N_15015,N_13817,N_14808);
or U15016 (N_15016,N_14739,N_14368);
nand U15017 (N_15017,N_14670,N_14387);
xor U15018 (N_15018,N_14674,N_14017);
and U15019 (N_15019,N_14942,N_14563);
xnor U15020 (N_15020,N_14223,N_14775);
xor U15021 (N_15021,N_14247,N_14367);
nand U15022 (N_15022,N_13999,N_14960);
and U15023 (N_15023,N_14847,N_14186);
xor U15024 (N_15024,N_14166,N_14526);
nor U15025 (N_15025,N_13946,N_14241);
xnor U15026 (N_15026,N_14492,N_14956);
nand U15027 (N_15027,N_14491,N_14213);
nor U15028 (N_15028,N_13859,N_14910);
and U15029 (N_15029,N_14962,N_14977);
and U15030 (N_15030,N_14198,N_13899);
nand U15031 (N_15031,N_14496,N_14647);
and U15032 (N_15032,N_14384,N_14628);
xnor U15033 (N_15033,N_13964,N_14542);
and U15034 (N_15034,N_14278,N_14197);
nand U15035 (N_15035,N_14081,N_14832);
nand U15036 (N_15036,N_14882,N_14583);
and U15037 (N_15037,N_14373,N_14702);
nor U15038 (N_15038,N_14677,N_14454);
nand U15039 (N_15039,N_14571,N_14614);
xnor U15040 (N_15040,N_13853,N_13888);
nor U15041 (N_15041,N_14917,N_14932);
and U15042 (N_15042,N_14435,N_14292);
and U15043 (N_15043,N_13870,N_14562);
nor U15044 (N_15044,N_14530,N_14477);
nor U15045 (N_15045,N_13789,N_14251);
nand U15046 (N_15046,N_14923,N_14124);
xor U15047 (N_15047,N_13778,N_14648);
nor U15048 (N_15048,N_14550,N_14554);
or U15049 (N_15049,N_14979,N_14837);
or U15050 (N_15050,N_14208,N_14729);
or U15051 (N_15051,N_14192,N_14595);
nor U15052 (N_15052,N_14823,N_14934);
and U15053 (N_15053,N_14645,N_14662);
nand U15054 (N_15054,N_14461,N_14844);
and U15055 (N_15055,N_14471,N_14753);
xor U15056 (N_15056,N_14850,N_14694);
nand U15057 (N_15057,N_14267,N_13761);
xnor U15058 (N_15058,N_14099,N_14833);
or U15059 (N_15059,N_14502,N_13944);
nand U15060 (N_15060,N_14743,N_14425);
or U15061 (N_15061,N_14681,N_13786);
xor U15062 (N_15062,N_14980,N_14868);
xor U15063 (N_15063,N_14861,N_13973);
xnor U15064 (N_15064,N_13994,N_14059);
nor U15065 (N_15065,N_14075,N_14196);
nand U15066 (N_15066,N_14481,N_14957);
xor U15067 (N_15067,N_14443,N_14524);
or U15068 (N_15068,N_14122,N_14774);
nor U15069 (N_15069,N_14570,N_14483);
or U15070 (N_15070,N_13928,N_13981);
xor U15071 (N_15071,N_14915,N_14782);
nand U15072 (N_15072,N_14306,N_14310);
xor U15073 (N_15073,N_14045,N_14079);
and U15074 (N_15074,N_13792,N_14133);
and U15075 (N_15075,N_14510,N_14708);
and U15076 (N_15076,N_14768,N_14544);
xor U15077 (N_15077,N_14061,N_14796);
and U15078 (N_15078,N_14812,N_13961);
nor U15079 (N_15079,N_14069,N_14943);
nand U15080 (N_15080,N_14027,N_14255);
xor U15081 (N_15081,N_14245,N_14324);
or U15082 (N_15082,N_14528,N_14233);
or U15083 (N_15083,N_13958,N_14888);
nand U15084 (N_15084,N_14394,N_14919);
and U15085 (N_15085,N_14288,N_14579);
or U15086 (N_15086,N_13919,N_14020);
and U15087 (N_15087,N_14236,N_14189);
xor U15088 (N_15088,N_14577,N_14553);
and U15089 (N_15089,N_14346,N_14063);
and U15090 (N_15090,N_14030,N_13871);
xor U15091 (N_15091,N_14220,N_14048);
nor U15092 (N_15092,N_14565,N_14918);
xor U15093 (N_15093,N_14127,N_14440);
or U15094 (N_15094,N_14449,N_14826);
and U15095 (N_15095,N_14938,N_13916);
and U15096 (N_15096,N_14884,N_13766);
nor U15097 (N_15097,N_14043,N_14723);
or U15098 (N_15098,N_14193,N_14347);
xnor U15099 (N_15099,N_14088,N_14684);
nor U15100 (N_15100,N_14871,N_14286);
nor U15101 (N_15101,N_13953,N_14916);
and U15102 (N_15102,N_14644,N_14839);
nor U15103 (N_15103,N_14037,N_14689);
nor U15104 (N_15104,N_14653,N_14005);
and U15105 (N_15105,N_14561,N_14931);
xnor U15106 (N_15106,N_14363,N_14200);
nor U15107 (N_15107,N_14448,N_14627);
and U15108 (N_15108,N_13765,N_14572);
or U15109 (N_15109,N_13816,N_14487);
or U15110 (N_15110,N_13767,N_14412);
nor U15111 (N_15111,N_14479,N_14770);
nor U15112 (N_15112,N_13950,N_14682);
nor U15113 (N_15113,N_14971,N_14110);
and U15114 (N_15114,N_14358,N_14569);
or U15115 (N_15115,N_14795,N_13863);
xor U15116 (N_15116,N_13759,N_13912);
nor U15117 (N_15117,N_14473,N_14285);
nor U15118 (N_15118,N_14246,N_14460);
nor U15119 (N_15119,N_14118,N_14700);
or U15120 (N_15120,N_14042,N_14187);
and U15121 (N_15121,N_14534,N_14108);
nand U15122 (N_15122,N_14361,N_14104);
or U15123 (N_15123,N_14873,N_14747);
and U15124 (N_15124,N_14096,N_13796);
xnor U15125 (N_15125,N_13827,N_14013);
nor U15126 (N_15126,N_13891,N_13934);
xor U15127 (N_15127,N_14704,N_14340);
and U15128 (N_15128,N_13830,N_13810);
xor U15129 (N_15129,N_13790,N_14863);
nand U15130 (N_15130,N_14312,N_14835);
nor U15131 (N_15131,N_14998,N_13972);
xnor U15132 (N_15132,N_14274,N_14378);
xnor U15133 (N_15133,N_14060,N_14764);
or U15134 (N_15134,N_13892,N_14854);
and U15135 (N_15135,N_13832,N_14556);
xor U15136 (N_15136,N_14411,N_14893);
and U15137 (N_15137,N_14777,N_14344);
xor U15138 (N_15138,N_14343,N_14986);
or U15139 (N_15139,N_13879,N_14325);
nand U15140 (N_15140,N_14589,N_14781);
nand U15141 (N_15141,N_14678,N_14867);
xor U15142 (N_15142,N_14194,N_14874);
or U15143 (N_15143,N_14121,N_13868);
nor U15144 (N_15144,N_14791,N_14800);
xor U15145 (N_15145,N_14172,N_13775);
and U15146 (N_15146,N_14876,N_14604);
nor U15147 (N_15147,N_14168,N_13997);
nand U15148 (N_15148,N_13940,N_14615);
or U15149 (N_15149,N_14984,N_14594);
xnor U15150 (N_15150,N_14687,N_13768);
nor U15151 (N_15151,N_13846,N_14907);
nand U15152 (N_15152,N_14203,N_14804);
or U15153 (N_15153,N_14933,N_14457);
or U15154 (N_15154,N_14276,N_14596);
nor U15155 (N_15155,N_14222,N_13809);
or U15156 (N_15156,N_14997,N_13758);
xor U15157 (N_15157,N_13908,N_14281);
and U15158 (N_15158,N_13931,N_14329);
xnor U15159 (N_15159,N_14319,N_14624);
and U15160 (N_15160,N_14388,N_14975);
and U15161 (N_15161,N_13776,N_13962);
and U15162 (N_15162,N_14925,N_14727);
nor U15163 (N_15163,N_14032,N_14629);
nor U15164 (N_15164,N_14031,N_14299);
or U15165 (N_15165,N_14607,N_14307);
nand U15166 (N_15166,N_13788,N_14398);
and U15167 (N_15167,N_13992,N_14654);
or U15168 (N_15168,N_14955,N_14283);
nor U15169 (N_15169,N_14982,N_14851);
nand U15170 (N_15170,N_14738,N_14153);
and U15171 (N_15171,N_14901,N_13866);
or U15172 (N_15172,N_14947,N_14406);
or U15173 (N_15173,N_14086,N_14191);
xnor U15174 (N_15174,N_14831,N_14146);
nand U15175 (N_15175,N_14183,N_14599);
and U15176 (N_15176,N_13894,N_14698);
or U15177 (N_15177,N_14951,N_13861);
nand U15178 (N_15178,N_14707,N_14869);
nor U15179 (N_15179,N_14545,N_14484);
xnor U15180 (N_15180,N_14778,N_14875);
and U15181 (N_15181,N_14602,N_14269);
or U15182 (N_15182,N_14459,N_14248);
and U15183 (N_15183,N_14590,N_13836);
nand U15184 (N_15184,N_13814,N_13925);
xor U15185 (N_15185,N_13967,N_14260);
and U15186 (N_15186,N_13904,N_13875);
xor U15187 (N_15187,N_13918,N_14294);
and U15188 (N_15188,N_13823,N_14452);
nand U15189 (N_15189,N_14547,N_13913);
and U15190 (N_15190,N_13865,N_14016);
and U15191 (N_15191,N_14098,N_13885);
xnor U15192 (N_15192,N_14143,N_14859);
nor U15193 (N_15193,N_14878,N_14315);
nand U15194 (N_15194,N_14639,N_14243);
xor U15195 (N_15195,N_14455,N_14488);
and U15196 (N_15196,N_13835,N_14410);
nand U15197 (N_15197,N_14828,N_13869);
xor U15198 (N_15198,N_14439,N_13771);
and U15199 (N_15199,N_14040,N_14848);
nor U15200 (N_15200,N_14320,N_14858);
nand U15201 (N_15201,N_14830,N_14620);
or U15202 (N_15202,N_14334,N_14752);
xor U15203 (N_15203,N_14428,N_13898);
or U15204 (N_15204,N_14621,N_13858);
nand U15205 (N_15205,N_14225,N_14478);
nor U15206 (N_15206,N_13848,N_14009);
and U15207 (N_15207,N_13808,N_13985);
xor U15208 (N_15208,N_14903,N_14497);
nand U15209 (N_15209,N_14806,N_13815);
nor U15210 (N_15210,N_14637,N_14877);
xnor U15211 (N_15211,N_14275,N_14055);
xor U15212 (N_15212,N_13797,N_14360);
and U15213 (N_15213,N_14817,N_14548);
and U15214 (N_15214,N_14807,N_13829);
xnor U15215 (N_15215,N_14789,N_14372);
nand U15216 (N_15216,N_14033,N_14675);
nand U15217 (N_15217,N_14619,N_14746);
xor U15218 (N_15218,N_14966,N_14963);
xor U15219 (N_15219,N_14287,N_13942);
nand U15220 (N_15220,N_14350,N_14612);
nand U15221 (N_15221,N_14772,N_14588);
nand U15222 (N_15222,N_13878,N_14935);
or U15223 (N_15223,N_14207,N_13837);
nor U15224 (N_15224,N_14002,N_13840);
xor U15225 (N_15225,N_14936,N_14083);
nand U15226 (N_15226,N_14638,N_14750);
xor U15227 (N_15227,N_14177,N_14018);
and U15228 (N_15228,N_14676,N_13939);
or U15229 (N_15229,N_14865,N_14761);
and U15230 (N_15230,N_13951,N_14685);
and U15231 (N_15231,N_14318,N_14610);
nand U15232 (N_15232,N_14890,N_14745);
xor U15233 (N_15233,N_14948,N_14149);
nor U15234 (N_15234,N_14190,N_14945);
and U15235 (N_15235,N_14231,N_14272);
nor U15236 (N_15236,N_14714,N_14580);
and U15237 (N_15237,N_14719,N_14541);
xor U15238 (N_15238,N_14365,N_14148);
xnor U15239 (N_15239,N_14311,N_14741);
or U15240 (N_15240,N_14924,N_13849);
or U15241 (N_15241,N_14516,N_13911);
xnor U15242 (N_15242,N_14995,N_14721);
nor U15243 (N_15243,N_14605,N_13791);
and U15244 (N_15244,N_14129,N_14001);
or U15245 (N_15245,N_14686,N_14463);
and U15246 (N_15246,N_14429,N_13847);
nor U15247 (N_15247,N_14843,N_13860);
xnor U15248 (N_15248,N_14558,N_14603);
xnor U15249 (N_15249,N_14493,N_14976);
and U15250 (N_15250,N_13993,N_14758);
xor U15251 (N_15251,N_14169,N_14337);
or U15252 (N_15252,N_13845,N_13872);
nor U15253 (N_15253,N_14392,N_14751);
or U15254 (N_15254,N_13965,N_14170);
nor U15255 (N_15255,N_14824,N_14038);
nand U15256 (N_15256,N_13757,N_14444);
nand U15257 (N_15257,N_14374,N_13924);
and U15258 (N_15258,N_13915,N_13754);
nor U15259 (N_15259,N_14180,N_14840);
nor U15260 (N_15260,N_14173,N_13784);
nand U15261 (N_15261,N_14887,N_14370);
or U15262 (N_15262,N_14116,N_14798);
and U15263 (N_15263,N_14206,N_14631);
xnor U15264 (N_15264,N_14134,N_14323);
nor U15265 (N_15265,N_14147,N_13976);
nor U15266 (N_15266,N_14703,N_14866);
xor U15267 (N_15267,N_14926,N_13864);
xor U15268 (N_15268,N_14505,N_14341);
or U15269 (N_15269,N_14717,N_14154);
nand U15270 (N_15270,N_14224,N_13900);
nand U15271 (N_15271,N_13983,N_13929);
nand U15272 (N_15272,N_14913,N_14262);
xor U15273 (N_15273,N_14242,N_13751);
nand U15274 (N_15274,N_14845,N_14691);
xor U15275 (N_15275,N_14762,N_14567);
or U15276 (N_15276,N_14386,N_14776);
nand U15277 (N_15277,N_14132,N_14280);
nor U15278 (N_15278,N_14298,N_14950);
nor U15279 (N_15279,N_14578,N_14423);
nor U15280 (N_15280,N_14852,N_14810);
nand U15281 (N_15281,N_14357,N_13977);
xor U15282 (N_15282,N_14065,N_14827);
nand U15283 (N_15283,N_14507,N_14765);
or U15284 (N_15284,N_14724,N_13881);
or U15285 (N_15285,N_13920,N_14073);
xor U15286 (N_15286,N_13980,N_14531);
or U15287 (N_15287,N_14176,N_14632);
nor U15288 (N_15288,N_14171,N_14238);
nor U15289 (N_15289,N_14862,N_14792);
nand U15290 (N_15290,N_14725,N_14606);
and U15291 (N_15291,N_14586,N_14829);
xnor U15292 (N_15292,N_14983,N_13782);
and U15293 (N_15293,N_14181,N_14585);
and U15294 (N_15294,N_14652,N_14097);
nand U15295 (N_15295,N_14517,N_14601);
nand U15296 (N_15296,N_13959,N_14633);
and U15297 (N_15297,N_14404,N_13851);
xor U15298 (N_15298,N_14201,N_13855);
xnor U15299 (N_15299,N_14515,N_14137);
or U15300 (N_15300,N_14399,N_13831);
and U15301 (N_15301,N_14119,N_13932);
nor U15302 (N_15302,N_14237,N_14266);
nand U15303 (N_15303,N_14113,N_13971);
nand U15304 (N_15304,N_14560,N_14611);
or U15305 (N_15305,N_14591,N_13753);
xnor U15306 (N_15306,N_14825,N_13905);
nand U15307 (N_15307,N_14911,N_14366);
xnor U15308 (N_15308,N_14513,N_13937);
nor U15309 (N_15309,N_13843,N_14905);
or U15310 (N_15310,N_14336,N_13818);
and U15311 (N_15311,N_14426,N_13807);
nand U15312 (N_15312,N_14369,N_13945);
or U15313 (N_15313,N_14634,N_13798);
nand U15314 (N_15314,N_14114,N_14939);
and U15315 (N_15315,N_14408,N_13780);
xnor U15316 (N_15316,N_13897,N_14989);
nor U15317 (N_15317,N_14141,N_13895);
nand U15318 (N_15318,N_14819,N_14785);
nor U15319 (N_15319,N_14195,N_14218);
or U15320 (N_15320,N_14927,N_14480);
xor U15321 (N_15321,N_13856,N_14179);
nand U15322 (N_15322,N_14872,N_14418);
or U15323 (N_15323,N_14749,N_14050);
xnor U15324 (N_15324,N_14023,N_13833);
nand U15325 (N_15325,N_14744,N_14068);
and U15326 (N_15326,N_14380,N_14103);
xor U15327 (N_15327,N_14351,N_14111);
or U15328 (N_15328,N_14811,N_13910);
or U15329 (N_15329,N_13794,N_14431);
and U15330 (N_15330,N_13922,N_14453);
nor U15331 (N_15331,N_14029,N_14420);
or U15332 (N_15332,N_14474,N_14209);
nor U15333 (N_15333,N_14093,N_14402);
xor U15334 (N_15334,N_13844,N_14978);
nor U15335 (N_15335,N_14150,N_14259);
nor U15336 (N_15336,N_14937,N_14462);
nor U15337 (N_15337,N_14080,N_14219);
xor U15338 (N_15338,N_14482,N_14472);
xnor U15339 (N_15339,N_14308,N_14291);
or U15340 (N_15340,N_14974,N_13986);
nand U15341 (N_15341,N_14036,N_13854);
xor U15342 (N_15342,N_13991,N_14450);
or U15343 (N_15343,N_14265,N_13862);
or U15344 (N_15344,N_14441,N_14159);
and U15345 (N_15345,N_13806,N_14886);
and U15346 (N_15346,N_14967,N_14089);
nor U15347 (N_15347,N_14834,N_13764);
and U15348 (N_15348,N_13963,N_14330);
or U15349 (N_15349,N_14519,N_14359);
and U15350 (N_15350,N_14309,N_14092);
xnor U15351 (N_15351,N_14232,N_13822);
xnor U15352 (N_15352,N_14688,N_14077);
nand U15353 (N_15353,N_13996,N_14381);
nor U15354 (N_15354,N_14658,N_14338);
nor U15355 (N_15355,N_14445,N_13874);
nor U15356 (N_15356,N_14379,N_13889);
nor U15357 (N_15357,N_14794,N_14897);
nand U15358 (N_15358,N_14635,N_13954);
nand U15359 (N_15359,N_13941,N_14314);
xnor U15360 (N_15360,N_14944,N_13795);
nor U15361 (N_15361,N_14434,N_13995);
or U15362 (N_15362,N_13850,N_14067);
xor U15363 (N_15363,N_14709,N_14102);
xnor U15364 (N_15364,N_14880,N_13783);
and U15365 (N_15365,N_14657,N_14417);
or U15366 (N_15366,N_14949,N_13909);
and U15367 (N_15367,N_13984,N_13756);
and U15368 (N_15368,N_14415,N_14609);
nand U15369 (N_15369,N_14718,N_14400);
nand U15370 (N_15370,N_14212,N_13752);
or U15371 (N_15371,N_14906,N_14458);
xnor U15372 (N_15372,N_14818,N_14349);
or U15373 (N_15373,N_14304,N_14053);
or U15374 (N_15374,N_14442,N_14742);
xnor U15375 (N_15375,N_14598,N_14740);
or U15376 (N_15376,N_14722,N_14712);
xor U15377 (N_15377,N_14049,N_14131);
or U15378 (N_15378,N_14522,N_14467);
or U15379 (N_15379,N_14640,N_13998);
nand U15380 (N_15380,N_14249,N_14991);
xor U15381 (N_15381,N_14814,N_14405);
or U15382 (N_15382,N_14221,N_14326);
nor U15383 (N_15383,N_13926,N_14870);
xnor U15384 (N_15384,N_14279,N_13821);
and U15385 (N_15385,N_14587,N_14904);
nand U15386 (N_15386,N_14205,N_14529);
nand U15387 (N_15387,N_14328,N_13811);
and U15388 (N_15388,N_14564,N_14074);
nand U15389 (N_15389,N_14566,N_14855);
xor U15390 (N_15390,N_13857,N_14115);
and U15391 (N_15391,N_14503,N_14779);
nor U15392 (N_15392,N_14885,N_13947);
xor U15393 (N_15393,N_14650,N_14557);
xor U15394 (N_15394,N_14470,N_13763);
nand U15395 (N_15395,N_14371,N_13828);
and U15396 (N_15396,N_14549,N_13907);
xor U15397 (N_15397,N_14625,N_14821);
nor U15398 (N_15398,N_14987,N_14123);
nand U15399 (N_15399,N_14446,N_13774);
or U15400 (N_15400,N_14856,N_14409);
nor U15401 (N_15401,N_14695,N_14403);
and U15402 (N_15402,N_14720,N_13988);
and U15403 (N_15403,N_14070,N_14297);
or U15404 (N_15404,N_14756,N_14052);
xor U15405 (N_15405,N_14864,N_14805);
xor U15406 (N_15406,N_14999,N_13884);
or U15407 (N_15407,N_14401,N_14552);
or U15408 (N_15408,N_14165,N_14921);
nor U15409 (N_15409,N_13873,N_14395);
or U15410 (N_15410,N_14575,N_14755);
and U15411 (N_15411,N_14651,N_14393);
xnor U15412 (N_15412,N_13772,N_14846);
nand U15413 (N_15413,N_14432,N_14706);
nor U15414 (N_15414,N_14282,N_14693);
nor U15415 (N_15415,N_14985,N_14801);
and U15416 (N_15416,N_14551,N_14316);
nand U15417 (N_15417,N_14214,N_14254);
nand U15418 (N_15418,N_14954,N_14626);
or U15419 (N_15419,N_14896,N_14574);
or U15420 (N_15420,N_14773,N_14797);
and U15421 (N_15421,N_14353,N_14382);
nor U15422 (N_15422,N_13969,N_14202);
nor U15423 (N_15423,N_14641,N_14289);
and U15424 (N_15424,N_14486,N_14229);
and U15425 (N_15425,N_14760,N_14041);
xnor U15426 (N_15426,N_14012,N_14414);
or U15427 (N_15427,N_14784,N_14385);
nand U15428 (N_15428,N_14623,N_14390);
or U15429 (N_15429,N_14815,N_14849);
and U15430 (N_15430,N_13877,N_14010);
or U15431 (N_15431,N_13979,N_14965);
or U15432 (N_15432,N_13803,N_14047);
nand U15433 (N_15433,N_14216,N_14174);
nand U15434 (N_15434,N_14489,N_13883);
and U15435 (N_15435,N_13970,N_14953);
nand U15436 (N_15436,N_14264,N_14961);
xor U15437 (N_15437,N_14696,N_13750);
nor U15438 (N_15438,N_14433,N_14930);
xnor U15439 (N_15439,N_14900,N_14252);
nand U15440 (N_15440,N_14771,N_14090);
or U15441 (N_15441,N_14754,N_14922);
xnor U15442 (N_15442,N_14535,N_14391);
nand U15443 (N_15443,N_14669,N_14780);
and U15444 (N_15444,N_13902,N_14451);
or U15445 (N_15445,N_13805,N_14107);
or U15446 (N_15446,N_14793,N_14284);
or U15447 (N_15447,N_13887,N_14485);
xnor U15448 (N_15448,N_14204,N_14523);
xnor U15449 (N_15449,N_14671,N_14759);
or U15450 (N_15450,N_14345,N_13930);
and U15451 (N_15451,N_14582,N_14790);
nor U15452 (N_15452,N_13957,N_14144);
or U15453 (N_15453,N_14271,N_14783);
nand U15454 (N_15454,N_14160,N_14022);
nor U15455 (N_15455,N_14164,N_14736);
nand U15456 (N_15456,N_14138,N_13839);
nor U15457 (N_15457,N_14539,N_14139);
xnor U15458 (N_15458,N_14397,N_14142);
or U15459 (N_15459,N_14665,N_14375);
nor U15460 (N_15460,N_14447,N_14716);
nor U15461 (N_15461,N_14014,N_13935);
xnor U15462 (N_15462,N_14199,N_13927);
xnor U15463 (N_15463,N_13812,N_14317);
nand U15464 (N_15464,N_14508,N_14407);
or U15465 (N_15465,N_13813,N_14655);
xnor U15466 (N_15466,N_14617,N_14973);
nor U15467 (N_15467,N_14051,N_14690);
nor U15468 (N_15468,N_13952,N_14642);
nor U15469 (N_15469,N_14568,N_13943);
or U15470 (N_15470,N_14813,N_14734);
xnor U15471 (N_15471,N_13799,N_13968);
and U15472 (N_15472,N_13914,N_14416);
and U15473 (N_15473,N_13901,N_14498);
or U15474 (N_15474,N_14732,N_14573);
nand U15475 (N_15475,N_14469,N_14841);
nor U15476 (N_15476,N_14711,N_14920);
xnor U15477 (N_15477,N_14091,N_13906);
nand U15478 (N_15478,N_14664,N_14889);
nand U15479 (N_15479,N_14763,N_14348);
xor U15480 (N_15480,N_14333,N_13826);
xnor U15481 (N_15481,N_14842,N_14659);
or U15482 (N_15482,N_14618,N_14125);
nor U15483 (N_15483,N_13800,N_13755);
nand U15484 (N_15484,N_13989,N_14256);
and U15485 (N_15485,N_14699,N_14737);
nand U15486 (N_15486,N_14799,N_14940);
or U15487 (N_15487,N_14071,N_14364);
nand U15488 (N_15488,N_13867,N_14438);
nand U15489 (N_15489,N_14185,N_14680);
nor U15490 (N_15490,N_14543,N_13777);
nor U15491 (N_15491,N_14518,N_14015);
and U15492 (N_15492,N_13876,N_14354);
nor U15493 (N_15493,N_14769,N_13842);
or U15494 (N_15494,N_13933,N_14993);
or U15495 (N_15495,N_14511,N_14581);
or U15496 (N_15496,N_14057,N_14475);
nand U15497 (N_15497,N_14733,N_14273);
nand U15498 (N_15498,N_14321,N_14019);
nand U15499 (N_15499,N_14085,N_14056);
and U15500 (N_15500,N_14158,N_14305);
xnor U15501 (N_15501,N_14035,N_14342);
nand U15502 (N_15502,N_13974,N_14094);
nand U15503 (N_15503,N_14234,N_14217);
and U15504 (N_15504,N_14902,N_14101);
or U15505 (N_15505,N_14836,N_14257);
or U15506 (N_15506,N_13779,N_14046);
or U15507 (N_15507,N_14263,N_14521);
nor U15508 (N_15508,N_14895,N_14100);
nand U15509 (N_15509,N_14235,N_14788);
nor U15510 (N_15510,N_14356,N_14468);
or U15511 (N_15511,N_14383,N_14476);
nand U15512 (N_15512,N_14820,N_14538);
nand U15513 (N_15513,N_13917,N_14649);
xnor U15514 (N_15514,N_14663,N_14167);
nand U15515 (N_15515,N_14490,N_14616);
nor U15516 (N_15516,N_14697,N_14994);
and U15517 (N_15517,N_14302,N_13921);
and U15518 (N_15518,N_14087,N_14853);
nor U15519 (N_15519,N_14593,N_14240);
nand U15520 (N_15520,N_14525,N_14182);
or U15521 (N_15521,N_13781,N_14728);
or U15522 (N_15522,N_13903,N_14301);
or U15523 (N_15523,N_14128,N_14152);
and U15524 (N_15524,N_14613,N_14026);
and U15525 (N_15525,N_14008,N_14514);
xor U15526 (N_15526,N_14226,N_14389);
nor U15527 (N_15527,N_14679,N_14003);
or U15528 (N_15528,N_14230,N_13787);
xor U15529 (N_15529,N_14105,N_13990);
or U15530 (N_15530,N_14816,N_14912);
and U15531 (N_15531,N_14968,N_14456);
and U15532 (N_15532,N_13825,N_14914);
nand U15533 (N_15533,N_14726,N_14120);
xnor U15534 (N_15534,N_13770,N_14891);
and U15535 (N_15535,N_13802,N_14546);
xnor U15536 (N_15536,N_14044,N_13834);
and U15537 (N_15537,N_14536,N_14430);
nand U15538 (N_15538,N_14715,N_14537);
or U15539 (N_15539,N_14767,N_13760);
xor U15540 (N_15540,N_14972,N_14290);
xnor U15541 (N_15541,N_14064,N_13923);
and U15542 (N_15542,N_14710,N_14066);
and U15543 (N_15543,N_14597,N_14970);
and U15544 (N_15544,N_13886,N_13841);
nor U15545 (N_15545,N_14188,N_14039);
and U15546 (N_15546,N_14660,N_14000);
nor U15547 (N_15547,N_14136,N_14058);
nand U15548 (N_15548,N_14028,N_14540);
xnor U15549 (N_15549,N_14178,N_14082);
xor U15550 (N_15550,N_14355,N_14929);
nor U15551 (N_15551,N_14054,N_14600);
and U15552 (N_15552,N_13960,N_14509);
nor U15553 (N_15553,N_14495,N_14163);
xnor U15554 (N_15554,N_14899,N_14946);
nor U15555 (N_15555,N_14809,N_13882);
xnor U15556 (N_15556,N_14270,N_14730);
or U15557 (N_15557,N_14084,N_14898);
nor U15558 (N_15558,N_14332,N_13852);
and U15559 (N_15559,N_14004,N_14731);
or U15560 (N_15560,N_14608,N_14135);
and U15561 (N_15561,N_14713,N_14668);
nor U15562 (N_15562,N_14112,N_13893);
nand U15563 (N_15563,N_14622,N_13793);
and U15564 (N_15564,N_14992,N_14928);
nand U15565 (N_15565,N_14559,N_14941);
nor U15566 (N_15566,N_14667,N_14883);
xnor U15567 (N_15567,N_14296,N_13819);
nand U15568 (N_15568,N_14261,N_14661);
or U15569 (N_15569,N_14860,N_14215);
and U15570 (N_15570,N_14145,N_14990);
nor U15571 (N_15571,N_14656,N_14175);
nand U15572 (N_15572,N_13762,N_13769);
nor U15573 (N_15573,N_14436,N_13838);
and U15574 (N_15574,N_14062,N_14157);
nand U15575 (N_15575,N_14024,N_14427);
nor U15576 (N_15576,N_14313,N_13987);
xnor U15577 (N_15577,N_14630,N_14211);
xnor U15578 (N_15578,N_13966,N_14838);
or U15579 (N_15579,N_14692,N_14636);
or U15580 (N_15580,N_14021,N_13936);
or U15581 (N_15581,N_14964,N_14421);
or U15582 (N_15582,N_14076,N_14437);
or U15583 (N_15583,N_14909,N_14646);
or U15584 (N_15584,N_14396,N_14424);
nand U15585 (N_15585,N_14705,N_14683);
nand U15586 (N_15586,N_14576,N_13804);
xnor U15587 (N_15587,N_14422,N_14555);
nand U15588 (N_15588,N_14464,N_14802);
and U15589 (N_15589,N_14504,N_14151);
and U15590 (N_15590,N_13896,N_13824);
nor U15591 (N_15591,N_14735,N_14025);
and U15592 (N_15592,N_14109,N_13955);
or U15593 (N_15593,N_14352,N_14757);
nor U15594 (N_15594,N_14162,N_14339);
or U15595 (N_15595,N_14584,N_14857);
or U15596 (N_15596,N_14533,N_14500);
or U15597 (N_15597,N_14499,N_14672);
and U15598 (N_15598,N_14981,N_14908);
or U15599 (N_15599,N_14952,N_14520);
nand U15600 (N_15600,N_14673,N_13956);
xnor U15601 (N_15601,N_14117,N_13948);
nand U15602 (N_15602,N_14293,N_13975);
or U15603 (N_15603,N_13890,N_14666);
xor U15604 (N_15604,N_14988,N_14268);
and U15605 (N_15605,N_14786,N_14007);
xor U15606 (N_15606,N_14295,N_14006);
nand U15607 (N_15607,N_14034,N_14494);
and U15608 (N_15608,N_14376,N_14465);
nor U15609 (N_15609,N_13982,N_13820);
xor U15610 (N_15610,N_14300,N_14210);
and U15611 (N_15611,N_14958,N_14184);
xnor U15612 (N_15612,N_14155,N_14419);
nor U15613 (N_15613,N_13978,N_14244);
and U15614 (N_15614,N_14532,N_14126);
nor U15615 (N_15615,N_14239,N_14362);
or U15616 (N_15616,N_14506,N_14701);
nand U15617 (N_15617,N_14258,N_14969);
nor U15618 (N_15618,N_14228,N_14881);
nor U15619 (N_15619,N_14277,N_14803);
or U15620 (N_15620,N_14322,N_14501);
and U15621 (N_15621,N_14787,N_14879);
xor U15622 (N_15622,N_14996,N_14592);
nand U15623 (N_15623,N_14140,N_14335);
nand U15624 (N_15624,N_14078,N_14894);
and U15625 (N_15625,N_14629,N_14760);
and U15626 (N_15626,N_14248,N_14851);
and U15627 (N_15627,N_13842,N_14028);
or U15628 (N_15628,N_14707,N_14938);
or U15629 (N_15629,N_13950,N_13994);
and U15630 (N_15630,N_14972,N_14639);
and U15631 (N_15631,N_14562,N_13874);
xnor U15632 (N_15632,N_14911,N_14770);
nor U15633 (N_15633,N_14016,N_14930);
or U15634 (N_15634,N_14086,N_14621);
or U15635 (N_15635,N_13977,N_14286);
or U15636 (N_15636,N_14296,N_14507);
nor U15637 (N_15637,N_14094,N_14272);
nand U15638 (N_15638,N_14477,N_14335);
or U15639 (N_15639,N_14171,N_14762);
xnor U15640 (N_15640,N_14922,N_14411);
and U15641 (N_15641,N_14560,N_14287);
or U15642 (N_15642,N_14325,N_13901);
and U15643 (N_15643,N_14088,N_14215);
nand U15644 (N_15644,N_14324,N_14192);
xnor U15645 (N_15645,N_14985,N_14818);
nand U15646 (N_15646,N_14326,N_14224);
nor U15647 (N_15647,N_13988,N_14864);
nor U15648 (N_15648,N_13952,N_14122);
and U15649 (N_15649,N_13796,N_14845);
nand U15650 (N_15650,N_14030,N_14798);
or U15651 (N_15651,N_14562,N_14717);
and U15652 (N_15652,N_13766,N_14851);
or U15653 (N_15653,N_14416,N_14172);
nor U15654 (N_15654,N_14790,N_13752);
nor U15655 (N_15655,N_14953,N_14339);
nor U15656 (N_15656,N_14301,N_14658);
xor U15657 (N_15657,N_14590,N_14145);
or U15658 (N_15658,N_14772,N_14786);
xnor U15659 (N_15659,N_14268,N_14552);
xnor U15660 (N_15660,N_14554,N_14224);
or U15661 (N_15661,N_13854,N_14786);
nor U15662 (N_15662,N_14374,N_14859);
xnor U15663 (N_15663,N_14603,N_14658);
and U15664 (N_15664,N_13995,N_14017);
or U15665 (N_15665,N_14795,N_14052);
nand U15666 (N_15666,N_14938,N_14817);
and U15667 (N_15667,N_14144,N_14280);
and U15668 (N_15668,N_13946,N_14038);
nor U15669 (N_15669,N_13982,N_14676);
nor U15670 (N_15670,N_14408,N_13796);
and U15671 (N_15671,N_14920,N_14367);
nor U15672 (N_15672,N_14435,N_14617);
xor U15673 (N_15673,N_14653,N_13795);
or U15674 (N_15674,N_14049,N_13864);
nand U15675 (N_15675,N_14030,N_14511);
nor U15676 (N_15676,N_14343,N_14429);
or U15677 (N_15677,N_14075,N_14615);
xnor U15678 (N_15678,N_14160,N_14370);
xor U15679 (N_15679,N_14810,N_14617);
and U15680 (N_15680,N_14682,N_14823);
or U15681 (N_15681,N_14818,N_14078);
nor U15682 (N_15682,N_14659,N_14905);
xnor U15683 (N_15683,N_14411,N_13947);
nor U15684 (N_15684,N_13836,N_13835);
nor U15685 (N_15685,N_13911,N_14899);
and U15686 (N_15686,N_14844,N_14985);
or U15687 (N_15687,N_14481,N_14723);
nand U15688 (N_15688,N_14203,N_14102);
nand U15689 (N_15689,N_14971,N_14579);
and U15690 (N_15690,N_14110,N_13957);
nor U15691 (N_15691,N_14345,N_14442);
xnor U15692 (N_15692,N_14816,N_14254);
or U15693 (N_15693,N_14723,N_14017);
and U15694 (N_15694,N_14605,N_13912);
xor U15695 (N_15695,N_14958,N_14131);
nand U15696 (N_15696,N_13929,N_14452);
xor U15697 (N_15697,N_14372,N_13999);
xnor U15698 (N_15698,N_14427,N_14470);
nand U15699 (N_15699,N_14564,N_14982);
or U15700 (N_15700,N_14365,N_14092);
and U15701 (N_15701,N_14100,N_14364);
nor U15702 (N_15702,N_13873,N_13851);
or U15703 (N_15703,N_14207,N_13909);
nor U15704 (N_15704,N_14704,N_14382);
or U15705 (N_15705,N_14535,N_14520);
or U15706 (N_15706,N_14882,N_14107);
or U15707 (N_15707,N_14854,N_14243);
nand U15708 (N_15708,N_14148,N_14286);
nor U15709 (N_15709,N_14991,N_14620);
nor U15710 (N_15710,N_13991,N_14981);
nor U15711 (N_15711,N_14634,N_14408);
nand U15712 (N_15712,N_13983,N_14451);
nor U15713 (N_15713,N_14846,N_14717);
and U15714 (N_15714,N_13842,N_13825);
nor U15715 (N_15715,N_14218,N_14030);
nor U15716 (N_15716,N_14010,N_13964);
and U15717 (N_15717,N_14786,N_14109);
nand U15718 (N_15718,N_13969,N_14041);
and U15719 (N_15719,N_14295,N_14791);
xnor U15720 (N_15720,N_14807,N_14634);
xnor U15721 (N_15721,N_14450,N_13930);
or U15722 (N_15722,N_14952,N_14747);
and U15723 (N_15723,N_14591,N_13907);
xor U15724 (N_15724,N_14101,N_14031);
nor U15725 (N_15725,N_14268,N_14309);
xnor U15726 (N_15726,N_14758,N_14190);
xor U15727 (N_15727,N_14244,N_13996);
and U15728 (N_15728,N_14625,N_13940);
and U15729 (N_15729,N_14055,N_14625);
and U15730 (N_15730,N_14337,N_14531);
nand U15731 (N_15731,N_13793,N_14058);
nand U15732 (N_15732,N_14343,N_14992);
or U15733 (N_15733,N_14430,N_14743);
and U15734 (N_15734,N_14175,N_14181);
xnor U15735 (N_15735,N_14607,N_14030);
nor U15736 (N_15736,N_14481,N_13953);
or U15737 (N_15737,N_13962,N_13910);
nand U15738 (N_15738,N_14219,N_14289);
nand U15739 (N_15739,N_14897,N_14024);
xnor U15740 (N_15740,N_14466,N_13757);
or U15741 (N_15741,N_13793,N_13965);
nor U15742 (N_15742,N_14789,N_14809);
nor U15743 (N_15743,N_13920,N_14752);
nand U15744 (N_15744,N_14136,N_14701);
or U15745 (N_15745,N_13859,N_14989);
or U15746 (N_15746,N_14930,N_14546);
and U15747 (N_15747,N_14350,N_14460);
nor U15748 (N_15748,N_14580,N_13927);
xnor U15749 (N_15749,N_13869,N_14781);
and U15750 (N_15750,N_14874,N_14441);
and U15751 (N_15751,N_14568,N_13936);
and U15752 (N_15752,N_13761,N_14431);
xor U15753 (N_15753,N_14723,N_14160);
or U15754 (N_15754,N_14064,N_14484);
and U15755 (N_15755,N_14553,N_14709);
nand U15756 (N_15756,N_14691,N_14950);
nand U15757 (N_15757,N_13924,N_14969);
or U15758 (N_15758,N_14486,N_14445);
or U15759 (N_15759,N_14182,N_13832);
and U15760 (N_15760,N_14535,N_14594);
nor U15761 (N_15761,N_14084,N_14923);
nand U15762 (N_15762,N_13991,N_14945);
and U15763 (N_15763,N_13924,N_14547);
nand U15764 (N_15764,N_14809,N_14181);
or U15765 (N_15765,N_14426,N_14840);
nand U15766 (N_15766,N_13940,N_14091);
and U15767 (N_15767,N_14663,N_13750);
nor U15768 (N_15768,N_14825,N_14196);
nand U15769 (N_15769,N_14465,N_13764);
xnor U15770 (N_15770,N_14077,N_13865);
xnor U15771 (N_15771,N_14387,N_14907);
nor U15772 (N_15772,N_14598,N_14651);
nand U15773 (N_15773,N_14914,N_13870);
nor U15774 (N_15774,N_14328,N_14169);
xor U15775 (N_15775,N_14307,N_14811);
nor U15776 (N_15776,N_13964,N_14379);
and U15777 (N_15777,N_14361,N_13984);
nand U15778 (N_15778,N_14469,N_14020);
or U15779 (N_15779,N_14979,N_14043);
xnor U15780 (N_15780,N_13889,N_14404);
nor U15781 (N_15781,N_14841,N_14293);
nand U15782 (N_15782,N_14253,N_14410);
and U15783 (N_15783,N_13895,N_13933);
and U15784 (N_15784,N_14153,N_14871);
xnor U15785 (N_15785,N_14215,N_13927);
xnor U15786 (N_15786,N_14543,N_14217);
nand U15787 (N_15787,N_14007,N_13956);
xnor U15788 (N_15788,N_14862,N_13980);
nor U15789 (N_15789,N_13763,N_14217);
xor U15790 (N_15790,N_14940,N_13816);
and U15791 (N_15791,N_14802,N_13866);
and U15792 (N_15792,N_14097,N_14154);
nor U15793 (N_15793,N_13791,N_14997);
xor U15794 (N_15794,N_14499,N_14490);
nand U15795 (N_15795,N_13925,N_13943);
nor U15796 (N_15796,N_14442,N_13794);
xnor U15797 (N_15797,N_13781,N_14500);
or U15798 (N_15798,N_14272,N_14810);
nor U15799 (N_15799,N_14473,N_14518);
xnor U15800 (N_15800,N_14473,N_14332);
nor U15801 (N_15801,N_14181,N_14646);
nor U15802 (N_15802,N_14040,N_14987);
and U15803 (N_15803,N_13929,N_14836);
and U15804 (N_15804,N_14227,N_13878);
or U15805 (N_15805,N_14121,N_14974);
nand U15806 (N_15806,N_13995,N_14398);
nor U15807 (N_15807,N_14650,N_14115);
or U15808 (N_15808,N_14986,N_14783);
and U15809 (N_15809,N_14116,N_14716);
or U15810 (N_15810,N_13930,N_13982);
xnor U15811 (N_15811,N_14571,N_14842);
and U15812 (N_15812,N_13856,N_13863);
nand U15813 (N_15813,N_14212,N_14982);
and U15814 (N_15814,N_13758,N_14604);
xnor U15815 (N_15815,N_13881,N_13922);
or U15816 (N_15816,N_14396,N_13858);
nand U15817 (N_15817,N_14226,N_13894);
or U15818 (N_15818,N_14596,N_14667);
or U15819 (N_15819,N_14762,N_14451);
xnor U15820 (N_15820,N_14160,N_14010);
and U15821 (N_15821,N_14470,N_14887);
nor U15822 (N_15822,N_14765,N_14779);
nor U15823 (N_15823,N_13861,N_14579);
xor U15824 (N_15824,N_14182,N_14134);
xor U15825 (N_15825,N_14666,N_14632);
and U15826 (N_15826,N_14221,N_14076);
nand U15827 (N_15827,N_14553,N_14305);
or U15828 (N_15828,N_14055,N_14115);
nor U15829 (N_15829,N_14224,N_14181);
or U15830 (N_15830,N_14788,N_14764);
and U15831 (N_15831,N_14543,N_14474);
or U15832 (N_15832,N_14829,N_14510);
and U15833 (N_15833,N_14168,N_13758);
and U15834 (N_15834,N_14809,N_14123);
and U15835 (N_15835,N_14343,N_14570);
xor U15836 (N_15836,N_14834,N_14956);
nor U15837 (N_15837,N_14854,N_13955);
or U15838 (N_15838,N_14398,N_14030);
xnor U15839 (N_15839,N_14044,N_14181);
or U15840 (N_15840,N_14047,N_13824);
and U15841 (N_15841,N_13827,N_14864);
and U15842 (N_15842,N_14764,N_13773);
xnor U15843 (N_15843,N_14202,N_14317);
and U15844 (N_15844,N_14555,N_14089);
or U15845 (N_15845,N_14825,N_13893);
xor U15846 (N_15846,N_14964,N_13883);
nand U15847 (N_15847,N_14875,N_13813);
nand U15848 (N_15848,N_13930,N_14988);
xor U15849 (N_15849,N_14621,N_14972);
and U15850 (N_15850,N_14309,N_14551);
nand U15851 (N_15851,N_14424,N_14576);
nor U15852 (N_15852,N_14586,N_13800);
nor U15853 (N_15853,N_14215,N_13896);
nor U15854 (N_15854,N_14211,N_13805);
or U15855 (N_15855,N_13829,N_14404);
nor U15856 (N_15856,N_14470,N_14048);
and U15857 (N_15857,N_14561,N_13978);
or U15858 (N_15858,N_14994,N_14653);
nand U15859 (N_15859,N_14191,N_14624);
xnor U15860 (N_15860,N_13863,N_14220);
nor U15861 (N_15861,N_14399,N_13832);
or U15862 (N_15862,N_14468,N_14407);
xnor U15863 (N_15863,N_13851,N_14922);
xnor U15864 (N_15864,N_13870,N_14272);
or U15865 (N_15865,N_14880,N_14268);
or U15866 (N_15866,N_13947,N_14837);
nor U15867 (N_15867,N_14399,N_14405);
nand U15868 (N_15868,N_14457,N_14484);
xor U15869 (N_15869,N_14084,N_14097);
and U15870 (N_15870,N_14449,N_14552);
nor U15871 (N_15871,N_14949,N_14501);
nor U15872 (N_15872,N_14059,N_14859);
nor U15873 (N_15873,N_14182,N_14246);
nor U15874 (N_15874,N_14383,N_14142);
and U15875 (N_15875,N_14375,N_14209);
nand U15876 (N_15876,N_13932,N_14617);
xnor U15877 (N_15877,N_14549,N_13852);
and U15878 (N_15878,N_14844,N_14924);
and U15879 (N_15879,N_14424,N_13888);
xor U15880 (N_15880,N_14441,N_14356);
xor U15881 (N_15881,N_14664,N_14969);
or U15882 (N_15882,N_14299,N_14129);
nand U15883 (N_15883,N_14664,N_14385);
nand U15884 (N_15884,N_14826,N_14728);
nor U15885 (N_15885,N_14850,N_14287);
or U15886 (N_15886,N_14466,N_14867);
xor U15887 (N_15887,N_14361,N_14633);
nand U15888 (N_15888,N_14797,N_14320);
or U15889 (N_15889,N_14098,N_13762);
nand U15890 (N_15890,N_14820,N_14753);
or U15891 (N_15891,N_14360,N_13816);
and U15892 (N_15892,N_14765,N_13869);
xnor U15893 (N_15893,N_14368,N_14016);
or U15894 (N_15894,N_13812,N_14697);
or U15895 (N_15895,N_14160,N_14852);
nand U15896 (N_15896,N_14595,N_14269);
or U15897 (N_15897,N_14410,N_14040);
nand U15898 (N_15898,N_14063,N_14340);
and U15899 (N_15899,N_14740,N_14007);
and U15900 (N_15900,N_13908,N_14447);
or U15901 (N_15901,N_14411,N_14539);
nand U15902 (N_15902,N_13854,N_14666);
and U15903 (N_15903,N_13820,N_14118);
and U15904 (N_15904,N_14381,N_14798);
nor U15905 (N_15905,N_14997,N_14796);
and U15906 (N_15906,N_14925,N_14976);
nand U15907 (N_15907,N_14562,N_14568);
and U15908 (N_15908,N_14752,N_14357);
xor U15909 (N_15909,N_13938,N_14036);
nor U15910 (N_15910,N_13998,N_13872);
nor U15911 (N_15911,N_14297,N_14002);
nand U15912 (N_15912,N_14479,N_14270);
xor U15913 (N_15913,N_14643,N_13839);
xor U15914 (N_15914,N_14972,N_14788);
nor U15915 (N_15915,N_14631,N_14596);
or U15916 (N_15916,N_14713,N_14959);
nor U15917 (N_15917,N_14368,N_14745);
and U15918 (N_15918,N_14315,N_14690);
or U15919 (N_15919,N_13820,N_14731);
nand U15920 (N_15920,N_14248,N_13781);
nand U15921 (N_15921,N_14246,N_14795);
xnor U15922 (N_15922,N_14520,N_14691);
xor U15923 (N_15923,N_14497,N_13902);
nor U15924 (N_15924,N_13977,N_14249);
and U15925 (N_15925,N_14108,N_14987);
nand U15926 (N_15926,N_14758,N_14849);
xor U15927 (N_15927,N_13777,N_14938);
and U15928 (N_15928,N_14026,N_14278);
nand U15929 (N_15929,N_14857,N_14883);
xor U15930 (N_15930,N_14766,N_14186);
and U15931 (N_15931,N_14349,N_13778);
nand U15932 (N_15932,N_14309,N_14607);
or U15933 (N_15933,N_14618,N_14307);
nand U15934 (N_15934,N_14331,N_14589);
nor U15935 (N_15935,N_13906,N_14869);
nor U15936 (N_15936,N_13966,N_14630);
and U15937 (N_15937,N_14153,N_13999);
nor U15938 (N_15938,N_14376,N_14036);
or U15939 (N_15939,N_14747,N_14338);
or U15940 (N_15940,N_14522,N_14348);
xnor U15941 (N_15941,N_13864,N_14816);
nand U15942 (N_15942,N_14108,N_14795);
nand U15943 (N_15943,N_14210,N_13861);
nor U15944 (N_15944,N_14654,N_14242);
or U15945 (N_15945,N_14684,N_14272);
nand U15946 (N_15946,N_13881,N_13798);
xnor U15947 (N_15947,N_13946,N_14179);
xor U15948 (N_15948,N_14840,N_14344);
nand U15949 (N_15949,N_14368,N_14141);
nor U15950 (N_15950,N_14603,N_14650);
or U15951 (N_15951,N_14054,N_14489);
or U15952 (N_15952,N_14699,N_14724);
or U15953 (N_15953,N_14432,N_14851);
nand U15954 (N_15954,N_14266,N_14731);
xnor U15955 (N_15955,N_14136,N_14685);
and U15956 (N_15956,N_14150,N_14366);
and U15957 (N_15957,N_14628,N_14356);
or U15958 (N_15958,N_14906,N_14204);
or U15959 (N_15959,N_14434,N_14815);
nor U15960 (N_15960,N_14893,N_14646);
nand U15961 (N_15961,N_14052,N_14963);
and U15962 (N_15962,N_14713,N_14936);
nor U15963 (N_15963,N_14432,N_14345);
nand U15964 (N_15964,N_14252,N_14918);
xor U15965 (N_15965,N_14816,N_13906);
xor U15966 (N_15966,N_13766,N_14702);
or U15967 (N_15967,N_14672,N_14327);
xnor U15968 (N_15968,N_14988,N_14250);
xor U15969 (N_15969,N_14266,N_13775);
xnor U15970 (N_15970,N_14077,N_14131);
xnor U15971 (N_15971,N_14204,N_14017);
or U15972 (N_15972,N_14491,N_14708);
nor U15973 (N_15973,N_14559,N_14276);
nor U15974 (N_15974,N_13939,N_14281);
and U15975 (N_15975,N_14193,N_14798);
nand U15976 (N_15976,N_14023,N_14304);
and U15977 (N_15977,N_14604,N_14515);
xor U15978 (N_15978,N_14576,N_13771);
xnor U15979 (N_15979,N_14914,N_14972);
and U15980 (N_15980,N_14530,N_13862);
nand U15981 (N_15981,N_13923,N_14859);
xor U15982 (N_15982,N_14010,N_14256);
xnor U15983 (N_15983,N_14690,N_13823);
xnor U15984 (N_15984,N_14010,N_14063);
nand U15985 (N_15985,N_14971,N_14444);
and U15986 (N_15986,N_14273,N_14557);
or U15987 (N_15987,N_14851,N_14132);
and U15988 (N_15988,N_14762,N_14729);
xor U15989 (N_15989,N_14732,N_14388);
nand U15990 (N_15990,N_14413,N_14919);
and U15991 (N_15991,N_13930,N_14124);
nand U15992 (N_15992,N_14940,N_13769);
or U15993 (N_15993,N_14396,N_14320);
or U15994 (N_15994,N_14600,N_14407);
nand U15995 (N_15995,N_13834,N_13800);
or U15996 (N_15996,N_14839,N_14859);
or U15997 (N_15997,N_14511,N_13772);
nor U15998 (N_15998,N_14040,N_14403);
and U15999 (N_15999,N_14505,N_14189);
and U16000 (N_16000,N_13856,N_13920);
xor U16001 (N_16001,N_14269,N_13837);
nor U16002 (N_16002,N_14664,N_14887);
xnor U16003 (N_16003,N_14886,N_14128);
nor U16004 (N_16004,N_13880,N_14437);
and U16005 (N_16005,N_13812,N_14778);
and U16006 (N_16006,N_13797,N_14376);
nand U16007 (N_16007,N_14041,N_13833);
or U16008 (N_16008,N_14532,N_14882);
or U16009 (N_16009,N_14352,N_14802);
nor U16010 (N_16010,N_13894,N_13920);
and U16011 (N_16011,N_14592,N_14003);
nand U16012 (N_16012,N_14456,N_14278);
xor U16013 (N_16013,N_14454,N_14599);
nand U16014 (N_16014,N_13988,N_14066);
nor U16015 (N_16015,N_14056,N_13944);
nand U16016 (N_16016,N_14551,N_14083);
or U16017 (N_16017,N_14347,N_14737);
nand U16018 (N_16018,N_14458,N_14452);
nand U16019 (N_16019,N_13877,N_13754);
nor U16020 (N_16020,N_14249,N_14092);
or U16021 (N_16021,N_14216,N_14721);
nand U16022 (N_16022,N_14527,N_14343);
or U16023 (N_16023,N_14267,N_14483);
or U16024 (N_16024,N_14529,N_14526);
xnor U16025 (N_16025,N_14835,N_14999);
nand U16026 (N_16026,N_13962,N_14482);
or U16027 (N_16027,N_14965,N_14497);
and U16028 (N_16028,N_14982,N_14744);
nor U16029 (N_16029,N_14143,N_14987);
and U16030 (N_16030,N_13994,N_14230);
or U16031 (N_16031,N_13968,N_14727);
xor U16032 (N_16032,N_14775,N_14312);
nand U16033 (N_16033,N_14862,N_14079);
nand U16034 (N_16034,N_14094,N_14815);
and U16035 (N_16035,N_14041,N_14563);
and U16036 (N_16036,N_14677,N_14663);
xnor U16037 (N_16037,N_13941,N_14838);
and U16038 (N_16038,N_13935,N_13888);
nand U16039 (N_16039,N_14821,N_14520);
nand U16040 (N_16040,N_14712,N_14647);
xor U16041 (N_16041,N_13828,N_14418);
nor U16042 (N_16042,N_13850,N_13980);
xnor U16043 (N_16043,N_14781,N_14339);
nor U16044 (N_16044,N_14831,N_14304);
and U16045 (N_16045,N_14045,N_14341);
xor U16046 (N_16046,N_14163,N_14986);
nand U16047 (N_16047,N_14787,N_13826);
and U16048 (N_16048,N_14396,N_14699);
or U16049 (N_16049,N_14218,N_13786);
xnor U16050 (N_16050,N_13762,N_14676);
nor U16051 (N_16051,N_14390,N_14986);
nor U16052 (N_16052,N_14411,N_14886);
and U16053 (N_16053,N_14338,N_14535);
nor U16054 (N_16054,N_13817,N_14752);
and U16055 (N_16055,N_14624,N_14934);
and U16056 (N_16056,N_14100,N_14465);
nor U16057 (N_16057,N_13977,N_14981);
and U16058 (N_16058,N_14665,N_14561);
and U16059 (N_16059,N_14513,N_14971);
xor U16060 (N_16060,N_14251,N_14000);
and U16061 (N_16061,N_14294,N_14339);
nand U16062 (N_16062,N_14861,N_14194);
nand U16063 (N_16063,N_14339,N_14349);
nand U16064 (N_16064,N_14565,N_14949);
xor U16065 (N_16065,N_14430,N_14541);
or U16066 (N_16066,N_14600,N_14412);
xnor U16067 (N_16067,N_14641,N_13925);
or U16068 (N_16068,N_14099,N_14827);
or U16069 (N_16069,N_13771,N_14592);
nor U16070 (N_16070,N_14703,N_14969);
nand U16071 (N_16071,N_14623,N_14334);
nand U16072 (N_16072,N_14243,N_14554);
and U16073 (N_16073,N_14056,N_14130);
and U16074 (N_16074,N_13797,N_14166);
nand U16075 (N_16075,N_14264,N_14138);
xor U16076 (N_16076,N_14391,N_14000);
or U16077 (N_16077,N_13821,N_14741);
or U16078 (N_16078,N_14950,N_14334);
nor U16079 (N_16079,N_13918,N_14876);
and U16080 (N_16080,N_13858,N_14449);
and U16081 (N_16081,N_14177,N_14699);
nor U16082 (N_16082,N_13820,N_14282);
nor U16083 (N_16083,N_14555,N_14437);
nor U16084 (N_16084,N_14089,N_14964);
or U16085 (N_16085,N_13997,N_14949);
nor U16086 (N_16086,N_14059,N_14865);
or U16087 (N_16087,N_13962,N_14329);
or U16088 (N_16088,N_14952,N_14224);
nor U16089 (N_16089,N_14601,N_14991);
nand U16090 (N_16090,N_14461,N_14000);
xnor U16091 (N_16091,N_14200,N_14817);
xnor U16092 (N_16092,N_14983,N_14757);
or U16093 (N_16093,N_14927,N_14206);
nor U16094 (N_16094,N_14457,N_14131);
or U16095 (N_16095,N_14940,N_14948);
nor U16096 (N_16096,N_14751,N_13774);
nor U16097 (N_16097,N_14461,N_14353);
and U16098 (N_16098,N_14237,N_14624);
nand U16099 (N_16099,N_14304,N_14966);
nor U16100 (N_16100,N_14855,N_13975);
xnor U16101 (N_16101,N_14057,N_14629);
nand U16102 (N_16102,N_14132,N_14094);
nor U16103 (N_16103,N_13961,N_14090);
or U16104 (N_16104,N_13770,N_13937);
xor U16105 (N_16105,N_14991,N_14589);
xnor U16106 (N_16106,N_14269,N_13756);
and U16107 (N_16107,N_13841,N_14049);
xnor U16108 (N_16108,N_14100,N_14878);
nor U16109 (N_16109,N_14278,N_14609);
xor U16110 (N_16110,N_14668,N_14297);
xor U16111 (N_16111,N_14807,N_14083);
nand U16112 (N_16112,N_14564,N_14978);
xnor U16113 (N_16113,N_14843,N_14104);
or U16114 (N_16114,N_14249,N_14320);
xor U16115 (N_16115,N_14191,N_14271);
nand U16116 (N_16116,N_13752,N_14351);
xor U16117 (N_16117,N_14888,N_13889);
or U16118 (N_16118,N_14102,N_14701);
or U16119 (N_16119,N_14971,N_14053);
and U16120 (N_16120,N_14701,N_14131);
or U16121 (N_16121,N_14353,N_13855);
nor U16122 (N_16122,N_14939,N_14481);
xnor U16123 (N_16123,N_14714,N_14724);
nor U16124 (N_16124,N_14570,N_13976);
or U16125 (N_16125,N_13972,N_13990);
nor U16126 (N_16126,N_14048,N_13960);
or U16127 (N_16127,N_14203,N_14048);
nor U16128 (N_16128,N_13803,N_14404);
or U16129 (N_16129,N_14008,N_14668);
xor U16130 (N_16130,N_14453,N_13855);
nor U16131 (N_16131,N_14217,N_14000);
xnor U16132 (N_16132,N_14217,N_14488);
and U16133 (N_16133,N_14757,N_14937);
or U16134 (N_16134,N_14067,N_13825);
xnor U16135 (N_16135,N_14730,N_14214);
nand U16136 (N_16136,N_13907,N_14101);
or U16137 (N_16137,N_13818,N_14099);
or U16138 (N_16138,N_14752,N_13761);
xor U16139 (N_16139,N_13837,N_14127);
nor U16140 (N_16140,N_14465,N_14045);
nand U16141 (N_16141,N_14487,N_14176);
nand U16142 (N_16142,N_14534,N_13918);
nor U16143 (N_16143,N_14755,N_14220);
or U16144 (N_16144,N_14548,N_14254);
or U16145 (N_16145,N_14394,N_14864);
nor U16146 (N_16146,N_13753,N_14302);
and U16147 (N_16147,N_14659,N_14591);
nor U16148 (N_16148,N_14975,N_14804);
xor U16149 (N_16149,N_14072,N_13870);
nand U16150 (N_16150,N_14859,N_14581);
and U16151 (N_16151,N_14705,N_14924);
nand U16152 (N_16152,N_14297,N_13810);
nand U16153 (N_16153,N_14647,N_14795);
and U16154 (N_16154,N_14206,N_13828);
and U16155 (N_16155,N_14566,N_14964);
nand U16156 (N_16156,N_14464,N_14229);
nor U16157 (N_16157,N_14872,N_13833);
and U16158 (N_16158,N_14709,N_14072);
xor U16159 (N_16159,N_14195,N_13791);
nand U16160 (N_16160,N_14197,N_14227);
xnor U16161 (N_16161,N_14965,N_14078);
xor U16162 (N_16162,N_14403,N_13913);
nor U16163 (N_16163,N_14593,N_14105);
nor U16164 (N_16164,N_13934,N_14495);
and U16165 (N_16165,N_14136,N_13910);
xnor U16166 (N_16166,N_14381,N_14254);
and U16167 (N_16167,N_14608,N_14269);
and U16168 (N_16168,N_13917,N_14223);
or U16169 (N_16169,N_14652,N_13994);
xor U16170 (N_16170,N_14712,N_14164);
nand U16171 (N_16171,N_14425,N_14341);
nand U16172 (N_16172,N_14495,N_14678);
xnor U16173 (N_16173,N_14828,N_14143);
and U16174 (N_16174,N_14983,N_14947);
xnor U16175 (N_16175,N_14891,N_14474);
and U16176 (N_16176,N_14101,N_14182);
xnor U16177 (N_16177,N_14374,N_14097);
xor U16178 (N_16178,N_13768,N_14481);
or U16179 (N_16179,N_14614,N_14638);
nor U16180 (N_16180,N_14879,N_14112);
nor U16181 (N_16181,N_14207,N_13923);
or U16182 (N_16182,N_14132,N_14521);
nand U16183 (N_16183,N_14459,N_14272);
or U16184 (N_16184,N_14497,N_14887);
and U16185 (N_16185,N_13773,N_14226);
xnor U16186 (N_16186,N_14089,N_14005);
nor U16187 (N_16187,N_14871,N_14022);
or U16188 (N_16188,N_14458,N_14727);
or U16189 (N_16189,N_13921,N_14887);
nand U16190 (N_16190,N_14999,N_14002);
nor U16191 (N_16191,N_14922,N_14223);
xnor U16192 (N_16192,N_14119,N_14435);
xor U16193 (N_16193,N_14344,N_14625);
and U16194 (N_16194,N_14264,N_14210);
xor U16195 (N_16195,N_14563,N_14206);
and U16196 (N_16196,N_14335,N_14933);
or U16197 (N_16197,N_14034,N_14720);
or U16198 (N_16198,N_14096,N_14875);
nand U16199 (N_16199,N_14451,N_13859);
and U16200 (N_16200,N_13956,N_13978);
xnor U16201 (N_16201,N_14304,N_14642);
xor U16202 (N_16202,N_14894,N_14414);
nand U16203 (N_16203,N_14168,N_14494);
or U16204 (N_16204,N_13987,N_14221);
or U16205 (N_16205,N_14609,N_14498);
nand U16206 (N_16206,N_14733,N_14483);
nand U16207 (N_16207,N_14391,N_14708);
and U16208 (N_16208,N_13902,N_14653);
and U16209 (N_16209,N_14005,N_13906);
and U16210 (N_16210,N_14575,N_13753);
and U16211 (N_16211,N_14157,N_14591);
nand U16212 (N_16212,N_14482,N_14721);
xor U16213 (N_16213,N_14913,N_14676);
or U16214 (N_16214,N_14907,N_14213);
nor U16215 (N_16215,N_14894,N_14150);
nand U16216 (N_16216,N_14350,N_14845);
nand U16217 (N_16217,N_14573,N_13882);
and U16218 (N_16218,N_14424,N_14324);
nand U16219 (N_16219,N_14350,N_14309);
and U16220 (N_16220,N_14555,N_14619);
xnor U16221 (N_16221,N_13852,N_14056);
xor U16222 (N_16222,N_14499,N_14688);
xor U16223 (N_16223,N_13928,N_13786);
nor U16224 (N_16224,N_14155,N_14224);
xnor U16225 (N_16225,N_14609,N_14374);
nand U16226 (N_16226,N_14182,N_14562);
nor U16227 (N_16227,N_14978,N_14867);
or U16228 (N_16228,N_14736,N_14722);
xor U16229 (N_16229,N_14435,N_14141);
nand U16230 (N_16230,N_14365,N_14323);
nand U16231 (N_16231,N_14213,N_14324);
nand U16232 (N_16232,N_13901,N_13913);
xor U16233 (N_16233,N_14557,N_14807);
nand U16234 (N_16234,N_14314,N_14633);
nor U16235 (N_16235,N_13935,N_14034);
nor U16236 (N_16236,N_14082,N_14747);
nor U16237 (N_16237,N_13961,N_14215);
nor U16238 (N_16238,N_14878,N_13760);
and U16239 (N_16239,N_14156,N_14280);
and U16240 (N_16240,N_14840,N_13857);
or U16241 (N_16241,N_14030,N_14841);
nor U16242 (N_16242,N_14265,N_14917);
and U16243 (N_16243,N_13980,N_14752);
xor U16244 (N_16244,N_14059,N_14209);
or U16245 (N_16245,N_14103,N_14829);
and U16246 (N_16246,N_14350,N_13891);
nor U16247 (N_16247,N_14438,N_14286);
or U16248 (N_16248,N_14895,N_13826);
nor U16249 (N_16249,N_14431,N_13784);
xnor U16250 (N_16250,N_15584,N_15056);
and U16251 (N_16251,N_15358,N_15490);
and U16252 (N_16252,N_16039,N_16216);
xnor U16253 (N_16253,N_15247,N_15261);
nand U16254 (N_16254,N_15688,N_16156);
or U16255 (N_16255,N_15025,N_15124);
and U16256 (N_16256,N_15405,N_15646);
or U16257 (N_16257,N_15648,N_15686);
and U16258 (N_16258,N_16153,N_15181);
and U16259 (N_16259,N_15845,N_16158);
nand U16260 (N_16260,N_15757,N_15432);
nor U16261 (N_16261,N_15211,N_15875);
nor U16262 (N_16262,N_15925,N_15359);
and U16263 (N_16263,N_15240,N_15416);
or U16264 (N_16264,N_15929,N_15833);
and U16265 (N_16265,N_15420,N_15699);
xor U16266 (N_16266,N_15488,N_15203);
and U16267 (N_16267,N_15243,N_15778);
xnor U16268 (N_16268,N_15909,N_15252);
or U16269 (N_16269,N_15012,N_15070);
xor U16270 (N_16270,N_15924,N_15858);
nand U16271 (N_16271,N_15720,N_15919);
xor U16272 (N_16272,N_15384,N_15861);
xor U16273 (N_16273,N_15456,N_15849);
or U16274 (N_16274,N_16249,N_15886);
nand U16275 (N_16275,N_15602,N_15714);
nand U16276 (N_16276,N_15910,N_15156);
nand U16277 (N_16277,N_15661,N_15161);
and U16278 (N_16278,N_15402,N_15524);
xnor U16279 (N_16279,N_15186,N_16217);
xnor U16280 (N_16280,N_15217,N_15689);
and U16281 (N_16281,N_15489,N_16131);
or U16282 (N_16282,N_15447,N_16229);
xor U16283 (N_16283,N_15841,N_15296);
xor U16284 (N_16284,N_15760,N_16182);
and U16285 (N_16285,N_15483,N_15640);
nor U16286 (N_16286,N_15491,N_15262);
xor U16287 (N_16287,N_16148,N_16135);
or U16288 (N_16288,N_15383,N_15257);
nor U16289 (N_16289,N_15703,N_15277);
or U16290 (N_16290,N_15768,N_16165);
and U16291 (N_16291,N_15905,N_15641);
nor U16292 (N_16292,N_15639,N_15556);
xnor U16293 (N_16293,N_16241,N_15476);
nor U16294 (N_16294,N_16002,N_15658);
or U16295 (N_16295,N_15855,N_15902);
nor U16296 (N_16296,N_15835,N_15058);
nand U16297 (N_16297,N_15694,N_16010);
and U16298 (N_16298,N_15246,N_16031);
xnor U16299 (N_16299,N_15749,N_16108);
xor U16300 (N_16300,N_15266,N_15659);
nand U16301 (N_16301,N_15063,N_15995);
xnor U16302 (N_16302,N_15946,N_16093);
xor U16303 (N_16303,N_15064,N_15282);
or U16304 (N_16304,N_15014,N_15285);
nor U16305 (N_16305,N_16020,N_15588);
or U16306 (N_16306,N_15469,N_15040);
nor U16307 (N_16307,N_15140,N_15942);
and U16308 (N_16308,N_15687,N_16151);
nand U16309 (N_16309,N_16197,N_15137);
nand U16310 (N_16310,N_15196,N_15348);
nor U16311 (N_16311,N_15616,N_15985);
nor U16312 (N_16312,N_15957,N_15001);
or U16313 (N_16313,N_15113,N_16027);
or U16314 (N_16314,N_15599,N_15250);
nor U16315 (N_16315,N_15133,N_15604);
xor U16316 (N_16316,N_15430,N_16003);
xnor U16317 (N_16317,N_15182,N_15783);
nor U16318 (N_16318,N_15236,N_15242);
nand U16319 (N_16319,N_15275,N_15174);
nor U16320 (N_16320,N_15042,N_16237);
xor U16321 (N_16321,N_15000,N_15832);
nor U16322 (N_16322,N_16211,N_15429);
nand U16323 (N_16323,N_16170,N_16068);
xnor U16324 (N_16324,N_15756,N_15139);
nor U16325 (N_16325,N_15668,N_15276);
and U16326 (N_16326,N_15700,N_15461);
xnor U16327 (N_16327,N_16188,N_15312);
nor U16328 (N_16328,N_15082,N_15869);
and U16329 (N_16329,N_15517,N_15870);
or U16330 (N_16330,N_15074,N_15656);
and U16331 (N_16331,N_15928,N_15162);
nor U16332 (N_16332,N_15958,N_15825);
and U16333 (N_16333,N_15560,N_15309);
or U16334 (N_16334,N_15854,N_15673);
nor U16335 (N_16335,N_15620,N_16048);
and U16336 (N_16336,N_15607,N_16001);
nand U16337 (N_16337,N_15459,N_15727);
nor U16338 (N_16338,N_15866,N_15787);
nor U16339 (N_16339,N_16240,N_16018);
and U16340 (N_16340,N_15593,N_16190);
and U16341 (N_16341,N_15547,N_15590);
xor U16342 (N_16342,N_16232,N_15600);
nor U16343 (N_16343,N_15479,N_15435);
nand U16344 (N_16344,N_15824,N_15346);
xor U16345 (N_16345,N_15531,N_15759);
nor U16346 (N_16346,N_16198,N_15004);
and U16347 (N_16347,N_15449,N_16009);
nand U16348 (N_16348,N_16126,N_15976);
and U16349 (N_16349,N_15844,N_15422);
xor U16350 (N_16350,N_15138,N_15041);
nor U16351 (N_16351,N_16037,N_15318);
xor U16352 (N_16352,N_15453,N_15375);
nor U16353 (N_16353,N_15219,N_15800);
nand U16354 (N_16354,N_15322,N_15486);
nor U16355 (N_16355,N_16120,N_15540);
nand U16356 (N_16356,N_15685,N_15372);
and U16357 (N_16357,N_16201,N_15998);
and U16358 (N_16358,N_15008,N_15896);
xnor U16359 (N_16359,N_15934,N_15200);
or U16360 (N_16360,N_15290,N_16053);
nor U16361 (N_16361,N_15274,N_15210);
and U16362 (N_16362,N_15736,N_15951);
xnor U16363 (N_16363,N_15884,N_15305);
nand U16364 (N_16364,N_15015,N_15592);
or U16365 (N_16365,N_15024,N_15104);
nand U16366 (N_16366,N_15520,N_15363);
nand U16367 (N_16367,N_15956,N_15894);
nand U16368 (N_16368,N_15766,N_15513);
and U16369 (N_16369,N_15626,N_15379);
nor U16370 (N_16370,N_16043,N_15707);
nand U16371 (N_16371,N_15795,N_15831);
and U16372 (N_16372,N_15650,N_15698);
xnor U16373 (N_16373,N_15895,N_15734);
or U16374 (N_16374,N_15235,N_15681);
nor U16375 (N_16375,N_15974,N_16200);
nand U16376 (N_16376,N_15349,N_15011);
nand U16377 (N_16377,N_15779,N_15049);
nand U16378 (N_16378,N_15750,N_15549);
or U16379 (N_16379,N_15380,N_15514);
nand U16380 (N_16380,N_16087,N_15912);
nor U16381 (N_16381,N_15546,N_15207);
nand U16382 (N_16382,N_15569,N_15791);
nand U16383 (N_16383,N_15804,N_15353);
or U16384 (N_16384,N_15580,N_15053);
or U16385 (N_16385,N_16060,N_15173);
xor U16386 (N_16386,N_15733,N_15330);
or U16387 (N_16387,N_16008,N_15722);
nand U16388 (N_16388,N_16011,N_16086);
or U16389 (N_16389,N_15392,N_15997);
nor U16390 (N_16390,N_15630,N_16052);
or U16391 (N_16391,N_15007,N_15502);
and U16392 (N_16392,N_15117,N_15904);
nand U16393 (N_16393,N_15153,N_15898);
nor U16394 (N_16394,N_15415,N_15529);
xnor U16395 (N_16395,N_15087,N_16074);
nor U16396 (N_16396,N_15829,N_15992);
or U16397 (N_16397,N_16144,N_15037);
and U16398 (N_16398,N_15935,N_15280);
xor U16399 (N_16399,N_15079,N_15744);
and U16400 (N_16400,N_15785,N_15177);
nor U16401 (N_16401,N_15081,N_16112);
and U16402 (N_16402,N_15554,N_15206);
nor U16403 (N_16403,N_15442,N_15194);
nand U16404 (N_16404,N_15899,N_15819);
xnor U16405 (N_16405,N_15273,N_15860);
xor U16406 (N_16406,N_15188,N_15678);
or U16407 (N_16407,N_15792,N_16004);
xor U16408 (N_16408,N_15164,N_15059);
or U16409 (N_16409,N_16171,N_15323);
nand U16410 (N_16410,N_15692,N_15971);
or U16411 (N_16411,N_15765,N_15562);
and U16412 (N_16412,N_15631,N_15506);
nand U16413 (N_16413,N_15767,N_15370);
xnor U16414 (N_16414,N_15334,N_15959);
and U16415 (N_16415,N_15283,N_15227);
xnor U16416 (N_16416,N_16129,N_15538);
or U16417 (N_16417,N_15615,N_15916);
and U16418 (N_16418,N_15999,N_15726);
and U16419 (N_16419,N_15216,N_15851);
nor U16420 (N_16420,N_15477,N_15255);
nor U16421 (N_16421,N_15613,N_15594);
nand U16422 (N_16422,N_15980,N_15473);
xnor U16423 (N_16423,N_15048,N_16017);
or U16424 (N_16424,N_15103,N_15047);
and U16425 (N_16425,N_15019,N_16032);
and U16426 (N_16426,N_15657,N_16176);
nand U16427 (N_16427,N_15545,N_15126);
and U16428 (N_16428,N_15633,N_15728);
nor U16429 (N_16429,N_15180,N_15862);
and U16430 (N_16430,N_16036,N_15316);
and U16431 (N_16431,N_16161,N_15628);
nand U16432 (N_16432,N_15150,N_16209);
and U16433 (N_16433,N_15611,N_15598);
or U16434 (N_16434,N_15705,N_15339);
and U16435 (N_16435,N_15143,N_15035);
or U16436 (N_16436,N_15263,N_15706);
nand U16437 (N_16437,N_15654,N_15184);
xor U16438 (N_16438,N_15121,N_15239);
xor U16439 (N_16439,N_15676,N_15621);
or U16440 (N_16440,N_16231,N_15932);
and U16441 (N_16441,N_15347,N_15664);
or U16442 (N_16442,N_15146,N_16166);
nor U16443 (N_16443,N_15834,N_15101);
or U16444 (N_16444,N_15399,N_15943);
and U16445 (N_16445,N_15608,N_15256);
nand U16446 (N_16446,N_15625,N_15494);
xor U16447 (N_16447,N_15328,N_15403);
nor U16448 (N_16448,N_15267,N_15417);
and U16449 (N_16449,N_15578,N_16234);
nor U16450 (N_16450,N_15268,N_15947);
nor U16451 (N_16451,N_15762,N_16105);
and U16452 (N_16452,N_15637,N_15474);
or U16453 (N_16453,N_15465,N_15357);
and U16454 (N_16454,N_15542,N_15470);
nand U16455 (N_16455,N_16245,N_15623);
nor U16456 (N_16456,N_15409,N_16083);
nor U16457 (N_16457,N_15222,N_16085);
and U16458 (N_16458,N_15536,N_15135);
nor U16459 (N_16459,N_16092,N_15108);
xnor U16460 (N_16460,N_15497,N_16062);
and U16461 (N_16461,N_16212,N_15033);
or U16462 (N_16462,N_15893,N_15237);
or U16463 (N_16463,N_15890,N_15311);
nand U16464 (N_16464,N_16168,N_15045);
nor U16465 (N_16465,N_16244,N_15903);
nor U16466 (N_16466,N_15002,N_15292);
and U16467 (N_16467,N_15709,N_16167);
xor U16468 (N_16468,N_16186,N_15125);
nor U16469 (N_16469,N_16067,N_15365);
xnor U16470 (N_16470,N_15345,N_15565);
xor U16471 (N_16471,N_15682,N_15986);
or U16472 (N_16472,N_15333,N_15404);
nand U16473 (N_16473,N_15746,N_15589);
and U16474 (N_16474,N_15710,N_15026);
xnor U16475 (N_16475,N_15291,N_15289);
nor U16476 (N_16476,N_15675,N_15923);
xor U16477 (N_16477,N_16119,N_16169);
nor U16478 (N_16478,N_16081,N_15526);
xnor U16479 (N_16479,N_16050,N_15208);
xnor U16480 (N_16480,N_15737,N_15649);
nor U16481 (N_16481,N_16128,N_15134);
and U16482 (N_16482,N_15109,N_15360);
xor U16483 (N_16483,N_15114,N_15798);
or U16484 (N_16484,N_15663,N_15455);
xor U16485 (N_16485,N_15391,N_15444);
or U16486 (N_16486,N_15102,N_15577);
nor U16487 (N_16487,N_16118,N_16044);
or U16488 (N_16488,N_15350,N_15094);
nand U16489 (N_16489,N_15982,N_15010);
xor U16490 (N_16490,N_15900,N_15475);
xnor U16491 (N_16491,N_15201,N_15367);
or U16492 (N_16492,N_15293,N_15670);
and U16493 (N_16493,N_15773,N_15234);
nor U16494 (N_16494,N_15300,N_15907);
xor U16495 (N_16495,N_16015,N_15828);
or U16496 (N_16496,N_15583,N_15511);
nand U16497 (N_16497,N_15882,N_15695);
nor U16498 (N_16498,N_15128,N_15572);
xnor U16499 (N_16499,N_15189,N_16012);
nor U16500 (N_16500,N_16065,N_15771);
nor U16501 (N_16501,N_16103,N_15813);
and U16502 (N_16502,N_16090,N_15541);
nor U16503 (N_16503,N_15098,N_16046);
nor U16504 (N_16504,N_15665,N_15763);
nor U16505 (N_16505,N_16045,N_15721);
or U16506 (N_16506,N_15374,N_15448);
nor U16507 (N_16507,N_15232,N_15642);
or U16508 (N_16508,N_16056,N_15610);
nor U16509 (N_16509,N_15095,N_15651);
or U16510 (N_16510,N_15467,N_16159);
nor U16511 (N_16511,N_15776,N_15669);
or U16512 (N_16512,N_15810,N_15249);
and U16513 (N_16513,N_15454,N_15185);
xor U16514 (N_16514,N_15426,N_15226);
xor U16515 (N_16515,N_15635,N_15732);
nand U16516 (N_16516,N_16130,N_15826);
nand U16517 (N_16517,N_15761,N_16084);
and U16518 (N_16518,N_16183,N_16236);
nand U16519 (N_16519,N_15803,N_16248);
nor U16520 (N_16520,N_16088,N_16069);
xor U16521 (N_16521,N_15075,N_15815);
nand U16522 (N_16522,N_15843,N_16204);
nor U16523 (N_16523,N_15319,N_15752);
xor U16524 (N_16524,N_15362,N_15119);
nor U16525 (N_16525,N_16145,N_15597);
and U16526 (N_16526,N_15144,N_15751);
nor U16527 (N_16527,N_15696,N_15122);
nand U16528 (N_16528,N_15505,N_15050);
and U16529 (N_16529,N_15166,N_15865);
xor U16530 (N_16530,N_16006,N_15361);
or U16531 (N_16531,N_15425,N_15571);
or U16532 (N_16532,N_15179,N_15788);
and U16533 (N_16533,N_15191,N_15410);
xor U16534 (N_16534,N_15299,N_15717);
or U16535 (N_16535,N_15738,N_15557);
nor U16536 (N_16536,N_15655,N_15215);
xor U16537 (N_16537,N_16189,N_15155);
and U16538 (N_16538,N_15881,N_15495);
xnor U16539 (N_16539,N_15500,N_15984);
nand U16540 (N_16540,N_16016,N_16177);
nand U16541 (N_16541,N_15424,N_15199);
and U16542 (N_16542,N_15463,N_16040);
xor U16543 (N_16543,N_15614,N_15585);
nor U16544 (N_16544,N_15922,N_15627);
and U16545 (N_16545,N_15820,N_15743);
or U16546 (N_16546,N_15065,N_16138);
nand U16547 (N_16547,N_15874,N_15013);
and U16548 (N_16548,N_15034,N_15945);
nand U16549 (N_16549,N_16114,N_15739);
nor U16550 (N_16550,N_15794,N_15619);
nor U16551 (N_16551,N_16226,N_15989);
or U16552 (N_16552,N_15559,N_15202);
nand U16553 (N_16553,N_15725,N_15754);
nand U16554 (N_16554,N_15428,N_15084);
xor U16555 (N_16555,N_16137,N_15386);
nor U16556 (N_16556,N_15777,N_15018);
and U16557 (N_16557,N_15111,N_16149);
nand U16558 (N_16558,N_15458,N_16123);
and U16559 (N_16559,N_15068,N_15638);
and U16560 (N_16560,N_15933,N_15438);
nor U16561 (N_16561,N_16025,N_15052);
xor U16562 (N_16562,N_15576,N_16164);
nand U16563 (N_16563,N_16213,N_15853);
xnor U16564 (N_16564,N_15634,N_15419);
xnor U16565 (N_16565,N_15937,N_16133);
nor U16566 (N_16566,N_15806,N_16094);
or U16567 (N_16567,N_15774,N_15931);
nand U16568 (N_16568,N_16054,N_16098);
nor U16569 (N_16569,N_15431,N_15006);
nor U16570 (N_16570,N_15662,N_16035);
and U16571 (N_16571,N_16192,N_15786);
or U16572 (N_16572,N_15660,N_15214);
xnor U16573 (N_16573,N_15272,N_15555);
and U16574 (N_16574,N_15814,N_15209);
xnor U16575 (N_16575,N_15867,N_15512);
nor U16576 (N_16576,N_15534,N_15413);
xnor U16577 (N_16577,N_15969,N_16091);
xor U16578 (N_16578,N_15537,N_15434);
and U16579 (N_16579,N_15645,N_16063);
nand U16580 (N_16580,N_15452,N_16173);
nand U16581 (N_16581,N_15622,N_15516);
xor U16582 (N_16582,N_15652,N_15248);
or U16583 (N_16583,N_15667,N_15677);
and U16584 (N_16584,N_15582,N_15238);
xor U16585 (N_16585,N_15069,N_15187);
nand U16586 (N_16586,N_15618,N_15755);
xor U16587 (N_16587,N_15741,N_16076);
and U16588 (N_16588,N_15802,N_15371);
and U16589 (N_16589,N_15229,N_15601);
and U16590 (N_16590,N_15204,N_15397);
nor U16591 (N_16591,N_15351,N_15228);
or U16592 (N_16592,N_15801,N_16034);
xnor U16593 (N_16593,N_15337,N_15878);
and U16594 (N_16594,N_15535,N_15325);
and U16595 (N_16595,N_15758,N_15724);
xor U16596 (N_16596,N_15287,N_15848);
xor U16597 (N_16597,N_15088,N_15901);
or U16598 (N_16598,N_16078,N_15480);
and U16599 (N_16599,N_15457,N_15072);
and U16600 (N_16600,N_15073,N_15770);
nor U16601 (N_16601,N_15106,N_16013);
or U16602 (N_16602,N_16042,N_15307);
nor U16603 (N_16603,N_15190,N_15983);
nand U16604 (N_16604,N_15857,N_15340);
or U16605 (N_16605,N_15877,N_15550);
or U16606 (N_16606,N_15057,N_15693);
nor U16607 (N_16607,N_15965,N_15519);
and U16608 (N_16608,N_15515,N_16223);
and U16609 (N_16609,N_15286,N_15115);
xnor U16610 (N_16610,N_16141,N_16073);
and U16611 (N_16611,N_15224,N_15889);
xnor U16612 (N_16612,N_16194,N_15281);
xor U16613 (N_16613,N_16233,N_15341);
xnor U16614 (N_16614,N_15451,N_15054);
xor U16615 (N_16615,N_15532,N_15259);
or U16616 (N_16616,N_15716,N_15501);
or U16617 (N_16617,N_16005,N_15149);
or U16618 (N_16618,N_15988,N_15888);
and U16619 (N_16619,N_15836,N_15544);
nor U16620 (N_16620,N_16242,N_15930);
and U16621 (N_16621,N_15690,N_15464);
nand U16622 (N_16622,N_15543,N_15394);
nand U16623 (N_16623,N_15918,N_15715);
nor U16624 (N_16624,N_16109,N_15342);
xnor U16625 (N_16625,N_15807,N_15492);
nand U16626 (N_16626,N_15440,N_15671);
nand U16627 (N_16627,N_15023,N_15533);
nand U16628 (N_16628,N_15955,N_15443);
nand U16629 (N_16629,N_15172,N_15271);
nor U16630 (N_16630,N_15913,N_15433);
or U16631 (N_16631,N_15132,N_15478);
nor U16632 (N_16632,N_15218,N_16079);
or U16633 (N_16633,N_15089,N_15927);
and U16634 (N_16634,N_15643,N_15817);
nor U16635 (N_16635,N_16154,N_15326);
or U16636 (N_16636,N_15376,N_15784);
nor U16637 (N_16637,N_15044,N_15387);
and U16638 (N_16638,N_16122,N_15418);
and U16639 (N_16639,N_15027,N_15987);
nor U16640 (N_16640,N_15329,N_15003);
xor U16641 (N_16641,N_15879,N_16041);
and U16642 (N_16642,N_15936,N_15868);
nand U16643 (N_16643,N_16066,N_15278);
or U16644 (N_16644,N_15016,N_15586);
and U16645 (N_16645,N_15644,N_15436);
nand U16646 (N_16646,N_15568,N_16205);
nor U16647 (N_16647,N_15223,N_15366);
nor U16648 (N_16648,N_15527,N_16101);
nand U16649 (N_16649,N_15887,N_16104);
and U16650 (N_16650,N_15521,N_15412);
nand U16651 (N_16651,N_15175,N_15028);
or U16652 (N_16652,N_15968,N_15863);
or U16653 (N_16653,N_16082,N_15609);
xor U16654 (N_16654,N_15244,N_15498);
nand U16655 (N_16655,N_15051,N_15827);
xor U16656 (N_16656,N_15225,N_15279);
xnor U16657 (N_16657,N_15395,N_15183);
and U16658 (N_16658,N_16247,N_15704);
nand U16659 (N_16659,N_16191,N_15624);
xnor U16660 (N_16660,N_16111,N_15352);
nor U16661 (N_16661,N_15388,N_15892);
xnor U16662 (N_16662,N_15852,N_15310);
and U16663 (N_16663,N_15398,N_15169);
nand U16664 (N_16664,N_15876,N_16181);
or U16665 (N_16665,N_15120,N_15730);
or U16666 (N_16666,N_16070,N_15039);
or U16667 (N_16667,N_15636,N_15508);
or U16668 (N_16668,N_15295,N_15096);
nand U16669 (N_16669,N_15270,N_15195);
and U16670 (N_16670,N_15205,N_15136);
nor U16671 (N_16671,N_15030,N_16215);
nand U16672 (N_16672,N_15294,N_15575);
or U16673 (N_16673,N_15996,N_15908);
and U16674 (N_16674,N_16038,N_15332);
nand U16675 (N_16675,N_15493,N_15067);
nand U16676 (N_16676,N_16208,N_15548);
xnor U16677 (N_16677,N_15812,N_15712);
nand U16678 (N_16678,N_15321,N_15790);
and U16679 (N_16679,N_16140,N_15085);
or U16680 (N_16680,N_15157,N_15029);
nand U16681 (N_16681,N_15612,N_15129);
and U16682 (N_16682,N_15579,N_15967);
xnor U16683 (N_16683,N_15158,N_15847);
xnor U16684 (N_16684,N_16220,N_16214);
or U16685 (N_16685,N_15856,N_15245);
or U16686 (N_16686,N_15864,N_15260);
xor U16687 (N_16687,N_15303,N_15629);
nor U16688 (N_16688,N_15837,N_16230);
nor U16689 (N_16689,N_16146,N_16100);
and U16690 (N_16690,N_15423,N_15883);
and U16691 (N_16691,N_16089,N_15154);
xnor U16692 (N_16692,N_15100,N_16024);
xnor U16693 (N_16693,N_15163,N_15466);
nand U16694 (N_16694,N_15396,N_15308);
nand U16695 (N_16695,N_15414,N_15141);
xor U16696 (N_16696,N_16160,N_15369);
nor U16697 (N_16697,N_16000,N_15816);
xor U16698 (N_16698,N_16175,N_16157);
or U16699 (N_16699,N_16219,N_15167);
xnor U16700 (N_16700,N_15911,N_16218);
nand U16701 (N_16701,N_15960,N_15719);
or U16702 (N_16702,N_16075,N_15343);
and U16703 (N_16703,N_16180,N_15566);
and U16704 (N_16704,N_15605,N_15977);
nand U16705 (N_16705,N_15302,N_15897);
and U16706 (N_16706,N_15344,N_15269);
xor U16707 (N_16707,N_15021,N_15702);
and U16708 (N_16708,N_15481,N_15797);
nor U16709 (N_16709,N_15439,N_15253);
and U16710 (N_16710,N_15994,N_15830);
nand U16711 (N_16711,N_15966,N_15921);
and U16712 (N_16712,N_15504,N_15406);
xor U16713 (N_16713,N_15723,N_15471);
xor U16714 (N_16714,N_16014,N_15389);
and U16715 (N_16715,N_15306,N_15324);
or U16716 (N_16716,N_15680,N_15020);
nor U16717 (N_16717,N_16195,N_15530);
xnor U16718 (N_16718,N_16102,N_16150);
or U16719 (N_16719,N_15840,N_16225);
xor U16720 (N_16720,N_15729,N_16022);
xor U16721 (N_16721,N_15407,N_15080);
nand U16722 (N_16722,N_15327,N_16127);
and U16723 (N_16723,N_16033,N_15846);
and U16724 (N_16724,N_15711,N_15595);
or U16725 (N_16725,N_15811,N_15975);
nand U16726 (N_16726,N_16064,N_15684);
nand U16727 (N_16727,N_16071,N_15221);
and U16728 (N_16728,N_16227,N_15948);
and U16729 (N_16729,N_15872,N_15666);
nand U16730 (N_16730,N_15031,N_15781);
or U16731 (N_16731,N_15220,N_16026);
or U16732 (N_16732,N_15441,N_15091);
or U16733 (N_16733,N_15304,N_15450);
or U16734 (N_16734,N_16095,N_15796);
nor U16735 (N_16735,N_15775,N_15873);
and U16736 (N_16736,N_16143,N_15920);
nand U16737 (N_16737,N_15265,N_15198);
xnor U16738 (N_16738,N_15617,N_15382);
or U16739 (N_16739,N_15926,N_16049);
xnor U16740 (N_16740,N_15046,N_15178);
nor U16741 (N_16741,N_15891,N_15558);
or U16742 (N_16742,N_15510,N_15487);
xnor U16743 (N_16743,N_15077,N_15944);
xnor U16744 (N_16744,N_16021,N_15385);
or U16745 (N_16745,N_15764,N_15954);
and U16746 (N_16746,N_16179,N_16099);
nand U16747 (N_16747,N_15780,N_15991);
xor U16748 (N_16748,N_15468,N_15962);
and U16749 (N_16749,N_15148,N_15197);
xor U16750 (N_16750,N_15496,N_15674);
xnor U16751 (N_16751,N_15401,N_15708);
nand U16752 (N_16752,N_15672,N_15147);
or U16753 (N_16753,N_15950,N_15381);
xor U16754 (N_16754,N_15145,N_15142);
nor U16755 (N_16755,N_16019,N_15799);
nor U16756 (N_16756,N_15338,N_15408);
nand U16757 (N_16757,N_16059,N_15906);
or U16758 (N_16758,N_16136,N_15264);
xor U16759 (N_16759,N_16239,N_15939);
nor U16760 (N_16760,N_15009,N_16061);
or U16761 (N_16761,N_15446,N_15254);
and U16762 (N_16762,N_15171,N_15885);
and U16763 (N_16763,N_16080,N_15964);
nor U16764 (N_16764,N_15563,N_15850);
and U16765 (N_16765,N_16055,N_15503);
nand U16766 (N_16766,N_15314,N_15573);
or U16767 (N_16767,N_15963,N_16125);
or U16768 (N_16768,N_15038,N_16238);
and U16769 (N_16769,N_15427,N_15822);
and U16770 (N_16770,N_15606,N_16246);
nor U16771 (N_16771,N_15523,N_15509);
or U16772 (N_16772,N_16117,N_15152);
xor U16773 (N_16773,N_15097,N_15301);
or U16774 (N_16774,N_15697,N_16072);
xor U16775 (N_16775,N_15335,N_15043);
nor U16776 (N_16776,N_15683,N_15355);
nand U16777 (N_16777,N_15017,N_15151);
nor U16778 (N_16778,N_15821,N_15123);
nor U16779 (N_16779,N_15701,N_15978);
and U16780 (N_16780,N_15528,N_16221);
and U16781 (N_16781,N_15679,N_16047);
or U16782 (N_16782,N_16210,N_15336);
nor U16783 (N_16783,N_16184,N_15567);
nor U16784 (N_16784,N_15789,N_15160);
nand U16785 (N_16785,N_15742,N_16106);
xor U16786 (N_16786,N_16124,N_15485);
xnor U16787 (N_16787,N_15284,N_15317);
nand U16788 (N_16788,N_15460,N_15231);
nor U16789 (N_16789,N_15241,N_15740);
and U16790 (N_16790,N_16228,N_15165);
or U16791 (N_16791,N_15005,N_15981);
xor U16792 (N_16792,N_15632,N_16132);
xor U16793 (N_16793,N_15809,N_15076);
xor U16794 (N_16794,N_16113,N_16163);
and U16795 (N_16795,N_15356,N_15062);
xnor U16796 (N_16796,N_15105,N_16121);
nor U16797 (N_16797,N_16235,N_15518);
and U16798 (N_16798,N_15110,N_15061);
or U16799 (N_16799,N_15390,N_15230);
nor U16800 (N_16800,N_15564,N_16178);
nor U16801 (N_16801,N_15731,N_16110);
xor U16802 (N_16802,N_15083,N_16162);
or U16803 (N_16803,N_16207,N_15251);
and U16804 (N_16804,N_15525,N_15078);
nor U16805 (N_16805,N_16058,N_16206);
xor U16806 (N_16806,N_15647,N_15574);
or U16807 (N_16807,N_16023,N_15596);
or U16808 (N_16808,N_15331,N_16155);
and U16809 (N_16809,N_15745,N_15972);
xnor U16810 (N_16810,N_16116,N_15482);
nor U16811 (N_16811,N_15297,N_15823);
nand U16812 (N_16812,N_16142,N_15990);
nor U16813 (N_16813,N_15373,N_16222);
or U16814 (N_16814,N_15805,N_16202);
nand U16815 (N_16815,N_16172,N_15112);
xor U16816 (N_16816,N_15093,N_16147);
nand U16817 (N_16817,N_15938,N_15354);
nand U16818 (N_16818,N_15377,N_15170);
or U16819 (N_16819,N_16174,N_15772);
nor U16820 (N_16820,N_16097,N_15192);
xnor U16821 (N_16821,N_15949,N_15769);
or U16822 (N_16822,N_15871,N_15973);
nand U16823 (N_16823,N_15066,N_15168);
and U16824 (N_16824,N_15472,N_15116);
and U16825 (N_16825,N_15484,N_15298);
nand U16826 (N_16826,N_15591,N_15970);
or U16827 (N_16827,N_15288,N_15941);
nor U16828 (N_16828,N_15979,N_16193);
or U16829 (N_16829,N_15859,N_15735);
nand U16830 (N_16830,N_15099,N_16203);
nand U16831 (N_16831,N_16187,N_16007);
xnor U16832 (N_16832,N_16077,N_15917);
and U16833 (N_16833,N_15320,N_15060);
and U16834 (N_16834,N_15176,N_16139);
nand U16835 (N_16835,N_15808,N_15842);
and U16836 (N_16836,N_15499,N_16029);
or U16837 (N_16837,N_15130,N_15092);
xor U16838 (N_16838,N_16185,N_15553);
or U16839 (N_16839,N_15961,N_15071);
nor U16840 (N_16840,N_15090,N_16107);
or U16841 (N_16841,N_15552,N_15313);
or U16842 (N_16842,N_15818,N_15411);
xor U16843 (N_16843,N_15570,N_15213);
xnor U16844 (N_16844,N_16028,N_15364);
nand U16845 (N_16845,N_15587,N_15718);
xor U16846 (N_16846,N_15539,N_15748);
nor U16847 (N_16847,N_15393,N_15233);
nand U16848 (N_16848,N_16243,N_15159);
nand U16849 (N_16849,N_15782,N_16096);
nand U16850 (N_16850,N_15212,N_15691);
or U16851 (N_16851,N_15445,N_15378);
xnor U16852 (N_16852,N_15653,N_15118);
and U16853 (N_16853,N_15522,N_15953);
xor U16854 (N_16854,N_16224,N_15315);
nand U16855 (N_16855,N_15107,N_15581);
and U16856 (N_16856,N_16030,N_15993);
nor U16857 (N_16857,N_15368,N_16196);
nand U16858 (N_16858,N_15915,N_15839);
nor U16859 (N_16859,N_15747,N_16051);
xor U16860 (N_16860,N_15713,N_15603);
nor U16861 (N_16861,N_15131,N_15952);
nor U16862 (N_16862,N_15880,N_15551);
nor U16863 (N_16863,N_16057,N_15753);
xnor U16864 (N_16864,N_15258,N_15036);
nor U16865 (N_16865,N_15462,N_15400);
or U16866 (N_16866,N_15561,N_15022);
nor U16867 (N_16867,N_15055,N_15086);
xor U16868 (N_16868,N_15914,N_15793);
and U16869 (N_16869,N_15940,N_15507);
and U16870 (N_16870,N_15193,N_16115);
or U16871 (N_16871,N_15838,N_15437);
nor U16872 (N_16872,N_16152,N_16134);
and U16873 (N_16873,N_16199,N_15421);
nand U16874 (N_16874,N_15032,N_15127);
or U16875 (N_16875,N_15905,N_16169);
xnor U16876 (N_16876,N_15519,N_16240);
nand U16877 (N_16877,N_16123,N_15800);
and U16878 (N_16878,N_15363,N_15142);
xor U16879 (N_16879,N_15403,N_15623);
or U16880 (N_16880,N_15235,N_15355);
nor U16881 (N_16881,N_15000,N_15581);
or U16882 (N_16882,N_15654,N_15987);
xnor U16883 (N_16883,N_15876,N_15516);
nand U16884 (N_16884,N_16027,N_15083);
or U16885 (N_16885,N_15738,N_16069);
or U16886 (N_16886,N_15208,N_15488);
or U16887 (N_16887,N_15753,N_15165);
xor U16888 (N_16888,N_16239,N_15238);
nand U16889 (N_16889,N_15437,N_15555);
nand U16890 (N_16890,N_16109,N_15724);
xnor U16891 (N_16891,N_16124,N_15609);
nor U16892 (N_16892,N_15276,N_15870);
and U16893 (N_16893,N_15810,N_15503);
nand U16894 (N_16894,N_15112,N_15161);
xor U16895 (N_16895,N_16085,N_15656);
nor U16896 (N_16896,N_15396,N_16134);
and U16897 (N_16897,N_15644,N_15092);
nand U16898 (N_16898,N_15723,N_15470);
nor U16899 (N_16899,N_15504,N_15814);
nor U16900 (N_16900,N_15938,N_15525);
or U16901 (N_16901,N_15462,N_15023);
xor U16902 (N_16902,N_15465,N_15591);
and U16903 (N_16903,N_15456,N_15968);
xor U16904 (N_16904,N_15454,N_15432);
xnor U16905 (N_16905,N_15661,N_15293);
xor U16906 (N_16906,N_15184,N_15115);
nand U16907 (N_16907,N_15122,N_15960);
and U16908 (N_16908,N_15249,N_15133);
nand U16909 (N_16909,N_15388,N_15781);
and U16910 (N_16910,N_15615,N_15763);
nor U16911 (N_16911,N_15300,N_15717);
nand U16912 (N_16912,N_15306,N_15269);
nand U16913 (N_16913,N_15560,N_15335);
nand U16914 (N_16914,N_16000,N_15524);
and U16915 (N_16915,N_15259,N_16089);
and U16916 (N_16916,N_15164,N_15812);
nand U16917 (N_16917,N_15552,N_15214);
xor U16918 (N_16918,N_16126,N_15521);
nand U16919 (N_16919,N_15057,N_15511);
xor U16920 (N_16920,N_16101,N_15170);
and U16921 (N_16921,N_15325,N_15301);
nand U16922 (N_16922,N_15398,N_16070);
nor U16923 (N_16923,N_16151,N_15036);
or U16924 (N_16924,N_15039,N_15479);
or U16925 (N_16925,N_15120,N_15741);
nand U16926 (N_16926,N_15721,N_15803);
nor U16927 (N_16927,N_15310,N_15276);
xor U16928 (N_16928,N_16187,N_15221);
xor U16929 (N_16929,N_15713,N_15353);
or U16930 (N_16930,N_15958,N_15761);
or U16931 (N_16931,N_15545,N_15981);
nand U16932 (N_16932,N_15641,N_15752);
or U16933 (N_16933,N_15599,N_15556);
nand U16934 (N_16934,N_16036,N_15122);
and U16935 (N_16935,N_15001,N_15649);
or U16936 (N_16936,N_15661,N_15278);
nor U16937 (N_16937,N_15426,N_15294);
and U16938 (N_16938,N_15284,N_15064);
or U16939 (N_16939,N_15864,N_16065);
nor U16940 (N_16940,N_15877,N_15854);
or U16941 (N_16941,N_15760,N_15631);
or U16942 (N_16942,N_15605,N_15639);
nand U16943 (N_16943,N_15916,N_15725);
or U16944 (N_16944,N_15386,N_15296);
nor U16945 (N_16945,N_15564,N_15485);
xnor U16946 (N_16946,N_15444,N_15712);
or U16947 (N_16947,N_15632,N_15020);
and U16948 (N_16948,N_15468,N_15945);
nand U16949 (N_16949,N_15992,N_15588);
or U16950 (N_16950,N_15131,N_16125);
or U16951 (N_16951,N_15844,N_16112);
and U16952 (N_16952,N_15112,N_15197);
nand U16953 (N_16953,N_15158,N_15670);
or U16954 (N_16954,N_15300,N_16241);
or U16955 (N_16955,N_15853,N_15067);
nor U16956 (N_16956,N_16082,N_15336);
or U16957 (N_16957,N_15885,N_16230);
xnor U16958 (N_16958,N_15560,N_16063);
or U16959 (N_16959,N_15903,N_15382);
and U16960 (N_16960,N_16050,N_15119);
nand U16961 (N_16961,N_16064,N_15222);
xor U16962 (N_16962,N_15821,N_15135);
nand U16963 (N_16963,N_16048,N_15512);
nor U16964 (N_16964,N_15803,N_15771);
nand U16965 (N_16965,N_15909,N_15349);
nor U16966 (N_16966,N_15020,N_15213);
nor U16967 (N_16967,N_15282,N_15673);
and U16968 (N_16968,N_16178,N_15651);
xor U16969 (N_16969,N_15761,N_15396);
nand U16970 (N_16970,N_15927,N_15926);
nand U16971 (N_16971,N_15929,N_15245);
or U16972 (N_16972,N_16202,N_16072);
xnor U16973 (N_16973,N_15414,N_16220);
and U16974 (N_16974,N_15053,N_15541);
nand U16975 (N_16975,N_15357,N_15270);
nand U16976 (N_16976,N_15384,N_15229);
xor U16977 (N_16977,N_16098,N_15132);
nand U16978 (N_16978,N_15456,N_15624);
xor U16979 (N_16979,N_15310,N_15617);
xor U16980 (N_16980,N_15298,N_15817);
or U16981 (N_16981,N_15453,N_16189);
nor U16982 (N_16982,N_15754,N_15566);
xnor U16983 (N_16983,N_15275,N_15212);
xnor U16984 (N_16984,N_16229,N_15099);
xnor U16985 (N_16985,N_15352,N_15842);
nor U16986 (N_16986,N_16204,N_15515);
or U16987 (N_16987,N_16226,N_16090);
xor U16988 (N_16988,N_15180,N_15365);
and U16989 (N_16989,N_15676,N_15861);
and U16990 (N_16990,N_15735,N_15179);
nor U16991 (N_16991,N_15198,N_15904);
nand U16992 (N_16992,N_15785,N_15864);
xnor U16993 (N_16993,N_15130,N_15838);
xnor U16994 (N_16994,N_16215,N_15005);
nor U16995 (N_16995,N_15360,N_15924);
or U16996 (N_16996,N_16001,N_15268);
nor U16997 (N_16997,N_15645,N_15506);
nor U16998 (N_16998,N_15178,N_15926);
or U16999 (N_16999,N_15660,N_15794);
xnor U17000 (N_17000,N_16032,N_16022);
xor U17001 (N_17001,N_15246,N_15159);
nor U17002 (N_17002,N_15999,N_15822);
xor U17003 (N_17003,N_15959,N_15851);
xor U17004 (N_17004,N_16137,N_15376);
nand U17005 (N_17005,N_15012,N_15267);
nor U17006 (N_17006,N_15704,N_16003);
or U17007 (N_17007,N_15972,N_15548);
nor U17008 (N_17008,N_15878,N_16105);
xnor U17009 (N_17009,N_15494,N_15956);
and U17010 (N_17010,N_15077,N_15254);
or U17011 (N_17011,N_15503,N_15984);
xor U17012 (N_17012,N_15059,N_16249);
nor U17013 (N_17013,N_15588,N_15999);
or U17014 (N_17014,N_15837,N_16006);
nor U17015 (N_17015,N_15884,N_15363);
or U17016 (N_17016,N_15163,N_16138);
or U17017 (N_17017,N_15133,N_15343);
and U17018 (N_17018,N_15742,N_15481);
xor U17019 (N_17019,N_15616,N_15921);
nand U17020 (N_17020,N_15283,N_15819);
nand U17021 (N_17021,N_16050,N_15715);
nor U17022 (N_17022,N_15661,N_15686);
nor U17023 (N_17023,N_15559,N_15849);
and U17024 (N_17024,N_16129,N_15376);
nand U17025 (N_17025,N_15662,N_15516);
xor U17026 (N_17026,N_15969,N_15043);
and U17027 (N_17027,N_15469,N_15822);
nor U17028 (N_17028,N_15675,N_16167);
or U17029 (N_17029,N_15498,N_15994);
and U17030 (N_17030,N_15808,N_15017);
or U17031 (N_17031,N_15782,N_15016);
nor U17032 (N_17032,N_15422,N_16101);
nor U17033 (N_17033,N_15511,N_15145);
nand U17034 (N_17034,N_15418,N_15902);
xor U17035 (N_17035,N_15936,N_15975);
nand U17036 (N_17036,N_15916,N_16078);
xor U17037 (N_17037,N_16048,N_15348);
or U17038 (N_17038,N_15167,N_16169);
and U17039 (N_17039,N_15968,N_15261);
or U17040 (N_17040,N_15994,N_15186);
and U17041 (N_17041,N_15710,N_15754);
or U17042 (N_17042,N_15022,N_15852);
or U17043 (N_17043,N_15853,N_15377);
nor U17044 (N_17044,N_15228,N_15713);
or U17045 (N_17045,N_15470,N_15086);
or U17046 (N_17046,N_15738,N_15884);
xnor U17047 (N_17047,N_15248,N_15653);
nor U17048 (N_17048,N_15764,N_15924);
nand U17049 (N_17049,N_16081,N_15948);
or U17050 (N_17050,N_15624,N_15801);
or U17051 (N_17051,N_15662,N_16226);
nor U17052 (N_17052,N_15375,N_15311);
nand U17053 (N_17053,N_15958,N_16096);
nor U17054 (N_17054,N_15452,N_15011);
nor U17055 (N_17055,N_15409,N_16148);
and U17056 (N_17056,N_15073,N_15183);
or U17057 (N_17057,N_16022,N_15993);
xnor U17058 (N_17058,N_15342,N_15637);
or U17059 (N_17059,N_15680,N_15206);
or U17060 (N_17060,N_15798,N_15158);
xnor U17061 (N_17061,N_16235,N_15404);
nor U17062 (N_17062,N_15429,N_15857);
xnor U17063 (N_17063,N_15201,N_16084);
xor U17064 (N_17064,N_16212,N_15370);
nand U17065 (N_17065,N_16141,N_16006);
or U17066 (N_17066,N_15757,N_16125);
or U17067 (N_17067,N_15355,N_16245);
nor U17068 (N_17068,N_15975,N_15639);
or U17069 (N_17069,N_15345,N_16154);
nand U17070 (N_17070,N_15397,N_15024);
and U17071 (N_17071,N_15550,N_15584);
xnor U17072 (N_17072,N_15457,N_15068);
nor U17073 (N_17073,N_15941,N_15895);
or U17074 (N_17074,N_16129,N_15299);
or U17075 (N_17075,N_15843,N_15993);
and U17076 (N_17076,N_15146,N_16083);
xnor U17077 (N_17077,N_15528,N_16236);
nor U17078 (N_17078,N_15935,N_15638);
nand U17079 (N_17079,N_15907,N_15565);
and U17080 (N_17080,N_15463,N_15839);
nand U17081 (N_17081,N_16139,N_16082);
and U17082 (N_17082,N_15293,N_15192);
nor U17083 (N_17083,N_16228,N_15127);
or U17084 (N_17084,N_15772,N_16181);
or U17085 (N_17085,N_15443,N_16248);
and U17086 (N_17086,N_15862,N_15285);
xor U17087 (N_17087,N_16009,N_15049);
and U17088 (N_17088,N_15958,N_16197);
nor U17089 (N_17089,N_16069,N_15238);
or U17090 (N_17090,N_15972,N_16052);
and U17091 (N_17091,N_15657,N_15781);
or U17092 (N_17092,N_15590,N_15408);
or U17093 (N_17093,N_15812,N_15923);
xnor U17094 (N_17094,N_15016,N_15139);
xnor U17095 (N_17095,N_15111,N_16194);
nand U17096 (N_17096,N_15303,N_15238);
nor U17097 (N_17097,N_15508,N_15536);
xor U17098 (N_17098,N_15582,N_15209);
nand U17099 (N_17099,N_15172,N_15306);
nand U17100 (N_17100,N_15252,N_15302);
or U17101 (N_17101,N_15677,N_15758);
nor U17102 (N_17102,N_16003,N_15570);
xnor U17103 (N_17103,N_15229,N_15507);
nor U17104 (N_17104,N_15361,N_15521);
nand U17105 (N_17105,N_15924,N_15667);
and U17106 (N_17106,N_15204,N_16012);
xnor U17107 (N_17107,N_15034,N_15484);
nor U17108 (N_17108,N_16063,N_15344);
and U17109 (N_17109,N_15588,N_15199);
nand U17110 (N_17110,N_16100,N_15335);
nand U17111 (N_17111,N_16165,N_15812);
nand U17112 (N_17112,N_15875,N_16143);
xor U17113 (N_17113,N_15049,N_15317);
nor U17114 (N_17114,N_15839,N_15041);
nand U17115 (N_17115,N_15254,N_16161);
or U17116 (N_17116,N_15633,N_16183);
nor U17117 (N_17117,N_16022,N_15041);
or U17118 (N_17118,N_15233,N_15367);
nand U17119 (N_17119,N_15722,N_15505);
nor U17120 (N_17120,N_15847,N_15253);
and U17121 (N_17121,N_16117,N_15865);
nor U17122 (N_17122,N_15328,N_15144);
nor U17123 (N_17123,N_15357,N_16006);
nor U17124 (N_17124,N_16215,N_15982);
and U17125 (N_17125,N_15770,N_15847);
nand U17126 (N_17126,N_16171,N_15547);
nor U17127 (N_17127,N_15102,N_15154);
and U17128 (N_17128,N_15994,N_15237);
nor U17129 (N_17129,N_16172,N_15555);
and U17130 (N_17130,N_15711,N_15058);
and U17131 (N_17131,N_15077,N_15160);
xnor U17132 (N_17132,N_15897,N_15148);
or U17133 (N_17133,N_16244,N_15144);
or U17134 (N_17134,N_15334,N_15594);
nand U17135 (N_17135,N_15128,N_16080);
nor U17136 (N_17136,N_15776,N_15321);
nand U17137 (N_17137,N_16108,N_15788);
nor U17138 (N_17138,N_15400,N_15244);
and U17139 (N_17139,N_16105,N_15260);
and U17140 (N_17140,N_16115,N_15282);
xor U17141 (N_17141,N_15643,N_15822);
xor U17142 (N_17142,N_15866,N_15628);
xor U17143 (N_17143,N_15210,N_15359);
or U17144 (N_17144,N_15824,N_15091);
or U17145 (N_17145,N_15289,N_15472);
xnor U17146 (N_17146,N_15662,N_15502);
nor U17147 (N_17147,N_16082,N_15146);
and U17148 (N_17148,N_15914,N_15014);
nand U17149 (N_17149,N_15028,N_15643);
xor U17150 (N_17150,N_15560,N_15272);
and U17151 (N_17151,N_15700,N_16126);
nor U17152 (N_17152,N_15284,N_15624);
or U17153 (N_17153,N_15896,N_15738);
nand U17154 (N_17154,N_15192,N_15493);
or U17155 (N_17155,N_16054,N_15755);
and U17156 (N_17156,N_16087,N_15402);
nor U17157 (N_17157,N_16180,N_15876);
or U17158 (N_17158,N_16085,N_15460);
nor U17159 (N_17159,N_15227,N_15085);
or U17160 (N_17160,N_16229,N_15981);
nor U17161 (N_17161,N_15816,N_15866);
xnor U17162 (N_17162,N_15183,N_15776);
nor U17163 (N_17163,N_15760,N_15578);
xnor U17164 (N_17164,N_15096,N_15353);
nand U17165 (N_17165,N_15692,N_15930);
or U17166 (N_17166,N_15225,N_15039);
and U17167 (N_17167,N_16194,N_15787);
or U17168 (N_17168,N_16010,N_15592);
xnor U17169 (N_17169,N_16195,N_15405);
or U17170 (N_17170,N_16176,N_15371);
nand U17171 (N_17171,N_15926,N_15747);
nand U17172 (N_17172,N_15170,N_15051);
nor U17173 (N_17173,N_15378,N_16188);
xnor U17174 (N_17174,N_16175,N_16136);
nand U17175 (N_17175,N_15338,N_16229);
xor U17176 (N_17176,N_15967,N_15292);
nand U17177 (N_17177,N_16030,N_16234);
and U17178 (N_17178,N_16191,N_15271);
and U17179 (N_17179,N_16057,N_15583);
and U17180 (N_17180,N_15850,N_15178);
and U17181 (N_17181,N_15472,N_15176);
xor U17182 (N_17182,N_15834,N_15284);
nor U17183 (N_17183,N_15945,N_15240);
nand U17184 (N_17184,N_15654,N_15985);
or U17185 (N_17185,N_15979,N_15090);
and U17186 (N_17186,N_15378,N_15107);
xnor U17187 (N_17187,N_15702,N_15646);
nor U17188 (N_17188,N_16094,N_15270);
or U17189 (N_17189,N_15281,N_15856);
or U17190 (N_17190,N_15271,N_15734);
xnor U17191 (N_17191,N_15819,N_15695);
and U17192 (N_17192,N_15485,N_15994);
nand U17193 (N_17193,N_15494,N_15535);
and U17194 (N_17194,N_15448,N_15591);
xnor U17195 (N_17195,N_15026,N_15661);
or U17196 (N_17196,N_15245,N_15681);
xnor U17197 (N_17197,N_15713,N_15934);
and U17198 (N_17198,N_15228,N_15412);
xnor U17199 (N_17199,N_15723,N_15217);
or U17200 (N_17200,N_15854,N_15585);
or U17201 (N_17201,N_15730,N_15533);
nand U17202 (N_17202,N_15429,N_15381);
or U17203 (N_17203,N_15282,N_15418);
or U17204 (N_17204,N_15930,N_15706);
nand U17205 (N_17205,N_15561,N_15456);
or U17206 (N_17206,N_16189,N_15881);
nand U17207 (N_17207,N_16041,N_15937);
and U17208 (N_17208,N_15802,N_15360);
xnor U17209 (N_17209,N_15107,N_15529);
nor U17210 (N_17210,N_15751,N_15481);
nand U17211 (N_17211,N_15350,N_15330);
nor U17212 (N_17212,N_15363,N_15771);
and U17213 (N_17213,N_16172,N_15369);
nor U17214 (N_17214,N_16219,N_15597);
or U17215 (N_17215,N_15038,N_15961);
nand U17216 (N_17216,N_15458,N_15562);
and U17217 (N_17217,N_15612,N_15991);
nor U17218 (N_17218,N_16150,N_16133);
nand U17219 (N_17219,N_15333,N_15177);
or U17220 (N_17220,N_15096,N_15302);
xor U17221 (N_17221,N_15966,N_15021);
xnor U17222 (N_17222,N_16211,N_15761);
nand U17223 (N_17223,N_15617,N_15730);
and U17224 (N_17224,N_15476,N_15992);
and U17225 (N_17225,N_15014,N_15056);
xor U17226 (N_17226,N_15456,N_15758);
xor U17227 (N_17227,N_15814,N_15201);
or U17228 (N_17228,N_15892,N_15576);
nor U17229 (N_17229,N_15855,N_16130);
and U17230 (N_17230,N_16055,N_16224);
nor U17231 (N_17231,N_15342,N_15210);
or U17232 (N_17232,N_16163,N_15944);
nor U17233 (N_17233,N_15120,N_15098);
xnor U17234 (N_17234,N_16056,N_16106);
xnor U17235 (N_17235,N_16046,N_15235);
or U17236 (N_17236,N_15908,N_16052);
nand U17237 (N_17237,N_16176,N_15521);
nor U17238 (N_17238,N_15298,N_16049);
nor U17239 (N_17239,N_15313,N_15813);
nand U17240 (N_17240,N_15069,N_15439);
or U17241 (N_17241,N_16090,N_15017);
nor U17242 (N_17242,N_15351,N_16155);
and U17243 (N_17243,N_16123,N_16007);
nor U17244 (N_17244,N_15277,N_15691);
xor U17245 (N_17245,N_15799,N_15931);
or U17246 (N_17246,N_15250,N_15940);
nor U17247 (N_17247,N_16079,N_15550);
xor U17248 (N_17248,N_15763,N_15631);
or U17249 (N_17249,N_15824,N_16239);
or U17250 (N_17250,N_15234,N_15523);
and U17251 (N_17251,N_15097,N_15385);
or U17252 (N_17252,N_16127,N_15725);
nor U17253 (N_17253,N_15007,N_16209);
xnor U17254 (N_17254,N_15116,N_15034);
and U17255 (N_17255,N_15715,N_15974);
and U17256 (N_17256,N_15603,N_15532);
nand U17257 (N_17257,N_15650,N_16063);
and U17258 (N_17258,N_15426,N_15707);
and U17259 (N_17259,N_16025,N_15429);
xor U17260 (N_17260,N_15475,N_15290);
xor U17261 (N_17261,N_16097,N_15865);
nand U17262 (N_17262,N_15492,N_16056);
xnor U17263 (N_17263,N_15077,N_15492);
nand U17264 (N_17264,N_15748,N_15190);
or U17265 (N_17265,N_15483,N_16246);
nor U17266 (N_17266,N_15275,N_16018);
and U17267 (N_17267,N_15037,N_15138);
or U17268 (N_17268,N_15241,N_15360);
xor U17269 (N_17269,N_16166,N_15340);
nor U17270 (N_17270,N_15541,N_15629);
nor U17271 (N_17271,N_15730,N_15804);
nand U17272 (N_17272,N_15225,N_15124);
or U17273 (N_17273,N_15466,N_15592);
nor U17274 (N_17274,N_16156,N_15188);
and U17275 (N_17275,N_15443,N_15189);
nand U17276 (N_17276,N_15447,N_15689);
or U17277 (N_17277,N_15730,N_15261);
xor U17278 (N_17278,N_15578,N_15143);
nand U17279 (N_17279,N_15483,N_15698);
and U17280 (N_17280,N_15902,N_15787);
xnor U17281 (N_17281,N_16106,N_16059);
or U17282 (N_17282,N_16158,N_15324);
nand U17283 (N_17283,N_15434,N_15734);
or U17284 (N_17284,N_15861,N_15729);
nor U17285 (N_17285,N_16034,N_15224);
or U17286 (N_17286,N_15298,N_15057);
xnor U17287 (N_17287,N_16028,N_16169);
nand U17288 (N_17288,N_16058,N_15003);
or U17289 (N_17289,N_15254,N_16047);
nand U17290 (N_17290,N_15538,N_15040);
nand U17291 (N_17291,N_15026,N_16148);
nand U17292 (N_17292,N_16235,N_15596);
or U17293 (N_17293,N_15102,N_15758);
or U17294 (N_17294,N_15947,N_15207);
nand U17295 (N_17295,N_15864,N_15727);
nand U17296 (N_17296,N_15855,N_16046);
nor U17297 (N_17297,N_15763,N_15285);
nor U17298 (N_17298,N_15126,N_15612);
and U17299 (N_17299,N_15833,N_16169);
nor U17300 (N_17300,N_15787,N_15162);
xor U17301 (N_17301,N_15138,N_15062);
or U17302 (N_17302,N_16220,N_15968);
nor U17303 (N_17303,N_15518,N_15879);
nand U17304 (N_17304,N_16232,N_15406);
xor U17305 (N_17305,N_15561,N_15859);
xnor U17306 (N_17306,N_16034,N_15711);
or U17307 (N_17307,N_15183,N_15463);
xor U17308 (N_17308,N_15144,N_15539);
and U17309 (N_17309,N_15482,N_15810);
or U17310 (N_17310,N_15275,N_15689);
xor U17311 (N_17311,N_16053,N_15111);
or U17312 (N_17312,N_15496,N_15841);
and U17313 (N_17313,N_15047,N_15710);
nand U17314 (N_17314,N_15172,N_16221);
nor U17315 (N_17315,N_15051,N_15666);
and U17316 (N_17316,N_16249,N_15177);
or U17317 (N_17317,N_15481,N_15037);
nand U17318 (N_17318,N_16017,N_15594);
or U17319 (N_17319,N_16117,N_15239);
and U17320 (N_17320,N_15877,N_15282);
nand U17321 (N_17321,N_15634,N_16038);
or U17322 (N_17322,N_16241,N_15709);
or U17323 (N_17323,N_16243,N_15378);
nor U17324 (N_17324,N_16100,N_16197);
and U17325 (N_17325,N_15775,N_15864);
nand U17326 (N_17326,N_15480,N_15203);
nand U17327 (N_17327,N_16031,N_15414);
or U17328 (N_17328,N_15830,N_16025);
nand U17329 (N_17329,N_15559,N_16178);
and U17330 (N_17330,N_15208,N_15735);
xor U17331 (N_17331,N_15908,N_15928);
nand U17332 (N_17332,N_16094,N_15055);
and U17333 (N_17333,N_15465,N_15606);
or U17334 (N_17334,N_15326,N_16023);
xnor U17335 (N_17335,N_15320,N_15401);
xor U17336 (N_17336,N_15018,N_15545);
nand U17337 (N_17337,N_15249,N_15990);
xnor U17338 (N_17338,N_15878,N_15422);
nor U17339 (N_17339,N_16141,N_15415);
nand U17340 (N_17340,N_15866,N_15844);
nor U17341 (N_17341,N_15057,N_16168);
and U17342 (N_17342,N_16060,N_15059);
or U17343 (N_17343,N_15447,N_15892);
and U17344 (N_17344,N_15824,N_15034);
and U17345 (N_17345,N_15500,N_15394);
xnor U17346 (N_17346,N_15588,N_15461);
or U17347 (N_17347,N_16139,N_15269);
nand U17348 (N_17348,N_16136,N_15856);
or U17349 (N_17349,N_16138,N_15215);
and U17350 (N_17350,N_15502,N_15791);
xnor U17351 (N_17351,N_15438,N_15535);
xnor U17352 (N_17352,N_15133,N_15390);
nor U17353 (N_17353,N_15019,N_15574);
nand U17354 (N_17354,N_15268,N_15091);
nand U17355 (N_17355,N_15818,N_15602);
nor U17356 (N_17356,N_16248,N_15853);
nor U17357 (N_17357,N_15145,N_16073);
xor U17358 (N_17358,N_15106,N_15467);
nor U17359 (N_17359,N_15626,N_15795);
xor U17360 (N_17360,N_15043,N_15783);
and U17361 (N_17361,N_15292,N_15822);
xor U17362 (N_17362,N_16181,N_15140);
nand U17363 (N_17363,N_15727,N_15656);
nor U17364 (N_17364,N_15003,N_15350);
and U17365 (N_17365,N_15419,N_15380);
nand U17366 (N_17366,N_15471,N_15413);
xnor U17367 (N_17367,N_15633,N_16102);
and U17368 (N_17368,N_16130,N_16011);
nor U17369 (N_17369,N_15694,N_15874);
nand U17370 (N_17370,N_15106,N_15729);
or U17371 (N_17371,N_15951,N_15255);
nand U17372 (N_17372,N_15245,N_16122);
and U17373 (N_17373,N_15588,N_16146);
nand U17374 (N_17374,N_16060,N_15232);
or U17375 (N_17375,N_15907,N_16193);
and U17376 (N_17376,N_15618,N_15962);
and U17377 (N_17377,N_15986,N_15869);
or U17378 (N_17378,N_15958,N_15270);
and U17379 (N_17379,N_15801,N_15360);
nor U17380 (N_17380,N_15041,N_16128);
or U17381 (N_17381,N_16244,N_15341);
and U17382 (N_17382,N_16151,N_15941);
or U17383 (N_17383,N_16168,N_15873);
nand U17384 (N_17384,N_15626,N_15163);
nor U17385 (N_17385,N_15176,N_15005);
nand U17386 (N_17386,N_15559,N_16203);
or U17387 (N_17387,N_15059,N_15169);
nand U17388 (N_17388,N_15566,N_15880);
or U17389 (N_17389,N_15069,N_15247);
xnor U17390 (N_17390,N_15501,N_16188);
nand U17391 (N_17391,N_15574,N_15600);
nor U17392 (N_17392,N_15402,N_15958);
or U17393 (N_17393,N_16223,N_15718);
xor U17394 (N_17394,N_16228,N_16176);
xor U17395 (N_17395,N_15692,N_15963);
and U17396 (N_17396,N_15485,N_16094);
or U17397 (N_17397,N_16189,N_15049);
and U17398 (N_17398,N_16053,N_15864);
or U17399 (N_17399,N_15029,N_16053);
nand U17400 (N_17400,N_16243,N_16017);
nand U17401 (N_17401,N_15300,N_16062);
nand U17402 (N_17402,N_15039,N_15592);
xor U17403 (N_17403,N_15547,N_16231);
xnor U17404 (N_17404,N_15698,N_16058);
nor U17405 (N_17405,N_15423,N_16083);
xnor U17406 (N_17406,N_15568,N_15843);
nand U17407 (N_17407,N_15146,N_15864);
xnor U17408 (N_17408,N_15848,N_15874);
xnor U17409 (N_17409,N_15766,N_15054);
nor U17410 (N_17410,N_16225,N_15579);
xnor U17411 (N_17411,N_15649,N_15656);
or U17412 (N_17412,N_15191,N_15360);
or U17413 (N_17413,N_15762,N_16211);
and U17414 (N_17414,N_15753,N_15206);
nor U17415 (N_17415,N_16189,N_15803);
and U17416 (N_17416,N_15685,N_15041);
or U17417 (N_17417,N_15217,N_15299);
or U17418 (N_17418,N_15201,N_15251);
nand U17419 (N_17419,N_15904,N_15415);
xor U17420 (N_17420,N_16062,N_16031);
or U17421 (N_17421,N_15370,N_15504);
or U17422 (N_17422,N_15503,N_15298);
nand U17423 (N_17423,N_15720,N_15267);
and U17424 (N_17424,N_15709,N_15571);
and U17425 (N_17425,N_15664,N_15115);
xnor U17426 (N_17426,N_15322,N_15567);
nor U17427 (N_17427,N_15047,N_15233);
or U17428 (N_17428,N_15049,N_16176);
xor U17429 (N_17429,N_15178,N_15724);
or U17430 (N_17430,N_15671,N_15141);
or U17431 (N_17431,N_15927,N_15332);
or U17432 (N_17432,N_15390,N_15141);
nand U17433 (N_17433,N_16205,N_16070);
and U17434 (N_17434,N_15237,N_15321);
nand U17435 (N_17435,N_15404,N_15633);
and U17436 (N_17436,N_16212,N_16041);
nor U17437 (N_17437,N_15490,N_15785);
nor U17438 (N_17438,N_15633,N_15961);
or U17439 (N_17439,N_15275,N_15088);
nor U17440 (N_17440,N_15421,N_16226);
xor U17441 (N_17441,N_15339,N_15595);
nand U17442 (N_17442,N_15050,N_15336);
nor U17443 (N_17443,N_15913,N_16064);
and U17444 (N_17444,N_15014,N_16200);
nand U17445 (N_17445,N_15733,N_15179);
xnor U17446 (N_17446,N_15085,N_15178);
or U17447 (N_17447,N_15692,N_15395);
nand U17448 (N_17448,N_15596,N_15742);
or U17449 (N_17449,N_15003,N_15231);
nor U17450 (N_17450,N_16162,N_15115);
and U17451 (N_17451,N_16209,N_15925);
or U17452 (N_17452,N_15814,N_16060);
and U17453 (N_17453,N_15576,N_15321);
xnor U17454 (N_17454,N_15861,N_16079);
xnor U17455 (N_17455,N_15925,N_15326);
or U17456 (N_17456,N_15280,N_15851);
and U17457 (N_17457,N_15409,N_15341);
xor U17458 (N_17458,N_15928,N_15745);
xnor U17459 (N_17459,N_15454,N_15748);
and U17460 (N_17460,N_16053,N_16046);
nor U17461 (N_17461,N_15892,N_15244);
and U17462 (N_17462,N_15474,N_15112);
xor U17463 (N_17463,N_15921,N_15612);
nor U17464 (N_17464,N_15885,N_15032);
or U17465 (N_17465,N_15143,N_15550);
or U17466 (N_17466,N_16073,N_15439);
and U17467 (N_17467,N_15992,N_15548);
xor U17468 (N_17468,N_15398,N_15783);
xor U17469 (N_17469,N_15541,N_15264);
xor U17470 (N_17470,N_15702,N_15081);
xor U17471 (N_17471,N_15306,N_15126);
nor U17472 (N_17472,N_15535,N_15869);
nor U17473 (N_17473,N_15320,N_15300);
xor U17474 (N_17474,N_15220,N_15460);
xnor U17475 (N_17475,N_16114,N_15615);
and U17476 (N_17476,N_16103,N_15546);
and U17477 (N_17477,N_15528,N_15325);
and U17478 (N_17478,N_15096,N_16197);
or U17479 (N_17479,N_15570,N_15107);
nand U17480 (N_17480,N_15834,N_15408);
nand U17481 (N_17481,N_15682,N_15779);
nand U17482 (N_17482,N_15727,N_15185);
nand U17483 (N_17483,N_15398,N_16107);
xnor U17484 (N_17484,N_15408,N_16104);
nand U17485 (N_17485,N_15175,N_15699);
and U17486 (N_17486,N_15925,N_15121);
and U17487 (N_17487,N_15837,N_15595);
and U17488 (N_17488,N_16207,N_15993);
nand U17489 (N_17489,N_15437,N_16181);
nor U17490 (N_17490,N_15682,N_15819);
nor U17491 (N_17491,N_15437,N_15187);
xnor U17492 (N_17492,N_15210,N_16157);
xnor U17493 (N_17493,N_16166,N_15118);
nor U17494 (N_17494,N_16209,N_15915);
xnor U17495 (N_17495,N_15263,N_15423);
xnor U17496 (N_17496,N_15266,N_15045);
nand U17497 (N_17497,N_15018,N_15399);
nor U17498 (N_17498,N_15037,N_16103);
nor U17499 (N_17499,N_15999,N_15916);
and U17500 (N_17500,N_16919,N_17249);
or U17501 (N_17501,N_16298,N_17258);
and U17502 (N_17502,N_17053,N_16261);
nor U17503 (N_17503,N_16567,N_17073);
nand U17504 (N_17504,N_16510,N_16425);
nor U17505 (N_17505,N_16702,N_17209);
and U17506 (N_17506,N_17194,N_17305);
nand U17507 (N_17507,N_16503,N_16630);
or U17508 (N_17508,N_16553,N_17479);
nand U17509 (N_17509,N_17114,N_17317);
or U17510 (N_17510,N_17267,N_17004);
xnor U17511 (N_17511,N_17302,N_17311);
nor U17512 (N_17512,N_16789,N_16308);
or U17513 (N_17513,N_17106,N_17374);
nor U17514 (N_17514,N_16356,N_17420);
or U17515 (N_17515,N_16421,N_16945);
nand U17516 (N_17516,N_17085,N_17163);
xor U17517 (N_17517,N_17191,N_17327);
nand U17518 (N_17518,N_16586,N_17307);
nor U17519 (N_17519,N_16722,N_17429);
xor U17520 (N_17520,N_16764,N_16451);
nand U17521 (N_17521,N_16666,N_17326);
nor U17522 (N_17522,N_17182,N_16832);
xor U17523 (N_17523,N_17202,N_16639);
and U17524 (N_17524,N_16924,N_17329);
and U17525 (N_17525,N_16416,N_17125);
nand U17526 (N_17526,N_17021,N_17160);
nand U17527 (N_17527,N_16342,N_17447);
and U17528 (N_17528,N_17104,N_16929);
xnor U17529 (N_17529,N_17487,N_16760);
or U17530 (N_17530,N_16754,N_16957);
xnor U17531 (N_17531,N_16500,N_16256);
and U17532 (N_17532,N_17460,N_17469);
and U17533 (N_17533,N_16437,N_17240);
or U17534 (N_17534,N_16881,N_16828);
xor U17535 (N_17535,N_16493,N_16858);
or U17536 (N_17536,N_17219,N_17224);
nor U17537 (N_17537,N_17483,N_16439);
and U17538 (N_17538,N_16662,N_16676);
nor U17539 (N_17539,N_17001,N_16649);
nand U17540 (N_17540,N_17471,N_16583);
and U17541 (N_17541,N_17366,N_16856);
and U17542 (N_17542,N_17150,N_16575);
nand U17543 (N_17543,N_16501,N_17410);
nor U17544 (N_17544,N_16885,N_16637);
or U17545 (N_17545,N_16732,N_16407);
or U17546 (N_17546,N_16449,N_17119);
nor U17547 (N_17547,N_16365,N_16391);
and U17548 (N_17548,N_17061,N_16867);
nor U17549 (N_17549,N_16375,N_17003);
and U17550 (N_17550,N_17454,N_16955);
nor U17551 (N_17551,N_16672,N_16737);
or U17552 (N_17552,N_16406,N_16580);
nand U17553 (N_17553,N_16530,N_17443);
and U17554 (N_17554,N_16681,N_17079);
nor U17555 (N_17555,N_16762,N_16515);
nand U17556 (N_17556,N_17264,N_17288);
xor U17557 (N_17557,N_17399,N_17072);
and U17558 (N_17558,N_16331,N_17415);
nand U17559 (N_17559,N_16875,N_17105);
xor U17560 (N_17560,N_16834,N_17455);
xor U17561 (N_17561,N_16922,N_16665);
xnor U17562 (N_17562,N_16829,N_16934);
nand U17563 (N_17563,N_16611,N_16804);
or U17564 (N_17564,N_17394,N_16748);
nor U17565 (N_17565,N_17017,N_16911);
nand U17566 (N_17566,N_17301,N_16673);
and U17567 (N_17567,N_17295,N_17041);
or U17568 (N_17568,N_16470,N_17115);
or U17569 (N_17569,N_16953,N_16276);
or U17570 (N_17570,N_16363,N_17364);
or U17571 (N_17571,N_17177,N_16593);
or U17572 (N_17572,N_16606,N_16374);
and U17573 (N_17573,N_17151,N_16733);
xor U17574 (N_17574,N_17395,N_17109);
nor U17575 (N_17575,N_16327,N_16688);
xor U17576 (N_17576,N_17449,N_16860);
or U17577 (N_17577,N_17344,N_17475);
nor U17578 (N_17578,N_16344,N_16967);
or U17579 (N_17579,N_16863,N_17051);
nor U17580 (N_17580,N_16976,N_17189);
or U17581 (N_17581,N_16284,N_17254);
nand U17582 (N_17582,N_17250,N_17405);
nor U17583 (N_17583,N_16488,N_16476);
xnor U17584 (N_17584,N_17430,N_17141);
nor U17585 (N_17585,N_17088,N_16660);
nand U17586 (N_17586,N_17083,N_16337);
and U17587 (N_17587,N_17232,N_16265);
and U17588 (N_17588,N_16800,N_17494);
or U17589 (N_17589,N_16694,N_16349);
nor U17590 (N_17590,N_16625,N_16559);
and U17591 (N_17591,N_16727,N_17108);
nor U17592 (N_17592,N_16290,N_17378);
nor U17593 (N_17593,N_16474,N_17368);
or U17594 (N_17594,N_16802,N_16358);
xor U17595 (N_17595,N_16378,N_16765);
or U17596 (N_17596,N_17414,N_16274);
xnor U17597 (N_17597,N_16752,N_16538);
nor U17598 (N_17598,N_16939,N_16490);
nand U17599 (N_17599,N_16835,N_16321);
nand U17600 (N_17600,N_17094,N_17229);
xnor U17601 (N_17601,N_16977,N_16706);
and U17602 (N_17602,N_16255,N_17300);
nor U17603 (N_17603,N_17486,N_17245);
nand U17604 (N_17604,N_16990,N_17413);
or U17605 (N_17605,N_17011,N_16844);
nor U17606 (N_17606,N_16669,N_16726);
nand U17607 (N_17607,N_16779,N_17318);
and U17608 (N_17608,N_17123,N_16289);
and U17609 (N_17609,N_16724,N_16352);
and U17610 (N_17610,N_16679,N_17193);
or U17611 (N_17611,N_16972,N_16292);
nand U17612 (N_17612,N_16277,N_16812);
or U17613 (N_17613,N_17116,N_16404);
nor U17614 (N_17614,N_16604,N_16560);
or U17615 (N_17615,N_16578,N_16790);
and U17616 (N_17616,N_16833,N_16279);
or U17617 (N_17617,N_17265,N_17183);
nor U17618 (N_17618,N_16591,N_17384);
nand U17619 (N_17619,N_16787,N_17101);
nand U17620 (N_17620,N_16808,N_16550);
xnor U17621 (N_17621,N_16565,N_16629);
xnor U17622 (N_17622,N_17392,N_16393);
or U17623 (N_17623,N_16302,N_16831);
xor U17624 (N_17624,N_16543,N_16545);
or U17625 (N_17625,N_17120,N_17274);
nor U17626 (N_17626,N_16661,N_17199);
nand U17627 (N_17627,N_17030,N_16433);
xnor U17628 (N_17628,N_17185,N_16896);
and U17629 (N_17629,N_17146,N_17165);
nand U17630 (N_17630,N_17338,N_16791);
nand U17631 (N_17631,N_16343,N_17018);
nor U17632 (N_17632,N_17337,N_17153);
and U17633 (N_17633,N_16264,N_17351);
nand U17634 (N_17634,N_16719,N_16315);
and U17635 (N_17635,N_16564,N_16674);
xnor U17636 (N_17636,N_17465,N_17349);
xnor U17637 (N_17637,N_17458,N_17196);
or U17638 (N_17638,N_16305,N_17381);
and U17639 (N_17639,N_16963,N_16778);
or U17640 (N_17640,N_16400,N_16506);
xnor U17641 (N_17641,N_16615,N_16784);
or U17642 (N_17642,N_16278,N_17498);
or U17643 (N_17643,N_16381,N_17331);
and U17644 (N_17644,N_16685,N_17000);
or U17645 (N_17645,N_17359,N_16857);
or U17646 (N_17646,N_16263,N_17304);
xnor U17647 (N_17647,N_16524,N_16462);
nor U17648 (N_17648,N_16577,N_16621);
or U17649 (N_17649,N_17316,N_17416);
nand U17650 (N_17650,N_16325,N_17169);
or U17651 (N_17651,N_16413,N_17371);
nor U17652 (N_17652,N_17157,N_17425);
or U17653 (N_17653,N_16979,N_16709);
nor U17654 (N_17654,N_16902,N_17480);
or U17655 (N_17655,N_16599,N_17323);
or U17656 (N_17656,N_17277,N_16392);
xor U17657 (N_17657,N_16909,N_16347);
or U17658 (N_17658,N_17499,N_17459);
nand U17659 (N_17659,N_16452,N_17409);
nor U17660 (N_17660,N_16521,N_16633);
xnor U17661 (N_17661,N_16584,N_16890);
nand U17662 (N_17662,N_17071,N_16923);
xor U17663 (N_17663,N_16539,N_16552);
nand U17664 (N_17664,N_16982,N_17358);
and U17665 (N_17665,N_17045,N_17043);
or U17666 (N_17666,N_16980,N_16956);
and U17667 (N_17667,N_16964,N_16382);
nor U17668 (N_17668,N_16253,N_16262);
nor U17669 (N_17669,N_17015,N_16782);
or U17670 (N_17670,N_16477,N_16431);
xnor U17671 (N_17671,N_17036,N_16288);
or U17672 (N_17672,N_16949,N_16542);
nor U17673 (N_17673,N_16683,N_17127);
nand U17674 (N_17674,N_17315,N_17291);
and U17675 (N_17675,N_16984,N_16974);
nor U17676 (N_17676,N_17067,N_16512);
nor U17677 (N_17677,N_17089,N_16489);
xnor U17678 (N_17678,N_16294,N_16950);
nand U17679 (N_17679,N_16386,N_16794);
xor U17680 (N_17680,N_16395,N_16655);
or U17681 (N_17681,N_16322,N_16658);
xor U17682 (N_17682,N_16721,N_17367);
nand U17683 (N_17683,N_17238,N_16314);
xor U17684 (N_17684,N_16941,N_16704);
nand U17685 (N_17685,N_17439,N_17333);
nor U17686 (N_17686,N_17027,N_16566);
or U17687 (N_17687,N_16952,N_16893);
or U17688 (N_17688,N_16817,N_17213);
nor U17689 (N_17689,N_17342,N_16320);
nor U17690 (N_17690,N_17350,N_16531);
and U17691 (N_17691,N_16642,N_16291);
nand U17692 (N_17692,N_16426,N_16366);
or U17693 (N_17693,N_17107,N_16275);
nand U17694 (N_17694,N_16297,N_17453);
nor U17695 (N_17695,N_16544,N_16364);
or U17696 (N_17696,N_17320,N_16464);
or U17697 (N_17697,N_17297,N_16485);
nor U17698 (N_17698,N_16991,N_16837);
xor U17699 (N_17699,N_16403,N_16745);
nor U17700 (N_17700,N_17222,N_16390);
xnor U17701 (N_17701,N_16852,N_17407);
or U17702 (N_17702,N_16914,N_16333);
nand U17703 (N_17703,N_17086,N_16409);
or U17704 (N_17704,N_16698,N_16851);
nand U17705 (N_17705,N_16269,N_17215);
xnor U17706 (N_17706,N_17248,N_16897);
nand U17707 (N_17707,N_17180,N_17275);
xor U17708 (N_17708,N_16329,N_17192);
nand U17709 (N_17709,N_16361,N_17207);
nor U17710 (N_17710,N_17226,N_17477);
nand U17711 (N_17711,N_17012,N_17048);
xor U17712 (N_17712,N_16626,N_17237);
nor U17713 (N_17713,N_17408,N_16747);
nor U17714 (N_17714,N_16995,N_17398);
and U17715 (N_17715,N_16346,N_17009);
and U17716 (N_17716,N_17314,N_16847);
xnor U17717 (N_17717,N_17322,N_16813);
or U17718 (N_17718,N_16594,N_16440);
and U17719 (N_17719,N_16855,N_16774);
and U17720 (N_17720,N_16958,N_17198);
nand U17721 (N_17721,N_16954,N_17122);
and U17722 (N_17722,N_17339,N_16609);
and U17723 (N_17723,N_16743,N_16285);
xnor U17724 (N_17724,N_16323,N_17039);
nand U17725 (N_17725,N_17375,N_16251);
xnor U17726 (N_17726,N_17336,N_17441);
and U17727 (N_17727,N_16635,N_16921);
nand U17728 (N_17728,N_17343,N_16551);
or U17729 (N_17729,N_16891,N_16799);
and U17730 (N_17730,N_16355,N_17357);
xnor U17731 (N_17731,N_16286,N_16648);
nor U17732 (N_17732,N_17485,N_17402);
nand U17733 (N_17733,N_17142,N_16898);
nand U17734 (N_17734,N_16751,N_17445);
and U17735 (N_17735,N_17247,N_17423);
nor U17736 (N_17736,N_17369,N_17093);
xor U17737 (N_17737,N_17286,N_17195);
nand U17738 (N_17738,N_17020,N_16418);
and U17739 (N_17739,N_16618,N_17493);
xnor U17740 (N_17740,N_16311,N_17280);
xnor U17741 (N_17741,N_17137,N_17260);
and U17742 (N_17742,N_16458,N_16427);
xnor U17743 (N_17743,N_16689,N_17034);
nand U17744 (N_17744,N_17065,N_17457);
xor U17745 (N_17745,N_16714,N_16496);
xor U17746 (N_17746,N_16519,N_17121);
and U17747 (N_17747,N_17404,N_16970);
xor U17748 (N_17748,N_17438,N_16708);
or U17749 (N_17749,N_16918,N_16492);
xnor U17750 (N_17750,N_17356,N_16874);
or U17751 (N_17751,N_17325,N_16613);
nand U17752 (N_17752,N_17396,N_17190);
or U17753 (N_17753,N_16870,N_16465);
and U17754 (N_17754,N_17411,N_16405);
nor U17755 (N_17755,N_16723,N_17118);
nand U17756 (N_17756,N_16917,N_16810);
nor U17757 (N_17757,N_16283,N_16394);
nor U17758 (N_17758,N_16942,N_16252);
nor U17759 (N_17759,N_17270,N_17095);
nand U17760 (N_17760,N_16818,N_16367);
and U17761 (N_17761,N_16450,N_16282);
nand U17762 (N_17762,N_17446,N_16482);
nand U17763 (N_17763,N_17383,N_16505);
and U17764 (N_17764,N_17138,N_17058);
or U17765 (N_17765,N_16534,N_16484);
nand U17766 (N_17766,N_16310,N_16650);
nand U17767 (N_17767,N_17059,N_17129);
or U17768 (N_17768,N_17289,N_16735);
and U17769 (N_17769,N_17225,N_17328);
nor U17770 (N_17770,N_17309,N_17484);
nor U17771 (N_17771,N_16581,N_16771);
and U17772 (N_17772,N_17023,N_16362);
and U17773 (N_17773,N_16697,N_16354);
nand U17774 (N_17774,N_17162,N_17388);
or U17775 (N_17775,N_17155,N_17126);
and U17776 (N_17776,N_16905,N_16792);
nand U17777 (N_17777,N_16775,N_16975);
or U17778 (N_17778,N_17397,N_16499);
or U17779 (N_17779,N_16461,N_16640);
and U17780 (N_17780,N_16785,N_17365);
nor U17781 (N_17781,N_16357,N_17296);
or U17782 (N_17782,N_17158,N_16563);
or U17783 (N_17783,N_16360,N_16827);
or U17784 (N_17784,N_17269,N_16997);
nand U17785 (N_17785,N_16925,N_17348);
nor U17786 (N_17786,N_17271,N_16260);
or U17787 (N_17787,N_17131,N_17178);
nor U17788 (N_17788,N_16987,N_16872);
xnor U17789 (N_17789,N_16595,N_17244);
nand U17790 (N_17790,N_16882,N_16861);
nor U17791 (N_17791,N_16610,N_17235);
nor U17792 (N_17792,N_16744,N_16809);
or U17793 (N_17793,N_16585,N_16388);
nand U17794 (N_17794,N_17252,N_16340);
and U17795 (N_17795,N_16444,N_17354);
xnor U17796 (N_17796,N_17451,N_17046);
nor U17797 (N_17797,N_17223,N_17102);
nand U17798 (N_17798,N_16466,N_17230);
or U17799 (N_17799,N_16996,N_17361);
xnor U17800 (N_17800,N_16836,N_17400);
nand U17801 (N_17801,N_16498,N_16372);
or U17802 (N_17802,N_17419,N_16823);
and U17803 (N_17803,N_16319,N_16687);
nor U17804 (N_17804,N_16756,N_16336);
nand U17805 (N_17805,N_16773,N_17171);
or U17806 (N_17806,N_16401,N_17139);
nand U17807 (N_17807,N_17170,N_16940);
xnor U17808 (N_17808,N_16371,N_17476);
and U17809 (N_17809,N_17426,N_16569);
and U17810 (N_17810,N_16700,N_16454);
or U17811 (N_17811,N_16713,N_16624);
nand U17812 (N_17812,N_16463,N_17172);
xnor U17813 (N_17813,N_16938,N_17389);
nor U17814 (N_17814,N_16522,N_17492);
or U17815 (N_17815,N_16259,N_17422);
xnor U17816 (N_17816,N_16717,N_17181);
and U17817 (N_17817,N_16258,N_16992);
and U17818 (N_17818,N_16758,N_16328);
or U17819 (N_17819,N_17303,N_16969);
or U17820 (N_17820,N_17334,N_17042);
and U17821 (N_17821,N_16478,N_16889);
and U17822 (N_17822,N_16888,N_17418);
xnor U17823 (N_17823,N_17208,N_16759);
nand U17824 (N_17824,N_17243,N_16845);
nand U17825 (N_17825,N_16541,N_17362);
or U17826 (N_17826,N_16561,N_16699);
or U17827 (N_17827,N_17332,N_16414);
nor U17828 (N_17828,N_16479,N_17294);
and U17829 (N_17829,N_16632,N_17062);
and U17830 (N_17830,N_16999,N_16616);
xnor U17831 (N_17831,N_16769,N_16816);
nand U17832 (N_17832,N_16307,N_16517);
nor U17833 (N_17833,N_17080,N_16623);
and U17834 (N_17834,N_16266,N_17002);
nand U17835 (N_17835,N_16849,N_16460);
or U17836 (N_17836,N_16312,N_16718);
and U17837 (N_17837,N_16965,N_16815);
and U17838 (N_17838,N_17482,N_16555);
xor U17839 (N_17839,N_16293,N_16304);
or U17840 (N_17840,N_16504,N_16537);
nand U17841 (N_17841,N_17214,N_16877);
nand U17842 (N_17842,N_16927,N_17149);
and U17843 (N_17843,N_17259,N_17112);
or U17844 (N_17844,N_17087,N_16664);
or U17845 (N_17845,N_16608,N_16494);
and U17846 (N_17846,N_16895,N_17014);
nor U17847 (N_17847,N_16518,N_16651);
and U17848 (N_17848,N_16430,N_17161);
and U17849 (N_17849,N_17006,N_16634);
and U17850 (N_17850,N_16830,N_16947);
or U17851 (N_17851,N_16273,N_16620);
and U17852 (N_17852,N_16571,N_16894);
nand U17853 (N_17853,N_16472,N_16600);
and U17854 (N_17854,N_17287,N_17273);
xnor U17855 (N_17855,N_17175,N_17033);
or U17856 (N_17856,N_17216,N_17013);
and U17857 (N_17857,N_16971,N_17231);
and U17858 (N_17858,N_17292,N_16840);
and U17859 (N_17859,N_17032,N_17052);
or U17860 (N_17860,N_16776,N_16267);
nor U17861 (N_17861,N_17204,N_16998);
and U17862 (N_17862,N_16842,N_16960);
or U17863 (N_17863,N_16481,N_16385);
nor U17864 (N_17864,N_16912,N_17421);
xor U17865 (N_17865,N_16767,N_17470);
nor U17866 (N_17866,N_16287,N_16904);
xor U17867 (N_17867,N_16422,N_16495);
nand U17868 (N_17868,N_16824,N_17187);
xor U17869 (N_17869,N_17372,N_17076);
nor U17870 (N_17870,N_16428,N_16766);
or U17871 (N_17871,N_16846,N_16369);
and U17872 (N_17872,N_17025,N_17074);
xnor U17873 (N_17873,N_17016,N_17424);
and U17874 (N_17874,N_16303,N_16738);
nor U17875 (N_17875,N_17377,N_17136);
nor U17876 (N_17876,N_17462,N_16468);
nand U17877 (N_17877,N_16690,N_17330);
nor U17878 (N_17878,N_17113,N_17444);
and U17879 (N_17879,N_17026,N_16734);
and U17880 (N_17880,N_17242,N_16497);
xnor U17881 (N_17881,N_16612,N_17463);
xnor U17882 (N_17882,N_16729,N_16777);
and U17883 (N_17883,N_16944,N_16602);
nor U17884 (N_17884,N_16408,N_16605);
and U17885 (N_17885,N_16254,N_16597);
nor U17886 (N_17886,N_16682,N_16926);
nor U17887 (N_17887,N_16350,N_16480);
nor U17888 (N_17888,N_17096,N_17263);
nand U17889 (N_17889,N_17154,N_16715);
or U17890 (N_17890,N_17346,N_17256);
xor U17891 (N_17891,N_17024,N_16712);
xor U17892 (N_17892,N_17128,N_16742);
and U17893 (N_17893,N_16380,N_16703);
nand U17894 (N_17894,N_16780,N_17452);
nor U17895 (N_17895,N_16410,N_16438);
and U17896 (N_17896,N_16788,N_16272);
xor U17897 (N_17897,N_17218,N_16839);
nand U17898 (N_17898,N_17220,N_16859);
nand U17899 (N_17899,N_16317,N_17272);
xor U17900 (N_17900,N_17166,N_16528);
nor U17901 (N_17901,N_17335,N_16508);
xnor U17902 (N_17902,N_16579,N_16707);
nor U17903 (N_17903,N_16959,N_16781);
xnor U17904 (N_17904,N_16384,N_16516);
and U17905 (N_17905,N_16486,N_17082);
and U17906 (N_17906,N_16985,N_17049);
nor U17907 (N_17907,N_16659,N_17246);
nor U17908 (N_17908,N_17491,N_16822);
or U17909 (N_17909,N_16526,N_16915);
and U17910 (N_17910,N_17077,N_17070);
nand U17911 (N_17911,N_16424,N_16736);
xnor U17912 (N_17912,N_16644,N_16843);
xor U17913 (N_17913,N_17437,N_16880);
or U17914 (N_17914,N_17047,N_17299);
nand U17915 (N_17915,N_17478,N_16383);
nor U17916 (N_17916,N_16653,N_17253);
nand U17917 (N_17917,N_16379,N_17037);
nand U17918 (N_17918,N_17075,N_17298);
nand U17919 (N_17919,N_16373,N_17210);
nor U17920 (N_17920,N_17063,N_17186);
or U17921 (N_17921,N_17417,N_16483);
or U17922 (N_17922,N_16436,N_17228);
xnor U17923 (N_17923,N_16692,N_16798);
nor U17924 (N_17924,N_16596,N_16368);
or U17925 (N_17925,N_17031,N_16740);
xor U17926 (N_17926,N_17393,N_16670);
nand U17927 (N_17927,N_16582,N_17261);
or U17928 (N_17928,N_16507,N_16749);
nand U17929 (N_17929,N_16806,N_16535);
nand U17930 (N_17930,N_17403,N_16547);
xor U17931 (N_17931,N_17436,N_17130);
and U17932 (N_17932,N_16901,N_17285);
or U17933 (N_17933,N_16351,N_16913);
xnor U17934 (N_17934,N_16533,N_16864);
xor U17935 (N_17935,N_16961,N_16930);
nand U17936 (N_17936,N_17290,N_16928);
xor U17937 (N_17937,N_16502,N_17467);
and U17938 (N_17938,N_17078,N_16614);
and U17939 (N_17939,N_16487,N_16441);
xor U17940 (N_17940,N_17255,N_17293);
xor U17941 (N_17941,N_16326,N_16455);
or U17942 (N_17942,N_16335,N_17352);
xnor U17943 (N_17943,N_17066,N_16932);
and U17944 (N_17944,N_16663,N_17283);
nand U17945 (N_17945,N_17321,N_16309);
xor U17946 (N_17946,N_16916,N_16948);
xor U17947 (N_17947,N_16467,N_16741);
nor U17948 (N_17948,N_17111,N_16617);
xnor U17949 (N_17949,N_16862,N_17200);
xnor U17950 (N_17950,N_17168,N_16257);
and U17951 (N_17951,N_16576,N_17188);
and U17952 (N_17952,N_16796,N_17466);
and U17953 (N_17953,N_16886,N_17308);
and U17954 (N_17954,N_17450,N_16590);
and U17955 (N_17955,N_17092,N_16803);
nand U17956 (N_17956,N_17100,N_16807);
nor U17957 (N_17957,N_17117,N_17488);
and U17958 (N_17958,N_16491,N_17347);
or U17959 (N_17959,N_16339,N_16429);
or U17960 (N_17960,N_16701,N_16968);
or U17961 (N_17961,N_17205,N_17028);
or U17962 (N_17962,N_17435,N_16962);
and U17963 (N_17963,N_17068,N_17373);
nand U17964 (N_17964,N_17167,N_16795);
and U17965 (N_17965,N_16471,N_17428);
or U17966 (N_17966,N_16819,N_16641);
or U17967 (N_17967,N_17135,N_17279);
xor U17968 (N_17968,N_16556,N_16281);
xor U17969 (N_17969,N_17174,N_17251);
xor U17970 (N_17970,N_16296,N_17029);
xor U17971 (N_17971,N_17145,N_16306);
nand U17972 (N_17972,N_16850,N_16873);
nand U17973 (N_17973,N_17490,N_16876);
nor U17974 (N_17974,N_17427,N_16983);
nor U17975 (N_17975,N_16443,N_17044);
nor U17976 (N_17976,N_16359,N_16562);
and U17977 (N_17977,N_17184,N_16448);
nor U17978 (N_17978,N_17412,N_16899);
nand U17979 (N_17979,N_16668,N_17211);
or U17980 (N_17980,N_16398,N_16509);
nor U17981 (N_17981,N_16417,N_17432);
nand U17982 (N_17982,N_17387,N_17098);
or U17983 (N_17983,N_16786,N_16270);
xnor U17984 (N_17984,N_16866,N_16667);
and U17985 (N_17985,N_17008,N_17440);
nor U17986 (N_17986,N_17081,N_17156);
and U17987 (N_17987,N_17266,N_17050);
xor U17988 (N_17988,N_16387,N_17313);
or U17989 (N_17989,N_16397,N_16936);
or U17990 (N_17990,N_16520,N_16447);
or U17991 (N_17991,N_17385,N_16946);
or U17992 (N_17992,N_16678,N_16989);
nor U17993 (N_17993,N_17110,N_17007);
xnor U17994 (N_17994,N_16636,N_17379);
nand U17995 (N_17995,N_17143,N_16299);
nor U17996 (N_17996,N_16783,N_16511);
and U17997 (N_17997,N_17091,N_17284);
or U17998 (N_17998,N_16432,N_17360);
nor U17999 (N_17999,N_16330,N_16601);
or U18000 (N_18000,N_16820,N_17281);
nor U18001 (N_18001,N_16825,N_16316);
or U18002 (N_18002,N_17084,N_16536);
and U18003 (N_18003,N_17464,N_16988);
nand U18004 (N_18004,N_17431,N_16838);
nor U18005 (N_18005,N_17386,N_17054);
xnor U18006 (N_18006,N_16973,N_16978);
xor U18007 (N_18007,N_16892,N_16592);
nor U18008 (N_18008,N_16710,N_17233);
or U18009 (N_18009,N_17495,N_16728);
or U18010 (N_18010,N_17282,N_17227);
nand U18011 (N_18011,N_17497,N_17234);
or U18012 (N_18012,N_16910,N_16341);
or U18013 (N_18013,N_17134,N_16768);
xor U18014 (N_18014,N_16772,N_16402);
xor U18015 (N_18015,N_16572,N_16933);
or U18016 (N_18016,N_17433,N_16295);
nand U18017 (N_18017,N_16514,N_17148);
xor U18018 (N_18018,N_17345,N_16419);
xor U18019 (N_18019,N_16525,N_16456);
or U18020 (N_18020,N_17097,N_17064);
or U18021 (N_18021,N_16628,N_16684);
and U18022 (N_18022,N_17221,N_16412);
nand U18023 (N_18023,N_16469,N_16652);
nand U18024 (N_18024,N_17391,N_16841);
and U18025 (N_18025,N_17319,N_16868);
nand U18026 (N_18026,N_16280,N_17236);
and U18027 (N_18027,N_16473,N_16523);
and U18028 (N_18028,N_17132,N_16731);
and U18029 (N_18029,N_16589,N_17353);
nor U18030 (N_18030,N_16761,N_16966);
xor U18031 (N_18031,N_17241,N_16931);
nor U18032 (N_18032,N_16457,N_17099);
nor U18033 (N_18033,N_17069,N_16631);
or U18034 (N_18034,N_16370,N_16755);
or U18035 (N_18035,N_16570,N_17461);
and U18036 (N_18036,N_16513,N_16643);
xnor U18037 (N_18037,N_16399,N_17010);
xor U18038 (N_18038,N_16603,N_16376);
nand U18039 (N_18039,N_16446,N_17038);
or U18040 (N_18040,N_17406,N_16935);
nand U18041 (N_18041,N_16607,N_17035);
nand U18042 (N_18042,N_16313,N_17473);
or U18043 (N_18043,N_17217,N_17363);
or U18044 (N_18044,N_16348,N_16332);
or U18045 (N_18045,N_17022,N_17179);
nand U18046 (N_18046,N_16445,N_16301);
nand U18047 (N_18047,N_17005,N_16420);
nand U18048 (N_18048,N_16720,N_16527);
or U18049 (N_18049,N_16801,N_17103);
and U18050 (N_18050,N_16677,N_16557);
xor U18051 (N_18051,N_16338,N_17057);
nand U18052 (N_18052,N_17133,N_16548);
nand U18053 (N_18053,N_17257,N_16377);
xor U18054 (N_18054,N_16906,N_16554);
nand U18055 (N_18055,N_17489,N_16908);
or U18056 (N_18056,N_16415,N_17201);
and U18057 (N_18057,N_16848,N_17152);
and U18058 (N_18058,N_17164,N_16568);
nand U18059 (N_18059,N_17456,N_17147);
nand U18060 (N_18060,N_16691,N_17376);
and U18061 (N_18061,N_16675,N_16994);
nor U18062 (N_18062,N_16869,N_16903);
or U18063 (N_18063,N_16475,N_16671);
and U18064 (N_18064,N_16318,N_16730);
or U18065 (N_18065,N_16739,N_17370);
nand U18066 (N_18066,N_17060,N_16878);
nor U18067 (N_18067,N_16716,N_17380);
and U18068 (N_18068,N_17306,N_17262);
nand U18069 (N_18069,N_16920,N_17481);
or U18070 (N_18070,N_16532,N_17090);
or U18071 (N_18071,N_17124,N_16705);
nand U18072 (N_18072,N_17239,N_16943);
nand U18073 (N_18073,N_16883,N_17434);
or U18074 (N_18074,N_16647,N_16654);
or U18075 (N_18075,N_17472,N_16770);
or U18076 (N_18076,N_16573,N_16442);
and U18077 (N_18077,N_16588,N_16300);
and U18078 (N_18078,N_17382,N_16854);
xnor U18079 (N_18079,N_16656,N_16797);
xnor U18080 (N_18080,N_17474,N_17324);
or U18081 (N_18081,N_16853,N_16879);
nor U18082 (N_18082,N_16750,N_17442);
and U18083 (N_18083,N_16627,N_17203);
nand U18084 (N_18084,N_16250,N_17276);
xnor U18085 (N_18085,N_16574,N_16811);
nor U18086 (N_18086,N_17355,N_16711);
nor U18087 (N_18087,N_16805,N_17496);
xnor U18088 (N_18088,N_16645,N_17040);
nand U18089 (N_18089,N_17468,N_16435);
and U18090 (N_18090,N_16696,N_17159);
nand U18091 (N_18091,N_16900,N_16981);
and U18092 (N_18092,N_16622,N_16725);
nor U18093 (N_18093,N_16549,N_17173);
nand U18094 (N_18094,N_17341,N_16814);
nand U18095 (N_18095,N_16937,N_17055);
xor U18096 (N_18096,N_17310,N_17278);
nand U18097 (N_18097,N_17390,N_16753);
nand U18098 (N_18098,N_17056,N_16453);
nand U18099 (N_18099,N_16558,N_17401);
xor U18100 (N_18100,N_16345,N_16746);
nand U18101 (N_18101,N_16793,N_16587);
nor U18102 (N_18102,N_16638,N_16423);
or U18103 (N_18103,N_16619,N_16693);
or U18104 (N_18104,N_16657,N_16757);
nor U18105 (N_18105,N_16951,N_17140);
and U18106 (N_18106,N_16324,N_16389);
and U18107 (N_18107,N_17197,N_16411);
and U18108 (N_18108,N_16540,N_16459);
or U18109 (N_18109,N_16434,N_17206);
xor U18110 (N_18110,N_16268,N_16334);
nor U18111 (N_18111,N_16821,N_16986);
xnor U18112 (N_18112,N_17448,N_16763);
nor U18113 (N_18113,N_16826,N_17144);
or U18114 (N_18114,N_16907,N_16396);
or U18115 (N_18115,N_16871,N_16884);
xnor U18116 (N_18116,N_16865,N_17312);
or U18117 (N_18117,N_16271,N_16546);
and U18118 (N_18118,N_16680,N_16646);
and U18119 (N_18119,N_16353,N_16993);
and U18120 (N_18120,N_17019,N_17268);
xor U18121 (N_18121,N_16686,N_16529);
xnor U18122 (N_18122,N_17340,N_17176);
nor U18123 (N_18123,N_16598,N_16887);
nand U18124 (N_18124,N_16695,N_17212);
or U18125 (N_18125,N_17267,N_17398);
and U18126 (N_18126,N_17126,N_16590);
nor U18127 (N_18127,N_17057,N_17230);
and U18128 (N_18128,N_16345,N_17132);
and U18129 (N_18129,N_16761,N_17221);
or U18130 (N_18130,N_16471,N_16833);
xnor U18131 (N_18131,N_16912,N_16961);
xnor U18132 (N_18132,N_16289,N_17329);
xnor U18133 (N_18133,N_17110,N_17296);
or U18134 (N_18134,N_16796,N_17349);
xor U18135 (N_18135,N_17266,N_17424);
nor U18136 (N_18136,N_16720,N_16925);
xnor U18137 (N_18137,N_16392,N_17207);
nor U18138 (N_18138,N_16426,N_17185);
and U18139 (N_18139,N_16932,N_17337);
or U18140 (N_18140,N_16307,N_17262);
nor U18141 (N_18141,N_17118,N_17399);
nor U18142 (N_18142,N_16459,N_16252);
and U18143 (N_18143,N_17292,N_16678);
or U18144 (N_18144,N_17059,N_16648);
nand U18145 (N_18145,N_16963,N_17154);
nor U18146 (N_18146,N_16833,N_16458);
nor U18147 (N_18147,N_16490,N_17028);
xnor U18148 (N_18148,N_17249,N_16296);
xnor U18149 (N_18149,N_17271,N_16458);
xor U18150 (N_18150,N_16331,N_16997);
or U18151 (N_18151,N_17040,N_17460);
nand U18152 (N_18152,N_16611,N_17277);
or U18153 (N_18153,N_16718,N_17162);
nand U18154 (N_18154,N_16659,N_16514);
or U18155 (N_18155,N_16528,N_16981);
and U18156 (N_18156,N_17229,N_16582);
xnor U18157 (N_18157,N_16755,N_17147);
xnor U18158 (N_18158,N_17082,N_16382);
and U18159 (N_18159,N_16859,N_17134);
and U18160 (N_18160,N_16403,N_17078);
and U18161 (N_18161,N_16389,N_17322);
xnor U18162 (N_18162,N_17211,N_16322);
nand U18163 (N_18163,N_16847,N_16762);
nor U18164 (N_18164,N_16427,N_16588);
and U18165 (N_18165,N_16980,N_17128);
and U18166 (N_18166,N_16980,N_17218);
or U18167 (N_18167,N_16451,N_16913);
and U18168 (N_18168,N_16672,N_16396);
and U18169 (N_18169,N_17288,N_17204);
nand U18170 (N_18170,N_16452,N_17337);
nand U18171 (N_18171,N_16880,N_16750);
nor U18172 (N_18172,N_17155,N_17259);
and U18173 (N_18173,N_16693,N_16814);
or U18174 (N_18174,N_16902,N_17481);
and U18175 (N_18175,N_17280,N_17074);
nand U18176 (N_18176,N_16780,N_17463);
xnor U18177 (N_18177,N_16535,N_16347);
or U18178 (N_18178,N_16640,N_16845);
xnor U18179 (N_18179,N_16643,N_16767);
nand U18180 (N_18180,N_16704,N_17451);
nand U18181 (N_18181,N_17401,N_16761);
nor U18182 (N_18182,N_17082,N_17172);
or U18183 (N_18183,N_17268,N_17246);
nor U18184 (N_18184,N_16557,N_17180);
nand U18185 (N_18185,N_17211,N_16344);
or U18186 (N_18186,N_17455,N_17186);
nand U18187 (N_18187,N_17380,N_16440);
nand U18188 (N_18188,N_16829,N_16574);
nor U18189 (N_18189,N_16806,N_17041);
nor U18190 (N_18190,N_16789,N_17355);
nand U18191 (N_18191,N_16463,N_16439);
or U18192 (N_18192,N_17132,N_16601);
nor U18193 (N_18193,N_17133,N_17194);
nor U18194 (N_18194,N_16553,N_17233);
and U18195 (N_18195,N_16518,N_17391);
nor U18196 (N_18196,N_16655,N_16924);
or U18197 (N_18197,N_17325,N_17451);
nand U18198 (N_18198,N_17377,N_17135);
nand U18199 (N_18199,N_17172,N_16425);
xnor U18200 (N_18200,N_17419,N_16936);
nand U18201 (N_18201,N_16764,N_16460);
nand U18202 (N_18202,N_16993,N_17310);
nand U18203 (N_18203,N_16596,N_17447);
xnor U18204 (N_18204,N_16276,N_17072);
nor U18205 (N_18205,N_16278,N_16602);
and U18206 (N_18206,N_17420,N_17025);
nor U18207 (N_18207,N_16425,N_16498);
xor U18208 (N_18208,N_16903,N_16402);
and U18209 (N_18209,N_17339,N_17465);
nor U18210 (N_18210,N_16455,N_16321);
nor U18211 (N_18211,N_17018,N_17146);
nand U18212 (N_18212,N_16706,N_17464);
nor U18213 (N_18213,N_16831,N_16383);
or U18214 (N_18214,N_17468,N_16317);
and U18215 (N_18215,N_16870,N_16926);
or U18216 (N_18216,N_17017,N_16448);
and U18217 (N_18217,N_17168,N_17405);
xnor U18218 (N_18218,N_16818,N_16733);
nand U18219 (N_18219,N_16773,N_17037);
nor U18220 (N_18220,N_17180,N_17067);
nor U18221 (N_18221,N_17177,N_17492);
and U18222 (N_18222,N_16737,N_16883);
nor U18223 (N_18223,N_16338,N_16497);
and U18224 (N_18224,N_17241,N_16669);
nand U18225 (N_18225,N_17058,N_16484);
and U18226 (N_18226,N_16898,N_17469);
nor U18227 (N_18227,N_16873,N_16634);
nand U18228 (N_18228,N_16615,N_16492);
nor U18229 (N_18229,N_16961,N_16989);
and U18230 (N_18230,N_17394,N_16723);
or U18231 (N_18231,N_16534,N_16770);
nor U18232 (N_18232,N_16869,N_17455);
nor U18233 (N_18233,N_16911,N_16319);
and U18234 (N_18234,N_16824,N_16697);
nand U18235 (N_18235,N_17161,N_16533);
xor U18236 (N_18236,N_16813,N_17049);
or U18237 (N_18237,N_17119,N_16780);
xor U18238 (N_18238,N_17031,N_16282);
nand U18239 (N_18239,N_16662,N_16862);
xor U18240 (N_18240,N_17004,N_17482);
or U18241 (N_18241,N_16995,N_16333);
xnor U18242 (N_18242,N_16738,N_16594);
xnor U18243 (N_18243,N_16902,N_17039);
nor U18244 (N_18244,N_17159,N_17120);
or U18245 (N_18245,N_16937,N_17355);
or U18246 (N_18246,N_16283,N_16392);
nand U18247 (N_18247,N_17478,N_17333);
or U18248 (N_18248,N_16383,N_16469);
or U18249 (N_18249,N_17009,N_16269);
nor U18250 (N_18250,N_16411,N_16998);
nor U18251 (N_18251,N_16904,N_17025);
and U18252 (N_18252,N_16328,N_16268);
or U18253 (N_18253,N_16768,N_16992);
or U18254 (N_18254,N_17392,N_16925);
xnor U18255 (N_18255,N_16628,N_16984);
and U18256 (N_18256,N_16520,N_17186);
and U18257 (N_18257,N_16543,N_16309);
xnor U18258 (N_18258,N_16263,N_17483);
or U18259 (N_18259,N_16326,N_16566);
or U18260 (N_18260,N_16982,N_17485);
or U18261 (N_18261,N_17365,N_16467);
or U18262 (N_18262,N_16824,N_16999);
and U18263 (N_18263,N_16258,N_16461);
or U18264 (N_18264,N_16547,N_16457);
nand U18265 (N_18265,N_16674,N_16694);
and U18266 (N_18266,N_16580,N_17302);
or U18267 (N_18267,N_16358,N_16862);
nand U18268 (N_18268,N_16749,N_16875);
nand U18269 (N_18269,N_16747,N_16571);
and U18270 (N_18270,N_17244,N_16648);
nand U18271 (N_18271,N_17337,N_16532);
or U18272 (N_18272,N_16962,N_16482);
or U18273 (N_18273,N_17008,N_17337);
nor U18274 (N_18274,N_17377,N_16441);
or U18275 (N_18275,N_16642,N_16278);
nor U18276 (N_18276,N_16370,N_16598);
xor U18277 (N_18277,N_17087,N_16395);
or U18278 (N_18278,N_16323,N_17274);
nand U18279 (N_18279,N_17155,N_16646);
nor U18280 (N_18280,N_16823,N_16464);
or U18281 (N_18281,N_17166,N_16471);
xnor U18282 (N_18282,N_17499,N_16798);
xor U18283 (N_18283,N_16667,N_17439);
nor U18284 (N_18284,N_16492,N_16992);
nor U18285 (N_18285,N_16898,N_17102);
xnor U18286 (N_18286,N_16820,N_17116);
nand U18287 (N_18287,N_17022,N_17261);
nor U18288 (N_18288,N_16759,N_17065);
xnor U18289 (N_18289,N_16829,N_16986);
nor U18290 (N_18290,N_17453,N_16494);
xnor U18291 (N_18291,N_16699,N_16975);
or U18292 (N_18292,N_16851,N_16552);
and U18293 (N_18293,N_17239,N_16386);
xor U18294 (N_18294,N_16521,N_16293);
and U18295 (N_18295,N_16712,N_17429);
nand U18296 (N_18296,N_16595,N_16870);
nand U18297 (N_18297,N_17463,N_16562);
xnor U18298 (N_18298,N_17447,N_17244);
or U18299 (N_18299,N_16695,N_17033);
nor U18300 (N_18300,N_17027,N_17130);
nand U18301 (N_18301,N_17058,N_16846);
or U18302 (N_18302,N_16785,N_16282);
or U18303 (N_18303,N_16565,N_16589);
nand U18304 (N_18304,N_16965,N_16910);
xor U18305 (N_18305,N_17177,N_16441);
nand U18306 (N_18306,N_16566,N_17050);
nor U18307 (N_18307,N_16394,N_16597);
or U18308 (N_18308,N_16642,N_17313);
xnor U18309 (N_18309,N_16538,N_16882);
or U18310 (N_18310,N_17201,N_17269);
nor U18311 (N_18311,N_16927,N_16809);
or U18312 (N_18312,N_16934,N_17236);
or U18313 (N_18313,N_17024,N_16791);
nand U18314 (N_18314,N_17310,N_16894);
nand U18315 (N_18315,N_17142,N_17373);
or U18316 (N_18316,N_16878,N_17138);
or U18317 (N_18317,N_17445,N_16756);
or U18318 (N_18318,N_17025,N_16619);
nand U18319 (N_18319,N_16872,N_16548);
nand U18320 (N_18320,N_17222,N_17320);
xnor U18321 (N_18321,N_16883,N_17377);
nand U18322 (N_18322,N_16587,N_16377);
and U18323 (N_18323,N_16519,N_16323);
xnor U18324 (N_18324,N_17410,N_16477);
nand U18325 (N_18325,N_17378,N_17197);
and U18326 (N_18326,N_16463,N_16865);
xnor U18327 (N_18327,N_16558,N_17405);
xnor U18328 (N_18328,N_16518,N_16477);
or U18329 (N_18329,N_16598,N_17287);
xnor U18330 (N_18330,N_17319,N_17447);
or U18331 (N_18331,N_17111,N_17363);
xnor U18332 (N_18332,N_17447,N_16647);
and U18333 (N_18333,N_16978,N_16801);
or U18334 (N_18334,N_16689,N_16688);
xnor U18335 (N_18335,N_17010,N_16915);
or U18336 (N_18336,N_16251,N_17036);
and U18337 (N_18337,N_16889,N_16502);
or U18338 (N_18338,N_16283,N_17153);
xor U18339 (N_18339,N_16624,N_17087);
xnor U18340 (N_18340,N_16887,N_16611);
and U18341 (N_18341,N_17233,N_16496);
or U18342 (N_18342,N_16482,N_17129);
nor U18343 (N_18343,N_16620,N_16738);
or U18344 (N_18344,N_16351,N_17164);
and U18345 (N_18345,N_16442,N_17486);
and U18346 (N_18346,N_16347,N_17493);
xnor U18347 (N_18347,N_17056,N_17136);
nand U18348 (N_18348,N_17080,N_17376);
or U18349 (N_18349,N_16258,N_16748);
xnor U18350 (N_18350,N_16475,N_16371);
or U18351 (N_18351,N_17085,N_16342);
nand U18352 (N_18352,N_16673,N_16750);
nor U18353 (N_18353,N_17289,N_16692);
or U18354 (N_18354,N_17216,N_16993);
and U18355 (N_18355,N_17364,N_16433);
nand U18356 (N_18356,N_16739,N_16790);
or U18357 (N_18357,N_17185,N_17337);
nand U18358 (N_18358,N_16714,N_16776);
or U18359 (N_18359,N_16390,N_16295);
or U18360 (N_18360,N_16529,N_16399);
xnor U18361 (N_18361,N_16284,N_16778);
xor U18362 (N_18362,N_16456,N_17128);
nor U18363 (N_18363,N_16569,N_16882);
or U18364 (N_18364,N_16996,N_17399);
nand U18365 (N_18365,N_16975,N_17358);
nand U18366 (N_18366,N_17439,N_16469);
xnor U18367 (N_18367,N_16408,N_16568);
nand U18368 (N_18368,N_17197,N_17250);
xnor U18369 (N_18369,N_16826,N_16463);
nand U18370 (N_18370,N_16947,N_16870);
and U18371 (N_18371,N_16307,N_16326);
and U18372 (N_18372,N_16974,N_16715);
and U18373 (N_18373,N_16659,N_17327);
nor U18374 (N_18374,N_16449,N_16978);
nand U18375 (N_18375,N_16740,N_16920);
nor U18376 (N_18376,N_16783,N_16922);
and U18377 (N_18377,N_16393,N_16961);
and U18378 (N_18378,N_16833,N_16425);
nor U18379 (N_18379,N_16718,N_16579);
and U18380 (N_18380,N_17085,N_16767);
xor U18381 (N_18381,N_16488,N_17197);
xnor U18382 (N_18382,N_17431,N_17465);
and U18383 (N_18383,N_16368,N_17157);
nor U18384 (N_18384,N_17064,N_16549);
nor U18385 (N_18385,N_16646,N_17285);
xnor U18386 (N_18386,N_16350,N_17323);
or U18387 (N_18387,N_17269,N_16712);
nor U18388 (N_18388,N_17286,N_16295);
nor U18389 (N_18389,N_17395,N_17322);
and U18390 (N_18390,N_17047,N_17250);
or U18391 (N_18391,N_17290,N_17413);
or U18392 (N_18392,N_17172,N_16506);
and U18393 (N_18393,N_16668,N_16750);
and U18394 (N_18394,N_16542,N_16399);
nand U18395 (N_18395,N_16506,N_16422);
and U18396 (N_18396,N_17417,N_16625);
xor U18397 (N_18397,N_16795,N_17169);
nor U18398 (N_18398,N_17395,N_17411);
xor U18399 (N_18399,N_17297,N_16451);
and U18400 (N_18400,N_17293,N_16873);
xnor U18401 (N_18401,N_17204,N_17060);
or U18402 (N_18402,N_17129,N_17051);
or U18403 (N_18403,N_17146,N_17432);
or U18404 (N_18404,N_16576,N_16824);
nor U18405 (N_18405,N_17077,N_16596);
xnor U18406 (N_18406,N_17397,N_16567);
and U18407 (N_18407,N_16765,N_16396);
and U18408 (N_18408,N_16787,N_17032);
nor U18409 (N_18409,N_17103,N_17107);
xor U18410 (N_18410,N_16383,N_16558);
or U18411 (N_18411,N_17074,N_17497);
and U18412 (N_18412,N_17202,N_16761);
and U18413 (N_18413,N_17340,N_16962);
nand U18414 (N_18414,N_16467,N_17263);
or U18415 (N_18415,N_16310,N_17367);
and U18416 (N_18416,N_16381,N_17008);
nand U18417 (N_18417,N_17436,N_16763);
xnor U18418 (N_18418,N_17152,N_16599);
xnor U18419 (N_18419,N_16756,N_17100);
xor U18420 (N_18420,N_17234,N_16479);
nand U18421 (N_18421,N_16567,N_16480);
nand U18422 (N_18422,N_16984,N_17326);
and U18423 (N_18423,N_17123,N_16767);
xor U18424 (N_18424,N_16803,N_16743);
nand U18425 (N_18425,N_17474,N_16531);
nand U18426 (N_18426,N_16725,N_16657);
and U18427 (N_18427,N_17150,N_17069);
nand U18428 (N_18428,N_16578,N_16705);
or U18429 (N_18429,N_16376,N_17325);
nand U18430 (N_18430,N_16420,N_16450);
nand U18431 (N_18431,N_17128,N_17213);
and U18432 (N_18432,N_16346,N_17344);
nor U18433 (N_18433,N_16253,N_16994);
or U18434 (N_18434,N_17456,N_16972);
xnor U18435 (N_18435,N_16932,N_17154);
and U18436 (N_18436,N_17483,N_17499);
or U18437 (N_18437,N_17181,N_16843);
and U18438 (N_18438,N_16511,N_16500);
nand U18439 (N_18439,N_16528,N_16980);
xor U18440 (N_18440,N_16707,N_16850);
nor U18441 (N_18441,N_17486,N_16359);
or U18442 (N_18442,N_16336,N_16659);
and U18443 (N_18443,N_16494,N_16971);
xor U18444 (N_18444,N_17305,N_16825);
nor U18445 (N_18445,N_16761,N_16583);
nor U18446 (N_18446,N_16645,N_17080);
xnor U18447 (N_18447,N_16948,N_17321);
and U18448 (N_18448,N_16933,N_17135);
xor U18449 (N_18449,N_17012,N_16833);
xnor U18450 (N_18450,N_16836,N_16355);
nand U18451 (N_18451,N_17084,N_16791);
nor U18452 (N_18452,N_16756,N_17387);
or U18453 (N_18453,N_17230,N_16297);
xnor U18454 (N_18454,N_17398,N_16779);
or U18455 (N_18455,N_16379,N_16355);
xor U18456 (N_18456,N_16764,N_17214);
xor U18457 (N_18457,N_16545,N_16363);
xor U18458 (N_18458,N_17263,N_17323);
and U18459 (N_18459,N_17194,N_17365);
and U18460 (N_18460,N_17405,N_17273);
xor U18461 (N_18461,N_17212,N_17024);
xor U18462 (N_18462,N_16718,N_17365);
nand U18463 (N_18463,N_16495,N_16940);
xor U18464 (N_18464,N_17189,N_16383);
xor U18465 (N_18465,N_17029,N_16617);
xor U18466 (N_18466,N_16828,N_16918);
xnor U18467 (N_18467,N_16453,N_16376);
xnor U18468 (N_18468,N_16832,N_16889);
xor U18469 (N_18469,N_17354,N_16500);
or U18470 (N_18470,N_16282,N_16519);
and U18471 (N_18471,N_17267,N_16446);
or U18472 (N_18472,N_16370,N_16771);
and U18473 (N_18473,N_16925,N_16390);
xor U18474 (N_18474,N_16984,N_16291);
or U18475 (N_18475,N_17060,N_16767);
nand U18476 (N_18476,N_16921,N_17404);
or U18477 (N_18477,N_17092,N_16511);
nand U18478 (N_18478,N_17096,N_17145);
nand U18479 (N_18479,N_17418,N_16991);
and U18480 (N_18480,N_16571,N_17004);
xor U18481 (N_18481,N_17381,N_16952);
xor U18482 (N_18482,N_16488,N_16482);
nand U18483 (N_18483,N_17306,N_16347);
or U18484 (N_18484,N_16576,N_16428);
or U18485 (N_18485,N_17111,N_17172);
nand U18486 (N_18486,N_17101,N_16445);
or U18487 (N_18487,N_17207,N_16872);
nor U18488 (N_18488,N_17373,N_16990);
and U18489 (N_18489,N_16403,N_16335);
nor U18490 (N_18490,N_16261,N_17270);
or U18491 (N_18491,N_16713,N_17079);
or U18492 (N_18492,N_16892,N_17477);
nand U18493 (N_18493,N_17027,N_17305);
xnor U18494 (N_18494,N_17144,N_16268);
nor U18495 (N_18495,N_16928,N_16426);
or U18496 (N_18496,N_17344,N_17187);
xnor U18497 (N_18497,N_17112,N_17451);
or U18498 (N_18498,N_16323,N_17376);
xnor U18499 (N_18499,N_16264,N_16675);
xor U18500 (N_18500,N_17042,N_16852);
nand U18501 (N_18501,N_16408,N_16555);
and U18502 (N_18502,N_16313,N_17320);
xnor U18503 (N_18503,N_16295,N_16862);
nand U18504 (N_18504,N_16823,N_16653);
nor U18505 (N_18505,N_16965,N_16483);
nand U18506 (N_18506,N_16282,N_16629);
or U18507 (N_18507,N_17302,N_16595);
nand U18508 (N_18508,N_16868,N_16738);
or U18509 (N_18509,N_16990,N_16782);
and U18510 (N_18510,N_16487,N_17093);
xor U18511 (N_18511,N_16294,N_16728);
nand U18512 (N_18512,N_16878,N_17053);
or U18513 (N_18513,N_16986,N_17151);
and U18514 (N_18514,N_17266,N_16392);
nor U18515 (N_18515,N_16608,N_17118);
or U18516 (N_18516,N_16333,N_16933);
or U18517 (N_18517,N_17039,N_16684);
or U18518 (N_18518,N_16999,N_16716);
nor U18519 (N_18519,N_16620,N_17189);
nand U18520 (N_18520,N_16541,N_17101);
nor U18521 (N_18521,N_17324,N_17349);
nor U18522 (N_18522,N_16407,N_17016);
or U18523 (N_18523,N_16728,N_16458);
xnor U18524 (N_18524,N_17007,N_17073);
or U18525 (N_18525,N_17421,N_16881);
and U18526 (N_18526,N_16382,N_16888);
nor U18527 (N_18527,N_16320,N_16469);
nor U18528 (N_18528,N_16373,N_16725);
or U18529 (N_18529,N_17225,N_16884);
nor U18530 (N_18530,N_16603,N_16695);
or U18531 (N_18531,N_16856,N_17419);
or U18532 (N_18532,N_16892,N_16539);
or U18533 (N_18533,N_16411,N_16321);
or U18534 (N_18534,N_16472,N_17204);
nand U18535 (N_18535,N_17371,N_16270);
and U18536 (N_18536,N_16504,N_17441);
nand U18537 (N_18537,N_17176,N_17386);
or U18538 (N_18538,N_16655,N_16415);
xor U18539 (N_18539,N_16253,N_16573);
nor U18540 (N_18540,N_17047,N_16863);
or U18541 (N_18541,N_16827,N_16667);
nand U18542 (N_18542,N_16414,N_17434);
and U18543 (N_18543,N_17429,N_16787);
nor U18544 (N_18544,N_17078,N_16652);
or U18545 (N_18545,N_17107,N_17077);
nor U18546 (N_18546,N_17121,N_17310);
nand U18547 (N_18547,N_17351,N_16647);
and U18548 (N_18548,N_16303,N_17045);
nor U18549 (N_18549,N_16779,N_17249);
and U18550 (N_18550,N_17497,N_16626);
or U18551 (N_18551,N_16444,N_17379);
nor U18552 (N_18552,N_17468,N_17423);
nor U18553 (N_18553,N_17219,N_17173);
or U18554 (N_18554,N_16700,N_17350);
xor U18555 (N_18555,N_16570,N_17344);
and U18556 (N_18556,N_16369,N_16842);
nand U18557 (N_18557,N_17330,N_16489);
and U18558 (N_18558,N_16460,N_16607);
and U18559 (N_18559,N_17376,N_16390);
or U18560 (N_18560,N_16263,N_17123);
xnor U18561 (N_18561,N_17441,N_16802);
and U18562 (N_18562,N_16641,N_17051);
nor U18563 (N_18563,N_16707,N_17324);
and U18564 (N_18564,N_17295,N_17310);
nand U18565 (N_18565,N_16542,N_16712);
or U18566 (N_18566,N_17266,N_17182);
nor U18567 (N_18567,N_16512,N_16780);
xor U18568 (N_18568,N_16912,N_16361);
nand U18569 (N_18569,N_16783,N_16666);
and U18570 (N_18570,N_16708,N_16621);
nor U18571 (N_18571,N_16995,N_16352);
or U18572 (N_18572,N_16645,N_16974);
and U18573 (N_18573,N_17453,N_16823);
or U18574 (N_18574,N_16548,N_17454);
nand U18575 (N_18575,N_16764,N_16847);
or U18576 (N_18576,N_16718,N_16536);
nor U18577 (N_18577,N_16605,N_16403);
nand U18578 (N_18578,N_17009,N_17194);
nand U18579 (N_18579,N_16762,N_17262);
or U18580 (N_18580,N_16849,N_16373);
and U18581 (N_18581,N_16785,N_17343);
or U18582 (N_18582,N_16834,N_16351);
nor U18583 (N_18583,N_16639,N_17222);
xnor U18584 (N_18584,N_17422,N_16723);
or U18585 (N_18585,N_17229,N_16751);
or U18586 (N_18586,N_16998,N_17446);
and U18587 (N_18587,N_16891,N_17330);
nor U18588 (N_18588,N_16851,N_16437);
or U18589 (N_18589,N_17245,N_17380);
nand U18590 (N_18590,N_16764,N_16965);
nand U18591 (N_18591,N_16570,N_16829);
nor U18592 (N_18592,N_16999,N_17481);
and U18593 (N_18593,N_16674,N_16614);
or U18594 (N_18594,N_16781,N_16620);
or U18595 (N_18595,N_16372,N_16657);
and U18596 (N_18596,N_17022,N_17070);
nand U18597 (N_18597,N_17306,N_17373);
or U18598 (N_18598,N_17217,N_17438);
xnor U18599 (N_18599,N_16304,N_17448);
or U18600 (N_18600,N_16652,N_17243);
xor U18601 (N_18601,N_16951,N_17011);
xnor U18602 (N_18602,N_17425,N_16773);
nor U18603 (N_18603,N_16893,N_17050);
nand U18604 (N_18604,N_16517,N_17464);
nand U18605 (N_18605,N_17472,N_16836);
nor U18606 (N_18606,N_17311,N_16403);
and U18607 (N_18607,N_17361,N_17093);
and U18608 (N_18608,N_16400,N_17332);
xnor U18609 (N_18609,N_16693,N_17075);
xor U18610 (N_18610,N_16454,N_16818);
nor U18611 (N_18611,N_17001,N_16827);
nor U18612 (N_18612,N_17219,N_16811);
and U18613 (N_18613,N_17255,N_16911);
xnor U18614 (N_18614,N_16598,N_16708);
or U18615 (N_18615,N_17210,N_16274);
nor U18616 (N_18616,N_17164,N_16303);
nor U18617 (N_18617,N_16724,N_17038);
or U18618 (N_18618,N_17243,N_16836);
nor U18619 (N_18619,N_17377,N_16342);
or U18620 (N_18620,N_16474,N_17431);
or U18621 (N_18621,N_16864,N_16991);
and U18622 (N_18622,N_17291,N_17231);
or U18623 (N_18623,N_16942,N_17116);
xnor U18624 (N_18624,N_17374,N_17128);
nand U18625 (N_18625,N_16923,N_17125);
nor U18626 (N_18626,N_16755,N_16613);
and U18627 (N_18627,N_17209,N_16445);
nor U18628 (N_18628,N_16752,N_16567);
xnor U18629 (N_18629,N_16989,N_16333);
xnor U18630 (N_18630,N_17207,N_17136);
xor U18631 (N_18631,N_17421,N_16338);
nor U18632 (N_18632,N_16942,N_16945);
nor U18633 (N_18633,N_16720,N_16735);
nor U18634 (N_18634,N_17290,N_17111);
xnor U18635 (N_18635,N_16413,N_16429);
and U18636 (N_18636,N_17438,N_16635);
and U18637 (N_18637,N_16752,N_16258);
nor U18638 (N_18638,N_16873,N_16595);
and U18639 (N_18639,N_16591,N_17111);
or U18640 (N_18640,N_17224,N_17279);
and U18641 (N_18641,N_17497,N_16693);
and U18642 (N_18642,N_16406,N_16463);
nand U18643 (N_18643,N_16614,N_16749);
or U18644 (N_18644,N_16554,N_17094);
nor U18645 (N_18645,N_17281,N_17041);
nor U18646 (N_18646,N_17133,N_17132);
xor U18647 (N_18647,N_17033,N_16937);
or U18648 (N_18648,N_16502,N_16419);
nor U18649 (N_18649,N_16802,N_17496);
nand U18650 (N_18650,N_16770,N_16998);
xor U18651 (N_18651,N_17025,N_16473);
xor U18652 (N_18652,N_16729,N_16521);
or U18653 (N_18653,N_17245,N_17447);
xor U18654 (N_18654,N_17481,N_17229);
nor U18655 (N_18655,N_16436,N_17237);
or U18656 (N_18656,N_16889,N_16885);
and U18657 (N_18657,N_16454,N_16788);
and U18658 (N_18658,N_17454,N_16851);
or U18659 (N_18659,N_17237,N_17242);
or U18660 (N_18660,N_16361,N_16362);
and U18661 (N_18661,N_17311,N_16445);
nor U18662 (N_18662,N_17023,N_17236);
xor U18663 (N_18663,N_16632,N_17358);
or U18664 (N_18664,N_16525,N_16549);
and U18665 (N_18665,N_16358,N_17100);
nand U18666 (N_18666,N_17168,N_16316);
nand U18667 (N_18667,N_17287,N_16298);
or U18668 (N_18668,N_17296,N_17486);
nand U18669 (N_18669,N_16337,N_17229);
nor U18670 (N_18670,N_16409,N_16581);
nor U18671 (N_18671,N_16470,N_16688);
and U18672 (N_18672,N_16563,N_16694);
nand U18673 (N_18673,N_16292,N_16548);
nor U18674 (N_18674,N_16779,N_16510);
or U18675 (N_18675,N_17239,N_16272);
or U18676 (N_18676,N_17027,N_17128);
and U18677 (N_18677,N_17084,N_16481);
or U18678 (N_18678,N_16417,N_16324);
xor U18679 (N_18679,N_17365,N_17097);
nor U18680 (N_18680,N_16434,N_16536);
nand U18681 (N_18681,N_16914,N_16928);
xor U18682 (N_18682,N_16318,N_16982);
nor U18683 (N_18683,N_16540,N_16864);
and U18684 (N_18684,N_16824,N_16413);
and U18685 (N_18685,N_16410,N_16658);
and U18686 (N_18686,N_16637,N_17312);
nand U18687 (N_18687,N_16315,N_16774);
nand U18688 (N_18688,N_16876,N_16753);
and U18689 (N_18689,N_16427,N_17051);
nand U18690 (N_18690,N_16879,N_16307);
nor U18691 (N_18691,N_17358,N_17084);
and U18692 (N_18692,N_17476,N_17463);
xor U18693 (N_18693,N_17247,N_16658);
nor U18694 (N_18694,N_16262,N_17113);
nor U18695 (N_18695,N_17224,N_17452);
and U18696 (N_18696,N_17017,N_16656);
and U18697 (N_18697,N_16301,N_17337);
or U18698 (N_18698,N_16501,N_16413);
and U18699 (N_18699,N_16410,N_17248);
or U18700 (N_18700,N_17291,N_17107);
or U18701 (N_18701,N_16710,N_16333);
nand U18702 (N_18702,N_16320,N_16282);
nor U18703 (N_18703,N_16711,N_17393);
xnor U18704 (N_18704,N_16692,N_16859);
and U18705 (N_18705,N_16641,N_16806);
or U18706 (N_18706,N_17433,N_16911);
xor U18707 (N_18707,N_17078,N_16331);
nand U18708 (N_18708,N_16336,N_17436);
and U18709 (N_18709,N_17287,N_17272);
xor U18710 (N_18710,N_17092,N_16878);
or U18711 (N_18711,N_16842,N_16990);
nand U18712 (N_18712,N_16621,N_16256);
or U18713 (N_18713,N_16474,N_16761);
and U18714 (N_18714,N_17195,N_16390);
and U18715 (N_18715,N_16359,N_16754);
xor U18716 (N_18716,N_17443,N_16857);
nor U18717 (N_18717,N_16596,N_16389);
nor U18718 (N_18718,N_17333,N_16736);
xor U18719 (N_18719,N_16388,N_17423);
or U18720 (N_18720,N_16638,N_16753);
and U18721 (N_18721,N_16315,N_16412);
nor U18722 (N_18722,N_16384,N_16511);
or U18723 (N_18723,N_17209,N_17250);
nand U18724 (N_18724,N_17256,N_16767);
nand U18725 (N_18725,N_17156,N_16623);
or U18726 (N_18726,N_16556,N_16574);
and U18727 (N_18727,N_16676,N_16802);
xor U18728 (N_18728,N_17131,N_16691);
nand U18729 (N_18729,N_16361,N_16906);
and U18730 (N_18730,N_16706,N_17414);
xnor U18731 (N_18731,N_17096,N_16958);
xor U18732 (N_18732,N_16864,N_17054);
or U18733 (N_18733,N_16844,N_16325);
or U18734 (N_18734,N_16684,N_16542);
nor U18735 (N_18735,N_17464,N_16347);
xnor U18736 (N_18736,N_17439,N_16525);
or U18737 (N_18737,N_16771,N_17124);
nand U18738 (N_18738,N_17225,N_17070);
nor U18739 (N_18739,N_16560,N_17495);
nand U18740 (N_18740,N_17341,N_17265);
xnor U18741 (N_18741,N_17220,N_16560);
and U18742 (N_18742,N_17459,N_16926);
nand U18743 (N_18743,N_17479,N_17152);
xor U18744 (N_18744,N_17125,N_16573);
or U18745 (N_18745,N_16405,N_16455);
or U18746 (N_18746,N_17183,N_16478);
and U18747 (N_18747,N_17223,N_16503);
xor U18748 (N_18748,N_17435,N_17009);
nor U18749 (N_18749,N_16562,N_17405);
and U18750 (N_18750,N_17691,N_18103);
nand U18751 (N_18751,N_17989,N_17692);
or U18752 (N_18752,N_17811,N_18070);
nand U18753 (N_18753,N_18465,N_17815);
or U18754 (N_18754,N_18629,N_18019);
nor U18755 (N_18755,N_17714,N_18570);
nand U18756 (N_18756,N_18273,N_18327);
nor U18757 (N_18757,N_17615,N_17818);
or U18758 (N_18758,N_18374,N_18049);
nand U18759 (N_18759,N_18315,N_17908);
xnor U18760 (N_18760,N_17630,N_18297);
xnor U18761 (N_18761,N_17530,N_17761);
and U18762 (N_18762,N_17794,N_17546);
xor U18763 (N_18763,N_18602,N_18302);
and U18764 (N_18764,N_17995,N_18488);
and U18765 (N_18765,N_18169,N_18742);
or U18766 (N_18766,N_17817,N_17913);
and U18767 (N_18767,N_18523,N_17592);
or U18768 (N_18768,N_18368,N_17551);
and U18769 (N_18769,N_18216,N_18240);
nor U18770 (N_18770,N_18094,N_18402);
nor U18771 (N_18771,N_18228,N_17788);
xor U18772 (N_18772,N_18609,N_17897);
and U18773 (N_18773,N_17735,N_18125);
or U18774 (N_18774,N_17825,N_17736);
nand U18775 (N_18775,N_17965,N_17520);
nor U18776 (N_18776,N_17614,N_18028);
and U18777 (N_18777,N_18110,N_17547);
or U18778 (N_18778,N_18238,N_18280);
xnor U18779 (N_18779,N_17977,N_17536);
nor U18780 (N_18780,N_17524,N_18007);
nand U18781 (N_18781,N_18058,N_18385);
or U18782 (N_18782,N_17964,N_18642);
or U18783 (N_18783,N_18362,N_18226);
and U18784 (N_18784,N_18383,N_18243);
and U18785 (N_18785,N_18709,N_17993);
nand U18786 (N_18786,N_18355,N_18571);
or U18787 (N_18787,N_18391,N_18396);
nand U18788 (N_18788,N_18694,N_18406);
nor U18789 (N_18789,N_18587,N_17729);
or U18790 (N_18790,N_18156,N_17888);
xnor U18791 (N_18791,N_18418,N_17588);
nand U18792 (N_18792,N_18444,N_17838);
xnor U18793 (N_18793,N_18260,N_17983);
nor U18794 (N_18794,N_18463,N_18670);
nand U18795 (N_18795,N_17875,N_17997);
xnor U18796 (N_18796,N_17861,N_18469);
xnor U18797 (N_18797,N_17512,N_17747);
nand U18798 (N_18798,N_18213,N_18295);
xnor U18799 (N_18799,N_18697,N_17601);
nor U18800 (N_18800,N_18118,N_17722);
and U18801 (N_18801,N_17912,N_18598);
nand U18802 (N_18802,N_18707,N_17771);
and U18803 (N_18803,N_17947,N_18056);
nor U18804 (N_18804,N_17962,N_18230);
or U18805 (N_18805,N_18205,N_18721);
nor U18806 (N_18806,N_17593,N_17883);
xor U18807 (N_18807,N_17847,N_18036);
nor U18808 (N_18808,N_18664,N_17523);
or U18809 (N_18809,N_17981,N_17905);
nand U18810 (N_18810,N_18274,N_18290);
xor U18811 (N_18811,N_18384,N_18453);
or U18812 (N_18812,N_18161,N_18566);
and U18813 (N_18813,N_18720,N_18660);
nand U18814 (N_18814,N_18092,N_18533);
nor U18815 (N_18815,N_18364,N_18509);
or U18816 (N_18816,N_17662,N_17585);
and U18817 (N_18817,N_18320,N_17621);
xor U18818 (N_18818,N_18404,N_17743);
and U18819 (N_18819,N_18155,N_17949);
nand U18820 (N_18820,N_17954,N_18063);
nor U18821 (N_18821,N_17996,N_17918);
or U18822 (N_18822,N_17707,N_17541);
xnor U18823 (N_18823,N_18180,N_18378);
or U18824 (N_18824,N_17784,N_18628);
and U18825 (N_18825,N_17974,N_18310);
nand U18826 (N_18826,N_17539,N_18481);
nand U18827 (N_18827,N_17748,N_18151);
or U18828 (N_18828,N_17782,N_18003);
and U18829 (N_18829,N_18080,N_18505);
xor U18830 (N_18830,N_18654,N_18254);
xor U18831 (N_18831,N_18365,N_18442);
xor U18832 (N_18832,N_18564,N_18076);
or U18833 (N_18833,N_18042,N_17644);
xor U18834 (N_18834,N_17865,N_17936);
nor U18835 (N_18835,N_18666,N_17646);
nand U18836 (N_18836,N_17935,N_18543);
xnor U18837 (N_18837,N_18485,N_18329);
and U18838 (N_18838,N_17766,N_18634);
and U18839 (N_18839,N_18127,N_18207);
nor U18840 (N_18840,N_17940,N_18575);
nand U18841 (N_18841,N_17559,N_17705);
nand U18842 (N_18842,N_18136,N_18287);
nand U18843 (N_18843,N_18426,N_18291);
nor U18844 (N_18844,N_18684,N_17719);
xor U18845 (N_18845,N_18328,N_18342);
or U18846 (N_18846,N_18500,N_18112);
and U18847 (N_18847,N_18168,N_17603);
and U18848 (N_18848,N_18578,N_17677);
nand U18849 (N_18849,N_17952,N_18589);
and U18850 (N_18850,N_18229,N_17851);
or U18851 (N_18851,N_18296,N_18746);
xor U18852 (N_18852,N_18519,N_18231);
nand U18853 (N_18853,N_18511,N_18167);
nand U18854 (N_18854,N_18235,N_18148);
nand U18855 (N_18855,N_17931,N_18350);
nor U18856 (N_18856,N_18210,N_18282);
or U18857 (N_18857,N_17521,N_18120);
nand U18858 (N_18858,N_18474,N_18106);
or U18859 (N_18859,N_17939,N_18663);
nor U18860 (N_18860,N_18071,N_17823);
nand U18861 (N_18861,N_17683,N_18347);
or U18862 (N_18862,N_17634,N_17645);
nor U18863 (N_18863,N_17690,N_18489);
nand U18864 (N_18864,N_18584,N_18527);
nand U18865 (N_18865,N_17801,N_18066);
and U18866 (N_18866,N_18114,N_18673);
xnor U18867 (N_18867,N_17830,N_17657);
xnor U18868 (N_18868,N_18253,N_17697);
and U18869 (N_18869,N_18083,N_17558);
xnor U18870 (N_18870,N_18281,N_17573);
or U18871 (N_18871,N_18192,N_18445);
nor U18872 (N_18872,N_18536,N_18032);
and U18873 (N_18873,N_18464,N_18479);
or U18874 (N_18874,N_17724,N_18069);
nor U18875 (N_18875,N_17879,N_18194);
nor U18876 (N_18876,N_17655,N_18470);
xnor U18877 (N_18877,N_18191,N_18093);
xor U18878 (N_18878,N_18560,N_18460);
nand U18879 (N_18879,N_18659,N_17597);
and U18880 (N_18880,N_18567,N_17768);
nand U18881 (N_18881,N_17700,N_18102);
nor U18882 (N_18882,N_18137,N_17650);
and U18883 (N_18883,N_18193,N_17901);
and U18884 (N_18884,N_18539,N_18215);
nor U18885 (N_18885,N_17653,N_18308);
nand U18886 (N_18886,N_18438,N_18504);
or U18887 (N_18887,N_18305,N_17552);
xor U18888 (N_18888,N_18717,N_17968);
and U18889 (N_18889,N_18214,N_18409);
xnor U18890 (N_18890,N_18269,N_18405);
or U18891 (N_18891,N_17742,N_17658);
nor U18892 (N_18892,N_18633,N_18345);
nor U18893 (N_18893,N_18645,N_18119);
nand U18894 (N_18894,N_18288,N_18528);
xnor U18895 (N_18895,N_17793,N_18441);
nand U18896 (N_18896,N_18221,N_18727);
or U18897 (N_18897,N_17928,N_18594);
nor U18898 (N_18898,N_17575,N_17850);
or U18899 (N_18899,N_18419,N_18576);
or U18900 (N_18900,N_17737,N_17513);
nand U18901 (N_18901,N_18572,N_17703);
and U18902 (N_18902,N_18436,N_18565);
and U18903 (N_18903,N_18580,N_18644);
nand U18904 (N_18904,N_18611,N_18692);
nand U18905 (N_18905,N_18531,N_18201);
or U18906 (N_18906,N_18175,N_18002);
xnor U18907 (N_18907,N_17626,N_17797);
or U18908 (N_18908,N_18486,N_18706);
nand U18909 (N_18909,N_18104,N_17946);
and U18910 (N_18910,N_18407,N_18250);
xor U18911 (N_18911,N_17919,N_17622);
and U18912 (N_18912,N_17607,N_17660);
and U18913 (N_18913,N_17859,N_18105);
xnor U18914 (N_18914,N_17792,N_18714);
or U18915 (N_18915,N_17911,N_18448);
xnor U18916 (N_18916,N_18552,N_17746);
or U18917 (N_18917,N_18512,N_17759);
and U18918 (N_18918,N_18462,N_17591);
or U18919 (N_18919,N_18217,N_17980);
and U18920 (N_18920,N_17544,N_18200);
xnor U18921 (N_18921,N_18181,N_18245);
nand U18922 (N_18922,N_18503,N_18074);
nand U18923 (N_18923,N_17517,N_18595);
nor U18924 (N_18924,N_18187,N_18577);
nor U18925 (N_18925,N_17772,N_17730);
or U18926 (N_18926,N_18283,N_17620);
nand U18927 (N_18927,N_17625,N_18625);
xnor U18928 (N_18928,N_18499,N_18557);
nor U18929 (N_18929,N_18467,N_17608);
and U18930 (N_18930,N_18735,N_18592);
or U18931 (N_18931,N_18023,N_18331);
nor U18932 (N_18932,N_18427,N_18001);
nor U18933 (N_18933,N_18255,N_17550);
or U18934 (N_18934,N_18284,N_17606);
nor U18935 (N_18935,N_18332,N_18683);
nand U18936 (N_18936,N_18731,N_17890);
nand U18937 (N_18937,N_17702,N_18321);
and U18938 (N_18938,N_18492,N_17893);
or U18939 (N_18939,N_17877,N_18473);
or U18940 (N_18940,N_18428,N_18468);
and U18941 (N_18941,N_17929,N_18524);
xnor U18942 (N_18942,N_18554,N_18067);
nand U18943 (N_18943,N_17574,N_18237);
nand U18944 (N_18944,N_18537,N_18730);
xor U18945 (N_18945,N_18160,N_18154);
and U18946 (N_18946,N_17846,N_18636);
nor U18947 (N_18947,N_17986,N_17755);
nor U18948 (N_18948,N_18691,N_18157);
nor U18949 (N_18949,N_18198,N_18437);
or U18950 (N_18950,N_18233,N_18725);
or U18951 (N_18951,N_17813,N_17843);
nor U18952 (N_18952,N_18084,N_17616);
or U18953 (N_18953,N_17833,N_18712);
xnor U18954 (N_18954,N_18624,N_18520);
and U18955 (N_18955,N_18627,N_18696);
nor U18956 (N_18956,N_18037,N_17698);
nand U18957 (N_18957,N_18053,N_18190);
xnor U18958 (N_18958,N_18701,N_18265);
nand U18959 (N_18959,N_18621,N_17648);
nand U18960 (N_18960,N_18346,N_17501);
nand U18961 (N_18961,N_17583,N_18062);
and U18962 (N_18962,N_18650,N_17640);
or U18963 (N_18963,N_18241,N_17810);
nor U18964 (N_18964,N_17674,N_17824);
and U18965 (N_18965,N_18425,N_17921);
nor U18966 (N_18966,N_18361,N_18422);
nor U18967 (N_18967,N_18719,N_17687);
xnor U18968 (N_18968,N_18574,N_18451);
nor U18969 (N_18969,N_17762,N_17679);
nor U18970 (N_18970,N_17581,N_18360);
xor U18971 (N_18971,N_18669,N_17510);
and U18972 (N_18972,N_18612,N_17745);
or U18973 (N_18973,N_18113,N_18555);
nor U18974 (N_18974,N_18335,N_18232);
nand U18975 (N_18975,N_18546,N_17545);
or U18976 (N_18976,N_18487,N_18729);
nor U18977 (N_18977,N_18741,N_18568);
nand U18978 (N_18978,N_18197,N_18130);
and U18979 (N_18979,N_18204,N_18220);
or U18980 (N_18980,N_17923,N_18144);
nand U18981 (N_18981,N_18304,N_18292);
and U18982 (N_18982,N_17509,N_17560);
xor U18983 (N_18983,N_17958,N_18208);
nand U18984 (N_18984,N_17854,N_18583);
nand U18985 (N_18985,N_18548,N_18606);
nand U18986 (N_18986,N_18632,N_18591);
or U18987 (N_18987,N_18421,N_18738);
or U18988 (N_18988,N_17582,N_17578);
and U18989 (N_18989,N_18506,N_17773);
or U18990 (N_18990,N_17696,N_18048);
or U18991 (N_18991,N_17990,N_18024);
nand U18992 (N_18992,N_18652,N_18185);
nor U18993 (N_18993,N_18025,N_18604);
xnor U18994 (N_18994,N_18619,N_17710);
and U18995 (N_18995,N_17665,N_18330);
xor U18996 (N_18996,N_17820,N_18150);
and U18997 (N_18997,N_17945,N_17540);
nand U18998 (N_18998,N_18239,N_18618);
and U18999 (N_18999,N_17862,N_18620);
and U19000 (N_19000,N_18247,N_17699);
and U19001 (N_19001,N_18146,N_18597);
nor U19002 (N_19002,N_18339,N_17994);
nor U19003 (N_19003,N_18410,N_18457);
nor U19004 (N_19004,N_18685,N_17503);
xnor U19005 (N_19005,N_17579,N_18563);
nand U19006 (N_19006,N_17987,N_18242);
or U19007 (N_19007,N_18072,N_17508);
nand U19008 (N_19008,N_17694,N_18510);
nor U19009 (N_19009,N_18373,N_18248);
xor U19010 (N_19010,N_17834,N_18517);
and U19011 (N_19011,N_18411,N_18482);
nand U19012 (N_19012,N_18224,N_17880);
nand U19013 (N_19013,N_17631,N_18165);
nor U19014 (N_19014,N_18188,N_18158);
or U19015 (N_19015,N_18159,N_18529);
nand U19016 (N_19016,N_18679,N_17926);
and U19017 (N_19017,N_18672,N_18277);
nand U19018 (N_19018,N_18086,N_17602);
and U19019 (N_19019,N_18454,N_18675);
nor U19020 (N_19020,N_18458,N_17519);
or U19021 (N_19021,N_18432,N_18635);
nor U19022 (N_19022,N_18262,N_18021);
nand U19023 (N_19023,N_17749,N_18401);
nor U19024 (N_19024,N_18413,N_18375);
xnor U19025 (N_19025,N_18140,N_17769);
nor U19026 (N_19026,N_17878,N_18513);
and U19027 (N_19027,N_17978,N_18099);
xor U19028 (N_19028,N_17953,N_18678);
xor U19029 (N_19029,N_18090,N_17955);
or U19030 (N_19030,N_17542,N_18525);
nand U19031 (N_19031,N_18206,N_17909);
and U19032 (N_19032,N_18153,N_18275);
xor U19033 (N_19033,N_17543,N_17957);
xnor U19034 (N_19034,N_17887,N_18324);
xor U19035 (N_19035,N_17537,N_17569);
xnor U19036 (N_19036,N_17505,N_18390);
nand U19037 (N_19037,N_17561,N_18266);
xnor U19038 (N_19038,N_17731,N_18055);
xor U19039 (N_19039,N_18211,N_17638);
nor U19040 (N_19040,N_17984,N_17991);
and U19041 (N_19041,N_17734,N_17902);
nand U19042 (N_19042,N_17584,N_17654);
and U19043 (N_19043,N_17709,N_17874);
and U19044 (N_19044,N_18736,N_18507);
or U19045 (N_19045,N_18170,N_18162);
or U19046 (N_19046,N_17774,N_17717);
or U19047 (N_19047,N_17872,N_18147);
nand U19048 (N_19048,N_17500,N_18585);
nor U19049 (N_19049,N_17627,N_18466);
nand U19050 (N_19050,N_18294,N_18008);
and U19051 (N_19051,N_17739,N_18276);
xnor U19052 (N_19052,N_17516,N_18073);
or U19053 (N_19053,N_18256,N_18455);
and U19054 (N_19054,N_17889,N_18212);
or U19055 (N_19055,N_17979,N_17549);
nor U19056 (N_19056,N_17808,N_17618);
or U19057 (N_19057,N_18225,N_17971);
nand U19058 (N_19058,N_17867,N_17763);
nand U19059 (N_19059,N_18749,N_18416);
xor U19060 (N_19060,N_18098,N_18562);
nor U19061 (N_19061,N_18496,N_17816);
nor U19062 (N_19062,N_17619,N_18371);
and U19063 (N_19063,N_18252,N_17706);
xnor U19064 (N_19064,N_17898,N_18223);
or U19065 (N_19065,N_18082,N_17882);
nand U19066 (N_19066,N_17688,N_17868);
nor U19067 (N_19067,N_18271,N_18034);
nor U19068 (N_19068,N_17985,N_17885);
nand U19069 (N_19069,N_17917,N_18388);
xor U19070 (N_19070,N_18423,N_17806);
or U19071 (N_19071,N_18091,N_17845);
or U19072 (N_19072,N_18301,N_17807);
and U19073 (N_19073,N_18312,N_18651);
xor U19074 (N_19074,N_18703,N_17628);
nor U19075 (N_19075,N_17840,N_17666);
or U19076 (N_19076,N_18397,N_17798);
xnor U19077 (N_19077,N_18348,N_17812);
nand U19078 (N_19078,N_17999,N_18057);
nor U19079 (N_19079,N_18480,N_18439);
xnor U19080 (N_19080,N_17779,N_18268);
nor U19081 (N_19081,N_18559,N_18195);
or U19082 (N_19082,N_18077,N_18688);
nor U19083 (N_19083,N_18354,N_18122);
and U19084 (N_19084,N_18178,N_17831);
nand U19085 (N_19085,N_18545,N_18363);
nand U19086 (N_19086,N_17775,N_18251);
or U19087 (N_19087,N_18440,N_18234);
and U19088 (N_19088,N_17675,N_18616);
and U19089 (N_19089,N_18009,N_18471);
and U19090 (N_19090,N_17756,N_18051);
nor U19091 (N_19091,N_17891,N_17960);
nand U19092 (N_19092,N_18186,N_18227);
nand U19093 (N_19093,N_17992,N_18096);
and U19094 (N_19094,N_17760,N_18734);
or U19095 (N_19095,N_18377,N_18088);
and U19096 (N_19096,N_18108,N_18740);
nor U19097 (N_19097,N_17857,N_18089);
nor U19098 (N_19098,N_17656,N_18521);
nor U19099 (N_19099,N_17783,N_18026);
and U19100 (N_19100,N_18526,N_18199);
and U19101 (N_19101,N_17944,N_17659);
or U19102 (N_19102,N_18267,N_18544);
and U19103 (N_19103,N_17809,N_17751);
xnor U19104 (N_19104,N_18420,N_17934);
or U19105 (N_19105,N_18382,N_17790);
or U19106 (N_19106,N_17556,N_18498);
nor U19107 (N_19107,N_18316,N_18588);
nand U19108 (N_19108,N_18038,N_18323);
or U19109 (N_19109,N_18075,N_18638);
xor U19110 (N_19110,N_17670,N_18298);
xor U19111 (N_19111,N_17982,N_17522);
xor U19112 (N_19112,N_18152,N_18249);
xor U19113 (N_19113,N_17529,N_18293);
nor U19114 (N_19114,N_17836,N_18647);
xnor U19115 (N_19115,N_17721,N_18733);
nand U19116 (N_19116,N_17594,N_17951);
nor U19117 (N_19117,N_18184,N_17827);
or U19118 (N_19118,N_17571,N_18522);
or U19119 (N_19119,N_17723,N_17672);
and U19120 (N_19120,N_18639,N_18012);
xor U19121 (N_19121,N_18497,N_18314);
and U19122 (N_19122,N_17711,N_18713);
or U19123 (N_19123,N_17750,N_18030);
nor U19124 (N_19124,N_17832,N_17924);
xor U19125 (N_19125,N_17533,N_17639);
nand U19126 (N_19126,N_18270,N_18433);
nor U19127 (N_19127,N_18033,N_17564);
or U19128 (N_19128,N_17577,N_18236);
nor U19129 (N_19129,N_18264,N_17701);
or U19130 (N_19130,N_17693,N_17829);
xor U19131 (N_19131,N_17532,N_17998);
xnor U19132 (N_19132,N_18417,N_18626);
nand U19133 (N_19133,N_17642,N_18472);
nor U19134 (N_19134,N_17689,N_18414);
or U19135 (N_19135,N_18174,N_17595);
and U19136 (N_19136,N_18556,N_18747);
nor U19137 (N_19137,N_17643,N_18728);
and U19138 (N_19138,N_18484,N_17632);
nand U19139 (N_19139,N_18311,N_18662);
and U19140 (N_19140,N_18286,N_18586);
or U19141 (N_19141,N_17844,N_17916);
nand U19142 (N_19142,N_17870,N_17727);
or U19143 (N_19143,N_18358,N_17966);
or U19144 (N_19144,N_18538,N_17531);
nor U19145 (N_19145,N_17972,N_18689);
xnor U19146 (N_19146,N_17791,N_17895);
or U19147 (N_19147,N_18461,N_17967);
nor U19148 (N_19148,N_17611,N_17789);
xor U19149 (N_19149,N_17681,N_17837);
nand U19150 (N_19150,N_18593,N_18476);
nor U19151 (N_19151,N_17787,N_17617);
xnor U19152 (N_19152,N_17514,N_18743);
and U19153 (N_19153,N_18022,N_17765);
nor U19154 (N_19154,N_17527,N_18325);
nor U19155 (N_19155,N_18605,N_17961);
and U19156 (N_19156,N_17927,N_18015);
nor U19157 (N_19157,N_18176,N_17515);
nand U19158 (N_19158,N_18044,N_17596);
nor U19159 (N_19159,N_18349,N_18643);
nor U19160 (N_19160,N_18501,N_17695);
or U19161 (N_19161,N_18333,N_17805);
and U19162 (N_19162,N_18549,N_18558);
or U19163 (N_19163,N_17770,N_18299);
and U19164 (N_19164,N_17821,N_18435);
or U19165 (N_19165,N_18340,N_18029);
and U19166 (N_19166,N_18341,N_18017);
and U19167 (N_19167,N_17685,N_17652);
or U19168 (N_19168,N_17959,N_17732);
and U19169 (N_19169,N_18387,N_18351);
and U19170 (N_19170,N_18711,N_18258);
nor U19171 (N_19171,N_18434,N_17680);
or U19172 (N_19172,N_18690,N_18613);
or U19173 (N_19173,N_17506,N_18343);
and U19174 (N_19174,N_17969,N_17828);
and U19175 (N_19175,N_17623,N_17933);
nor U19176 (N_19176,N_18244,N_17651);
or U19177 (N_19177,N_17973,N_18648);
xnor U19178 (N_19178,N_18123,N_18117);
nor U19179 (N_19179,N_18392,N_17752);
xnor U19180 (N_19180,N_18542,N_18547);
or U19181 (N_19181,N_18516,N_18142);
nor U19182 (N_19182,N_17906,N_18357);
and U19183 (N_19183,N_17892,N_18353);
or U19184 (N_19184,N_17786,N_18367);
nor U19185 (N_19185,N_18478,N_17855);
nor U19186 (N_19186,N_17896,N_17598);
xor U19187 (N_19187,N_17976,N_17563);
nand U19188 (N_19188,N_18138,N_18004);
xnor U19189 (N_19189,N_17803,N_18705);
and U19190 (N_19190,N_17518,N_18686);
nor U19191 (N_19191,N_18630,N_17567);
nor U19192 (N_19192,N_17557,N_18319);
and U19193 (N_19193,N_18579,N_17884);
nor U19194 (N_19194,N_17841,N_18370);
and U19195 (N_19195,N_18202,N_18064);
xnor U19196 (N_19196,N_18059,N_17568);
xor U19197 (N_19197,N_18430,N_17842);
nand U19198 (N_19198,N_17757,N_18681);
and U19199 (N_19199,N_17555,N_17852);
xnor U19200 (N_19200,N_17526,N_18682);
xor U19201 (N_19201,N_18352,N_18322);
xnor U19202 (N_19202,N_18366,N_18610);
nor U19203 (N_19203,N_17671,N_17720);
nor U19204 (N_19204,N_18540,N_18737);
or U19205 (N_19205,N_18700,N_18475);
nand U19206 (N_19206,N_17538,N_17605);
xnor U19207 (N_19207,N_17780,N_18656);
or U19208 (N_19208,N_18111,N_18196);
nand U19209 (N_19209,N_18502,N_18376);
and U19210 (N_19210,N_17920,N_18313);
xor U19211 (N_19211,N_17572,N_17886);
xnor U19212 (N_19212,N_18261,N_17863);
xor U19213 (N_19213,N_18745,N_18131);
nor U19214 (N_19214,N_18653,N_17586);
xor U19215 (N_19215,N_18581,N_17726);
xor U19216 (N_19216,N_18561,N_17600);
nor U19217 (N_19217,N_17848,N_18189);
nor U19218 (N_19218,N_17580,N_18041);
nor U19219 (N_19219,N_17930,N_18303);
xor U19220 (N_19220,N_18164,N_18014);
or U19221 (N_19221,N_18424,N_18450);
or U19222 (N_19222,N_18166,N_17511);
nor U19223 (N_19223,N_18655,N_18631);
and U19224 (N_19224,N_18035,N_17778);
or U19225 (N_19225,N_18000,N_17881);
nor U19226 (N_19226,N_18447,N_17610);
and U19227 (N_19227,N_17754,N_18209);
nor U19228 (N_19228,N_17637,N_17860);
and U19229 (N_19229,N_17725,N_17609);
nor U19230 (N_19230,N_18135,N_18710);
or U19231 (N_19231,N_18443,N_17562);
or U19232 (N_19232,N_18637,N_17668);
or U19233 (N_19233,N_17948,N_18534);
nand U19234 (N_19234,N_18622,N_17647);
nand U19235 (N_19235,N_18657,N_18338);
nand U19236 (N_19236,N_17604,N_18027);
and U19237 (N_19237,N_18116,N_18490);
nor U19238 (N_19238,N_17819,N_18087);
or U19239 (N_19239,N_18278,N_18600);
nand U19240 (N_19240,N_17667,N_18179);
and U19241 (N_19241,N_18607,N_18129);
nor U19242 (N_19242,N_18603,N_18722);
or U19243 (N_19243,N_18412,N_18046);
xnor U19244 (N_19244,N_18039,N_18726);
nand U19245 (N_19245,N_18641,N_18222);
nor U19246 (N_19246,N_18326,N_18623);
nand U19247 (N_19247,N_17856,N_17716);
nor U19248 (N_19248,N_17678,N_18541);
or U19249 (N_19249,N_17504,N_18495);
nand U19250 (N_19250,N_17873,N_17764);
nor U19251 (N_19251,N_18698,N_17849);
nand U19252 (N_19252,N_18550,N_18133);
nor U19253 (N_19253,N_17738,N_17894);
and U19254 (N_19254,N_18372,N_17970);
nand U19255 (N_19255,N_18121,N_18658);
xor U19256 (N_19256,N_17744,N_18219);
and U19257 (N_19257,N_17963,N_18045);
nand U19258 (N_19258,N_17502,N_17590);
and U19259 (N_19259,N_18379,N_18081);
and U19260 (N_19260,N_17941,N_18010);
nor U19261 (N_19261,N_18408,N_17858);
and U19262 (N_19262,N_18415,N_17612);
or U19263 (N_19263,N_18115,N_18344);
and U19264 (N_19264,N_17800,N_18601);
xor U19265 (N_19265,N_18723,N_17776);
xnor U19266 (N_19266,N_18515,N_18309);
nor U19267 (N_19267,N_17799,N_17871);
or U19268 (N_19268,N_17661,N_18608);
or U19269 (N_19269,N_18050,N_18061);
nand U19270 (N_19270,N_17853,N_18739);
and U19271 (N_19271,N_18553,N_18272);
or U19272 (N_19272,N_18095,N_17781);
nand U19273 (N_19273,N_18005,N_17525);
nand U19274 (N_19274,N_18139,N_18596);
nor U19275 (N_19275,N_18307,N_18100);
or U19276 (N_19276,N_17587,N_18446);
nand U19277 (N_19277,N_18569,N_18699);
xor U19278 (N_19278,N_18013,N_17624);
nor U19279 (N_19279,N_18532,N_18514);
nand U19280 (N_19280,N_18744,N_18182);
xor U19281 (N_19281,N_17988,N_18334);
and U19282 (N_19282,N_18317,N_18398);
or U19283 (N_19283,N_17534,N_17684);
or U19284 (N_19284,N_18393,N_18665);
or U19285 (N_19285,N_17570,N_18163);
xnor U19286 (N_19286,N_18614,N_18399);
nand U19287 (N_19287,N_17589,N_17907);
nand U19288 (N_19288,N_18693,N_18016);
xor U19289 (N_19289,N_17915,N_18097);
xnor U19290 (N_19290,N_18126,N_18667);
or U19291 (N_19291,N_18718,N_18289);
or U19292 (N_19292,N_18748,N_17796);
nor U19293 (N_19293,N_17554,N_18680);
nor U19294 (N_19294,N_18132,N_18369);
and U19295 (N_19295,N_17636,N_18124);
and U19296 (N_19296,N_17673,N_17804);
nor U19297 (N_19297,N_17733,N_18040);
xnor U19298 (N_19298,N_17553,N_18671);
and U19299 (N_19299,N_17950,N_17943);
or U19300 (N_19300,N_17899,N_17866);
nand U19301 (N_19301,N_18101,N_17613);
xnor U19302 (N_19302,N_17715,N_17676);
or U19303 (N_19303,N_17664,N_18702);
and U19304 (N_19304,N_18400,N_17925);
nand U19305 (N_19305,N_18649,N_18279);
nand U19306 (N_19306,N_18687,N_17633);
xnor U19307 (N_19307,N_18109,N_18617);
nand U19308 (N_19308,N_18456,N_18079);
or U19309 (N_19309,N_18107,N_18695);
nand U19310 (N_19310,N_18640,N_18300);
or U19311 (N_19311,N_18518,N_17777);
or U19312 (N_19312,N_18306,N_17864);
or U19313 (N_19313,N_17835,N_18661);
nand U19314 (N_19314,N_18052,N_18337);
nor U19315 (N_19315,N_17741,N_18493);
nand U19316 (N_19316,N_17629,N_18704);
or U19317 (N_19317,N_17712,N_17718);
nand U19318 (N_19318,N_17914,N_18459);
nor U19319 (N_19319,N_18065,N_17713);
nor U19320 (N_19320,N_18677,N_18674);
and U19321 (N_19321,N_18394,N_18177);
and U19322 (N_19322,N_18020,N_17802);
and U19323 (N_19323,N_18732,N_18615);
nand U19324 (N_19324,N_18429,N_18573);
xnor U19325 (N_19325,N_18491,N_18395);
and U19326 (N_19326,N_17635,N_17876);
or U19327 (N_19327,N_17663,N_17869);
or U19328 (N_19328,N_17904,N_18285);
or U19329 (N_19329,N_18006,N_18494);
xnor U19330 (N_19330,N_18031,N_18380);
xnor U19331 (N_19331,N_18183,N_18668);
nand U19332 (N_19332,N_18143,N_18452);
nand U19333 (N_19333,N_17822,N_18218);
xor U19334 (N_19334,N_17932,N_17566);
or U19335 (N_19335,N_17535,N_18060);
or U19336 (N_19336,N_18359,N_18134);
nand U19337 (N_19337,N_18203,N_18172);
xnor U19338 (N_19338,N_17900,N_17669);
nand U19339 (N_19339,N_18477,N_18483);
or U19340 (N_19340,N_18068,N_18171);
nor U19341 (N_19341,N_18389,N_17528);
xnor U19342 (N_19342,N_17956,N_17922);
and U19343 (N_19343,N_17649,N_17839);
and U19344 (N_19344,N_18582,N_18011);
xor U19345 (N_19345,N_17704,N_18386);
or U19346 (N_19346,N_18551,N_18590);
and U19347 (N_19347,N_18149,N_17937);
or U19348 (N_19348,N_17938,N_17826);
and U19349 (N_19349,N_18716,N_17785);
and U19350 (N_19350,N_18085,N_18246);
nor U19351 (N_19351,N_17682,N_18128);
nand U19352 (N_19352,N_17767,N_17507);
or U19353 (N_19353,N_17903,N_18530);
or U19354 (N_19354,N_18381,N_18257);
or U19355 (N_19355,N_18724,N_18336);
nor U19356 (N_19356,N_18356,N_18141);
nand U19357 (N_19357,N_18535,N_18259);
or U19358 (N_19358,N_17708,N_18449);
or U19359 (N_19359,N_17910,N_18173);
xnor U19360 (N_19360,N_18403,N_17942);
or U19361 (N_19361,N_17740,N_18078);
or U19362 (N_19362,N_18646,N_18043);
or U19363 (N_19363,N_18318,N_17686);
or U19364 (N_19364,N_17795,N_18599);
xnor U19365 (N_19365,N_18708,N_17565);
and U19366 (N_19366,N_18263,N_17641);
and U19367 (N_19367,N_18508,N_18676);
nand U19368 (N_19368,N_17548,N_17758);
xor U19369 (N_19369,N_17599,N_17753);
nor U19370 (N_19370,N_18715,N_18145);
xnor U19371 (N_19371,N_17975,N_18047);
and U19372 (N_19372,N_18054,N_17814);
or U19373 (N_19373,N_18431,N_18018);
nand U19374 (N_19374,N_17728,N_17576);
nor U19375 (N_19375,N_18224,N_17729);
and U19376 (N_19376,N_17797,N_17792);
xor U19377 (N_19377,N_18043,N_18484);
or U19378 (N_19378,N_17656,N_18274);
or U19379 (N_19379,N_17655,N_17569);
xor U19380 (N_19380,N_18735,N_18432);
or U19381 (N_19381,N_18236,N_17816);
or U19382 (N_19382,N_18603,N_18149);
nor U19383 (N_19383,N_18462,N_18159);
or U19384 (N_19384,N_17689,N_18330);
nor U19385 (N_19385,N_17609,N_18146);
nand U19386 (N_19386,N_17583,N_18385);
and U19387 (N_19387,N_18338,N_17581);
or U19388 (N_19388,N_18071,N_17816);
or U19389 (N_19389,N_17593,N_18276);
and U19390 (N_19390,N_18160,N_17756);
xor U19391 (N_19391,N_18584,N_18564);
and U19392 (N_19392,N_17800,N_17922);
or U19393 (N_19393,N_17907,N_17517);
and U19394 (N_19394,N_17898,N_17969);
nor U19395 (N_19395,N_18712,N_18327);
nand U19396 (N_19396,N_17643,N_17521);
and U19397 (N_19397,N_18043,N_18510);
nand U19398 (N_19398,N_17870,N_18314);
xnor U19399 (N_19399,N_18289,N_18058);
and U19400 (N_19400,N_17909,N_18379);
nand U19401 (N_19401,N_17983,N_18128);
or U19402 (N_19402,N_18386,N_17625);
nand U19403 (N_19403,N_17679,N_18271);
nand U19404 (N_19404,N_18019,N_18461);
or U19405 (N_19405,N_17522,N_17895);
nand U19406 (N_19406,N_18654,N_17686);
xnor U19407 (N_19407,N_18413,N_18574);
nor U19408 (N_19408,N_18051,N_17822);
and U19409 (N_19409,N_18023,N_18640);
nor U19410 (N_19410,N_17594,N_18719);
or U19411 (N_19411,N_17776,N_18689);
nor U19412 (N_19412,N_18376,N_18308);
and U19413 (N_19413,N_17910,N_18028);
and U19414 (N_19414,N_18395,N_17832);
nor U19415 (N_19415,N_18483,N_18353);
nand U19416 (N_19416,N_18366,N_18420);
or U19417 (N_19417,N_17571,N_18444);
and U19418 (N_19418,N_17988,N_18456);
xnor U19419 (N_19419,N_17878,N_18115);
or U19420 (N_19420,N_18251,N_18205);
xnor U19421 (N_19421,N_17870,N_17576);
or U19422 (N_19422,N_17770,N_18151);
nand U19423 (N_19423,N_18267,N_17684);
xor U19424 (N_19424,N_17784,N_18326);
nor U19425 (N_19425,N_17524,N_17956);
nor U19426 (N_19426,N_17956,N_18265);
xor U19427 (N_19427,N_17544,N_17844);
or U19428 (N_19428,N_18283,N_17604);
and U19429 (N_19429,N_18362,N_18407);
xnor U19430 (N_19430,N_17777,N_17560);
xnor U19431 (N_19431,N_18045,N_18466);
or U19432 (N_19432,N_18261,N_18546);
nand U19433 (N_19433,N_18702,N_18352);
and U19434 (N_19434,N_17873,N_17540);
or U19435 (N_19435,N_18419,N_18312);
xor U19436 (N_19436,N_17603,N_18089);
xnor U19437 (N_19437,N_18298,N_18395);
xnor U19438 (N_19438,N_17584,N_18017);
xnor U19439 (N_19439,N_18558,N_17992);
nand U19440 (N_19440,N_18425,N_17783);
nor U19441 (N_19441,N_18467,N_17894);
and U19442 (N_19442,N_18625,N_17692);
xnor U19443 (N_19443,N_17908,N_18063);
xnor U19444 (N_19444,N_17794,N_17985);
nand U19445 (N_19445,N_17917,N_18423);
nor U19446 (N_19446,N_18644,N_17509);
or U19447 (N_19447,N_18747,N_17852);
and U19448 (N_19448,N_18126,N_18463);
xor U19449 (N_19449,N_17703,N_17721);
xor U19450 (N_19450,N_18473,N_18120);
nand U19451 (N_19451,N_18579,N_18638);
nor U19452 (N_19452,N_18500,N_18737);
or U19453 (N_19453,N_17642,N_17912);
or U19454 (N_19454,N_18063,N_18423);
and U19455 (N_19455,N_17838,N_17927);
or U19456 (N_19456,N_18453,N_18685);
nand U19457 (N_19457,N_18437,N_17656);
xor U19458 (N_19458,N_18098,N_18587);
or U19459 (N_19459,N_17915,N_18306);
nand U19460 (N_19460,N_18283,N_18514);
nor U19461 (N_19461,N_17748,N_17690);
nor U19462 (N_19462,N_18035,N_18137);
nor U19463 (N_19463,N_18088,N_17685);
and U19464 (N_19464,N_18477,N_18188);
nand U19465 (N_19465,N_18434,N_17869);
nand U19466 (N_19466,N_17778,N_17620);
and U19467 (N_19467,N_17565,N_18163);
xor U19468 (N_19468,N_18295,N_17822);
and U19469 (N_19469,N_17838,N_18636);
nor U19470 (N_19470,N_18454,N_18469);
and U19471 (N_19471,N_18668,N_18605);
nand U19472 (N_19472,N_18207,N_18031);
or U19473 (N_19473,N_18351,N_18558);
nor U19474 (N_19474,N_18276,N_18723);
or U19475 (N_19475,N_18083,N_18341);
nor U19476 (N_19476,N_17906,N_17870);
nand U19477 (N_19477,N_17793,N_18429);
nor U19478 (N_19478,N_18494,N_18596);
xnor U19479 (N_19479,N_18605,N_18322);
xnor U19480 (N_19480,N_18136,N_18394);
and U19481 (N_19481,N_17506,N_17740);
or U19482 (N_19482,N_17610,N_18600);
nor U19483 (N_19483,N_18517,N_17909);
and U19484 (N_19484,N_17532,N_17756);
and U19485 (N_19485,N_17831,N_17917);
nand U19486 (N_19486,N_17640,N_18132);
xor U19487 (N_19487,N_17925,N_17659);
nor U19488 (N_19488,N_17552,N_18115);
nor U19489 (N_19489,N_18747,N_18619);
or U19490 (N_19490,N_17742,N_18411);
and U19491 (N_19491,N_18072,N_17655);
and U19492 (N_19492,N_17914,N_18547);
and U19493 (N_19493,N_18545,N_17983);
and U19494 (N_19494,N_17853,N_18694);
nor U19495 (N_19495,N_18723,N_18612);
and U19496 (N_19496,N_18538,N_17538);
or U19497 (N_19497,N_17872,N_18444);
nand U19498 (N_19498,N_18748,N_18714);
or U19499 (N_19499,N_18745,N_17573);
xnor U19500 (N_19500,N_18386,N_18324);
nand U19501 (N_19501,N_17685,N_17918);
xnor U19502 (N_19502,N_17769,N_17995);
nand U19503 (N_19503,N_17988,N_17667);
xnor U19504 (N_19504,N_18509,N_18603);
nor U19505 (N_19505,N_17875,N_18036);
or U19506 (N_19506,N_18121,N_17546);
xor U19507 (N_19507,N_18677,N_17989);
nand U19508 (N_19508,N_18665,N_18233);
xor U19509 (N_19509,N_17582,N_18538);
nand U19510 (N_19510,N_17635,N_17787);
xor U19511 (N_19511,N_17946,N_18007);
and U19512 (N_19512,N_17791,N_17549);
nor U19513 (N_19513,N_17825,N_18261);
nand U19514 (N_19514,N_18579,N_18538);
and U19515 (N_19515,N_18208,N_17631);
nand U19516 (N_19516,N_17784,N_18248);
nor U19517 (N_19517,N_17534,N_17750);
and U19518 (N_19518,N_18498,N_17743);
nand U19519 (N_19519,N_17869,N_18021);
xnor U19520 (N_19520,N_17942,N_18191);
and U19521 (N_19521,N_18609,N_18156);
nand U19522 (N_19522,N_17586,N_18294);
xnor U19523 (N_19523,N_18626,N_17511);
nor U19524 (N_19524,N_18574,N_18328);
nor U19525 (N_19525,N_18179,N_18336);
nand U19526 (N_19526,N_18093,N_17898);
and U19527 (N_19527,N_18336,N_18613);
or U19528 (N_19528,N_18403,N_17882);
and U19529 (N_19529,N_18261,N_18028);
nand U19530 (N_19530,N_18113,N_18530);
and U19531 (N_19531,N_18222,N_18432);
or U19532 (N_19532,N_18117,N_17941);
or U19533 (N_19533,N_18743,N_18502);
xor U19534 (N_19534,N_17504,N_18340);
or U19535 (N_19535,N_18397,N_17610);
xor U19536 (N_19536,N_18623,N_17723);
xnor U19537 (N_19537,N_17650,N_18716);
nor U19538 (N_19538,N_17953,N_18178);
or U19539 (N_19539,N_17834,N_17859);
xor U19540 (N_19540,N_18259,N_18095);
nand U19541 (N_19541,N_18067,N_18096);
nor U19542 (N_19542,N_17779,N_18556);
nor U19543 (N_19543,N_18566,N_17546);
nor U19544 (N_19544,N_17826,N_18006);
or U19545 (N_19545,N_18029,N_17957);
nand U19546 (N_19546,N_18506,N_17559);
nor U19547 (N_19547,N_17823,N_18244);
or U19548 (N_19548,N_18474,N_18415);
or U19549 (N_19549,N_18399,N_18544);
or U19550 (N_19550,N_18642,N_18285);
and U19551 (N_19551,N_18633,N_18132);
nand U19552 (N_19552,N_17975,N_17545);
or U19553 (N_19553,N_17615,N_18117);
nand U19554 (N_19554,N_18365,N_18585);
nor U19555 (N_19555,N_17983,N_18591);
or U19556 (N_19556,N_18376,N_18511);
and U19557 (N_19557,N_18367,N_18284);
nand U19558 (N_19558,N_18692,N_17786);
nand U19559 (N_19559,N_18557,N_18521);
nand U19560 (N_19560,N_18578,N_18098);
and U19561 (N_19561,N_17861,N_18248);
xnor U19562 (N_19562,N_18056,N_18417);
nor U19563 (N_19563,N_18419,N_18231);
nor U19564 (N_19564,N_18055,N_18135);
nand U19565 (N_19565,N_18211,N_18164);
and U19566 (N_19566,N_17684,N_18325);
xor U19567 (N_19567,N_18576,N_17758);
xnor U19568 (N_19568,N_17632,N_17786);
nor U19569 (N_19569,N_17656,N_18075);
or U19570 (N_19570,N_18691,N_17559);
nor U19571 (N_19571,N_18722,N_18564);
and U19572 (N_19572,N_18464,N_17599);
nor U19573 (N_19573,N_17976,N_18475);
or U19574 (N_19574,N_18116,N_18717);
and U19575 (N_19575,N_17561,N_18110);
nand U19576 (N_19576,N_18629,N_17728);
nor U19577 (N_19577,N_17820,N_18222);
or U19578 (N_19578,N_18716,N_18693);
or U19579 (N_19579,N_18441,N_18307);
and U19580 (N_19580,N_18617,N_17668);
xnor U19581 (N_19581,N_17708,N_17688);
xor U19582 (N_19582,N_18351,N_18456);
xor U19583 (N_19583,N_17789,N_18122);
nand U19584 (N_19584,N_17893,N_17576);
and U19585 (N_19585,N_17677,N_18425);
and U19586 (N_19586,N_18370,N_17782);
nor U19587 (N_19587,N_17822,N_18675);
and U19588 (N_19588,N_18405,N_18154);
xnor U19589 (N_19589,N_17742,N_18197);
or U19590 (N_19590,N_17741,N_17767);
nand U19591 (N_19591,N_17951,N_17567);
nor U19592 (N_19592,N_17625,N_18164);
and U19593 (N_19593,N_18128,N_17796);
or U19594 (N_19594,N_17614,N_18697);
or U19595 (N_19595,N_18260,N_18596);
nor U19596 (N_19596,N_17518,N_18044);
xnor U19597 (N_19597,N_18105,N_17544);
or U19598 (N_19598,N_17771,N_18345);
nand U19599 (N_19599,N_17856,N_18661);
xnor U19600 (N_19600,N_18657,N_18706);
nand U19601 (N_19601,N_17616,N_18188);
nand U19602 (N_19602,N_18182,N_18299);
nor U19603 (N_19603,N_18527,N_18148);
and U19604 (N_19604,N_17655,N_18223);
nand U19605 (N_19605,N_18680,N_17767);
nor U19606 (N_19606,N_17739,N_17917);
and U19607 (N_19607,N_17866,N_17763);
xnor U19608 (N_19608,N_17814,N_18282);
nor U19609 (N_19609,N_17820,N_18487);
and U19610 (N_19610,N_18253,N_18678);
or U19611 (N_19611,N_18234,N_18531);
nand U19612 (N_19612,N_18698,N_18311);
nand U19613 (N_19613,N_18461,N_18302);
and U19614 (N_19614,N_17723,N_17501);
or U19615 (N_19615,N_18531,N_18293);
and U19616 (N_19616,N_17751,N_17883);
and U19617 (N_19617,N_18499,N_17830);
nor U19618 (N_19618,N_18678,N_18303);
nand U19619 (N_19619,N_18104,N_17527);
nand U19620 (N_19620,N_17766,N_17959);
or U19621 (N_19621,N_17838,N_17978);
or U19622 (N_19622,N_18614,N_18196);
or U19623 (N_19623,N_18170,N_18561);
or U19624 (N_19624,N_18013,N_17999);
nand U19625 (N_19625,N_18720,N_17648);
nor U19626 (N_19626,N_17766,N_18555);
or U19627 (N_19627,N_18585,N_18023);
xnor U19628 (N_19628,N_18668,N_18014);
and U19629 (N_19629,N_18222,N_18331);
or U19630 (N_19630,N_18016,N_17611);
nor U19631 (N_19631,N_17643,N_17519);
and U19632 (N_19632,N_18382,N_18725);
or U19633 (N_19633,N_18017,N_18290);
nand U19634 (N_19634,N_18360,N_18465);
nand U19635 (N_19635,N_17671,N_17902);
and U19636 (N_19636,N_17779,N_18458);
nand U19637 (N_19637,N_18051,N_18724);
or U19638 (N_19638,N_17729,N_18671);
xor U19639 (N_19639,N_18358,N_18659);
and U19640 (N_19640,N_18215,N_18468);
and U19641 (N_19641,N_18237,N_18648);
nor U19642 (N_19642,N_18432,N_18454);
nand U19643 (N_19643,N_18028,N_17544);
or U19644 (N_19644,N_17933,N_17656);
nand U19645 (N_19645,N_18418,N_18413);
nand U19646 (N_19646,N_17676,N_18508);
xor U19647 (N_19647,N_17767,N_17790);
nand U19648 (N_19648,N_18029,N_18154);
nand U19649 (N_19649,N_17535,N_17888);
nor U19650 (N_19650,N_17505,N_18541);
or U19651 (N_19651,N_18064,N_17757);
or U19652 (N_19652,N_17709,N_18043);
and U19653 (N_19653,N_18559,N_18705);
xor U19654 (N_19654,N_18432,N_17843);
nor U19655 (N_19655,N_17554,N_18587);
nor U19656 (N_19656,N_17744,N_17795);
and U19657 (N_19657,N_17742,N_17752);
nand U19658 (N_19658,N_18103,N_18165);
or U19659 (N_19659,N_18291,N_18476);
nor U19660 (N_19660,N_18655,N_18195);
nand U19661 (N_19661,N_18426,N_18674);
and U19662 (N_19662,N_17768,N_17569);
xnor U19663 (N_19663,N_17575,N_18102);
or U19664 (N_19664,N_18623,N_18533);
xor U19665 (N_19665,N_17570,N_18514);
and U19666 (N_19666,N_17580,N_18364);
nor U19667 (N_19667,N_18188,N_17694);
nor U19668 (N_19668,N_17749,N_18381);
nor U19669 (N_19669,N_18079,N_18233);
nor U19670 (N_19670,N_18283,N_17546);
nor U19671 (N_19671,N_18688,N_18173);
or U19672 (N_19672,N_17886,N_18264);
nor U19673 (N_19673,N_18134,N_18495);
nor U19674 (N_19674,N_18376,N_18239);
nor U19675 (N_19675,N_18736,N_18460);
or U19676 (N_19676,N_17905,N_17910);
and U19677 (N_19677,N_18738,N_18655);
or U19678 (N_19678,N_18623,N_17679);
nand U19679 (N_19679,N_18305,N_17830);
and U19680 (N_19680,N_18540,N_17732);
nand U19681 (N_19681,N_17686,N_18282);
nand U19682 (N_19682,N_17735,N_17899);
nand U19683 (N_19683,N_18424,N_18179);
nand U19684 (N_19684,N_18509,N_18440);
or U19685 (N_19685,N_17924,N_18075);
and U19686 (N_19686,N_17835,N_18695);
nand U19687 (N_19687,N_18259,N_18593);
nand U19688 (N_19688,N_17690,N_17788);
and U19689 (N_19689,N_17800,N_18457);
xnor U19690 (N_19690,N_18715,N_17641);
and U19691 (N_19691,N_18702,N_18119);
nor U19692 (N_19692,N_17589,N_18224);
or U19693 (N_19693,N_18121,N_18067);
nor U19694 (N_19694,N_18476,N_18688);
xnor U19695 (N_19695,N_18226,N_18251);
and U19696 (N_19696,N_18262,N_18025);
xnor U19697 (N_19697,N_18300,N_18713);
nor U19698 (N_19698,N_17841,N_18578);
nor U19699 (N_19699,N_18690,N_17900);
or U19700 (N_19700,N_18168,N_17756);
nand U19701 (N_19701,N_18094,N_18110);
nor U19702 (N_19702,N_18332,N_17516);
xor U19703 (N_19703,N_18158,N_18516);
nor U19704 (N_19704,N_18363,N_18669);
xor U19705 (N_19705,N_18379,N_18622);
xnor U19706 (N_19706,N_18475,N_18591);
nand U19707 (N_19707,N_18487,N_17621);
and U19708 (N_19708,N_18191,N_18334);
or U19709 (N_19709,N_18053,N_18073);
or U19710 (N_19710,N_17584,N_17755);
and U19711 (N_19711,N_17606,N_17735);
or U19712 (N_19712,N_17762,N_17994);
and U19713 (N_19713,N_17566,N_18746);
and U19714 (N_19714,N_18431,N_17612);
and U19715 (N_19715,N_17647,N_18413);
nand U19716 (N_19716,N_18390,N_17654);
nand U19717 (N_19717,N_17830,N_17710);
or U19718 (N_19718,N_18081,N_18174);
and U19719 (N_19719,N_17604,N_17661);
xor U19720 (N_19720,N_18546,N_18568);
nand U19721 (N_19721,N_17511,N_17578);
or U19722 (N_19722,N_18332,N_18538);
nor U19723 (N_19723,N_18074,N_18517);
xnor U19724 (N_19724,N_18250,N_17694);
nor U19725 (N_19725,N_18148,N_17673);
nand U19726 (N_19726,N_18353,N_18231);
and U19727 (N_19727,N_18396,N_17591);
xnor U19728 (N_19728,N_18351,N_18597);
xor U19729 (N_19729,N_18647,N_18054);
nor U19730 (N_19730,N_18244,N_18050);
or U19731 (N_19731,N_18265,N_18337);
nor U19732 (N_19732,N_18473,N_18223);
or U19733 (N_19733,N_18331,N_18202);
or U19734 (N_19734,N_18199,N_17738);
nor U19735 (N_19735,N_17972,N_17890);
or U19736 (N_19736,N_17591,N_17965);
and U19737 (N_19737,N_18732,N_18215);
or U19738 (N_19738,N_18635,N_18146);
nand U19739 (N_19739,N_18559,N_17773);
xnor U19740 (N_19740,N_18528,N_17880);
xnor U19741 (N_19741,N_18124,N_18613);
and U19742 (N_19742,N_17520,N_18599);
nand U19743 (N_19743,N_17904,N_17656);
and U19744 (N_19744,N_18456,N_17966);
and U19745 (N_19745,N_17869,N_18548);
or U19746 (N_19746,N_18191,N_18193);
or U19747 (N_19747,N_17885,N_17750);
nand U19748 (N_19748,N_17779,N_18125);
and U19749 (N_19749,N_18689,N_18640);
nand U19750 (N_19750,N_18109,N_18693);
or U19751 (N_19751,N_17747,N_17875);
or U19752 (N_19752,N_18388,N_17567);
and U19753 (N_19753,N_18180,N_17991);
xor U19754 (N_19754,N_18329,N_18061);
nand U19755 (N_19755,N_18527,N_18108);
nand U19756 (N_19756,N_18609,N_17653);
or U19757 (N_19757,N_18100,N_17638);
or U19758 (N_19758,N_17662,N_17749);
nand U19759 (N_19759,N_17505,N_18668);
nand U19760 (N_19760,N_17585,N_17738);
xnor U19761 (N_19761,N_17703,N_18334);
nor U19762 (N_19762,N_18065,N_18667);
nor U19763 (N_19763,N_17646,N_17706);
or U19764 (N_19764,N_18683,N_18618);
or U19765 (N_19765,N_18410,N_18318);
or U19766 (N_19766,N_17752,N_18527);
xor U19767 (N_19767,N_18659,N_18344);
nor U19768 (N_19768,N_18316,N_17713);
xor U19769 (N_19769,N_17635,N_17739);
xor U19770 (N_19770,N_18301,N_18145);
and U19771 (N_19771,N_18513,N_18294);
nand U19772 (N_19772,N_18215,N_17869);
nand U19773 (N_19773,N_18343,N_17863);
or U19774 (N_19774,N_17803,N_18263);
nor U19775 (N_19775,N_18125,N_18290);
and U19776 (N_19776,N_18100,N_18189);
nor U19777 (N_19777,N_18669,N_18051);
nand U19778 (N_19778,N_17755,N_17559);
xor U19779 (N_19779,N_18380,N_17539);
xnor U19780 (N_19780,N_18278,N_18737);
and U19781 (N_19781,N_18040,N_17619);
or U19782 (N_19782,N_17731,N_17897);
and U19783 (N_19783,N_17863,N_17841);
nor U19784 (N_19784,N_17556,N_18560);
xnor U19785 (N_19785,N_18607,N_17886);
xnor U19786 (N_19786,N_17717,N_18653);
or U19787 (N_19787,N_17606,N_18156);
or U19788 (N_19788,N_17989,N_17508);
or U19789 (N_19789,N_18005,N_18136);
or U19790 (N_19790,N_17702,N_18083);
nand U19791 (N_19791,N_18475,N_18325);
and U19792 (N_19792,N_18123,N_18186);
nor U19793 (N_19793,N_18294,N_17620);
and U19794 (N_19794,N_17699,N_18741);
nor U19795 (N_19795,N_17686,N_18553);
or U19796 (N_19796,N_17609,N_18140);
xor U19797 (N_19797,N_18378,N_18614);
or U19798 (N_19798,N_17633,N_18645);
nand U19799 (N_19799,N_18530,N_18719);
nand U19800 (N_19800,N_18417,N_18169);
or U19801 (N_19801,N_18121,N_17828);
or U19802 (N_19802,N_18587,N_17907);
nor U19803 (N_19803,N_17963,N_18538);
and U19804 (N_19804,N_17994,N_18326);
nor U19805 (N_19805,N_18239,N_18131);
nand U19806 (N_19806,N_18140,N_18522);
or U19807 (N_19807,N_18678,N_18640);
nor U19808 (N_19808,N_18440,N_17628);
and U19809 (N_19809,N_17766,N_17942);
and U19810 (N_19810,N_17634,N_18077);
nand U19811 (N_19811,N_17887,N_18686);
and U19812 (N_19812,N_18002,N_18612);
nor U19813 (N_19813,N_18527,N_18487);
or U19814 (N_19814,N_18453,N_18373);
nor U19815 (N_19815,N_18697,N_18287);
xnor U19816 (N_19816,N_18051,N_17964);
xnor U19817 (N_19817,N_18644,N_18117);
xor U19818 (N_19818,N_17684,N_18617);
nand U19819 (N_19819,N_18550,N_18727);
xnor U19820 (N_19820,N_18481,N_17906);
nand U19821 (N_19821,N_17948,N_18734);
nand U19822 (N_19822,N_18085,N_17584);
nor U19823 (N_19823,N_18664,N_18710);
and U19824 (N_19824,N_17800,N_18607);
and U19825 (N_19825,N_17821,N_18066);
nand U19826 (N_19826,N_17672,N_18337);
xor U19827 (N_19827,N_17999,N_18487);
or U19828 (N_19828,N_18589,N_18258);
or U19829 (N_19829,N_17555,N_18707);
xnor U19830 (N_19830,N_18225,N_17718);
and U19831 (N_19831,N_18054,N_18656);
nand U19832 (N_19832,N_17870,N_17711);
nor U19833 (N_19833,N_17689,N_18108);
xnor U19834 (N_19834,N_17927,N_18245);
nor U19835 (N_19835,N_18598,N_18627);
and U19836 (N_19836,N_18259,N_18403);
and U19837 (N_19837,N_18128,N_18571);
and U19838 (N_19838,N_18235,N_17708);
nor U19839 (N_19839,N_17552,N_17765);
nor U19840 (N_19840,N_17887,N_18678);
or U19841 (N_19841,N_17867,N_18400);
nand U19842 (N_19842,N_18243,N_18106);
and U19843 (N_19843,N_18501,N_17600);
and U19844 (N_19844,N_18145,N_17850);
and U19845 (N_19845,N_17989,N_17781);
xor U19846 (N_19846,N_18280,N_18324);
xnor U19847 (N_19847,N_17998,N_18662);
xor U19848 (N_19848,N_18232,N_18460);
nand U19849 (N_19849,N_18678,N_17702);
nor U19850 (N_19850,N_18024,N_18250);
nor U19851 (N_19851,N_18283,N_17530);
xor U19852 (N_19852,N_18658,N_18490);
or U19853 (N_19853,N_17657,N_18609);
xnor U19854 (N_19854,N_18140,N_18331);
nand U19855 (N_19855,N_18098,N_18177);
nor U19856 (N_19856,N_17573,N_17636);
or U19857 (N_19857,N_18178,N_17580);
nand U19858 (N_19858,N_18720,N_18363);
nand U19859 (N_19859,N_17835,N_18678);
nor U19860 (N_19860,N_17948,N_17543);
nor U19861 (N_19861,N_18321,N_18642);
and U19862 (N_19862,N_18174,N_18437);
xor U19863 (N_19863,N_18541,N_18644);
xnor U19864 (N_19864,N_18142,N_18057);
or U19865 (N_19865,N_18168,N_17749);
nor U19866 (N_19866,N_17759,N_18536);
xnor U19867 (N_19867,N_17791,N_18703);
nor U19868 (N_19868,N_18117,N_17817);
and U19869 (N_19869,N_18280,N_17730);
nor U19870 (N_19870,N_18592,N_17652);
nor U19871 (N_19871,N_17931,N_17838);
or U19872 (N_19872,N_18040,N_18522);
xnor U19873 (N_19873,N_18150,N_18574);
xor U19874 (N_19874,N_17790,N_17669);
nor U19875 (N_19875,N_18703,N_18654);
and U19876 (N_19876,N_18484,N_18029);
nor U19877 (N_19877,N_18220,N_18637);
nor U19878 (N_19878,N_17608,N_17512);
or U19879 (N_19879,N_17781,N_17553);
nor U19880 (N_19880,N_17987,N_18226);
xor U19881 (N_19881,N_18698,N_17766);
nor U19882 (N_19882,N_18027,N_18132);
and U19883 (N_19883,N_17875,N_18402);
nor U19884 (N_19884,N_17901,N_18093);
xor U19885 (N_19885,N_18445,N_17870);
nand U19886 (N_19886,N_17521,N_17628);
xor U19887 (N_19887,N_18634,N_18366);
nand U19888 (N_19888,N_18703,N_17849);
or U19889 (N_19889,N_18585,N_18429);
nand U19890 (N_19890,N_18302,N_17594);
xor U19891 (N_19891,N_17773,N_17750);
nor U19892 (N_19892,N_18184,N_18102);
or U19893 (N_19893,N_17918,N_18737);
or U19894 (N_19894,N_17904,N_17653);
and U19895 (N_19895,N_18092,N_18233);
and U19896 (N_19896,N_17828,N_18510);
and U19897 (N_19897,N_18703,N_17534);
or U19898 (N_19898,N_17825,N_18292);
nor U19899 (N_19899,N_17524,N_18586);
xnor U19900 (N_19900,N_18487,N_17798);
xor U19901 (N_19901,N_17516,N_18421);
xnor U19902 (N_19902,N_18266,N_18230);
nor U19903 (N_19903,N_18740,N_18102);
nand U19904 (N_19904,N_18523,N_17751);
nand U19905 (N_19905,N_17866,N_18707);
or U19906 (N_19906,N_18155,N_17930);
or U19907 (N_19907,N_18732,N_17939);
xnor U19908 (N_19908,N_18594,N_18690);
or U19909 (N_19909,N_18171,N_17607);
xor U19910 (N_19910,N_18494,N_18553);
and U19911 (N_19911,N_17866,N_18173);
xor U19912 (N_19912,N_18512,N_17609);
or U19913 (N_19913,N_18063,N_17527);
nand U19914 (N_19914,N_18495,N_18441);
xor U19915 (N_19915,N_17687,N_18149);
xor U19916 (N_19916,N_18553,N_18673);
xnor U19917 (N_19917,N_17942,N_18619);
nand U19918 (N_19918,N_18575,N_17842);
and U19919 (N_19919,N_18210,N_18681);
and U19920 (N_19920,N_18215,N_18284);
nor U19921 (N_19921,N_18567,N_18193);
or U19922 (N_19922,N_17831,N_18627);
or U19923 (N_19923,N_18705,N_18354);
nor U19924 (N_19924,N_18458,N_17592);
nand U19925 (N_19925,N_17624,N_18743);
xnor U19926 (N_19926,N_18255,N_18192);
or U19927 (N_19927,N_17756,N_17847);
or U19928 (N_19928,N_18214,N_17932);
nand U19929 (N_19929,N_17885,N_18229);
nor U19930 (N_19930,N_18086,N_17937);
xor U19931 (N_19931,N_18616,N_18639);
xnor U19932 (N_19932,N_17888,N_18690);
nor U19933 (N_19933,N_17646,N_17617);
nand U19934 (N_19934,N_17556,N_18143);
xnor U19935 (N_19935,N_17665,N_18132);
and U19936 (N_19936,N_18093,N_18163);
nand U19937 (N_19937,N_17558,N_18048);
nor U19938 (N_19938,N_18440,N_18327);
xnor U19939 (N_19939,N_18440,N_18426);
nor U19940 (N_19940,N_18186,N_18352);
nand U19941 (N_19941,N_18566,N_18723);
xor U19942 (N_19942,N_17763,N_17944);
or U19943 (N_19943,N_17622,N_17714);
and U19944 (N_19944,N_18726,N_18053);
nand U19945 (N_19945,N_18321,N_18594);
nor U19946 (N_19946,N_18714,N_17821);
or U19947 (N_19947,N_18283,N_17929);
and U19948 (N_19948,N_18351,N_18120);
nand U19949 (N_19949,N_18044,N_18431);
and U19950 (N_19950,N_18279,N_17560);
or U19951 (N_19951,N_18574,N_18701);
and U19952 (N_19952,N_17798,N_18663);
nor U19953 (N_19953,N_17972,N_17921);
nand U19954 (N_19954,N_18570,N_17733);
nor U19955 (N_19955,N_17506,N_17684);
nor U19956 (N_19956,N_17552,N_18266);
or U19957 (N_19957,N_18695,N_17806);
and U19958 (N_19958,N_17854,N_18100);
or U19959 (N_19959,N_17759,N_18228);
and U19960 (N_19960,N_18352,N_18453);
and U19961 (N_19961,N_18683,N_18411);
and U19962 (N_19962,N_18399,N_18697);
or U19963 (N_19963,N_18467,N_18357);
nand U19964 (N_19964,N_18300,N_17511);
and U19965 (N_19965,N_18649,N_17584);
xnor U19966 (N_19966,N_17586,N_18345);
nor U19967 (N_19967,N_18029,N_17995);
nand U19968 (N_19968,N_18174,N_18588);
and U19969 (N_19969,N_18132,N_18321);
or U19970 (N_19970,N_18195,N_18448);
xor U19971 (N_19971,N_18719,N_17890);
nand U19972 (N_19972,N_18677,N_17597);
and U19973 (N_19973,N_17604,N_18363);
nor U19974 (N_19974,N_18453,N_18401);
and U19975 (N_19975,N_18327,N_17720);
xnor U19976 (N_19976,N_18682,N_17838);
and U19977 (N_19977,N_17961,N_18119);
nand U19978 (N_19978,N_17519,N_17615);
and U19979 (N_19979,N_18233,N_18392);
xor U19980 (N_19980,N_17778,N_18142);
nand U19981 (N_19981,N_17790,N_18391);
and U19982 (N_19982,N_18742,N_17699);
nand U19983 (N_19983,N_18548,N_18634);
xnor U19984 (N_19984,N_18310,N_17916);
and U19985 (N_19985,N_18044,N_17751);
xor U19986 (N_19986,N_17909,N_18019);
nor U19987 (N_19987,N_17791,N_18391);
or U19988 (N_19988,N_18296,N_18570);
nand U19989 (N_19989,N_18376,N_18473);
nor U19990 (N_19990,N_17959,N_17772);
nor U19991 (N_19991,N_18304,N_17999);
and U19992 (N_19992,N_18402,N_17739);
and U19993 (N_19993,N_18057,N_18648);
xnor U19994 (N_19994,N_18171,N_18042);
and U19995 (N_19995,N_18153,N_17651);
or U19996 (N_19996,N_18631,N_17702);
nand U19997 (N_19997,N_18592,N_17994);
or U19998 (N_19998,N_17780,N_17994);
and U19999 (N_19999,N_17794,N_17901);
and U20000 (N_20000,N_19102,N_18964);
nor U20001 (N_20001,N_19080,N_19321);
or U20002 (N_20002,N_18795,N_19050);
nand U20003 (N_20003,N_19827,N_19900);
and U20004 (N_20004,N_19870,N_19352);
and U20005 (N_20005,N_19366,N_19519);
nor U20006 (N_20006,N_18948,N_19271);
and U20007 (N_20007,N_18918,N_19540);
nor U20008 (N_20008,N_19190,N_19318);
xor U20009 (N_20009,N_19263,N_19220);
nand U20010 (N_20010,N_18826,N_19511);
or U20011 (N_20011,N_19162,N_19226);
nor U20012 (N_20012,N_19430,N_18860);
and U20013 (N_20013,N_18876,N_19817);
or U20014 (N_20014,N_19360,N_18784);
and U20015 (N_20015,N_18898,N_19811);
and U20016 (N_20016,N_19041,N_19640);
nor U20017 (N_20017,N_19347,N_19187);
nand U20018 (N_20018,N_19735,N_18956);
nor U20019 (N_20019,N_19335,N_18854);
or U20020 (N_20020,N_19393,N_19935);
nor U20021 (N_20021,N_19128,N_19895);
and U20022 (N_20022,N_18924,N_19867);
or U20023 (N_20023,N_19968,N_18996);
and U20024 (N_20024,N_19259,N_19548);
and U20025 (N_20025,N_18851,N_19500);
and U20026 (N_20026,N_18940,N_19490);
or U20027 (N_20027,N_19242,N_18849);
and U20028 (N_20028,N_19921,N_19672);
nor U20029 (N_20029,N_19876,N_19576);
nor U20030 (N_20030,N_19937,N_19032);
or U20031 (N_20031,N_18847,N_19744);
or U20032 (N_20032,N_19552,N_19353);
and U20033 (N_20033,N_19378,N_19067);
xnor U20034 (N_20034,N_18926,N_19916);
and U20035 (N_20035,N_19238,N_19816);
nand U20036 (N_20036,N_19083,N_19905);
xor U20037 (N_20037,N_19699,N_19858);
nor U20038 (N_20038,N_19855,N_19244);
nor U20039 (N_20039,N_18885,N_18982);
nand U20040 (N_20040,N_19336,N_19790);
nor U20041 (N_20041,N_19865,N_19773);
nor U20042 (N_20042,N_19119,N_18962);
or U20043 (N_20043,N_19651,N_19704);
nand U20044 (N_20044,N_18821,N_19230);
nand U20045 (N_20045,N_19141,N_19369);
and U20046 (N_20046,N_19068,N_19303);
or U20047 (N_20047,N_19301,N_19415);
nor U20048 (N_20048,N_19154,N_19554);
nand U20049 (N_20049,N_19262,N_19587);
and U20050 (N_20050,N_19962,N_19583);
nand U20051 (N_20051,N_19908,N_19869);
nor U20052 (N_20052,N_19240,N_18949);
nand U20053 (N_20053,N_19581,N_19355);
xnor U20054 (N_20054,N_19175,N_19326);
nor U20055 (N_20055,N_19887,N_19974);
xor U20056 (N_20056,N_19470,N_19088);
or U20057 (N_20057,N_19372,N_19086);
xor U20058 (N_20058,N_18978,N_19542);
or U20059 (N_20059,N_19479,N_19243);
xor U20060 (N_20060,N_19523,N_19342);
or U20061 (N_20061,N_19024,N_19623);
or U20062 (N_20062,N_19434,N_19433);
and U20063 (N_20063,N_19034,N_19108);
nor U20064 (N_20064,N_19718,N_19823);
or U20065 (N_20065,N_19142,N_19498);
or U20066 (N_20066,N_18803,N_19401);
nand U20067 (N_20067,N_19406,N_19105);
and U20068 (N_20068,N_19466,N_19741);
nor U20069 (N_20069,N_19755,N_18779);
nand U20070 (N_20070,N_18767,N_19530);
and U20071 (N_20071,N_18910,N_19103);
xnor U20072 (N_20072,N_18947,N_18959);
or U20073 (N_20073,N_18950,N_19345);
nand U20074 (N_20074,N_19517,N_19566);
or U20075 (N_20075,N_19666,N_19524);
xnor U20076 (N_20076,N_18764,N_19099);
and U20077 (N_20077,N_19450,N_18961);
xor U20078 (N_20078,N_19201,N_19348);
and U20079 (N_20079,N_19743,N_19012);
nand U20080 (N_20080,N_19821,N_19632);
and U20081 (N_20081,N_19997,N_19953);
xor U20082 (N_20082,N_19714,N_19673);
nand U20083 (N_20083,N_19081,N_19197);
xor U20084 (N_20084,N_19987,N_19915);
nand U20085 (N_20085,N_19904,N_19487);
or U20086 (N_20086,N_19385,N_19489);
or U20087 (N_20087,N_18966,N_19638);
xnor U20088 (N_20088,N_19733,N_19996);
nand U20089 (N_20089,N_19531,N_19155);
nor U20090 (N_20090,N_18832,N_19562);
nor U20091 (N_20091,N_19590,N_19747);
nor U20092 (N_20092,N_19693,N_19398);
or U20093 (N_20093,N_19338,N_19302);
nand U20094 (N_20094,N_18893,N_19943);
and U20095 (N_20095,N_19717,N_19216);
nor U20096 (N_20096,N_19859,N_19346);
nand U20097 (N_20097,N_19465,N_18807);
nand U20098 (N_20098,N_19341,N_18873);
nand U20099 (N_20099,N_19866,N_19443);
or U20100 (N_20100,N_19715,N_18823);
or U20101 (N_20101,N_19092,N_18973);
or U20102 (N_20102,N_19025,N_19655);
or U20103 (N_20103,N_19309,N_19028);
and U20104 (N_20104,N_19290,N_19113);
and U20105 (N_20105,N_19471,N_18886);
nand U20106 (N_20106,N_18867,N_19316);
and U20107 (N_20107,N_18974,N_18925);
xor U20108 (N_20108,N_19826,N_19245);
xor U20109 (N_20109,N_19351,N_19188);
xor U20110 (N_20110,N_18993,N_18912);
nor U20111 (N_20111,N_19898,N_19782);
xor U20112 (N_20112,N_19624,N_19793);
or U20113 (N_20113,N_19875,N_19535);
nor U20114 (N_20114,N_19284,N_19629);
and U20115 (N_20115,N_18987,N_19365);
xnor U20116 (N_20116,N_19927,N_19759);
and U20117 (N_20117,N_19878,N_19986);
xor U20118 (N_20118,N_19789,N_19634);
xnor U20119 (N_20119,N_18916,N_19973);
nor U20120 (N_20120,N_19438,N_18887);
or U20121 (N_20121,N_19368,N_19204);
nor U20122 (N_20122,N_19662,N_18980);
xnor U20123 (N_20123,N_18889,N_19384);
nand U20124 (N_20124,N_18969,N_18985);
nor U20125 (N_20125,N_18880,N_19971);
nand U20126 (N_20126,N_18883,N_19594);
and U20127 (N_20127,N_19277,N_19757);
xor U20128 (N_20128,N_19665,N_19250);
nand U20129 (N_20129,N_18968,N_19173);
or U20130 (N_20130,N_19070,N_19392);
nor U20131 (N_20131,N_19998,N_18894);
nor U20132 (N_20132,N_19445,N_18967);
and U20133 (N_20133,N_19031,N_18776);
nor U20134 (N_20134,N_19006,N_19745);
xnor U20135 (N_20135,N_19224,N_19502);
or U20136 (N_20136,N_19044,N_19558);
nor U20137 (N_20137,N_19258,N_19791);
and U20138 (N_20138,N_19181,N_19178);
and U20139 (N_20139,N_19721,N_19425);
or U20140 (N_20140,N_19657,N_19950);
or U20141 (N_20141,N_19192,N_19538);
xnor U20142 (N_20142,N_19059,N_19215);
nor U20143 (N_20143,N_19320,N_19681);
nor U20144 (N_20144,N_19608,N_19850);
nor U20145 (N_20145,N_19480,N_19809);
xor U20146 (N_20146,N_19712,N_19003);
nor U20147 (N_20147,N_19628,N_18970);
and U20148 (N_20148,N_19196,N_19289);
nor U20149 (N_20149,N_19097,N_19537);
nand U20150 (N_20150,N_19136,N_18919);
nand U20151 (N_20151,N_19846,N_19127);
nor U20152 (N_20152,N_18900,N_19988);
and U20153 (N_20153,N_18899,N_19222);
nand U20154 (N_20154,N_19169,N_19779);
or U20155 (N_20155,N_19602,N_19093);
nor U20156 (N_20156,N_19007,N_19004);
xor U20157 (N_20157,N_19993,N_19476);
or U20158 (N_20158,N_19896,N_19929);
nor U20159 (N_20159,N_19209,N_18976);
or U20160 (N_20160,N_18763,N_19061);
and U20161 (N_20161,N_19435,N_19112);
or U20162 (N_20162,N_19256,N_19146);
and U20163 (N_20163,N_19970,N_19952);
or U20164 (N_20164,N_19229,N_19379);
and U20165 (N_20165,N_18802,N_19404);
or U20166 (N_20166,N_19899,N_19884);
and U20167 (N_20167,N_19926,N_19567);
or U20168 (N_20168,N_18778,N_19674);
nor U20169 (N_20169,N_19444,N_19189);
and U20170 (N_20170,N_19765,N_19736);
xnor U20171 (N_20171,N_19893,N_18853);
nand U20172 (N_20172,N_18935,N_19491);
or U20173 (N_20173,N_19446,N_18836);
or U20174 (N_20174,N_19218,N_19436);
nand U20175 (N_20175,N_19930,N_19292);
and U20176 (N_20176,N_19056,N_19701);
nand U20177 (N_20177,N_19603,N_19889);
or U20178 (N_20178,N_19231,N_18822);
and U20179 (N_20179,N_19270,N_19668);
and U20180 (N_20180,N_18951,N_19076);
nand U20181 (N_20181,N_19453,N_19417);
nand U20182 (N_20182,N_19077,N_18874);
and U20183 (N_20183,N_18942,N_19903);
and U20184 (N_20184,N_19268,N_19233);
nand U20185 (N_20185,N_19688,N_19239);
nand U20186 (N_20186,N_19257,N_19891);
or U20187 (N_20187,N_19000,N_19002);
nand U20188 (N_20188,N_19052,N_19315);
or U20189 (N_20189,N_18769,N_19575);
or U20190 (N_20190,N_18988,N_19545);
nor U20191 (N_20191,N_19650,N_18788);
xnor U20192 (N_20192,N_19664,N_18932);
nor U20193 (N_20193,N_19473,N_19593);
nand U20194 (N_20194,N_19026,N_19123);
nand U20195 (N_20195,N_19913,N_19225);
or U20196 (N_20196,N_19199,N_18891);
nor U20197 (N_20197,N_19994,N_19685);
nand U20198 (N_20198,N_18813,N_19788);
nand U20199 (N_20199,N_18793,N_19403);
nand U20200 (N_20200,N_19265,N_19675);
or U20201 (N_20201,N_19011,N_18920);
xnor U20202 (N_20202,N_19472,N_19228);
xor U20203 (N_20203,N_19330,N_18859);
nand U20204 (N_20204,N_19932,N_19496);
nand U20205 (N_20205,N_19768,N_19104);
or U20206 (N_20206,N_19084,N_19754);
xnor U20207 (N_20207,N_18998,N_19340);
nor U20208 (N_20208,N_19048,N_19276);
or U20209 (N_20209,N_19588,N_19247);
xnor U20210 (N_20210,N_19122,N_19098);
xnor U20211 (N_20211,N_19095,N_19163);
and U20212 (N_20212,N_19728,N_19945);
nor U20213 (N_20213,N_18986,N_19582);
or U20214 (N_20214,N_19854,N_19770);
nor U20215 (N_20215,N_19047,N_19621);
xnor U20216 (N_20216,N_18991,N_19515);
nor U20217 (N_20217,N_19591,N_19864);
and U20218 (N_20218,N_19419,N_19038);
nand U20219 (N_20219,N_19138,N_19022);
nand U20220 (N_20220,N_19264,N_19604);
xnor U20221 (N_20221,N_19422,N_19800);
nor U20222 (N_20222,N_19750,N_19710);
nor U20223 (N_20223,N_19615,N_19559);
or U20224 (N_20224,N_18852,N_19729);
and U20225 (N_20225,N_19328,N_19058);
and U20226 (N_20226,N_19395,N_19079);
nand U20227 (N_20227,N_19111,N_19692);
nor U20228 (N_20228,N_19475,N_19663);
xnor U20229 (N_20229,N_19758,N_19839);
and U20230 (N_20230,N_18827,N_19881);
or U20231 (N_20231,N_18914,N_19402);
and U20232 (N_20232,N_19888,N_19234);
or U20233 (N_20233,N_19090,N_19172);
nand U20234 (N_20234,N_19117,N_19574);
xnor U20235 (N_20235,N_18936,N_19280);
and U20236 (N_20236,N_19543,N_19984);
and U20237 (N_20237,N_18865,N_19771);
and U20238 (N_20238,N_18820,N_19956);
nand U20239 (N_20239,N_18977,N_19509);
nor U20240 (N_20240,N_19087,N_19795);
nor U20241 (N_20241,N_19357,N_19802);
and U20242 (N_20242,N_19359,N_19397);
or U20243 (N_20243,N_18983,N_19720);
and U20244 (N_20244,N_18957,N_19948);
or U20245 (N_20245,N_19428,N_19001);
or U20246 (N_20246,N_19687,N_18879);
nand U20247 (N_20247,N_19505,N_18917);
nand U20248 (N_20248,N_18750,N_19804);
and U20249 (N_20249,N_19461,N_19920);
and U20250 (N_20250,N_19999,N_19828);
nor U20251 (N_20251,N_19391,N_19849);
xor U20252 (N_20252,N_19462,N_19652);
nand U20253 (N_20253,N_19907,N_18811);
xnor U20254 (N_20254,N_19787,N_19644);
nor U20255 (N_20255,N_19168,N_19705);
nor U20256 (N_20256,N_19620,N_18770);
or U20257 (N_20257,N_18835,N_19483);
or U20258 (N_20258,N_19008,N_19852);
nand U20259 (N_20259,N_19989,N_19570);
and U20260 (N_20260,N_19214,N_18828);
nand U20261 (N_20261,N_19711,N_19286);
nand U20262 (N_20262,N_19622,N_19253);
nor U20263 (N_20263,N_19539,N_18845);
nor U20264 (N_20264,N_19738,N_19860);
and U20265 (N_20265,N_19957,N_19585);
or U20266 (N_20266,N_19868,N_19317);
nor U20267 (N_20267,N_19798,N_18955);
or U20268 (N_20268,N_19641,N_19333);
and U20269 (N_20269,N_19296,N_19626);
xor U20270 (N_20270,N_19153,N_19746);
and U20271 (N_20271,N_18801,N_19383);
and U20272 (N_20272,N_19703,N_19769);
xor U20273 (N_20273,N_19390,N_19260);
and U20274 (N_20274,N_19844,N_19775);
and U20275 (N_20275,N_19293,N_19497);
nand U20276 (N_20276,N_19825,N_19246);
xnor U20277 (N_20277,N_19100,N_19646);
nand U20278 (N_20278,N_19958,N_19808);
nor U20279 (N_20279,N_18830,N_19504);
xor U20280 (N_20280,N_19017,N_19394);
xor U20281 (N_20281,N_19033,N_19167);
nor U20282 (N_20282,N_18752,N_19579);
and U20283 (N_20283,N_19835,N_19429);
or U20284 (N_20284,N_19931,N_19845);
and U20285 (N_20285,N_19563,N_19707);
and U20286 (N_20286,N_18785,N_19812);
nand U20287 (N_20287,N_18971,N_18902);
and U20288 (N_20288,N_19255,N_19857);
xnor U20289 (N_20289,N_19492,N_19906);
or U20290 (N_20290,N_19577,N_19124);
or U20291 (N_20291,N_19306,N_19556);
xor U20292 (N_20292,N_19831,N_18884);
nor U20293 (N_20293,N_18923,N_19269);
or U20294 (N_20294,N_19521,N_19294);
nand U20295 (N_20295,N_19129,N_19427);
nand U20296 (N_20296,N_19902,N_19980);
xnor U20297 (N_20297,N_19376,N_19726);
xnor U20298 (N_20298,N_19308,N_19132);
xnor U20299 (N_20299,N_19514,N_19633);
or U20300 (N_20300,N_18848,N_19740);
xnor U20301 (N_20301,N_19202,N_18938);
nor U20302 (N_20302,N_18759,N_19659);
xnor U20303 (N_20303,N_19995,N_19251);
and U20304 (N_20304,N_19323,N_19761);
and U20305 (N_20305,N_19021,N_19085);
nand U20306 (N_20306,N_19396,N_19416);
or U20307 (N_20307,N_18979,N_19830);
nand U20308 (N_20308,N_19358,N_19571);
xor U20309 (N_20309,N_18773,N_19182);
nand U20310 (N_20310,N_19314,N_18943);
nand U20311 (N_20311,N_19503,N_19334);
nand U20312 (N_20312,N_19049,N_19065);
or U20313 (N_20313,N_19546,N_18846);
xor U20314 (N_20314,N_19171,N_19299);
nor U20315 (N_20315,N_19518,N_18929);
nand U20316 (N_20316,N_19612,N_19046);
xnor U20317 (N_20317,N_19727,N_19607);
nand U20318 (N_20318,N_19964,N_19606);
or U20319 (N_20319,N_19933,N_18995);
nor U20320 (N_20320,N_19520,N_19671);
xnor U20321 (N_20321,N_19170,N_19580);
or U20322 (N_20322,N_19670,N_19990);
or U20323 (N_20323,N_18843,N_18870);
nor U20324 (N_20324,N_19039,N_19135);
nand U20325 (N_20325,N_19074,N_19073);
xnor U20326 (N_20326,N_18877,N_18939);
nand U20327 (N_20327,N_19840,N_19227);
or U20328 (N_20328,N_19649,N_19512);
nand U20329 (N_20329,N_18922,N_19824);
and U20330 (N_20330,N_19423,N_19985);
nor U20331 (N_20331,N_19658,N_19506);
or U20332 (N_20332,N_19695,N_19847);
nand U20333 (N_20333,N_19249,N_19861);
nand U20334 (N_20334,N_19078,N_19619);
and U20335 (N_20335,N_19753,N_18799);
or U20336 (N_20336,N_19448,N_19572);
nand U20337 (N_20337,N_19942,N_18800);
and U20338 (N_20338,N_19731,N_19149);
and U20339 (N_20339,N_18765,N_19329);
or U20340 (N_20340,N_19459,N_18897);
or U20341 (N_20341,N_18782,N_19778);
nor U20342 (N_20342,N_19709,N_19139);
or U20343 (N_20343,N_19837,N_19918);
and U20344 (N_20344,N_19478,N_19424);
xor U20345 (N_20345,N_19040,N_19356);
nor U20346 (N_20346,N_19069,N_19130);
or U20347 (N_20347,N_19797,N_19118);
and U20348 (N_20348,N_19045,N_18818);
nor U20349 (N_20349,N_18812,N_19116);
or U20350 (N_20350,N_19210,N_19643);
nand U20351 (N_20351,N_18994,N_18907);
nand U20352 (N_20352,N_19669,N_19454);
xnor U20353 (N_20353,N_19730,N_19421);
or U20354 (N_20354,N_18755,N_18871);
and U20355 (N_20355,N_19557,N_18850);
nand U20356 (N_20356,N_18958,N_19035);
xor U20357 (N_20357,N_19057,N_19439);
and U20358 (N_20358,N_19151,N_18927);
xnor U20359 (N_20359,N_19617,N_18796);
xnor U20360 (N_20360,N_19982,N_19555);
xor U20361 (N_20361,N_18774,N_19803);
nor U20362 (N_20362,N_19873,N_19332);
xnor U20363 (N_20363,N_19786,N_19613);
xor U20364 (N_20364,N_19946,N_19568);
xor U20365 (N_20365,N_19614,N_19109);
or U20366 (N_20366,N_19179,N_18808);
or U20367 (N_20367,N_19322,N_18839);
and U20368 (N_20368,N_19781,N_19185);
xnor U20369 (N_20369,N_19922,N_19654);
and U20370 (N_20370,N_19560,N_19221);
or U20371 (N_20371,N_19460,N_18760);
xor U20372 (N_20372,N_19295,N_19550);
or U20373 (N_20373,N_19140,N_19618);
nand U20374 (N_20374,N_18933,N_19955);
and U20375 (N_20375,N_19300,N_18772);
nand U20376 (N_20376,N_19683,N_19969);
xnor U20377 (N_20377,N_19451,N_18913);
and U20378 (N_20378,N_18863,N_19051);
nor U20379 (N_20379,N_19125,N_19637);
or U20380 (N_20380,N_19205,N_18999);
or U20381 (N_20381,N_19018,N_19036);
nand U20382 (N_20382,N_19785,N_19311);
and U20383 (N_20383,N_19133,N_19508);
nand U20384 (N_20384,N_19679,N_19213);
nor U20385 (N_20385,N_19331,N_19194);
nand U20386 (N_20386,N_19883,N_19019);
or U20387 (N_20387,N_19014,N_19941);
nand U20388 (N_20388,N_19507,N_19157);
or U20389 (N_20389,N_18780,N_19967);
and U20390 (N_20390,N_19596,N_18963);
and U20391 (N_20391,N_19647,N_19174);
nor U20392 (N_20392,N_19183,N_19541);
nor U20393 (N_20393,N_19807,N_19949);
or U20394 (N_20394,N_19690,N_19836);
and U20395 (N_20395,N_19241,N_19925);
or U20396 (N_20396,N_19337,N_19408);
xor U20397 (N_20397,N_19400,N_18965);
xnor U20398 (N_20398,N_19371,N_18794);
or U20399 (N_20399,N_18946,N_19186);
and U20400 (N_20400,N_19879,N_18869);
nand U20401 (N_20401,N_19616,N_19737);
nand U20402 (N_20402,N_18931,N_19983);
nand U20403 (N_20403,N_19200,N_18882);
nand U20404 (N_20404,N_19121,N_19834);
xnor U20405 (N_20405,N_19732,N_19410);
nor U20406 (N_20406,N_19600,N_18783);
nor U20407 (N_20407,N_19660,N_19965);
nand U20408 (N_20408,N_18903,N_19147);
or U20409 (N_20409,N_18901,N_19776);
xor U20410 (N_20410,N_19248,N_18798);
and U20411 (N_20411,N_19193,N_19015);
and U20412 (N_20412,N_19283,N_19742);
or U20413 (N_20413,N_19842,N_18944);
and U20414 (N_20414,N_19960,N_19437);
nor U20415 (N_20415,N_19464,N_19431);
nor U20416 (N_20416,N_19474,N_19091);
nand U20417 (N_20417,N_19164,N_18814);
xor U20418 (N_20418,N_19783,N_19344);
xnor U20419 (N_20419,N_19938,N_19959);
or U20420 (N_20420,N_18888,N_19592);
nor U20421 (N_20421,N_19288,N_19534);
nor U20422 (N_20422,N_19784,N_19305);
xnor U20423 (N_20423,N_19885,N_19739);
or U20424 (N_20424,N_19037,N_18766);
xor U20425 (N_20425,N_19976,N_18781);
and U20426 (N_20426,N_19029,N_18840);
nand U20427 (N_20427,N_19691,N_19533);
xor U20428 (N_20428,N_18930,N_19274);
xor U20429 (N_20429,N_19206,N_19578);
and U20430 (N_20430,N_19426,N_19405);
xor U20431 (N_20431,N_18824,N_19605);
nand U20432 (N_20432,N_18857,N_19635);
nand U20433 (N_20433,N_19380,N_19697);
nor U20434 (N_20434,N_19934,N_19528);
nor U20435 (N_20435,N_19447,N_19413);
nor U20436 (N_20436,N_19066,N_19853);
nand U20437 (N_20437,N_19696,N_18909);
xor U20438 (N_20438,N_19682,N_19180);
nand U20439 (N_20439,N_19648,N_19752);
or U20440 (N_20440,N_19777,N_18945);
nand U20441 (N_20441,N_19304,N_19748);
nor U20442 (N_20442,N_19477,N_19107);
nand U20443 (N_20443,N_19734,N_18833);
nor U20444 (N_20444,N_18997,N_19805);
nand U20445 (N_20445,N_19799,N_19680);
and U20446 (N_20446,N_19254,N_19838);
nand U20447 (N_20447,N_19463,N_19547);
nor U20448 (N_20448,N_18751,N_19219);
nor U20449 (N_20449,N_19525,N_19645);
and U20450 (N_20450,N_18858,N_19005);
or U20451 (N_20451,N_19526,N_19820);
nor U20452 (N_20452,N_19325,N_19882);
or U20453 (N_20453,N_19678,N_18953);
nor U20454 (N_20454,N_19467,N_18792);
nand U20455 (N_20455,N_19420,N_19856);
xor U20456 (N_20456,N_19706,N_19832);
xnor U20457 (N_20457,N_18804,N_18834);
nand U20458 (N_20458,N_18906,N_19549);
or U20459 (N_20459,N_18805,N_19106);
nand U20460 (N_20460,N_18758,N_18791);
and U20461 (N_20461,N_18989,N_19414);
nor U20462 (N_20462,N_19126,N_19252);
xor U20463 (N_20463,N_19829,N_19917);
and U20464 (N_20464,N_19708,N_18904);
and U20465 (N_20465,N_19966,N_19412);
and U20466 (N_20466,N_19909,N_19944);
or U20467 (N_20467,N_19488,N_19862);
xnor U20468 (N_20468,N_19716,N_18815);
nand U20469 (N_20469,N_19458,N_19702);
nor U20470 (N_20470,N_19774,N_19236);
nand U20471 (N_20471,N_18864,N_19940);
and U20472 (N_20472,N_19851,N_18838);
xnor U20473 (N_20473,N_19055,N_19924);
or U20474 (N_20474,N_19661,N_18875);
nor U20475 (N_20475,N_19364,N_19725);
nor U20476 (N_20476,N_19114,N_19527);
nand U20477 (N_20477,N_19610,N_19016);
xnor U20478 (N_20478,N_19096,N_19792);
nor U20479 (N_20479,N_19894,N_19760);
nor U20480 (N_20480,N_18844,N_19310);
xor U20481 (N_20481,N_19597,N_19386);
nor U20482 (N_20482,N_19382,N_19780);
and U20483 (N_20483,N_18809,N_18757);
and U20484 (N_20484,N_19493,N_19367);
and U20485 (N_20485,N_18928,N_19134);
nand U20486 (N_20486,N_18866,N_19486);
nand U20487 (N_20487,N_19598,N_19806);
nand U20488 (N_20488,N_19569,N_19684);
or U20489 (N_20489,N_19027,N_19631);
xor U20490 (N_20490,N_19979,N_19232);
and U20491 (N_20491,N_19810,N_18753);
and U20492 (N_20492,N_19553,N_19963);
nor U20493 (N_20493,N_18829,N_19159);
nor U20494 (N_20494,N_18789,N_19625);
and U20495 (N_20495,N_19686,N_18896);
and U20496 (N_20496,N_18855,N_19137);
and U20497 (N_20497,N_19601,N_19217);
and U20498 (N_20498,N_19282,N_19818);
xnor U20499 (N_20499,N_19307,N_19455);
nor U20500 (N_20500,N_19064,N_19407);
or U20501 (N_20501,N_19897,N_19452);
nand U20502 (N_20502,N_19235,N_18762);
nor U20503 (N_20503,N_18816,N_19266);
xor U20504 (N_20504,N_19072,N_19319);
and U20505 (N_20505,N_18756,N_19872);
xnor U20506 (N_20506,N_19919,N_18981);
and U20507 (N_20507,N_19532,N_19813);
nor U20508 (N_20508,N_19501,N_19143);
xnor U20509 (N_20509,N_19279,N_19544);
xnor U20510 (N_20510,N_18841,N_19536);
nand U20511 (N_20511,N_19992,N_19212);
xor U20512 (N_20512,N_19339,N_19261);
xor U20513 (N_20513,N_19054,N_19767);
nand U20514 (N_20514,N_19794,N_19009);
nand U20515 (N_20515,N_19723,N_19165);
nor U20516 (N_20516,N_19495,N_19120);
and U20517 (N_20517,N_19981,N_19298);
and U20518 (N_20518,N_18941,N_19287);
nand U20519 (N_20519,N_19203,N_19374);
nand U20520 (N_20520,N_18861,N_19529);
nand U20521 (N_20521,N_19485,N_18819);
nand U20522 (N_20522,N_19694,N_19890);
nor U20523 (N_20523,N_18895,N_19101);
and U20524 (N_20524,N_19561,N_19237);
and U20525 (N_20525,N_19469,N_18992);
nand U20526 (N_20526,N_19698,N_18984);
xnor U20527 (N_20527,N_18960,N_19564);
nor U20528 (N_20528,N_19833,N_19184);
nor U20529 (N_20529,N_19978,N_18890);
nand U20530 (N_20530,N_18972,N_19551);
nor U20531 (N_20531,N_19763,N_19375);
nor U20532 (N_20532,N_19145,N_19363);
nand U20533 (N_20533,N_19354,N_19874);
nand U20534 (N_20534,N_19060,N_19312);
and U20535 (N_20535,N_19766,N_19043);
xor U20536 (N_20536,N_19131,N_19667);
xnor U20537 (N_20537,N_19177,N_18881);
nor U20538 (N_20538,N_18817,N_19158);
nand U20539 (N_20539,N_18934,N_19432);
or U20540 (N_20540,N_18908,N_19161);
or U20541 (N_20541,N_19972,N_18761);
or U20542 (N_20542,N_19627,N_19042);
nand U20543 (N_20543,N_19749,N_19063);
and U20544 (N_20544,N_19499,N_19272);
or U20545 (N_20545,N_19267,N_19841);
xnor U20546 (N_20546,N_19150,N_19910);
nor U20547 (N_20547,N_18937,N_19822);
nand U20548 (N_20548,N_19814,N_19947);
or U20549 (N_20549,N_19457,N_18786);
and U20550 (N_20550,N_19291,N_19208);
nor U20551 (N_20551,N_18825,N_19089);
and U20552 (N_20552,N_19565,N_19751);
or U20553 (N_20553,N_19494,N_19075);
or U20554 (N_20554,N_19442,N_19361);
and U20555 (N_20555,N_19689,N_19642);
nand U20556 (N_20556,N_19418,N_19327);
nor U20557 (N_20557,N_19343,N_19848);
nand U20558 (N_20558,N_19722,N_19901);
and U20559 (N_20559,N_18856,N_19991);
nand U20560 (N_20560,N_19440,N_18837);
nor U20561 (N_20561,N_18797,N_19062);
nor U20562 (N_20562,N_19484,N_18915);
xnor U20563 (N_20563,N_19510,N_18831);
nor U20564 (N_20564,N_19456,N_19482);
and U20565 (N_20565,N_19273,N_18954);
or U20566 (N_20566,N_19324,N_18862);
nor U20567 (N_20567,N_19639,N_19522);
or U20568 (N_20568,N_19796,N_18768);
nor U20569 (N_20569,N_19939,N_19819);
nor U20570 (N_20570,N_19772,N_19152);
nand U20571 (N_20571,N_19677,N_19595);
and U20572 (N_20572,N_18990,N_19166);
or U20573 (N_20573,N_19700,N_19144);
nand U20574 (N_20574,N_19815,N_19281);
nand U20575 (N_20575,N_19911,N_19713);
nor U20576 (N_20576,N_19513,N_19441);
and U20577 (N_20577,N_19914,N_19223);
nor U20578 (N_20578,N_19297,N_19912);
xnor U20579 (N_20579,N_19762,N_19030);
xor U20580 (N_20580,N_19954,N_19013);
nor U20581 (N_20581,N_19756,N_19148);
or U20582 (N_20582,N_19370,N_19160);
xnor U20583 (N_20583,N_19676,N_18771);
or U20584 (N_20584,N_18905,N_19801);
or U20585 (N_20585,N_18842,N_18868);
nor U20586 (N_20586,N_19589,N_19719);
and U20587 (N_20587,N_19449,N_19110);
nand U20588 (N_20588,N_18775,N_19020);
xor U20589 (N_20589,N_19880,N_18810);
xor U20590 (N_20590,N_19278,N_19156);
nor U20591 (N_20591,N_19653,N_18790);
nor U20592 (N_20592,N_19481,N_19656);
and U20593 (N_20593,N_19977,N_19389);
or U20594 (N_20594,N_19082,N_19071);
or U20595 (N_20595,N_19115,N_18777);
and U20596 (N_20596,N_19764,N_19285);
nor U20597 (N_20597,N_19468,N_19573);
xnor U20598 (N_20598,N_19387,N_19176);
and U20599 (N_20599,N_19388,N_19362);
nand U20600 (N_20600,N_19599,N_18975);
and U20601 (N_20601,N_19951,N_19961);
or U20602 (N_20602,N_19975,N_18806);
and U20603 (N_20603,N_19871,N_19724);
or U20604 (N_20604,N_19373,N_19381);
nand U20605 (N_20605,N_19207,N_18892);
and U20606 (N_20606,N_18911,N_19609);
or U20607 (N_20607,N_19010,N_19377);
and U20608 (N_20608,N_19313,N_19586);
nand U20609 (N_20609,N_19349,N_19936);
xor U20610 (N_20610,N_19843,N_19877);
or U20611 (N_20611,N_19191,N_19636);
and U20612 (N_20612,N_19584,N_18952);
xor U20613 (N_20613,N_19630,N_18878);
nor U20614 (N_20614,N_19863,N_19023);
nand U20615 (N_20615,N_18754,N_19094);
nand U20616 (N_20616,N_19409,N_19275);
or U20617 (N_20617,N_19516,N_19211);
nor U20618 (N_20618,N_18787,N_19892);
xor U20619 (N_20619,N_19350,N_19195);
and U20620 (N_20620,N_19928,N_19923);
nand U20621 (N_20621,N_18921,N_19399);
and U20622 (N_20622,N_19198,N_18872);
and U20623 (N_20623,N_19611,N_19053);
xor U20624 (N_20624,N_19886,N_19411);
xor U20625 (N_20625,N_19319,N_19084);
xor U20626 (N_20626,N_19975,N_19971);
and U20627 (N_20627,N_19736,N_19774);
nand U20628 (N_20628,N_19872,N_19178);
nand U20629 (N_20629,N_18996,N_19875);
or U20630 (N_20630,N_19531,N_19321);
nor U20631 (N_20631,N_19314,N_19792);
and U20632 (N_20632,N_19045,N_19893);
xnor U20633 (N_20633,N_19990,N_19207);
nor U20634 (N_20634,N_19989,N_18942);
nor U20635 (N_20635,N_19534,N_19696);
nor U20636 (N_20636,N_19796,N_19759);
nor U20637 (N_20637,N_19555,N_18789);
nor U20638 (N_20638,N_19727,N_19047);
xor U20639 (N_20639,N_19165,N_19080);
nor U20640 (N_20640,N_19382,N_19004);
xor U20641 (N_20641,N_19042,N_19078);
or U20642 (N_20642,N_19753,N_19748);
and U20643 (N_20643,N_19634,N_18817);
and U20644 (N_20644,N_19761,N_18955);
and U20645 (N_20645,N_19442,N_19438);
and U20646 (N_20646,N_19627,N_19630);
or U20647 (N_20647,N_19586,N_18800);
xor U20648 (N_20648,N_19397,N_19143);
and U20649 (N_20649,N_18824,N_19418);
nor U20650 (N_20650,N_19904,N_19932);
xor U20651 (N_20651,N_19280,N_19684);
or U20652 (N_20652,N_19761,N_19753);
and U20653 (N_20653,N_19964,N_19862);
and U20654 (N_20654,N_19065,N_19554);
nor U20655 (N_20655,N_19815,N_19208);
and U20656 (N_20656,N_18823,N_19443);
and U20657 (N_20657,N_19054,N_19725);
nor U20658 (N_20658,N_19115,N_19164);
xnor U20659 (N_20659,N_19648,N_19293);
xnor U20660 (N_20660,N_19348,N_19286);
nor U20661 (N_20661,N_18981,N_19802);
or U20662 (N_20662,N_19078,N_19194);
and U20663 (N_20663,N_19277,N_19056);
nand U20664 (N_20664,N_19227,N_18894);
and U20665 (N_20665,N_19496,N_18775);
and U20666 (N_20666,N_18990,N_19422);
nor U20667 (N_20667,N_19241,N_19943);
xnor U20668 (N_20668,N_18775,N_19933);
nor U20669 (N_20669,N_19318,N_19986);
nand U20670 (N_20670,N_19260,N_19815);
xor U20671 (N_20671,N_19599,N_19513);
and U20672 (N_20672,N_19324,N_19520);
and U20673 (N_20673,N_19727,N_19622);
and U20674 (N_20674,N_19304,N_19529);
nand U20675 (N_20675,N_18833,N_19279);
and U20676 (N_20676,N_19659,N_19474);
xor U20677 (N_20677,N_19670,N_18997);
and U20678 (N_20678,N_19392,N_19768);
or U20679 (N_20679,N_19355,N_19667);
nor U20680 (N_20680,N_19504,N_19482);
nand U20681 (N_20681,N_19908,N_19496);
or U20682 (N_20682,N_19811,N_19424);
or U20683 (N_20683,N_19416,N_19436);
nand U20684 (N_20684,N_19890,N_18996);
xor U20685 (N_20685,N_19510,N_18968);
or U20686 (N_20686,N_19663,N_19488);
nand U20687 (N_20687,N_19744,N_19502);
and U20688 (N_20688,N_18784,N_18758);
or U20689 (N_20689,N_19210,N_19186);
and U20690 (N_20690,N_18800,N_19974);
xnor U20691 (N_20691,N_19659,N_19333);
nand U20692 (N_20692,N_19537,N_19397);
nand U20693 (N_20693,N_19134,N_19541);
xnor U20694 (N_20694,N_19202,N_19470);
xnor U20695 (N_20695,N_19475,N_19147);
and U20696 (N_20696,N_19569,N_19852);
xor U20697 (N_20697,N_19203,N_18762);
or U20698 (N_20698,N_19757,N_19519);
nor U20699 (N_20699,N_19768,N_19337);
nand U20700 (N_20700,N_19703,N_18773);
nor U20701 (N_20701,N_18894,N_19675);
nand U20702 (N_20702,N_19252,N_19851);
nand U20703 (N_20703,N_19695,N_19398);
xnor U20704 (N_20704,N_19949,N_19549);
nand U20705 (N_20705,N_19531,N_19433);
nor U20706 (N_20706,N_18878,N_19534);
or U20707 (N_20707,N_19898,N_19119);
xor U20708 (N_20708,N_19894,N_19968);
xnor U20709 (N_20709,N_19267,N_18905);
xor U20710 (N_20710,N_19214,N_18989);
xor U20711 (N_20711,N_19391,N_19283);
and U20712 (N_20712,N_19294,N_19255);
xnor U20713 (N_20713,N_19476,N_19544);
or U20714 (N_20714,N_19575,N_18785);
or U20715 (N_20715,N_19863,N_19625);
nor U20716 (N_20716,N_19092,N_18777);
xor U20717 (N_20717,N_19210,N_19003);
and U20718 (N_20718,N_19238,N_19870);
xor U20719 (N_20719,N_19141,N_19997);
or U20720 (N_20720,N_18773,N_19569);
or U20721 (N_20721,N_18788,N_19776);
nand U20722 (N_20722,N_19033,N_19022);
nor U20723 (N_20723,N_19518,N_19314);
or U20724 (N_20724,N_19475,N_19329);
xnor U20725 (N_20725,N_18784,N_19240);
nor U20726 (N_20726,N_19609,N_19315);
or U20727 (N_20727,N_19948,N_18873);
or U20728 (N_20728,N_19977,N_19585);
nand U20729 (N_20729,N_19605,N_19822);
and U20730 (N_20730,N_19252,N_18968);
nor U20731 (N_20731,N_19119,N_19298);
nand U20732 (N_20732,N_19112,N_19717);
nor U20733 (N_20733,N_19366,N_19760);
and U20734 (N_20734,N_19381,N_19420);
nor U20735 (N_20735,N_19549,N_19127);
nor U20736 (N_20736,N_19242,N_19805);
nor U20737 (N_20737,N_19987,N_18796);
nand U20738 (N_20738,N_18767,N_19141);
and U20739 (N_20739,N_19274,N_19982);
nor U20740 (N_20740,N_18851,N_19225);
or U20741 (N_20741,N_19780,N_19965);
or U20742 (N_20742,N_19724,N_19776);
nor U20743 (N_20743,N_19591,N_19937);
or U20744 (N_20744,N_19457,N_19089);
nand U20745 (N_20745,N_19175,N_19409);
xnor U20746 (N_20746,N_18844,N_18759);
xnor U20747 (N_20747,N_19787,N_19170);
xor U20748 (N_20748,N_19878,N_19305);
or U20749 (N_20749,N_18805,N_18941);
nor U20750 (N_20750,N_19399,N_19819);
xnor U20751 (N_20751,N_19183,N_18905);
xor U20752 (N_20752,N_18764,N_19990);
nor U20753 (N_20753,N_19031,N_19870);
and U20754 (N_20754,N_19014,N_19033);
or U20755 (N_20755,N_19415,N_19916);
and U20756 (N_20756,N_19246,N_19673);
xnor U20757 (N_20757,N_19860,N_19711);
xnor U20758 (N_20758,N_19494,N_19536);
nor U20759 (N_20759,N_18780,N_19629);
and U20760 (N_20760,N_19948,N_19897);
and U20761 (N_20761,N_19939,N_19166);
nand U20762 (N_20762,N_19739,N_19569);
or U20763 (N_20763,N_19677,N_19151);
nand U20764 (N_20764,N_19653,N_18766);
nor U20765 (N_20765,N_19892,N_19297);
and U20766 (N_20766,N_19549,N_18796);
and U20767 (N_20767,N_19007,N_19280);
xnor U20768 (N_20768,N_19273,N_19705);
and U20769 (N_20769,N_19581,N_19122);
nand U20770 (N_20770,N_19739,N_19324);
xor U20771 (N_20771,N_19593,N_19804);
nor U20772 (N_20772,N_19142,N_19603);
nor U20773 (N_20773,N_18835,N_19518);
or U20774 (N_20774,N_19185,N_18994);
nand U20775 (N_20775,N_19098,N_19432);
or U20776 (N_20776,N_19254,N_19408);
nand U20777 (N_20777,N_18822,N_19988);
nand U20778 (N_20778,N_19763,N_18833);
and U20779 (N_20779,N_19371,N_19139);
nor U20780 (N_20780,N_19453,N_19135);
and U20781 (N_20781,N_18789,N_19547);
and U20782 (N_20782,N_19207,N_19969);
nand U20783 (N_20783,N_19350,N_19657);
nand U20784 (N_20784,N_19824,N_19023);
and U20785 (N_20785,N_19706,N_19904);
xor U20786 (N_20786,N_18786,N_18901);
nor U20787 (N_20787,N_19595,N_19513);
xor U20788 (N_20788,N_19953,N_19331);
xnor U20789 (N_20789,N_19064,N_19181);
xor U20790 (N_20790,N_19979,N_19403);
and U20791 (N_20791,N_19884,N_19397);
nand U20792 (N_20792,N_19246,N_19364);
nor U20793 (N_20793,N_19169,N_19383);
and U20794 (N_20794,N_19906,N_19699);
nor U20795 (N_20795,N_18840,N_19374);
xor U20796 (N_20796,N_19418,N_18992);
xnor U20797 (N_20797,N_19835,N_19643);
xnor U20798 (N_20798,N_19222,N_19100);
nand U20799 (N_20799,N_19314,N_19291);
xor U20800 (N_20800,N_19791,N_18835);
nand U20801 (N_20801,N_19684,N_18768);
xnor U20802 (N_20802,N_19327,N_19778);
xor U20803 (N_20803,N_19048,N_19870);
or U20804 (N_20804,N_19823,N_18796);
nor U20805 (N_20805,N_19968,N_19546);
and U20806 (N_20806,N_18936,N_19132);
xor U20807 (N_20807,N_18885,N_19049);
or U20808 (N_20808,N_19237,N_19899);
nor U20809 (N_20809,N_18879,N_19783);
xor U20810 (N_20810,N_19376,N_19174);
or U20811 (N_20811,N_19203,N_18831);
nand U20812 (N_20812,N_18816,N_19565);
nand U20813 (N_20813,N_18818,N_19081);
or U20814 (N_20814,N_19245,N_19046);
nor U20815 (N_20815,N_19882,N_18851);
and U20816 (N_20816,N_19515,N_18825);
and U20817 (N_20817,N_19333,N_19770);
or U20818 (N_20818,N_19923,N_19904);
and U20819 (N_20819,N_19620,N_19468);
and U20820 (N_20820,N_19502,N_19289);
or U20821 (N_20821,N_19492,N_19672);
nand U20822 (N_20822,N_19810,N_18933);
or U20823 (N_20823,N_19293,N_19631);
and U20824 (N_20824,N_19571,N_18763);
nor U20825 (N_20825,N_19469,N_19575);
or U20826 (N_20826,N_19150,N_19398);
nand U20827 (N_20827,N_19677,N_19278);
nor U20828 (N_20828,N_19739,N_19368);
nor U20829 (N_20829,N_19758,N_18982);
or U20830 (N_20830,N_19508,N_18813);
and U20831 (N_20831,N_19777,N_19220);
or U20832 (N_20832,N_19150,N_19863);
xnor U20833 (N_20833,N_19844,N_19949);
or U20834 (N_20834,N_19016,N_19938);
nand U20835 (N_20835,N_19838,N_18826);
nand U20836 (N_20836,N_19373,N_19652);
nand U20837 (N_20837,N_18935,N_19759);
nand U20838 (N_20838,N_19107,N_18914);
or U20839 (N_20839,N_19063,N_19059);
nor U20840 (N_20840,N_19038,N_19012);
and U20841 (N_20841,N_19514,N_18902);
or U20842 (N_20842,N_19718,N_19847);
nand U20843 (N_20843,N_18847,N_18819);
nand U20844 (N_20844,N_19463,N_19303);
xnor U20845 (N_20845,N_19122,N_19220);
xnor U20846 (N_20846,N_19579,N_19561);
nor U20847 (N_20847,N_19919,N_19815);
nand U20848 (N_20848,N_19636,N_19904);
and U20849 (N_20849,N_19728,N_18784);
and U20850 (N_20850,N_19919,N_19082);
or U20851 (N_20851,N_19056,N_19310);
and U20852 (N_20852,N_19502,N_18768);
xor U20853 (N_20853,N_18985,N_19156);
nor U20854 (N_20854,N_19176,N_19824);
nand U20855 (N_20855,N_19684,N_19572);
nand U20856 (N_20856,N_19898,N_19835);
or U20857 (N_20857,N_19094,N_19139);
and U20858 (N_20858,N_19090,N_19911);
or U20859 (N_20859,N_19753,N_19451);
nor U20860 (N_20860,N_19440,N_19004);
and U20861 (N_20861,N_19092,N_19890);
xor U20862 (N_20862,N_19778,N_19192);
xor U20863 (N_20863,N_19879,N_18898);
or U20864 (N_20864,N_19479,N_19914);
nor U20865 (N_20865,N_19147,N_19841);
and U20866 (N_20866,N_19971,N_18766);
nand U20867 (N_20867,N_19693,N_19076);
xor U20868 (N_20868,N_19099,N_19702);
nor U20869 (N_20869,N_19410,N_19931);
and U20870 (N_20870,N_19788,N_19722);
nand U20871 (N_20871,N_19233,N_19853);
nand U20872 (N_20872,N_19027,N_18840);
nand U20873 (N_20873,N_19305,N_19278);
xor U20874 (N_20874,N_19695,N_19352);
nand U20875 (N_20875,N_19397,N_19619);
nor U20876 (N_20876,N_19824,N_19603);
or U20877 (N_20877,N_18962,N_18758);
nand U20878 (N_20878,N_19999,N_19719);
nor U20879 (N_20879,N_18754,N_19377);
nor U20880 (N_20880,N_19410,N_18887);
nand U20881 (N_20881,N_19698,N_18759);
xnor U20882 (N_20882,N_19652,N_19854);
nand U20883 (N_20883,N_19459,N_19349);
nand U20884 (N_20884,N_19089,N_19870);
xnor U20885 (N_20885,N_19827,N_18988);
xor U20886 (N_20886,N_18820,N_19216);
nand U20887 (N_20887,N_18992,N_19868);
xnor U20888 (N_20888,N_19300,N_19079);
nor U20889 (N_20889,N_18753,N_19656);
nor U20890 (N_20890,N_19604,N_19161);
or U20891 (N_20891,N_19983,N_19470);
nor U20892 (N_20892,N_18813,N_18942);
nand U20893 (N_20893,N_19919,N_19759);
nand U20894 (N_20894,N_19803,N_19479);
nor U20895 (N_20895,N_18858,N_18863);
xor U20896 (N_20896,N_18981,N_19782);
nand U20897 (N_20897,N_19614,N_19034);
or U20898 (N_20898,N_19056,N_18814);
and U20899 (N_20899,N_19512,N_19822);
or U20900 (N_20900,N_19567,N_19813);
nor U20901 (N_20901,N_18825,N_19666);
and U20902 (N_20902,N_19759,N_19979);
xnor U20903 (N_20903,N_18856,N_19656);
or U20904 (N_20904,N_19060,N_19434);
xor U20905 (N_20905,N_18904,N_19872);
or U20906 (N_20906,N_18853,N_18802);
nor U20907 (N_20907,N_19763,N_18942);
xor U20908 (N_20908,N_18983,N_19329);
or U20909 (N_20909,N_19494,N_18857);
or U20910 (N_20910,N_19302,N_19224);
nor U20911 (N_20911,N_19992,N_19648);
nor U20912 (N_20912,N_19242,N_19952);
nor U20913 (N_20913,N_19330,N_19415);
or U20914 (N_20914,N_19912,N_19258);
or U20915 (N_20915,N_19465,N_19541);
or U20916 (N_20916,N_19712,N_18816);
and U20917 (N_20917,N_19544,N_19746);
or U20918 (N_20918,N_18861,N_19198);
and U20919 (N_20919,N_19175,N_19023);
xor U20920 (N_20920,N_19887,N_19044);
and U20921 (N_20921,N_19314,N_19981);
and U20922 (N_20922,N_19578,N_19575);
or U20923 (N_20923,N_18771,N_18946);
nor U20924 (N_20924,N_18784,N_19898);
xor U20925 (N_20925,N_18843,N_19336);
xnor U20926 (N_20926,N_18807,N_18752);
or U20927 (N_20927,N_18823,N_19015);
xor U20928 (N_20928,N_19812,N_19890);
nor U20929 (N_20929,N_18895,N_19469);
or U20930 (N_20930,N_19287,N_19870);
nor U20931 (N_20931,N_18955,N_19774);
nor U20932 (N_20932,N_19175,N_19756);
nor U20933 (N_20933,N_19413,N_19287);
or U20934 (N_20934,N_19549,N_19689);
xnor U20935 (N_20935,N_19159,N_19000);
xor U20936 (N_20936,N_19839,N_18916);
or U20937 (N_20937,N_19276,N_19865);
xnor U20938 (N_20938,N_19139,N_18765);
or U20939 (N_20939,N_19512,N_19644);
and U20940 (N_20940,N_19443,N_19643);
or U20941 (N_20941,N_19042,N_19153);
xnor U20942 (N_20942,N_18940,N_18970);
xnor U20943 (N_20943,N_19878,N_19243);
nand U20944 (N_20944,N_18838,N_19681);
or U20945 (N_20945,N_19475,N_19615);
nor U20946 (N_20946,N_19186,N_19993);
and U20947 (N_20947,N_18839,N_19664);
nand U20948 (N_20948,N_19612,N_19137);
and U20949 (N_20949,N_19353,N_19626);
xnor U20950 (N_20950,N_19919,N_19272);
nand U20951 (N_20951,N_19537,N_18902);
nand U20952 (N_20952,N_19824,N_18816);
nand U20953 (N_20953,N_19812,N_19920);
nor U20954 (N_20954,N_19352,N_19009);
and U20955 (N_20955,N_19691,N_19111);
nor U20956 (N_20956,N_18995,N_18907);
nor U20957 (N_20957,N_19530,N_18966);
or U20958 (N_20958,N_19281,N_19895);
nand U20959 (N_20959,N_19485,N_18917);
nand U20960 (N_20960,N_19691,N_19102);
nor U20961 (N_20961,N_19170,N_19570);
nand U20962 (N_20962,N_19262,N_19274);
and U20963 (N_20963,N_19206,N_19174);
nand U20964 (N_20964,N_19579,N_19454);
nor U20965 (N_20965,N_18963,N_18952);
or U20966 (N_20966,N_19855,N_19759);
and U20967 (N_20967,N_19997,N_19097);
nand U20968 (N_20968,N_19258,N_19309);
nand U20969 (N_20969,N_19068,N_18926);
nor U20970 (N_20970,N_19324,N_19853);
xor U20971 (N_20971,N_19736,N_19318);
or U20972 (N_20972,N_19263,N_19989);
xnor U20973 (N_20973,N_18818,N_18908);
xnor U20974 (N_20974,N_18986,N_19349);
nand U20975 (N_20975,N_19017,N_19998);
or U20976 (N_20976,N_19621,N_19000);
nand U20977 (N_20977,N_19364,N_19223);
or U20978 (N_20978,N_19876,N_18841);
xnor U20979 (N_20979,N_19468,N_19289);
nand U20980 (N_20980,N_19448,N_18798);
nor U20981 (N_20981,N_19707,N_19889);
nand U20982 (N_20982,N_19722,N_19313);
xor U20983 (N_20983,N_19913,N_19206);
nor U20984 (N_20984,N_18999,N_19381);
nor U20985 (N_20985,N_19508,N_19833);
or U20986 (N_20986,N_19922,N_19804);
xnor U20987 (N_20987,N_19511,N_18898);
or U20988 (N_20988,N_19440,N_19740);
nand U20989 (N_20989,N_19613,N_19541);
nor U20990 (N_20990,N_19633,N_19077);
or U20991 (N_20991,N_19534,N_19550);
nand U20992 (N_20992,N_19799,N_19667);
or U20993 (N_20993,N_19971,N_19866);
or U20994 (N_20994,N_19014,N_19836);
nor U20995 (N_20995,N_19280,N_19686);
nand U20996 (N_20996,N_19702,N_18995);
and U20997 (N_20997,N_19578,N_18875);
nor U20998 (N_20998,N_19674,N_19057);
nand U20999 (N_20999,N_19494,N_19795);
nor U21000 (N_21000,N_19960,N_18796);
xor U21001 (N_21001,N_19363,N_19849);
nand U21002 (N_21002,N_19600,N_19509);
nand U21003 (N_21003,N_19636,N_18963);
or U21004 (N_21004,N_18763,N_19864);
nor U21005 (N_21005,N_19999,N_19667);
nand U21006 (N_21006,N_19291,N_19135);
and U21007 (N_21007,N_19424,N_18987);
and U21008 (N_21008,N_18975,N_18964);
and U21009 (N_21009,N_19718,N_19434);
and U21010 (N_21010,N_18767,N_19600);
xor U21011 (N_21011,N_18857,N_19146);
and U21012 (N_21012,N_19406,N_19296);
xor U21013 (N_21013,N_19034,N_19601);
nor U21014 (N_21014,N_19920,N_19104);
and U21015 (N_21015,N_19141,N_19095);
or U21016 (N_21016,N_19500,N_19402);
nand U21017 (N_21017,N_18803,N_18940);
nand U21018 (N_21018,N_18933,N_19787);
or U21019 (N_21019,N_19391,N_19988);
nand U21020 (N_21020,N_18973,N_18969);
nand U21021 (N_21021,N_19415,N_19868);
nand U21022 (N_21022,N_19950,N_19884);
nand U21023 (N_21023,N_19784,N_19458);
or U21024 (N_21024,N_19018,N_19464);
xnor U21025 (N_21025,N_19201,N_19757);
nand U21026 (N_21026,N_19285,N_18900);
or U21027 (N_21027,N_19429,N_19359);
xnor U21028 (N_21028,N_19469,N_18935);
or U21029 (N_21029,N_19171,N_19259);
nand U21030 (N_21030,N_19341,N_19588);
and U21031 (N_21031,N_19808,N_19636);
xnor U21032 (N_21032,N_18959,N_19403);
xor U21033 (N_21033,N_19477,N_18824);
nor U21034 (N_21034,N_19784,N_19413);
xnor U21035 (N_21035,N_18757,N_19885);
xnor U21036 (N_21036,N_19025,N_19145);
or U21037 (N_21037,N_18997,N_19390);
nor U21038 (N_21038,N_19023,N_19820);
nor U21039 (N_21039,N_18914,N_19663);
xor U21040 (N_21040,N_19531,N_19981);
nand U21041 (N_21041,N_19316,N_19689);
nand U21042 (N_21042,N_19475,N_18935);
xnor U21043 (N_21043,N_19934,N_19287);
nand U21044 (N_21044,N_19067,N_19195);
nor U21045 (N_21045,N_19223,N_19180);
or U21046 (N_21046,N_19993,N_19970);
xnor U21047 (N_21047,N_19107,N_19943);
xnor U21048 (N_21048,N_19065,N_19467);
nor U21049 (N_21049,N_19721,N_19786);
nand U21050 (N_21050,N_19384,N_19562);
and U21051 (N_21051,N_19972,N_19966);
nand U21052 (N_21052,N_19124,N_19186);
or U21053 (N_21053,N_19198,N_19344);
or U21054 (N_21054,N_18793,N_19529);
xnor U21055 (N_21055,N_19651,N_19956);
xnor U21056 (N_21056,N_19317,N_19095);
xor U21057 (N_21057,N_19792,N_19134);
and U21058 (N_21058,N_19925,N_18892);
and U21059 (N_21059,N_19850,N_19966);
nor U21060 (N_21060,N_19315,N_19083);
nor U21061 (N_21061,N_18984,N_19838);
and U21062 (N_21062,N_19507,N_19828);
nor U21063 (N_21063,N_19041,N_19620);
nand U21064 (N_21064,N_19409,N_19317);
xnor U21065 (N_21065,N_19373,N_18995);
and U21066 (N_21066,N_19238,N_19200);
or U21067 (N_21067,N_19078,N_19794);
nor U21068 (N_21068,N_18897,N_19998);
or U21069 (N_21069,N_19111,N_19766);
nand U21070 (N_21070,N_19553,N_19024);
xnor U21071 (N_21071,N_19817,N_19857);
or U21072 (N_21072,N_19158,N_19702);
nor U21073 (N_21073,N_19417,N_18806);
nor U21074 (N_21074,N_18996,N_19770);
nor U21075 (N_21075,N_19813,N_19579);
nand U21076 (N_21076,N_19308,N_19718);
and U21077 (N_21077,N_18847,N_18905);
and U21078 (N_21078,N_19705,N_18767);
nor U21079 (N_21079,N_19806,N_19964);
xnor U21080 (N_21080,N_19573,N_18777);
nand U21081 (N_21081,N_19604,N_19402);
nand U21082 (N_21082,N_18964,N_18829);
nor U21083 (N_21083,N_18865,N_19748);
or U21084 (N_21084,N_18834,N_18790);
xor U21085 (N_21085,N_19467,N_19639);
xnor U21086 (N_21086,N_19630,N_18916);
and U21087 (N_21087,N_19632,N_19683);
and U21088 (N_21088,N_19173,N_19136);
or U21089 (N_21089,N_19362,N_19355);
nor U21090 (N_21090,N_19245,N_19192);
or U21091 (N_21091,N_19448,N_19380);
nand U21092 (N_21092,N_19466,N_19384);
nand U21093 (N_21093,N_19612,N_19144);
or U21094 (N_21094,N_19020,N_19438);
nor U21095 (N_21095,N_19038,N_19593);
nand U21096 (N_21096,N_19720,N_19138);
nand U21097 (N_21097,N_19258,N_19011);
and U21098 (N_21098,N_19900,N_19526);
nor U21099 (N_21099,N_19868,N_19134);
xor U21100 (N_21100,N_19011,N_19270);
and U21101 (N_21101,N_18812,N_19694);
and U21102 (N_21102,N_19368,N_19892);
nand U21103 (N_21103,N_18879,N_19175);
nand U21104 (N_21104,N_19717,N_19036);
xor U21105 (N_21105,N_19442,N_19449);
nand U21106 (N_21106,N_19129,N_19781);
xnor U21107 (N_21107,N_19410,N_18905);
and U21108 (N_21108,N_19380,N_19140);
nand U21109 (N_21109,N_19257,N_19955);
nand U21110 (N_21110,N_19380,N_19215);
xnor U21111 (N_21111,N_19352,N_19978);
nand U21112 (N_21112,N_19596,N_19691);
nor U21113 (N_21113,N_18784,N_19525);
nand U21114 (N_21114,N_19472,N_19884);
nor U21115 (N_21115,N_18964,N_19084);
or U21116 (N_21116,N_19595,N_19126);
or U21117 (N_21117,N_18778,N_19439);
nand U21118 (N_21118,N_19426,N_19770);
nand U21119 (N_21119,N_19806,N_19471);
or U21120 (N_21120,N_19643,N_19829);
xnor U21121 (N_21121,N_18818,N_19885);
xnor U21122 (N_21122,N_19744,N_19727);
nand U21123 (N_21123,N_19972,N_19904);
xor U21124 (N_21124,N_19466,N_19529);
nor U21125 (N_21125,N_19452,N_19083);
nor U21126 (N_21126,N_18926,N_19287);
nand U21127 (N_21127,N_19947,N_19550);
nor U21128 (N_21128,N_18770,N_19765);
nor U21129 (N_21129,N_19593,N_19547);
and U21130 (N_21130,N_19295,N_19462);
and U21131 (N_21131,N_19650,N_19138);
nand U21132 (N_21132,N_18919,N_19344);
or U21133 (N_21133,N_19882,N_19445);
nand U21134 (N_21134,N_19670,N_19413);
nor U21135 (N_21135,N_19241,N_19273);
nor U21136 (N_21136,N_19562,N_18785);
or U21137 (N_21137,N_19592,N_19867);
nand U21138 (N_21138,N_19496,N_19546);
nand U21139 (N_21139,N_19488,N_19472);
xor U21140 (N_21140,N_19289,N_19279);
nor U21141 (N_21141,N_19796,N_19360);
nand U21142 (N_21142,N_19171,N_19087);
nand U21143 (N_21143,N_19816,N_19189);
or U21144 (N_21144,N_18875,N_18980);
or U21145 (N_21145,N_19789,N_18797);
or U21146 (N_21146,N_18820,N_19371);
nor U21147 (N_21147,N_19723,N_19789);
xor U21148 (N_21148,N_19710,N_19444);
xnor U21149 (N_21149,N_19826,N_19098);
nor U21150 (N_21150,N_19277,N_19312);
and U21151 (N_21151,N_19843,N_19453);
nand U21152 (N_21152,N_18850,N_19028);
nand U21153 (N_21153,N_19243,N_19619);
nor U21154 (N_21154,N_19465,N_19798);
and U21155 (N_21155,N_19283,N_19626);
nand U21156 (N_21156,N_19824,N_19026);
nand U21157 (N_21157,N_19601,N_19679);
nand U21158 (N_21158,N_18798,N_19163);
and U21159 (N_21159,N_18806,N_19721);
xor U21160 (N_21160,N_19575,N_19357);
nand U21161 (N_21161,N_19598,N_19292);
and U21162 (N_21162,N_19029,N_18882);
nor U21163 (N_21163,N_18755,N_19981);
nand U21164 (N_21164,N_19106,N_18924);
and U21165 (N_21165,N_19244,N_18862);
or U21166 (N_21166,N_19655,N_19538);
or U21167 (N_21167,N_19884,N_18783);
and U21168 (N_21168,N_19658,N_18981);
nor U21169 (N_21169,N_19665,N_19379);
xnor U21170 (N_21170,N_19926,N_19839);
nor U21171 (N_21171,N_19409,N_19959);
nor U21172 (N_21172,N_19672,N_19392);
and U21173 (N_21173,N_19957,N_19420);
nand U21174 (N_21174,N_19484,N_19576);
xnor U21175 (N_21175,N_19120,N_19140);
and U21176 (N_21176,N_19151,N_19299);
and U21177 (N_21177,N_18901,N_19400);
or U21178 (N_21178,N_18944,N_19403);
nor U21179 (N_21179,N_18874,N_18877);
nor U21180 (N_21180,N_18821,N_19227);
nand U21181 (N_21181,N_18921,N_19090);
or U21182 (N_21182,N_19574,N_19717);
or U21183 (N_21183,N_19004,N_19735);
and U21184 (N_21184,N_19266,N_19743);
nor U21185 (N_21185,N_19221,N_19079);
or U21186 (N_21186,N_18904,N_19189);
nand U21187 (N_21187,N_19348,N_19360);
nand U21188 (N_21188,N_19733,N_18847);
xor U21189 (N_21189,N_19041,N_18945);
xnor U21190 (N_21190,N_19409,N_19144);
nand U21191 (N_21191,N_19085,N_19261);
or U21192 (N_21192,N_19992,N_19791);
xor U21193 (N_21193,N_19049,N_19069);
or U21194 (N_21194,N_18834,N_18840);
nand U21195 (N_21195,N_19826,N_19304);
nor U21196 (N_21196,N_19573,N_19508);
or U21197 (N_21197,N_19533,N_18802);
nor U21198 (N_21198,N_19940,N_19905);
nor U21199 (N_21199,N_19467,N_19469);
or U21200 (N_21200,N_18785,N_18870);
and U21201 (N_21201,N_19852,N_18848);
nor U21202 (N_21202,N_19723,N_19944);
xor U21203 (N_21203,N_19891,N_19373);
nor U21204 (N_21204,N_18813,N_19139);
nor U21205 (N_21205,N_18800,N_19184);
nor U21206 (N_21206,N_19603,N_19825);
nand U21207 (N_21207,N_19222,N_19575);
and U21208 (N_21208,N_19978,N_19117);
xor U21209 (N_21209,N_19343,N_19109);
and U21210 (N_21210,N_19266,N_19175);
xor U21211 (N_21211,N_19878,N_18996);
xnor U21212 (N_21212,N_19005,N_19762);
and U21213 (N_21213,N_18780,N_19845);
or U21214 (N_21214,N_19087,N_19737);
nand U21215 (N_21215,N_19492,N_19107);
xor U21216 (N_21216,N_19383,N_19426);
nor U21217 (N_21217,N_19060,N_19408);
nand U21218 (N_21218,N_19438,N_18767);
xor U21219 (N_21219,N_19717,N_19258);
nand U21220 (N_21220,N_19408,N_19281);
nor U21221 (N_21221,N_19801,N_18808);
and U21222 (N_21222,N_19954,N_18995);
and U21223 (N_21223,N_18968,N_19265);
or U21224 (N_21224,N_19472,N_18827);
xor U21225 (N_21225,N_19983,N_19812);
nand U21226 (N_21226,N_19867,N_18771);
nor U21227 (N_21227,N_19981,N_19267);
or U21228 (N_21228,N_19074,N_18873);
nand U21229 (N_21229,N_19577,N_19616);
or U21230 (N_21230,N_19200,N_18908);
nand U21231 (N_21231,N_19325,N_19611);
nand U21232 (N_21232,N_19947,N_19030);
and U21233 (N_21233,N_19573,N_19240);
and U21234 (N_21234,N_19422,N_18806);
nand U21235 (N_21235,N_19332,N_19524);
xor U21236 (N_21236,N_19467,N_19316);
and U21237 (N_21237,N_19510,N_19680);
nor U21238 (N_21238,N_19513,N_19939);
nor U21239 (N_21239,N_19742,N_19443);
nor U21240 (N_21240,N_19373,N_19368);
xor U21241 (N_21241,N_18999,N_19195);
nor U21242 (N_21242,N_19574,N_19169);
and U21243 (N_21243,N_19227,N_19866);
or U21244 (N_21244,N_19864,N_18881);
nand U21245 (N_21245,N_19233,N_19087);
xnor U21246 (N_21246,N_19643,N_19476);
xnor U21247 (N_21247,N_19149,N_18797);
and U21248 (N_21248,N_19003,N_18750);
nor U21249 (N_21249,N_18832,N_18897);
nor U21250 (N_21250,N_20050,N_20999);
xnor U21251 (N_21251,N_20422,N_20771);
and U21252 (N_21252,N_20402,N_20926);
or U21253 (N_21253,N_20161,N_20718);
or U21254 (N_21254,N_20469,N_20737);
xor U21255 (N_21255,N_21229,N_20272);
and U21256 (N_21256,N_20073,N_21001);
and U21257 (N_21257,N_20363,N_21117);
nor U21258 (N_21258,N_20724,N_20957);
or U21259 (N_21259,N_20768,N_20406);
nand U21260 (N_21260,N_20747,N_20896);
or U21261 (N_21261,N_20556,N_20792);
and U21262 (N_21262,N_20893,N_20357);
nand U21263 (N_21263,N_20485,N_21058);
or U21264 (N_21264,N_21177,N_20965);
and U21265 (N_21265,N_20269,N_21221);
and U21266 (N_21266,N_21029,N_21031);
or U21267 (N_21267,N_21243,N_21174);
nand U21268 (N_21268,N_20389,N_20544);
or U21269 (N_21269,N_20317,N_20876);
and U21270 (N_21270,N_20902,N_20000);
xnor U21271 (N_21271,N_20477,N_20150);
nor U21272 (N_21272,N_20114,N_20750);
nand U21273 (N_21273,N_20882,N_20763);
or U21274 (N_21274,N_20894,N_20250);
and U21275 (N_21275,N_20419,N_20142);
nand U21276 (N_21276,N_20734,N_20978);
xor U21277 (N_21277,N_21152,N_20887);
and U21278 (N_21278,N_20171,N_20910);
and U21279 (N_21279,N_20574,N_20232);
and U21280 (N_21280,N_20351,N_20971);
xor U21281 (N_21281,N_20413,N_20968);
and U21282 (N_21282,N_20020,N_20289);
xor U21283 (N_21283,N_20921,N_20502);
or U21284 (N_21284,N_20738,N_20546);
and U21285 (N_21285,N_20381,N_20671);
nor U21286 (N_21286,N_20519,N_20811);
and U21287 (N_21287,N_20658,N_20683);
xor U21288 (N_21288,N_20342,N_20677);
and U21289 (N_21289,N_20157,N_20547);
and U21290 (N_21290,N_20636,N_20437);
nor U21291 (N_21291,N_20529,N_20935);
nand U21292 (N_21292,N_20789,N_20576);
nor U21293 (N_21293,N_21018,N_20487);
nand U21294 (N_21294,N_21138,N_20909);
nor U21295 (N_21295,N_20878,N_20613);
or U21296 (N_21296,N_20224,N_20135);
nand U21297 (N_21297,N_20091,N_20620);
and U21298 (N_21298,N_20949,N_20831);
xnor U21299 (N_21299,N_21139,N_20640);
nand U21300 (N_21300,N_21013,N_20726);
and U21301 (N_21301,N_20065,N_20056);
and U21302 (N_21302,N_20031,N_20879);
or U21303 (N_21303,N_20537,N_20324);
nand U21304 (N_21304,N_21072,N_20967);
xor U21305 (N_21305,N_21151,N_20781);
xnor U21306 (N_21306,N_20542,N_20992);
xor U21307 (N_21307,N_20815,N_20264);
nand U21308 (N_21308,N_21027,N_20594);
nor U21309 (N_21309,N_20390,N_20454);
and U21310 (N_21310,N_20047,N_20665);
nand U21311 (N_21311,N_21154,N_20805);
xor U21312 (N_21312,N_20943,N_20557);
nor U21313 (N_21313,N_20731,N_20818);
and U21314 (N_21314,N_20849,N_20609);
and U21315 (N_21315,N_21225,N_20757);
or U21316 (N_21316,N_20721,N_20581);
nand U21317 (N_21317,N_20470,N_21180);
or U21318 (N_21318,N_20281,N_20712);
nand U21319 (N_21319,N_20039,N_21047);
nand U21320 (N_21320,N_21066,N_20223);
or U21321 (N_21321,N_20693,N_20072);
xnor U21322 (N_21322,N_20941,N_20361);
and U21323 (N_21323,N_20848,N_20146);
or U21324 (N_21324,N_20570,N_21220);
nor U21325 (N_21325,N_20472,N_20797);
and U21326 (N_21326,N_20899,N_21133);
xor U21327 (N_21327,N_20467,N_20139);
or U21328 (N_21328,N_21218,N_20503);
nor U21329 (N_21329,N_20372,N_21040);
xor U21330 (N_21330,N_20687,N_20365);
and U21331 (N_21331,N_20134,N_21006);
nand U21332 (N_21332,N_21135,N_20641);
nand U21333 (N_21333,N_20074,N_20951);
and U21334 (N_21334,N_20932,N_20486);
xor U21335 (N_21335,N_21217,N_20707);
nand U21336 (N_21336,N_20117,N_20204);
or U21337 (N_21337,N_20830,N_21056);
nand U21338 (N_21338,N_20776,N_21216);
nor U21339 (N_21339,N_20456,N_20458);
nand U21340 (N_21340,N_20660,N_21140);
nor U21341 (N_21341,N_21231,N_21237);
or U21342 (N_21342,N_20858,N_21089);
and U21343 (N_21343,N_20220,N_20990);
and U21344 (N_21344,N_20037,N_20447);
xor U21345 (N_21345,N_20698,N_20307);
and U21346 (N_21346,N_21012,N_20144);
nor U21347 (N_21347,N_20685,N_20551);
xor U21348 (N_21348,N_20748,N_21239);
or U21349 (N_21349,N_21205,N_20082);
or U21350 (N_21350,N_20780,N_20730);
and U21351 (N_21351,N_20398,N_20042);
nor U21352 (N_21352,N_21008,N_20309);
or U21353 (N_21353,N_20975,N_20610);
nor U21354 (N_21354,N_20643,N_20137);
or U21355 (N_21355,N_20178,N_20661);
nand U21356 (N_21356,N_21079,N_21141);
nor U21357 (N_21357,N_21175,N_21094);
or U21358 (N_21358,N_20828,N_20233);
and U21359 (N_21359,N_20931,N_20060);
or U21360 (N_21360,N_20121,N_21044);
nor U21361 (N_21361,N_20913,N_20038);
and U21362 (N_21362,N_20517,N_20350);
or U21363 (N_21363,N_20639,N_20782);
nor U21364 (N_21364,N_20918,N_21041);
nand U21365 (N_21365,N_20187,N_21145);
xor U21366 (N_21366,N_21198,N_20235);
or U21367 (N_21367,N_20754,N_20369);
or U21368 (N_21368,N_20206,N_21105);
nand U21369 (N_21369,N_20010,N_21214);
nand U21370 (N_21370,N_21063,N_20428);
nand U21371 (N_21371,N_20339,N_20623);
nand U21372 (N_21372,N_20680,N_20778);
xor U21373 (N_21373,N_20638,N_20521);
and U21374 (N_21374,N_20430,N_21017);
nor U21375 (N_21375,N_20238,N_20790);
and U21376 (N_21376,N_20938,N_20153);
xor U21377 (N_21377,N_20802,N_20567);
nor U21378 (N_21378,N_20656,N_20328);
and U21379 (N_21379,N_21093,N_20262);
xnor U21380 (N_21380,N_20572,N_20159);
nand U21381 (N_21381,N_20291,N_20268);
xor U21382 (N_21382,N_20714,N_20504);
and U21383 (N_21383,N_20032,N_20427);
or U21384 (N_21384,N_20842,N_21202);
or U21385 (N_21385,N_20579,N_21206);
or U21386 (N_21386,N_20490,N_20118);
and U21387 (N_21387,N_20961,N_21087);
nand U21388 (N_21388,N_20482,N_20588);
xor U21389 (N_21389,N_20801,N_20761);
or U21390 (N_21390,N_20431,N_20966);
nor U21391 (N_21391,N_20319,N_20024);
nand U21392 (N_21392,N_20426,N_20884);
or U21393 (N_21393,N_20548,N_20699);
and U21394 (N_21394,N_20285,N_20225);
nand U21395 (N_21395,N_20922,N_21098);
and U21396 (N_21396,N_20435,N_20634);
nand U21397 (N_21397,N_20892,N_20322);
and U21398 (N_21398,N_20555,N_20930);
or U21399 (N_21399,N_20933,N_20956);
and U21400 (N_21400,N_20676,N_21197);
and U21401 (N_21401,N_21023,N_20253);
nor U21402 (N_21402,N_20559,N_20786);
nor U21403 (N_21403,N_21025,N_20071);
and U21404 (N_21404,N_21156,N_20360);
xor U21405 (N_21405,N_21115,N_20051);
or U21406 (N_21406,N_20822,N_20258);
nor U21407 (N_21407,N_20785,N_20596);
nand U21408 (N_21408,N_20181,N_20464);
or U21409 (N_21409,N_20382,N_20147);
or U21410 (N_21410,N_20334,N_20649);
xor U21411 (N_21411,N_20563,N_20260);
nand U21412 (N_21412,N_20217,N_20314);
nor U21413 (N_21413,N_21035,N_20216);
nor U21414 (N_21414,N_20948,N_20564);
nor U21415 (N_21415,N_20702,N_20173);
xor U21416 (N_21416,N_20531,N_21132);
xnor U21417 (N_21417,N_20982,N_20799);
and U21418 (N_21418,N_20923,N_20720);
nor U21419 (N_21419,N_20937,N_20580);
nor U21420 (N_21420,N_20380,N_20344);
nor U21421 (N_21421,N_20222,N_21245);
nand U21422 (N_21422,N_21061,N_20424);
xor U21423 (N_21423,N_20346,N_20195);
nor U21424 (N_21424,N_20190,N_20652);
or U21425 (N_21425,N_20608,N_21074);
nand U21426 (N_21426,N_20078,N_20199);
nor U21427 (N_21427,N_20908,N_21034);
nor U21428 (N_21428,N_20343,N_20688);
or U21429 (N_21429,N_21130,N_20906);
or U21430 (N_21430,N_20098,N_20626);
nor U21431 (N_21431,N_20851,N_20697);
nand U21432 (N_21432,N_21182,N_20311);
and U21433 (N_21433,N_20023,N_20664);
and U21434 (N_21434,N_21129,N_21149);
nor U21435 (N_21435,N_20535,N_20184);
xor U21436 (N_21436,N_21199,N_20777);
nand U21437 (N_21437,N_20501,N_20434);
xor U21438 (N_21438,N_21172,N_21136);
and U21439 (N_21439,N_21230,N_20293);
xor U21440 (N_21440,N_21187,N_20871);
nand U21441 (N_21441,N_20586,N_20500);
xnor U21442 (N_21442,N_20227,N_20617);
or U21443 (N_21443,N_20874,N_20340);
or U21444 (N_21444,N_20616,N_20306);
nand U21445 (N_21445,N_20527,N_21084);
and U21446 (N_21446,N_20138,N_20973);
or U21447 (N_21447,N_20854,N_20226);
nor U21448 (N_21448,N_20300,N_21071);
or U21449 (N_21449,N_20415,N_20296);
nor U21450 (N_21450,N_20847,N_21178);
nand U21451 (N_21451,N_20280,N_21113);
and U21452 (N_21452,N_20077,N_21015);
xnor U21453 (N_21453,N_20104,N_21030);
xnor U21454 (N_21454,N_20409,N_20468);
nor U21455 (N_21455,N_20585,N_20455);
nor U21456 (N_21456,N_20614,N_20888);
xor U21457 (N_21457,N_20094,N_20928);
xnor U21458 (N_21458,N_21110,N_20651);
and U21459 (N_21459,N_20857,N_21192);
nor U21460 (N_21460,N_20189,N_20516);
nand U21461 (N_21461,N_20662,N_21165);
xor U21462 (N_21462,N_20920,N_20653);
xor U21463 (N_21463,N_20566,N_20067);
or U21464 (N_21464,N_20393,N_20686);
xor U21465 (N_21465,N_20550,N_21005);
or U21466 (N_21466,N_20259,N_21224);
nor U21467 (N_21467,N_21143,N_20678);
or U21468 (N_21468,N_21236,N_20043);
nor U21469 (N_21469,N_20715,N_21091);
or U21470 (N_21470,N_20940,N_20116);
nor U21471 (N_21471,N_21007,N_20758);
xor U21472 (N_21472,N_20997,N_20299);
xnor U21473 (N_21473,N_21150,N_20331);
nor U21474 (N_21474,N_20944,N_20185);
and U21475 (N_21475,N_21200,N_20095);
nor U21476 (N_21476,N_20635,N_20998);
and U21477 (N_21477,N_21026,N_20110);
nand U21478 (N_21478,N_20645,N_21060);
nand U21479 (N_21479,N_20945,N_20080);
or U21480 (N_21480,N_20420,N_20592);
and U21481 (N_21481,N_20606,N_20993);
nor U21482 (N_21482,N_20582,N_21184);
or U21483 (N_21483,N_20995,N_21123);
nor U21484 (N_21484,N_20001,N_20618);
or U21485 (N_21485,N_20341,N_21168);
nand U21486 (N_21486,N_20076,N_21042);
and U21487 (N_21487,N_21137,N_20081);
xor U21488 (N_21488,N_21109,N_20362);
nand U21489 (N_21489,N_20172,N_20079);
or U21490 (N_21490,N_20006,N_20979);
or U21491 (N_21491,N_20727,N_20283);
xor U21492 (N_21492,N_21191,N_20611);
or U21493 (N_21493,N_21088,N_21002);
or U21494 (N_21494,N_20191,N_21037);
nor U21495 (N_21495,N_20182,N_21083);
and U21496 (N_21496,N_20347,N_21104);
or U21497 (N_21497,N_20637,N_20353);
and U21498 (N_21498,N_20866,N_20773);
or U21499 (N_21499,N_20087,N_20549);
xor U21500 (N_21500,N_21022,N_20495);
and U21501 (N_21501,N_20621,N_21227);
nor U21502 (N_21502,N_20140,N_20729);
and U21503 (N_21503,N_20439,N_20751);
nand U21504 (N_21504,N_20700,N_20392);
xnor U21505 (N_21505,N_20929,N_20725);
and U21506 (N_21506,N_20479,N_20925);
xnor U21507 (N_21507,N_20105,N_20348);
nand U21508 (N_21508,N_21166,N_20807);
nor U21509 (N_21509,N_20880,N_20524);
and U21510 (N_21510,N_20543,N_20463);
nand U21511 (N_21511,N_20946,N_20732);
or U21512 (N_21512,N_20248,N_20112);
and U21513 (N_21513,N_20744,N_21046);
and U21514 (N_21514,N_20119,N_20212);
or U21515 (N_21515,N_20532,N_21102);
xnor U21516 (N_21516,N_20765,N_21121);
or U21517 (N_21517,N_20452,N_20667);
and U21518 (N_21518,N_20320,N_20958);
or U21519 (N_21519,N_20863,N_20852);
nand U21520 (N_21520,N_20193,N_20101);
and U21521 (N_21521,N_20775,N_20959);
xnor U21522 (N_21522,N_20453,N_20826);
and U21523 (N_21523,N_21081,N_21064);
xnor U21524 (N_21524,N_20666,N_20924);
or U21525 (N_21525,N_20845,N_21226);
and U21526 (N_21526,N_20728,N_20048);
and U21527 (N_21527,N_21235,N_20229);
nor U21528 (N_21528,N_20861,N_20249);
xnor U21529 (N_21529,N_20009,N_20230);
or U21530 (N_21530,N_20312,N_20093);
nor U21531 (N_21531,N_20890,N_20411);
nand U21532 (N_21532,N_21055,N_20399);
or U21533 (N_21533,N_20113,N_20241);
nor U21534 (N_21534,N_20027,N_20040);
nor U21535 (N_21535,N_20021,N_20286);
nor U21536 (N_21536,N_20901,N_21167);
nor U21537 (N_21537,N_20525,N_21107);
nand U21538 (N_21538,N_20266,N_20461);
nor U21539 (N_21539,N_20867,N_20236);
or U21540 (N_21540,N_21067,N_21096);
nand U21541 (N_21541,N_20917,N_20602);
nand U21542 (N_21542,N_20630,N_21033);
nand U21543 (N_21543,N_20597,N_20141);
or U21544 (N_21544,N_21114,N_20962);
nor U21545 (N_21545,N_21201,N_20376);
nor U21546 (N_21546,N_20298,N_20425);
and U21547 (N_21547,N_21085,N_20203);
and U21548 (N_21548,N_20210,N_20265);
nand U21549 (N_21549,N_21103,N_20629);
xnor U21550 (N_21550,N_20335,N_21157);
or U21551 (N_21551,N_20476,N_20569);
nand U21552 (N_21552,N_20315,N_20005);
and U21553 (N_21553,N_20459,N_20267);
xor U21554 (N_21554,N_21119,N_20766);
and U21555 (N_21555,N_20862,N_20974);
or U21556 (N_21556,N_20939,N_20841);
and U21557 (N_21557,N_20796,N_20070);
or U21558 (N_21558,N_20374,N_20791);
nor U21559 (N_21559,N_20183,N_21000);
nor U21560 (N_21560,N_20905,N_20457);
nor U21561 (N_21561,N_20814,N_20247);
nor U21562 (N_21562,N_21124,N_21050);
nor U21563 (N_21563,N_20528,N_20762);
xnor U21564 (N_21564,N_20970,N_20568);
and U21565 (N_21565,N_20631,N_21173);
nor U21566 (N_21566,N_20274,N_20231);
nor U21567 (N_21567,N_20397,N_20752);
or U21568 (N_21568,N_21241,N_21128);
and U21569 (N_21569,N_20869,N_21122);
nor U21570 (N_21570,N_20745,N_21024);
nand U21571 (N_21571,N_20221,N_20994);
nor U21572 (N_21572,N_20451,N_20131);
xor U21573 (N_21573,N_20615,N_20240);
nand U21574 (N_21574,N_20130,N_21045);
xnor U21575 (N_21575,N_20478,N_20349);
xor U21576 (N_21576,N_20211,N_20462);
and U21577 (N_21577,N_20981,N_20207);
nor U21578 (N_21578,N_20154,N_20513);
nor U21579 (N_21579,N_20214,N_20875);
or U21580 (N_21580,N_20522,N_21126);
and U21581 (N_21581,N_21032,N_20625);
or U21582 (N_21582,N_20446,N_20064);
and U21583 (N_21583,N_20192,N_20642);
and U21584 (N_21584,N_20607,N_20689);
xor U21585 (N_21585,N_20488,N_20804);
and U21586 (N_21586,N_20175,N_20739);
and U21587 (N_21587,N_20491,N_20800);
and U21588 (N_21588,N_20986,N_20261);
xnor U21589 (N_21589,N_20953,N_20332);
xnor U21590 (N_21590,N_20165,N_20254);
nor U21591 (N_21591,N_20701,N_20716);
or U21592 (N_21592,N_21171,N_20126);
or U21593 (N_21593,N_21059,N_21207);
or U21594 (N_21594,N_20395,N_20989);
or U21595 (N_21595,N_20659,N_20252);
or U21596 (N_21596,N_20045,N_20520);
or U21597 (N_21597,N_21194,N_20086);
and U21598 (N_21598,N_20885,N_21213);
and U21599 (N_21599,N_20497,N_20041);
nand U21600 (N_21600,N_20684,N_20275);
xnor U21601 (N_21601,N_20417,N_20108);
nand U21602 (N_21602,N_20976,N_21010);
xnor U21603 (N_21603,N_20494,N_20035);
and U21604 (N_21604,N_20595,N_20410);
nand U21605 (N_21605,N_20764,N_20090);
nand U21606 (N_21606,N_21080,N_20234);
nand U21607 (N_21607,N_21147,N_20152);
xnor U21608 (N_21608,N_20736,N_20449);
and U21609 (N_21609,N_21228,N_20011);
nand U21610 (N_21610,N_20242,N_20205);
nor U21611 (N_21611,N_20554,N_20375);
xor U21612 (N_21612,N_20273,N_21065);
nor U21613 (N_21613,N_20075,N_21004);
and U21614 (N_21614,N_20418,N_21208);
or U21615 (N_21615,N_20471,N_21232);
nand U21616 (N_21616,N_20442,N_20534);
and U21617 (N_21617,N_20168,N_21222);
and U21618 (N_21618,N_20012,N_20584);
or U21619 (N_21619,N_20429,N_20954);
and U21620 (N_21620,N_21131,N_20237);
nand U21621 (N_21621,N_21125,N_20466);
xor U21622 (N_21622,N_20870,N_20578);
or U21623 (N_21623,N_21164,N_21011);
and U21624 (N_21624,N_20336,N_20166);
or U21625 (N_21625,N_20278,N_20558);
and U21626 (N_21626,N_20806,N_21193);
xor U21627 (N_21627,N_20359,N_20681);
or U21628 (N_21628,N_20433,N_20808);
or U21629 (N_21629,N_20167,N_20004);
nand U21630 (N_21630,N_20379,N_20279);
nand U21631 (N_21631,N_21210,N_20624);
or U21632 (N_21632,N_20255,N_20028);
or U21633 (N_21633,N_20988,N_20018);
nor U21634 (N_21634,N_20912,N_20565);
nor U21635 (N_21635,N_20384,N_20895);
xor U21636 (N_21636,N_20628,N_21153);
nand U21637 (N_21637,N_21248,N_20352);
nand U21638 (N_21638,N_20391,N_21116);
nand U21639 (N_21639,N_21036,N_20632);
xor U21640 (N_21640,N_20577,N_20277);
xnor U21641 (N_21641,N_20016,N_20834);
or U21642 (N_21642,N_20955,N_21118);
xnor U21643 (N_21643,N_20900,N_20294);
and U21644 (N_21644,N_20052,N_20288);
xor U21645 (N_21645,N_20914,N_21209);
nand U21646 (N_21646,N_20837,N_20002);
nand U21647 (N_21647,N_20819,N_20304);
and U21648 (N_21648,N_20396,N_20904);
or U21649 (N_21649,N_20475,N_20096);
xnor U21650 (N_21650,N_20903,N_21097);
or U21651 (N_21651,N_20784,N_20019);
and U21652 (N_21652,N_20263,N_20129);
nor U21653 (N_21653,N_20526,N_20889);
or U21654 (N_21654,N_21057,N_20936);
nand U21655 (N_21655,N_20062,N_20877);
nor U21656 (N_21656,N_20136,N_20333);
nand U21657 (N_21657,N_21108,N_20151);
nand U21658 (N_21658,N_21204,N_20036);
xnor U21659 (N_21659,N_21038,N_21095);
xor U21660 (N_21660,N_20423,N_20492);
or U21661 (N_21661,N_20239,N_20977);
nand U21662 (N_21662,N_20984,N_20017);
nand U21663 (N_21663,N_21051,N_21048);
or U21664 (N_21664,N_21075,N_20753);
xor U21665 (N_21665,N_20364,N_20741);
nand U21666 (N_21666,N_20155,N_20102);
nor U21667 (N_21667,N_20600,N_20703);
nor U21668 (N_21668,N_20985,N_21043);
nor U21669 (N_21669,N_20633,N_20313);
nor U21670 (N_21670,N_20650,N_20509);
or U21671 (N_21671,N_20125,N_20599);
xor U21672 (N_21672,N_20836,N_20327);
and U21673 (N_21673,N_21092,N_20111);
nand U21674 (N_21674,N_20326,N_20886);
nor U21675 (N_21675,N_20055,N_20746);
xnor U21676 (N_21676,N_20496,N_20589);
and U21677 (N_21677,N_20044,N_20068);
and U21678 (N_21678,N_20827,N_20169);
nand U21679 (N_21679,N_20832,N_20162);
or U21680 (N_21680,N_20186,N_20106);
and U21681 (N_21681,N_20561,N_20257);
and U21682 (N_21682,N_21238,N_20619);
nor U21683 (N_21683,N_20856,N_21019);
nand U21684 (N_21684,N_20323,N_20194);
nand U21685 (N_21685,N_20270,N_20646);
xnor U21686 (N_21686,N_21016,N_20530);
nor U21687 (N_21687,N_21069,N_20541);
xor U21688 (N_21688,N_20156,N_20694);
nor U21689 (N_21689,N_20934,N_20759);
xor U21690 (N_21690,N_20829,N_20123);
nor U21691 (N_21691,N_20755,N_20163);
or U21692 (N_21692,N_20403,N_20545);
and U21693 (N_21693,N_20601,N_20246);
or U21694 (N_21694,N_20622,N_20860);
and U21695 (N_21695,N_20907,N_20122);
xnor U21696 (N_21696,N_20083,N_20838);
xor U21697 (N_21697,N_21195,N_20059);
nor U21698 (N_21698,N_20404,N_20089);
or U21699 (N_21699,N_21106,N_20927);
and U21700 (N_21700,N_20711,N_20085);
xnor U21701 (N_21701,N_20627,N_20612);
or U21702 (N_21702,N_20813,N_20603);
nor U21703 (N_21703,N_21134,N_20505);
or U21704 (N_21704,N_20911,N_20109);
nand U21705 (N_21705,N_20243,N_20881);
nand U21706 (N_21706,N_20305,N_20180);
xnor U21707 (N_21707,N_21052,N_20049);
or U21708 (N_21708,N_21158,N_20450);
and U21709 (N_21709,N_20713,N_21176);
and U21710 (N_21710,N_20321,N_20355);
and U21711 (N_21711,N_21247,N_20803);
nand U21712 (N_21712,N_20164,N_20710);
or U21713 (N_21713,N_21127,N_20473);
and U21714 (N_21714,N_20919,N_20378);
xor U21715 (N_21715,N_20795,N_20061);
or U21716 (N_21716,N_20124,N_20760);
nor U21717 (N_21717,N_20007,N_20480);
nor U21718 (N_21718,N_20682,N_20891);
and U21719 (N_21719,N_21021,N_20969);
and U21720 (N_21720,N_20740,N_20810);
or U21721 (N_21721,N_20358,N_20432);
xnor U21722 (N_21722,N_20174,N_20510);
or U21723 (N_21723,N_21185,N_20950);
or U21724 (N_21724,N_20952,N_20735);
xnor U21725 (N_21725,N_21028,N_21146);
and U21726 (N_21726,N_20663,N_20850);
and U21727 (N_21727,N_20297,N_20996);
nor U21728 (N_21728,N_20014,N_20514);
nor U21729 (N_21729,N_20722,N_21183);
nand U21730 (N_21730,N_20026,N_20244);
xnor U21731 (N_21731,N_20499,N_20282);
nor U21732 (N_21732,N_20583,N_20844);
xnor U21733 (N_21733,N_20460,N_20394);
nor U21734 (N_21734,N_20657,N_20506);
or U21735 (N_21735,N_20654,N_21120);
and U21736 (N_21736,N_20388,N_20817);
nand U21737 (N_21737,N_21162,N_20148);
xnor U21738 (N_21738,N_20201,N_21219);
or U21739 (N_21739,N_20987,N_20655);
xor U21740 (N_21740,N_20809,N_21234);
nand U21741 (N_21741,N_20103,N_20198);
and U21742 (N_21742,N_20295,N_20587);
xnor U21743 (N_21743,N_20916,N_20318);
xor U21744 (N_21744,N_20915,N_21070);
nand U21745 (N_21745,N_20675,N_20046);
or U21746 (N_21746,N_21144,N_20251);
or U21747 (N_21747,N_21039,N_21163);
nor U21748 (N_21748,N_20839,N_20679);
nand U21749 (N_21749,N_20245,N_21196);
nand U21750 (N_21750,N_20143,N_20213);
nand U21751 (N_21751,N_20196,N_20772);
xnor U21752 (N_21752,N_20414,N_20825);
and U21753 (N_21753,N_20387,N_20128);
nor U21754 (N_21754,N_20864,N_20115);
or U21755 (N_21755,N_20408,N_20824);
or U21756 (N_21756,N_20030,N_20107);
and U21757 (N_21757,N_20717,N_21240);
xnor U21758 (N_21758,N_20821,N_20648);
nor U21759 (N_21759,N_20840,N_21161);
and U21760 (N_21760,N_20448,N_20539);
and U21761 (N_21761,N_20942,N_20573);
or U21762 (N_21762,N_20668,N_20533);
xor U21763 (N_21763,N_20742,N_21014);
nor U21764 (N_21764,N_20575,N_20100);
xor U21765 (N_21765,N_20644,N_21233);
and U21766 (N_21766,N_20022,N_21160);
nor U21767 (N_21767,N_20385,N_20843);
xor U21768 (N_21768,N_20063,N_21062);
nand U21769 (N_21769,N_20383,N_20444);
nand U21770 (N_21770,N_20883,N_20672);
or U21771 (N_21771,N_21203,N_20176);
and U21772 (N_21772,N_20188,N_20092);
or U21773 (N_21773,N_20438,N_20033);
or U21774 (N_21774,N_20366,N_20058);
or U21775 (N_21775,N_20498,N_20704);
xor U21776 (N_21776,N_20647,N_20256);
and U21777 (N_21777,N_20345,N_20310);
nor U21778 (N_21778,N_20695,N_20066);
and U21779 (N_21779,N_21076,N_21181);
nand U21780 (N_21780,N_20846,N_20540);
nor U21781 (N_21781,N_21003,N_21068);
and U21782 (N_21782,N_20330,N_20793);
nand U21783 (N_21783,N_20593,N_20590);
or U21784 (N_21784,N_20960,N_20538);
or U21785 (N_21785,N_20407,N_20003);
and U21786 (N_21786,N_20972,N_20301);
nor U21787 (N_21787,N_20898,N_21009);
nor U21788 (N_21788,N_20794,N_21190);
nor U21789 (N_21789,N_21223,N_20571);
and U21790 (N_21790,N_20099,N_20177);
nor U21791 (N_21791,N_21054,N_21169);
nand U21792 (N_21792,N_21179,N_20057);
nand U21793 (N_21793,N_20370,N_20440);
and U21794 (N_21794,N_20287,N_20228);
or U21795 (N_21795,N_20474,N_21215);
nand U21796 (N_21796,N_20964,N_21086);
and U21797 (N_21797,N_20855,N_20054);
or U21798 (N_21798,N_20405,N_20692);
nand U21799 (N_21799,N_20511,N_20149);
or U21800 (N_21800,N_20508,N_20709);
and U21801 (N_21801,N_20674,N_21211);
or U21802 (N_21802,N_20316,N_20013);
xor U21803 (N_21803,N_20756,N_20401);
nand U21804 (N_21804,N_21186,N_20133);
xor U21805 (N_21805,N_20980,N_20512);
nor U21806 (N_21806,N_21049,N_20897);
or U21807 (N_21807,N_20088,N_20605);
or U21808 (N_21808,N_20276,N_20025);
xnor U21809 (N_21809,N_21170,N_21078);
and U21810 (N_21810,N_20158,N_20356);
or U21811 (N_21811,N_20489,N_20767);
or U21812 (N_21812,N_20493,N_20271);
or U21813 (N_21813,N_20481,N_20197);
nand U21814 (N_21814,N_20354,N_20484);
xor U21815 (N_21815,N_20373,N_20127);
nand U21816 (N_21816,N_20719,N_20284);
nor U21817 (N_21817,N_20367,N_20873);
and U21818 (N_21818,N_20769,N_20669);
or U21819 (N_21819,N_20436,N_20338);
nor U21820 (N_21820,N_20591,N_20868);
and U21821 (N_21821,N_20812,N_21082);
and U21822 (N_21822,N_21112,N_20069);
and U21823 (N_21823,N_20743,N_21142);
xnor U21824 (N_21824,N_20145,N_21246);
or U21825 (N_21825,N_20816,N_20084);
nor U21826 (N_21826,N_20303,N_20308);
and U21827 (N_21827,N_20292,N_20823);
or U21828 (N_21828,N_20218,N_20859);
nor U21829 (N_21829,N_20337,N_20788);
nor U21830 (N_21830,N_21099,N_20445);
nand U21831 (N_21831,N_20290,N_20733);
nor U21832 (N_21832,N_20723,N_20015);
and U21833 (N_21833,N_20783,N_21242);
xor U21834 (N_21834,N_20691,N_20787);
and U21835 (N_21835,N_20132,N_20518);
or U21836 (N_21836,N_20673,N_21073);
nand U21837 (N_21837,N_20421,N_21100);
nor U21838 (N_21838,N_20400,N_20779);
xnor U21839 (N_21839,N_20325,N_21090);
or U21840 (N_21840,N_20416,N_21053);
nor U21841 (N_21841,N_20329,N_20209);
nand U21842 (N_21842,N_20386,N_20412);
or U21843 (N_21843,N_21148,N_20552);
nand U21844 (N_21844,N_21249,N_21188);
xor U21845 (N_21845,N_20872,N_20368);
xnor U21846 (N_21846,N_20553,N_20983);
nand U21847 (N_21847,N_20200,N_21101);
nand U21848 (N_21848,N_20705,N_20604);
nand U21849 (N_21849,N_20523,N_20696);
or U21850 (N_21850,N_20706,N_20598);
nor U21851 (N_21851,N_20170,N_20536);
nand U21852 (N_21852,N_20215,N_20219);
xnor U21853 (N_21853,N_20820,N_20202);
nand U21854 (N_21854,N_20835,N_20441);
nor U21855 (N_21855,N_21159,N_20947);
nand U21856 (N_21856,N_20515,N_20774);
and U21857 (N_21857,N_20853,N_20008);
nand U21858 (N_21858,N_20833,N_20562);
nand U21859 (N_21859,N_20034,N_21189);
or U21860 (N_21860,N_20963,N_21212);
or U21861 (N_21861,N_21020,N_20798);
nand U21862 (N_21862,N_20029,N_20208);
nor U21863 (N_21863,N_20670,N_20443);
xor U21864 (N_21864,N_20302,N_20560);
and U21865 (N_21865,N_20749,N_21077);
or U21866 (N_21866,N_20097,N_20179);
nand U21867 (N_21867,N_21155,N_20053);
nor U21868 (N_21868,N_20483,N_20465);
xnor U21869 (N_21869,N_20160,N_20371);
xor U21870 (N_21870,N_21111,N_21244);
xor U21871 (N_21871,N_20708,N_20865);
and U21872 (N_21872,N_20770,N_20377);
and U21873 (N_21873,N_20120,N_20690);
nand U21874 (N_21874,N_20507,N_20991);
nand U21875 (N_21875,N_21207,N_20812);
xnor U21876 (N_21876,N_20303,N_20668);
and U21877 (N_21877,N_20232,N_20691);
or U21878 (N_21878,N_20056,N_20216);
xnor U21879 (N_21879,N_20393,N_20188);
xor U21880 (N_21880,N_20293,N_20991);
nor U21881 (N_21881,N_20275,N_20534);
xnor U21882 (N_21882,N_20414,N_20419);
and U21883 (N_21883,N_20769,N_20695);
nor U21884 (N_21884,N_20922,N_21202);
or U21885 (N_21885,N_20600,N_20956);
nor U21886 (N_21886,N_20006,N_20151);
or U21887 (N_21887,N_20416,N_20201);
or U21888 (N_21888,N_21106,N_21200);
xnor U21889 (N_21889,N_20648,N_20333);
nor U21890 (N_21890,N_20169,N_20148);
or U21891 (N_21891,N_21101,N_21209);
xor U21892 (N_21892,N_20418,N_21059);
or U21893 (N_21893,N_20114,N_20009);
and U21894 (N_21894,N_20220,N_21031);
xor U21895 (N_21895,N_20118,N_20730);
and U21896 (N_21896,N_20003,N_20355);
nand U21897 (N_21897,N_20752,N_20627);
and U21898 (N_21898,N_20195,N_20915);
and U21899 (N_21899,N_21082,N_20767);
nor U21900 (N_21900,N_20124,N_20140);
nor U21901 (N_21901,N_20854,N_20641);
nor U21902 (N_21902,N_20224,N_20889);
nor U21903 (N_21903,N_20347,N_20733);
nor U21904 (N_21904,N_20196,N_20859);
and U21905 (N_21905,N_20662,N_20756);
xnor U21906 (N_21906,N_20294,N_21096);
and U21907 (N_21907,N_20029,N_20307);
nand U21908 (N_21908,N_21239,N_21075);
and U21909 (N_21909,N_20770,N_20431);
nand U21910 (N_21910,N_20070,N_20221);
or U21911 (N_21911,N_20910,N_20794);
xnor U21912 (N_21912,N_20515,N_20174);
or U21913 (N_21913,N_20922,N_20056);
nor U21914 (N_21914,N_21108,N_20382);
xor U21915 (N_21915,N_20023,N_21140);
xor U21916 (N_21916,N_20181,N_21066);
nor U21917 (N_21917,N_20970,N_20149);
xnor U21918 (N_21918,N_21029,N_20224);
and U21919 (N_21919,N_20302,N_20296);
and U21920 (N_21920,N_21022,N_20913);
xnor U21921 (N_21921,N_20266,N_21046);
xnor U21922 (N_21922,N_20567,N_20255);
nand U21923 (N_21923,N_20993,N_21061);
xor U21924 (N_21924,N_20338,N_20576);
and U21925 (N_21925,N_21020,N_20275);
nor U21926 (N_21926,N_20084,N_20516);
or U21927 (N_21927,N_20439,N_21079);
and U21928 (N_21928,N_20560,N_20286);
nor U21929 (N_21929,N_20914,N_20347);
xor U21930 (N_21930,N_21208,N_20778);
and U21931 (N_21931,N_20616,N_20727);
and U21932 (N_21932,N_21033,N_20120);
nand U21933 (N_21933,N_21125,N_20420);
nand U21934 (N_21934,N_20547,N_20569);
nand U21935 (N_21935,N_20049,N_21213);
and U21936 (N_21936,N_21218,N_21190);
and U21937 (N_21937,N_20567,N_20512);
and U21938 (N_21938,N_21121,N_20301);
xor U21939 (N_21939,N_21011,N_21168);
xor U21940 (N_21940,N_20343,N_20065);
xor U21941 (N_21941,N_20026,N_21141);
nor U21942 (N_21942,N_20865,N_20016);
and U21943 (N_21943,N_21224,N_20641);
or U21944 (N_21944,N_20466,N_20865);
and U21945 (N_21945,N_20911,N_20893);
xnor U21946 (N_21946,N_20501,N_20930);
and U21947 (N_21947,N_20696,N_21090);
or U21948 (N_21948,N_20002,N_20921);
nor U21949 (N_21949,N_20842,N_20316);
nor U21950 (N_21950,N_21053,N_20702);
xor U21951 (N_21951,N_20434,N_20648);
xor U21952 (N_21952,N_20122,N_20581);
or U21953 (N_21953,N_20287,N_21122);
nor U21954 (N_21954,N_20823,N_20649);
nor U21955 (N_21955,N_21156,N_20462);
or U21956 (N_21956,N_20084,N_20069);
nand U21957 (N_21957,N_20479,N_20662);
and U21958 (N_21958,N_20596,N_20750);
nor U21959 (N_21959,N_20423,N_21247);
or U21960 (N_21960,N_21116,N_20986);
nand U21961 (N_21961,N_21087,N_20220);
nor U21962 (N_21962,N_20332,N_20458);
nor U21963 (N_21963,N_20087,N_20917);
or U21964 (N_21964,N_20550,N_20993);
nand U21965 (N_21965,N_20903,N_20626);
xor U21966 (N_21966,N_20717,N_20067);
or U21967 (N_21967,N_20974,N_20391);
nor U21968 (N_21968,N_20215,N_21000);
or U21969 (N_21969,N_20950,N_20863);
or U21970 (N_21970,N_20149,N_20110);
or U21971 (N_21971,N_21133,N_21248);
or U21972 (N_21972,N_20758,N_20265);
and U21973 (N_21973,N_21044,N_20892);
nand U21974 (N_21974,N_20204,N_20119);
and U21975 (N_21975,N_21161,N_21165);
and U21976 (N_21976,N_20167,N_20959);
or U21977 (N_21977,N_20721,N_20080);
or U21978 (N_21978,N_21072,N_20712);
nor U21979 (N_21979,N_20114,N_20261);
xnor U21980 (N_21980,N_20655,N_20196);
nor U21981 (N_21981,N_21043,N_21015);
nand U21982 (N_21982,N_21242,N_20375);
and U21983 (N_21983,N_21128,N_21099);
nand U21984 (N_21984,N_20749,N_20187);
xnor U21985 (N_21985,N_20419,N_20070);
nor U21986 (N_21986,N_21191,N_20126);
or U21987 (N_21987,N_20779,N_21152);
nor U21988 (N_21988,N_20507,N_20688);
or U21989 (N_21989,N_21063,N_20122);
nor U21990 (N_21990,N_21116,N_20174);
nor U21991 (N_21991,N_21170,N_20415);
or U21992 (N_21992,N_20110,N_20257);
xnor U21993 (N_21993,N_20907,N_20321);
xnor U21994 (N_21994,N_20999,N_20038);
nand U21995 (N_21995,N_20088,N_21072);
and U21996 (N_21996,N_20488,N_20463);
xnor U21997 (N_21997,N_20016,N_20019);
xnor U21998 (N_21998,N_20182,N_20215);
nand U21999 (N_21999,N_20751,N_20199);
nor U22000 (N_22000,N_20556,N_20605);
and U22001 (N_22001,N_20730,N_20368);
xor U22002 (N_22002,N_20452,N_20713);
or U22003 (N_22003,N_20133,N_20646);
xor U22004 (N_22004,N_21102,N_20426);
or U22005 (N_22005,N_20113,N_20880);
or U22006 (N_22006,N_20838,N_21016);
or U22007 (N_22007,N_20042,N_20946);
nor U22008 (N_22008,N_20091,N_20393);
and U22009 (N_22009,N_20747,N_20730);
and U22010 (N_22010,N_20218,N_20578);
or U22011 (N_22011,N_20146,N_20065);
xnor U22012 (N_22012,N_20244,N_20069);
and U22013 (N_22013,N_20969,N_20617);
xnor U22014 (N_22014,N_20415,N_21129);
or U22015 (N_22015,N_20586,N_20041);
nor U22016 (N_22016,N_20270,N_20493);
nor U22017 (N_22017,N_20430,N_20136);
nor U22018 (N_22018,N_21105,N_20527);
or U22019 (N_22019,N_20898,N_21015);
nor U22020 (N_22020,N_20143,N_20543);
xor U22021 (N_22021,N_20989,N_20584);
nand U22022 (N_22022,N_21054,N_20247);
xnor U22023 (N_22023,N_20983,N_20905);
or U22024 (N_22024,N_20229,N_20655);
nand U22025 (N_22025,N_20246,N_21100);
or U22026 (N_22026,N_20592,N_21152);
and U22027 (N_22027,N_20495,N_20221);
and U22028 (N_22028,N_20073,N_20107);
nand U22029 (N_22029,N_21144,N_20052);
nand U22030 (N_22030,N_20292,N_20137);
and U22031 (N_22031,N_20346,N_21150);
or U22032 (N_22032,N_20465,N_20807);
xor U22033 (N_22033,N_20049,N_20398);
and U22034 (N_22034,N_20536,N_20728);
or U22035 (N_22035,N_21204,N_20467);
xnor U22036 (N_22036,N_20915,N_20163);
nand U22037 (N_22037,N_20928,N_20204);
nand U22038 (N_22038,N_20050,N_21206);
nor U22039 (N_22039,N_21188,N_20334);
and U22040 (N_22040,N_21043,N_20190);
nand U22041 (N_22041,N_20374,N_20779);
xor U22042 (N_22042,N_21065,N_20916);
or U22043 (N_22043,N_20565,N_20011);
and U22044 (N_22044,N_20936,N_20462);
nor U22045 (N_22045,N_20354,N_20223);
nand U22046 (N_22046,N_21016,N_21128);
and U22047 (N_22047,N_20954,N_20503);
or U22048 (N_22048,N_20219,N_20002);
nor U22049 (N_22049,N_20504,N_20838);
nand U22050 (N_22050,N_20462,N_20388);
nor U22051 (N_22051,N_20803,N_20426);
or U22052 (N_22052,N_21036,N_20684);
nand U22053 (N_22053,N_20268,N_20203);
xnor U22054 (N_22054,N_20249,N_20568);
and U22055 (N_22055,N_20255,N_20160);
nor U22056 (N_22056,N_20481,N_20661);
and U22057 (N_22057,N_20827,N_20327);
and U22058 (N_22058,N_20891,N_20944);
nor U22059 (N_22059,N_20076,N_20141);
nand U22060 (N_22060,N_20037,N_21123);
and U22061 (N_22061,N_20379,N_20129);
or U22062 (N_22062,N_20096,N_20338);
or U22063 (N_22063,N_20056,N_21212);
nor U22064 (N_22064,N_20035,N_20090);
or U22065 (N_22065,N_20871,N_21051);
nand U22066 (N_22066,N_20841,N_21106);
or U22067 (N_22067,N_20829,N_20993);
nand U22068 (N_22068,N_20321,N_20544);
or U22069 (N_22069,N_20199,N_20931);
xnor U22070 (N_22070,N_21176,N_21143);
nor U22071 (N_22071,N_21060,N_20349);
nand U22072 (N_22072,N_20035,N_21144);
nor U22073 (N_22073,N_20434,N_20859);
nand U22074 (N_22074,N_20640,N_20053);
or U22075 (N_22075,N_20357,N_20788);
nor U22076 (N_22076,N_20768,N_20401);
nor U22077 (N_22077,N_20545,N_20827);
xor U22078 (N_22078,N_20304,N_20094);
nor U22079 (N_22079,N_20985,N_20096);
or U22080 (N_22080,N_21064,N_20051);
nand U22081 (N_22081,N_20194,N_20696);
nand U22082 (N_22082,N_20233,N_20157);
xor U22083 (N_22083,N_20799,N_20846);
xnor U22084 (N_22084,N_20350,N_20771);
and U22085 (N_22085,N_20341,N_20136);
or U22086 (N_22086,N_20029,N_21060);
and U22087 (N_22087,N_20734,N_20101);
nand U22088 (N_22088,N_20522,N_21149);
xnor U22089 (N_22089,N_20554,N_21237);
and U22090 (N_22090,N_20032,N_20775);
and U22091 (N_22091,N_21027,N_20077);
or U22092 (N_22092,N_20954,N_20894);
or U22093 (N_22093,N_21045,N_21096);
xor U22094 (N_22094,N_20966,N_20706);
nor U22095 (N_22095,N_20285,N_20955);
xor U22096 (N_22096,N_20025,N_21039);
xnor U22097 (N_22097,N_20860,N_20249);
or U22098 (N_22098,N_20543,N_20165);
nand U22099 (N_22099,N_20295,N_20397);
or U22100 (N_22100,N_20067,N_20858);
or U22101 (N_22101,N_20875,N_20833);
and U22102 (N_22102,N_20844,N_20556);
nor U22103 (N_22103,N_20376,N_20071);
nand U22104 (N_22104,N_20629,N_20591);
and U22105 (N_22105,N_20378,N_20032);
xnor U22106 (N_22106,N_20879,N_20657);
and U22107 (N_22107,N_20210,N_20116);
and U22108 (N_22108,N_20030,N_20018);
nand U22109 (N_22109,N_20588,N_20016);
nand U22110 (N_22110,N_20158,N_20459);
nor U22111 (N_22111,N_21114,N_21188);
nand U22112 (N_22112,N_21023,N_21099);
nand U22113 (N_22113,N_20344,N_20147);
and U22114 (N_22114,N_21027,N_20879);
nand U22115 (N_22115,N_21096,N_21066);
or U22116 (N_22116,N_20109,N_20065);
and U22117 (N_22117,N_20026,N_20357);
xnor U22118 (N_22118,N_21129,N_20123);
and U22119 (N_22119,N_20465,N_20134);
nand U22120 (N_22120,N_21010,N_20527);
nor U22121 (N_22121,N_21107,N_20416);
xnor U22122 (N_22122,N_20876,N_20590);
nand U22123 (N_22123,N_20035,N_20808);
xnor U22124 (N_22124,N_21036,N_20901);
xor U22125 (N_22125,N_21041,N_20197);
or U22126 (N_22126,N_20325,N_20534);
xor U22127 (N_22127,N_20923,N_20938);
xor U22128 (N_22128,N_21006,N_20344);
and U22129 (N_22129,N_20542,N_20618);
xor U22130 (N_22130,N_20380,N_20437);
xnor U22131 (N_22131,N_20107,N_21079);
and U22132 (N_22132,N_21184,N_21213);
and U22133 (N_22133,N_20434,N_20973);
or U22134 (N_22134,N_20866,N_20682);
nand U22135 (N_22135,N_20597,N_20266);
nor U22136 (N_22136,N_20718,N_20900);
xor U22137 (N_22137,N_20090,N_20301);
or U22138 (N_22138,N_20717,N_20819);
or U22139 (N_22139,N_20376,N_20864);
nand U22140 (N_22140,N_20903,N_20958);
and U22141 (N_22141,N_20939,N_21167);
nand U22142 (N_22142,N_20933,N_20975);
nand U22143 (N_22143,N_21207,N_20132);
xnor U22144 (N_22144,N_20441,N_20616);
or U22145 (N_22145,N_20877,N_20772);
nor U22146 (N_22146,N_20088,N_20795);
nand U22147 (N_22147,N_20139,N_20464);
or U22148 (N_22148,N_20369,N_20094);
xnor U22149 (N_22149,N_20737,N_21046);
nand U22150 (N_22150,N_20098,N_21189);
xnor U22151 (N_22151,N_20390,N_20264);
and U22152 (N_22152,N_20827,N_20845);
xnor U22153 (N_22153,N_21025,N_20320);
nor U22154 (N_22154,N_21158,N_20912);
nor U22155 (N_22155,N_20519,N_20959);
or U22156 (N_22156,N_20809,N_20692);
xor U22157 (N_22157,N_20313,N_20998);
nor U22158 (N_22158,N_20247,N_20121);
nor U22159 (N_22159,N_20866,N_20129);
nor U22160 (N_22160,N_21136,N_20508);
or U22161 (N_22161,N_20332,N_21245);
and U22162 (N_22162,N_20338,N_20521);
or U22163 (N_22163,N_21192,N_20155);
and U22164 (N_22164,N_20722,N_20665);
nor U22165 (N_22165,N_20973,N_21026);
nand U22166 (N_22166,N_20504,N_21009);
nor U22167 (N_22167,N_21157,N_20470);
nor U22168 (N_22168,N_20404,N_20490);
xor U22169 (N_22169,N_20000,N_20011);
and U22170 (N_22170,N_20820,N_20726);
nand U22171 (N_22171,N_21193,N_21243);
nand U22172 (N_22172,N_20477,N_20799);
nor U22173 (N_22173,N_20397,N_20930);
or U22174 (N_22174,N_20346,N_20649);
or U22175 (N_22175,N_21151,N_20814);
or U22176 (N_22176,N_20908,N_20680);
nor U22177 (N_22177,N_21236,N_20971);
xor U22178 (N_22178,N_21118,N_20347);
nand U22179 (N_22179,N_21116,N_21057);
nor U22180 (N_22180,N_21116,N_20476);
nor U22181 (N_22181,N_20385,N_20127);
xnor U22182 (N_22182,N_21138,N_21104);
and U22183 (N_22183,N_20950,N_20977);
nor U22184 (N_22184,N_20583,N_20581);
or U22185 (N_22185,N_20113,N_21069);
nand U22186 (N_22186,N_20147,N_21187);
nand U22187 (N_22187,N_21081,N_20115);
or U22188 (N_22188,N_20030,N_21003);
or U22189 (N_22189,N_20343,N_21028);
and U22190 (N_22190,N_20973,N_20128);
and U22191 (N_22191,N_21059,N_20592);
xor U22192 (N_22192,N_20639,N_20965);
nor U22193 (N_22193,N_20652,N_20620);
or U22194 (N_22194,N_20226,N_20748);
nand U22195 (N_22195,N_20094,N_20350);
and U22196 (N_22196,N_20163,N_20559);
nor U22197 (N_22197,N_20905,N_20242);
and U22198 (N_22198,N_20692,N_20523);
nor U22199 (N_22199,N_20215,N_20089);
nand U22200 (N_22200,N_20728,N_20894);
nor U22201 (N_22201,N_20747,N_20635);
and U22202 (N_22202,N_20877,N_20959);
nand U22203 (N_22203,N_20613,N_20022);
or U22204 (N_22204,N_20814,N_20318);
nand U22205 (N_22205,N_20854,N_20225);
nand U22206 (N_22206,N_20821,N_20936);
nand U22207 (N_22207,N_21194,N_20682);
and U22208 (N_22208,N_20032,N_20186);
nor U22209 (N_22209,N_21030,N_20314);
nor U22210 (N_22210,N_20072,N_20233);
nand U22211 (N_22211,N_20783,N_20987);
xor U22212 (N_22212,N_20737,N_20175);
and U22213 (N_22213,N_20217,N_21074);
or U22214 (N_22214,N_20200,N_20251);
and U22215 (N_22215,N_20597,N_20743);
nor U22216 (N_22216,N_20130,N_20395);
xnor U22217 (N_22217,N_20795,N_20377);
nand U22218 (N_22218,N_20959,N_20888);
nor U22219 (N_22219,N_20768,N_21001);
nand U22220 (N_22220,N_20817,N_20231);
or U22221 (N_22221,N_20461,N_20644);
nor U22222 (N_22222,N_20253,N_20416);
nor U22223 (N_22223,N_20371,N_20979);
xor U22224 (N_22224,N_20743,N_20144);
nor U22225 (N_22225,N_20748,N_20408);
nand U22226 (N_22226,N_20024,N_20675);
xnor U22227 (N_22227,N_20012,N_20042);
nand U22228 (N_22228,N_20386,N_20451);
and U22229 (N_22229,N_20953,N_20094);
or U22230 (N_22230,N_20338,N_20654);
and U22231 (N_22231,N_20797,N_21054);
and U22232 (N_22232,N_20825,N_20978);
nor U22233 (N_22233,N_20213,N_20060);
or U22234 (N_22234,N_21076,N_20687);
nand U22235 (N_22235,N_20349,N_20034);
nand U22236 (N_22236,N_20978,N_20020);
or U22237 (N_22237,N_20522,N_20588);
nand U22238 (N_22238,N_20225,N_20153);
or U22239 (N_22239,N_20443,N_21038);
nand U22240 (N_22240,N_21058,N_21037);
or U22241 (N_22241,N_21187,N_21163);
nor U22242 (N_22242,N_20461,N_20810);
nand U22243 (N_22243,N_21135,N_20015);
xor U22244 (N_22244,N_20195,N_20344);
or U22245 (N_22245,N_21205,N_20600);
and U22246 (N_22246,N_20400,N_20427);
nor U22247 (N_22247,N_20180,N_20139);
xnor U22248 (N_22248,N_20449,N_20991);
or U22249 (N_22249,N_21219,N_20416);
nand U22250 (N_22250,N_20494,N_20231);
and U22251 (N_22251,N_21059,N_20918);
nor U22252 (N_22252,N_20425,N_20285);
xor U22253 (N_22253,N_21247,N_20765);
nand U22254 (N_22254,N_20967,N_21151);
nand U22255 (N_22255,N_21030,N_20675);
or U22256 (N_22256,N_20365,N_20465);
nor U22257 (N_22257,N_20168,N_20810);
nor U22258 (N_22258,N_21003,N_20292);
or U22259 (N_22259,N_20343,N_20831);
and U22260 (N_22260,N_20399,N_20557);
and U22261 (N_22261,N_20543,N_20627);
nand U22262 (N_22262,N_20434,N_20791);
nor U22263 (N_22263,N_20994,N_20659);
nand U22264 (N_22264,N_20357,N_21179);
and U22265 (N_22265,N_20705,N_20278);
nor U22266 (N_22266,N_20702,N_20142);
or U22267 (N_22267,N_20261,N_20167);
xor U22268 (N_22268,N_20689,N_20927);
xor U22269 (N_22269,N_20364,N_20956);
nand U22270 (N_22270,N_20622,N_20177);
nor U22271 (N_22271,N_20779,N_20729);
nand U22272 (N_22272,N_20993,N_20928);
nor U22273 (N_22273,N_21191,N_20924);
and U22274 (N_22274,N_20009,N_20181);
and U22275 (N_22275,N_20349,N_20635);
or U22276 (N_22276,N_21139,N_20708);
nand U22277 (N_22277,N_21201,N_20985);
nor U22278 (N_22278,N_20969,N_21003);
and U22279 (N_22279,N_20439,N_20820);
xnor U22280 (N_22280,N_20077,N_20314);
or U22281 (N_22281,N_20225,N_21231);
or U22282 (N_22282,N_20374,N_20328);
and U22283 (N_22283,N_20962,N_20125);
and U22284 (N_22284,N_21184,N_20016);
xnor U22285 (N_22285,N_21231,N_20308);
or U22286 (N_22286,N_20655,N_21151);
nor U22287 (N_22287,N_21213,N_20303);
nand U22288 (N_22288,N_20360,N_20022);
or U22289 (N_22289,N_20731,N_20917);
nor U22290 (N_22290,N_20293,N_20496);
xor U22291 (N_22291,N_21088,N_20141);
nand U22292 (N_22292,N_20346,N_20508);
xor U22293 (N_22293,N_20260,N_21195);
xor U22294 (N_22294,N_20971,N_20976);
or U22295 (N_22295,N_20339,N_20821);
xor U22296 (N_22296,N_21162,N_21166);
or U22297 (N_22297,N_20847,N_20888);
or U22298 (N_22298,N_21119,N_20460);
nand U22299 (N_22299,N_21172,N_21033);
xor U22300 (N_22300,N_20074,N_20730);
nand U22301 (N_22301,N_20047,N_20807);
and U22302 (N_22302,N_20679,N_20600);
nand U22303 (N_22303,N_20196,N_20525);
nand U22304 (N_22304,N_21199,N_20288);
nor U22305 (N_22305,N_20442,N_20225);
xnor U22306 (N_22306,N_20942,N_20291);
nand U22307 (N_22307,N_21036,N_21242);
or U22308 (N_22308,N_20068,N_21188);
xnor U22309 (N_22309,N_20924,N_20161);
xnor U22310 (N_22310,N_20447,N_20524);
nand U22311 (N_22311,N_20767,N_21058);
and U22312 (N_22312,N_20234,N_21163);
xnor U22313 (N_22313,N_20856,N_20858);
nor U22314 (N_22314,N_20714,N_20512);
and U22315 (N_22315,N_20057,N_20101);
nand U22316 (N_22316,N_20963,N_20453);
xor U22317 (N_22317,N_20345,N_20530);
and U22318 (N_22318,N_20129,N_20647);
and U22319 (N_22319,N_20797,N_20979);
nand U22320 (N_22320,N_20667,N_20212);
xor U22321 (N_22321,N_20390,N_20125);
nor U22322 (N_22322,N_20273,N_20640);
or U22323 (N_22323,N_20777,N_21095);
or U22324 (N_22324,N_20374,N_20431);
or U22325 (N_22325,N_21227,N_21012);
and U22326 (N_22326,N_20293,N_20995);
xor U22327 (N_22327,N_20922,N_20464);
and U22328 (N_22328,N_20737,N_20591);
or U22329 (N_22329,N_20785,N_20206);
nand U22330 (N_22330,N_20144,N_21219);
and U22331 (N_22331,N_20015,N_21133);
and U22332 (N_22332,N_21152,N_20822);
and U22333 (N_22333,N_21107,N_21204);
nand U22334 (N_22334,N_20266,N_20603);
or U22335 (N_22335,N_20963,N_20688);
xor U22336 (N_22336,N_20849,N_20130);
nor U22337 (N_22337,N_20881,N_20062);
nor U22338 (N_22338,N_20916,N_20428);
or U22339 (N_22339,N_20637,N_20538);
nand U22340 (N_22340,N_20597,N_20474);
nand U22341 (N_22341,N_20138,N_20284);
nand U22342 (N_22342,N_20390,N_20438);
nor U22343 (N_22343,N_21135,N_20912);
and U22344 (N_22344,N_20255,N_20091);
or U22345 (N_22345,N_20427,N_20148);
or U22346 (N_22346,N_20660,N_20640);
or U22347 (N_22347,N_21249,N_20410);
and U22348 (N_22348,N_20826,N_20599);
nor U22349 (N_22349,N_20104,N_20628);
nor U22350 (N_22350,N_20074,N_20686);
nand U22351 (N_22351,N_20473,N_20275);
xnor U22352 (N_22352,N_20408,N_20943);
nand U22353 (N_22353,N_20529,N_20279);
xor U22354 (N_22354,N_20560,N_20200);
nand U22355 (N_22355,N_20728,N_20413);
xnor U22356 (N_22356,N_20906,N_20541);
xnor U22357 (N_22357,N_21206,N_21004);
xor U22358 (N_22358,N_20136,N_20816);
and U22359 (N_22359,N_21218,N_20918);
and U22360 (N_22360,N_20670,N_20449);
xor U22361 (N_22361,N_20174,N_20524);
nor U22362 (N_22362,N_20300,N_20055);
nor U22363 (N_22363,N_20521,N_21110);
nor U22364 (N_22364,N_20956,N_20790);
nand U22365 (N_22365,N_21184,N_21003);
or U22366 (N_22366,N_20492,N_20882);
xnor U22367 (N_22367,N_20944,N_21194);
xor U22368 (N_22368,N_20259,N_21087);
xor U22369 (N_22369,N_20345,N_20910);
and U22370 (N_22370,N_20729,N_20131);
or U22371 (N_22371,N_20872,N_20583);
and U22372 (N_22372,N_20430,N_20289);
and U22373 (N_22373,N_20672,N_20309);
nand U22374 (N_22374,N_21069,N_20994);
or U22375 (N_22375,N_20597,N_20027);
xor U22376 (N_22376,N_21055,N_20269);
and U22377 (N_22377,N_20882,N_20489);
or U22378 (N_22378,N_20213,N_21235);
and U22379 (N_22379,N_20349,N_20373);
xnor U22380 (N_22380,N_20585,N_20362);
or U22381 (N_22381,N_20517,N_20115);
xnor U22382 (N_22382,N_20491,N_20479);
or U22383 (N_22383,N_21034,N_21189);
nor U22384 (N_22384,N_20983,N_20320);
or U22385 (N_22385,N_20474,N_20093);
or U22386 (N_22386,N_21233,N_20453);
nor U22387 (N_22387,N_20766,N_21085);
nor U22388 (N_22388,N_20527,N_20824);
nor U22389 (N_22389,N_21010,N_20654);
nor U22390 (N_22390,N_20886,N_20557);
and U22391 (N_22391,N_20583,N_20164);
and U22392 (N_22392,N_20971,N_20881);
nand U22393 (N_22393,N_21208,N_20625);
xor U22394 (N_22394,N_20559,N_20483);
nor U22395 (N_22395,N_20583,N_21120);
or U22396 (N_22396,N_20895,N_21234);
and U22397 (N_22397,N_21183,N_20425);
and U22398 (N_22398,N_20296,N_21088);
nor U22399 (N_22399,N_20114,N_20318);
and U22400 (N_22400,N_20650,N_20529);
nor U22401 (N_22401,N_20147,N_20500);
or U22402 (N_22402,N_20977,N_20206);
nand U22403 (N_22403,N_20045,N_20484);
or U22404 (N_22404,N_21038,N_20811);
nor U22405 (N_22405,N_20252,N_20698);
nand U22406 (N_22406,N_20865,N_20964);
nor U22407 (N_22407,N_20646,N_21129);
nand U22408 (N_22408,N_20848,N_20275);
and U22409 (N_22409,N_20691,N_20291);
xnor U22410 (N_22410,N_20530,N_20951);
and U22411 (N_22411,N_20764,N_20967);
nand U22412 (N_22412,N_21234,N_20859);
or U22413 (N_22413,N_20837,N_20122);
and U22414 (N_22414,N_20097,N_20144);
or U22415 (N_22415,N_21210,N_20320);
and U22416 (N_22416,N_21010,N_21056);
nand U22417 (N_22417,N_20218,N_20579);
xnor U22418 (N_22418,N_21246,N_20281);
and U22419 (N_22419,N_20439,N_20966);
nand U22420 (N_22420,N_20495,N_21116);
or U22421 (N_22421,N_20091,N_20970);
and U22422 (N_22422,N_20471,N_20557);
nand U22423 (N_22423,N_20588,N_20948);
nor U22424 (N_22424,N_20234,N_20509);
nand U22425 (N_22425,N_21132,N_20831);
and U22426 (N_22426,N_20892,N_21104);
and U22427 (N_22427,N_20953,N_20984);
and U22428 (N_22428,N_20930,N_20950);
xnor U22429 (N_22429,N_20192,N_20804);
nand U22430 (N_22430,N_20437,N_20504);
and U22431 (N_22431,N_20306,N_20243);
xor U22432 (N_22432,N_20385,N_21224);
nand U22433 (N_22433,N_20908,N_20875);
nor U22434 (N_22434,N_20758,N_20554);
xnor U22435 (N_22435,N_20380,N_20806);
or U22436 (N_22436,N_20925,N_21062);
or U22437 (N_22437,N_21101,N_20783);
xnor U22438 (N_22438,N_21129,N_20744);
or U22439 (N_22439,N_21236,N_20906);
xor U22440 (N_22440,N_20999,N_20876);
nand U22441 (N_22441,N_20373,N_21232);
nand U22442 (N_22442,N_21244,N_20599);
and U22443 (N_22443,N_21166,N_20713);
nor U22444 (N_22444,N_20268,N_20014);
and U22445 (N_22445,N_20480,N_20477);
and U22446 (N_22446,N_20252,N_20357);
xnor U22447 (N_22447,N_20033,N_20149);
nor U22448 (N_22448,N_20990,N_20794);
xor U22449 (N_22449,N_20858,N_20766);
nor U22450 (N_22450,N_20551,N_20554);
xor U22451 (N_22451,N_21116,N_20955);
xnor U22452 (N_22452,N_20117,N_20542);
and U22453 (N_22453,N_20423,N_20058);
or U22454 (N_22454,N_20894,N_21079);
xor U22455 (N_22455,N_20956,N_20544);
or U22456 (N_22456,N_21039,N_20918);
xor U22457 (N_22457,N_20514,N_20649);
or U22458 (N_22458,N_20044,N_20578);
and U22459 (N_22459,N_20494,N_21039);
nor U22460 (N_22460,N_20372,N_20401);
nor U22461 (N_22461,N_20965,N_20651);
nor U22462 (N_22462,N_20404,N_20102);
nor U22463 (N_22463,N_20800,N_20003);
and U22464 (N_22464,N_21013,N_20099);
xnor U22465 (N_22465,N_20368,N_20688);
xnor U22466 (N_22466,N_20626,N_21176);
or U22467 (N_22467,N_21161,N_20151);
xnor U22468 (N_22468,N_20305,N_21059);
and U22469 (N_22469,N_20697,N_20304);
nor U22470 (N_22470,N_20808,N_20780);
xor U22471 (N_22471,N_20849,N_20653);
or U22472 (N_22472,N_21084,N_20959);
and U22473 (N_22473,N_20936,N_20855);
xnor U22474 (N_22474,N_20262,N_21222);
or U22475 (N_22475,N_20151,N_20891);
or U22476 (N_22476,N_21151,N_20787);
nor U22477 (N_22477,N_21197,N_20561);
xor U22478 (N_22478,N_20676,N_20041);
nand U22479 (N_22479,N_20505,N_21192);
nor U22480 (N_22480,N_20510,N_20211);
and U22481 (N_22481,N_21040,N_20774);
xnor U22482 (N_22482,N_21188,N_20836);
or U22483 (N_22483,N_20250,N_20176);
xnor U22484 (N_22484,N_20032,N_21212);
or U22485 (N_22485,N_21192,N_20588);
and U22486 (N_22486,N_21064,N_20193);
and U22487 (N_22487,N_21091,N_20240);
nand U22488 (N_22488,N_20086,N_21145);
xor U22489 (N_22489,N_20449,N_20788);
xor U22490 (N_22490,N_20118,N_20714);
nand U22491 (N_22491,N_20950,N_20067);
and U22492 (N_22492,N_20974,N_20541);
nand U22493 (N_22493,N_21154,N_20487);
xor U22494 (N_22494,N_20808,N_20265);
nand U22495 (N_22495,N_20079,N_20686);
nand U22496 (N_22496,N_20222,N_20572);
xnor U22497 (N_22497,N_21119,N_20828);
and U22498 (N_22498,N_20198,N_21049);
xor U22499 (N_22499,N_20573,N_20114);
nor U22500 (N_22500,N_21815,N_21601);
or U22501 (N_22501,N_22291,N_22445);
nand U22502 (N_22502,N_21623,N_22127);
nand U22503 (N_22503,N_22134,N_21403);
xnor U22504 (N_22504,N_22397,N_22155);
nand U22505 (N_22505,N_22376,N_21955);
and U22506 (N_22506,N_21859,N_22130);
or U22507 (N_22507,N_22411,N_21832);
or U22508 (N_22508,N_22432,N_21582);
xnor U22509 (N_22509,N_21747,N_22153);
and U22510 (N_22510,N_22164,N_22324);
and U22511 (N_22511,N_21847,N_21373);
nand U22512 (N_22512,N_22296,N_21417);
nor U22513 (N_22513,N_21502,N_22298);
xnor U22514 (N_22514,N_22096,N_21897);
xnor U22515 (N_22515,N_21345,N_21267);
nor U22516 (N_22516,N_22193,N_22477);
and U22517 (N_22517,N_22160,N_22489);
nand U22518 (N_22518,N_21740,N_22143);
and U22519 (N_22519,N_21867,N_22207);
nand U22520 (N_22520,N_21387,N_21394);
or U22521 (N_22521,N_22255,N_22354);
nor U22522 (N_22522,N_21320,N_21351);
xor U22523 (N_22523,N_21324,N_21588);
and U22524 (N_22524,N_21951,N_21873);
nor U22525 (N_22525,N_22105,N_21457);
and U22526 (N_22526,N_21608,N_22034);
nor U22527 (N_22527,N_22108,N_21471);
and U22528 (N_22528,N_22450,N_22212);
xor U22529 (N_22529,N_22389,N_21923);
and U22530 (N_22530,N_21722,N_21377);
or U22531 (N_22531,N_21359,N_21280);
or U22532 (N_22532,N_21657,N_21890);
or U22533 (N_22533,N_21789,N_21906);
nand U22534 (N_22534,N_21428,N_22455);
xnor U22535 (N_22535,N_22236,N_22433);
or U22536 (N_22536,N_22270,N_21975);
and U22537 (N_22537,N_22112,N_21449);
or U22538 (N_22538,N_22006,N_21261);
and U22539 (N_22539,N_21574,N_21983);
or U22540 (N_22540,N_21704,N_22303);
xnor U22541 (N_22541,N_22037,N_21754);
and U22542 (N_22542,N_21928,N_21777);
or U22543 (N_22543,N_22073,N_22075);
nand U22544 (N_22544,N_21609,N_21396);
nor U22545 (N_22545,N_22356,N_21862);
nor U22546 (N_22546,N_22222,N_21468);
or U22547 (N_22547,N_22008,N_22497);
xnor U22548 (N_22548,N_22406,N_22196);
and U22549 (N_22549,N_21452,N_22003);
xnor U22550 (N_22550,N_22259,N_21697);
nand U22551 (N_22551,N_22069,N_22430);
xor U22552 (N_22552,N_22007,N_22090);
nor U22553 (N_22553,N_22474,N_21826);
xnor U22554 (N_22554,N_22024,N_21378);
xnor U22555 (N_22555,N_21593,N_22307);
or U22556 (N_22556,N_21968,N_21866);
xor U22557 (N_22557,N_21986,N_21820);
and U22558 (N_22558,N_22272,N_22465);
and U22559 (N_22559,N_22436,N_22391);
or U22560 (N_22560,N_21773,N_22039);
or U22561 (N_22561,N_22103,N_22152);
or U22562 (N_22562,N_22056,N_22388);
and U22563 (N_22563,N_21446,N_22149);
nor U22564 (N_22564,N_21413,N_21605);
nand U22565 (N_22565,N_21656,N_21993);
xnor U22566 (N_22566,N_22263,N_22125);
nor U22567 (N_22567,N_22161,N_21586);
and U22568 (N_22568,N_21361,N_22137);
nand U22569 (N_22569,N_22215,N_22329);
xor U22570 (N_22570,N_22022,N_22343);
and U22571 (N_22571,N_21627,N_21891);
nor U22572 (N_22572,N_21776,N_21271);
nor U22573 (N_22573,N_22363,N_21505);
or U22574 (N_22574,N_21520,N_21333);
nor U22575 (N_22575,N_21787,N_21762);
xnor U22576 (N_22576,N_22361,N_21684);
or U22577 (N_22577,N_21870,N_22079);
nor U22578 (N_22578,N_21444,N_21934);
nand U22579 (N_22579,N_21781,N_22029);
nor U22580 (N_22580,N_22490,N_21901);
and U22581 (N_22581,N_21381,N_21801);
or U22582 (N_22582,N_22439,N_22470);
nor U22583 (N_22583,N_21759,N_22114);
xor U22584 (N_22584,N_22131,N_22216);
or U22585 (N_22585,N_22063,N_21878);
nor U22586 (N_22586,N_22262,N_22309);
and U22587 (N_22587,N_21827,N_22086);
xor U22588 (N_22588,N_22281,N_22087);
nand U22589 (N_22589,N_21569,N_21472);
nor U22590 (N_22590,N_21648,N_22081);
nor U22591 (N_22591,N_21914,N_22248);
nor U22592 (N_22592,N_21994,N_22026);
nand U22593 (N_22593,N_21304,N_21598);
nand U22594 (N_22594,N_22239,N_22488);
or U22595 (N_22595,N_21370,N_21407);
xor U22596 (N_22596,N_21703,N_22032);
or U22597 (N_22597,N_21539,N_21688);
nand U22598 (N_22598,N_22060,N_22165);
or U22599 (N_22599,N_22288,N_22448);
and U22600 (N_22600,N_21291,N_21322);
nand U22601 (N_22601,N_22487,N_21455);
nor U22602 (N_22602,N_22254,N_21990);
xor U22603 (N_22603,N_21266,N_22364);
nor U22604 (N_22604,N_22118,N_21872);
and U22605 (N_22605,N_21343,N_21474);
nand U22606 (N_22606,N_22201,N_21695);
or U22607 (N_22607,N_21786,N_21985);
nand U22608 (N_22608,N_21888,N_21828);
nor U22609 (N_22609,N_21745,N_21255);
nor U22610 (N_22610,N_22192,N_21876);
and U22611 (N_22611,N_22300,N_21426);
and U22612 (N_22612,N_22396,N_21950);
and U22613 (N_22613,N_22195,N_21450);
xor U22614 (N_22614,N_21479,N_21699);
or U22615 (N_22615,N_22355,N_22325);
and U22616 (N_22616,N_21709,N_21963);
and U22617 (N_22617,N_22018,N_21935);
or U22618 (N_22618,N_22269,N_22171);
and U22619 (N_22619,N_21356,N_21433);
and U22620 (N_22620,N_22419,N_21431);
xor U22621 (N_22621,N_21738,N_21250);
or U22622 (N_22622,N_22250,N_22413);
nor U22623 (N_22623,N_21438,N_21631);
xor U22624 (N_22624,N_21701,N_21440);
nand U22625 (N_22625,N_22338,N_22326);
nand U22626 (N_22626,N_21743,N_21830);
and U22627 (N_22627,N_21554,N_21253);
nand U22628 (N_22628,N_21655,N_21865);
and U22629 (N_22629,N_21406,N_21547);
nor U22630 (N_22630,N_21264,N_21691);
nand U22631 (N_22631,N_22228,N_21595);
and U22632 (N_22632,N_21354,N_21382);
nand U22633 (N_22633,N_21578,N_21780);
nand U22634 (N_22634,N_21817,N_22030);
nand U22635 (N_22635,N_21819,N_21682);
xnor U22636 (N_22636,N_22418,N_21422);
and U22637 (N_22637,N_21590,N_21610);
xnor U22638 (N_22638,N_21947,N_22074);
and U22639 (N_22639,N_22457,N_22144);
and U22640 (N_22640,N_21760,N_21334);
nand U22641 (N_22641,N_21685,N_21721);
and U22642 (N_22642,N_21362,N_22374);
or U22643 (N_22643,N_21849,N_22206);
nor U22644 (N_22644,N_21638,N_21579);
xnor U22645 (N_22645,N_21366,N_21969);
xor U22646 (N_22646,N_22186,N_22466);
and U22647 (N_22647,N_21339,N_21730);
and U22648 (N_22648,N_22264,N_21690);
nor U22649 (N_22649,N_21411,N_22452);
or U22650 (N_22650,N_22234,N_21957);
or U22651 (N_22651,N_21725,N_22058);
or U22652 (N_22652,N_22014,N_21643);
nand U22653 (N_22653,N_22182,N_21739);
xnor U22654 (N_22654,N_22187,N_21272);
nand U22655 (N_22655,N_21924,N_22252);
nor U22656 (N_22656,N_22221,N_21309);
or U22657 (N_22657,N_21812,N_21880);
nand U22658 (N_22658,N_22438,N_22481);
nor U22659 (N_22659,N_22210,N_21400);
nand U22660 (N_22660,N_22282,N_22373);
xnor U22661 (N_22661,N_22240,N_21732);
or U22662 (N_22662,N_21645,N_22175);
or U22663 (N_22663,N_21348,N_21278);
nand U22664 (N_22664,N_21894,N_21907);
nor U22665 (N_22665,N_21537,N_21794);
xnor U22666 (N_22666,N_21713,N_21485);
and U22667 (N_22667,N_21622,N_22100);
and U22668 (N_22668,N_21296,N_21774);
and U22669 (N_22669,N_22181,N_22398);
nand U22670 (N_22670,N_21613,N_22168);
xnor U22671 (N_22671,N_22395,N_22021);
and U22672 (N_22672,N_21338,N_22336);
xor U22673 (N_22673,N_22287,N_21617);
nor U22674 (N_22674,N_22004,N_21825);
nand U22675 (N_22675,N_22279,N_21599);
or U22676 (N_22676,N_22468,N_21409);
xor U22677 (N_22677,N_22019,N_21821);
nor U22678 (N_22678,N_21669,N_21911);
xnor U22679 (N_22679,N_21534,N_21694);
xnor U22680 (N_22680,N_21629,N_21757);
xnor U22681 (N_22681,N_22478,N_21833);
or U22682 (N_22682,N_22121,N_21735);
xor U22683 (N_22683,N_22486,N_21602);
or U22684 (N_22684,N_21842,N_21478);
nand U22685 (N_22685,N_21681,N_22484);
nor U22686 (N_22686,N_22188,N_22244);
and U22687 (N_22687,N_22273,N_22495);
or U22688 (N_22688,N_22491,N_21712);
and U22689 (N_22689,N_22426,N_21458);
nor U22690 (N_22690,N_21503,N_21494);
nand U22691 (N_22691,N_22253,N_21767);
and U22692 (N_22692,N_22427,N_21900);
and U22693 (N_22693,N_21480,N_22237);
or U22694 (N_22694,N_22015,N_22055);
xor U22695 (N_22695,N_21270,N_22463);
nand U22696 (N_22696,N_21380,N_21427);
or U22697 (N_22697,N_22294,N_21625);
and U22698 (N_22698,N_22315,N_21606);
xnor U22699 (N_22699,N_21672,N_22367);
and U22700 (N_22700,N_21414,N_21649);
or U22701 (N_22701,N_22095,N_21577);
nand U22702 (N_22702,N_21654,N_21966);
or U22703 (N_22703,N_21670,N_22337);
and U22704 (N_22704,N_21429,N_21834);
or U22705 (N_22705,N_21949,N_22366);
nor U22706 (N_22706,N_22459,N_22229);
or U22707 (N_22707,N_21453,N_22085);
xor U22708 (N_22708,N_22099,N_21557);
or U22709 (N_22709,N_22425,N_21932);
nand U22710 (N_22710,N_21904,N_22010);
or U22711 (N_22711,N_21799,N_21254);
xor U22712 (N_22712,N_21916,N_21889);
nor U22713 (N_22713,N_22328,N_22214);
and U22714 (N_22714,N_21504,N_21368);
nand U22715 (N_22715,N_22046,N_22173);
and U22716 (N_22716,N_21424,N_21899);
or U22717 (N_22717,N_22375,N_21528);
xnor U22718 (N_22718,N_22322,N_21954);
nor U22719 (N_22719,N_22286,N_21829);
nor U22720 (N_22720,N_22381,N_21437);
xor U22721 (N_22721,N_21727,N_21441);
nand U22722 (N_22722,N_22483,N_22176);
nand U22723 (N_22723,N_21972,N_22041);
nor U22724 (N_22724,N_22423,N_21328);
xnor U22725 (N_22725,N_21553,N_22265);
xnor U22726 (N_22726,N_21882,N_21454);
xnor U22727 (N_22727,N_21555,N_21813);
or U22728 (N_22728,N_21715,N_21410);
or U22729 (N_22729,N_21665,N_21663);
or U22730 (N_22730,N_22156,N_22128);
nor U22731 (N_22731,N_21772,N_21807);
nor U22732 (N_22732,N_21519,N_22420);
and U22733 (N_22733,N_22437,N_21252);
nor U22734 (N_22734,N_21319,N_22399);
or U22735 (N_22735,N_22382,N_21848);
nor U22736 (N_22736,N_22431,N_21310);
xnor U22737 (N_22737,N_21383,N_21895);
nand U22738 (N_22738,N_21615,N_21942);
nand U22739 (N_22739,N_21967,N_21439);
or U22740 (N_22740,N_21290,N_21512);
or U22741 (N_22741,N_22005,N_21775);
or U22742 (N_22742,N_22219,N_21768);
nor U22743 (N_22743,N_22313,N_21293);
and U22744 (N_22744,N_22059,N_21415);
xnor U22745 (N_22745,N_21784,N_21265);
nor U22746 (N_22746,N_22368,N_22461);
and U22747 (N_22747,N_22429,N_21612);
xor U22748 (N_22748,N_22049,N_22480);
and U22749 (N_22749,N_22141,N_21341);
or U22750 (N_22750,N_21477,N_22482);
nand U22751 (N_22751,N_21536,N_22362);
nor U22752 (N_22752,N_22306,N_22327);
xnor U22753 (N_22753,N_21347,N_21281);
xnor U22754 (N_22754,N_21525,N_22302);
xnor U22755 (N_22755,N_22353,N_21560);
nor U22756 (N_22756,N_22148,N_22068);
nor U22757 (N_22757,N_22401,N_21896);
and U22758 (N_22758,N_21771,N_22280);
nand U22759 (N_22759,N_21482,N_22017);
xor U22760 (N_22760,N_22054,N_21596);
nand U22761 (N_22761,N_21822,N_21918);
and U22762 (N_22762,N_22066,N_22077);
and U22763 (N_22763,N_22124,N_21447);
xor U22764 (N_22764,N_21902,N_21552);
or U22765 (N_22765,N_21311,N_21700);
nor U22766 (N_22766,N_22135,N_22371);
nand U22767 (N_22767,N_21836,N_21506);
nor U22768 (N_22768,N_22479,N_21679);
xnor U22769 (N_22769,N_22405,N_22276);
or U22770 (N_22770,N_22251,N_22266);
xor U22771 (N_22771,N_21929,N_22347);
and U22772 (N_22772,N_22205,N_22035);
or U22773 (N_22773,N_21464,N_21706);
or U22774 (N_22774,N_21761,N_21524);
xor U22775 (N_22775,N_21943,N_22416);
and U22776 (N_22776,N_21289,N_21515);
nand U22777 (N_22777,N_21435,N_21332);
or U22778 (N_22778,N_21877,N_21997);
nor U22779 (N_22779,N_21542,N_22258);
or U22780 (N_22780,N_21999,N_21869);
and U22781 (N_22781,N_21910,N_21664);
nand U22782 (N_22782,N_21687,N_22123);
and U22783 (N_22783,N_22238,N_22031);
xnor U22784 (N_22784,N_22136,N_22002);
nor U22785 (N_22785,N_21353,N_22417);
nor U22786 (N_22786,N_22047,N_21941);
nand U22787 (N_22787,N_21750,N_22027);
or U22788 (N_22788,N_21499,N_21667);
xnor U22789 (N_22789,N_22352,N_21755);
nand U22790 (N_22790,N_21445,N_21979);
and U22791 (N_22791,N_21329,N_22456);
xor U22792 (N_22792,N_21974,N_22412);
nor U22793 (N_22793,N_21920,N_21418);
nor U22794 (N_22794,N_21840,N_21260);
or U22795 (N_22795,N_21589,N_22045);
and U22796 (N_22796,N_21874,N_21591);
nor U22797 (N_22797,N_22267,N_22292);
nand U22798 (N_22798,N_22284,N_21634);
xor U22799 (N_22799,N_22320,N_22089);
nor U22800 (N_22800,N_21996,N_21526);
nor U22801 (N_22801,N_21374,N_21970);
and U22802 (N_22802,N_21484,N_21719);
xor U22803 (N_22803,N_21714,N_21850);
nor U22804 (N_22804,N_22469,N_21611);
or U22805 (N_22805,N_22076,N_21321);
or U22806 (N_22806,N_22393,N_22243);
xnor U22807 (N_22807,N_21973,N_21733);
nand U22808 (N_22808,N_22458,N_22183);
and U22809 (N_22809,N_22211,N_22194);
and U22810 (N_22810,N_21731,N_22370);
nor U22811 (N_22811,N_21548,N_21887);
nor U22812 (N_22812,N_21393,N_21386);
and U22813 (N_22813,N_21742,N_21436);
and U22814 (N_22814,N_21769,N_22120);
nand U22815 (N_22815,N_21395,N_21313);
or U22816 (N_22816,N_22138,N_21269);
nand U22817 (N_22817,N_22116,N_22231);
xnor U22818 (N_22818,N_21335,N_22422);
and U22819 (N_22819,N_21937,N_21442);
and U22820 (N_22820,N_21371,N_21259);
xor U22821 (N_22821,N_21841,N_22177);
xnor U22822 (N_22822,N_21856,N_22312);
xor U22823 (N_22823,N_21300,N_22051);
or U22824 (N_22824,N_21718,N_21987);
nor U22825 (N_22825,N_21603,N_22330);
nor U22826 (N_22826,N_21984,N_21823);
nand U22827 (N_22827,N_21401,N_22033);
or U22828 (N_22828,N_21746,N_21563);
nand U22829 (N_22829,N_21388,N_22295);
and U22830 (N_22830,N_21274,N_22385);
nor U22831 (N_22831,N_21758,N_22072);
nor U22832 (N_22832,N_21469,N_22308);
nand U22833 (N_22833,N_21340,N_21675);
nor U22834 (N_22834,N_21922,N_22208);
and U22835 (N_22835,N_21342,N_21948);
nand U22836 (N_22836,N_22434,N_21831);
and U22837 (N_22837,N_22174,N_22224);
xor U22838 (N_22838,N_21953,N_22394);
nor U22839 (N_22839,N_21796,N_21299);
nor U22840 (N_22840,N_21898,N_21544);
nor U22841 (N_22841,N_21276,N_21778);
nand U22842 (N_22842,N_21964,N_21488);
or U22843 (N_22843,N_21297,N_22189);
or U22844 (N_22844,N_21470,N_21496);
nor U22845 (N_22845,N_21462,N_21500);
nor U22846 (N_22846,N_21302,N_21365);
nand U22847 (N_22847,N_22092,N_21282);
xnor U22848 (N_22848,N_21835,N_21360);
or U22849 (N_22849,N_21931,N_21369);
xnor U22850 (N_22850,N_22197,N_21573);
nand U22851 (N_22851,N_21881,N_22129);
nand U22852 (N_22852,N_22365,N_21692);
nand U22853 (N_22853,N_21392,N_21710);
and U22854 (N_22854,N_22345,N_21845);
nand U22855 (N_22855,N_21811,N_21644);
nor U22856 (N_22856,N_21419,N_22159);
nor U22857 (N_22857,N_21491,N_21521);
and U22858 (N_22858,N_22335,N_21952);
nor U22859 (N_22859,N_22256,N_22453);
nor U22860 (N_22860,N_22157,N_22191);
nor U22861 (N_22861,N_21977,N_22261);
xor U22862 (N_22862,N_22475,N_21884);
xnor U22863 (N_22863,N_22245,N_21465);
and U22864 (N_22864,N_21661,N_22146);
and U22865 (N_22865,N_22400,N_21459);
nand U22866 (N_22866,N_21337,N_21284);
or U22867 (N_22867,N_21683,N_22492);
nor U22868 (N_22868,N_21531,N_21632);
or U22869 (N_22869,N_21398,N_21614);
or U22870 (N_22870,N_22223,N_21618);
nand U22871 (N_22871,N_21782,N_22443);
and U22872 (N_22872,N_21513,N_22025);
and U22873 (N_22873,N_21391,N_21666);
and U22874 (N_22874,N_22467,N_22064);
or U22875 (N_22875,N_22209,N_22299);
or U22876 (N_22876,N_21346,N_21995);
nand U22877 (N_22877,N_22233,N_21273);
nand U22878 (N_22878,N_21641,N_21660);
and U22879 (N_22879,N_22106,N_21998);
or U22880 (N_22880,N_21808,N_22230);
nand U22881 (N_22881,N_22020,N_21844);
or U22882 (N_22882,N_21938,N_22053);
nor U22883 (N_22883,N_22369,N_21853);
and U22884 (N_22884,N_21514,N_21893);
xnor U22885 (N_22885,N_22304,N_21567);
xor U22886 (N_22886,N_21659,N_21860);
xor U22887 (N_22887,N_21662,N_22257);
and U22888 (N_22888,N_21357,N_21384);
or U22889 (N_22889,N_21716,N_22318);
nor U22890 (N_22890,N_22036,N_22204);
and U22891 (N_22891,N_22009,N_22331);
nand U22892 (N_22892,N_21909,N_21568);
nor U22893 (N_22893,N_21420,N_21456);
or U22894 (N_22894,N_21564,N_22428);
and U22895 (N_22895,N_21508,N_21723);
xnor U22896 (N_22896,N_21978,N_22494);
nor U22897 (N_22897,N_22050,N_21795);
and U22898 (N_22898,N_22260,N_22088);
and U22899 (N_22899,N_21432,N_21779);
nand U22900 (N_22900,N_21314,N_22408);
or U22901 (N_22901,N_21763,N_22104);
or U22902 (N_22902,N_21676,N_21805);
nor U22903 (N_22903,N_21298,N_21961);
nand U22904 (N_22904,N_21275,N_21301);
or U22905 (N_22905,N_22000,N_22348);
or U22906 (N_22906,N_21336,N_22150);
or U22907 (N_22907,N_21358,N_21792);
or U22908 (N_22908,N_21650,N_21770);
or U22909 (N_22909,N_22132,N_21594);
xnor U22910 (N_22910,N_21855,N_21803);
xnor U22911 (N_22911,N_21868,N_21425);
or U22912 (N_22912,N_21277,N_21863);
nor U22913 (N_22913,N_21824,N_21389);
or U22914 (N_22914,N_21326,N_22349);
nand U22915 (N_22915,N_21570,N_21495);
or U22916 (N_22916,N_22140,N_21646);
nand U22917 (N_22917,N_22323,N_22390);
xor U22918 (N_22918,N_21892,N_22093);
and U22919 (N_22919,N_21680,N_21652);
nand U22920 (N_22920,N_21405,N_22246);
nand U22921 (N_22921,N_21604,N_21693);
xnor U22922 (N_22922,N_21698,N_21636);
nand U22923 (N_22923,N_21330,N_22440);
xor U22924 (N_22924,N_22447,N_21621);
nor U22925 (N_22925,N_21858,N_22271);
and U22926 (N_22926,N_22070,N_22464);
xor U22927 (N_22927,N_21487,N_21905);
or U22928 (N_22928,N_22115,N_22359);
nand U22929 (N_22929,N_21489,N_21734);
nand U22930 (N_22930,N_22065,N_22200);
or U22931 (N_22931,N_21546,N_22091);
and U22932 (N_22932,N_21635,N_22471);
xnor U22933 (N_22933,N_22111,N_21592);
nand U22934 (N_22934,N_22454,N_22451);
nand U22935 (N_22935,N_21535,N_21790);
nor U22936 (N_22936,N_21283,N_22179);
xor U22937 (N_22937,N_22344,N_21989);
and U22938 (N_22938,N_22442,N_21375);
and U22939 (N_22939,N_21965,N_21559);
xnor U22940 (N_22940,N_22167,N_21286);
and U22941 (N_22941,N_21992,N_21507);
nand U22942 (N_22942,N_22071,N_22202);
nor U22943 (N_22943,N_21885,N_21466);
nand U22944 (N_22944,N_22225,N_21268);
nor U22945 (N_22945,N_22218,N_22380);
nand U22946 (N_22946,N_21443,N_21558);
and U22947 (N_22947,N_21527,N_22403);
and U22948 (N_22948,N_21331,N_21960);
or U22949 (N_22949,N_22404,N_22162);
xor U22950 (N_22950,N_21363,N_22184);
nand U22951 (N_22951,N_21809,N_21658);
or U22952 (N_22952,N_21344,N_22078);
nand U22953 (N_22953,N_21571,N_21350);
nor U22954 (N_22954,N_21587,N_21430);
and U22955 (N_22955,N_21944,N_21279);
or U22956 (N_22956,N_21736,N_22449);
or U22957 (N_22957,N_21251,N_21707);
nor U22958 (N_22958,N_21945,N_22067);
or U22959 (N_22959,N_21461,N_22379);
or U22960 (N_22960,N_21483,N_22460);
or U22961 (N_22961,N_22415,N_21919);
nor U22962 (N_22962,N_22158,N_22062);
xor U22963 (N_22963,N_22473,N_21633);
or U22964 (N_22964,N_21473,N_21257);
or U22965 (N_22965,N_22305,N_21843);
nand U22966 (N_22966,N_22274,N_22057);
or U22967 (N_22967,N_21543,N_21991);
or U22968 (N_22968,N_22061,N_22317);
nand U22969 (N_22969,N_21576,N_21448);
xor U22970 (N_22970,N_21616,N_21785);
xnor U22971 (N_22971,N_21864,N_21915);
or U22972 (N_22972,N_21501,N_21753);
nand U22973 (N_22973,N_21263,N_21804);
nand U22974 (N_22974,N_21946,N_21256);
or U22975 (N_22975,N_21674,N_21717);
and U22976 (N_22976,N_22082,N_21791);
nand U22977 (N_22977,N_22185,N_21705);
xor U22978 (N_22978,N_21741,N_22247);
or U22979 (N_22979,N_21620,N_22145);
xnor U22980 (N_22980,N_21533,N_21562);
and U22981 (N_22981,N_21421,N_22122);
or U22982 (N_22982,N_21810,N_21390);
and U22983 (N_22983,N_21886,N_22113);
xnor U22984 (N_22984,N_22316,N_21797);
nor U22985 (N_22985,N_21726,N_21653);
nor U22986 (N_22986,N_22444,N_21308);
xor U22987 (N_22987,N_22048,N_21729);
xor U22988 (N_22988,N_21399,N_21538);
or U22989 (N_22989,N_21285,N_21316);
xor U22990 (N_22990,N_22169,N_22285);
xnor U22991 (N_22991,N_21737,N_22384);
xor U22992 (N_22992,N_21800,N_21630);
xnor U22993 (N_22993,N_21352,N_21486);
nor U22994 (N_22994,N_21581,N_21982);
nand U22995 (N_22995,N_21883,N_22038);
or U22996 (N_22996,N_22203,N_22383);
xnor U22997 (N_22997,N_22232,N_21522);
and U22998 (N_22998,N_21541,N_21903);
or U22999 (N_22999,N_22098,N_22341);
or U23000 (N_23000,N_22042,N_21323);
or U23001 (N_23001,N_22342,N_21492);
nand U23002 (N_23002,N_22283,N_21305);
and U23003 (N_23003,N_21379,N_21476);
xor U23004 (N_23004,N_22346,N_21565);
xor U23005 (N_23005,N_21940,N_21327);
nor U23006 (N_23006,N_22275,N_21958);
and U23007 (N_23007,N_21756,N_22297);
nand U23008 (N_23008,N_22499,N_22339);
or U23009 (N_23009,N_21798,N_22217);
and U23010 (N_23010,N_22407,N_21258);
xnor U23011 (N_23011,N_21921,N_21561);
xnor U23012 (N_23012,N_22154,N_21397);
nand U23013 (N_23013,N_22377,N_21956);
nand U23014 (N_23014,N_22441,N_21871);
nor U23015 (N_23015,N_21981,N_22314);
xor U23016 (N_23016,N_21639,N_21510);
nor U23017 (N_23017,N_21765,N_22166);
or U23018 (N_23018,N_22110,N_21744);
and U23019 (N_23019,N_22301,N_21708);
nor U23020 (N_23020,N_21600,N_21303);
or U23021 (N_23021,N_21939,N_21678);
and U23022 (N_23022,N_22139,N_21619);
nor U23023 (N_23023,N_22311,N_21404);
nand U23024 (N_23024,N_21529,N_22028);
nor U23025 (N_23025,N_22001,N_22040);
and U23026 (N_23026,N_21402,N_22351);
nor U23027 (N_23027,N_21434,N_22151);
and U23028 (N_23028,N_22350,N_21580);
xnor U23029 (N_23029,N_21748,N_22213);
or U23030 (N_23030,N_21980,N_22278);
nor U23031 (N_23031,N_21962,N_22249);
nand U23032 (N_23032,N_21846,N_21936);
nand U23033 (N_23033,N_22052,N_22293);
nand U23034 (N_23034,N_22357,N_21294);
xnor U23035 (N_23035,N_21724,N_22220);
nor U23036 (N_23036,N_22172,N_22012);
nand U23037 (N_23037,N_21607,N_21412);
xnor U23038 (N_23038,N_21312,N_21518);
or U23039 (N_23039,N_22117,N_21497);
and U23040 (N_23040,N_21408,N_21861);
and U23041 (N_23041,N_21481,N_21689);
nor U23042 (N_23042,N_21637,N_21673);
or U23043 (N_23043,N_21566,N_22424);
nor U23044 (N_23044,N_21686,N_21367);
nor U23045 (N_23045,N_22101,N_22289);
nor U23046 (N_23046,N_21416,N_22387);
nand U23047 (N_23047,N_21927,N_22392);
xor U23048 (N_23048,N_22094,N_21463);
xnor U23049 (N_23049,N_21493,N_22319);
or U23050 (N_23050,N_21818,N_21879);
and U23051 (N_23051,N_21925,N_22016);
nand U23052 (N_23052,N_21930,N_21728);
nor U23053 (N_23053,N_21839,N_21583);
nand U23054 (N_23054,N_21959,N_21788);
or U23055 (N_23055,N_22190,N_21475);
nor U23056 (N_23056,N_21292,N_22358);
and U23057 (N_23057,N_21749,N_22310);
and U23058 (N_23058,N_21647,N_21545);
and U23059 (N_23059,N_22340,N_21288);
or U23060 (N_23060,N_21551,N_21372);
nor U23061 (N_23061,N_21764,N_21875);
or U23062 (N_23062,N_22180,N_21317);
nor U23063 (N_23063,N_22023,N_22402);
nand U23064 (N_23064,N_21852,N_22277);
nand U23065 (N_23065,N_22198,N_22119);
nand U23066 (N_23066,N_21385,N_21295);
nor U23067 (N_23067,N_22386,N_22226);
and U23068 (N_23068,N_21677,N_21325);
xor U23069 (N_23069,N_22084,N_21509);
or U23070 (N_23070,N_21516,N_21597);
nand U23071 (N_23071,N_21532,N_22410);
xnor U23072 (N_23072,N_22414,N_21572);
or U23073 (N_23073,N_21315,N_21854);
nor U23074 (N_23074,N_21751,N_21783);
nor U23075 (N_23075,N_22199,N_21802);
nor U23076 (N_23076,N_22107,N_22498);
xnor U23077 (N_23077,N_21626,N_21467);
and U23078 (N_23078,N_21926,N_21556);
and U23079 (N_23079,N_22372,N_21451);
xor U23080 (N_23080,N_21912,N_21696);
xor U23081 (N_23081,N_21752,N_22011);
and U23082 (N_23082,N_21640,N_21490);
and U23083 (N_23083,N_21584,N_21720);
xnor U23084 (N_23084,N_22290,N_22333);
or U23085 (N_23085,N_21814,N_22334);
nand U23086 (N_23086,N_22472,N_21498);
and U23087 (N_23087,N_22080,N_21550);
xor U23088 (N_23088,N_22485,N_21624);
nand U23089 (N_23089,N_21523,N_22242);
xor U23090 (N_23090,N_22435,N_21766);
and U23091 (N_23091,N_21376,N_22409);
and U23092 (N_23092,N_22446,N_22462);
nand U23093 (N_23093,N_21806,N_21917);
nor U23094 (N_23094,N_22476,N_22360);
or U23095 (N_23095,N_22332,N_22044);
nand U23096 (N_23096,N_21530,N_22013);
nor U23097 (N_23097,N_21460,N_22227);
xnor U23098 (N_23098,N_21628,N_21307);
or U23099 (N_23099,N_21517,N_21549);
nand U23100 (N_23100,N_21585,N_21355);
or U23101 (N_23101,N_21988,N_22083);
nor U23102 (N_23102,N_22126,N_21711);
nor U23103 (N_23103,N_21851,N_21423);
xor U23104 (N_23104,N_22321,N_21933);
or U23105 (N_23105,N_21671,N_22133);
nand U23106 (N_23106,N_22378,N_21651);
or U23107 (N_23107,N_21976,N_22097);
and U23108 (N_23108,N_21349,N_22235);
or U23109 (N_23109,N_21793,N_21318);
nor U23110 (N_23110,N_21837,N_22493);
nor U23111 (N_23111,N_22102,N_21816);
nor U23112 (N_23112,N_21702,N_22241);
xnor U23113 (N_23113,N_21575,N_21511);
or U23114 (N_23114,N_21857,N_21364);
or U23115 (N_23115,N_22421,N_21306);
and U23116 (N_23116,N_21971,N_21908);
xnor U23117 (N_23117,N_22147,N_22109);
nand U23118 (N_23118,N_22170,N_21262);
nor U23119 (N_23119,N_21642,N_22043);
and U23120 (N_23120,N_22163,N_21913);
nor U23121 (N_23121,N_22496,N_21540);
nand U23122 (N_23122,N_22142,N_22268);
xnor U23123 (N_23123,N_21838,N_21668);
or U23124 (N_23124,N_21287,N_22178);
or U23125 (N_23125,N_21744,N_22444);
xnor U23126 (N_23126,N_22247,N_21518);
and U23127 (N_23127,N_21268,N_22244);
nor U23128 (N_23128,N_21880,N_21561);
nand U23129 (N_23129,N_21700,N_21542);
xor U23130 (N_23130,N_21441,N_21998);
nand U23131 (N_23131,N_21491,N_21808);
and U23132 (N_23132,N_21667,N_21494);
nand U23133 (N_23133,N_21350,N_22425);
nor U23134 (N_23134,N_22109,N_21994);
and U23135 (N_23135,N_21527,N_21912);
nor U23136 (N_23136,N_22382,N_21382);
xnor U23137 (N_23137,N_21786,N_21986);
nor U23138 (N_23138,N_21911,N_21608);
xnor U23139 (N_23139,N_22132,N_21883);
nand U23140 (N_23140,N_22024,N_21300);
nand U23141 (N_23141,N_21656,N_22216);
nand U23142 (N_23142,N_21883,N_22032);
xnor U23143 (N_23143,N_22342,N_21490);
xor U23144 (N_23144,N_21456,N_21341);
nand U23145 (N_23145,N_22098,N_22362);
or U23146 (N_23146,N_21371,N_22342);
and U23147 (N_23147,N_21593,N_22301);
nand U23148 (N_23148,N_21469,N_22270);
xor U23149 (N_23149,N_22150,N_21663);
and U23150 (N_23150,N_22455,N_21885);
and U23151 (N_23151,N_21544,N_22154);
xnor U23152 (N_23152,N_21402,N_22037);
and U23153 (N_23153,N_22321,N_21265);
xor U23154 (N_23154,N_22243,N_21722);
nor U23155 (N_23155,N_21529,N_22262);
nor U23156 (N_23156,N_21633,N_22018);
or U23157 (N_23157,N_21870,N_22160);
or U23158 (N_23158,N_22303,N_21419);
or U23159 (N_23159,N_22041,N_21710);
nor U23160 (N_23160,N_21488,N_22063);
and U23161 (N_23161,N_21512,N_22360);
nor U23162 (N_23162,N_21582,N_22126);
nor U23163 (N_23163,N_22077,N_21872);
and U23164 (N_23164,N_21582,N_21436);
nor U23165 (N_23165,N_22045,N_21724);
nand U23166 (N_23166,N_22249,N_22107);
nor U23167 (N_23167,N_21965,N_21503);
and U23168 (N_23168,N_22386,N_21697);
nand U23169 (N_23169,N_21349,N_22042);
or U23170 (N_23170,N_21905,N_21583);
and U23171 (N_23171,N_21340,N_22421);
or U23172 (N_23172,N_22361,N_21769);
or U23173 (N_23173,N_22431,N_22038);
and U23174 (N_23174,N_21328,N_21934);
xor U23175 (N_23175,N_22083,N_21521);
and U23176 (N_23176,N_22425,N_22088);
xnor U23177 (N_23177,N_21352,N_21426);
nor U23178 (N_23178,N_22200,N_21992);
and U23179 (N_23179,N_21844,N_22079);
nor U23180 (N_23180,N_21799,N_22444);
nand U23181 (N_23181,N_21267,N_21488);
xor U23182 (N_23182,N_22329,N_21428);
and U23183 (N_23183,N_21755,N_22124);
xor U23184 (N_23184,N_22026,N_21315);
nand U23185 (N_23185,N_21945,N_22387);
xor U23186 (N_23186,N_21466,N_21708);
or U23187 (N_23187,N_21447,N_21435);
or U23188 (N_23188,N_21382,N_21960);
xor U23189 (N_23189,N_21357,N_21483);
xnor U23190 (N_23190,N_22152,N_21990);
or U23191 (N_23191,N_21895,N_21275);
nand U23192 (N_23192,N_21449,N_22023);
or U23193 (N_23193,N_21646,N_21281);
or U23194 (N_23194,N_21461,N_21651);
nand U23195 (N_23195,N_21484,N_21907);
or U23196 (N_23196,N_21629,N_22088);
or U23197 (N_23197,N_21731,N_21763);
and U23198 (N_23198,N_22121,N_22419);
nand U23199 (N_23199,N_22211,N_21628);
or U23200 (N_23200,N_21328,N_21272);
xnor U23201 (N_23201,N_22206,N_21386);
and U23202 (N_23202,N_22401,N_21372);
nor U23203 (N_23203,N_22284,N_22302);
and U23204 (N_23204,N_22465,N_22310);
nand U23205 (N_23205,N_21560,N_22033);
nor U23206 (N_23206,N_21789,N_21990);
or U23207 (N_23207,N_21329,N_22381);
and U23208 (N_23208,N_21915,N_22073);
nand U23209 (N_23209,N_21310,N_22115);
nor U23210 (N_23210,N_22004,N_21395);
and U23211 (N_23211,N_22183,N_22256);
and U23212 (N_23212,N_21503,N_21921);
nor U23213 (N_23213,N_21576,N_22215);
nand U23214 (N_23214,N_21363,N_22011);
and U23215 (N_23215,N_22079,N_22372);
or U23216 (N_23216,N_21780,N_21656);
xnor U23217 (N_23217,N_21802,N_21966);
xor U23218 (N_23218,N_21853,N_21574);
nand U23219 (N_23219,N_21665,N_22198);
or U23220 (N_23220,N_21594,N_22196);
xor U23221 (N_23221,N_21264,N_21286);
and U23222 (N_23222,N_22418,N_22029);
or U23223 (N_23223,N_22030,N_21906);
xnor U23224 (N_23224,N_22086,N_22215);
xor U23225 (N_23225,N_21922,N_21287);
nor U23226 (N_23226,N_21982,N_21393);
or U23227 (N_23227,N_22145,N_22253);
nor U23228 (N_23228,N_22193,N_21749);
nand U23229 (N_23229,N_22083,N_22446);
nor U23230 (N_23230,N_22296,N_21510);
nor U23231 (N_23231,N_22308,N_21814);
nor U23232 (N_23232,N_22231,N_21804);
and U23233 (N_23233,N_22231,N_21842);
and U23234 (N_23234,N_22405,N_21995);
nor U23235 (N_23235,N_21445,N_22216);
nor U23236 (N_23236,N_22427,N_22494);
xor U23237 (N_23237,N_22309,N_21939);
and U23238 (N_23238,N_21912,N_21701);
xor U23239 (N_23239,N_21608,N_21768);
nor U23240 (N_23240,N_21736,N_22222);
and U23241 (N_23241,N_22168,N_22289);
nand U23242 (N_23242,N_21917,N_21308);
nand U23243 (N_23243,N_21932,N_22475);
nor U23244 (N_23244,N_21717,N_21348);
nand U23245 (N_23245,N_21336,N_22091);
and U23246 (N_23246,N_22311,N_22328);
nor U23247 (N_23247,N_21872,N_21735);
or U23248 (N_23248,N_22004,N_21545);
or U23249 (N_23249,N_21910,N_21689);
nand U23250 (N_23250,N_21830,N_22175);
nand U23251 (N_23251,N_21436,N_21389);
or U23252 (N_23252,N_21610,N_21545);
nor U23253 (N_23253,N_21331,N_21314);
nand U23254 (N_23254,N_22298,N_22027);
and U23255 (N_23255,N_21463,N_21885);
nor U23256 (N_23256,N_22207,N_21787);
and U23257 (N_23257,N_21318,N_22016);
xor U23258 (N_23258,N_21649,N_21912);
nand U23259 (N_23259,N_21814,N_21509);
and U23260 (N_23260,N_21841,N_22046);
nand U23261 (N_23261,N_21986,N_21671);
or U23262 (N_23262,N_21655,N_22088);
xor U23263 (N_23263,N_21448,N_22343);
or U23264 (N_23264,N_21294,N_22120);
nor U23265 (N_23265,N_22223,N_21351);
or U23266 (N_23266,N_22406,N_21556);
xor U23267 (N_23267,N_22318,N_22435);
nand U23268 (N_23268,N_22099,N_22388);
nand U23269 (N_23269,N_21716,N_22015);
nand U23270 (N_23270,N_21477,N_22118);
or U23271 (N_23271,N_21340,N_21705);
or U23272 (N_23272,N_21552,N_21939);
or U23273 (N_23273,N_21332,N_22160);
and U23274 (N_23274,N_22388,N_21505);
or U23275 (N_23275,N_22358,N_21544);
nor U23276 (N_23276,N_21895,N_21586);
and U23277 (N_23277,N_22053,N_21338);
and U23278 (N_23278,N_21451,N_21705);
nand U23279 (N_23279,N_21376,N_22320);
nand U23280 (N_23280,N_21936,N_21333);
nor U23281 (N_23281,N_22379,N_22263);
or U23282 (N_23282,N_21689,N_21367);
and U23283 (N_23283,N_22248,N_21503);
nor U23284 (N_23284,N_21739,N_21948);
xor U23285 (N_23285,N_22271,N_21495);
nand U23286 (N_23286,N_22431,N_21922);
xnor U23287 (N_23287,N_21783,N_21477);
xor U23288 (N_23288,N_21926,N_21560);
or U23289 (N_23289,N_21511,N_21348);
and U23290 (N_23290,N_21374,N_21316);
nor U23291 (N_23291,N_21295,N_21300);
nor U23292 (N_23292,N_21889,N_22013);
xor U23293 (N_23293,N_21494,N_21295);
nor U23294 (N_23294,N_21612,N_22406);
xor U23295 (N_23295,N_22204,N_21561);
and U23296 (N_23296,N_21298,N_21951);
nand U23297 (N_23297,N_22203,N_21479);
and U23298 (N_23298,N_21488,N_22081);
nand U23299 (N_23299,N_21887,N_21600);
xnor U23300 (N_23300,N_22233,N_22226);
or U23301 (N_23301,N_22312,N_21306);
or U23302 (N_23302,N_21290,N_21616);
nor U23303 (N_23303,N_22333,N_21519);
xor U23304 (N_23304,N_21753,N_21470);
xnor U23305 (N_23305,N_22238,N_21986);
nand U23306 (N_23306,N_22011,N_21595);
nor U23307 (N_23307,N_22206,N_21960);
xor U23308 (N_23308,N_22434,N_21323);
nand U23309 (N_23309,N_21639,N_21273);
and U23310 (N_23310,N_21764,N_22370);
or U23311 (N_23311,N_22330,N_21852);
nor U23312 (N_23312,N_22153,N_21559);
and U23313 (N_23313,N_22444,N_21343);
xor U23314 (N_23314,N_21284,N_22185);
nor U23315 (N_23315,N_22325,N_22494);
and U23316 (N_23316,N_22417,N_22431);
or U23317 (N_23317,N_22351,N_22312);
xor U23318 (N_23318,N_21494,N_22012);
xor U23319 (N_23319,N_21382,N_21626);
nor U23320 (N_23320,N_22192,N_22121);
nand U23321 (N_23321,N_22431,N_21381);
xor U23322 (N_23322,N_21966,N_21948);
nor U23323 (N_23323,N_22121,N_21443);
and U23324 (N_23324,N_21287,N_22029);
and U23325 (N_23325,N_21942,N_21822);
xor U23326 (N_23326,N_21515,N_22262);
and U23327 (N_23327,N_22286,N_22136);
and U23328 (N_23328,N_22006,N_22485);
nor U23329 (N_23329,N_21455,N_21693);
nor U23330 (N_23330,N_22311,N_22275);
nand U23331 (N_23331,N_21767,N_21519);
nand U23332 (N_23332,N_21649,N_21722);
nor U23333 (N_23333,N_21291,N_22115);
nand U23334 (N_23334,N_22058,N_21810);
nand U23335 (N_23335,N_21263,N_22097);
or U23336 (N_23336,N_21404,N_22471);
and U23337 (N_23337,N_21734,N_21675);
nor U23338 (N_23338,N_21335,N_21741);
nand U23339 (N_23339,N_21873,N_21341);
nand U23340 (N_23340,N_22132,N_21509);
xnor U23341 (N_23341,N_21390,N_21424);
nor U23342 (N_23342,N_22081,N_22498);
nand U23343 (N_23343,N_22341,N_21511);
xor U23344 (N_23344,N_22178,N_22465);
nand U23345 (N_23345,N_22332,N_22392);
or U23346 (N_23346,N_21558,N_21928);
xor U23347 (N_23347,N_21748,N_21591);
xnor U23348 (N_23348,N_22431,N_21652);
nor U23349 (N_23349,N_21874,N_22305);
or U23350 (N_23350,N_22337,N_21429);
nand U23351 (N_23351,N_22382,N_22030);
nand U23352 (N_23352,N_21768,N_21459);
nor U23353 (N_23353,N_22094,N_22415);
or U23354 (N_23354,N_22023,N_21989);
and U23355 (N_23355,N_21338,N_21375);
xnor U23356 (N_23356,N_21988,N_21791);
xor U23357 (N_23357,N_22113,N_22035);
or U23358 (N_23358,N_21901,N_22414);
nor U23359 (N_23359,N_21313,N_22205);
and U23360 (N_23360,N_21303,N_21804);
and U23361 (N_23361,N_21628,N_21385);
or U23362 (N_23362,N_21628,N_22137);
or U23363 (N_23363,N_21614,N_21843);
or U23364 (N_23364,N_21767,N_21659);
xor U23365 (N_23365,N_21754,N_21655);
and U23366 (N_23366,N_22117,N_21334);
xnor U23367 (N_23367,N_22355,N_21686);
and U23368 (N_23368,N_21817,N_22055);
nand U23369 (N_23369,N_22406,N_22180);
xor U23370 (N_23370,N_21256,N_22328);
nand U23371 (N_23371,N_21740,N_21616);
and U23372 (N_23372,N_22338,N_21313);
nor U23373 (N_23373,N_22441,N_22017);
or U23374 (N_23374,N_21742,N_22432);
xor U23375 (N_23375,N_21374,N_22156);
nand U23376 (N_23376,N_21678,N_22187);
or U23377 (N_23377,N_21930,N_22467);
and U23378 (N_23378,N_21465,N_22072);
nor U23379 (N_23379,N_21469,N_22255);
and U23380 (N_23380,N_21713,N_21726);
xor U23381 (N_23381,N_21595,N_22025);
nor U23382 (N_23382,N_22200,N_21945);
and U23383 (N_23383,N_22032,N_22327);
xor U23384 (N_23384,N_21379,N_21607);
nand U23385 (N_23385,N_22370,N_21260);
xor U23386 (N_23386,N_22438,N_21562);
nor U23387 (N_23387,N_22034,N_21414);
and U23388 (N_23388,N_21861,N_22014);
nand U23389 (N_23389,N_22098,N_21466);
nor U23390 (N_23390,N_22187,N_22219);
nor U23391 (N_23391,N_22275,N_21976);
nor U23392 (N_23392,N_21445,N_21911);
nand U23393 (N_23393,N_21932,N_21421);
xor U23394 (N_23394,N_22177,N_22190);
nand U23395 (N_23395,N_21491,N_21311);
nand U23396 (N_23396,N_21459,N_21253);
nand U23397 (N_23397,N_21733,N_21847);
and U23398 (N_23398,N_21779,N_21267);
or U23399 (N_23399,N_21705,N_21950);
xor U23400 (N_23400,N_21791,N_22435);
or U23401 (N_23401,N_21736,N_21505);
and U23402 (N_23402,N_21653,N_21627);
nand U23403 (N_23403,N_21398,N_21743);
nand U23404 (N_23404,N_21957,N_22059);
and U23405 (N_23405,N_22359,N_21265);
nand U23406 (N_23406,N_21900,N_21500);
nand U23407 (N_23407,N_21535,N_22299);
nor U23408 (N_23408,N_21293,N_22195);
and U23409 (N_23409,N_21753,N_22460);
xnor U23410 (N_23410,N_22490,N_21973);
nand U23411 (N_23411,N_21572,N_21907);
and U23412 (N_23412,N_22332,N_21453);
xor U23413 (N_23413,N_21340,N_21550);
and U23414 (N_23414,N_21641,N_22435);
and U23415 (N_23415,N_21741,N_21931);
or U23416 (N_23416,N_21539,N_21926);
nor U23417 (N_23417,N_21661,N_21787);
nor U23418 (N_23418,N_21853,N_21663);
xnor U23419 (N_23419,N_21711,N_22423);
nor U23420 (N_23420,N_21750,N_22180);
xor U23421 (N_23421,N_22464,N_22102);
or U23422 (N_23422,N_21909,N_21275);
nand U23423 (N_23423,N_21405,N_22278);
xnor U23424 (N_23424,N_22080,N_21478);
nor U23425 (N_23425,N_22078,N_21715);
or U23426 (N_23426,N_22225,N_22399);
nor U23427 (N_23427,N_22270,N_22083);
nor U23428 (N_23428,N_21945,N_21397);
or U23429 (N_23429,N_22176,N_21780);
nand U23430 (N_23430,N_21498,N_21991);
xnor U23431 (N_23431,N_21330,N_21462);
and U23432 (N_23432,N_22145,N_22126);
xnor U23433 (N_23433,N_21656,N_22132);
nand U23434 (N_23434,N_21642,N_21727);
and U23435 (N_23435,N_22032,N_21604);
nand U23436 (N_23436,N_22443,N_22159);
xor U23437 (N_23437,N_21626,N_21929);
nand U23438 (N_23438,N_22042,N_22264);
or U23439 (N_23439,N_22259,N_22037);
and U23440 (N_23440,N_21648,N_22328);
nor U23441 (N_23441,N_22129,N_22072);
nor U23442 (N_23442,N_21956,N_21362);
nor U23443 (N_23443,N_21657,N_22481);
or U23444 (N_23444,N_21372,N_22298);
nand U23445 (N_23445,N_21727,N_21865);
xnor U23446 (N_23446,N_21547,N_21765);
or U23447 (N_23447,N_21491,N_21976);
and U23448 (N_23448,N_21874,N_21976);
and U23449 (N_23449,N_22272,N_22150);
nand U23450 (N_23450,N_21763,N_21714);
and U23451 (N_23451,N_21376,N_22122);
nand U23452 (N_23452,N_21833,N_21921);
or U23453 (N_23453,N_21573,N_22161);
or U23454 (N_23454,N_22213,N_21329);
xor U23455 (N_23455,N_21551,N_22452);
nand U23456 (N_23456,N_21581,N_22370);
and U23457 (N_23457,N_21363,N_21830);
xnor U23458 (N_23458,N_21731,N_21592);
xnor U23459 (N_23459,N_21421,N_21928);
or U23460 (N_23460,N_22419,N_21512);
or U23461 (N_23461,N_21659,N_22069);
nor U23462 (N_23462,N_21946,N_21425);
nor U23463 (N_23463,N_22142,N_21864);
or U23464 (N_23464,N_22262,N_21702);
nand U23465 (N_23465,N_22183,N_22491);
nand U23466 (N_23466,N_21780,N_21506);
nand U23467 (N_23467,N_21570,N_21349);
nor U23468 (N_23468,N_22398,N_21819);
nor U23469 (N_23469,N_21379,N_21295);
nand U23470 (N_23470,N_21762,N_21637);
or U23471 (N_23471,N_22105,N_22282);
and U23472 (N_23472,N_21357,N_21577);
xor U23473 (N_23473,N_21519,N_21729);
and U23474 (N_23474,N_21579,N_21676);
and U23475 (N_23475,N_21277,N_21416);
and U23476 (N_23476,N_22122,N_22488);
xnor U23477 (N_23477,N_21466,N_21651);
or U23478 (N_23478,N_21939,N_22341);
nor U23479 (N_23479,N_21991,N_22409);
and U23480 (N_23480,N_21294,N_21934);
nand U23481 (N_23481,N_21913,N_21355);
xor U23482 (N_23482,N_22249,N_21976);
or U23483 (N_23483,N_21285,N_21576);
nor U23484 (N_23484,N_22305,N_21494);
or U23485 (N_23485,N_22233,N_21440);
nor U23486 (N_23486,N_21445,N_22317);
xor U23487 (N_23487,N_21905,N_21720);
xor U23488 (N_23488,N_22479,N_22164);
nand U23489 (N_23489,N_22366,N_22145);
xnor U23490 (N_23490,N_21766,N_21797);
nor U23491 (N_23491,N_22338,N_21864);
xor U23492 (N_23492,N_21707,N_21445);
and U23493 (N_23493,N_22124,N_21378);
and U23494 (N_23494,N_21934,N_22252);
nand U23495 (N_23495,N_21713,N_21822);
xnor U23496 (N_23496,N_21944,N_21857);
nand U23497 (N_23497,N_21596,N_21640);
nor U23498 (N_23498,N_21890,N_22158);
or U23499 (N_23499,N_21792,N_21870);
and U23500 (N_23500,N_21444,N_21652);
or U23501 (N_23501,N_21879,N_21712);
xnor U23502 (N_23502,N_21485,N_21609);
nor U23503 (N_23503,N_21558,N_21875);
xnor U23504 (N_23504,N_22191,N_22348);
nor U23505 (N_23505,N_21790,N_22456);
xor U23506 (N_23506,N_21330,N_21899);
and U23507 (N_23507,N_21471,N_21987);
nor U23508 (N_23508,N_21914,N_21443);
or U23509 (N_23509,N_21608,N_21953);
nand U23510 (N_23510,N_22494,N_21693);
nor U23511 (N_23511,N_21381,N_22216);
or U23512 (N_23512,N_21707,N_21415);
nand U23513 (N_23513,N_22445,N_21541);
nand U23514 (N_23514,N_22117,N_21670);
xor U23515 (N_23515,N_22340,N_21706);
or U23516 (N_23516,N_22087,N_21672);
nand U23517 (N_23517,N_21860,N_21985);
or U23518 (N_23518,N_22026,N_21954);
or U23519 (N_23519,N_21853,N_21313);
nor U23520 (N_23520,N_21295,N_22176);
or U23521 (N_23521,N_21863,N_21384);
or U23522 (N_23522,N_21706,N_21329);
nor U23523 (N_23523,N_21364,N_22276);
nand U23524 (N_23524,N_21767,N_21704);
and U23525 (N_23525,N_21682,N_21987);
nand U23526 (N_23526,N_21654,N_21819);
and U23527 (N_23527,N_22171,N_21659);
or U23528 (N_23528,N_21861,N_22483);
and U23529 (N_23529,N_21930,N_21568);
or U23530 (N_23530,N_22169,N_21872);
or U23531 (N_23531,N_21253,N_22180);
or U23532 (N_23532,N_21538,N_21947);
and U23533 (N_23533,N_21839,N_21735);
or U23534 (N_23534,N_21502,N_22043);
or U23535 (N_23535,N_22254,N_21964);
and U23536 (N_23536,N_22027,N_22127);
or U23537 (N_23537,N_21670,N_21982);
nor U23538 (N_23538,N_21506,N_22480);
and U23539 (N_23539,N_22220,N_22408);
nor U23540 (N_23540,N_21863,N_22480);
and U23541 (N_23541,N_21507,N_21463);
nand U23542 (N_23542,N_21783,N_22116);
xnor U23543 (N_23543,N_22016,N_22203);
nand U23544 (N_23544,N_22143,N_22053);
or U23545 (N_23545,N_21368,N_21257);
xnor U23546 (N_23546,N_22443,N_21776);
xor U23547 (N_23547,N_21423,N_22018);
or U23548 (N_23548,N_22133,N_21337);
or U23549 (N_23549,N_21821,N_21574);
nand U23550 (N_23550,N_22147,N_22377);
nor U23551 (N_23551,N_21517,N_21435);
xor U23552 (N_23552,N_21664,N_21914);
nor U23553 (N_23553,N_22166,N_21449);
nand U23554 (N_23554,N_22351,N_21258);
and U23555 (N_23555,N_21642,N_21357);
xnor U23556 (N_23556,N_21333,N_21971);
or U23557 (N_23557,N_22019,N_22097);
or U23558 (N_23558,N_22350,N_22068);
nand U23559 (N_23559,N_21766,N_22423);
or U23560 (N_23560,N_21447,N_21535);
xor U23561 (N_23561,N_22172,N_21771);
and U23562 (N_23562,N_21340,N_22237);
nor U23563 (N_23563,N_21447,N_21625);
xor U23564 (N_23564,N_21714,N_21266);
or U23565 (N_23565,N_21633,N_21275);
nor U23566 (N_23566,N_22288,N_21853);
nor U23567 (N_23567,N_21437,N_22122);
or U23568 (N_23568,N_22363,N_22095);
xnor U23569 (N_23569,N_21689,N_21765);
nand U23570 (N_23570,N_21978,N_22459);
or U23571 (N_23571,N_22168,N_22325);
and U23572 (N_23572,N_21467,N_22296);
or U23573 (N_23573,N_21990,N_21790);
nor U23574 (N_23574,N_21376,N_22131);
xor U23575 (N_23575,N_21447,N_21831);
nand U23576 (N_23576,N_21852,N_22171);
nand U23577 (N_23577,N_22255,N_21552);
and U23578 (N_23578,N_22402,N_22417);
or U23579 (N_23579,N_21579,N_22481);
or U23580 (N_23580,N_21867,N_21445);
or U23581 (N_23581,N_21648,N_21924);
and U23582 (N_23582,N_21349,N_21541);
xnor U23583 (N_23583,N_21977,N_21432);
or U23584 (N_23584,N_21282,N_22235);
or U23585 (N_23585,N_21485,N_21303);
or U23586 (N_23586,N_21561,N_22470);
nor U23587 (N_23587,N_22331,N_22456);
xor U23588 (N_23588,N_21524,N_21629);
or U23589 (N_23589,N_21827,N_22422);
xnor U23590 (N_23590,N_21617,N_21624);
nand U23591 (N_23591,N_22104,N_22444);
xor U23592 (N_23592,N_22134,N_22247);
xnor U23593 (N_23593,N_21635,N_21924);
or U23594 (N_23594,N_22313,N_21873);
nor U23595 (N_23595,N_22087,N_22165);
and U23596 (N_23596,N_21472,N_22324);
xor U23597 (N_23597,N_21914,N_21281);
and U23598 (N_23598,N_21416,N_21395);
or U23599 (N_23599,N_21639,N_21693);
xnor U23600 (N_23600,N_22490,N_21757);
or U23601 (N_23601,N_22198,N_21469);
nand U23602 (N_23602,N_22195,N_21264);
nor U23603 (N_23603,N_22432,N_21886);
nand U23604 (N_23604,N_22105,N_22063);
nand U23605 (N_23605,N_21320,N_22344);
nand U23606 (N_23606,N_21607,N_21826);
xor U23607 (N_23607,N_22388,N_22441);
xnor U23608 (N_23608,N_21265,N_22158);
and U23609 (N_23609,N_21328,N_22307);
and U23610 (N_23610,N_21454,N_21491);
or U23611 (N_23611,N_21814,N_21444);
and U23612 (N_23612,N_21928,N_22049);
and U23613 (N_23613,N_21911,N_21330);
xor U23614 (N_23614,N_21536,N_21871);
nand U23615 (N_23615,N_22453,N_22483);
nor U23616 (N_23616,N_22319,N_21923);
nand U23617 (N_23617,N_22314,N_21647);
nor U23618 (N_23618,N_21941,N_21602);
nand U23619 (N_23619,N_22433,N_21287);
xor U23620 (N_23620,N_21342,N_21956);
and U23621 (N_23621,N_22368,N_21730);
nor U23622 (N_23622,N_22053,N_21859);
nor U23623 (N_23623,N_21391,N_22076);
nor U23624 (N_23624,N_21628,N_22034);
nor U23625 (N_23625,N_21262,N_22337);
and U23626 (N_23626,N_21337,N_21746);
nand U23627 (N_23627,N_21341,N_22074);
and U23628 (N_23628,N_21820,N_22411);
or U23629 (N_23629,N_21527,N_22252);
nand U23630 (N_23630,N_21451,N_22155);
or U23631 (N_23631,N_22357,N_22042);
nand U23632 (N_23632,N_22399,N_21645);
or U23633 (N_23633,N_22024,N_21898);
xor U23634 (N_23634,N_22238,N_22013);
nor U23635 (N_23635,N_21586,N_22242);
or U23636 (N_23636,N_21439,N_21595);
nand U23637 (N_23637,N_22239,N_22128);
nand U23638 (N_23638,N_21407,N_21453);
and U23639 (N_23639,N_21651,N_21590);
nand U23640 (N_23640,N_22293,N_21946);
xor U23641 (N_23641,N_21918,N_21726);
or U23642 (N_23642,N_21729,N_21803);
nor U23643 (N_23643,N_21576,N_21518);
and U23644 (N_23644,N_21714,N_21459);
xnor U23645 (N_23645,N_21358,N_21841);
xor U23646 (N_23646,N_22033,N_21479);
nand U23647 (N_23647,N_22227,N_22486);
nor U23648 (N_23648,N_21390,N_21809);
and U23649 (N_23649,N_22428,N_21377);
xor U23650 (N_23650,N_21269,N_21811);
or U23651 (N_23651,N_21291,N_21312);
and U23652 (N_23652,N_22057,N_21340);
and U23653 (N_23653,N_21621,N_22013);
nor U23654 (N_23654,N_22198,N_22241);
or U23655 (N_23655,N_22204,N_21438);
or U23656 (N_23656,N_21714,N_21888);
and U23657 (N_23657,N_22005,N_21910);
nand U23658 (N_23658,N_21368,N_21876);
or U23659 (N_23659,N_21313,N_21268);
and U23660 (N_23660,N_21451,N_21368);
nand U23661 (N_23661,N_22238,N_21425);
and U23662 (N_23662,N_21773,N_21429);
and U23663 (N_23663,N_22351,N_21452);
and U23664 (N_23664,N_21628,N_22485);
or U23665 (N_23665,N_21908,N_22116);
and U23666 (N_23666,N_21788,N_21557);
and U23667 (N_23667,N_22335,N_22361);
nand U23668 (N_23668,N_21309,N_22030);
nand U23669 (N_23669,N_21916,N_21880);
or U23670 (N_23670,N_22381,N_22311);
and U23671 (N_23671,N_22462,N_22448);
and U23672 (N_23672,N_21638,N_21811);
nor U23673 (N_23673,N_21807,N_21798);
nand U23674 (N_23674,N_21628,N_22147);
xor U23675 (N_23675,N_21565,N_21547);
xor U23676 (N_23676,N_22317,N_21948);
nand U23677 (N_23677,N_22358,N_21907);
xnor U23678 (N_23678,N_21266,N_21671);
or U23679 (N_23679,N_21358,N_22444);
and U23680 (N_23680,N_21881,N_21509);
nor U23681 (N_23681,N_21561,N_22017);
or U23682 (N_23682,N_22320,N_21432);
or U23683 (N_23683,N_21477,N_21277);
xor U23684 (N_23684,N_21366,N_21650);
nor U23685 (N_23685,N_22033,N_22445);
nand U23686 (N_23686,N_22268,N_21908);
or U23687 (N_23687,N_21878,N_22383);
and U23688 (N_23688,N_22489,N_22421);
nand U23689 (N_23689,N_22191,N_22313);
nor U23690 (N_23690,N_22126,N_21302);
or U23691 (N_23691,N_22146,N_22340);
nand U23692 (N_23692,N_22175,N_22306);
nand U23693 (N_23693,N_21859,N_22490);
and U23694 (N_23694,N_21411,N_21516);
and U23695 (N_23695,N_22435,N_21658);
or U23696 (N_23696,N_21522,N_21342);
and U23697 (N_23697,N_22440,N_21869);
nand U23698 (N_23698,N_21589,N_21524);
nor U23699 (N_23699,N_22196,N_21750);
or U23700 (N_23700,N_21660,N_21570);
and U23701 (N_23701,N_22335,N_22285);
or U23702 (N_23702,N_21396,N_22426);
nor U23703 (N_23703,N_21587,N_22026);
nor U23704 (N_23704,N_22337,N_21741);
nor U23705 (N_23705,N_21960,N_21488);
nand U23706 (N_23706,N_22238,N_21488);
nor U23707 (N_23707,N_21256,N_22104);
or U23708 (N_23708,N_21935,N_21503);
nand U23709 (N_23709,N_21748,N_22059);
xnor U23710 (N_23710,N_22238,N_21542);
xnor U23711 (N_23711,N_22267,N_21470);
nand U23712 (N_23712,N_22277,N_22364);
nor U23713 (N_23713,N_22039,N_21737);
xor U23714 (N_23714,N_21779,N_21708);
and U23715 (N_23715,N_21272,N_21363);
or U23716 (N_23716,N_21853,N_22276);
xnor U23717 (N_23717,N_21782,N_22091);
or U23718 (N_23718,N_21262,N_21833);
and U23719 (N_23719,N_22048,N_21718);
nand U23720 (N_23720,N_21531,N_21620);
xnor U23721 (N_23721,N_22315,N_21598);
nand U23722 (N_23722,N_22477,N_22121);
and U23723 (N_23723,N_22468,N_21367);
nor U23724 (N_23724,N_22312,N_22348);
or U23725 (N_23725,N_21685,N_21812);
or U23726 (N_23726,N_21421,N_21666);
nor U23727 (N_23727,N_22110,N_22392);
nor U23728 (N_23728,N_21491,N_21299);
nand U23729 (N_23729,N_21784,N_22241);
nor U23730 (N_23730,N_22249,N_22325);
nand U23731 (N_23731,N_21479,N_22229);
or U23732 (N_23732,N_22454,N_21438);
or U23733 (N_23733,N_21870,N_22275);
and U23734 (N_23734,N_21471,N_21614);
nor U23735 (N_23735,N_22112,N_21582);
and U23736 (N_23736,N_22121,N_21832);
or U23737 (N_23737,N_22219,N_21414);
nor U23738 (N_23738,N_21530,N_22423);
or U23739 (N_23739,N_21296,N_21573);
nand U23740 (N_23740,N_21254,N_22402);
nor U23741 (N_23741,N_22259,N_21602);
and U23742 (N_23742,N_21884,N_21680);
and U23743 (N_23743,N_21521,N_21613);
nand U23744 (N_23744,N_21977,N_21743);
or U23745 (N_23745,N_22008,N_21534);
xnor U23746 (N_23746,N_21919,N_22254);
and U23747 (N_23747,N_21715,N_22144);
nor U23748 (N_23748,N_21925,N_21864);
nor U23749 (N_23749,N_22093,N_21489);
and U23750 (N_23750,N_22928,N_22952);
or U23751 (N_23751,N_23221,N_22690);
nor U23752 (N_23752,N_22877,N_22678);
nand U23753 (N_23753,N_22541,N_22940);
xor U23754 (N_23754,N_23631,N_22552);
nor U23755 (N_23755,N_22626,N_22797);
and U23756 (N_23756,N_22676,N_23580);
and U23757 (N_23757,N_23538,N_23430);
and U23758 (N_23758,N_23032,N_22549);
or U23759 (N_23759,N_23099,N_22779);
xnor U23760 (N_23760,N_23306,N_23127);
nor U23761 (N_23761,N_22686,N_23448);
or U23762 (N_23762,N_23096,N_23201);
and U23763 (N_23763,N_23482,N_22646);
or U23764 (N_23764,N_23675,N_23647);
nor U23765 (N_23765,N_22879,N_22926);
nor U23766 (N_23766,N_22974,N_22675);
xnor U23767 (N_23767,N_22592,N_23077);
nor U23768 (N_23768,N_22531,N_23266);
and U23769 (N_23769,N_23704,N_22898);
and U23770 (N_23770,N_23052,N_23334);
nand U23771 (N_23771,N_23125,N_22593);
nor U23772 (N_23772,N_22874,N_22743);
xor U23773 (N_23773,N_23340,N_22757);
nor U23774 (N_23774,N_23173,N_23595);
xor U23775 (N_23775,N_23472,N_22643);
xor U23776 (N_23776,N_22808,N_22510);
xnor U23777 (N_23777,N_23263,N_23058);
nor U23778 (N_23778,N_22941,N_23092);
nand U23779 (N_23779,N_22931,N_22939);
or U23780 (N_23780,N_23449,N_22783);
nor U23781 (N_23781,N_22614,N_23514);
nand U23782 (N_23782,N_22768,N_23024);
nand U23783 (N_23783,N_23153,N_22681);
and U23784 (N_23784,N_23682,N_22766);
nor U23785 (N_23785,N_22540,N_22884);
or U23786 (N_23786,N_23387,N_23367);
nor U23787 (N_23787,N_22912,N_23332);
or U23788 (N_23788,N_22845,N_23039);
or U23789 (N_23789,N_22883,N_22658);
nand U23790 (N_23790,N_22753,N_23346);
xnor U23791 (N_23791,N_22633,N_22617);
nor U23792 (N_23792,N_23229,N_23107);
xor U23793 (N_23793,N_22839,N_22594);
nor U23794 (N_23794,N_23445,N_22764);
nand U23795 (N_23795,N_23660,N_23484);
nand U23796 (N_23796,N_22615,N_23276);
and U23797 (N_23797,N_23667,N_22554);
and U23798 (N_23798,N_22992,N_23275);
nand U23799 (N_23799,N_23343,N_23509);
or U23800 (N_23800,N_23703,N_23572);
or U23801 (N_23801,N_22842,N_23313);
xnor U23802 (N_23802,N_22989,N_22721);
or U23803 (N_23803,N_23042,N_23676);
nand U23804 (N_23804,N_23217,N_23004);
and U23805 (N_23805,N_22848,N_23303);
nor U23806 (N_23806,N_23150,N_22508);
xor U23807 (N_23807,N_22630,N_23728);
nand U23808 (N_23808,N_23624,N_23573);
nand U23809 (N_23809,N_22968,N_23167);
xnor U23810 (N_23810,N_23139,N_22668);
and U23811 (N_23811,N_23486,N_22698);
or U23812 (N_23812,N_22837,N_23634);
or U23813 (N_23813,N_23112,N_23249);
xor U23814 (N_23814,N_23239,N_23274);
or U23815 (N_23815,N_23318,N_23286);
xnor U23816 (N_23816,N_23529,N_22702);
and U23817 (N_23817,N_23132,N_23267);
or U23818 (N_23818,N_22920,N_22502);
nand U23819 (N_23819,N_22609,N_23129);
nor U23820 (N_23820,N_22752,N_23191);
nor U23821 (N_23821,N_22907,N_23015);
and U23822 (N_23822,N_23498,N_23088);
nor U23823 (N_23823,N_23557,N_23105);
xnor U23824 (N_23824,N_23335,N_22910);
or U23825 (N_23825,N_22555,N_23065);
nand U23826 (N_23826,N_23307,N_22534);
xor U23827 (N_23827,N_23135,N_23045);
xnor U23828 (N_23828,N_23713,N_23431);
xnor U23829 (N_23829,N_22737,N_23358);
or U23830 (N_23830,N_23568,N_23464);
xnor U23831 (N_23831,N_23567,N_23465);
and U23832 (N_23832,N_22880,N_22684);
xor U23833 (N_23833,N_23301,N_23578);
or U23834 (N_23834,N_23607,N_23501);
xnor U23835 (N_23835,N_23694,N_22695);
xor U23836 (N_23836,N_22760,N_23064);
nor U23837 (N_23837,N_23271,N_23025);
and U23838 (N_23838,N_22544,N_23216);
nand U23839 (N_23839,N_22929,N_23087);
or U23840 (N_23840,N_23493,N_22785);
or U23841 (N_23841,N_22951,N_22769);
and U23842 (N_23842,N_23026,N_23622);
nor U23843 (N_23843,N_23468,N_23606);
and U23844 (N_23844,N_22551,N_22997);
nand U23845 (N_23845,N_23337,N_22784);
nor U23846 (N_23846,N_22889,N_23666);
nor U23847 (N_23847,N_23451,N_23355);
or U23848 (N_23848,N_23463,N_23238);
or U23849 (N_23849,N_23097,N_22921);
nor U23850 (N_23850,N_22978,N_22663);
nand U23851 (N_23851,N_22582,N_22810);
or U23852 (N_23852,N_23053,N_22836);
xnor U23853 (N_23853,N_23657,N_22607);
nand U23854 (N_23854,N_23527,N_23550);
nand U23855 (N_23855,N_23178,N_23446);
or U23856 (N_23856,N_23198,N_22805);
and U23857 (N_23857,N_22747,N_22616);
and U23858 (N_23858,N_23688,N_22868);
and U23859 (N_23859,N_23021,N_22944);
nor U23860 (N_23860,N_23645,N_22699);
xnor U23861 (N_23861,N_22774,N_23426);
nand U23862 (N_23862,N_23709,N_23535);
nand U23863 (N_23863,N_22542,N_22801);
xor U23864 (N_23864,N_23215,N_23040);
and U23865 (N_23865,N_22644,N_22982);
nor U23866 (N_23866,N_23587,N_23461);
and U23867 (N_23867,N_23084,N_22969);
and U23868 (N_23868,N_22556,N_23192);
nand U23869 (N_23869,N_22826,N_23735);
or U23870 (N_23870,N_23590,N_23636);
and U23871 (N_23871,N_23700,N_22703);
nor U23872 (N_23872,N_22525,N_23711);
or U23873 (N_23873,N_22621,N_23503);
nand U23874 (N_23874,N_22949,N_23067);
nand U23875 (N_23875,N_23487,N_23723);
or U23876 (N_23876,N_22905,N_22962);
nor U23877 (N_23877,N_23166,N_23511);
nand U23878 (N_23878,N_22807,N_23546);
nand U23879 (N_23879,N_23554,N_22577);
xnor U23880 (N_23880,N_23491,N_23328);
xor U23881 (N_23881,N_23653,N_23627);
or U23882 (N_23882,N_22843,N_22528);
or U23883 (N_23883,N_22741,N_22563);
xnor U23884 (N_23884,N_22831,N_22682);
or U23885 (N_23885,N_22565,N_22995);
or U23886 (N_23886,N_23725,N_22948);
nor U23887 (N_23887,N_23197,N_23291);
or U23888 (N_23888,N_23278,N_23476);
or U23889 (N_23889,N_23670,N_23179);
and U23890 (N_23890,N_22538,N_23686);
nor U23891 (N_23891,N_22707,N_23441);
and U23892 (N_23892,N_22840,N_22543);
or U23893 (N_23893,N_22787,N_23050);
xor U23894 (N_23894,N_22767,N_22763);
nand U23895 (N_23895,N_23394,N_22586);
xnor U23896 (N_23896,N_23012,N_23341);
nand U23897 (N_23897,N_23734,N_22590);
nand U23898 (N_23898,N_23231,N_22895);
xor U23899 (N_23899,N_23499,N_23663);
nor U23900 (N_23900,N_23327,N_23220);
xnor U23901 (N_23901,N_22574,N_22622);
nand U23902 (N_23902,N_22624,N_23038);
nand U23903 (N_23903,N_22853,N_23471);
and U23904 (N_23904,N_22581,N_23162);
nand U23905 (N_23905,N_22778,N_23111);
or U23906 (N_23906,N_23420,N_22829);
nor U23907 (N_23907,N_22572,N_22657);
nor U23908 (N_23908,N_22712,N_22794);
and U23909 (N_23909,N_23749,N_22745);
and U23910 (N_23910,N_23022,N_22570);
nand U23911 (N_23911,N_22720,N_23424);
and U23912 (N_23912,N_23692,N_23621);
xnor U23913 (N_23913,N_23458,N_23268);
xor U23914 (N_23914,N_22838,N_22793);
nor U23915 (N_23915,N_23017,N_23669);
xnor U23916 (N_23916,N_23413,N_23410);
xor U23917 (N_23917,N_23226,N_22685);
xnor U23918 (N_23918,N_22786,N_22571);
nand U23919 (N_23919,N_23134,N_22927);
and U23920 (N_23920,N_22820,N_23262);
nand U23921 (N_23921,N_23223,N_22738);
nor U23922 (N_23922,N_23157,N_22611);
nand U23923 (N_23923,N_23322,N_23364);
xor U23924 (N_23924,N_23722,N_23679);
xor U23925 (N_23925,N_23143,N_23611);
or U23926 (N_23926,N_23057,N_23746);
xor U23927 (N_23927,N_22819,N_23289);
nand U23928 (N_23928,N_23001,N_22864);
xor U23929 (N_23929,N_22813,N_22535);
nand U23930 (N_23930,N_22674,N_22985);
nor U23931 (N_23931,N_22956,N_23365);
xnor U23932 (N_23932,N_23361,N_23395);
xnor U23933 (N_23933,N_23247,N_23385);
xnor U23934 (N_23934,N_22524,N_23730);
and U23935 (N_23935,N_23641,N_23377);
nand U23936 (N_23936,N_23460,N_23436);
nand U23937 (N_23937,N_22850,N_23649);
and U23938 (N_23938,N_23727,N_23495);
nand U23939 (N_23939,N_23138,N_22990);
nor U23940 (N_23940,N_23048,N_22830);
xor U23941 (N_23941,N_23095,N_23044);
nand U23942 (N_23942,N_23011,N_23222);
and U23943 (N_23943,N_23121,N_22645);
and U23944 (N_23944,N_23380,N_22585);
and U23945 (N_23945,N_23626,N_22601);
or U23946 (N_23946,N_22847,N_23594);
or U23947 (N_23947,N_22629,N_23715);
or U23948 (N_23948,N_22970,N_22824);
xnor U23949 (N_23949,N_23251,N_23685);
or U23950 (N_23950,N_22650,N_23681);
nand U23951 (N_23951,N_23654,N_22608);
nand U23952 (N_23952,N_23672,N_22517);
nor U23953 (N_23953,N_23388,N_23156);
and U23954 (N_23954,N_22655,N_22934);
nand U23955 (N_23955,N_23103,N_22724);
xor U23956 (N_23956,N_23299,N_22567);
or U23957 (N_23957,N_22892,N_23599);
and U23958 (N_23958,N_23211,N_23731);
or U23959 (N_23959,N_23183,N_23601);
xnor U23960 (N_23960,N_22885,N_23331);
nand U23961 (N_23961,N_23591,N_23193);
xor U23962 (N_23962,N_23287,N_22727);
or U23963 (N_23963,N_23515,N_23579);
nand U23964 (N_23964,N_23349,N_23210);
or U23965 (N_23965,N_23282,N_23080);
or U23966 (N_23966,N_23063,N_23284);
xor U23967 (N_23967,N_23507,N_23309);
and U23968 (N_23968,N_22602,N_23598);
or U23969 (N_23969,N_23644,N_22876);
nand U23970 (N_23970,N_22893,N_22746);
and U23971 (N_23971,N_23613,N_23540);
nor U23972 (N_23972,N_22569,N_23733);
nand U23973 (N_23973,N_22965,N_23524);
nor U23974 (N_23974,N_23148,N_23541);
and U23975 (N_23975,N_22548,N_23158);
nand U23976 (N_23976,N_23230,N_23585);
nand U23977 (N_23977,N_22566,N_22613);
and U23978 (N_23978,N_23200,N_22780);
xor U23979 (N_23979,N_23706,N_23565);
nand U23980 (N_23980,N_23240,N_22664);
or U23981 (N_23981,N_23311,N_23429);
nand U23982 (N_23982,N_23124,N_23610);
nor U23983 (N_23983,N_23130,N_23202);
nor U23984 (N_23984,N_23623,N_23297);
xnor U23985 (N_23985,N_23574,N_23551);
or U23986 (N_23986,N_23504,N_22964);
xor U23987 (N_23987,N_22589,N_23374);
xor U23988 (N_23988,N_22976,N_23142);
and U23989 (N_23989,N_22692,N_23633);
nand U23990 (N_23990,N_23650,N_22800);
or U23991 (N_23991,N_23292,N_23227);
nor U23992 (N_23992,N_23533,N_22661);
xnor U23993 (N_23993,N_22762,N_22665);
xnor U23994 (N_23994,N_23416,N_23225);
xnor U23995 (N_23995,N_22537,N_23205);
or U23996 (N_23996,N_23566,N_23705);
nand U23997 (N_23997,N_22722,N_22963);
and U23998 (N_23998,N_23242,N_23505);
or U23999 (N_23999,N_23656,N_23444);
nor U24000 (N_24000,N_22873,N_23028);
xor U24001 (N_24001,N_23141,N_23639);
xor U24002 (N_24002,N_22715,N_23145);
and U24003 (N_24003,N_22993,N_23072);
xnor U24004 (N_24004,N_23712,N_22803);
and U24005 (N_24005,N_23203,N_22642);
or U24006 (N_24006,N_23433,N_23090);
nor U24007 (N_24007,N_22708,N_22687);
nor U24008 (N_24008,N_23018,N_23213);
xnor U24009 (N_24009,N_22798,N_22716);
and U24010 (N_24010,N_23720,N_22790);
nor U24011 (N_24011,N_23593,N_23483);
nand U24012 (N_24012,N_23002,N_22732);
or U24013 (N_24013,N_23272,N_23204);
and U24014 (N_24014,N_23386,N_22546);
nor U24015 (N_24015,N_23481,N_22849);
nand U24016 (N_24016,N_23399,N_22811);
nand U24017 (N_24017,N_22938,N_22587);
and U24018 (N_24018,N_23724,N_23008);
xor U24019 (N_24019,N_23133,N_23592);
xnor U24020 (N_24020,N_23455,N_23473);
or U24021 (N_24021,N_23224,N_22886);
nand U24022 (N_24022,N_23339,N_23294);
and U24023 (N_24023,N_23698,N_22960);
and U24024 (N_24024,N_23739,N_23005);
and U24025 (N_24025,N_23693,N_23646);
nand U24026 (N_24026,N_23652,N_23630);
and U24027 (N_24027,N_22771,N_23360);
or U24028 (N_24028,N_22575,N_22863);
and U24029 (N_24029,N_23070,N_23047);
or U24030 (N_24030,N_23403,N_23408);
or U24031 (N_24031,N_23181,N_22730);
or U24032 (N_24032,N_23014,N_23747);
nand U24033 (N_24033,N_22636,N_22717);
nand U24034 (N_24034,N_22919,N_22855);
and U24035 (N_24035,N_23236,N_23432);
xor U24036 (N_24036,N_23100,N_23561);
nand U24037 (N_24037,N_23617,N_22670);
nor U24038 (N_24038,N_22792,N_23575);
xnor U24039 (N_24039,N_23516,N_23397);
nor U24040 (N_24040,N_22875,N_22667);
nor U24041 (N_24041,N_22651,N_23659);
and U24042 (N_24042,N_23396,N_23625);
or U24043 (N_24043,N_22711,N_22709);
nor U24044 (N_24044,N_23312,N_22844);
nor U24045 (N_24045,N_22754,N_23319);
or U24046 (N_24046,N_23683,N_23402);
or U24047 (N_24047,N_23061,N_22529);
and U24048 (N_24048,N_23638,N_23632);
nand U24049 (N_24049,N_22823,N_22532);
xor U24050 (N_24050,N_23400,N_22694);
or U24051 (N_24051,N_22922,N_23308);
nor U24052 (N_24052,N_23326,N_23640);
nand U24053 (N_24053,N_22740,N_23147);
nor U24054 (N_24054,N_23317,N_23036);
xor U24055 (N_24055,N_23583,N_23154);
nand U24056 (N_24056,N_23467,N_23673);
xnor U24057 (N_24057,N_22911,N_23494);
nand U24058 (N_24058,N_23175,N_23165);
or U24059 (N_24059,N_23415,N_23212);
xor U24060 (N_24060,N_23207,N_23547);
nor U24061 (N_24061,N_22719,N_22924);
or U24062 (N_24062,N_23532,N_22882);
nor U24063 (N_24063,N_22598,N_22896);
xnor U24064 (N_24064,N_22662,N_23003);
nor U24065 (N_24065,N_22671,N_23259);
and U24066 (N_24066,N_23648,N_23006);
nor U24067 (N_24067,N_23122,N_23356);
or U24068 (N_24068,N_23745,N_23544);
xnor U24069 (N_24069,N_23152,N_22827);
and U24070 (N_24070,N_23701,N_22765);
nor U24071 (N_24071,N_23373,N_22782);
nor U24072 (N_24072,N_23543,N_23500);
xor U24073 (N_24073,N_23717,N_23577);
nand U24074 (N_24074,N_22520,N_22862);
nor U24075 (N_24075,N_22507,N_22937);
and U24076 (N_24076,N_23104,N_22943);
and U24077 (N_24077,N_23016,N_23440);
nand U24078 (N_24078,N_23558,N_23252);
or U24079 (N_24079,N_22726,N_23078);
and U24080 (N_24080,N_23674,N_23082);
nor U24081 (N_24081,N_23300,N_22576);
xor U24082 (N_24082,N_23665,N_23062);
or U24083 (N_24083,N_22913,N_22986);
xor U24084 (N_24084,N_22713,N_23697);
nor U24085 (N_24085,N_23506,N_22806);
xor U24086 (N_24086,N_22867,N_23219);
or U24087 (N_24087,N_23159,N_23741);
and U24088 (N_24088,N_22610,N_23405);
and U24089 (N_24089,N_23513,N_22553);
nor U24090 (N_24090,N_23160,N_22890);
xor U24091 (N_24091,N_22739,N_23545);
nand U24092 (N_24092,N_22828,N_22523);
or U24093 (N_24093,N_22533,N_23214);
and U24094 (N_24094,N_23019,N_22729);
and U24095 (N_24095,N_22513,N_22799);
xnor U24096 (N_24096,N_23462,N_23114);
or U24097 (N_24097,N_23512,N_22846);
or U24098 (N_24098,N_22888,N_23371);
and U24099 (N_24099,N_23571,N_23283);
and U24100 (N_24100,N_23684,N_22936);
nor U24101 (N_24101,N_23384,N_22639);
and U24102 (N_24102,N_23244,N_23174);
or U24103 (N_24103,N_23270,N_22858);
or U24104 (N_24104,N_23559,N_23423);
xnor U24105 (N_24105,N_22878,N_23180);
nor U24106 (N_24106,N_22526,N_23277);
and U24107 (N_24107,N_23280,N_23362);
nor U24108 (N_24108,N_23176,N_22761);
xnor U24109 (N_24109,N_22802,N_22979);
xor U24110 (N_24110,N_23253,N_23155);
xnor U24111 (N_24111,N_23323,N_23428);
and U24112 (N_24112,N_22984,N_22700);
or U24113 (N_24113,N_23246,N_22908);
nor U24114 (N_24114,N_22603,N_22683);
and U24115 (N_24115,N_23196,N_23389);
nor U24116 (N_24116,N_23168,N_22856);
and U24117 (N_24117,N_23391,N_22514);
or U24118 (N_24118,N_22748,N_23170);
xnor U24119 (N_24119,N_22558,N_23116);
and U24120 (N_24120,N_23195,N_23469);
nand U24121 (N_24121,N_23293,N_22854);
nand U24122 (N_24122,N_22530,N_23620);
nand U24123 (N_24123,N_23342,N_23049);
nand U24124 (N_24124,N_23379,N_22625);
nor U24125 (N_24125,N_23117,N_23074);
or U24126 (N_24126,N_22975,N_23298);
or U24127 (N_24127,N_23699,N_23316);
or U24128 (N_24128,N_23151,N_23066);
xor U24129 (N_24129,N_23690,N_23081);
or U24130 (N_24130,N_23031,N_23108);
and U24131 (N_24131,N_22597,N_23051);
nor U24132 (N_24132,N_23605,N_22775);
and U24133 (N_24133,N_23055,N_23398);
xor U24134 (N_24134,N_23378,N_22947);
and U24135 (N_24135,N_22641,N_23136);
or U24136 (N_24136,N_23586,N_23563);
xnor U24137 (N_24137,N_22909,N_22942);
nor U24138 (N_24138,N_23110,N_22701);
xnor U24139 (N_24139,N_23250,N_22519);
nor U24140 (N_24140,N_22731,N_23442);
or U24141 (N_24141,N_22623,N_22987);
or U24142 (N_24142,N_22891,N_22584);
xnor U24143 (N_24143,N_23459,N_22756);
or U24144 (N_24144,N_23260,N_23140);
nor U24145 (N_24145,N_23046,N_22710);
xnor U24146 (N_24146,N_22638,N_23354);
nand U24147 (N_24147,N_22718,N_23474);
nand U24148 (N_24148,N_22817,N_22689);
nand U24149 (N_24149,N_22559,N_22834);
nor U24150 (N_24150,N_23126,N_23496);
nor U24151 (N_24151,N_22916,N_23518);
nor U24152 (N_24152,N_23671,N_23553);
nor U24153 (N_24153,N_23344,N_23421);
xor U24154 (N_24154,N_23737,N_23414);
or U24155 (N_24155,N_23329,N_23086);
xor U24156 (N_24156,N_22773,N_22900);
and U24157 (N_24157,N_23119,N_23600);
and U24158 (N_24158,N_23655,N_22677);
and U24159 (N_24159,N_23366,N_23526);
and U24160 (N_24160,N_22812,N_23732);
or U24161 (N_24161,N_23248,N_23708);
nand U24162 (N_24162,N_22899,N_22777);
nand U24163 (N_24163,N_22501,N_23273);
nor U24164 (N_24164,N_23079,N_22573);
xnor U24165 (N_24165,N_23404,N_23186);
nor U24166 (N_24166,N_22871,N_23736);
and U24167 (N_24167,N_22509,N_22515);
or U24168 (N_24168,N_22696,N_22612);
xnor U24169 (N_24169,N_23321,N_23034);
and U24170 (N_24170,N_23614,N_23534);
xor U24171 (N_24171,N_22620,N_23035);
nand U24172 (N_24172,N_22946,N_23190);
nand U24173 (N_24173,N_23023,N_22894);
or U24174 (N_24174,N_23542,N_22961);
nor U24175 (N_24175,N_23615,N_23390);
nor U24176 (N_24176,N_23285,N_23696);
or U24177 (N_24177,N_23199,N_22500);
or U24178 (N_24178,N_23562,N_22632);
nor U24179 (N_24179,N_22832,N_23368);
nor U24180 (N_24180,N_22688,N_22770);
or U24181 (N_24181,N_23480,N_23375);
nor U24182 (N_24182,N_23581,N_23457);
xor U24183 (N_24183,N_22971,N_22857);
or U24184 (N_24184,N_22562,N_23241);
and U24185 (N_24185,N_23453,N_22669);
or U24186 (N_24186,N_23020,N_23537);
xor U24187 (N_24187,N_23629,N_23643);
or U24188 (N_24188,N_22973,N_23296);
nor U24189 (N_24189,N_22918,N_23691);
or U24190 (N_24190,N_23596,N_22728);
and U24191 (N_24191,N_22666,N_22672);
xor U24192 (N_24192,N_22742,N_23407);
and U24193 (N_24193,N_23680,N_23560);
xor U24194 (N_24194,N_23376,N_22635);
or U24195 (N_24195,N_23490,N_22536);
xnor U24196 (N_24196,N_23628,N_23409);
and U24197 (N_24197,N_23555,N_22522);
or U24198 (N_24198,N_23075,N_22568);
nand U24199 (N_24199,N_23258,N_23678);
or U24200 (N_24200,N_23609,N_22547);
and U24201 (N_24201,N_23548,N_22637);
xnor U24202 (N_24202,N_22744,N_23556);
xor U24203 (N_24203,N_22861,N_22950);
or U24204 (N_24204,N_22628,N_23668);
and U24205 (N_24205,N_23604,N_23662);
xnor U24206 (N_24206,N_22705,N_23447);
nand U24207 (N_24207,N_23608,N_23350);
xor U24208 (N_24208,N_23101,N_23422);
or U24209 (N_24209,N_23071,N_22967);
or U24210 (N_24210,N_23485,N_23492);
nand U24211 (N_24211,N_23576,N_22656);
or U24212 (N_24212,N_23128,N_22935);
or U24213 (N_24213,N_23564,N_23161);
and U24214 (N_24214,N_22545,N_23602);
or U24215 (N_24215,N_23456,N_22580);
or U24216 (N_24216,N_22869,N_22560);
xnor U24217 (N_24217,N_23120,N_22591);
nor U24218 (N_24218,N_22640,N_23164);
nor U24219 (N_24219,N_22679,N_23333);
nand U24220 (N_24220,N_22704,N_23041);
nor U24221 (N_24221,N_23177,N_23091);
nand U24222 (N_24222,N_23094,N_23406);
xor U24223 (N_24223,N_22822,N_22660);
nor U24224 (N_24224,N_23489,N_22564);
nor U24225 (N_24225,N_23519,N_23584);
xnor U24226 (N_24226,N_23163,N_23658);
and U24227 (N_24227,N_23411,N_23118);
or U24228 (N_24228,N_23589,N_23302);
or U24229 (N_24229,N_23522,N_23233);
xnor U24230 (N_24230,N_23642,N_23281);
xnor U24231 (N_24231,N_23714,N_23304);
xnor U24232 (N_24232,N_23208,N_22994);
xor U24233 (N_24233,N_23603,N_23677);
nor U24234 (N_24234,N_22561,N_22825);
nand U24235 (N_24235,N_23619,N_23470);
nor U24236 (N_24236,N_22966,N_22596);
or U24237 (N_24237,N_23073,N_22914);
and U24238 (N_24238,N_22915,N_23027);
nand U24239 (N_24239,N_22599,N_23254);
or U24240 (N_24240,N_23452,N_23245);
and U24241 (N_24241,N_23412,N_23106);
or U24242 (N_24242,N_22983,N_22816);
nor U24243 (N_24243,N_23726,N_22516);
or U24244 (N_24244,N_23616,N_23232);
nor U24245 (N_24245,N_23149,N_23478);
nor U24246 (N_24246,N_22977,N_23418);
xor U24247 (N_24247,N_23288,N_23382);
and U24248 (N_24248,N_22917,N_23169);
or U24249 (N_24249,N_22680,N_23552);
nand U24250 (N_24250,N_22795,N_22796);
xnor U24251 (N_24251,N_23109,N_23363);
xnor U24252 (N_24252,N_23076,N_22991);
xor U24253 (N_24253,N_23068,N_23184);
nand U24254 (N_24254,N_22578,N_23085);
or U24255 (N_24255,N_22521,N_22653);
and U24256 (N_24256,N_23521,N_22998);
xnor U24257 (N_24257,N_22583,N_23146);
or U24258 (N_24258,N_23325,N_23718);
nor U24259 (N_24259,N_22619,N_22604);
nand U24260 (N_24260,N_23475,N_23054);
and U24261 (N_24261,N_23393,N_23570);
or U24262 (N_24262,N_23218,N_22772);
xnor U24263 (N_24263,N_23098,N_23520);
xnor U24264 (N_24264,N_23687,N_23443);
xor U24265 (N_24265,N_22595,N_22673);
nand U24266 (N_24266,N_22904,N_22733);
and U24267 (N_24267,N_23113,N_23477);
and U24268 (N_24268,N_23651,N_23330);
nor U24269 (N_24269,N_22648,N_23359);
xnor U24270 (N_24270,N_23261,N_22600);
xor U24271 (N_24271,N_23206,N_22841);
nor U24272 (N_24272,N_23437,N_23000);
and U24273 (N_24273,N_22693,N_23417);
and U24274 (N_24274,N_23264,N_23123);
or U24275 (N_24275,N_23536,N_23702);
xor U24276 (N_24276,N_22902,N_23352);
nand U24277 (N_24277,N_22860,N_23030);
xor U24278 (N_24278,N_22999,N_23255);
xor U24279 (N_24279,N_22821,N_22809);
nor U24280 (N_24280,N_23265,N_23401);
and U24281 (N_24281,N_23425,N_22872);
xnor U24282 (N_24282,N_23010,N_22789);
nand U24283 (N_24283,N_22659,N_23305);
nand U24284 (N_24284,N_23348,N_22723);
nand U24285 (N_24285,N_23172,N_22887);
and U24286 (N_24286,N_22981,N_22749);
nand U24287 (N_24287,N_23182,N_22958);
or U24288 (N_24288,N_23235,N_22512);
nor U24289 (N_24289,N_22901,N_23748);
nor U24290 (N_24290,N_23209,N_23618);
or U24291 (N_24291,N_23531,N_22903);
xnor U24292 (N_24292,N_23740,N_22627);
or U24293 (N_24293,N_23372,N_23338);
nand U24294 (N_24294,N_23256,N_23320);
and U24295 (N_24295,N_23189,N_22634);
nor U24296 (N_24296,N_22954,N_22758);
xor U24297 (N_24297,N_23102,N_22851);
nor U24298 (N_24298,N_23597,N_22505);
nand U24299 (N_24299,N_22815,N_22605);
xnor U24300 (N_24300,N_23439,N_22751);
xor U24301 (N_24301,N_23037,N_23549);
or U24302 (N_24302,N_23582,N_22735);
nand U24303 (N_24303,N_22955,N_22833);
xnor U24304 (N_24304,N_22631,N_23695);
nor U24305 (N_24305,N_22933,N_22511);
nand U24306 (N_24306,N_23369,N_22959);
and U24307 (N_24307,N_23523,N_23588);
nand U24308 (N_24308,N_23710,N_23324);
nor U24309 (N_24309,N_23007,N_23488);
nor U24310 (N_24310,N_22865,N_23059);
or U24311 (N_24311,N_22691,N_23419);
or U24312 (N_24312,N_22897,N_23093);
or U24313 (N_24313,N_22804,N_22791);
nor U24314 (N_24314,N_23450,N_22814);
nor U24315 (N_24315,N_22835,N_22957);
nand U24316 (N_24316,N_22852,N_22618);
nor U24317 (N_24317,N_22881,N_23661);
nand U24318 (N_24318,N_23187,N_23228);
nand U24319 (N_24319,N_23171,N_22996);
or U24320 (N_24320,N_23502,N_22818);
xor U24321 (N_24321,N_22932,N_23347);
xnor U24322 (N_24322,N_22788,N_22866);
or U24323 (N_24323,N_23357,N_23089);
nand U24324 (N_24324,N_22988,N_23188);
nor U24325 (N_24325,N_23497,N_23131);
nor U24326 (N_24326,N_23664,N_22906);
nand U24327 (N_24327,N_22859,N_23083);
xor U24328 (N_24328,N_22557,N_23237);
xor U24329 (N_24329,N_22776,N_22504);
nor U24330 (N_24330,N_22606,N_23069);
or U24331 (N_24331,N_23185,N_22550);
and U24332 (N_24332,N_23033,N_23569);
xnor U24333 (N_24333,N_23517,N_23479);
or U24334 (N_24334,N_22736,N_22539);
xor U24335 (N_24335,N_23295,N_23013);
or U24336 (N_24336,N_22925,N_23115);
nand U24337 (N_24337,N_22647,N_22980);
xor U24338 (N_24338,N_23612,N_23525);
nor U24339 (N_24339,N_23043,N_23637);
or U24340 (N_24340,N_23290,N_23454);
or U24341 (N_24341,N_22755,N_23508);
xnor U24342 (N_24342,N_22506,N_22518);
nand U24343 (N_24343,N_23716,N_22930);
or U24344 (N_24344,N_23742,N_22714);
nand U24345 (N_24345,N_23689,N_23635);
xnor U24346 (N_24346,N_22972,N_23370);
and U24347 (N_24347,N_23315,N_22759);
xnor U24348 (N_24348,N_23510,N_22725);
xnor U24349 (N_24349,N_23438,N_23721);
nand U24350 (N_24350,N_23336,N_23392);
nand U24351 (N_24351,N_22870,N_23729);
and U24352 (N_24352,N_23194,N_22652);
nand U24353 (N_24353,N_22953,N_22923);
xor U24354 (N_24354,N_23719,N_22654);
nor U24355 (N_24355,N_22503,N_22579);
xnor U24356 (N_24356,N_23009,N_23137);
and U24357 (N_24357,N_22588,N_23738);
and U24358 (N_24358,N_23314,N_23269);
or U24359 (N_24359,N_23029,N_23528);
or U24360 (N_24360,N_23466,N_23381);
nor U24361 (N_24361,N_23345,N_22945);
or U24362 (N_24362,N_23427,N_23056);
nand U24363 (N_24363,N_23743,N_23434);
nand U24364 (N_24364,N_22750,N_23234);
or U24365 (N_24365,N_22706,N_22649);
nand U24366 (N_24366,N_23279,N_23144);
nor U24367 (N_24367,N_23257,N_22697);
xor U24368 (N_24368,N_23744,N_23353);
nor U24369 (N_24369,N_22734,N_22527);
xnor U24370 (N_24370,N_23351,N_23530);
xnor U24371 (N_24371,N_23310,N_23060);
nand U24372 (N_24372,N_23539,N_23383);
and U24373 (N_24373,N_23707,N_23243);
and U24374 (N_24374,N_22781,N_23435);
nor U24375 (N_24375,N_23140,N_23736);
nor U24376 (N_24376,N_22547,N_23353);
and U24377 (N_24377,N_23654,N_22923);
nand U24378 (N_24378,N_23124,N_23415);
and U24379 (N_24379,N_22752,N_23625);
or U24380 (N_24380,N_23412,N_23660);
or U24381 (N_24381,N_22905,N_22863);
xor U24382 (N_24382,N_23386,N_23445);
and U24383 (N_24383,N_23731,N_22915);
and U24384 (N_24384,N_23041,N_23566);
or U24385 (N_24385,N_22724,N_23509);
or U24386 (N_24386,N_23093,N_22577);
or U24387 (N_24387,N_23414,N_22997);
nor U24388 (N_24388,N_23043,N_23388);
xor U24389 (N_24389,N_23633,N_22500);
nor U24390 (N_24390,N_22950,N_22584);
and U24391 (N_24391,N_22699,N_23339);
and U24392 (N_24392,N_23175,N_23578);
or U24393 (N_24393,N_23054,N_23614);
or U24394 (N_24394,N_22725,N_22985);
xnor U24395 (N_24395,N_23121,N_22942);
nand U24396 (N_24396,N_23701,N_22776);
or U24397 (N_24397,N_23714,N_23246);
and U24398 (N_24398,N_23514,N_22620);
and U24399 (N_24399,N_23441,N_22654);
nor U24400 (N_24400,N_23234,N_22856);
xnor U24401 (N_24401,N_23208,N_22781);
nor U24402 (N_24402,N_23336,N_22898);
nand U24403 (N_24403,N_23679,N_23293);
xnor U24404 (N_24404,N_23662,N_23203);
xnor U24405 (N_24405,N_23168,N_23223);
and U24406 (N_24406,N_22892,N_22944);
nand U24407 (N_24407,N_22543,N_22783);
and U24408 (N_24408,N_23503,N_23293);
and U24409 (N_24409,N_22736,N_23499);
and U24410 (N_24410,N_23273,N_23724);
xor U24411 (N_24411,N_23052,N_23579);
and U24412 (N_24412,N_22715,N_23511);
or U24413 (N_24413,N_22635,N_23358);
xor U24414 (N_24414,N_22842,N_23257);
xor U24415 (N_24415,N_23034,N_23651);
xnor U24416 (N_24416,N_22972,N_23041);
nand U24417 (N_24417,N_22524,N_23718);
and U24418 (N_24418,N_22941,N_23596);
nand U24419 (N_24419,N_23108,N_22763);
and U24420 (N_24420,N_22916,N_22875);
and U24421 (N_24421,N_23622,N_23576);
xor U24422 (N_24422,N_23604,N_22794);
or U24423 (N_24423,N_23171,N_23346);
xor U24424 (N_24424,N_23188,N_23274);
and U24425 (N_24425,N_22830,N_23114);
xnor U24426 (N_24426,N_23312,N_23098);
and U24427 (N_24427,N_23382,N_22782);
nand U24428 (N_24428,N_22836,N_23217);
and U24429 (N_24429,N_23182,N_22622);
nand U24430 (N_24430,N_23717,N_22946);
nand U24431 (N_24431,N_22846,N_23192);
xnor U24432 (N_24432,N_22709,N_23362);
nor U24433 (N_24433,N_23200,N_23369);
xor U24434 (N_24434,N_23616,N_23514);
nor U24435 (N_24435,N_22559,N_22929);
and U24436 (N_24436,N_23653,N_23304);
and U24437 (N_24437,N_23024,N_22574);
nand U24438 (N_24438,N_23301,N_23509);
nand U24439 (N_24439,N_23545,N_22520);
nor U24440 (N_24440,N_23501,N_23378);
and U24441 (N_24441,N_23536,N_22553);
or U24442 (N_24442,N_22871,N_23733);
nor U24443 (N_24443,N_23574,N_23290);
nand U24444 (N_24444,N_22913,N_23358);
nand U24445 (N_24445,N_22756,N_23744);
and U24446 (N_24446,N_22996,N_23252);
and U24447 (N_24447,N_23540,N_23030);
nor U24448 (N_24448,N_23709,N_22515);
and U24449 (N_24449,N_23479,N_22864);
nand U24450 (N_24450,N_23268,N_22745);
nand U24451 (N_24451,N_22649,N_22945);
or U24452 (N_24452,N_23393,N_23489);
nand U24453 (N_24453,N_23726,N_23030);
nand U24454 (N_24454,N_22784,N_23399);
nand U24455 (N_24455,N_23176,N_22862);
and U24456 (N_24456,N_23199,N_23608);
nand U24457 (N_24457,N_23157,N_23293);
nor U24458 (N_24458,N_23468,N_23190);
and U24459 (N_24459,N_23672,N_23453);
nor U24460 (N_24460,N_23105,N_23082);
nor U24461 (N_24461,N_23044,N_22834);
or U24462 (N_24462,N_23440,N_23507);
nand U24463 (N_24463,N_23095,N_23031);
or U24464 (N_24464,N_23008,N_23575);
xor U24465 (N_24465,N_23036,N_23000);
xnor U24466 (N_24466,N_23018,N_23439);
xor U24467 (N_24467,N_23678,N_22556);
or U24468 (N_24468,N_22867,N_22530);
nor U24469 (N_24469,N_23465,N_22605);
nor U24470 (N_24470,N_22662,N_23082);
or U24471 (N_24471,N_22801,N_23729);
and U24472 (N_24472,N_23020,N_22580);
or U24473 (N_24473,N_22823,N_23297);
xnor U24474 (N_24474,N_22876,N_23439);
nor U24475 (N_24475,N_23242,N_23391);
and U24476 (N_24476,N_23287,N_22910);
or U24477 (N_24477,N_22640,N_22996);
nand U24478 (N_24478,N_22816,N_23306);
and U24479 (N_24479,N_22799,N_23180);
nand U24480 (N_24480,N_23447,N_23086);
or U24481 (N_24481,N_23279,N_23471);
or U24482 (N_24482,N_23681,N_22670);
or U24483 (N_24483,N_23540,N_22729);
nand U24484 (N_24484,N_23325,N_23368);
and U24485 (N_24485,N_22551,N_23414);
or U24486 (N_24486,N_23500,N_23459);
xnor U24487 (N_24487,N_23713,N_23014);
or U24488 (N_24488,N_22650,N_23408);
nand U24489 (N_24489,N_22763,N_23744);
or U24490 (N_24490,N_23367,N_22957);
xnor U24491 (N_24491,N_23536,N_22761);
or U24492 (N_24492,N_22584,N_23650);
nand U24493 (N_24493,N_23209,N_22707);
or U24494 (N_24494,N_22880,N_22953);
nand U24495 (N_24495,N_22881,N_22969);
xnor U24496 (N_24496,N_23141,N_23379);
or U24497 (N_24497,N_22662,N_22971);
and U24498 (N_24498,N_23460,N_23626);
nor U24499 (N_24499,N_22733,N_23636);
xor U24500 (N_24500,N_23257,N_23503);
nor U24501 (N_24501,N_22617,N_23127);
xor U24502 (N_24502,N_23190,N_23252);
or U24503 (N_24503,N_23298,N_22805);
xnor U24504 (N_24504,N_23621,N_22868);
and U24505 (N_24505,N_23737,N_22762);
xnor U24506 (N_24506,N_22890,N_23534);
or U24507 (N_24507,N_23324,N_22587);
and U24508 (N_24508,N_22810,N_22993);
nor U24509 (N_24509,N_23483,N_23338);
or U24510 (N_24510,N_22927,N_23736);
nor U24511 (N_24511,N_23625,N_22829);
nor U24512 (N_24512,N_22933,N_22921);
and U24513 (N_24513,N_23068,N_22979);
nand U24514 (N_24514,N_23381,N_23622);
or U24515 (N_24515,N_23483,N_23211);
nand U24516 (N_24516,N_22504,N_22765);
nand U24517 (N_24517,N_22644,N_23061);
nor U24518 (N_24518,N_23135,N_22594);
or U24519 (N_24519,N_22511,N_23166);
and U24520 (N_24520,N_23257,N_23301);
and U24521 (N_24521,N_22856,N_23019);
nor U24522 (N_24522,N_23477,N_22500);
or U24523 (N_24523,N_22825,N_23024);
xnor U24524 (N_24524,N_23344,N_23624);
nor U24525 (N_24525,N_23413,N_23179);
xnor U24526 (N_24526,N_23285,N_23170);
or U24527 (N_24527,N_23298,N_22609);
nor U24528 (N_24528,N_22585,N_22707);
nor U24529 (N_24529,N_23516,N_23532);
xor U24530 (N_24530,N_22647,N_22716);
xor U24531 (N_24531,N_23628,N_22517);
nand U24532 (N_24532,N_22587,N_23405);
nor U24533 (N_24533,N_22659,N_22707);
nor U24534 (N_24534,N_22965,N_23359);
and U24535 (N_24535,N_22788,N_23100);
or U24536 (N_24536,N_23352,N_23447);
xor U24537 (N_24537,N_23620,N_23550);
or U24538 (N_24538,N_23238,N_23462);
xnor U24539 (N_24539,N_23012,N_23616);
xor U24540 (N_24540,N_23592,N_23120);
and U24541 (N_24541,N_23180,N_22757);
and U24542 (N_24542,N_23437,N_23635);
nand U24543 (N_24543,N_22718,N_23107);
or U24544 (N_24544,N_23366,N_23472);
xnor U24545 (N_24545,N_23644,N_23373);
xor U24546 (N_24546,N_23674,N_23596);
and U24547 (N_24547,N_23335,N_23078);
nand U24548 (N_24548,N_23435,N_22856);
and U24549 (N_24549,N_22959,N_23143);
nand U24550 (N_24550,N_23419,N_22705);
and U24551 (N_24551,N_23562,N_23342);
or U24552 (N_24552,N_22650,N_23098);
or U24553 (N_24553,N_23278,N_23237);
and U24554 (N_24554,N_23485,N_23354);
nor U24555 (N_24555,N_22544,N_23595);
and U24556 (N_24556,N_23428,N_23303);
nor U24557 (N_24557,N_23432,N_23282);
or U24558 (N_24558,N_23609,N_23340);
xnor U24559 (N_24559,N_23146,N_22627);
xnor U24560 (N_24560,N_22989,N_23330);
nand U24561 (N_24561,N_23084,N_23639);
and U24562 (N_24562,N_23227,N_23697);
nor U24563 (N_24563,N_22710,N_23294);
xor U24564 (N_24564,N_23131,N_22630);
nor U24565 (N_24565,N_22518,N_23102);
nand U24566 (N_24566,N_22605,N_22642);
nor U24567 (N_24567,N_23099,N_23714);
or U24568 (N_24568,N_23431,N_23376);
or U24569 (N_24569,N_22661,N_22736);
xnor U24570 (N_24570,N_22529,N_23181);
nand U24571 (N_24571,N_23037,N_23072);
or U24572 (N_24572,N_23376,N_23551);
and U24573 (N_24573,N_22648,N_23484);
and U24574 (N_24574,N_23053,N_23474);
or U24575 (N_24575,N_23590,N_23367);
or U24576 (N_24576,N_22648,N_22895);
nand U24577 (N_24577,N_23524,N_23014);
nor U24578 (N_24578,N_22528,N_22878);
nor U24579 (N_24579,N_23161,N_22778);
nand U24580 (N_24580,N_22949,N_22815);
nand U24581 (N_24581,N_22945,N_23556);
and U24582 (N_24582,N_22997,N_23101);
nor U24583 (N_24583,N_23479,N_22571);
and U24584 (N_24584,N_22680,N_23611);
or U24585 (N_24585,N_23209,N_22783);
nand U24586 (N_24586,N_22728,N_23036);
nor U24587 (N_24587,N_23634,N_23703);
xor U24588 (N_24588,N_23304,N_22893);
xor U24589 (N_24589,N_23495,N_23427);
xnor U24590 (N_24590,N_23056,N_22591);
or U24591 (N_24591,N_23441,N_23431);
or U24592 (N_24592,N_23325,N_22950);
nor U24593 (N_24593,N_23501,N_22792);
and U24594 (N_24594,N_22783,N_22706);
nor U24595 (N_24595,N_22630,N_22634);
xor U24596 (N_24596,N_22599,N_22978);
nand U24597 (N_24597,N_22628,N_23469);
or U24598 (N_24598,N_22666,N_23559);
or U24599 (N_24599,N_22628,N_22831);
xnor U24600 (N_24600,N_22545,N_22919);
or U24601 (N_24601,N_22929,N_23294);
nand U24602 (N_24602,N_23078,N_22661);
nand U24603 (N_24603,N_22944,N_23664);
nor U24604 (N_24604,N_23734,N_23261);
xnor U24605 (N_24605,N_22797,N_23097);
and U24606 (N_24606,N_23146,N_23346);
nor U24607 (N_24607,N_23243,N_23153);
nand U24608 (N_24608,N_23419,N_23424);
or U24609 (N_24609,N_23586,N_23025);
xor U24610 (N_24610,N_23375,N_23654);
nand U24611 (N_24611,N_22875,N_22752);
or U24612 (N_24612,N_23657,N_23647);
and U24613 (N_24613,N_23735,N_22724);
or U24614 (N_24614,N_23394,N_22715);
xnor U24615 (N_24615,N_23016,N_23271);
and U24616 (N_24616,N_23556,N_22576);
or U24617 (N_24617,N_23661,N_22601);
and U24618 (N_24618,N_23345,N_23500);
nor U24619 (N_24619,N_23326,N_23255);
nand U24620 (N_24620,N_23391,N_22778);
and U24621 (N_24621,N_22822,N_23541);
or U24622 (N_24622,N_23298,N_22513);
nor U24623 (N_24623,N_22846,N_22868);
xor U24624 (N_24624,N_23489,N_23683);
xnor U24625 (N_24625,N_22583,N_23692);
xor U24626 (N_24626,N_23152,N_22775);
and U24627 (N_24627,N_23628,N_22968);
nand U24628 (N_24628,N_22557,N_23310);
nor U24629 (N_24629,N_23162,N_22972);
or U24630 (N_24630,N_23546,N_23313);
or U24631 (N_24631,N_23725,N_22947);
nor U24632 (N_24632,N_23694,N_22511);
xor U24633 (N_24633,N_23033,N_23176);
or U24634 (N_24634,N_22613,N_23093);
or U24635 (N_24635,N_22897,N_23630);
or U24636 (N_24636,N_22968,N_22867);
nand U24637 (N_24637,N_22535,N_23184);
or U24638 (N_24638,N_23058,N_23099);
nor U24639 (N_24639,N_23527,N_23317);
nand U24640 (N_24640,N_23611,N_23105);
or U24641 (N_24641,N_22850,N_22724);
or U24642 (N_24642,N_22958,N_23414);
and U24643 (N_24643,N_22904,N_23488);
xor U24644 (N_24644,N_23566,N_23215);
or U24645 (N_24645,N_22603,N_22779);
nor U24646 (N_24646,N_23105,N_23443);
xor U24647 (N_24647,N_23203,N_23012);
and U24648 (N_24648,N_22796,N_22820);
nand U24649 (N_24649,N_23716,N_23543);
or U24650 (N_24650,N_23161,N_23424);
and U24651 (N_24651,N_23347,N_23349);
nand U24652 (N_24652,N_22608,N_23554);
xnor U24653 (N_24653,N_22814,N_22922);
xnor U24654 (N_24654,N_23518,N_23122);
or U24655 (N_24655,N_23240,N_22583);
and U24656 (N_24656,N_22570,N_23492);
nor U24657 (N_24657,N_22612,N_22572);
nor U24658 (N_24658,N_22532,N_22782);
nand U24659 (N_24659,N_22956,N_23508);
nor U24660 (N_24660,N_23318,N_23640);
nor U24661 (N_24661,N_23204,N_23103);
or U24662 (N_24662,N_23632,N_23689);
xor U24663 (N_24663,N_22712,N_22610);
or U24664 (N_24664,N_23177,N_23141);
or U24665 (N_24665,N_22956,N_23104);
or U24666 (N_24666,N_22948,N_23119);
or U24667 (N_24667,N_23476,N_23146);
xnor U24668 (N_24668,N_23153,N_23681);
nor U24669 (N_24669,N_22647,N_22503);
nand U24670 (N_24670,N_23012,N_23227);
nor U24671 (N_24671,N_22743,N_23192);
and U24672 (N_24672,N_22990,N_22952);
nor U24673 (N_24673,N_23702,N_22949);
nand U24674 (N_24674,N_23434,N_23527);
or U24675 (N_24675,N_22882,N_22787);
and U24676 (N_24676,N_23084,N_23727);
nor U24677 (N_24677,N_22769,N_22510);
or U24678 (N_24678,N_23719,N_22540);
nand U24679 (N_24679,N_22537,N_22894);
nand U24680 (N_24680,N_22786,N_22972);
and U24681 (N_24681,N_23165,N_22947);
or U24682 (N_24682,N_23673,N_23595);
nor U24683 (N_24683,N_23593,N_23183);
nor U24684 (N_24684,N_23084,N_22926);
nor U24685 (N_24685,N_23456,N_23498);
xor U24686 (N_24686,N_22736,N_23545);
or U24687 (N_24687,N_23297,N_23409);
nor U24688 (N_24688,N_23156,N_22825);
or U24689 (N_24689,N_22800,N_23733);
xor U24690 (N_24690,N_23479,N_23660);
nor U24691 (N_24691,N_23449,N_23427);
or U24692 (N_24692,N_23697,N_23362);
nand U24693 (N_24693,N_22895,N_22608);
and U24694 (N_24694,N_23044,N_23396);
and U24695 (N_24695,N_22744,N_23273);
nor U24696 (N_24696,N_22741,N_23485);
nand U24697 (N_24697,N_22716,N_23280);
or U24698 (N_24698,N_22780,N_23636);
nor U24699 (N_24699,N_22818,N_22558);
nand U24700 (N_24700,N_22865,N_23735);
nand U24701 (N_24701,N_23553,N_23258);
and U24702 (N_24702,N_22546,N_23573);
nor U24703 (N_24703,N_23654,N_22563);
nor U24704 (N_24704,N_22693,N_23659);
nand U24705 (N_24705,N_23643,N_23247);
xnor U24706 (N_24706,N_23535,N_23429);
and U24707 (N_24707,N_23312,N_22620);
or U24708 (N_24708,N_23346,N_23135);
and U24709 (N_24709,N_22969,N_23699);
or U24710 (N_24710,N_22843,N_22703);
and U24711 (N_24711,N_22540,N_23642);
nand U24712 (N_24712,N_23271,N_23418);
xnor U24713 (N_24713,N_23287,N_22501);
and U24714 (N_24714,N_23159,N_23190);
and U24715 (N_24715,N_22752,N_23591);
or U24716 (N_24716,N_23676,N_22733);
xor U24717 (N_24717,N_22582,N_23237);
xor U24718 (N_24718,N_22561,N_23322);
nand U24719 (N_24719,N_23246,N_23690);
and U24720 (N_24720,N_22847,N_22702);
or U24721 (N_24721,N_23296,N_23175);
xor U24722 (N_24722,N_22857,N_23534);
xnor U24723 (N_24723,N_23599,N_23440);
xnor U24724 (N_24724,N_22797,N_22551);
nand U24725 (N_24725,N_23297,N_22585);
nor U24726 (N_24726,N_23072,N_23024);
nand U24727 (N_24727,N_22715,N_23427);
or U24728 (N_24728,N_23183,N_23096);
and U24729 (N_24729,N_23742,N_23042);
nor U24730 (N_24730,N_23365,N_23227);
nand U24731 (N_24731,N_23145,N_23335);
nand U24732 (N_24732,N_23003,N_23576);
or U24733 (N_24733,N_22570,N_22725);
and U24734 (N_24734,N_22923,N_23184);
or U24735 (N_24735,N_23618,N_23320);
and U24736 (N_24736,N_22834,N_22632);
nor U24737 (N_24737,N_23149,N_22832);
xnor U24738 (N_24738,N_23078,N_23265);
nand U24739 (N_24739,N_23307,N_23155);
or U24740 (N_24740,N_23030,N_23365);
xor U24741 (N_24741,N_23161,N_23642);
nand U24742 (N_24742,N_22507,N_22626);
and U24743 (N_24743,N_23424,N_23407);
or U24744 (N_24744,N_23272,N_22555);
nand U24745 (N_24745,N_23712,N_23567);
or U24746 (N_24746,N_23741,N_22622);
xor U24747 (N_24747,N_23150,N_23087);
nand U24748 (N_24748,N_22908,N_22662);
nor U24749 (N_24749,N_22951,N_23686);
or U24750 (N_24750,N_23089,N_23659);
nor U24751 (N_24751,N_23109,N_22843);
nor U24752 (N_24752,N_23526,N_22863);
or U24753 (N_24753,N_23525,N_23586);
and U24754 (N_24754,N_23303,N_22868);
nor U24755 (N_24755,N_22840,N_23005);
nand U24756 (N_24756,N_22517,N_23365);
nor U24757 (N_24757,N_23369,N_23502);
nor U24758 (N_24758,N_23121,N_23341);
nor U24759 (N_24759,N_23234,N_22718);
and U24760 (N_24760,N_23609,N_22890);
nor U24761 (N_24761,N_22972,N_23531);
and U24762 (N_24762,N_22682,N_22595);
nand U24763 (N_24763,N_22786,N_23417);
xnor U24764 (N_24764,N_23720,N_22579);
nand U24765 (N_24765,N_22792,N_23303);
nor U24766 (N_24766,N_22831,N_23259);
nor U24767 (N_24767,N_22887,N_22700);
nor U24768 (N_24768,N_22961,N_23390);
or U24769 (N_24769,N_23739,N_23021);
and U24770 (N_24770,N_23359,N_23048);
nand U24771 (N_24771,N_23169,N_22935);
nor U24772 (N_24772,N_23147,N_23017);
nor U24773 (N_24773,N_23506,N_23284);
nor U24774 (N_24774,N_23567,N_23380);
and U24775 (N_24775,N_22542,N_22675);
nand U24776 (N_24776,N_23569,N_22704);
and U24777 (N_24777,N_22913,N_22727);
nor U24778 (N_24778,N_22915,N_23558);
or U24779 (N_24779,N_23139,N_23454);
or U24780 (N_24780,N_23152,N_22852);
xor U24781 (N_24781,N_23350,N_22768);
and U24782 (N_24782,N_23263,N_22825);
xor U24783 (N_24783,N_22976,N_23235);
and U24784 (N_24784,N_22591,N_23080);
xor U24785 (N_24785,N_23694,N_23652);
nand U24786 (N_24786,N_23449,N_23267);
nand U24787 (N_24787,N_22901,N_23214);
xnor U24788 (N_24788,N_23581,N_23651);
nor U24789 (N_24789,N_23743,N_23004);
or U24790 (N_24790,N_22926,N_23663);
and U24791 (N_24791,N_22512,N_23137);
xnor U24792 (N_24792,N_22930,N_23067);
nor U24793 (N_24793,N_23545,N_23688);
or U24794 (N_24794,N_22574,N_22868);
nor U24795 (N_24795,N_22876,N_22797);
or U24796 (N_24796,N_23185,N_23485);
nand U24797 (N_24797,N_23286,N_23524);
and U24798 (N_24798,N_22795,N_23282);
or U24799 (N_24799,N_23639,N_23002);
nor U24800 (N_24800,N_22556,N_23566);
nand U24801 (N_24801,N_23165,N_22776);
or U24802 (N_24802,N_23683,N_23695);
or U24803 (N_24803,N_22992,N_22872);
nor U24804 (N_24804,N_23533,N_23686);
xnor U24805 (N_24805,N_22724,N_23408);
nand U24806 (N_24806,N_22601,N_23598);
xor U24807 (N_24807,N_22847,N_23329);
or U24808 (N_24808,N_22855,N_23467);
nand U24809 (N_24809,N_23034,N_23451);
or U24810 (N_24810,N_22923,N_22726);
nand U24811 (N_24811,N_22547,N_22930);
xor U24812 (N_24812,N_23088,N_23665);
nand U24813 (N_24813,N_22676,N_22732);
or U24814 (N_24814,N_22790,N_22550);
nand U24815 (N_24815,N_22519,N_23587);
xor U24816 (N_24816,N_23496,N_23019);
or U24817 (N_24817,N_23408,N_22686);
xor U24818 (N_24818,N_23266,N_22553);
and U24819 (N_24819,N_23274,N_22723);
nand U24820 (N_24820,N_23138,N_22665);
and U24821 (N_24821,N_22695,N_22702);
and U24822 (N_24822,N_23251,N_23565);
xor U24823 (N_24823,N_22951,N_23715);
nor U24824 (N_24824,N_23450,N_22658);
nand U24825 (N_24825,N_23574,N_22668);
nor U24826 (N_24826,N_22898,N_22611);
xnor U24827 (N_24827,N_22837,N_22527);
xor U24828 (N_24828,N_23160,N_22659);
xnor U24829 (N_24829,N_23274,N_23480);
and U24830 (N_24830,N_23307,N_22558);
nor U24831 (N_24831,N_22751,N_23113);
or U24832 (N_24832,N_22514,N_22970);
nor U24833 (N_24833,N_23666,N_23098);
nor U24834 (N_24834,N_22985,N_23739);
and U24835 (N_24835,N_22649,N_23747);
xnor U24836 (N_24836,N_22672,N_22905);
nor U24837 (N_24837,N_23351,N_22999);
nor U24838 (N_24838,N_22927,N_23591);
nand U24839 (N_24839,N_23628,N_22889);
nor U24840 (N_24840,N_23113,N_23323);
nand U24841 (N_24841,N_22554,N_22535);
or U24842 (N_24842,N_23669,N_23731);
nor U24843 (N_24843,N_22763,N_23508);
and U24844 (N_24844,N_23691,N_23049);
nor U24845 (N_24845,N_22756,N_22824);
and U24846 (N_24846,N_23701,N_23410);
or U24847 (N_24847,N_23544,N_23272);
xnor U24848 (N_24848,N_23118,N_23390);
xor U24849 (N_24849,N_23588,N_23351);
nand U24850 (N_24850,N_23464,N_22867);
and U24851 (N_24851,N_23707,N_22903);
nor U24852 (N_24852,N_22713,N_22633);
nor U24853 (N_24853,N_22545,N_23116);
or U24854 (N_24854,N_22687,N_23324);
and U24855 (N_24855,N_23551,N_23589);
and U24856 (N_24856,N_23420,N_23664);
nor U24857 (N_24857,N_23214,N_23441);
and U24858 (N_24858,N_23201,N_22507);
nand U24859 (N_24859,N_23263,N_23276);
and U24860 (N_24860,N_23689,N_22937);
nand U24861 (N_24861,N_23152,N_23044);
nand U24862 (N_24862,N_22835,N_23419);
xor U24863 (N_24863,N_23551,N_23697);
xor U24864 (N_24864,N_23298,N_22620);
xor U24865 (N_24865,N_23521,N_22772);
or U24866 (N_24866,N_23087,N_22701);
or U24867 (N_24867,N_23610,N_23482);
xor U24868 (N_24868,N_22679,N_23245);
nand U24869 (N_24869,N_23662,N_22977);
nand U24870 (N_24870,N_22798,N_22773);
xor U24871 (N_24871,N_22884,N_23653);
xnor U24872 (N_24872,N_22785,N_23038);
or U24873 (N_24873,N_23512,N_22786);
nand U24874 (N_24874,N_23385,N_23457);
nor U24875 (N_24875,N_23648,N_22733);
or U24876 (N_24876,N_23393,N_23000);
nor U24877 (N_24877,N_22662,N_22716);
or U24878 (N_24878,N_23434,N_23368);
nand U24879 (N_24879,N_22831,N_23454);
or U24880 (N_24880,N_23069,N_23194);
and U24881 (N_24881,N_22946,N_23220);
and U24882 (N_24882,N_23046,N_23711);
nor U24883 (N_24883,N_22841,N_23459);
xor U24884 (N_24884,N_22884,N_23498);
and U24885 (N_24885,N_23566,N_23527);
or U24886 (N_24886,N_23678,N_23072);
or U24887 (N_24887,N_23501,N_22636);
nand U24888 (N_24888,N_22520,N_22988);
nor U24889 (N_24889,N_23209,N_22858);
or U24890 (N_24890,N_23417,N_23568);
nand U24891 (N_24891,N_22921,N_23138);
nor U24892 (N_24892,N_23578,N_23312);
or U24893 (N_24893,N_23126,N_22903);
and U24894 (N_24894,N_23203,N_23559);
xor U24895 (N_24895,N_22845,N_22924);
or U24896 (N_24896,N_23101,N_22676);
and U24897 (N_24897,N_22830,N_22989);
or U24898 (N_24898,N_23266,N_23559);
xnor U24899 (N_24899,N_23527,N_22787);
and U24900 (N_24900,N_22796,N_23731);
or U24901 (N_24901,N_22713,N_22821);
and U24902 (N_24902,N_23153,N_22660);
xor U24903 (N_24903,N_22500,N_23665);
and U24904 (N_24904,N_22926,N_23379);
and U24905 (N_24905,N_23662,N_23041);
or U24906 (N_24906,N_23022,N_23668);
and U24907 (N_24907,N_23189,N_23582);
and U24908 (N_24908,N_23060,N_23164);
xor U24909 (N_24909,N_22653,N_22733);
or U24910 (N_24910,N_23079,N_22822);
xnor U24911 (N_24911,N_23552,N_22986);
nor U24912 (N_24912,N_22789,N_23585);
or U24913 (N_24913,N_22649,N_22910);
nand U24914 (N_24914,N_23691,N_23652);
nand U24915 (N_24915,N_23500,N_22541);
xnor U24916 (N_24916,N_23445,N_23735);
or U24917 (N_24917,N_23718,N_22954);
and U24918 (N_24918,N_23010,N_22935);
or U24919 (N_24919,N_22824,N_23004);
and U24920 (N_24920,N_23712,N_22906);
or U24921 (N_24921,N_23487,N_22971);
and U24922 (N_24922,N_23202,N_22761);
xnor U24923 (N_24923,N_23517,N_22589);
nor U24924 (N_24924,N_23258,N_23153);
and U24925 (N_24925,N_22658,N_23327);
or U24926 (N_24926,N_23189,N_22573);
xnor U24927 (N_24927,N_23683,N_22941);
or U24928 (N_24928,N_23725,N_22874);
xor U24929 (N_24929,N_22880,N_23613);
xnor U24930 (N_24930,N_23202,N_23481);
xnor U24931 (N_24931,N_23086,N_23376);
nor U24932 (N_24932,N_23174,N_22853);
or U24933 (N_24933,N_22759,N_23144);
xnor U24934 (N_24934,N_23583,N_23090);
and U24935 (N_24935,N_22841,N_22550);
nand U24936 (N_24936,N_23687,N_23100);
xnor U24937 (N_24937,N_22767,N_23395);
xnor U24938 (N_24938,N_22703,N_22852);
xnor U24939 (N_24939,N_23749,N_23656);
and U24940 (N_24940,N_22693,N_22797);
xnor U24941 (N_24941,N_22933,N_23073);
and U24942 (N_24942,N_22863,N_22516);
nor U24943 (N_24943,N_22614,N_22772);
or U24944 (N_24944,N_23404,N_23066);
or U24945 (N_24945,N_23060,N_22871);
or U24946 (N_24946,N_22655,N_23205);
xor U24947 (N_24947,N_23091,N_22798);
and U24948 (N_24948,N_23112,N_22587);
nor U24949 (N_24949,N_23257,N_23266);
xor U24950 (N_24950,N_22886,N_22847);
nor U24951 (N_24951,N_22697,N_22719);
xnor U24952 (N_24952,N_23714,N_23010);
or U24953 (N_24953,N_23674,N_23084);
nor U24954 (N_24954,N_23492,N_23117);
nand U24955 (N_24955,N_23440,N_22662);
nand U24956 (N_24956,N_22864,N_23733);
or U24957 (N_24957,N_22813,N_22549);
xor U24958 (N_24958,N_23742,N_23623);
or U24959 (N_24959,N_23240,N_22938);
xor U24960 (N_24960,N_23713,N_23631);
and U24961 (N_24961,N_23091,N_23502);
or U24962 (N_24962,N_22557,N_23395);
xor U24963 (N_24963,N_23720,N_23113);
or U24964 (N_24964,N_23374,N_22671);
nor U24965 (N_24965,N_23528,N_23730);
xnor U24966 (N_24966,N_22724,N_23181);
nand U24967 (N_24967,N_22617,N_22956);
nor U24968 (N_24968,N_23036,N_22925);
and U24969 (N_24969,N_22695,N_22650);
nand U24970 (N_24970,N_23673,N_23244);
nor U24971 (N_24971,N_23412,N_23291);
or U24972 (N_24972,N_22897,N_23012);
xnor U24973 (N_24973,N_22696,N_23509);
nor U24974 (N_24974,N_22777,N_23704);
and U24975 (N_24975,N_22853,N_23280);
xnor U24976 (N_24976,N_22789,N_23390);
and U24977 (N_24977,N_23445,N_23579);
xnor U24978 (N_24978,N_23632,N_23509);
nand U24979 (N_24979,N_22937,N_23179);
nor U24980 (N_24980,N_23003,N_22530);
or U24981 (N_24981,N_22821,N_23334);
or U24982 (N_24982,N_22957,N_23511);
and U24983 (N_24983,N_22552,N_22742);
nor U24984 (N_24984,N_23425,N_23308);
nor U24985 (N_24985,N_23736,N_23123);
nand U24986 (N_24986,N_22718,N_23155);
nor U24987 (N_24987,N_23012,N_22648);
nand U24988 (N_24988,N_23681,N_22914);
or U24989 (N_24989,N_22646,N_22950);
or U24990 (N_24990,N_23710,N_22925);
nand U24991 (N_24991,N_22827,N_22951);
nand U24992 (N_24992,N_22520,N_22871);
and U24993 (N_24993,N_22748,N_23524);
nand U24994 (N_24994,N_23234,N_22937);
xor U24995 (N_24995,N_22863,N_22500);
nor U24996 (N_24996,N_23086,N_22799);
and U24997 (N_24997,N_23290,N_23221);
or U24998 (N_24998,N_23687,N_23189);
and U24999 (N_24999,N_23692,N_23151);
xor UO_0 (O_0,N_24603,N_23932);
nand UO_1 (O_1,N_24365,N_23802);
nor UO_2 (O_2,N_24640,N_24025);
nor UO_3 (O_3,N_24285,N_24691);
or UO_4 (O_4,N_24490,N_24489);
nor UO_5 (O_5,N_24755,N_24429);
nand UO_6 (O_6,N_24065,N_24628);
nand UO_7 (O_7,N_24898,N_24487);
nor UO_8 (O_8,N_24103,N_24060);
nor UO_9 (O_9,N_24602,N_24294);
nand UO_10 (O_10,N_24350,N_24889);
nor UO_11 (O_11,N_24968,N_24099);
or UO_12 (O_12,N_23976,N_24195);
nor UO_13 (O_13,N_24237,N_24380);
or UO_14 (O_14,N_24581,N_24054);
nand UO_15 (O_15,N_24770,N_24960);
nor UO_16 (O_16,N_24647,N_24503);
nor UO_17 (O_17,N_23903,N_23828);
nor UO_18 (O_18,N_24062,N_24921);
xnor UO_19 (O_19,N_24355,N_24605);
and UO_20 (O_20,N_24506,N_24582);
nand UO_21 (O_21,N_24068,N_23959);
and UO_22 (O_22,N_24318,N_24008);
xor UO_23 (O_23,N_24979,N_24223);
xor UO_24 (O_24,N_24533,N_24679);
nand UO_25 (O_25,N_23982,N_24173);
xor UO_26 (O_26,N_24416,N_24015);
xor UO_27 (O_27,N_24336,N_23837);
and UO_28 (O_28,N_24729,N_24048);
nand UO_29 (O_29,N_23852,N_24804);
or UO_30 (O_30,N_23908,N_24807);
and UO_31 (O_31,N_24041,N_24282);
xnor UO_32 (O_32,N_23930,N_24609);
or UO_33 (O_33,N_24904,N_24480);
and UO_34 (O_34,N_24808,N_24090);
or UO_35 (O_35,N_23783,N_23896);
xor UO_36 (O_36,N_24732,N_24339);
or UO_37 (O_37,N_23769,N_23818);
nand UO_38 (O_38,N_24585,N_24089);
and UO_39 (O_39,N_24984,N_24427);
xor UO_40 (O_40,N_24034,N_24678);
or UO_41 (O_41,N_24649,N_24391);
nor UO_42 (O_42,N_24822,N_23919);
and UO_43 (O_43,N_24112,N_24353);
xor UO_44 (O_44,N_24337,N_24650);
and UO_45 (O_45,N_24295,N_24915);
nor UO_46 (O_46,N_24660,N_24164);
nand UO_47 (O_47,N_24159,N_24162);
or UO_48 (O_48,N_24619,N_24593);
or UO_49 (O_49,N_24260,N_24875);
nand UO_50 (O_50,N_23934,N_24606);
nor UO_51 (O_51,N_23822,N_24927);
and UO_52 (O_52,N_24109,N_24406);
xnor UO_53 (O_53,N_24283,N_23833);
xnor UO_54 (O_54,N_24956,N_24623);
nor UO_55 (O_55,N_24893,N_24987);
or UO_56 (O_56,N_24839,N_24202);
or UO_57 (O_57,N_24706,N_24188);
or UO_58 (O_58,N_24595,N_24111);
or UO_59 (O_59,N_24727,N_24645);
xor UO_60 (O_60,N_23878,N_24363);
or UO_61 (O_61,N_23964,N_24383);
nand UO_62 (O_62,N_24870,N_24996);
nor UO_63 (O_63,N_24771,N_24307);
or UO_64 (O_64,N_23801,N_24346);
xor UO_65 (O_65,N_24936,N_24723);
and UO_66 (O_66,N_24475,N_24305);
nor UO_67 (O_67,N_24180,N_24107);
xor UO_68 (O_68,N_24143,N_24241);
nand UO_69 (O_69,N_24174,N_24097);
nand UO_70 (O_70,N_24478,N_24254);
xor UO_71 (O_71,N_24855,N_24695);
xor UO_72 (O_72,N_24117,N_24945);
xor UO_73 (O_73,N_24995,N_24952);
or UO_74 (O_74,N_23840,N_24273);
nor UO_75 (O_75,N_24354,N_24638);
xor UO_76 (O_76,N_24183,N_23827);
nand UO_77 (O_77,N_24539,N_24262);
nor UO_78 (O_78,N_23987,N_24953);
nand UO_79 (O_79,N_24309,N_24287);
nand UO_80 (O_80,N_23891,N_24225);
nand UO_81 (O_81,N_24063,N_24018);
xor UO_82 (O_82,N_24738,N_24409);
nor UO_83 (O_83,N_24447,N_24950);
nand UO_84 (O_84,N_24718,N_23963);
nor UO_85 (O_85,N_24516,N_23948);
or UO_86 (O_86,N_23916,N_24269);
xor UO_87 (O_87,N_24786,N_24003);
nor UO_88 (O_88,N_24308,N_24127);
nor UO_89 (O_89,N_24298,N_24525);
or UO_90 (O_90,N_23800,N_24209);
nand UO_91 (O_91,N_23753,N_23944);
or UO_92 (O_92,N_23792,N_24526);
or UO_93 (O_93,N_24425,N_24395);
xor UO_94 (O_94,N_24630,N_24458);
xor UO_95 (O_95,N_24887,N_24163);
or UO_96 (O_96,N_24121,N_23933);
nand UO_97 (O_97,N_24890,N_24378);
and UO_98 (O_98,N_24256,N_24027);
nor UO_99 (O_99,N_24876,N_24873);
nor UO_100 (O_100,N_24912,N_23847);
xor UO_101 (O_101,N_24798,N_24944);
xnor UO_102 (O_102,N_24144,N_24083);
and UO_103 (O_103,N_23914,N_24922);
nor UO_104 (O_104,N_24125,N_24930);
and UO_105 (O_105,N_24423,N_23907);
or UO_106 (O_106,N_23756,N_23813);
xor UO_107 (O_107,N_24126,N_24325);
nand UO_108 (O_108,N_24087,N_24926);
xnor UO_109 (O_109,N_24049,N_24712);
nor UO_110 (O_110,N_23971,N_24001);
nand UO_111 (O_111,N_24080,N_24999);
nor UO_112 (O_112,N_24805,N_24150);
and UO_113 (O_113,N_24499,N_24179);
or UO_114 (O_114,N_24574,N_24819);
and UO_115 (O_115,N_24616,N_24779);
and UO_116 (O_116,N_24741,N_24633);
nand UO_117 (O_117,N_24370,N_24171);
or UO_118 (O_118,N_24374,N_24253);
nand UO_119 (O_119,N_24698,N_24338);
and UO_120 (O_120,N_24055,N_23946);
nor UO_121 (O_121,N_24651,N_24730);
nor UO_122 (O_122,N_24643,N_24009);
and UO_123 (O_123,N_24219,N_23968);
nand UO_124 (O_124,N_24787,N_24056);
nor UO_125 (O_125,N_24737,N_24011);
or UO_126 (O_126,N_24459,N_24834);
or UO_127 (O_127,N_24542,N_24557);
nand UO_128 (O_128,N_24705,N_24497);
xnor UO_129 (O_129,N_23758,N_23863);
and UO_130 (O_130,N_24994,N_24841);
xor UO_131 (O_131,N_23879,N_24428);
xnor UO_132 (O_132,N_24182,N_23862);
nor UO_133 (O_133,N_24012,N_24369);
xnor UO_134 (O_134,N_24498,N_24147);
nand UO_135 (O_135,N_24572,N_24803);
and UO_136 (O_136,N_24884,N_23777);
nand UO_137 (O_137,N_24275,N_24442);
and UO_138 (O_138,N_23767,N_24563);
nand UO_139 (O_139,N_24991,N_24510);
nand UO_140 (O_140,N_23811,N_24797);
and UO_141 (O_141,N_24733,N_24684);
nor UO_142 (O_142,N_23877,N_24760);
and UO_143 (O_143,N_24594,N_24371);
nor UO_144 (O_144,N_24659,N_23956);
nand UO_145 (O_145,N_24666,N_23958);
and UO_146 (O_146,N_23868,N_24512);
xnor UO_147 (O_147,N_24972,N_24907);
xnor UO_148 (O_148,N_24813,N_24045);
nand UO_149 (O_149,N_24610,N_24746);
or UO_150 (O_150,N_24096,N_24064);
nor UO_151 (O_151,N_24997,N_23803);
xnor UO_152 (O_152,N_24006,N_24982);
nor UO_153 (O_153,N_24983,N_23910);
xor UO_154 (O_154,N_23771,N_24759);
nor UO_155 (O_155,N_24550,N_24719);
or UO_156 (O_156,N_24901,N_24686);
or UO_157 (O_157,N_24569,N_24985);
nor UO_158 (O_158,N_24024,N_23804);
nor UO_159 (O_159,N_24270,N_24136);
or UO_160 (O_160,N_24030,N_23761);
nand UO_161 (O_161,N_24743,N_24883);
and UO_162 (O_162,N_24035,N_24867);
nand UO_163 (O_163,N_23760,N_23839);
nor UO_164 (O_164,N_24522,N_24840);
or UO_165 (O_165,N_24830,N_24251);
or UO_166 (O_166,N_24992,N_24675);
nand UO_167 (O_167,N_24359,N_24820);
or UO_168 (O_168,N_24233,N_23940);
xnor UO_169 (O_169,N_24259,N_23764);
xor UO_170 (O_170,N_23941,N_24155);
xnor UO_171 (O_171,N_24860,N_24192);
and UO_172 (O_172,N_23843,N_24702);
xor UO_173 (O_173,N_23985,N_24778);
xnor UO_174 (O_174,N_24361,N_24925);
and UO_175 (O_175,N_24366,N_23989);
and UO_176 (O_176,N_24198,N_24614);
nor UO_177 (O_177,N_24485,N_24507);
or UO_178 (O_178,N_24882,N_24909);
nor UO_179 (O_179,N_23966,N_23912);
xnor UO_180 (O_180,N_24468,N_24796);
nand UO_181 (O_181,N_24954,N_24976);
and UO_182 (O_182,N_24026,N_24440);
and UO_183 (O_183,N_23766,N_23781);
xnor UO_184 (O_184,N_24313,N_24848);
nor UO_185 (O_185,N_24343,N_24946);
or UO_186 (O_186,N_24123,N_24288);
nor UO_187 (O_187,N_24250,N_23816);
and UO_188 (O_188,N_24078,N_24340);
nor UO_189 (O_189,N_24652,N_24599);
or UO_190 (O_190,N_24825,N_24948);
and UO_191 (O_191,N_24239,N_24501);
or UO_192 (O_192,N_23913,N_24735);
nand UO_193 (O_193,N_24553,N_23911);
xnor UO_194 (O_194,N_24443,N_24810);
nor UO_195 (O_195,N_24221,N_23820);
nand UO_196 (O_196,N_24959,N_23943);
nor UO_197 (O_197,N_23750,N_24433);
nand UO_198 (O_198,N_24981,N_24879);
and UO_199 (O_199,N_24693,N_24415);
nand UO_200 (O_200,N_23988,N_24407);
or UO_201 (O_201,N_24410,N_24726);
or UO_202 (O_202,N_24524,N_24680);
nand UO_203 (O_203,N_24128,N_24255);
nor UO_204 (O_204,N_24878,N_23845);
and UO_205 (O_205,N_24265,N_24627);
xor UO_206 (O_206,N_24894,N_24583);
and UO_207 (O_207,N_24906,N_24913);
nor UO_208 (O_208,N_24677,N_23817);
or UO_209 (O_209,N_24687,N_23876);
nand UO_210 (O_210,N_24213,N_23775);
nor UO_211 (O_211,N_24281,N_24364);
nand UO_212 (O_212,N_23901,N_24699);
and UO_213 (O_213,N_24276,N_24607);
or UO_214 (O_214,N_24767,N_24296);
xor UO_215 (O_215,N_24271,N_24314);
nand UO_216 (O_216,N_24775,N_24604);
or UO_217 (O_217,N_24036,N_24788);
or UO_218 (O_218,N_24465,N_23762);
or UO_219 (O_219,N_23978,N_23857);
and UO_220 (O_220,N_24509,N_24621);
or UO_221 (O_221,N_23854,N_24432);
and UO_222 (O_222,N_24812,N_24216);
nand UO_223 (O_223,N_23942,N_24717);
nor UO_224 (O_224,N_24935,N_24115);
xnor UO_225 (O_225,N_24360,N_23994);
and UO_226 (O_226,N_24491,N_24838);
nand UO_227 (O_227,N_24843,N_24244);
and UO_228 (O_228,N_24849,N_24851);
and UO_229 (O_229,N_24565,N_24561);
or UO_230 (O_230,N_24790,N_24301);
and UO_231 (O_231,N_24257,N_24093);
nor UO_232 (O_232,N_23888,N_24709);
or UO_233 (O_233,N_24701,N_24274);
nor UO_234 (O_234,N_24757,N_24508);
nand UO_235 (O_235,N_24937,N_24158);
nand UO_236 (O_236,N_24148,N_24249);
nor UO_237 (O_237,N_24368,N_24100);
and UO_238 (O_238,N_24502,N_24302);
nor UO_239 (O_239,N_24470,N_24362);
or UO_240 (O_240,N_24777,N_24279);
and UO_241 (O_241,N_24082,N_23751);
and UO_242 (O_242,N_24654,N_23905);
and UO_243 (O_243,N_24773,N_23929);
nand UO_244 (O_244,N_23979,N_23961);
nor UO_245 (O_245,N_24153,N_24341);
nor UO_246 (O_246,N_24005,N_24869);
nor UO_247 (O_247,N_24940,N_23794);
xor UO_248 (O_248,N_24505,N_24970);
nand UO_249 (O_249,N_24205,N_24208);
xor UO_250 (O_250,N_24092,N_24450);
and UO_251 (O_251,N_24020,N_23831);
nor UO_252 (O_252,N_24801,N_24449);
nand UO_253 (O_253,N_23779,N_24392);
or UO_254 (O_254,N_24232,N_23938);
xor UO_255 (O_255,N_24795,N_24220);
nor UO_256 (O_256,N_24031,N_24792);
nand UO_257 (O_257,N_24028,N_24306);
nor UO_258 (O_258,N_23830,N_24891);
nand UO_259 (O_259,N_24817,N_24769);
xor UO_260 (O_260,N_24567,N_24226);
and UO_261 (O_261,N_24844,N_24685);
or UO_262 (O_262,N_24245,N_24242);
xnor UO_263 (O_263,N_23990,N_24334);
or UO_264 (O_264,N_23995,N_24897);
and UO_265 (O_265,N_23867,N_24004);
nor UO_266 (O_266,N_24067,N_23898);
or UO_267 (O_267,N_24529,N_23873);
and UO_268 (O_268,N_24856,N_24289);
nor UO_269 (O_269,N_24311,N_24218);
and UO_270 (O_270,N_24696,N_24038);
nand UO_271 (O_271,N_23834,N_24070);
and UO_272 (O_272,N_24482,N_24157);
nor UO_273 (O_273,N_24942,N_24077);
xnor UO_274 (O_274,N_24439,N_24472);
xnor UO_275 (O_275,N_24133,N_24412);
nand UO_276 (O_276,N_23759,N_24231);
and UO_277 (O_277,N_24895,N_24486);
nand UO_278 (O_278,N_23928,N_24765);
xnor UO_279 (O_279,N_24168,N_23962);
and UO_280 (O_280,N_24252,N_24980);
nor UO_281 (O_281,N_24629,N_24978);
nor UO_282 (O_282,N_24227,N_24931);
nor UO_283 (O_283,N_24074,N_23795);
nand UO_284 (O_284,N_24784,N_23974);
nor UO_285 (O_285,N_24170,N_24632);
and UO_286 (O_286,N_24753,N_23814);
nor UO_287 (O_287,N_24929,N_24248);
and UO_288 (O_288,N_24319,N_23780);
and UO_289 (O_289,N_23874,N_24347);
xnor UO_290 (O_290,N_24105,N_24880);
or UO_291 (O_291,N_24393,N_24124);
and UO_292 (O_292,N_24246,N_24664);
nand UO_293 (O_293,N_24356,N_23782);
and UO_294 (O_294,N_24731,N_24961);
and UO_295 (O_295,N_24555,N_24258);
nor UO_296 (O_296,N_24417,N_24419);
or UO_297 (O_297,N_24010,N_24332);
xnor UO_298 (O_298,N_24612,N_23846);
xnor UO_299 (O_299,N_24642,N_24513);
nor UO_300 (O_300,N_24772,N_24998);
or UO_301 (O_301,N_24016,N_24175);
xor UO_302 (O_302,N_24426,N_24923);
nor UO_303 (O_303,N_23784,N_24591);
or UO_304 (O_304,N_23860,N_23824);
and UO_305 (O_305,N_24973,N_23778);
nand UO_306 (O_306,N_23810,N_24316);
or UO_307 (O_307,N_24816,N_24530);
nand UO_308 (O_308,N_24580,N_24665);
and UO_309 (O_309,N_23980,N_24694);
or UO_310 (O_310,N_24492,N_23981);
nor UO_311 (O_311,N_23895,N_24655);
nor UO_312 (O_312,N_24920,N_24613);
or UO_313 (O_313,N_23773,N_24657);
or UO_314 (O_314,N_24310,N_24578);
and UO_315 (O_315,N_24754,N_24333);
and UO_316 (O_316,N_23832,N_24079);
nor UO_317 (O_317,N_24413,N_24545);
nand UO_318 (O_318,N_24152,N_24800);
or UO_319 (O_319,N_24908,N_24634);
nor UO_320 (O_320,N_24763,N_24540);
nand UO_321 (O_321,N_24520,N_24431);
and UO_322 (O_322,N_24191,N_24918);
nor UO_323 (O_323,N_24794,N_24290);
nand UO_324 (O_324,N_24683,N_24877);
nand UO_325 (O_325,N_24046,N_24871);
or UO_326 (O_326,N_24326,N_24137);
xnor UO_327 (O_327,N_24076,N_24674);
nor UO_328 (O_328,N_24536,N_24688);
nor UO_329 (O_329,N_23902,N_23972);
nor UO_330 (O_330,N_24139,N_23836);
or UO_331 (O_331,N_24955,N_24352);
and UO_332 (O_332,N_24385,N_24791);
nand UO_333 (O_333,N_23806,N_24892);
and UO_334 (O_334,N_23937,N_24806);
and UO_335 (O_335,N_24002,N_24943);
and UO_336 (O_336,N_24330,N_24405);
xnor UO_337 (O_337,N_24297,N_24122);
nand UO_338 (O_338,N_24905,N_24132);
xor UO_339 (O_339,N_23787,N_24761);
nand UO_340 (O_340,N_23848,N_23996);
nor UO_341 (O_341,N_24853,N_24019);
xor UO_342 (O_342,N_24543,N_24900);
and UO_343 (O_343,N_24783,N_24521);
nand UO_344 (O_344,N_24451,N_24858);
nand UO_345 (O_345,N_24456,N_24881);
nor UO_346 (O_346,N_24776,N_24689);
nand UO_347 (O_347,N_24750,N_24764);
nand UO_348 (O_348,N_24455,N_24528);
and UO_349 (O_349,N_24663,N_23993);
nor UO_350 (O_350,N_24514,N_24420);
nor UO_351 (O_351,N_24061,N_24044);
or UO_352 (O_352,N_24444,N_24495);
and UO_353 (O_353,N_23886,N_24592);
or UO_354 (O_354,N_24989,N_23998);
and UO_355 (O_355,N_24401,N_24094);
or UO_356 (O_356,N_23909,N_23859);
and UO_357 (O_357,N_24230,N_23973);
and UO_358 (O_358,N_24351,N_24146);
and UO_359 (O_359,N_24547,N_24344);
nand UO_360 (O_360,N_24007,N_24481);
or UO_361 (O_361,N_24704,N_24934);
or UO_362 (O_362,N_24477,N_23797);
and UO_363 (O_363,N_24211,N_24375);
xor UO_364 (O_364,N_24430,N_23881);
or UO_365 (O_365,N_24398,N_24197);
nor UO_366 (O_366,N_24466,N_24032);
or UO_367 (O_367,N_23880,N_24571);
nand UO_368 (O_368,N_23997,N_24672);
nand UO_369 (O_369,N_24414,N_24224);
or UO_370 (O_370,N_24720,N_24165);
xnor UO_371 (O_371,N_24990,N_24404);
nand UO_372 (O_372,N_24329,N_24102);
and UO_373 (O_373,N_23935,N_24728);
nor UO_374 (O_374,N_24824,N_24247);
and UO_375 (O_375,N_24899,N_24462);
or UO_376 (O_376,N_23922,N_24228);
nand UO_377 (O_377,N_23798,N_24831);
xor UO_378 (O_378,N_24865,N_23918);
or UO_379 (O_379,N_23768,N_24418);
or UO_380 (O_380,N_24399,N_24130);
xor UO_381 (O_381,N_24902,N_24559);
xor UO_382 (O_382,N_24268,N_24129);
or UO_383 (O_383,N_23788,N_24039);
nand UO_384 (O_384,N_24110,N_23936);
xnor UO_385 (O_385,N_24322,N_24053);
or UO_386 (O_386,N_24671,N_24071);
or UO_387 (O_387,N_24681,N_24312);
xnor UO_388 (O_388,N_24747,N_24185);
xor UO_389 (O_389,N_23844,N_24138);
xnor UO_390 (O_390,N_23849,N_24859);
or UO_391 (O_391,N_24267,N_23821);
xnor UO_392 (O_392,N_24742,N_24119);
and UO_393 (O_393,N_24300,N_24161);
nand UO_394 (O_394,N_24888,N_24240);
and UO_395 (O_395,N_23893,N_23770);
nor UO_396 (O_396,N_24957,N_23950);
nand UO_397 (O_397,N_24331,N_24091);
nand UO_398 (O_398,N_24217,N_23900);
or UO_399 (O_399,N_24386,N_24264);
or UO_400 (O_400,N_24676,N_24377);
or UO_401 (O_401,N_24611,N_24075);
and UO_402 (O_402,N_24552,N_24966);
nor UO_403 (O_403,N_24656,N_24523);
xor UO_404 (O_404,N_24641,N_24903);
nand UO_405 (O_405,N_24141,N_24172);
nand UO_406 (O_406,N_24780,N_24852);
nor UO_407 (O_407,N_24022,N_24376);
or UO_408 (O_408,N_24199,N_23957);
nor UO_409 (O_409,N_24722,N_24342);
xnor UO_410 (O_410,N_24328,N_24573);
and UO_411 (O_411,N_23960,N_24500);
and UO_412 (O_412,N_24846,N_24568);
xnor UO_413 (O_413,N_24367,N_24081);
nand UO_414 (O_414,N_24394,N_24639);
or UO_415 (O_415,N_24176,N_24445);
or UO_416 (O_416,N_24789,N_24716);
or UO_417 (O_417,N_23838,N_24734);
nor UO_418 (O_418,N_23842,N_24886);
xor UO_419 (O_419,N_24304,N_24828);
nand UO_420 (O_420,N_23815,N_24280);
or UO_421 (O_421,N_24673,N_24043);
or UO_422 (O_422,N_24739,N_24584);
nor UO_423 (O_423,N_24622,N_24668);
nand UO_424 (O_424,N_23986,N_24576);
nand UO_425 (O_425,N_24988,N_24842);
or UO_426 (O_426,N_24452,N_24919);
xor UO_427 (O_427,N_23789,N_24626);
nor UO_428 (O_428,N_23765,N_24862);
xor UO_429 (O_429,N_23931,N_23864);
nand UO_430 (O_430,N_24118,N_24758);
or UO_431 (O_431,N_24448,N_24947);
nand UO_432 (O_432,N_23984,N_23920);
nand UO_433 (O_433,N_24600,N_24597);
nor UO_434 (O_434,N_24924,N_24013);
xor UO_435 (O_435,N_24203,N_24204);
nand UO_436 (O_436,N_24186,N_24042);
nor UO_437 (O_437,N_24424,N_24740);
nor UO_438 (O_438,N_23927,N_24184);
or UO_439 (O_439,N_24400,N_24864);
or UO_440 (O_440,N_23808,N_23826);
or UO_441 (O_441,N_24177,N_23865);
or UO_442 (O_442,N_24169,N_24151);
nand UO_443 (O_443,N_24167,N_24964);
and UO_444 (O_444,N_23917,N_24537);
nand UO_445 (O_445,N_23897,N_24637);
nor UO_446 (O_446,N_24558,N_24751);
and UO_447 (O_447,N_24857,N_24744);
xnor UO_448 (O_448,N_24471,N_24236);
and UO_449 (O_449,N_24562,N_24190);
nand UO_450 (O_450,N_24166,N_24261);
xnor UO_451 (O_451,N_24636,N_23921);
and UO_452 (O_452,N_24993,N_23870);
or UO_453 (O_453,N_23882,N_24598);
and UO_454 (O_454,N_24441,N_24653);
or UO_455 (O_455,N_24560,N_24483);
nand UO_456 (O_456,N_24617,N_24238);
nand UO_457 (O_457,N_24135,N_23969);
and UO_458 (O_458,N_24963,N_24866);
nor UO_459 (O_459,N_24396,N_24464);
and UO_460 (O_460,N_24615,N_23850);
or UO_461 (O_461,N_24868,N_24662);
or UO_462 (O_462,N_23899,N_24974);
nand UO_463 (O_463,N_24212,N_24863);
nor UO_464 (O_464,N_23774,N_24762);
and UO_465 (O_465,N_23786,N_23871);
or UO_466 (O_466,N_24620,N_24736);
xor UO_467 (O_467,N_24434,N_24278);
and UO_468 (O_468,N_24785,N_24818);
nand UO_469 (O_469,N_23755,N_24967);
or UO_470 (O_470,N_24140,N_23977);
xnor UO_471 (O_471,N_23796,N_23752);
nand UO_472 (O_472,N_24476,N_23809);
xnor UO_473 (O_473,N_24835,N_24711);
or UO_474 (O_474,N_23992,N_24057);
xor UO_475 (O_475,N_23866,N_24291);
and UO_476 (O_476,N_23965,N_24896);
nor UO_477 (O_477,N_24021,N_24201);
xnor UO_478 (O_478,N_24544,N_24682);
nor UO_479 (O_479,N_24234,N_24799);
and UO_480 (O_480,N_24293,N_24323);
and UO_481 (O_481,N_24532,N_24531);
xnor UO_482 (O_482,N_24556,N_24658);
nor UO_483 (O_483,N_24874,N_24390);
nor UO_484 (O_484,N_24131,N_23835);
nand UO_485 (O_485,N_24387,N_24348);
nand UO_486 (O_486,N_23875,N_24266);
or UO_487 (O_487,N_24335,N_24910);
or UO_488 (O_488,N_24469,N_24134);
and UO_489 (O_489,N_24721,N_24535);
or UO_490 (O_490,N_24541,N_24749);
nand UO_491 (O_491,N_24040,N_24949);
or UO_492 (O_492,N_24527,N_24850);
or UO_493 (O_493,N_24768,N_23772);
nand UO_494 (O_494,N_24411,N_24029);
nor UO_495 (O_495,N_24814,N_23904);
and UO_496 (O_496,N_24670,N_23791);
nor UO_497 (O_497,N_24938,N_24194);
nor UO_498 (O_498,N_24579,N_24460);
or UO_499 (O_499,N_24854,N_24113);
nor UO_500 (O_500,N_23999,N_24518);
and UO_501 (O_501,N_24690,N_23967);
xor UO_502 (O_502,N_23812,N_24725);
xnor UO_503 (O_503,N_24618,N_23953);
and UO_504 (O_504,N_24088,N_24590);
and UO_505 (O_505,N_24206,N_23885);
nor UO_506 (O_506,N_24292,N_24815);
xnor UO_507 (O_507,N_24454,N_24037);
xnor UO_508 (O_508,N_24023,N_23819);
nor UO_509 (O_509,N_24971,N_23952);
nor UO_510 (O_510,N_24085,N_23858);
and UO_511 (O_511,N_24120,N_24108);
or UO_512 (O_512,N_24145,N_24357);
and UO_513 (O_513,N_24154,N_23841);
and UO_514 (O_514,N_24534,N_24832);
xor UO_515 (O_515,N_24086,N_24000);
and UO_516 (O_516,N_23757,N_24193);
or UO_517 (O_517,N_24517,N_23872);
xor UO_518 (O_518,N_24697,N_24916);
nor UO_519 (O_519,N_24210,N_23763);
nand UO_520 (O_520,N_24149,N_24546);
or UO_521 (O_521,N_24207,N_24229);
or UO_522 (O_522,N_23855,N_24969);
nand UO_523 (O_523,N_24243,N_24836);
nor UO_524 (O_524,N_24438,N_24667);
nor UO_525 (O_525,N_24435,N_24802);
xnor UO_526 (O_526,N_23861,N_24885);
or UO_527 (O_527,N_23851,N_24504);
nand UO_528 (O_528,N_24196,N_24284);
and UO_529 (O_529,N_24457,N_24461);
xor UO_530 (O_530,N_24975,N_24700);
nand UO_531 (O_531,N_23939,N_24845);
and UO_532 (O_532,N_24017,N_24277);
or UO_533 (O_533,N_24084,N_24811);
and UO_534 (O_534,N_24156,N_24631);
nand UO_535 (O_535,N_24554,N_24837);
nor UO_536 (O_536,N_24511,N_24272);
nand UO_537 (O_537,N_23776,N_23951);
and UO_538 (O_538,N_24928,N_24349);
and UO_539 (O_539,N_24382,N_24826);
nor UO_540 (O_540,N_24214,N_24625);
or UO_541 (O_541,N_24479,N_24977);
nand UO_542 (O_542,N_24601,N_24463);
xor UO_543 (O_543,N_24847,N_24315);
or UO_544 (O_544,N_23923,N_23975);
xor UO_545 (O_545,N_24317,N_24958);
nor UO_546 (O_546,N_24745,N_23829);
nand UO_547 (O_547,N_24648,N_24069);
nand UO_548 (O_548,N_23869,N_24200);
xor UO_549 (O_549,N_24821,N_24187);
nor UO_550 (O_550,N_24493,N_24809);
or UO_551 (O_551,N_24379,N_24951);
xnor UO_552 (O_552,N_24570,N_24488);
xor UO_553 (O_553,N_24421,N_24713);
nand UO_554 (O_554,N_23954,N_24095);
and UO_555 (O_555,N_24566,N_23856);
xor UO_556 (O_556,N_23906,N_23884);
xor UO_557 (O_557,N_24575,N_24756);
xor UO_558 (O_558,N_24752,N_23925);
xnor UO_559 (O_559,N_24917,N_24872);
nor UO_560 (O_560,N_23754,N_24014);
and UO_561 (O_561,N_24608,N_24446);
xnor UO_562 (O_562,N_24793,N_24047);
nand UO_563 (O_563,N_24646,N_24321);
nor UO_564 (O_564,N_24827,N_24299);
xor UO_565 (O_565,N_24714,N_23915);
nand UO_566 (O_566,N_24515,N_23947);
nand UO_567 (O_567,N_24710,N_24072);
nand UO_568 (O_568,N_24933,N_24703);
xnor UO_569 (O_569,N_24235,N_24474);
xor UO_570 (O_570,N_24829,N_24327);
or UO_571 (O_571,N_24101,N_23892);
nand UO_572 (O_572,N_23883,N_23983);
nand UO_573 (O_573,N_24104,N_23887);
or UO_574 (O_574,N_24624,N_24986);
or UO_575 (O_575,N_24467,N_23853);
or UO_576 (O_576,N_23823,N_24436);
nor UO_577 (O_577,N_23799,N_23924);
nor UO_578 (O_578,N_24589,N_24833);
and UO_579 (O_579,N_24222,N_23949);
nand UO_580 (O_580,N_24781,N_24052);
xnor UO_581 (O_581,N_24437,N_23991);
xnor UO_582 (O_582,N_24033,N_24402);
or UO_583 (O_583,N_24669,N_24911);
xnor UO_584 (O_584,N_24774,N_24098);
and UO_585 (O_585,N_24381,N_23785);
nand UO_586 (O_586,N_24538,N_24941);
xnor UO_587 (O_587,N_24932,N_23825);
and UO_588 (O_588,N_24484,N_24058);
or UO_589 (O_589,N_24050,N_24116);
nor UO_590 (O_590,N_24707,N_24596);
nor UO_591 (O_591,N_24708,N_24142);
and UO_592 (O_592,N_24051,N_24586);
xnor UO_593 (O_593,N_23894,N_24408);
and UO_594 (O_594,N_23790,N_24473);
nor UO_595 (O_595,N_23807,N_24962);
or UO_596 (O_596,N_24215,N_24114);
and UO_597 (O_597,N_24320,N_24066);
xnor UO_598 (O_598,N_24453,N_24661);
nand UO_599 (O_599,N_24388,N_23970);
xnor UO_600 (O_600,N_24303,N_24160);
and UO_601 (O_601,N_23926,N_24715);
nand UO_602 (O_602,N_24564,N_24587);
or UO_603 (O_603,N_24384,N_23945);
xor UO_604 (O_604,N_24766,N_24372);
and UO_605 (O_605,N_24549,N_24724);
or UO_606 (O_606,N_24422,N_24389);
and UO_607 (O_607,N_24519,N_24551);
or UO_608 (O_608,N_23955,N_24635);
nor UO_609 (O_609,N_24782,N_24106);
nor UO_610 (O_610,N_24914,N_24286);
nand UO_611 (O_611,N_24748,N_23890);
and UO_612 (O_612,N_24644,N_24403);
nor UO_613 (O_613,N_24939,N_24692);
xor UO_614 (O_614,N_24588,N_24345);
xnor UO_615 (O_615,N_24823,N_24178);
and UO_616 (O_616,N_24059,N_24373);
xor UO_617 (O_617,N_24189,N_24073);
nand UO_618 (O_618,N_24494,N_24263);
or UO_619 (O_619,N_24965,N_23805);
or UO_620 (O_620,N_24397,N_24577);
nor UO_621 (O_621,N_24181,N_24861);
nand UO_622 (O_622,N_23889,N_23793);
or UO_623 (O_623,N_24496,N_24324);
nor UO_624 (O_624,N_24358,N_24548);
or UO_625 (O_625,N_24452,N_23918);
nand UO_626 (O_626,N_24715,N_24738);
xor UO_627 (O_627,N_24224,N_24943);
nand UO_628 (O_628,N_23814,N_24356);
xor UO_629 (O_629,N_23919,N_24568);
and UO_630 (O_630,N_23795,N_24135);
xnor UO_631 (O_631,N_24728,N_23756);
xnor UO_632 (O_632,N_24729,N_24730);
nand UO_633 (O_633,N_24167,N_24263);
or UO_634 (O_634,N_24770,N_23836);
or UO_635 (O_635,N_24430,N_23760);
nor UO_636 (O_636,N_24640,N_24847);
nor UO_637 (O_637,N_24772,N_24988);
or UO_638 (O_638,N_24888,N_24580);
xnor UO_639 (O_639,N_24175,N_24580);
nand UO_640 (O_640,N_24914,N_23755);
xnor UO_641 (O_641,N_24674,N_24322);
xnor UO_642 (O_642,N_24145,N_24140);
or UO_643 (O_643,N_23851,N_24437);
nor UO_644 (O_644,N_24950,N_24952);
xor UO_645 (O_645,N_24671,N_23955);
and UO_646 (O_646,N_24255,N_23948);
xnor UO_647 (O_647,N_24869,N_24872);
and UO_648 (O_648,N_23905,N_24112);
and UO_649 (O_649,N_23985,N_24428);
or UO_650 (O_650,N_24869,N_24888);
nor UO_651 (O_651,N_24447,N_24755);
nand UO_652 (O_652,N_24488,N_24865);
nor UO_653 (O_653,N_24033,N_23974);
or UO_654 (O_654,N_24673,N_24905);
nor UO_655 (O_655,N_24409,N_24656);
xor UO_656 (O_656,N_24866,N_24165);
nor UO_657 (O_657,N_24114,N_24897);
xnor UO_658 (O_658,N_24267,N_24783);
and UO_659 (O_659,N_24350,N_24242);
xor UO_660 (O_660,N_23851,N_24761);
nand UO_661 (O_661,N_24861,N_24960);
or UO_662 (O_662,N_24226,N_24414);
xor UO_663 (O_663,N_24129,N_24291);
xor UO_664 (O_664,N_24100,N_24522);
and UO_665 (O_665,N_24587,N_24814);
nor UO_666 (O_666,N_23957,N_24164);
nor UO_667 (O_667,N_23970,N_24611);
and UO_668 (O_668,N_24993,N_23772);
and UO_669 (O_669,N_24480,N_24138);
or UO_670 (O_670,N_24515,N_23979);
or UO_671 (O_671,N_24576,N_24619);
nand UO_672 (O_672,N_24009,N_24538);
nand UO_673 (O_673,N_24976,N_24861);
nand UO_674 (O_674,N_24406,N_24373);
or UO_675 (O_675,N_24444,N_24552);
nand UO_676 (O_676,N_24625,N_24172);
nand UO_677 (O_677,N_24612,N_24667);
and UO_678 (O_678,N_24185,N_24699);
xor UO_679 (O_679,N_24643,N_24957);
and UO_680 (O_680,N_24820,N_23940);
or UO_681 (O_681,N_23888,N_24773);
or UO_682 (O_682,N_24644,N_24468);
nand UO_683 (O_683,N_24342,N_24336);
nand UO_684 (O_684,N_24082,N_24104);
nand UO_685 (O_685,N_24716,N_23850);
nor UO_686 (O_686,N_24630,N_24057);
xor UO_687 (O_687,N_24665,N_23763);
nor UO_688 (O_688,N_24909,N_24121);
nor UO_689 (O_689,N_24202,N_24889);
nor UO_690 (O_690,N_24528,N_24709);
and UO_691 (O_691,N_24273,N_24385);
nor UO_692 (O_692,N_24779,N_23895);
nor UO_693 (O_693,N_24202,N_24966);
nor UO_694 (O_694,N_24088,N_24892);
nor UO_695 (O_695,N_23866,N_24508);
and UO_696 (O_696,N_23974,N_24624);
nand UO_697 (O_697,N_23887,N_24789);
xor UO_698 (O_698,N_23885,N_24496);
xor UO_699 (O_699,N_24944,N_23951);
nand UO_700 (O_700,N_24897,N_24543);
nor UO_701 (O_701,N_24429,N_24790);
xor UO_702 (O_702,N_24917,N_24654);
xor UO_703 (O_703,N_24448,N_23946);
nand UO_704 (O_704,N_23874,N_24246);
and UO_705 (O_705,N_23824,N_24688);
nand UO_706 (O_706,N_24963,N_24787);
nand UO_707 (O_707,N_24382,N_24218);
nor UO_708 (O_708,N_24246,N_23787);
xnor UO_709 (O_709,N_24928,N_23974);
xnor UO_710 (O_710,N_24726,N_24801);
and UO_711 (O_711,N_24334,N_24806);
nand UO_712 (O_712,N_24741,N_24587);
nor UO_713 (O_713,N_24312,N_24137);
or UO_714 (O_714,N_24886,N_23792);
nor UO_715 (O_715,N_23969,N_23864);
and UO_716 (O_716,N_24896,N_23763);
nor UO_717 (O_717,N_24062,N_24792);
nor UO_718 (O_718,N_24834,N_23818);
or UO_719 (O_719,N_24266,N_24959);
xor UO_720 (O_720,N_24917,N_24011);
or UO_721 (O_721,N_24234,N_24696);
nand UO_722 (O_722,N_24452,N_24769);
nor UO_723 (O_723,N_24020,N_24191);
xor UO_724 (O_724,N_24396,N_24012);
xor UO_725 (O_725,N_24996,N_24151);
and UO_726 (O_726,N_23980,N_24665);
or UO_727 (O_727,N_24840,N_23930);
nor UO_728 (O_728,N_24451,N_24768);
xor UO_729 (O_729,N_24880,N_23779);
or UO_730 (O_730,N_23928,N_24983);
and UO_731 (O_731,N_24256,N_23802);
nor UO_732 (O_732,N_24521,N_24127);
nand UO_733 (O_733,N_23816,N_24642);
nand UO_734 (O_734,N_23851,N_24604);
nor UO_735 (O_735,N_24075,N_24643);
xor UO_736 (O_736,N_24462,N_24280);
nor UO_737 (O_737,N_23930,N_24941);
and UO_738 (O_738,N_24135,N_23810);
nand UO_739 (O_739,N_23907,N_23794);
nand UO_740 (O_740,N_24549,N_24540);
nor UO_741 (O_741,N_24152,N_23981);
nor UO_742 (O_742,N_24373,N_24804);
and UO_743 (O_743,N_24728,N_24691);
nand UO_744 (O_744,N_24306,N_24431);
xnor UO_745 (O_745,N_24543,N_24349);
or UO_746 (O_746,N_24400,N_24305);
nor UO_747 (O_747,N_24596,N_24362);
nand UO_748 (O_748,N_24823,N_24096);
nor UO_749 (O_749,N_24685,N_24809);
or UO_750 (O_750,N_23886,N_24383);
nor UO_751 (O_751,N_24794,N_24499);
and UO_752 (O_752,N_24409,N_24152);
nand UO_753 (O_753,N_24161,N_24760);
nor UO_754 (O_754,N_23763,N_23898);
and UO_755 (O_755,N_24146,N_24156);
or UO_756 (O_756,N_24330,N_24748);
nor UO_757 (O_757,N_24537,N_23897);
nand UO_758 (O_758,N_24632,N_24372);
and UO_759 (O_759,N_24352,N_24514);
xnor UO_760 (O_760,N_24968,N_24474);
or UO_761 (O_761,N_24270,N_24393);
or UO_762 (O_762,N_23952,N_24691);
or UO_763 (O_763,N_23834,N_24696);
xnor UO_764 (O_764,N_24753,N_24363);
and UO_765 (O_765,N_23756,N_24746);
and UO_766 (O_766,N_23898,N_24384);
nor UO_767 (O_767,N_23765,N_24484);
nand UO_768 (O_768,N_24096,N_24416);
or UO_769 (O_769,N_24881,N_23927);
xor UO_770 (O_770,N_24580,N_24893);
nand UO_771 (O_771,N_24940,N_23942);
and UO_772 (O_772,N_24282,N_23926);
xnor UO_773 (O_773,N_24209,N_24514);
or UO_774 (O_774,N_24409,N_24894);
nand UO_775 (O_775,N_24422,N_24037);
nor UO_776 (O_776,N_24848,N_23789);
nand UO_777 (O_777,N_23981,N_23914);
nor UO_778 (O_778,N_24738,N_24590);
nand UO_779 (O_779,N_23808,N_24330);
nor UO_780 (O_780,N_23791,N_23929);
xor UO_781 (O_781,N_24721,N_24962);
nor UO_782 (O_782,N_24049,N_24704);
and UO_783 (O_783,N_24139,N_24199);
or UO_784 (O_784,N_24503,N_24578);
nand UO_785 (O_785,N_23827,N_23901);
nor UO_786 (O_786,N_23889,N_24089);
nand UO_787 (O_787,N_24671,N_24872);
nor UO_788 (O_788,N_24130,N_24820);
nand UO_789 (O_789,N_24122,N_24088);
and UO_790 (O_790,N_24778,N_24953);
or UO_791 (O_791,N_24886,N_23946);
nand UO_792 (O_792,N_24133,N_24393);
xor UO_793 (O_793,N_24074,N_24647);
xnor UO_794 (O_794,N_24111,N_24673);
nand UO_795 (O_795,N_24837,N_24724);
xor UO_796 (O_796,N_24863,N_23915);
nor UO_797 (O_797,N_24650,N_23767);
or UO_798 (O_798,N_24488,N_24393);
nor UO_799 (O_799,N_24045,N_24937);
and UO_800 (O_800,N_23965,N_24326);
nor UO_801 (O_801,N_24780,N_24094);
xor UO_802 (O_802,N_24580,N_24435);
or UO_803 (O_803,N_24352,N_24966);
and UO_804 (O_804,N_24433,N_24606);
nand UO_805 (O_805,N_23989,N_23902);
and UO_806 (O_806,N_24574,N_24278);
and UO_807 (O_807,N_24448,N_23814);
xnor UO_808 (O_808,N_24848,N_24320);
nand UO_809 (O_809,N_24868,N_24417);
xor UO_810 (O_810,N_24642,N_24195);
or UO_811 (O_811,N_23957,N_23804);
nor UO_812 (O_812,N_24415,N_24525);
xnor UO_813 (O_813,N_23960,N_24565);
nand UO_814 (O_814,N_24531,N_24538);
nand UO_815 (O_815,N_24667,N_24752);
and UO_816 (O_816,N_24430,N_24157);
xnor UO_817 (O_817,N_24933,N_23901);
nor UO_818 (O_818,N_24687,N_23983);
or UO_819 (O_819,N_24439,N_24787);
xnor UO_820 (O_820,N_23889,N_23902);
and UO_821 (O_821,N_24371,N_24982);
and UO_822 (O_822,N_24825,N_24385);
xnor UO_823 (O_823,N_24831,N_23971);
or UO_824 (O_824,N_24166,N_24635);
nor UO_825 (O_825,N_24884,N_24612);
or UO_826 (O_826,N_24183,N_24273);
or UO_827 (O_827,N_24786,N_24683);
xor UO_828 (O_828,N_24854,N_24576);
nand UO_829 (O_829,N_24544,N_24804);
nand UO_830 (O_830,N_24541,N_24860);
nand UO_831 (O_831,N_24794,N_24873);
nor UO_832 (O_832,N_24623,N_23977);
nor UO_833 (O_833,N_23941,N_24554);
xor UO_834 (O_834,N_24094,N_24546);
nor UO_835 (O_835,N_24366,N_24973);
and UO_836 (O_836,N_23902,N_24730);
xnor UO_837 (O_837,N_24826,N_24092);
xor UO_838 (O_838,N_24040,N_24284);
xnor UO_839 (O_839,N_24358,N_24692);
nor UO_840 (O_840,N_24038,N_24194);
nor UO_841 (O_841,N_24368,N_24664);
and UO_842 (O_842,N_23955,N_24585);
or UO_843 (O_843,N_24078,N_24815);
xor UO_844 (O_844,N_23982,N_24831);
nor UO_845 (O_845,N_24201,N_24739);
or UO_846 (O_846,N_23846,N_24401);
nor UO_847 (O_847,N_24177,N_24161);
or UO_848 (O_848,N_24223,N_24957);
nand UO_849 (O_849,N_24096,N_24360);
xnor UO_850 (O_850,N_24497,N_24976);
and UO_851 (O_851,N_24402,N_24099);
nor UO_852 (O_852,N_24728,N_24276);
nand UO_853 (O_853,N_24480,N_24574);
xor UO_854 (O_854,N_24411,N_24117);
nor UO_855 (O_855,N_23904,N_24491);
nand UO_856 (O_856,N_24314,N_24872);
nor UO_857 (O_857,N_24198,N_24978);
nand UO_858 (O_858,N_24442,N_23788);
xor UO_859 (O_859,N_24986,N_24252);
and UO_860 (O_860,N_23753,N_24526);
nand UO_861 (O_861,N_23848,N_24003);
and UO_862 (O_862,N_24224,N_24978);
or UO_863 (O_863,N_24235,N_24478);
xnor UO_864 (O_864,N_24951,N_24651);
nor UO_865 (O_865,N_24737,N_24842);
nor UO_866 (O_866,N_24458,N_23801);
and UO_867 (O_867,N_23988,N_24158);
nor UO_868 (O_868,N_23938,N_24832);
nor UO_869 (O_869,N_24658,N_24145);
or UO_870 (O_870,N_24066,N_24371);
nor UO_871 (O_871,N_24151,N_24818);
and UO_872 (O_872,N_24867,N_24573);
nor UO_873 (O_873,N_24315,N_24186);
xnor UO_874 (O_874,N_24091,N_24086);
nor UO_875 (O_875,N_24037,N_23814);
nand UO_876 (O_876,N_24890,N_23933);
nor UO_877 (O_877,N_24424,N_23846);
xnor UO_878 (O_878,N_24238,N_24722);
and UO_879 (O_879,N_23824,N_23825);
or UO_880 (O_880,N_24686,N_24657);
nor UO_881 (O_881,N_24554,N_24477);
or UO_882 (O_882,N_24221,N_23839);
nor UO_883 (O_883,N_24630,N_24372);
nand UO_884 (O_884,N_24430,N_24754);
xnor UO_885 (O_885,N_24095,N_23995);
xnor UO_886 (O_886,N_23875,N_24022);
xor UO_887 (O_887,N_24149,N_24404);
and UO_888 (O_888,N_24321,N_24364);
or UO_889 (O_889,N_24242,N_24990);
nor UO_890 (O_890,N_24908,N_24423);
and UO_891 (O_891,N_24932,N_24990);
and UO_892 (O_892,N_24547,N_24404);
nand UO_893 (O_893,N_24461,N_24893);
nand UO_894 (O_894,N_24979,N_24545);
nand UO_895 (O_895,N_24645,N_24942);
or UO_896 (O_896,N_24029,N_24200);
and UO_897 (O_897,N_24686,N_24617);
nand UO_898 (O_898,N_24916,N_23874);
or UO_899 (O_899,N_24973,N_24505);
nor UO_900 (O_900,N_24252,N_24329);
nor UO_901 (O_901,N_24528,N_24367);
nor UO_902 (O_902,N_24223,N_24188);
or UO_903 (O_903,N_24404,N_24101);
and UO_904 (O_904,N_24610,N_24036);
nor UO_905 (O_905,N_24945,N_24536);
or UO_906 (O_906,N_24570,N_23888);
and UO_907 (O_907,N_24683,N_24500);
or UO_908 (O_908,N_23860,N_24095);
nand UO_909 (O_909,N_24983,N_24966);
nand UO_910 (O_910,N_24077,N_23865);
nor UO_911 (O_911,N_24685,N_24748);
and UO_912 (O_912,N_24228,N_24739);
xnor UO_913 (O_913,N_24409,N_23884);
or UO_914 (O_914,N_24241,N_24308);
or UO_915 (O_915,N_23790,N_24776);
nor UO_916 (O_916,N_24949,N_23878);
nor UO_917 (O_917,N_24032,N_24873);
xor UO_918 (O_918,N_24271,N_24701);
and UO_919 (O_919,N_24556,N_24651);
or UO_920 (O_920,N_24191,N_24444);
and UO_921 (O_921,N_24351,N_24141);
and UO_922 (O_922,N_23969,N_24403);
xor UO_923 (O_923,N_23970,N_24716);
nand UO_924 (O_924,N_24796,N_23995);
and UO_925 (O_925,N_24978,N_24254);
nand UO_926 (O_926,N_24169,N_23768);
or UO_927 (O_927,N_24220,N_24237);
xnor UO_928 (O_928,N_24475,N_23767);
or UO_929 (O_929,N_23951,N_24201);
nor UO_930 (O_930,N_24765,N_24118);
or UO_931 (O_931,N_24672,N_24131);
xnor UO_932 (O_932,N_24286,N_23920);
and UO_933 (O_933,N_24242,N_24315);
or UO_934 (O_934,N_24613,N_24747);
nand UO_935 (O_935,N_24869,N_24881);
nand UO_936 (O_936,N_24237,N_24649);
xnor UO_937 (O_937,N_23894,N_24582);
and UO_938 (O_938,N_24568,N_24265);
xnor UO_939 (O_939,N_24211,N_24667);
nand UO_940 (O_940,N_23982,N_24933);
xor UO_941 (O_941,N_24694,N_24659);
or UO_942 (O_942,N_23782,N_24307);
nand UO_943 (O_943,N_24833,N_24184);
nand UO_944 (O_944,N_24255,N_23888);
or UO_945 (O_945,N_23817,N_24414);
or UO_946 (O_946,N_24475,N_24476);
xor UO_947 (O_947,N_24614,N_24481);
or UO_948 (O_948,N_24274,N_24062);
and UO_949 (O_949,N_24250,N_24276);
xnor UO_950 (O_950,N_23992,N_24545);
nor UO_951 (O_951,N_24545,N_23837);
or UO_952 (O_952,N_23758,N_24426);
xor UO_953 (O_953,N_24935,N_24786);
nor UO_954 (O_954,N_24343,N_24016);
or UO_955 (O_955,N_24385,N_24412);
nor UO_956 (O_956,N_24578,N_24661);
and UO_957 (O_957,N_24145,N_24921);
nand UO_958 (O_958,N_24086,N_24886);
and UO_959 (O_959,N_23784,N_24891);
nand UO_960 (O_960,N_23997,N_23889);
nand UO_961 (O_961,N_24876,N_24647);
nor UO_962 (O_962,N_23937,N_23946);
xor UO_963 (O_963,N_23780,N_23841);
xor UO_964 (O_964,N_24367,N_23862);
or UO_965 (O_965,N_24439,N_24788);
xnor UO_966 (O_966,N_23954,N_24085);
xor UO_967 (O_967,N_24211,N_23785);
and UO_968 (O_968,N_24079,N_24439);
nand UO_969 (O_969,N_24007,N_23799);
nand UO_970 (O_970,N_24898,N_24590);
xor UO_971 (O_971,N_23964,N_24136);
nor UO_972 (O_972,N_24562,N_23811);
or UO_973 (O_973,N_23993,N_24139);
nor UO_974 (O_974,N_24501,N_24630);
nand UO_975 (O_975,N_24289,N_24930);
nand UO_976 (O_976,N_24210,N_23810);
or UO_977 (O_977,N_24268,N_24662);
xor UO_978 (O_978,N_24832,N_24572);
xnor UO_979 (O_979,N_24629,N_24206);
nor UO_980 (O_980,N_23972,N_24178);
and UO_981 (O_981,N_23836,N_23843);
nand UO_982 (O_982,N_24599,N_23963);
nor UO_983 (O_983,N_24393,N_24542);
nor UO_984 (O_984,N_24704,N_24351);
nand UO_985 (O_985,N_24260,N_24776);
nor UO_986 (O_986,N_24884,N_24279);
or UO_987 (O_987,N_24603,N_24183);
xnor UO_988 (O_988,N_24607,N_24688);
and UO_989 (O_989,N_23770,N_24854);
nor UO_990 (O_990,N_24976,N_23967);
nand UO_991 (O_991,N_23906,N_24426);
or UO_992 (O_992,N_24204,N_23853);
xnor UO_993 (O_993,N_24646,N_24909);
nor UO_994 (O_994,N_23975,N_23964);
nand UO_995 (O_995,N_24634,N_24382);
xor UO_996 (O_996,N_23786,N_24608);
nand UO_997 (O_997,N_24044,N_24535);
nor UO_998 (O_998,N_24672,N_24425);
and UO_999 (O_999,N_24470,N_24458);
nor UO_1000 (O_1000,N_23919,N_24159);
xor UO_1001 (O_1001,N_24986,N_24044);
and UO_1002 (O_1002,N_23754,N_24827);
or UO_1003 (O_1003,N_23843,N_23887);
and UO_1004 (O_1004,N_23804,N_24575);
and UO_1005 (O_1005,N_24557,N_24368);
xor UO_1006 (O_1006,N_24911,N_24316);
and UO_1007 (O_1007,N_24631,N_24957);
nor UO_1008 (O_1008,N_24490,N_23828);
nand UO_1009 (O_1009,N_24809,N_24633);
or UO_1010 (O_1010,N_24005,N_24277);
and UO_1011 (O_1011,N_24126,N_24213);
and UO_1012 (O_1012,N_23928,N_24080);
xor UO_1013 (O_1013,N_24698,N_24352);
xor UO_1014 (O_1014,N_24321,N_24356);
nand UO_1015 (O_1015,N_24259,N_23918);
xnor UO_1016 (O_1016,N_24162,N_23865);
or UO_1017 (O_1017,N_24607,N_24561);
or UO_1018 (O_1018,N_24009,N_24362);
or UO_1019 (O_1019,N_24743,N_24311);
nor UO_1020 (O_1020,N_24747,N_23951);
nand UO_1021 (O_1021,N_23829,N_24634);
nor UO_1022 (O_1022,N_24835,N_24282);
nand UO_1023 (O_1023,N_24766,N_24516);
or UO_1024 (O_1024,N_24320,N_24394);
and UO_1025 (O_1025,N_24040,N_23795);
and UO_1026 (O_1026,N_24175,N_24522);
nand UO_1027 (O_1027,N_24202,N_24206);
or UO_1028 (O_1028,N_24352,N_24757);
and UO_1029 (O_1029,N_23786,N_24386);
and UO_1030 (O_1030,N_24309,N_23779);
xor UO_1031 (O_1031,N_23992,N_24423);
nand UO_1032 (O_1032,N_24391,N_24734);
nor UO_1033 (O_1033,N_24566,N_23788);
or UO_1034 (O_1034,N_23916,N_24967);
xnor UO_1035 (O_1035,N_24567,N_24122);
nand UO_1036 (O_1036,N_24354,N_24814);
nand UO_1037 (O_1037,N_24461,N_24066);
nor UO_1038 (O_1038,N_24934,N_24863);
nand UO_1039 (O_1039,N_24246,N_24624);
or UO_1040 (O_1040,N_24978,N_23804);
and UO_1041 (O_1041,N_24027,N_23850);
xor UO_1042 (O_1042,N_23957,N_24852);
nor UO_1043 (O_1043,N_24484,N_24101);
nor UO_1044 (O_1044,N_24223,N_24422);
and UO_1045 (O_1045,N_23901,N_24055);
or UO_1046 (O_1046,N_24728,N_24752);
and UO_1047 (O_1047,N_24585,N_24734);
nand UO_1048 (O_1048,N_24661,N_24187);
xor UO_1049 (O_1049,N_23915,N_24448);
or UO_1050 (O_1050,N_24050,N_24990);
nor UO_1051 (O_1051,N_23874,N_24954);
and UO_1052 (O_1052,N_24139,N_24011);
nand UO_1053 (O_1053,N_24122,N_24249);
or UO_1054 (O_1054,N_24427,N_24693);
nand UO_1055 (O_1055,N_23897,N_24874);
nor UO_1056 (O_1056,N_23857,N_24534);
nand UO_1057 (O_1057,N_24790,N_24356);
xor UO_1058 (O_1058,N_24136,N_24823);
and UO_1059 (O_1059,N_23857,N_24850);
nor UO_1060 (O_1060,N_23795,N_24963);
nand UO_1061 (O_1061,N_23781,N_24570);
and UO_1062 (O_1062,N_24297,N_24666);
and UO_1063 (O_1063,N_24874,N_24360);
and UO_1064 (O_1064,N_24524,N_23985);
nand UO_1065 (O_1065,N_24666,N_23842);
nand UO_1066 (O_1066,N_24509,N_23774);
or UO_1067 (O_1067,N_24094,N_24018);
and UO_1068 (O_1068,N_24126,N_24186);
nand UO_1069 (O_1069,N_24207,N_24104);
nand UO_1070 (O_1070,N_24653,N_24243);
and UO_1071 (O_1071,N_24436,N_24741);
or UO_1072 (O_1072,N_24668,N_24227);
and UO_1073 (O_1073,N_24868,N_24088);
xor UO_1074 (O_1074,N_24691,N_24640);
and UO_1075 (O_1075,N_23875,N_24403);
or UO_1076 (O_1076,N_24449,N_24616);
nand UO_1077 (O_1077,N_24538,N_24723);
xnor UO_1078 (O_1078,N_24785,N_24937);
nor UO_1079 (O_1079,N_23856,N_23809);
nor UO_1080 (O_1080,N_24038,N_23893);
nor UO_1081 (O_1081,N_24473,N_24261);
nor UO_1082 (O_1082,N_23798,N_24486);
nor UO_1083 (O_1083,N_24747,N_24720);
or UO_1084 (O_1084,N_24690,N_24943);
and UO_1085 (O_1085,N_24452,N_24043);
and UO_1086 (O_1086,N_24684,N_24635);
nor UO_1087 (O_1087,N_24705,N_24265);
nand UO_1088 (O_1088,N_24035,N_23961);
and UO_1089 (O_1089,N_24337,N_24964);
or UO_1090 (O_1090,N_24669,N_24684);
nor UO_1091 (O_1091,N_23881,N_24393);
or UO_1092 (O_1092,N_24680,N_23942);
or UO_1093 (O_1093,N_24111,N_24295);
and UO_1094 (O_1094,N_24455,N_24202);
or UO_1095 (O_1095,N_24043,N_24723);
and UO_1096 (O_1096,N_24338,N_23765);
nand UO_1097 (O_1097,N_24337,N_24433);
nor UO_1098 (O_1098,N_24912,N_24631);
nand UO_1099 (O_1099,N_24079,N_24573);
and UO_1100 (O_1100,N_24521,N_24254);
nand UO_1101 (O_1101,N_24324,N_24292);
xnor UO_1102 (O_1102,N_24706,N_24482);
nand UO_1103 (O_1103,N_24376,N_24200);
nor UO_1104 (O_1104,N_24070,N_24235);
xnor UO_1105 (O_1105,N_24264,N_24904);
nand UO_1106 (O_1106,N_23898,N_23843);
and UO_1107 (O_1107,N_23971,N_24891);
xor UO_1108 (O_1108,N_24783,N_24440);
nor UO_1109 (O_1109,N_24693,N_24635);
nor UO_1110 (O_1110,N_24688,N_24417);
or UO_1111 (O_1111,N_24282,N_24296);
nor UO_1112 (O_1112,N_24175,N_24653);
xor UO_1113 (O_1113,N_24773,N_23755);
nand UO_1114 (O_1114,N_23909,N_23884);
nand UO_1115 (O_1115,N_24900,N_24398);
nor UO_1116 (O_1116,N_24358,N_24967);
and UO_1117 (O_1117,N_24854,N_24418);
xnor UO_1118 (O_1118,N_24827,N_24468);
or UO_1119 (O_1119,N_24326,N_23754);
nor UO_1120 (O_1120,N_24860,N_24165);
xor UO_1121 (O_1121,N_24271,N_24830);
nand UO_1122 (O_1122,N_23756,N_23887);
nor UO_1123 (O_1123,N_24086,N_24737);
nand UO_1124 (O_1124,N_24172,N_24340);
nand UO_1125 (O_1125,N_24115,N_24531);
nor UO_1126 (O_1126,N_24897,N_23834);
nand UO_1127 (O_1127,N_24743,N_24317);
nor UO_1128 (O_1128,N_24116,N_24121);
nand UO_1129 (O_1129,N_23841,N_24901);
nor UO_1130 (O_1130,N_24960,N_24638);
and UO_1131 (O_1131,N_23837,N_24084);
and UO_1132 (O_1132,N_24961,N_23841);
nand UO_1133 (O_1133,N_24030,N_23944);
nor UO_1134 (O_1134,N_24366,N_24872);
nor UO_1135 (O_1135,N_24211,N_24492);
nor UO_1136 (O_1136,N_24238,N_24015);
and UO_1137 (O_1137,N_23916,N_24461);
nor UO_1138 (O_1138,N_24697,N_24395);
and UO_1139 (O_1139,N_24801,N_24567);
xnor UO_1140 (O_1140,N_24267,N_24518);
or UO_1141 (O_1141,N_24212,N_24474);
or UO_1142 (O_1142,N_24130,N_24711);
or UO_1143 (O_1143,N_23915,N_24240);
xor UO_1144 (O_1144,N_24509,N_24759);
and UO_1145 (O_1145,N_24429,N_24275);
and UO_1146 (O_1146,N_24036,N_23968);
or UO_1147 (O_1147,N_23883,N_24098);
or UO_1148 (O_1148,N_24403,N_24320);
nand UO_1149 (O_1149,N_24570,N_24117);
xor UO_1150 (O_1150,N_24646,N_23925);
or UO_1151 (O_1151,N_24319,N_24368);
or UO_1152 (O_1152,N_24859,N_23830);
xnor UO_1153 (O_1153,N_24046,N_24057);
or UO_1154 (O_1154,N_24541,N_23975);
nand UO_1155 (O_1155,N_23832,N_24477);
nand UO_1156 (O_1156,N_24804,N_24888);
and UO_1157 (O_1157,N_24478,N_24643);
nor UO_1158 (O_1158,N_24662,N_24980);
and UO_1159 (O_1159,N_24600,N_23949);
xnor UO_1160 (O_1160,N_24332,N_24155);
nand UO_1161 (O_1161,N_23988,N_24856);
xnor UO_1162 (O_1162,N_23819,N_23785);
nor UO_1163 (O_1163,N_24326,N_24165);
or UO_1164 (O_1164,N_24131,N_24712);
nor UO_1165 (O_1165,N_24060,N_24977);
nor UO_1166 (O_1166,N_24088,N_24657);
nand UO_1167 (O_1167,N_23917,N_23768);
or UO_1168 (O_1168,N_24692,N_24864);
nand UO_1169 (O_1169,N_23819,N_24754);
nand UO_1170 (O_1170,N_24613,N_24644);
nor UO_1171 (O_1171,N_23837,N_24391);
xnor UO_1172 (O_1172,N_24992,N_24911);
nor UO_1173 (O_1173,N_24047,N_24652);
or UO_1174 (O_1174,N_24588,N_24911);
nand UO_1175 (O_1175,N_23800,N_24753);
or UO_1176 (O_1176,N_24799,N_24738);
xor UO_1177 (O_1177,N_24174,N_24107);
or UO_1178 (O_1178,N_24481,N_24440);
or UO_1179 (O_1179,N_23925,N_24774);
and UO_1180 (O_1180,N_24663,N_24748);
or UO_1181 (O_1181,N_24520,N_23763);
nand UO_1182 (O_1182,N_24877,N_24095);
and UO_1183 (O_1183,N_24940,N_24612);
nor UO_1184 (O_1184,N_23853,N_24992);
nor UO_1185 (O_1185,N_23924,N_23937);
xnor UO_1186 (O_1186,N_24570,N_24182);
and UO_1187 (O_1187,N_24185,N_23772);
nand UO_1188 (O_1188,N_24232,N_24245);
xnor UO_1189 (O_1189,N_24541,N_24167);
nand UO_1190 (O_1190,N_24461,N_23753);
xor UO_1191 (O_1191,N_24693,N_24273);
and UO_1192 (O_1192,N_24148,N_24319);
or UO_1193 (O_1193,N_23899,N_24463);
and UO_1194 (O_1194,N_24268,N_24081);
or UO_1195 (O_1195,N_24677,N_24366);
nand UO_1196 (O_1196,N_24787,N_24256);
nor UO_1197 (O_1197,N_24607,N_24657);
xor UO_1198 (O_1198,N_24971,N_24459);
nand UO_1199 (O_1199,N_24878,N_24229);
nand UO_1200 (O_1200,N_24003,N_23800);
or UO_1201 (O_1201,N_24836,N_23975);
nor UO_1202 (O_1202,N_24820,N_24623);
nand UO_1203 (O_1203,N_24161,N_24055);
nand UO_1204 (O_1204,N_24087,N_24447);
xnor UO_1205 (O_1205,N_24628,N_24242);
nor UO_1206 (O_1206,N_24414,N_23924);
or UO_1207 (O_1207,N_24926,N_24592);
or UO_1208 (O_1208,N_24990,N_24913);
nand UO_1209 (O_1209,N_24975,N_23861);
xnor UO_1210 (O_1210,N_23835,N_24695);
nand UO_1211 (O_1211,N_23780,N_24186);
or UO_1212 (O_1212,N_23911,N_23957);
xor UO_1213 (O_1213,N_24092,N_24993);
nor UO_1214 (O_1214,N_24587,N_24305);
nor UO_1215 (O_1215,N_24270,N_24825);
xor UO_1216 (O_1216,N_24164,N_24659);
or UO_1217 (O_1217,N_24506,N_24008);
nand UO_1218 (O_1218,N_23952,N_23780);
xor UO_1219 (O_1219,N_24135,N_24990);
xor UO_1220 (O_1220,N_24392,N_24143);
nor UO_1221 (O_1221,N_24016,N_24273);
or UO_1222 (O_1222,N_24533,N_23971);
and UO_1223 (O_1223,N_24606,N_24797);
nor UO_1224 (O_1224,N_24376,N_24931);
nor UO_1225 (O_1225,N_24147,N_24305);
and UO_1226 (O_1226,N_24552,N_23974);
and UO_1227 (O_1227,N_23960,N_24492);
xor UO_1228 (O_1228,N_23982,N_23852);
nand UO_1229 (O_1229,N_24525,N_24986);
nand UO_1230 (O_1230,N_24976,N_24826);
and UO_1231 (O_1231,N_23809,N_24197);
nand UO_1232 (O_1232,N_24853,N_23951);
nor UO_1233 (O_1233,N_24389,N_24011);
and UO_1234 (O_1234,N_24027,N_24664);
and UO_1235 (O_1235,N_24295,N_24326);
nor UO_1236 (O_1236,N_24244,N_24808);
xor UO_1237 (O_1237,N_24416,N_24135);
nand UO_1238 (O_1238,N_24681,N_24641);
xor UO_1239 (O_1239,N_24015,N_24468);
nor UO_1240 (O_1240,N_23883,N_24280);
nand UO_1241 (O_1241,N_24653,N_24676);
nand UO_1242 (O_1242,N_24689,N_24650);
or UO_1243 (O_1243,N_24446,N_24195);
or UO_1244 (O_1244,N_24639,N_24619);
nand UO_1245 (O_1245,N_24908,N_24824);
xor UO_1246 (O_1246,N_24399,N_24032);
and UO_1247 (O_1247,N_24825,N_23948);
and UO_1248 (O_1248,N_23767,N_24823);
and UO_1249 (O_1249,N_24961,N_24641);
nor UO_1250 (O_1250,N_24595,N_24580);
xnor UO_1251 (O_1251,N_24238,N_23773);
xor UO_1252 (O_1252,N_24726,N_24927);
nand UO_1253 (O_1253,N_23809,N_24064);
nor UO_1254 (O_1254,N_24561,N_24579);
and UO_1255 (O_1255,N_24694,N_24734);
xnor UO_1256 (O_1256,N_24925,N_24955);
nand UO_1257 (O_1257,N_23993,N_24158);
xnor UO_1258 (O_1258,N_24178,N_24166);
and UO_1259 (O_1259,N_24581,N_24897);
or UO_1260 (O_1260,N_24021,N_24713);
xnor UO_1261 (O_1261,N_24739,N_24056);
nor UO_1262 (O_1262,N_24007,N_24382);
nand UO_1263 (O_1263,N_24410,N_24656);
nor UO_1264 (O_1264,N_24717,N_24847);
nand UO_1265 (O_1265,N_24925,N_24742);
or UO_1266 (O_1266,N_23893,N_24304);
nor UO_1267 (O_1267,N_24043,N_24927);
nand UO_1268 (O_1268,N_24560,N_23766);
xor UO_1269 (O_1269,N_24078,N_23902);
xnor UO_1270 (O_1270,N_24908,N_23881);
or UO_1271 (O_1271,N_24266,N_24352);
or UO_1272 (O_1272,N_24602,N_24370);
nand UO_1273 (O_1273,N_24734,N_24559);
xnor UO_1274 (O_1274,N_24187,N_24445);
nor UO_1275 (O_1275,N_24335,N_24623);
nor UO_1276 (O_1276,N_23962,N_24967);
nand UO_1277 (O_1277,N_24403,N_24794);
or UO_1278 (O_1278,N_24917,N_24878);
nand UO_1279 (O_1279,N_24760,N_24112);
nor UO_1280 (O_1280,N_23757,N_24107);
nand UO_1281 (O_1281,N_23924,N_23988);
xnor UO_1282 (O_1282,N_24568,N_24582);
or UO_1283 (O_1283,N_24490,N_24328);
nand UO_1284 (O_1284,N_24613,N_24614);
nand UO_1285 (O_1285,N_24940,N_23997);
nor UO_1286 (O_1286,N_24102,N_24624);
nor UO_1287 (O_1287,N_24059,N_24891);
nand UO_1288 (O_1288,N_24883,N_24100);
and UO_1289 (O_1289,N_24531,N_24145);
and UO_1290 (O_1290,N_23760,N_23885);
or UO_1291 (O_1291,N_24346,N_24119);
or UO_1292 (O_1292,N_24059,N_23765);
nor UO_1293 (O_1293,N_24221,N_24619);
nor UO_1294 (O_1294,N_24109,N_23872);
or UO_1295 (O_1295,N_24290,N_24361);
nor UO_1296 (O_1296,N_24570,N_23790);
or UO_1297 (O_1297,N_24354,N_24418);
and UO_1298 (O_1298,N_24472,N_24616);
and UO_1299 (O_1299,N_24053,N_24583);
nand UO_1300 (O_1300,N_24304,N_24859);
and UO_1301 (O_1301,N_24932,N_24216);
and UO_1302 (O_1302,N_23894,N_24910);
and UO_1303 (O_1303,N_24486,N_24089);
or UO_1304 (O_1304,N_24700,N_24799);
or UO_1305 (O_1305,N_24915,N_24186);
nand UO_1306 (O_1306,N_24849,N_24358);
or UO_1307 (O_1307,N_24011,N_24464);
xnor UO_1308 (O_1308,N_24048,N_24719);
xnor UO_1309 (O_1309,N_24077,N_24994);
xnor UO_1310 (O_1310,N_24855,N_24503);
and UO_1311 (O_1311,N_24323,N_24416);
xnor UO_1312 (O_1312,N_24564,N_24238);
nor UO_1313 (O_1313,N_24493,N_24183);
xor UO_1314 (O_1314,N_23767,N_24692);
or UO_1315 (O_1315,N_24267,N_24665);
or UO_1316 (O_1316,N_24938,N_24826);
nor UO_1317 (O_1317,N_23944,N_23906);
or UO_1318 (O_1318,N_24364,N_23959);
xnor UO_1319 (O_1319,N_24325,N_24956);
nand UO_1320 (O_1320,N_24185,N_24638);
xor UO_1321 (O_1321,N_24454,N_24985);
and UO_1322 (O_1322,N_23848,N_24176);
nand UO_1323 (O_1323,N_24726,N_24021);
nand UO_1324 (O_1324,N_23815,N_24826);
or UO_1325 (O_1325,N_24252,N_23829);
nand UO_1326 (O_1326,N_24409,N_24141);
nor UO_1327 (O_1327,N_24369,N_24506);
nand UO_1328 (O_1328,N_24048,N_24291);
nand UO_1329 (O_1329,N_23908,N_24484);
and UO_1330 (O_1330,N_24250,N_24665);
and UO_1331 (O_1331,N_23825,N_23897);
or UO_1332 (O_1332,N_23967,N_24736);
and UO_1333 (O_1333,N_24725,N_24548);
xnor UO_1334 (O_1334,N_24754,N_24455);
nand UO_1335 (O_1335,N_24480,N_24651);
nor UO_1336 (O_1336,N_23905,N_24815);
or UO_1337 (O_1337,N_24919,N_23895);
nand UO_1338 (O_1338,N_24254,N_24582);
nor UO_1339 (O_1339,N_23878,N_24368);
and UO_1340 (O_1340,N_23964,N_24279);
and UO_1341 (O_1341,N_23758,N_23900);
nor UO_1342 (O_1342,N_24755,N_24860);
nor UO_1343 (O_1343,N_24884,N_24485);
nor UO_1344 (O_1344,N_23869,N_24286);
or UO_1345 (O_1345,N_24971,N_24045);
xor UO_1346 (O_1346,N_24213,N_24828);
xor UO_1347 (O_1347,N_24974,N_23880);
xnor UO_1348 (O_1348,N_24786,N_24687);
or UO_1349 (O_1349,N_23966,N_23861);
nor UO_1350 (O_1350,N_24172,N_24497);
nor UO_1351 (O_1351,N_24649,N_24642);
and UO_1352 (O_1352,N_24803,N_24902);
and UO_1353 (O_1353,N_24970,N_24729);
xnor UO_1354 (O_1354,N_23765,N_24078);
nand UO_1355 (O_1355,N_24537,N_24244);
nand UO_1356 (O_1356,N_24184,N_24228);
or UO_1357 (O_1357,N_23845,N_24662);
or UO_1358 (O_1358,N_24918,N_24592);
nand UO_1359 (O_1359,N_24040,N_24016);
or UO_1360 (O_1360,N_24846,N_24358);
xnor UO_1361 (O_1361,N_23829,N_24334);
xor UO_1362 (O_1362,N_24775,N_24357);
or UO_1363 (O_1363,N_24410,N_24980);
xnor UO_1364 (O_1364,N_24095,N_24368);
xnor UO_1365 (O_1365,N_24731,N_24359);
nor UO_1366 (O_1366,N_24568,N_24483);
nor UO_1367 (O_1367,N_23825,N_24964);
and UO_1368 (O_1368,N_24583,N_24389);
or UO_1369 (O_1369,N_24395,N_23774);
and UO_1370 (O_1370,N_23757,N_23960);
and UO_1371 (O_1371,N_24906,N_24327);
nor UO_1372 (O_1372,N_23786,N_24722);
nand UO_1373 (O_1373,N_24393,N_23923);
or UO_1374 (O_1374,N_24595,N_24527);
xor UO_1375 (O_1375,N_24843,N_24543);
nand UO_1376 (O_1376,N_24621,N_24472);
and UO_1377 (O_1377,N_24184,N_23838);
and UO_1378 (O_1378,N_24512,N_24783);
nand UO_1379 (O_1379,N_24992,N_24262);
nor UO_1380 (O_1380,N_23794,N_24547);
or UO_1381 (O_1381,N_24199,N_23871);
or UO_1382 (O_1382,N_24012,N_24094);
xnor UO_1383 (O_1383,N_24774,N_24020);
nand UO_1384 (O_1384,N_23759,N_23842);
nor UO_1385 (O_1385,N_24276,N_24806);
nor UO_1386 (O_1386,N_24043,N_24699);
xor UO_1387 (O_1387,N_24992,N_24663);
xor UO_1388 (O_1388,N_24225,N_24400);
or UO_1389 (O_1389,N_24225,N_24565);
xnor UO_1390 (O_1390,N_24866,N_24682);
nand UO_1391 (O_1391,N_24755,N_24849);
nor UO_1392 (O_1392,N_23986,N_24482);
nor UO_1393 (O_1393,N_24800,N_24300);
or UO_1394 (O_1394,N_24737,N_24800);
or UO_1395 (O_1395,N_24877,N_24944);
and UO_1396 (O_1396,N_24156,N_24819);
nor UO_1397 (O_1397,N_24622,N_24964);
nand UO_1398 (O_1398,N_23776,N_24290);
xor UO_1399 (O_1399,N_24757,N_24538);
or UO_1400 (O_1400,N_24950,N_24368);
and UO_1401 (O_1401,N_24014,N_24926);
or UO_1402 (O_1402,N_24404,N_24006);
xor UO_1403 (O_1403,N_24918,N_24949);
and UO_1404 (O_1404,N_24513,N_24070);
nor UO_1405 (O_1405,N_24733,N_24775);
or UO_1406 (O_1406,N_24902,N_24467);
and UO_1407 (O_1407,N_24972,N_24889);
or UO_1408 (O_1408,N_24557,N_24006);
nor UO_1409 (O_1409,N_24813,N_23919);
nor UO_1410 (O_1410,N_24580,N_24098);
nor UO_1411 (O_1411,N_23792,N_24598);
xor UO_1412 (O_1412,N_24642,N_24003);
and UO_1413 (O_1413,N_24976,N_24431);
or UO_1414 (O_1414,N_24103,N_23798);
nor UO_1415 (O_1415,N_23776,N_23837);
xnor UO_1416 (O_1416,N_24923,N_23948);
or UO_1417 (O_1417,N_24858,N_24068);
xnor UO_1418 (O_1418,N_24846,N_24543);
xor UO_1419 (O_1419,N_24453,N_24570);
or UO_1420 (O_1420,N_23987,N_23998);
nand UO_1421 (O_1421,N_24348,N_23832);
and UO_1422 (O_1422,N_24930,N_24724);
or UO_1423 (O_1423,N_24439,N_24507);
or UO_1424 (O_1424,N_24191,N_24539);
and UO_1425 (O_1425,N_24132,N_24748);
or UO_1426 (O_1426,N_24193,N_24880);
nor UO_1427 (O_1427,N_23902,N_23993);
nor UO_1428 (O_1428,N_24822,N_24152);
nand UO_1429 (O_1429,N_24876,N_24596);
nand UO_1430 (O_1430,N_24556,N_23923);
xor UO_1431 (O_1431,N_24362,N_24819);
or UO_1432 (O_1432,N_23925,N_24134);
and UO_1433 (O_1433,N_24007,N_24351);
or UO_1434 (O_1434,N_23756,N_24952);
nor UO_1435 (O_1435,N_24191,N_24123);
nor UO_1436 (O_1436,N_24931,N_23834);
nand UO_1437 (O_1437,N_24166,N_24391);
and UO_1438 (O_1438,N_24378,N_24474);
or UO_1439 (O_1439,N_24433,N_23926);
and UO_1440 (O_1440,N_23827,N_24285);
xnor UO_1441 (O_1441,N_24020,N_24751);
xnor UO_1442 (O_1442,N_24796,N_24310);
nor UO_1443 (O_1443,N_24608,N_24438);
xnor UO_1444 (O_1444,N_24049,N_24955);
or UO_1445 (O_1445,N_24014,N_24523);
and UO_1446 (O_1446,N_23811,N_24986);
nand UO_1447 (O_1447,N_23917,N_23853);
or UO_1448 (O_1448,N_24847,N_24689);
nand UO_1449 (O_1449,N_24484,N_24439);
and UO_1450 (O_1450,N_24656,N_23791);
nor UO_1451 (O_1451,N_24467,N_24236);
and UO_1452 (O_1452,N_24063,N_23974);
and UO_1453 (O_1453,N_24683,N_24197);
xor UO_1454 (O_1454,N_24876,N_24122);
and UO_1455 (O_1455,N_24639,N_24012);
or UO_1456 (O_1456,N_24844,N_24927);
nor UO_1457 (O_1457,N_24262,N_24122);
nor UO_1458 (O_1458,N_24068,N_23941);
nand UO_1459 (O_1459,N_24127,N_24022);
and UO_1460 (O_1460,N_24218,N_23845);
nor UO_1461 (O_1461,N_24549,N_23875);
or UO_1462 (O_1462,N_24295,N_24296);
xor UO_1463 (O_1463,N_23847,N_24466);
xnor UO_1464 (O_1464,N_24576,N_24385);
nor UO_1465 (O_1465,N_24792,N_24694);
nand UO_1466 (O_1466,N_23817,N_24122);
nor UO_1467 (O_1467,N_23947,N_24625);
nand UO_1468 (O_1468,N_23755,N_24547);
xnor UO_1469 (O_1469,N_24818,N_24789);
and UO_1470 (O_1470,N_24124,N_24821);
nor UO_1471 (O_1471,N_24104,N_24782);
nand UO_1472 (O_1472,N_23790,N_24454);
xor UO_1473 (O_1473,N_24074,N_24950);
nor UO_1474 (O_1474,N_23962,N_24414);
or UO_1475 (O_1475,N_24853,N_24708);
nor UO_1476 (O_1476,N_24464,N_23801);
and UO_1477 (O_1477,N_24900,N_24254);
nor UO_1478 (O_1478,N_24199,N_24483);
and UO_1479 (O_1479,N_23888,N_24820);
or UO_1480 (O_1480,N_24744,N_24750);
or UO_1481 (O_1481,N_24577,N_23888);
xor UO_1482 (O_1482,N_23816,N_24731);
nand UO_1483 (O_1483,N_24952,N_23998);
nand UO_1484 (O_1484,N_24289,N_24792);
xor UO_1485 (O_1485,N_24382,N_23834);
or UO_1486 (O_1486,N_24607,N_24042);
or UO_1487 (O_1487,N_23843,N_24183);
nor UO_1488 (O_1488,N_24418,N_24410);
xnor UO_1489 (O_1489,N_23814,N_24360);
and UO_1490 (O_1490,N_24362,N_24050);
and UO_1491 (O_1491,N_24802,N_24398);
nor UO_1492 (O_1492,N_24582,N_24290);
nand UO_1493 (O_1493,N_24432,N_24421);
or UO_1494 (O_1494,N_24071,N_24970);
xnor UO_1495 (O_1495,N_24536,N_24781);
xor UO_1496 (O_1496,N_24037,N_24770);
xor UO_1497 (O_1497,N_24362,N_24538);
xor UO_1498 (O_1498,N_24102,N_23867);
and UO_1499 (O_1499,N_24244,N_24770);
nand UO_1500 (O_1500,N_24246,N_23922);
nor UO_1501 (O_1501,N_23770,N_24004);
xor UO_1502 (O_1502,N_23932,N_24384);
and UO_1503 (O_1503,N_23989,N_24831);
xnor UO_1504 (O_1504,N_24160,N_24759);
nor UO_1505 (O_1505,N_24598,N_24752);
or UO_1506 (O_1506,N_24810,N_24920);
nand UO_1507 (O_1507,N_24047,N_23950);
nand UO_1508 (O_1508,N_24471,N_24434);
xor UO_1509 (O_1509,N_24052,N_24841);
and UO_1510 (O_1510,N_24254,N_24605);
nand UO_1511 (O_1511,N_24998,N_24405);
nand UO_1512 (O_1512,N_24238,N_24162);
and UO_1513 (O_1513,N_24382,N_24968);
xor UO_1514 (O_1514,N_24066,N_24885);
and UO_1515 (O_1515,N_24998,N_24421);
and UO_1516 (O_1516,N_23916,N_24593);
nand UO_1517 (O_1517,N_24046,N_24570);
nor UO_1518 (O_1518,N_24453,N_24827);
or UO_1519 (O_1519,N_24118,N_24490);
and UO_1520 (O_1520,N_24892,N_24334);
nand UO_1521 (O_1521,N_24877,N_23959);
and UO_1522 (O_1522,N_24423,N_24429);
or UO_1523 (O_1523,N_24840,N_23914);
or UO_1524 (O_1524,N_23796,N_23973);
xnor UO_1525 (O_1525,N_24144,N_23881);
and UO_1526 (O_1526,N_24381,N_24439);
or UO_1527 (O_1527,N_24051,N_24213);
and UO_1528 (O_1528,N_23846,N_23826);
nand UO_1529 (O_1529,N_24357,N_24617);
and UO_1530 (O_1530,N_24110,N_24301);
and UO_1531 (O_1531,N_24370,N_24354);
nor UO_1532 (O_1532,N_23770,N_24715);
nor UO_1533 (O_1533,N_23994,N_24671);
nor UO_1534 (O_1534,N_24712,N_24597);
xor UO_1535 (O_1535,N_24004,N_24199);
xor UO_1536 (O_1536,N_23960,N_23967);
xnor UO_1537 (O_1537,N_23844,N_24632);
nand UO_1538 (O_1538,N_23915,N_24618);
xor UO_1539 (O_1539,N_24035,N_24158);
nand UO_1540 (O_1540,N_23756,N_23993);
nor UO_1541 (O_1541,N_23996,N_24187);
or UO_1542 (O_1542,N_24107,N_24462);
and UO_1543 (O_1543,N_24016,N_24252);
nor UO_1544 (O_1544,N_24444,N_24592);
nand UO_1545 (O_1545,N_24387,N_24710);
nor UO_1546 (O_1546,N_24991,N_23927);
and UO_1547 (O_1547,N_24126,N_23792);
or UO_1548 (O_1548,N_24139,N_24935);
or UO_1549 (O_1549,N_24617,N_24597);
and UO_1550 (O_1550,N_24262,N_24164);
nor UO_1551 (O_1551,N_24028,N_24969);
nand UO_1552 (O_1552,N_24452,N_24986);
xor UO_1553 (O_1553,N_24938,N_24062);
or UO_1554 (O_1554,N_24472,N_24267);
nand UO_1555 (O_1555,N_24404,N_24668);
xnor UO_1556 (O_1556,N_24536,N_24828);
nand UO_1557 (O_1557,N_23789,N_24325);
nand UO_1558 (O_1558,N_24423,N_24147);
nor UO_1559 (O_1559,N_24805,N_23793);
nand UO_1560 (O_1560,N_24094,N_24387);
nand UO_1561 (O_1561,N_24314,N_24139);
and UO_1562 (O_1562,N_24508,N_24699);
xor UO_1563 (O_1563,N_24454,N_23819);
nor UO_1564 (O_1564,N_24506,N_24540);
and UO_1565 (O_1565,N_23892,N_24184);
nor UO_1566 (O_1566,N_24517,N_24952);
and UO_1567 (O_1567,N_23839,N_23828);
xnor UO_1568 (O_1568,N_24485,N_24555);
nand UO_1569 (O_1569,N_24856,N_24562);
xor UO_1570 (O_1570,N_24026,N_24304);
and UO_1571 (O_1571,N_24960,N_23949);
nand UO_1572 (O_1572,N_24559,N_24372);
or UO_1573 (O_1573,N_24460,N_24719);
nor UO_1574 (O_1574,N_24884,N_24158);
or UO_1575 (O_1575,N_24396,N_24398);
and UO_1576 (O_1576,N_24926,N_24972);
or UO_1577 (O_1577,N_24450,N_24114);
and UO_1578 (O_1578,N_23868,N_24961);
and UO_1579 (O_1579,N_24025,N_24328);
xor UO_1580 (O_1580,N_24433,N_24199);
nor UO_1581 (O_1581,N_23788,N_23809);
xor UO_1582 (O_1582,N_24449,N_24744);
and UO_1583 (O_1583,N_24388,N_23968);
nor UO_1584 (O_1584,N_24919,N_24003);
or UO_1585 (O_1585,N_24804,N_24083);
xor UO_1586 (O_1586,N_23829,N_24688);
or UO_1587 (O_1587,N_24333,N_24976);
or UO_1588 (O_1588,N_24861,N_24228);
xor UO_1589 (O_1589,N_24779,N_24752);
xnor UO_1590 (O_1590,N_24548,N_23988);
xnor UO_1591 (O_1591,N_24928,N_24377);
nand UO_1592 (O_1592,N_24142,N_24383);
or UO_1593 (O_1593,N_24693,N_24028);
and UO_1594 (O_1594,N_24758,N_24279);
xnor UO_1595 (O_1595,N_24710,N_23805);
and UO_1596 (O_1596,N_24949,N_24160);
and UO_1597 (O_1597,N_24174,N_24382);
xnor UO_1598 (O_1598,N_24245,N_24444);
nor UO_1599 (O_1599,N_24721,N_24082);
xor UO_1600 (O_1600,N_24003,N_23964);
nor UO_1601 (O_1601,N_24364,N_23901);
nand UO_1602 (O_1602,N_24040,N_24918);
or UO_1603 (O_1603,N_24492,N_24738);
or UO_1604 (O_1604,N_24053,N_23999);
xor UO_1605 (O_1605,N_24159,N_24178);
and UO_1606 (O_1606,N_24754,N_24236);
nor UO_1607 (O_1607,N_24827,N_24444);
xor UO_1608 (O_1608,N_24010,N_24616);
nand UO_1609 (O_1609,N_24574,N_24089);
and UO_1610 (O_1610,N_24255,N_24152);
nand UO_1611 (O_1611,N_24327,N_24608);
and UO_1612 (O_1612,N_24922,N_24444);
or UO_1613 (O_1613,N_24842,N_24503);
and UO_1614 (O_1614,N_24634,N_24606);
or UO_1615 (O_1615,N_24564,N_23817);
nor UO_1616 (O_1616,N_24541,N_23753);
nand UO_1617 (O_1617,N_24715,N_24515);
xor UO_1618 (O_1618,N_24527,N_24882);
nor UO_1619 (O_1619,N_24750,N_23756);
nand UO_1620 (O_1620,N_24340,N_24761);
and UO_1621 (O_1621,N_24773,N_24720);
nor UO_1622 (O_1622,N_24232,N_24683);
and UO_1623 (O_1623,N_23940,N_24279);
nand UO_1624 (O_1624,N_24646,N_23887);
and UO_1625 (O_1625,N_24635,N_24227);
nor UO_1626 (O_1626,N_23967,N_23979);
xnor UO_1627 (O_1627,N_23889,N_24680);
or UO_1628 (O_1628,N_24657,N_24393);
or UO_1629 (O_1629,N_24734,N_23950);
xnor UO_1630 (O_1630,N_24490,N_23838);
and UO_1631 (O_1631,N_24940,N_24909);
or UO_1632 (O_1632,N_24182,N_24222);
xnor UO_1633 (O_1633,N_24619,N_24944);
xnor UO_1634 (O_1634,N_24709,N_23968);
xor UO_1635 (O_1635,N_24599,N_23826);
or UO_1636 (O_1636,N_24492,N_24510);
xor UO_1637 (O_1637,N_24477,N_24344);
xnor UO_1638 (O_1638,N_24679,N_24526);
nor UO_1639 (O_1639,N_24519,N_23996);
or UO_1640 (O_1640,N_24956,N_23803);
nand UO_1641 (O_1641,N_24584,N_24601);
and UO_1642 (O_1642,N_24302,N_24289);
and UO_1643 (O_1643,N_23950,N_24427);
or UO_1644 (O_1644,N_24796,N_24776);
nor UO_1645 (O_1645,N_24103,N_23805);
and UO_1646 (O_1646,N_24694,N_24579);
or UO_1647 (O_1647,N_24644,N_24413);
nand UO_1648 (O_1648,N_24227,N_24066);
nand UO_1649 (O_1649,N_24384,N_23950);
and UO_1650 (O_1650,N_24437,N_23956);
xnor UO_1651 (O_1651,N_24679,N_24263);
and UO_1652 (O_1652,N_24353,N_24460);
and UO_1653 (O_1653,N_23771,N_23798);
xor UO_1654 (O_1654,N_24956,N_24252);
or UO_1655 (O_1655,N_24397,N_24508);
xor UO_1656 (O_1656,N_24324,N_24286);
nand UO_1657 (O_1657,N_24966,N_23822);
nand UO_1658 (O_1658,N_24142,N_24561);
and UO_1659 (O_1659,N_23780,N_24893);
nand UO_1660 (O_1660,N_24869,N_24311);
xor UO_1661 (O_1661,N_24887,N_23777);
nor UO_1662 (O_1662,N_24603,N_24120);
or UO_1663 (O_1663,N_24438,N_24895);
nor UO_1664 (O_1664,N_24252,N_24276);
nor UO_1665 (O_1665,N_24494,N_24637);
and UO_1666 (O_1666,N_24360,N_23971);
nand UO_1667 (O_1667,N_24960,N_24722);
and UO_1668 (O_1668,N_24016,N_24302);
or UO_1669 (O_1669,N_23853,N_24871);
nand UO_1670 (O_1670,N_24360,N_23772);
and UO_1671 (O_1671,N_24847,N_24385);
or UO_1672 (O_1672,N_24226,N_24948);
nor UO_1673 (O_1673,N_24092,N_24140);
xnor UO_1674 (O_1674,N_24960,N_24944);
and UO_1675 (O_1675,N_24248,N_24205);
nand UO_1676 (O_1676,N_23825,N_24075);
nor UO_1677 (O_1677,N_24698,N_24733);
nand UO_1678 (O_1678,N_24992,N_24277);
and UO_1679 (O_1679,N_24123,N_23920);
nand UO_1680 (O_1680,N_24157,N_23943);
nor UO_1681 (O_1681,N_24113,N_23953);
nand UO_1682 (O_1682,N_24026,N_24610);
nor UO_1683 (O_1683,N_24980,N_23754);
and UO_1684 (O_1684,N_24549,N_24396);
nand UO_1685 (O_1685,N_23867,N_24158);
or UO_1686 (O_1686,N_24388,N_24842);
xnor UO_1687 (O_1687,N_24676,N_24652);
and UO_1688 (O_1688,N_24404,N_24224);
xor UO_1689 (O_1689,N_23949,N_23923);
nand UO_1690 (O_1690,N_24576,N_23868);
or UO_1691 (O_1691,N_23854,N_24814);
and UO_1692 (O_1692,N_24326,N_24168);
and UO_1693 (O_1693,N_24955,N_24151);
and UO_1694 (O_1694,N_24699,N_23853);
nand UO_1695 (O_1695,N_23972,N_24332);
nor UO_1696 (O_1696,N_23800,N_24650);
xor UO_1697 (O_1697,N_24220,N_23998);
and UO_1698 (O_1698,N_24494,N_24026);
nand UO_1699 (O_1699,N_24405,N_24821);
xor UO_1700 (O_1700,N_24071,N_24385);
and UO_1701 (O_1701,N_24598,N_24537);
xnor UO_1702 (O_1702,N_24318,N_24107);
or UO_1703 (O_1703,N_24886,N_24151);
xor UO_1704 (O_1704,N_24515,N_24258);
xor UO_1705 (O_1705,N_24995,N_24663);
nand UO_1706 (O_1706,N_24404,N_24664);
xnor UO_1707 (O_1707,N_24921,N_24219);
nand UO_1708 (O_1708,N_24426,N_24582);
nand UO_1709 (O_1709,N_24996,N_24323);
nand UO_1710 (O_1710,N_24951,N_24322);
nor UO_1711 (O_1711,N_24147,N_23820);
xnor UO_1712 (O_1712,N_24455,N_24606);
or UO_1713 (O_1713,N_24813,N_23941);
nor UO_1714 (O_1714,N_24388,N_24726);
nand UO_1715 (O_1715,N_24996,N_24452);
and UO_1716 (O_1716,N_23772,N_23986);
and UO_1717 (O_1717,N_24774,N_24891);
nand UO_1718 (O_1718,N_24247,N_23775);
nand UO_1719 (O_1719,N_24886,N_24282);
nand UO_1720 (O_1720,N_23944,N_24388);
nor UO_1721 (O_1721,N_24916,N_24275);
xnor UO_1722 (O_1722,N_24268,N_24287);
and UO_1723 (O_1723,N_24065,N_24849);
nor UO_1724 (O_1724,N_24528,N_24202);
nor UO_1725 (O_1725,N_24352,N_23869);
or UO_1726 (O_1726,N_24376,N_23789);
or UO_1727 (O_1727,N_24841,N_24074);
and UO_1728 (O_1728,N_24164,N_23831);
nor UO_1729 (O_1729,N_24506,N_23841);
nor UO_1730 (O_1730,N_24527,N_23862);
xnor UO_1731 (O_1731,N_24478,N_23967);
xor UO_1732 (O_1732,N_23802,N_24825);
nor UO_1733 (O_1733,N_24496,N_24162);
xnor UO_1734 (O_1734,N_24683,N_24953);
or UO_1735 (O_1735,N_24311,N_24972);
or UO_1736 (O_1736,N_23866,N_23853);
or UO_1737 (O_1737,N_24243,N_24841);
and UO_1738 (O_1738,N_24015,N_24064);
and UO_1739 (O_1739,N_24378,N_24976);
nand UO_1740 (O_1740,N_24880,N_24609);
and UO_1741 (O_1741,N_24517,N_23836);
or UO_1742 (O_1742,N_24732,N_24635);
or UO_1743 (O_1743,N_24068,N_24330);
nand UO_1744 (O_1744,N_24525,N_23974);
or UO_1745 (O_1745,N_24330,N_24056);
or UO_1746 (O_1746,N_24093,N_24446);
and UO_1747 (O_1747,N_24685,N_24910);
nand UO_1748 (O_1748,N_24675,N_23763);
or UO_1749 (O_1749,N_24007,N_24554);
nor UO_1750 (O_1750,N_24963,N_23810);
xor UO_1751 (O_1751,N_24093,N_24507);
xor UO_1752 (O_1752,N_24058,N_23828);
or UO_1753 (O_1753,N_24679,N_23881);
xor UO_1754 (O_1754,N_24023,N_24204);
nand UO_1755 (O_1755,N_24525,N_24455);
and UO_1756 (O_1756,N_23879,N_24170);
xor UO_1757 (O_1757,N_23882,N_24168);
and UO_1758 (O_1758,N_23991,N_24832);
and UO_1759 (O_1759,N_24499,N_24459);
and UO_1760 (O_1760,N_23907,N_24463);
or UO_1761 (O_1761,N_24536,N_24038);
xor UO_1762 (O_1762,N_24236,N_24126);
and UO_1763 (O_1763,N_24539,N_23914);
nor UO_1764 (O_1764,N_23770,N_24738);
and UO_1765 (O_1765,N_24066,N_24204);
or UO_1766 (O_1766,N_24028,N_24425);
xnor UO_1767 (O_1767,N_24859,N_24911);
or UO_1768 (O_1768,N_23793,N_24571);
nand UO_1769 (O_1769,N_24067,N_24786);
or UO_1770 (O_1770,N_24306,N_24721);
xnor UO_1771 (O_1771,N_24550,N_24509);
or UO_1772 (O_1772,N_24807,N_24325);
and UO_1773 (O_1773,N_24326,N_24851);
xnor UO_1774 (O_1774,N_24463,N_24393);
nand UO_1775 (O_1775,N_24625,N_24446);
or UO_1776 (O_1776,N_24100,N_24041);
xor UO_1777 (O_1777,N_24391,N_24566);
nand UO_1778 (O_1778,N_24899,N_24379);
nand UO_1779 (O_1779,N_24818,N_24083);
and UO_1780 (O_1780,N_24013,N_24774);
xor UO_1781 (O_1781,N_24756,N_24844);
xnor UO_1782 (O_1782,N_24641,N_24231);
xnor UO_1783 (O_1783,N_24813,N_23822);
or UO_1784 (O_1784,N_24312,N_23950);
nor UO_1785 (O_1785,N_24864,N_24859);
nor UO_1786 (O_1786,N_24558,N_24514);
xnor UO_1787 (O_1787,N_24425,N_23999);
nor UO_1788 (O_1788,N_24204,N_24587);
xor UO_1789 (O_1789,N_24007,N_23928);
nand UO_1790 (O_1790,N_23801,N_23968);
nor UO_1791 (O_1791,N_24501,N_24785);
xnor UO_1792 (O_1792,N_23933,N_23909);
and UO_1793 (O_1793,N_23868,N_24119);
and UO_1794 (O_1794,N_23939,N_24030);
and UO_1795 (O_1795,N_24767,N_24967);
nor UO_1796 (O_1796,N_24066,N_24525);
or UO_1797 (O_1797,N_23978,N_24782);
nand UO_1798 (O_1798,N_24933,N_24063);
nand UO_1799 (O_1799,N_24132,N_24454);
or UO_1800 (O_1800,N_24625,N_23776);
nor UO_1801 (O_1801,N_24130,N_24324);
nand UO_1802 (O_1802,N_24615,N_24871);
or UO_1803 (O_1803,N_23756,N_24127);
or UO_1804 (O_1804,N_23918,N_23762);
nand UO_1805 (O_1805,N_24852,N_23859);
nor UO_1806 (O_1806,N_24702,N_23923);
and UO_1807 (O_1807,N_24968,N_24343);
or UO_1808 (O_1808,N_24708,N_24132);
or UO_1809 (O_1809,N_24843,N_24000);
nand UO_1810 (O_1810,N_24753,N_24923);
nor UO_1811 (O_1811,N_24631,N_24078);
nand UO_1812 (O_1812,N_24870,N_24124);
nand UO_1813 (O_1813,N_24381,N_23887);
or UO_1814 (O_1814,N_24064,N_24182);
nand UO_1815 (O_1815,N_24967,N_24421);
nand UO_1816 (O_1816,N_24370,N_24078);
and UO_1817 (O_1817,N_24505,N_23928);
xnor UO_1818 (O_1818,N_24784,N_23956);
nand UO_1819 (O_1819,N_24452,N_24263);
or UO_1820 (O_1820,N_24302,N_24172);
nor UO_1821 (O_1821,N_23997,N_24454);
xor UO_1822 (O_1822,N_24836,N_23871);
and UO_1823 (O_1823,N_24304,N_24789);
and UO_1824 (O_1824,N_24347,N_24284);
nor UO_1825 (O_1825,N_24463,N_24638);
and UO_1826 (O_1826,N_24938,N_24209);
and UO_1827 (O_1827,N_23964,N_24362);
or UO_1828 (O_1828,N_23812,N_24423);
xor UO_1829 (O_1829,N_24161,N_24814);
nand UO_1830 (O_1830,N_24567,N_24633);
xor UO_1831 (O_1831,N_24502,N_24528);
nand UO_1832 (O_1832,N_24656,N_24899);
nor UO_1833 (O_1833,N_24360,N_24104);
nand UO_1834 (O_1834,N_23841,N_24918);
and UO_1835 (O_1835,N_24030,N_24624);
nand UO_1836 (O_1836,N_24842,N_24716);
nand UO_1837 (O_1837,N_24340,N_24230);
nand UO_1838 (O_1838,N_24054,N_24213);
or UO_1839 (O_1839,N_24244,N_24627);
nor UO_1840 (O_1840,N_24795,N_23827);
and UO_1841 (O_1841,N_24714,N_23874);
and UO_1842 (O_1842,N_24457,N_24697);
nand UO_1843 (O_1843,N_24232,N_24765);
xnor UO_1844 (O_1844,N_24571,N_24556);
xor UO_1845 (O_1845,N_24721,N_23838);
xnor UO_1846 (O_1846,N_23939,N_24655);
xor UO_1847 (O_1847,N_24864,N_23911);
or UO_1848 (O_1848,N_24049,N_24432);
nor UO_1849 (O_1849,N_24624,N_24011);
xor UO_1850 (O_1850,N_24663,N_24556);
or UO_1851 (O_1851,N_24508,N_23918);
nand UO_1852 (O_1852,N_24122,N_24133);
xor UO_1853 (O_1853,N_23969,N_24969);
or UO_1854 (O_1854,N_24091,N_24184);
and UO_1855 (O_1855,N_24073,N_24075);
xnor UO_1856 (O_1856,N_24551,N_24532);
and UO_1857 (O_1857,N_24738,N_24682);
or UO_1858 (O_1858,N_23879,N_24588);
and UO_1859 (O_1859,N_24298,N_24369);
nor UO_1860 (O_1860,N_23901,N_24691);
nand UO_1861 (O_1861,N_24408,N_23985);
nand UO_1862 (O_1862,N_24747,N_23882);
nand UO_1863 (O_1863,N_24844,N_24303);
nor UO_1864 (O_1864,N_24907,N_23960);
nand UO_1865 (O_1865,N_24177,N_24526);
and UO_1866 (O_1866,N_24211,N_24114);
or UO_1867 (O_1867,N_23971,N_23801);
nand UO_1868 (O_1868,N_24422,N_24284);
or UO_1869 (O_1869,N_24493,N_24430);
nand UO_1870 (O_1870,N_24250,N_24606);
xor UO_1871 (O_1871,N_24461,N_24729);
and UO_1872 (O_1872,N_23839,N_23918);
and UO_1873 (O_1873,N_24370,N_24192);
nor UO_1874 (O_1874,N_24287,N_24829);
nor UO_1875 (O_1875,N_24706,N_23974);
and UO_1876 (O_1876,N_24667,N_24161);
xnor UO_1877 (O_1877,N_24653,N_24114);
or UO_1878 (O_1878,N_24373,N_24403);
xor UO_1879 (O_1879,N_23868,N_24572);
nand UO_1880 (O_1880,N_24564,N_24546);
nand UO_1881 (O_1881,N_24299,N_24124);
nand UO_1882 (O_1882,N_24319,N_24271);
and UO_1883 (O_1883,N_24077,N_24331);
xor UO_1884 (O_1884,N_24497,N_23833);
nor UO_1885 (O_1885,N_24372,N_23872);
nor UO_1886 (O_1886,N_24510,N_24958);
or UO_1887 (O_1887,N_24300,N_23751);
nand UO_1888 (O_1888,N_24773,N_24548);
xnor UO_1889 (O_1889,N_24582,N_24217);
nand UO_1890 (O_1890,N_24675,N_24293);
and UO_1891 (O_1891,N_24044,N_24010);
nor UO_1892 (O_1892,N_23831,N_24017);
and UO_1893 (O_1893,N_24956,N_24781);
nand UO_1894 (O_1894,N_23799,N_24372);
xnor UO_1895 (O_1895,N_24127,N_24992);
xnor UO_1896 (O_1896,N_24061,N_24263);
nand UO_1897 (O_1897,N_24086,N_24433);
xor UO_1898 (O_1898,N_24097,N_24022);
and UO_1899 (O_1899,N_24039,N_23849);
nand UO_1900 (O_1900,N_24998,N_24799);
xnor UO_1901 (O_1901,N_24098,N_24466);
xnor UO_1902 (O_1902,N_24369,N_24663);
or UO_1903 (O_1903,N_24299,N_24436);
xnor UO_1904 (O_1904,N_23796,N_24208);
nand UO_1905 (O_1905,N_24242,N_24635);
xor UO_1906 (O_1906,N_23777,N_23791);
nor UO_1907 (O_1907,N_23859,N_24297);
nor UO_1908 (O_1908,N_24850,N_24443);
nand UO_1909 (O_1909,N_23984,N_24738);
xor UO_1910 (O_1910,N_24634,N_23899);
nor UO_1911 (O_1911,N_23765,N_24340);
nand UO_1912 (O_1912,N_24043,N_24071);
and UO_1913 (O_1913,N_23818,N_24216);
nand UO_1914 (O_1914,N_24148,N_23815);
nor UO_1915 (O_1915,N_24835,N_23950);
nand UO_1916 (O_1916,N_24284,N_24673);
or UO_1917 (O_1917,N_24922,N_24979);
and UO_1918 (O_1918,N_24633,N_24916);
and UO_1919 (O_1919,N_24902,N_23968);
xnor UO_1920 (O_1920,N_24080,N_24297);
nand UO_1921 (O_1921,N_24892,N_24953);
nor UO_1922 (O_1922,N_24204,N_24222);
and UO_1923 (O_1923,N_24797,N_24607);
xnor UO_1924 (O_1924,N_24289,N_23933);
and UO_1925 (O_1925,N_24884,N_24347);
nor UO_1926 (O_1926,N_24393,N_24155);
xnor UO_1927 (O_1927,N_24899,N_24663);
or UO_1928 (O_1928,N_24159,N_24903);
or UO_1929 (O_1929,N_24701,N_24194);
nand UO_1930 (O_1930,N_24394,N_24438);
xor UO_1931 (O_1931,N_24939,N_24608);
xor UO_1932 (O_1932,N_24316,N_23875);
xnor UO_1933 (O_1933,N_24952,N_24688);
nand UO_1934 (O_1934,N_24892,N_23835);
or UO_1935 (O_1935,N_24408,N_24815);
xor UO_1936 (O_1936,N_24128,N_23833);
nand UO_1937 (O_1937,N_24629,N_24356);
or UO_1938 (O_1938,N_24820,N_24200);
and UO_1939 (O_1939,N_24155,N_24423);
nor UO_1940 (O_1940,N_24369,N_24659);
or UO_1941 (O_1941,N_24149,N_24491);
xor UO_1942 (O_1942,N_24552,N_24096);
xor UO_1943 (O_1943,N_24510,N_23985);
and UO_1944 (O_1944,N_24771,N_24323);
xnor UO_1945 (O_1945,N_24262,N_24771);
nor UO_1946 (O_1946,N_24889,N_24876);
nor UO_1947 (O_1947,N_24947,N_24109);
xor UO_1948 (O_1948,N_24984,N_23912);
nor UO_1949 (O_1949,N_24041,N_24628);
nor UO_1950 (O_1950,N_24775,N_24811);
or UO_1951 (O_1951,N_24901,N_24192);
or UO_1952 (O_1952,N_24093,N_24975);
or UO_1953 (O_1953,N_24954,N_24947);
nand UO_1954 (O_1954,N_24746,N_23954);
or UO_1955 (O_1955,N_24048,N_24457);
nand UO_1956 (O_1956,N_24056,N_24859);
or UO_1957 (O_1957,N_23816,N_24419);
nor UO_1958 (O_1958,N_23858,N_24363);
nand UO_1959 (O_1959,N_24771,N_24009);
or UO_1960 (O_1960,N_24084,N_24519);
nand UO_1961 (O_1961,N_24408,N_24590);
nand UO_1962 (O_1962,N_23755,N_24502);
and UO_1963 (O_1963,N_23985,N_23773);
or UO_1964 (O_1964,N_24152,N_24486);
and UO_1965 (O_1965,N_24862,N_23828);
nor UO_1966 (O_1966,N_24023,N_24515);
xor UO_1967 (O_1967,N_24885,N_24860);
nand UO_1968 (O_1968,N_24561,N_24328);
xnor UO_1969 (O_1969,N_24401,N_24673);
nor UO_1970 (O_1970,N_24971,N_24589);
nand UO_1971 (O_1971,N_24213,N_23812);
nor UO_1972 (O_1972,N_24044,N_24518);
nor UO_1973 (O_1973,N_24134,N_24157);
xor UO_1974 (O_1974,N_24212,N_24407);
or UO_1975 (O_1975,N_24524,N_24791);
or UO_1976 (O_1976,N_24812,N_24289);
and UO_1977 (O_1977,N_24502,N_24678);
or UO_1978 (O_1978,N_24942,N_24179);
nor UO_1979 (O_1979,N_24324,N_24727);
xor UO_1980 (O_1980,N_24712,N_24076);
and UO_1981 (O_1981,N_23948,N_23890);
nand UO_1982 (O_1982,N_24208,N_24993);
and UO_1983 (O_1983,N_23758,N_24003);
xor UO_1984 (O_1984,N_24722,N_23966);
or UO_1985 (O_1985,N_24965,N_24456);
or UO_1986 (O_1986,N_24933,N_24065);
and UO_1987 (O_1987,N_24316,N_24116);
nor UO_1988 (O_1988,N_24539,N_24374);
xnor UO_1989 (O_1989,N_24754,N_23996);
and UO_1990 (O_1990,N_24521,N_24954);
or UO_1991 (O_1991,N_24123,N_24968);
and UO_1992 (O_1992,N_24206,N_23919);
nor UO_1993 (O_1993,N_24622,N_23925);
and UO_1994 (O_1994,N_24520,N_23947);
and UO_1995 (O_1995,N_24878,N_24223);
and UO_1996 (O_1996,N_24489,N_23992);
nor UO_1997 (O_1997,N_23759,N_24602);
and UO_1998 (O_1998,N_24898,N_24511);
xor UO_1999 (O_1999,N_24246,N_24836);
xor UO_2000 (O_2000,N_24377,N_24869);
nor UO_2001 (O_2001,N_24704,N_24413);
or UO_2002 (O_2002,N_24365,N_24366);
or UO_2003 (O_2003,N_24208,N_23942);
nor UO_2004 (O_2004,N_23766,N_24333);
xor UO_2005 (O_2005,N_23816,N_24124);
or UO_2006 (O_2006,N_24816,N_24005);
xor UO_2007 (O_2007,N_24312,N_24157);
or UO_2008 (O_2008,N_24968,N_23907);
xor UO_2009 (O_2009,N_24750,N_23952);
nand UO_2010 (O_2010,N_23956,N_24259);
or UO_2011 (O_2011,N_23915,N_24701);
nand UO_2012 (O_2012,N_24563,N_24181);
nand UO_2013 (O_2013,N_24579,N_23905);
or UO_2014 (O_2014,N_24117,N_23918);
xnor UO_2015 (O_2015,N_24859,N_24550);
xnor UO_2016 (O_2016,N_24343,N_24634);
and UO_2017 (O_2017,N_24338,N_23766);
nor UO_2018 (O_2018,N_24042,N_24755);
and UO_2019 (O_2019,N_24050,N_24062);
xor UO_2020 (O_2020,N_24319,N_24870);
nand UO_2021 (O_2021,N_24768,N_24064);
xor UO_2022 (O_2022,N_23908,N_24329);
xnor UO_2023 (O_2023,N_23786,N_24869);
xnor UO_2024 (O_2024,N_24797,N_24636);
nand UO_2025 (O_2025,N_24953,N_24805);
and UO_2026 (O_2026,N_24274,N_23795);
nand UO_2027 (O_2027,N_24511,N_24838);
xnor UO_2028 (O_2028,N_24991,N_24672);
xor UO_2029 (O_2029,N_24989,N_23988);
or UO_2030 (O_2030,N_24773,N_24663);
or UO_2031 (O_2031,N_24756,N_24607);
and UO_2032 (O_2032,N_24946,N_23759);
xor UO_2033 (O_2033,N_24233,N_24830);
or UO_2034 (O_2034,N_23815,N_24614);
xnor UO_2035 (O_2035,N_24509,N_24092);
xor UO_2036 (O_2036,N_24924,N_24923);
nor UO_2037 (O_2037,N_24053,N_23814);
and UO_2038 (O_2038,N_24195,N_24962);
nor UO_2039 (O_2039,N_23999,N_24815);
or UO_2040 (O_2040,N_24008,N_24132);
nor UO_2041 (O_2041,N_24765,N_24855);
xor UO_2042 (O_2042,N_24755,N_24781);
xnor UO_2043 (O_2043,N_24091,N_24841);
xor UO_2044 (O_2044,N_24068,N_24849);
and UO_2045 (O_2045,N_23775,N_24272);
xor UO_2046 (O_2046,N_24194,N_24354);
and UO_2047 (O_2047,N_23893,N_24746);
or UO_2048 (O_2048,N_23870,N_23802);
nor UO_2049 (O_2049,N_24482,N_24483);
nor UO_2050 (O_2050,N_23750,N_23944);
and UO_2051 (O_2051,N_24479,N_24557);
or UO_2052 (O_2052,N_24883,N_24674);
xor UO_2053 (O_2053,N_24745,N_23949);
nand UO_2054 (O_2054,N_24035,N_24302);
nand UO_2055 (O_2055,N_24992,N_24129);
nand UO_2056 (O_2056,N_24801,N_24991);
or UO_2057 (O_2057,N_24739,N_24271);
or UO_2058 (O_2058,N_24267,N_24778);
and UO_2059 (O_2059,N_24422,N_24983);
nor UO_2060 (O_2060,N_24420,N_24238);
nand UO_2061 (O_2061,N_24361,N_24895);
nand UO_2062 (O_2062,N_24071,N_23862);
nand UO_2063 (O_2063,N_24698,N_23778);
nor UO_2064 (O_2064,N_23838,N_24809);
nand UO_2065 (O_2065,N_24498,N_24659);
xnor UO_2066 (O_2066,N_24723,N_24195);
xnor UO_2067 (O_2067,N_24663,N_23839);
or UO_2068 (O_2068,N_24164,N_24868);
or UO_2069 (O_2069,N_24789,N_24690);
and UO_2070 (O_2070,N_24850,N_24885);
nor UO_2071 (O_2071,N_24084,N_24347);
nand UO_2072 (O_2072,N_24614,N_24366);
xnor UO_2073 (O_2073,N_24780,N_24946);
nor UO_2074 (O_2074,N_24648,N_23901);
or UO_2075 (O_2075,N_24638,N_24759);
or UO_2076 (O_2076,N_23777,N_24076);
nor UO_2077 (O_2077,N_23896,N_24822);
nor UO_2078 (O_2078,N_24140,N_24224);
nand UO_2079 (O_2079,N_24625,N_24677);
xnor UO_2080 (O_2080,N_24204,N_24038);
nand UO_2081 (O_2081,N_23915,N_24900);
and UO_2082 (O_2082,N_23761,N_24290);
xnor UO_2083 (O_2083,N_24124,N_24082);
or UO_2084 (O_2084,N_24754,N_24551);
nor UO_2085 (O_2085,N_23831,N_24876);
nand UO_2086 (O_2086,N_24651,N_23953);
or UO_2087 (O_2087,N_23763,N_24102);
xor UO_2088 (O_2088,N_24278,N_24199);
and UO_2089 (O_2089,N_24918,N_24773);
or UO_2090 (O_2090,N_23951,N_24627);
xnor UO_2091 (O_2091,N_24208,N_24495);
nor UO_2092 (O_2092,N_24792,N_24580);
or UO_2093 (O_2093,N_24400,N_24553);
or UO_2094 (O_2094,N_24642,N_24564);
xor UO_2095 (O_2095,N_24917,N_24687);
xnor UO_2096 (O_2096,N_23966,N_24084);
nor UO_2097 (O_2097,N_23950,N_24594);
or UO_2098 (O_2098,N_24170,N_24746);
or UO_2099 (O_2099,N_24494,N_24511);
or UO_2100 (O_2100,N_24772,N_24660);
nor UO_2101 (O_2101,N_24034,N_24644);
xnor UO_2102 (O_2102,N_24939,N_24168);
nor UO_2103 (O_2103,N_24847,N_23916);
and UO_2104 (O_2104,N_23954,N_23827);
or UO_2105 (O_2105,N_24881,N_23781);
nand UO_2106 (O_2106,N_24058,N_23942);
and UO_2107 (O_2107,N_24067,N_24290);
nor UO_2108 (O_2108,N_24897,N_23782);
and UO_2109 (O_2109,N_24402,N_24700);
and UO_2110 (O_2110,N_24882,N_24628);
xnor UO_2111 (O_2111,N_24041,N_24053);
or UO_2112 (O_2112,N_24440,N_24781);
and UO_2113 (O_2113,N_23981,N_23753);
and UO_2114 (O_2114,N_23760,N_24050);
xnor UO_2115 (O_2115,N_24811,N_23823);
xnor UO_2116 (O_2116,N_23920,N_24958);
nor UO_2117 (O_2117,N_24301,N_23831);
and UO_2118 (O_2118,N_24875,N_24858);
nand UO_2119 (O_2119,N_24032,N_24795);
xor UO_2120 (O_2120,N_24474,N_24046);
xnor UO_2121 (O_2121,N_24470,N_24285);
and UO_2122 (O_2122,N_24493,N_23972);
and UO_2123 (O_2123,N_24560,N_24940);
or UO_2124 (O_2124,N_24629,N_24204);
or UO_2125 (O_2125,N_24493,N_24874);
and UO_2126 (O_2126,N_24135,N_24391);
or UO_2127 (O_2127,N_24986,N_23946);
xnor UO_2128 (O_2128,N_23792,N_24659);
nand UO_2129 (O_2129,N_24750,N_24590);
nand UO_2130 (O_2130,N_24225,N_23971);
nand UO_2131 (O_2131,N_24488,N_24007);
xnor UO_2132 (O_2132,N_24123,N_23776);
or UO_2133 (O_2133,N_24195,N_23983);
and UO_2134 (O_2134,N_23864,N_24636);
xor UO_2135 (O_2135,N_24105,N_24709);
xor UO_2136 (O_2136,N_24543,N_24090);
nand UO_2137 (O_2137,N_24520,N_24219);
or UO_2138 (O_2138,N_24957,N_24182);
nand UO_2139 (O_2139,N_24523,N_24755);
or UO_2140 (O_2140,N_24460,N_24067);
nand UO_2141 (O_2141,N_24053,N_24987);
or UO_2142 (O_2142,N_23767,N_24110);
or UO_2143 (O_2143,N_23829,N_24774);
nor UO_2144 (O_2144,N_24972,N_24949);
or UO_2145 (O_2145,N_24197,N_23882);
and UO_2146 (O_2146,N_24657,N_24293);
nor UO_2147 (O_2147,N_24274,N_24817);
nor UO_2148 (O_2148,N_24328,N_24791);
nor UO_2149 (O_2149,N_24739,N_24160);
nor UO_2150 (O_2150,N_24202,N_24497);
nor UO_2151 (O_2151,N_23870,N_24055);
xnor UO_2152 (O_2152,N_24773,N_23801);
xnor UO_2153 (O_2153,N_24353,N_24339);
nand UO_2154 (O_2154,N_24259,N_24758);
xnor UO_2155 (O_2155,N_24038,N_24582);
or UO_2156 (O_2156,N_24392,N_24785);
or UO_2157 (O_2157,N_24222,N_24395);
xnor UO_2158 (O_2158,N_24559,N_24207);
or UO_2159 (O_2159,N_24544,N_23910);
xor UO_2160 (O_2160,N_24110,N_24537);
nor UO_2161 (O_2161,N_24098,N_23798);
nand UO_2162 (O_2162,N_24117,N_24383);
or UO_2163 (O_2163,N_24211,N_23818);
or UO_2164 (O_2164,N_24820,N_24692);
nor UO_2165 (O_2165,N_24196,N_23754);
nor UO_2166 (O_2166,N_24435,N_24604);
and UO_2167 (O_2167,N_24939,N_24091);
nand UO_2168 (O_2168,N_24504,N_24421);
xor UO_2169 (O_2169,N_24445,N_24955);
nand UO_2170 (O_2170,N_24620,N_24353);
nor UO_2171 (O_2171,N_24022,N_24665);
or UO_2172 (O_2172,N_23980,N_24353);
nor UO_2173 (O_2173,N_24641,N_24613);
or UO_2174 (O_2174,N_24430,N_24041);
or UO_2175 (O_2175,N_24943,N_24868);
and UO_2176 (O_2176,N_24700,N_23889);
nand UO_2177 (O_2177,N_23895,N_24775);
and UO_2178 (O_2178,N_24124,N_24425);
or UO_2179 (O_2179,N_24551,N_24484);
nand UO_2180 (O_2180,N_24851,N_24107);
xor UO_2181 (O_2181,N_24553,N_23990);
nor UO_2182 (O_2182,N_24524,N_24872);
or UO_2183 (O_2183,N_24825,N_24968);
and UO_2184 (O_2184,N_23824,N_24790);
or UO_2185 (O_2185,N_24035,N_24150);
xor UO_2186 (O_2186,N_24318,N_24522);
and UO_2187 (O_2187,N_24200,N_24031);
xor UO_2188 (O_2188,N_24590,N_24633);
or UO_2189 (O_2189,N_24355,N_24348);
nand UO_2190 (O_2190,N_24393,N_24474);
and UO_2191 (O_2191,N_24027,N_24341);
or UO_2192 (O_2192,N_23982,N_24044);
or UO_2193 (O_2193,N_24356,N_24786);
nand UO_2194 (O_2194,N_24935,N_24505);
and UO_2195 (O_2195,N_24062,N_24098);
nand UO_2196 (O_2196,N_24541,N_23941);
xnor UO_2197 (O_2197,N_24810,N_24791);
and UO_2198 (O_2198,N_24503,N_24836);
xor UO_2199 (O_2199,N_24401,N_24040);
or UO_2200 (O_2200,N_23944,N_23804);
or UO_2201 (O_2201,N_23983,N_24554);
or UO_2202 (O_2202,N_24819,N_24171);
nand UO_2203 (O_2203,N_24174,N_24556);
nor UO_2204 (O_2204,N_24678,N_24268);
nor UO_2205 (O_2205,N_24303,N_24451);
nand UO_2206 (O_2206,N_24719,N_24040);
nor UO_2207 (O_2207,N_24934,N_23820);
xor UO_2208 (O_2208,N_24861,N_23974);
and UO_2209 (O_2209,N_23984,N_24618);
nand UO_2210 (O_2210,N_23836,N_24766);
and UO_2211 (O_2211,N_23853,N_24434);
and UO_2212 (O_2212,N_24877,N_24724);
nand UO_2213 (O_2213,N_24864,N_24811);
and UO_2214 (O_2214,N_24314,N_24989);
and UO_2215 (O_2215,N_24295,N_24455);
or UO_2216 (O_2216,N_24885,N_24341);
xnor UO_2217 (O_2217,N_24601,N_24524);
xnor UO_2218 (O_2218,N_24838,N_24476);
nand UO_2219 (O_2219,N_24017,N_24134);
xnor UO_2220 (O_2220,N_24940,N_24815);
nor UO_2221 (O_2221,N_24359,N_24913);
nand UO_2222 (O_2222,N_24846,N_24232);
nand UO_2223 (O_2223,N_24316,N_24960);
nor UO_2224 (O_2224,N_23841,N_23813);
xnor UO_2225 (O_2225,N_24184,N_24399);
and UO_2226 (O_2226,N_24104,N_24426);
and UO_2227 (O_2227,N_23899,N_24602);
xnor UO_2228 (O_2228,N_23788,N_24845);
nor UO_2229 (O_2229,N_24904,N_24162);
nand UO_2230 (O_2230,N_24664,N_23796);
nand UO_2231 (O_2231,N_23804,N_24244);
xnor UO_2232 (O_2232,N_24835,N_24979);
xnor UO_2233 (O_2233,N_24700,N_24501);
xnor UO_2234 (O_2234,N_24769,N_24233);
nor UO_2235 (O_2235,N_23768,N_24427);
and UO_2236 (O_2236,N_24284,N_24717);
or UO_2237 (O_2237,N_24180,N_24716);
nand UO_2238 (O_2238,N_23979,N_24624);
and UO_2239 (O_2239,N_24305,N_24495);
and UO_2240 (O_2240,N_24491,N_24889);
and UO_2241 (O_2241,N_24810,N_24850);
or UO_2242 (O_2242,N_24732,N_24045);
or UO_2243 (O_2243,N_23929,N_24183);
xnor UO_2244 (O_2244,N_24159,N_24122);
or UO_2245 (O_2245,N_23841,N_24635);
and UO_2246 (O_2246,N_24996,N_24687);
and UO_2247 (O_2247,N_23911,N_24011);
xnor UO_2248 (O_2248,N_24449,N_24310);
and UO_2249 (O_2249,N_24981,N_24017);
nor UO_2250 (O_2250,N_24882,N_24676);
or UO_2251 (O_2251,N_24002,N_24387);
nor UO_2252 (O_2252,N_24662,N_23919);
nand UO_2253 (O_2253,N_24881,N_24519);
nor UO_2254 (O_2254,N_23985,N_24673);
and UO_2255 (O_2255,N_24813,N_23792);
nand UO_2256 (O_2256,N_24544,N_24383);
nand UO_2257 (O_2257,N_24204,N_24630);
xor UO_2258 (O_2258,N_24640,N_24786);
and UO_2259 (O_2259,N_24478,N_23822);
and UO_2260 (O_2260,N_24158,N_24609);
or UO_2261 (O_2261,N_24952,N_24375);
xor UO_2262 (O_2262,N_23837,N_24360);
or UO_2263 (O_2263,N_24932,N_24644);
nor UO_2264 (O_2264,N_24567,N_24704);
nor UO_2265 (O_2265,N_24649,N_24684);
nor UO_2266 (O_2266,N_24579,N_23973);
or UO_2267 (O_2267,N_24100,N_24369);
nor UO_2268 (O_2268,N_24356,N_24249);
nor UO_2269 (O_2269,N_23764,N_24008);
nand UO_2270 (O_2270,N_24921,N_24681);
or UO_2271 (O_2271,N_24409,N_24540);
xor UO_2272 (O_2272,N_23821,N_23892);
nor UO_2273 (O_2273,N_24241,N_24804);
nor UO_2274 (O_2274,N_24936,N_24891);
and UO_2275 (O_2275,N_24377,N_24877);
xor UO_2276 (O_2276,N_24988,N_24876);
nand UO_2277 (O_2277,N_24472,N_24829);
nand UO_2278 (O_2278,N_24678,N_24413);
xnor UO_2279 (O_2279,N_23941,N_24373);
nand UO_2280 (O_2280,N_24047,N_23849);
or UO_2281 (O_2281,N_24957,N_24885);
or UO_2282 (O_2282,N_23890,N_24344);
and UO_2283 (O_2283,N_24552,N_23832);
and UO_2284 (O_2284,N_24099,N_24595);
nand UO_2285 (O_2285,N_24291,N_23864);
or UO_2286 (O_2286,N_24434,N_24086);
nand UO_2287 (O_2287,N_23933,N_23819);
nor UO_2288 (O_2288,N_24868,N_23771);
xnor UO_2289 (O_2289,N_24597,N_24235);
nand UO_2290 (O_2290,N_24855,N_23977);
nor UO_2291 (O_2291,N_24521,N_24724);
or UO_2292 (O_2292,N_24768,N_24890);
or UO_2293 (O_2293,N_24991,N_24484);
nor UO_2294 (O_2294,N_24950,N_24145);
xnor UO_2295 (O_2295,N_24819,N_24540);
or UO_2296 (O_2296,N_24437,N_24905);
xor UO_2297 (O_2297,N_23859,N_24300);
nand UO_2298 (O_2298,N_23900,N_24959);
or UO_2299 (O_2299,N_24929,N_23978);
and UO_2300 (O_2300,N_24463,N_23891);
or UO_2301 (O_2301,N_23867,N_24085);
nor UO_2302 (O_2302,N_24171,N_24367);
xor UO_2303 (O_2303,N_23993,N_24229);
nor UO_2304 (O_2304,N_23834,N_24167);
or UO_2305 (O_2305,N_23927,N_24297);
nand UO_2306 (O_2306,N_23848,N_24495);
and UO_2307 (O_2307,N_24404,N_24731);
and UO_2308 (O_2308,N_23910,N_24682);
xnor UO_2309 (O_2309,N_24343,N_24609);
nor UO_2310 (O_2310,N_24359,N_24076);
and UO_2311 (O_2311,N_24236,N_24967);
xnor UO_2312 (O_2312,N_24764,N_24425);
and UO_2313 (O_2313,N_23841,N_24703);
nand UO_2314 (O_2314,N_24127,N_24551);
nor UO_2315 (O_2315,N_24478,N_24002);
nand UO_2316 (O_2316,N_24476,N_24839);
nand UO_2317 (O_2317,N_24605,N_23980);
nor UO_2318 (O_2318,N_23819,N_24284);
nand UO_2319 (O_2319,N_24179,N_24982);
and UO_2320 (O_2320,N_23993,N_24457);
and UO_2321 (O_2321,N_23780,N_24087);
nor UO_2322 (O_2322,N_24825,N_24068);
or UO_2323 (O_2323,N_23828,N_24652);
xnor UO_2324 (O_2324,N_24636,N_24959);
xnor UO_2325 (O_2325,N_24167,N_23922);
nor UO_2326 (O_2326,N_24080,N_24342);
and UO_2327 (O_2327,N_24946,N_24334);
and UO_2328 (O_2328,N_23766,N_23767);
and UO_2329 (O_2329,N_24681,N_24133);
nand UO_2330 (O_2330,N_24706,N_24711);
or UO_2331 (O_2331,N_24220,N_24976);
nand UO_2332 (O_2332,N_24835,N_24151);
nand UO_2333 (O_2333,N_24704,N_23835);
and UO_2334 (O_2334,N_24664,N_24003);
nand UO_2335 (O_2335,N_24691,N_24515);
or UO_2336 (O_2336,N_24136,N_24847);
or UO_2337 (O_2337,N_24778,N_24346);
nor UO_2338 (O_2338,N_24711,N_24298);
or UO_2339 (O_2339,N_24775,N_24545);
or UO_2340 (O_2340,N_24694,N_24414);
nand UO_2341 (O_2341,N_24227,N_24037);
xor UO_2342 (O_2342,N_23880,N_24922);
nor UO_2343 (O_2343,N_23776,N_24621);
and UO_2344 (O_2344,N_24255,N_24518);
xor UO_2345 (O_2345,N_24604,N_24306);
and UO_2346 (O_2346,N_24521,N_23920);
and UO_2347 (O_2347,N_24043,N_23769);
or UO_2348 (O_2348,N_23773,N_24464);
and UO_2349 (O_2349,N_23868,N_24109);
xor UO_2350 (O_2350,N_24742,N_23913);
xor UO_2351 (O_2351,N_23795,N_24933);
xor UO_2352 (O_2352,N_24270,N_24506);
and UO_2353 (O_2353,N_24489,N_24734);
and UO_2354 (O_2354,N_24071,N_24196);
xnor UO_2355 (O_2355,N_24226,N_23898);
and UO_2356 (O_2356,N_24315,N_24939);
nor UO_2357 (O_2357,N_24713,N_24185);
xnor UO_2358 (O_2358,N_23859,N_23986);
or UO_2359 (O_2359,N_23854,N_24608);
or UO_2360 (O_2360,N_24143,N_24590);
or UO_2361 (O_2361,N_23980,N_24018);
xnor UO_2362 (O_2362,N_24584,N_24712);
xor UO_2363 (O_2363,N_24997,N_24588);
nor UO_2364 (O_2364,N_24513,N_24113);
nand UO_2365 (O_2365,N_23968,N_24282);
xor UO_2366 (O_2366,N_24090,N_24442);
or UO_2367 (O_2367,N_24128,N_23965);
nand UO_2368 (O_2368,N_24384,N_24409);
and UO_2369 (O_2369,N_23862,N_24636);
or UO_2370 (O_2370,N_24647,N_24323);
or UO_2371 (O_2371,N_24882,N_24370);
nand UO_2372 (O_2372,N_24019,N_24223);
nor UO_2373 (O_2373,N_24625,N_23772);
and UO_2374 (O_2374,N_24302,N_24488);
nor UO_2375 (O_2375,N_24444,N_24377);
or UO_2376 (O_2376,N_24601,N_24883);
xnor UO_2377 (O_2377,N_24378,N_24454);
xor UO_2378 (O_2378,N_24055,N_24252);
xnor UO_2379 (O_2379,N_23973,N_24241);
or UO_2380 (O_2380,N_23954,N_24828);
nor UO_2381 (O_2381,N_23892,N_24224);
or UO_2382 (O_2382,N_24239,N_24274);
xnor UO_2383 (O_2383,N_24594,N_24670);
or UO_2384 (O_2384,N_23931,N_24597);
nor UO_2385 (O_2385,N_24918,N_24516);
and UO_2386 (O_2386,N_24882,N_24785);
nand UO_2387 (O_2387,N_23841,N_24090);
or UO_2388 (O_2388,N_24763,N_24500);
or UO_2389 (O_2389,N_24984,N_24961);
nand UO_2390 (O_2390,N_24247,N_24979);
nand UO_2391 (O_2391,N_24827,N_24056);
xor UO_2392 (O_2392,N_24432,N_24547);
or UO_2393 (O_2393,N_24397,N_24403);
nor UO_2394 (O_2394,N_23983,N_24971);
or UO_2395 (O_2395,N_24876,N_24400);
xnor UO_2396 (O_2396,N_24788,N_23997);
xor UO_2397 (O_2397,N_24464,N_24466);
nand UO_2398 (O_2398,N_23921,N_24776);
or UO_2399 (O_2399,N_24561,N_24948);
xnor UO_2400 (O_2400,N_24624,N_24221);
nand UO_2401 (O_2401,N_24880,N_24222);
nand UO_2402 (O_2402,N_23813,N_24843);
and UO_2403 (O_2403,N_24985,N_24651);
and UO_2404 (O_2404,N_24860,N_24687);
nor UO_2405 (O_2405,N_24685,N_23808);
nand UO_2406 (O_2406,N_24418,N_24895);
xor UO_2407 (O_2407,N_24150,N_24593);
nand UO_2408 (O_2408,N_23861,N_24995);
xnor UO_2409 (O_2409,N_23979,N_24265);
nor UO_2410 (O_2410,N_24594,N_24491);
xor UO_2411 (O_2411,N_24732,N_24551);
nor UO_2412 (O_2412,N_24481,N_23956);
xnor UO_2413 (O_2413,N_23927,N_24898);
nor UO_2414 (O_2414,N_24420,N_24289);
nand UO_2415 (O_2415,N_23928,N_24217);
nor UO_2416 (O_2416,N_23789,N_24747);
xnor UO_2417 (O_2417,N_24837,N_24521);
nor UO_2418 (O_2418,N_24093,N_24452);
and UO_2419 (O_2419,N_24502,N_24087);
nor UO_2420 (O_2420,N_24223,N_24894);
and UO_2421 (O_2421,N_24642,N_23851);
and UO_2422 (O_2422,N_23841,N_23842);
nand UO_2423 (O_2423,N_24218,N_24067);
nand UO_2424 (O_2424,N_23975,N_24122);
nor UO_2425 (O_2425,N_23911,N_24803);
nor UO_2426 (O_2426,N_23991,N_24550);
nand UO_2427 (O_2427,N_24235,N_24768);
and UO_2428 (O_2428,N_24706,N_24030);
or UO_2429 (O_2429,N_23770,N_24654);
nand UO_2430 (O_2430,N_24487,N_24636);
or UO_2431 (O_2431,N_23794,N_24842);
nor UO_2432 (O_2432,N_24335,N_24169);
or UO_2433 (O_2433,N_24680,N_24646);
nor UO_2434 (O_2434,N_24864,N_23943);
nor UO_2435 (O_2435,N_24277,N_24553);
nand UO_2436 (O_2436,N_23888,N_24665);
nor UO_2437 (O_2437,N_24758,N_24645);
xor UO_2438 (O_2438,N_24515,N_24894);
nor UO_2439 (O_2439,N_24979,N_24677);
nand UO_2440 (O_2440,N_24147,N_24591);
or UO_2441 (O_2441,N_24083,N_24776);
or UO_2442 (O_2442,N_24062,N_24038);
nand UO_2443 (O_2443,N_23860,N_24986);
nand UO_2444 (O_2444,N_24883,N_24466);
and UO_2445 (O_2445,N_24219,N_24966);
nand UO_2446 (O_2446,N_23793,N_24776);
nor UO_2447 (O_2447,N_24814,N_24870);
and UO_2448 (O_2448,N_24868,N_24618);
and UO_2449 (O_2449,N_24528,N_24421);
and UO_2450 (O_2450,N_24194,N_23995);
or UO_2451 (O_2451,N_23908,N_24196);
nand UO_2452 (O_2452,N_24904,N_24444);
nor UO_2453 (O_2453,N_24882,N_23873);
or UO_2454 (O_2454,N_24521,N_24310);
nor UO_2455 (O_2455,N_23860,N_24547);
or UO_2456 (O_2456,N_24713,N_24461);
nor UO_2457 (O_2457,N_24040,N_23838);
and UO_2458 (O_2458,N_24846,N_23925);
or UO_2459 (O_2459,N_23919,N_24392);
nand UO_2460 (O_2460,N_24925,N_24653);
xnor UO_2461 (O_2461,N_24998,N_24471);
xor UO_2462 (O_2462,N_23801,N_24078);
and UO_2463 (O_2463,N_24417,N_24161);
xor UO_2464 (O_2464,N_23902,N_24831);
nor UO_2465 (O_2465,N_24468,N_23880);
or UO_2466 (O_2466,N_24966,N_24168);
and UO_2467 (O_2467,N_23764,N_23805);
or UO_2468 (O_2468,N_24498,N_24804);
nor UO_2469 (O_2469,N_24242,N_23826);
nand UO_2470 (O_2470,N_24420,N_24798);
nor UO_2471 (O_2471,N_24122,N_24003);
xnor UO_2472 (O_2472,N_24921,N_24118);
or UO_2473 (O_2473,N_23874,N_24867);
or UO_2474 (O_2474,N_24213,N_23752);
nor UO_2475 (O_2475,N_24426,N_24951);
and UO_2476 (O_2476,N_24236,N_24316);
or UO_2477 (O_2477,N_24985,N_23920);
and UO_2478 (O_2478,N_24312,N_23798);
or UO_2479 (O_2479,N_24458,N_24572);
xnor UO_2480 (O_2480,N_24341,N_24100);
and UO_2481 (O_2481,N_24665,N_24836);
nand UO_2482 (O_2482,N_23978,N_24723);
nor UO_2483 (O_2483,N_23877,N_24152);
nand UO_2484 (O_2484,N_24846,N_24869);
or UO_2485 (O_2485,N_24450,N_23976);
and UO_2486 (O_2486,N_24024,N_24794);
or UO_2487 (O_2487,N_24751,N_24554);
or UO_2488 (O_2488,N_24910,N_24604);
xor UO_2489 (O_2489,N_24952,N_24029);
nor UO_2490 (O_2490,N_24814,N_23758);
and UO_2491 (O_2491,N_23815,N_24423);
xnor UO_2492 (O_2492,N_24716,N_24222);
xnor UO_2493 (O_2493,N_24508,N_24162);
nor UO_2494 (O_2494,N_24097,N_23820);
nand UO_2495 (O_2495,N_23839,N_24713);
nor UO_2496 (O_2496,N_24636,N_24029);
nor UO_2497 (O_2497,N_24493,N_24772);
or UO_2498 (O_2498,N_24370,N_24226);
xor UO_2499 (O_2499,N_24812,N_24025);
nor UO_2500 (O_2500,N_24335,N_24511);
nand UO_2501 (O_2501,N_23889,N_24278);
nand UO_2502 (O_2502,N_24331,N_24368);
or UO_2503 (O_2503,N_24097,N_24033);
or UO_2504 (O_2504,N_24706,N_24029);
nor UO_2505 (O_2505,N_24892,N_24881);
nor UO_2506 (O_2506,N_24261,N_24491);
nor UO_2507 (O_2507,N_24419,N_24578);
nand UO_2508 (O_2508,N_23906,N_24939);
nand UO_2509 (O_2509,N_24859,N_24208);
nand UO_2510 (O_2510,N_23900,N_24309);
and UO_2511 (O_2511,N_23886,N_24019);
and UO_2512 (O_2512,N_23872,N_24566);
nor UO_2513 (O_2513,N_24754,N_24899);
xor UO_2514 (O_2514,N_24064,N_24544);
nand UO_2515 (O_2515,N_23791,N_24042);
or UO_2516 (O_2516,N_24702,N_24689);
and UO_2517 (O_2517,N_24922,N_24648);
xor UO_2518 (O_2518,N_23911,N_24020);
nor UO_2519 (O_2519,N_24007,N_24677);
nand UO_2520 (O_2520,N_24315,N_24337);
and UO_2521 (O_2521,N_24006,N_24961);
xnor UO_2522 (O_2522,N_24311,N_24238);
and UO_2523 (O_2523,N_24720,N_24026);
or UO_2524 (O_2524,N_24137,N_24139);
nor UO_2525 (O_2525,N_24479,N_24860);
or UO_2526 (O_2526,N_24010,N_24740);
nor UO_2527 (O_2527,N_23935,N_24577);
nand UO_2528 (O_2528,N_23753,N_24008);
or UO_2529 (O_2529,N_24465,N_24199);
xnor UO_2530 (O_2530,N_24346,N_24693);
or UO_2531 (O_2531,N_24496,N_24184);
xnor UO_2532 (O_2532,N_24216,N_24375);
nand UO_2533 (O_2533,N_24560,N_24665);
or UO_2534 (O_2534,N_23984,N_24755);
or UO_2535 (O_2535,N_24408,N_23885);
or UO_2536 (O_2536,N_24485,N_23818);
and UO_2537 (O_2537,N_24935,N_24345);
nor UO_2538 (O_2538,N_24576,N_24303);
nand UO_2539 (O_2539,N_24269,N_23896);
and UO_2540 (O_2540,N_24161,N_24919);
or UO_2541 (O_2541,N_24885,N_24842);
or UO_2542 (O_2542,N_24718,N_24915);
or UO_2543 (O_2543,N_23751,N_24229);
and UO_2544 (O_2544,N_24560,N_23916);
xor UO_2545 (O_2545,N_24130,N_24282);
or UO_2546 (O_2546,N_24358,N_24680);
nor UO_2547 (O_2547,N_24856,N_23898);
xor UO_2548 (O_2548,N_24833,N_24701);
nand UO_2549 (O_2549,N_24624,N_23868);
nor UO_2550 (O_2550,N_23820,N_24587);
xnor UO_2551 (O_2551,N_24860,N_24109);
or UO_2552 (O_2552,N_24365,N_24147);
nand UO_2553 (O_2553,N_24191,N_24471);
nor UO_2554 (O_2554,N_24826,N_24359);
nand UO_2555 (O_2555,N_24151,N_24802);
xor UO_2556 (O_2556,N_23790,N_24935);
xnor UO_2557 (O_2557,N_24409,N_24552);
or UO_2558 (O_2558,N_24748,N_23885);
xnor UO_2559 (O_2559,N_24077,N_24036);
xor UO_2560 (O_2560,N_24211,N_23829);
nor UO_2561 (O_2561,N_24389,N_23956);
nand UO_2562 (O_2562,N_24182,N_23794);
nand UO_2563 (O_2563,N_24979,N_24444);
or UO_2564 (O_2564,N_24662,N_24434);
nand UO_2565 (O_2565,N_24885,N_24429);
and UO_2566 (O_2566,N_24512,N_24335);
nand UO_2567 (O_2567,N_24996,N_24299);
xnor UO_2568 (O_2568,N_23876,N_24448);
nand UO_2569 (O_2569,N_24461,N_23791);
nand UO_2570 (O_2570,N_24862,N_24858);
nand UO_2571 (O_2571,N_24394,N_24979);
or UO_2572 (O_2572,N_24193,N_24873);
and UO_2573 (O_2573,N_24385,N_23849);
xor UO_2574 (O_2574,N_23832,N_24934);
or UO_2575 (O_2575,N_24534,N_24305);
nor UO_2576 (O_2576,N_24319,N_24016);
nand UO_2577 (O_2577,N_24470,N_24993);
xnor UO_2578 (O_2578,N_23752,N_24815);
nand UO_2579 (O_2579,N_24832,N_24520);
nand UO_2580 (O_2580,N_24922,N_24621);
nor UO_2581 (O_2581,N_24771,N_24754);
nor UO_2582 (O_2582,N_24039,N_24310);
and UO_2583 (O_2583,N_24095,N_24207);
and UO_2584 (O_2584,N_24467,N_24254);
or UO_2585 (O_2585,N_24375,N_24074);
xnor UO_2586 (O_2586,N_23751,N_24266);
nor UO_2587 (O_2587,N_24474,N_24664);
xnor UO_2588 (O_2588,N_24202,N_24399);
and UO_2589 (O_2589,N_24452,N_24233);
or UO_2590 (O_2590,N_24223,N_24590);
nand UO_2591 (O_2591,N_24751,N_24958);
nand UO_2592 (O_2592,N_24222,N_24728);
nor UO_2593 (O_2593,N_24845,N_24850);
xnor UO_2594 (O_2594,N_24088,N_24647);
and UO_2595 (O_2595,N_24061,N_24077);
nor UO_2596 (O_2596,N_23849,N_24242);
nor UO_2597 (O_2597,N_23925,N_24856);
and UO_2598 (O_2598,N_24744,N_24764);
nand UO_2599 (O_2599,N_23796,N_24281);
or UO_2600 (O_2600,N_24416,N_24958);
or UO_2601 (O_2601,N_23914,N_24155);
or UO_2602 (O_2602,N_24262,N_23847);
or UO_2603 (O_2603,N_24473,N_24859);
nand UO_2604 (O_2604,N_23843,N_24808);
or UO_2605 (O_2605,N_23759,N_23957);
nand UO_2606 (O_2606,N_24796,N_23843);
and UO_2607 (O_2607,N_24947,N_24909);
and UO_2608 (O_2608,N_24153,N_23850);
xor UO_2609 (O_2609,N_24796,N_24330);
nor UO_2610 (O_2610,N_24992,N_24432);
nand UO_2611 (O_2611,N_24710,N_23990);
xor UO_2612 (O_2612,N_24364,N_24935);
xnor UO_2613 (O_2613,N_24759,N_23951);
and UO_2614 (O_2614,N_23879,N_23764);
xnor UO_2615 (O_2615,N_24824,N_24058);
and UO_2616 (O_2616,N_24945,N_24024);
xor UO_2617 (O_2617,N_24219,N_24636);
and UO_2618 (O_2618,N_24730,N_24429);
xor UO_2619 (O_2619,N_23866,N_24338);
nor UO_2620 (O_2620,N_24733,N_24207);
xnor UO_2621 (O_2621,N_24027,N_23905);
or UO_2622 (O_2622,N_23902,N_24765);
and UO_2623 (O_2623,N_24597,N_24583);
or UO_2624 (O_2624,N_24113,N_23901);
nand UO_2625 (O_2625,N_24040,N_24128);
or UO_2626 (O_2626,N_24097,N_24276);
and UO_2627 (O_2627,N_24452,N_24948);
and UO_2628 (O_2628,N_24772,N_24064);
nor UO_2629 (O_2629,N_24716,N_24425);
nand UO_2630 (O_2630,N_24802,N_24695);
nor UO_2631 (O_2631,N_24736,N_24811);
xor UO_2632 (O_2632,N_24134,N_24281);
nand UO_2633 (O_2633,N_24599,N_24645);
xor UO_2634 (O_2634,N_23957,N_24406);
xnor UO_2635 (O_2635,N_24022,N_24356);
or UO_2636 (O_2636,N_24400,N_24719);
and UO_2637 (O_2637,N_23825,N_24550);
xor UO_2638 (O_2638,N_24052,N_24945);
nor UO_2639 (O_2639,N_24503,N_24230);
xnor UO_2640 (O_2640,N_23846,N_23820);
and UO_2641 (O_2641,N_23755,N_24739);
nand UO_2642 (O_2642,N_24104,N_24084);
xnor UO_2643 (O_2643,N_24736,N_24118);
nand UO_2644 (O_2644,N_24341,N_24600);
or UO_2645 (O_2645,N_24843,N_24937);
and UO_2646 (O_2646,N_24354,N_23772);
xnor UO_2647 (O_2647,N_24949,N_24993);
nor UO_2648 (O_2648,N_24561,N_24550);
nand UO_2649 (O_2649,N_24888,N_24112);
nand UO_2650 (O_2650,N_24632,N_24901);
nor UO_2651 (O_2651,N_24649,N_24715);
nand UO_2652 (O_2652,N_24049,N_23906);
xor UO_2653 (O_2653,N_24985,N_24769);
and UO_2654 (O_2654,N_24808,N_24878);
nand UO_2655 (O_2655,N_24039,N_24476);
xor UO_2656 (O_2656,N_23974,N_23852);
and UO_2657 (O_2657,N_24574,N_24823);
and UO_2658 (O_2658,N_24653,N_24525);
nand UO_2659 (O_2659,N_24745,N_24784);
nor UO_2660 (O_2660,N_24963,N_23786);
nor UO_2661 (O_2661,N_24739,N_24908);
or UO_2662 (O_2662,N_24938,N_24277);
nor UO_2663 (O_2663,N_24954,N_24082);
nor UO_2664 (O_2664,N_24989,N_23866);
or UO_2665 (O_2665,N_24008,N_23842);
nor UO_2666 (O_2666,N_24292,N_24362);
or UO_2667 (O_2667,N_23836,N_24526);
nand UO_2668 (O_2668,N_24621,N_24834);
nand UO_2669 (O_2669,N_24425,N_24731);
nor UO_2670 (O_2670,N_24667,N_24956);
or UO_2671 (O_2671,N_24623,N_24673);
nor UO_2672 (O_2672,N_24826,N_23784);
xor UO_2673 (O_2673,N_24833,N_24427);
and UO_2674 (O_2674,N_24434,N_24597);
or UO_2675 (O_2675,N_23931,N_23955);
nand UO_2676 (O_2676,N_24864,N_24646);
xor UO_2677 (O_2677,N_24497,N_23778);
nand UO_2678 (O_2678,N_23839,N_24984);
nand UO_2679 (O_2679,N_24545,N_24815);
xor UO_2680 (O_2680,N_24338,N_24069);
nand UO_2681 (O_2681,N_24198,N_24526);
or UO_2682 (O_2682,N_24619,N_24803);
nand UO_2683 (O_2683,N_24322,N_24331);
or UO_2684 (O_2684,N_24657,N_23885);
or UO_2685 (O_2685,N_24888,N_24373);
xor UO_2686 (O_2686,N_24979,N_24705);
nor UO_2687 (O_2687,N_24293,N_24262);
nor UO_2688 (O_2688,N_23824,N_24281);
or UO_2689 (O_2689,N_24080,N_23773);
and UO_2690 (O_2690,N_24867,N_24580);
xor UO_2691 (O_2691,N_24586,N_24790);
and UO_2692 (O_2692,N_24009,N_24290);
nand UO_2693 (O_2693,N_24240,N_24555);
or UO_2694 (O_2694,N_24689,N_24976);
or UO_2695 (O_2695,N_24269,N_24156);
xor UO_2696 (O_2696,N_24583,N_24888);
xor UO_2697 (O_2697,N_23904,N_24960);
xor UO_2698 (O_2698,N_24432,N_23945);
xor UO_2699 (O_2699,N_24486,N_24455);
nand UO_2700 (O_2700,N_23883,N_24946);
xor UO_2701 (O_2701,N_23915,N_24692);
xnor UO_2702 (O_2702,N_24343,N_24774);
nor UO_2703 (O_2703,N_23768,N_24278);
or UO_2704 (O_2704,N_23804,N_24279);
nand UO_2705 (O_2705,N_24456,N_24503);
nand UO_2706 (O_2706,N_24095,N_24260);
or UO_2707 (O_2707,N_24059,N_24927);
nand UO_2708 (O_2708,N_24231,N_23765);
or UO_2709 (O_2709,N_24954,N_24562);
xor UO_2710 (O_2710,N_24024,N_23793);
and UO_2711 (O_2711,N_24813,N_24260);
nand UO_2712 (O_2712,N_23923,N_24152);
or UO_2713 (O_2713,N_24964,N_24171);
nor UO_2714 (O_2714,N_24934,N_24236);
and UO_2715 (O_2715,N_24011,N_23897);
and UO_2716 (O_2716,N_24140,N_24872);
xnor UO_2717 (O_2717,N_24339,N_24674);
and UO_2718 (O_2718,N_24076,N_23920);
nand UO_2719 (O_2719,N_24881,N_24171);
nor UO_2720 (O_2720,N_24275,N_24574);
or UO_2721 (O_2721,N_24728,N_24374);
nand UO_2722 (O_2722,N_23899,N_24116);
and UO_2723 (O_2723,N_24930,N_23856);
nand UO_2724 (O_2724,N_24064,N_23816);
nand UO_2725 (O_2725,N_24839,N_23842);
or UO_2726 (O_2726,N_24502,N_24819);
nor UO_2727 (O_2727,N_23757,N_24463);
or UO_2728 (O_2728,N_24926,N_24736);
or UO_2729 (O_2729,N_24521,N_23857);
nand UO_2730 (O_2730,N_24018,N_24967);
or UO_2731 (O_2731,N_24840,N_24921);
and UO_2732 (O_2732,N_24393,N_24407);
and UO_2733 (O_2733,N_24375,N_24500);
nor UO_2734 (O_2734,N_24148,N_24756);
nor UO_2735 (O_2735,N_24771,N_23850);
or UO_2736 (O_2736,N_24687,N_24187);
and UO_2737 (O_2737,N_23882,N_24517);
and UO_2738 (O_2738,N_24160,N_24829);
nor UO_2739 (O_2739,N_24806,N_24404);
xnor UO_2740 (O_2740,N_24485,N_24274);
nand UO_2741 (O_2741,N_24280,N_24795);
and UO_2742 (O_2742,N_24823,N_24001);
xnor UO_2743 (O_2743,N_24964,N_23902);
nand UO_2744 (O_2744,N_24366,N_24211);
nand UO_2745 (O_2745,N_24640,N_24961);
or UO_2746 (O_2746,N_24407,N_24031);
nor UO_2747 (O_2747,N_23780,N_24842);
xnor UO_2748 (O_2748,N_24034,N_24370);
nor UO_2749 (O_2749,N_24753,N_24097);
nor UO_2750 (O_2750,N_23923,N_24633);
or UO_2751 (O_2751,N_24382,N_24550);
and UO_2752 (O_2752,N_24864,N_23928);
and UO_2753 (O_2753,N_24479,N_24153);
and UO_2754 (O_2754,N_24610,N_24790);
xor UO_2755 (O_2755,N_24459,N_24100);
and UO_2756 (O_2756,N_24157,N_24509);
nor UO_2757 (O_2757,N_24763,N_24774);
or UO_2758 (O_2758,N_24657,N_23874);
xor UO_2759 (O_2759,N_24921,N_24256);
nand UO_2760 (O_2760,N_24279,N_24122);
and UO_2761 (O_2761,N_24500,N_24563);
nand UO_2762 (O_2762,N_24415,N_23975);
or UO_2763 (O_2763,N_24508,N_24249);
nand UO_2764 (O_2764,N_24734,N_24990);
xor UO_2765 (O_2765,N_23928,N_24707);
nand UO_2766 (O_2766,N_24986,N_24914);
nor UO_2767 (O_2767,N_24163,N_24844);
nor UO_2768 (O_2768,N_24265,N_23860);
nor UO_2769 (O_2769,N_24042,N_24918);
xnor UO_2770 (O_2770,N_24805,N_23927);
nand UO_2771 (O_2771,N_23854,N_24939);
and UO_2772 (O_2772,N_24339,N_24776);
nor UO_2773 (O_2773,N_23871,N_24151);
nor UO_2774 (O_2774,N_24661,N_24551);
and UO_2775 (O_2775,N_24958,N_24212);
and UO_2776 (O_2776,N_24843,N_24477);
nor UO_2777 (O_2777,N_24236,N_24622);
xor UO_2778 (O_2778,N_23854,N_23859);
and UO_2779 (O_2779,N_24828,N_23996);
nor UO_2780 (O_2780,N_24001,N_24601);
xor UO_2781 (O_2781,N_24081,N_24782);
nand UO_2782 (O_2782,N_24106,N_24189);
xnor UO_2783 (O_2783,N_24126,N_23800);
xnor UO_2784 (O_2784,N_24607,N_23920);
nand UO_2785 (O_2785,N_24026,N_24315);
or UO_2786 (O_2786,N_24650,N_24980);
or UO_2787 (O_2787,N_23917,N_24342);
or UO_2788 (O_2788,N_24590,N_24943);
and UO_2789 (O_2789,N_23752,N_24302);
or UO_2790 (O_2790,N_24258,N_24262);
and UO_2791 (O_2791,N_24972,N_24038);
nand UO_2792 (O_2792,N_24471,N_24979);
and UO_2793 (O_2793,N_24527,N_24435);
and UO_2794 (O_2794,N_24642,N_24738);
xnor UO_2795 (O_2795,N_24847,N_24737);
nand UO_2796 (O_2796,N_24553,N_23772);
or UO_2797 (O_2797,N_24983,N_24442);
or UO_2798 (O_2798,N_23755,N_24326);
nor UO_2799 (O_2799,N_24612,N_24833);
xor UO_2800 (O_2800,N_24311,N_23831);
nand UO_2801 (O_2801,N_24135,N_24279);
nand UO_2802 (O_2802,N_24969,N_24843);
nor UO_2803 (O_2803,N_24599,N_24008);
xor UO_2804 (O_2804,N_24109,N_24099);
nor UO_2805 (O_2805,N_24464,N_24991);
xor UO_2806 (O_2806,N_24159,N_24625);
and UO_2807 (O_2807,N_24027,N_24460);
or UO_2808 (O_2808,N_24598,N_23851);
xnor UO_2809 (O_2809,N_24443,N_24752);
and UO_2810 (O_2810,N_23799,N_24675);
nor UO_2811 (O_2811,N_24767,N_23982);
xor UO_2812 (O_2812,N_23758,N_24424);
or UO_2813 (O_2813,N_23822,N_24196);
xnor UO_2814 (O_2814,N_24829,N_24803);
and UO_2815 (O_2815,N_24974,N_24413);
nor UO_2816 (O_2816,N_24879,N_24792);
xnor UO_2817 (O_2817,N_23916,N_23900);
nand UO_2818 (O_2818,N_24138,N_24154);
or UO_2819 (O_2819,N_24799,N_24827);
and UO_2820 (O_2820,N_24898,N_24489);
or UO_2821 (O_2821,N_24349,N_23808);
nand UO_2822 (O_2822,N_24929,N_24451);
and UO_2823 (O_2823,N_24031,N_24331);
or UO_2824 (O_2824,N_24988,N_24546);
nand UO_2825 (O_2825,N_23957,N_24025);
xor UO_2826 (O_2826,N_24389,N_24837);
nor UO_2827 (O_2827,N_24324,N_24262);
nor UO_2828 (O_2828,N_24851,N_24177);
nand UO_2829 (O_2829,N_24492,N_24188);
or UO_2830 (O_2830,N_24890,N_23989);
xnor UO_2831 (O_2831,N_23863,N_24096);
nand UO_2832 (O_2832,N_23763,N_24536);
or UO_2833 (O_2833,N_23987,N_24862);
nor UO_2834 (O_2834,N_24656,N_24040);
and UO_2835 (O_2835,N_23934,N_23905);
or UO_2836 (O_2836,N_23801,N_24457);
nand UO_2837 (O_2837,N_24832,N_24942);
nor UO_2838 (O_2838,N_24403,N_24331);
nor UO_2839 (O_2839,N_24009,N_23812);
xnor UO_2840 (O_2840,N_24091,N_23992);
and UO_2841 (O_2841,N_24289,N_23803);
or UO_2842 (O_2842,N_24971,N_23820);
nor UO_2843 (O_2843,N_24661,N_24197);
and UO_2844 (O_2844,N_24506,N_24110);
or UO_2845 (O_2845,N_24865,N_23921);
nor UO_2846 (O_2846,N_24525,N_24474);
nor UO_2847 (O_2847,N_24747,N_24484);
nand UO_2848 (O_2848,N_24738,N_24915);
xnor UO_2849 (O_2849,N_24616,N_23952);
and UO_2850 (O_2850,N_24183,N_24857);
nor UO_2851 (O_2851,N_24165,N_24551);
xor UO_2852 (O_2852,N_23905,N_23914);
nand UO_2853 (O_2853,N_24252,N_24637);
nor UO_2854 (O_2854,N_23965,N_24501);
xor UO_2855 (O_2855,N_24125,N_24909);
xor UO_2856 (O_2856,N_24827,N_24478);
xnor UO_2857 (O_2857,N_24763,N_24452);
nand UO_2858 (O_2858,N_23881,N_24160);
and UO_2859 (O_2859,N_24436,N_24883);
or UO_2860 (O_2860,N_24773,N_24292);
nor UO_2861 (O_2861,N_23792,N_24968);
nand UO_2862 (O_2862,N_24092,N_24516);
nand UO_2863 (O_2863,N_24703,N_24362);
nor UO_2864 (O_2864,N_24429,N_24211);
and UO_2865 (O_2865,N_24791,N_24806);
or UO_2866 (O_2866,N_23952,N_24587);
nor UO_2867 (O_2867,N_24840,N_24365);
and UO_2868 (O_2868,N_24323,N_24417);
nor UO_2869 (O_2869,N_24999,N_24889);
nor UO_2870 (O_2870,N_23844,N_24172);
xor UO_2871 (O_2871,N_24622,N_24552);
and UO_2872 (O_2872,N_24610,N_24530);
or UO_2873 (O_2873,N_24118,N_24639);
xnor UO_2874 (O_2874,N_24949,N_23886);
nor UO_2875 (O_2875,N_24370,N_23781);
or UO_2876 (O_2876,N_24094,N_23915);
xor UO_2877 (O_2877,N_24161,N_23939);
nor UO_2878 (O_2878,N_24592,N_23970);
xor UO_2879 (O_2879,N_24714,N_24899);
or UO_2880 (O_2880,N_24858,N_24040);
or UO_2881 (O_2881,N_24529,N_23921);
nor UO_2882 (O_2882,N_24588,N_24817);
nor UO_2883 (O_2883,N_24846,N_24714);
xnor UO_2884 (O_2884,N_24903,N_24676);
xor UO_2885 (O_2885,N_24236,N_24480);
xor UO_2886 (O_2886,N_24083,N_24296);
nand UO_2887 (O_2887,N_24234,N_24594);
nor UO_2888 (O_2888,N_24859,N_24894);
and UO_2889 (O_2889,N_24345,N_24383);
nor UO_2890 (O_2890,N_24951,N_24664);
xnor UO_2891 (O_2891,N_24831,N_24586);
and UO_2892 (O_2892,N_24176,N_24720);
and UO_2893 (O_2893,N_24842,N_23880);
xor UO_2894 (O_2894,N_24304,N_24972);
xnor UO_2895 (O_2895,N_24649,N_24906);
or UO_2896 (O_2896,N_24107,N_24778);
and UO_2897 (O_2897,N_24219,N_24708);
and UO_2898 (O_2898,N_23751,N_24760);
xnor UO_2899 (O_2899,N_24825,N_24689);
and UO_2900 (O_2900,N_24085,N_24079);
nor UO_2901 (O_2901,N_23952,N_24154);
nor UO_2902 (O_2902,N_24045,N_24392);
or UO_2903 (O_2903,N_24835,N_23784);
or UO_2904 (O_2904,N_24586,N_24638);
xnor UO_2905 (O_2905,N_23810,N_24824);
and UO_2906 (O_2906,N_24266,N_24013);
xor UO_2907 (O_2907,N_24840,N_24330);
xnor UO_2908 (O_2908,N_24389,N_24546);
xnor UO_2909 (O_2909,N_24392,N_23975);
nand UO_2910 (O_2910,N_24473,N_24885);
xnor UO_2911 (O_2911,N_24147,N_23986);
nand UO_2912 (O_2912,N_24601,N_24640);
nand UO_2913 (O_2913,N_24197,N_23985);
and UO_2914 (O_2914,N_24260,N_24221);
nand UO_2915 (O_2915,N_24370,N_23846);
nor UO_2916 (O_2916,N_23844,N_23957);
xor UO_2917 (O_2917,N_24153,N_24798);
or UO_2918 (O_2918,N_24244,N_24337);
nand UO_2919 (O_2919,N_24716,N_24089);
nand UO_2920 (O_2920,N_24160,N_24795);
nor UO_2921 (O_2921,N_24716,N_24554);
or UO_2922 (O_2922,N_24106,N_23911);
nand UO_2923 (O_2923,N_24811,N_24494);
xnor UO_2924 (O_2924,N_24804,N_24135);
and UO_2925 (O_2925,N_24384,N_24194);
nand UO_2926 (O_2926,N_24705,N_24289);
and UO_2927 (O_2927,N_24961,N_24639);
nand UO_2928 (O_2928,N_24685,N_24865);
xnor UO_2929 (O_2929,N_23844,N_24217);
nor UO_2930 (O_2930,N_24724,N_24928);
or UO_2931 (O_2931,N_24585,N_24036);
or UO_2932 (O_2932,N_24123,N_24470);
nand UO_2933 (O_2933,N_23978,N_24494);
nor UO_2934 (O_2934,N_24347,N_24863);
and UO_2935 (O_2935,N_24023,N_24744);
or UO_2936 (O_2936,N_23932,N_23867);
and UO_2937 (O_2937,N_24752,N_24816);
and UO_2938 (O_2938,N_23778,N_24934);
and UO_2939 (O_2939,N_23880,N_23820);
xor UO_2940 (O_2940,N_24829,N_23980);
nor UO_2941 (O_2941,N_24164,N_24762);
and UO_2942 (O_2942,N_24652,N_24640);
xnor UO_2943 (O_2943,N_24621,N_23797);
or UO_2944 (O_2944,N_24773,N_24942);
nor UO_2945 (O_2945,N_24719,N_23952);
nand UO_2946 (O_2946,N_24259,N_24084);
nor UO_2947 (O_2947,N_24007,N_24510);
nor UO_2948 (O_2948,N_23934,N_24666);
nor UO_2949 (O_2949,N_23803,N_24453);
and UO_2950 (O_2950,N_23879,N_23820);
nand UO_2951 (O_2951,N_24293,N_24228);
nor UO_2952 (O_2952,N_23865,N_23938);
nand UO_2953 (O_2953,N_24271,N_24730);
and UO_2954 (O_2954,N_24062,N_24271);
or UO_2955 (O_2955,N_24994,N_24274);
and UO_2956 (O_2956,N_23990,N_24599);
nor UO_2957 (O_2957,N_24183,N_24084);
or UO_2958 (O_2958,N_23895,N_24577);
xnor UO_2959 (O_2959,N_23811,N_24474);
or UO_2960 (O_2960,N_24636,N_24558);
nand UO_2961 (O_2961,N_23880,N_24700);
xnor UO_2962 (O_2962,N_23891,N_24656);
and UO_2963 (O_2963,N_24639,N_24285);
and UO_2964 (O_2964,N_24189,N_23782);
xor UO_2965 (O_2965,N_23846,N_24446);
and UO_2966 (O_2966,N_24259,N_23964);
and UO_2967 (O_2967,N_24960,N_24600);
or UO_2968 (O_2968,N_24845,N_24943);
xnor UO_2969 (O_2969,N_24294,N_24143);
and UO_2970 (O_2970,N_23918,N_24005);
and UO_2971 (O_2971,N_23841,N_24155);
and UO_2972 (O_2972,N_24123,N_24011);
xor UO_2973 (O_2973,N_23923,N_24026);
nor UO_2974 (O_2974,N_23845,N_23922);
or UO_2975 (O_2975,N_23761,N_24955);
and UO_2976 (O_2976,N_24246,N_24088);
and UO_2977 (O_2977,N_24118,N_24751);
nand UO_2978 (O_2978,N_24036,N_24656);
nor UO_2979 (O_2979,N_23990,N_24057);
or UO_2980 (O_2980,N_24772,N_24726);
nand UO_2981 (O_2981,N_24060,N_23799);
nor UO_2982 (O_2982,N_24917,N_24269);
or UO_2983 (O_2983,N_24552,N_24538);
nand UO_2984 (O_2984,N_24058,N_24907);
nand UO_2985 (O_2985,N_24204,N_24005);
xnor UO_2986 (O_2986,N_24799,N_24322);
or UO_2987 (O_2987,N_24999,N_24287);
nand UO_2988 (O_2988,N_24049,N_23782);
nand UO_2989 (O_2989,N_24000,N_24886);
xnor UO_2990 (O_2990,N_24224,N_24873);
nor UO_2991 (O_2991,N_24355,N_24326);
and UO_2992 (O_2992,N_24395,N_24569);
xor UO_2993 (O_2993,N_24331,N_23783);
nor UO_2994 (O_2994,N_24381,N_24241);
nor UO_2995 (O_2995,N_24474,N_23879);
and UO_2996 (O_2996,N_23886,N_24867);
xnor UO_2997 (O_2997,N_24369,N_24062);
and UO_2998 (O_2998,N_24865,N_24896);
and UO_2999 (O_2999,N_24299,N_24606);
endmodule