module basic_1000_10000_1500_4_levels_2xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999;
or U0 (N_0,In_1,In_657);
or U1 (N_1,In_794,In_685);
or U2 (N_2,In_579,In_842);
or U3 (N_3,In_783,In_379);
nor U4 (N_4,In_372,In_861);
nor U5 (N_5,In_325,In_145);
nor U6 (N_6,In_167,In_615);
and U7 (N_7,In_601,In_847);
or U8 (N_8,In_228,In_408);
nand U9 (N_9,In_7,In_698);
nor U10 (N_10,In_187,In_430);
and U11 (N_11,In_482,In_26);
or U12 (N_12,In_268,In_403);
and U13 (N_13,In_185,In_278);
nand U14 (N_14,In_581,In_911);
and U15 (N_15,In_557,In_37);
nor U16 (N_16,In_686,In_400);
and U17 (N_17,In_787,In_381);
nand U18 (N_18,In_518,In_417);
and U19 (N_19,In_376,In_186);
nor U20 (N_20,In_143,In_383);
or U21 (N_21,In_845,In_782);
and U22 (N_22,In_915,In_411);
nor U23 (N_23,In_282,In_129);
or U24 (N_24,In_62,In_933);
or U25 (N_25,In_97,In_875);
nor U26 (N_26,In_665,In_338);
nor U27 (N_27,In_548,In_814);
nand U28 (N_28,In_100,In_512);
and U29 (N_29,In_435,In_904);
or U30 (N_30,In_753,In_843);
or U31 (N_31,In_76,In_175);
nor U32 (N_32,In_336,In_350);
and U33 (N_33,In_744,In_922);
nand U34 (N_34,In_756,In_474);
or U35 (N_35,In_421,In_491);
and U36 (N_36,In_852,In_447);
or U37 (N_37,In_501,In_994);
nor U38 (N_38,In_429,In_680);
xor U39 (N_39,In_211,In_793);
or U40 (N_40,In_818,In_305);
or U41 (N_41,In_317,In_202);
nand U42 (N_42,In_469,In_738);
nor U43 (N_43,In_182,In_545);
or U44 (N_44,In_258,In_908);
nor U45 (N_45,In_356,In_266);
or U46 (N_46,In_983,In_807);
nor U47 (N_47,In_540,In_646);
and U48 (N_48,In_513,In_361);
and U49 (N_49,In_718,In_333);
and U50 (N_50,In_523,In_380);
nand U51 (N_51,In_583,In_844);
and U52 (N_52,In_197,In_878);
nor U53 (N_53,In_582,In_347);
and U54 (N_54,In_871,In_711);
nor U55 (N_55,In_757,In_624);
and U56 (N_56,In_496,In_590);
xor U57 (N_57,In_480,In_357);
and U58 (N_58,In_862,In_395);
nor U59 (N_59,In_571,In_900);
or U60 (N_60,In_728,In_355);
xor U61 (N_61,In_514,In_103);
nor U62 (N_62,In_378,In_959);
nand U63 (N_63,In_978,In_340);
xnor U64 (N_64,In_112,In_495);
nand U65 (N_65,In_633,In_54);
or U66 (N_66,In_947,In_311);
and U67 (N_67,In_882,In_731);
and U68 (N_68,In_991,In_797);
nand U69 (N_69,In_568,In_530);
or U70 (N_70,In_67,In_795);
nor U71 (N_71,In_106,In_988);
nand U72 (N_72,In_578,In_327);
or U73 (N_73,In_790,In_577);
nand U74 (N_74,In_385,In_17);
and U75 (N_75,In_640,In_763);
nand U76 (N_76,In_323,In_595);
or U77 (N_77,In_661,In_397);
or U78 (N_78,In_12,In_836);
and U79 (N_79,In_538,In_413);
nand U80 (N_80,In_606,In_257);
and U81 (N_81,In_440,In_517);
nand U82 (N_82,In_808,In_135);
nand U83 (N_83,In_260,In_954);
nor U84 (N_84,In_773,In_146);
nand U85 (N_85,In_85,In_344);
or U86 (N_86,In_774,In_527);
or U87 (N_87,In_580,In_454);
nand U88 (N_88,In_301,In_11);
or U89 (N_89,In_801,In_767);
nand U90 (N_90,In_800,In_302);
nand U91 (N_91,In_918,In_63);
nor U92 (N_92,In_286,In_910);
nor U93 (N_93,In_791,In_565);
nor U94 (N_94,In_218,In_865);
nand U95 (N_95,In_688,In_283);
and U96 (N_96,In_49,In_792);
nor U97 (N_97,In_89,In_990);
and U98 (N_98,In_93,In_53);
and U99 (N_99,In_856,In_414);
xnor U100 (N_100,In_598,In_939);
nand U101 (N_101,In_425,In_289);
and U102 (N_102,In_537,In_980);
and U103 (N_103,In_876,In_120);
or U104 (N_104,In_727,In_94);
nor U105 (N_105,In_168,In_424);
nor U106 (N_106,In_43,In_467);
nor U107 (N_107,In_860,In_901);
or U108 (N_108,In_883,In_367);
or U109 (N_109,In_236,In_764);
nand U110 (N_110,In_566,In_259);
nand U111 (N_111,In_997,In_623);
nand U112 (N_112,In_740,In_812);
nor U113 (N_113,In_310,In_872);
and U114 (N_114,In_99,In_353);
nand U115 (N_115,In_678,In_586);
and U116 (N_116,In_489,In_706);
and U117 (N_117,In_928,In_221);
nor U118 (N_118,In_976,In_499);
or U119 (N_119,In_820,In_989);
nor U120 (N_120,In_732,In_90);
nand U121 (N_121,In_511,In_897);
and U122 (N_122,In_198,In_789);
and U123 (N_123,In_359,In_230);
nand U124 (N_124,In_894,In_889);
or U125 (N_125,In_321,In_567);
and U126 (N_126,In_50,In_238);
and U127 (N_127,In_449,In_898);
nand U128 (N_128,In_734,In_377);
or U129 (N_129,In_293,In_161);
and U130 (N_130,In_451,In_374);
nor U131 (N_131,In_126,In_996);
and U132 (N_132,In_314,In_903);
or U133 (N_133,In_932,In_562);
nand U134 (N_134,In_751,In_817);
or U135 (N_135,In_243,In_895);
nor U136 (N_136,In_205,In_853);
nor U137 (N_137,In_674,In_250);
and U138 (N_138,In_927,In_949);
or U139 (N_139,In_556,In_490);
or U140 (N_140,In_504,In_365);
nand U141 (N_141,In_747,In_737);
and U142 (N_142,In_22,In_890);
nand U143 (N_143,In_925,In_475);
or U144 (N_144,In_885,In_290);
and U145 (N_145,In_761,In_341);
and U146 (N_146,In_893,In_216);
or U147 (N_147,In_609,In_368);
nor U148 (N_148,In_722,In_705);
and U149 (N_149,In_956,In_74);
or U150 (N_150,In_563,In_57);
nand U151 (N_151,In_655,In_245);
and U152 (N_152,In_448,In_470);
and U153 (N_153,In_999,In_637);
nand U154 (N_154,In_332,In_473);
nand U155 (N_155,In_735,In_799);
and U156 (N_156,In_938,In_240);
and U157 (N_157,In_673,In_522);
nor U158 (N_158,In_285,In_584);
nand U159 (N_159,In_144,In_196);
and U160 (N_160,In_140,In_950);
or U161 (N_161,In_253,In_275);
and U162 (N_162,In_329,In_941);
or U163 (N_163,In_668,In_730);
nand U164 (N_164,In_104,In_262);
and U165 (N_165,In_827,In_654);
or U166 (N_166,In_539,In_549);
nor U167 (N_167,In_546,In_47);
nand U168 (N_168,In_709,In_82);
and U169 (N_169,In_768,In_444);
or U170 (N_170,In_634,In_981);
and U171 (N_171,In_930,In_271);
nor U172 (N_172,In_973,In_252);
nand U173 (N_173,In_426,In_833);
or U174 (N_174,In_386,In_136);
nor U175 (N_175,In_739,In_46);
nand U176 (N_176,In_193,In_543);
nand U177 (N_177,In_274,In_551);
or U178 (N_178,In_977,In_445);
nor U179 (N_179,In_929,In_77);
nor U180 (N_180,In_859,In_339);
nor U181 (N_181,In_415,In_102);
nand U182 (N_182,In_651,In_36);
nor U183 (N_183,In_452,In_237);
and U184 (N_184,In_687,In_667);
nor U185 (N_185,In_92,In_535);
and U186 (N_186,In_946,In_472);
nand U187 (N_187,In_79,In_892);
nand U188 (N_188,In_707,In_916);
nand U189 (N_189,In_315,In_226);
or U190 (N_190,In_699,In_241);
nand U191 (N_191,In_128,In_117);
nor U192 (N_192,In_702,In_312);
nor U193 (N_193,In_811,In_834);
and U194 (N_194,In_868,In_460);
and U195 (N_195,In_300,In_822);
nand U196 (N_196,In_905,In_422);
or U197 (N_197,In_696,In_796);
and U198 (N_198,In_239,In_115);
and U199 (N_199,In_370,In_965);
nor U200 (N_200,In_294,In_169);
nor U201 (N_201,In_222,In_389);
nor U202 (N_202,In_715,In_78);
nand U203 (N_203,In_4,In_72);
and U204 (N_204,In_838,In_44);
or U205 (N_205,In_487,In_638);
or U206 (N_206,In_755,In_462);
nor U207 (N_207,In_635,In_724);
and U208 (N_208,In_387,In_560);
and U209 (N_209,In_453,In_199);
nand U210 (N_210,In_406,In_121);
nand U211 (N_211,In_648,In_455);
or U212 (N_212,In_249,In_779);
nor U213 (N_213,In_693,In_536);
nand U214 (N_214,In_206,In_320);
nor U215 (N_215,In_457,In_391);
nor U216 (N_216,In_388,In_91);
and U217 (N_217,In_213,In_384);
nand U218 (N_218,In_671,In_393);
nand U219 (N_219,In_131,In_488);
nand U220 (N_220,In_554,In_676);
or U221 (N_221,In_227,In_269);
or U222 (N_222,In_483,In_298);
or U223 (N_223,In_71,In_466);
and U224 (N_224,In_778,In_596);
nand U225 (N_225,In_18,In_410);
nor U226 (N_226,In_529,In_951);
nor U227 (N_227,In_645,In_124);
nand U228 (N_228,In_745,In_0);
nor U229 (N_229,In_208,In_364);
nor U230 (N_230,In_309,In_427);
or U231 (N_231,In_95,In_561);
and U232 (N_232,In_281,In_758);
and U233 (N_233,In_479,In_544);
or U234 (N_234,In_171,In_907);
and U235 (N_235,In_234,In_108);
or U236 (N_236,In_870,In_3);
nor U237 (N_237,In_974,In_653);
nand U238 (N_238,In_528,In_162);
and U239 (N_239,In_891,In_313);
or U240 (N_240,In_683,In_407);
and U241 (N_241,In_463,In_464);
and U242 (N_242,In_324,In_151);
xnor U243 (N_243,In_375,In_691);
nor U244 (N_244,In_142,In_630);
or U245 (N_245,In_247,In_178);
nor U246 (N_246,In_952,In_113);
nor U247 (N_247,In_101,In_334);
or U248 (N_248,In_975,In_316);
nand U249 (N_249,In_141,In_694);
or U250 (N_250,In_823,In_926);
nor U251 (N_251,In_593,In_41);
nor U252 (N_252,In_273,In_176);
nand U253 (N_253,In_29,In_840);
and U254 (N_254,In_179,In_815);
nand U255 (N_255,In_681,In_720);
or U256 (N_256,In_307,In_109);
or U257 (N_257,In_166,In_979);
or U258 (N_258,In_855,In_966);
nor U259 (N_259,In_498,In_899);
and U260 (N_260,In_912,In_292);
nand U261 (N_261,In_777,In_343);
nand U262 (N_262,In_960,In_231);
nand U263 (N_263,In_902,In_180);
nor U264 (N_264,In_627,In_813);
or U265 (N_265,In_215,In_442);
nand U266 (N_266,In_599,In_468);
or U267 (N_267,In_277,In_15);
and U268 (N_268,In_346,In_242);
nor U269 (N_269,In_839,In_138);
and U270 (N_270,In_158,In_888);
or U271 (N_271,In_119,In_360);
xnor U272 (N_272,In_958,In_746);
and U273 (N_273,In_992,In_957);
or U274 (N_274,In_118,In_345);
nor U275 (N_275,In_233,In_670);
nand U276 (N_276,In_366,In_851);
or U277 (N_277,In_729,In_986);
and U278 (N_278,In_98,In_848);
nand U279 (N_279,In_710,In_87);
or U280 (N_280,In_650,In_909);
and U281 (N_281,In_235,In_207);
xnor U282 (N_282,In_507,In_60);
nor U283 (N_283,In_936,In_212);
or U284 (N_284,In_214,In_219);
and U285 (N_285,In_471,In_880);
or U286 (N_286,In_114,In_485);
and U287 (N_287,In_520,In_806);
nor U288 (N_288,In_526,In_256);
xnor U289 (N_289,In_776,In_652);
and U290 (N_290,In_690,In_987);
or U291 (N_291,In_532,In_982);
and U292 (N_292,In_858,In_835);
or U293 (N_293,In_38,In_80);
or U294 (N_294,In_587,In_123);
nor U295 (N_295,In_195,In_625);
and U296 (N_296,In_420,In_461);
nor U297 (N_297,In_177,In_614);
nor U298 (N_298,In_438,In_780);
nand U299 (N_299,In_632,In_873);
nor U300 (N_300,In_267,In_358);
nand U301 (N_301,In_194,In_382);
nor U302 (N_302,In_86,In_669);
or U303 (N_303,In_945,In_255);
nor U304 (N_304,In_148,In_809);
or U305 (N_305,In_917,In_684);
nor U306 (N_306,In_644,In_84);
and U307 (N_307,In_399,In_704);
or U308 (N_308,In_749,In_409);
or U309 (N_309,In_510,In_944);
and U310 (N_310,In_953,In_433);
nand U311 (N_311,In_604,In_656);
nand U312 (N_312,In_152,In_857);
and U313 (N_313,In_304,In_884);
and U314 (N_314,In_363,In_846);
nand U315 (N_315,In_51,In_299);
and U316 (N_316,In_328,In_154);
xor U317 (N_317,In_432,In_819);
xnor U318 (N_318,In_181,In_318);
and U319 (N_319,In_502,In_766);
nand U320 (N_320,In_697,In_330);
nor U321 (N_321,In_967,In_295);
nor U322 (N_322,In_829,In_831);
and U323 (N_323,In_572,In_184);
nor U324 (N_324,In_920,In_45);
or U325 (N_325,In_431,In_133);
or U326 (N_326,In_264,In_147);
and U327 (N_327,In_810,In_866);
or U328 (N_328,In_484,In_712);
or U329 (N_329,In_209,In_30);
nand U330 (N_330,In_931,In_287);
or U331 (N_331,In_229,In_402);
nor U332 (N_332,In_984,In_284);
nor U333 (N_333,In_443,In_137);
nor U334 (N_334,In_509,In_20);
and U335 (N_335,In_19,In_352);
xnor U336 (N_336,In_937,In_547);
or U337 (N_337,In_816,In_405);
nand U338 (N_338,In_8,In_170);
nand U339 (N_339,In_626,In_594);
nor U340 (N_340,In_754,In_864);
nor U341 (N_341,In_164,In_642);
nor U342 (N_342,In_641,In_703);
and U343 (N_343,In_743,In_832);
or U344 (N_344,In_319,In_446);
nand U345 (N_345,In_963,In_879);
and U346 (N_346,In_263,In_664);
nand U347 (N_347,In_998,In_497);
nor U348 (N_348,In_428,In_486);
nor U349 (N_349,In_27,In_458);
nor U350 (N_350,In_628,In_28);
nor U351 (N_351,In_83,In_204);
and U352 (N_352,In_786,In_351);
and U353 (N_353,In_70,In_719);
or U354 (N_354,In_88,In_914);
nor U355 (N_355,In_130,In_66);
and U356 (N_356,In_224,In_759);
or U357 (N_357,In_156,In_349);
and U358 (N_358,In_701,In_660);
or U359 (N_359,In_643,In_769);
and U360 (N_360,In_303,In_476);
and U361 (N_361,In_798,In_675);
or U362 (N_362,In_75,In_585);
nand U363 (N_363,In_741,In_68);
nand U364 (N_364,In_52,In_765);
and U365 (N_365,In_564,In_962);
and U366 (N_366,In_16,In_525);
nor U367 (N_367,In_742,In_603);
or U368 (N_368,In_574,In_244);
nand U369 (N_369,In_804,In_348);
and U370 (N_370,In_830,In_576);
and U371 (N_371,In_969,In_217);
or U372 (N_372,In_760,In_968);
or U373 (N_373,In_192,In_919);
and U374 (N_374,In_553,In_172);
and U375 (N_375,In_639,In_508);
nor U376 (N_376,In_10,In_600);
nand U377 (N_377,In_401,In_516);
nand U378 (N_378,In_592,In_232);
or U379 (N_379,In_165,In_163);
or U380 (N_380,In_869,In_459);
and U381 (N_381,In_588,In_272);
and U382 (N_382,In_248,In_191);
nand U383 (N_383,In_552,In_726);
and U384 (N_384,In_770,In_608);
nand U385 (N_385,In_456,In_610);
nor U386 (N_386,In_940,In_748);
or U387 (N_387,In_506,In_31);
and U388 (N_388,In_591,In_437);
and U389 (N_389,In_478,In_296);
nor U390 (N_390,In_663,In_616);
nand U391 (N_391,In_906,In_612);
xnor U392 (N_392,In_935,In_841);
nand U393 (N_393,In_649,In_280);
and U394 (N_394,In_225,In_874);
and U395 (N_395,In_276,In_183);
nand U396 (N_396,In_270,In_921);
nand U397 (N_397,In_993,In_2);
nor U398 (N_398,In_110,In_73);
or U399 (N_399,In_826,In_629);
xor U400 (N_400,In_788,In_541);
nor U401 (N_401,In_725,In_404);
nor U402 (N_402,In_708,In_23);
or U403 (N_403,In_200,In_342);
and U404 (N_404,In_394,In_33);
and U405 (N_405,In_995,In_13);
or U406 (N_406,In_56,In_493);
and U407 (N_407,In_771,In_390);
or U408 (N_408,In_961,In_679);
and U409 (N_409,In_700,In_972);
nand U410 (N_410,In_854,In_534);
nand U411 (N_411,In_531,In_828);
or U412 (N_412,In_619,In_210);
nor U413 (N_413,In_721,In_896);
or U414 (N_414,In_436,In_418);
nand U415 (N_415,In_803,In_647);
and U416 (N_416,In_441,In_542);
or U417 (N_417,In_306,In_40);
or U418 (N_418,In_602,In_943);
nor U419 (N_419,In_331,In_775);
and U420 (N_420,In_105,In_188);
or U421 (N_421,In_419,In_613);
nor U422 (N_422,In_21,In_335);
nor U423 (N_423,In_481,In_736);
or U424 (N_424,In_555,In_689);
and U425 (N_425,In_558,In_573);
or U426 (N_426,In_713,In_308);
and U427 (N_427,In_631,In_850);
and U428 (N_428,In_666,In_14);
xor U429 (N_429,In_107,In_521);
or U430 (N_430,In_533,In_201);
and U431 (N_431,In_173,In_750);
and U432 (N_432,In_867,In_5);
nor U433 (N_433,In_849,In_326);
nand U434 (N_434,In_662,In_265);
nor U435 (N_435,In_189,In_570);
or U436 (N_436,In_971,In_524);
and U437 (N_437,In_416,In_622);
nor U438 (N_438,In_772,In_61);
and U439 (N_439,In_886,In_494);
nor U440 (N_440,In_220,In_157);
nor U441 (N_441,In_695,In_423);
nor U442 (N_442,In_9,In_64);
and U443 (N_443,In_223,In_677);
or U444 (N_444,In_781,In_559);
and U445 (N_445,In_948,In_439);
nor U446 (N_446,In_762,In_913);
or U447 (N_447,In_519,In_716);
nor U448 (N_448,In_59,In_934);
nor U449 (N_449,In_492,In_254);
nor U450 (N_450,In_34,In_337);
nor U451 (N_451,In_618,In_733);
nand U452 (N_452,In_174,In_837);
or U453 (N_453,In_159,In_69);
or U454 (N_454,In_605,In_32);
nand U455 (N_455,In_877,In_251);
or U456 (N_456,In_6,In_150);
nand U457 (N_457,In_122,In_132);
xnor U458 (N_458,In_160,In_515);
nor U459 (N_459,In_39,In_964);
nor U460 (N_460,In_785,In_203);
nor U461 (N_461,In_682,In_597);
and U462 (N_462,In_139,In_297);
and U463 (N_463,In_288,In_279);
nand U464 (N_464,In_24,In_714);
and U465 (N_465,In_881,In_127);
nand U466 (N_466,In_116,In_717);
nand U467 (N_467,In_620,In_134);
or U468 (N_468,In_149,In_569);
nand U469 (N_469,In_412,In_291);
nor U470 (N_470,In_500,In_955);
or U471 (N_471,In_465,In_111);
nor U472 (N_472,In_924,In_322);
nand U473 (N_473,In_450,In_802);
nor U474 (N_474,In_261,In_723);
nand U475 (N_475,In_550,In_369);
or U476 (N_476,In_659,In_81);
nor U477 (N_477,In_672,In_636);
and U478 (N_478,In_617,In_589);
nor U479 (N_479,In_503,In_887);
and U480 (N_480,In_434,In_65);
nand U481 (N_481,In_658,In_575);
nor U482 (N_482,In_863,In_362);
and U483 (N_483,In_396,In_985);
xor U484 (N_484,In_692,In_373);
nor U485 (N_485,In_923,In_155);
or U486 (N_486,In_190,In_611);
nor U487 (N_487,In_805,In_621);
and U488 (N_488,In_55,In_477);
nand U489 (N_489,In_58,In_942);
or U490 (N_490,In_505,In_35);
nand U491 (N_491,In_25,In_371);
and U492 (N_492,In_96,In_48);
nand U493 (N_493,In_824,In_246);
or U494 (N_494,In_821,In_392);
nand U495 (N_495,In_752,In_153);
and U496 (N_496,In_607,In_398);
or U497 (N_497,In_825,In_125);
and U498 (N_498,In_784,In_970);
nor U499 (N_499,In_42,In_354);
and U500 (N_500,In_944,In_992);
or U501 (N_501,In_525,In_977);
or U502 (N_502,In_720,In_805);
xor U503 (N_503,In_25,In_134);
nand U504 (N_504,In_342,In_332);
or U505 (N_505,In_327,In_954);
nor U506 (N_506,In_970,In_900);
nor U507 (N_507,In_132,In_779);
nor U508 (N_508,In_978,In_369);
nand U509 (N_509,In_656,In_893);
and U510 (N_510,In_947,In_117);
nand U511 (N_511,In_524,In_658);
xor U512 (N_512,In_723,In_470);
or U513 (N_513,In_948,In_888);
nor U514 (N_514,In_495,In_382);
nand U515 (N_515,In_275,In_313);
or U516 (N_516,In_329,In_362);
nor U517 (N_517,In_792,In_409);
nor U518 (N_518,In_726,In_697);
or U519 (N_519,In_201,In_622);
or U520 (N_520,In_53,In_256);
and U521 (N_521,In_656,In_727);
nor U522 (N_522,In_987,In_641);
nor U523 (N_523,In_47,In_365);
nand U524 (N_524,In_725,In_221);
nand U525 (N_525,In_404,In_93);
and U526 (N_526,In_146,In_672);
or U527 (N_527,In_982,In_181);
and U528 (N_528,In_671,In_478);
and U529 (N_529,In_722,In_63);
and U530 (N_530,In_680,In_839);
and U531 (N_531,In_576,In_731);
and U532 (N_532,In_897,In_682);
nor U533 (N_533,In_878,In_350);
and U534 (N_534,In_404,In_209);
and U535 (N_535,In_947,In_557);
xnor U536 (N_536,In_264,In_196);
xor U537 (N_537,In_114,In_146);
or U538 (N_538,In_973,In_828);
nor U539 (N_539,In_704,In_451);
nand U540 (N_540,In_330,In_91);
nand U541 (N_541,In_408,In_296);
or U542 (N_542,In_154,In_967);
and U543 (N_543,In_129,In_377);
nor U544 (N_544,In_280,In_920);
and U545 (N_545,In_698,In_210);
or U546 (N_546,In_87,In_851);
nand U547 (N_547,In_606,In_174);
and U548 (N_548,In_241,In_860);
or U549 (N_549,In_661,In_468);
nor U550 (N_550,In_869,In_617);
nand U551 (N_551,In_136,In_765);
nor U552 (N_552,In_292,In_197);
and U553 (N_553,In_283,In_292);
or U554 (N_554,In_854,In_786);
nand U555 (N_555,In_153,In_57);
and U556 (N_556,In_305,In_724);
nor U557 (N_557,In_535,In_892);
and U558 (N_558,In_510,In_680);
nor U559 (N_559,In_430,In_889);
nand U560 (N_560,In_565,In_129);
and U561 (N_561,In_957,In_738);
nor U562 (N_562,In_770,In_607);
nor U563 (N_563,In_652,In_182);
nor U564 (N_564,In_672,In_742);
or U565 (N_565,In_615,In_900);
or U566 (N_566,In_299,In_478);
nor U567 (N_567,In_588,In_624);
or U568 (N_568,In_55,In_495);
and U569 (N_569,In_821,In_487);
and U570 (N_570,In_354,In_635);
and U571 (N_571,In_899,In_304);
or U572 (N_572,In_316,In_678);
nor U573 (N_573,In_577,In_938);
nor U574 (N_574,In_44,In_221);
nand U575 (N_575,In_575,In_496);
nor U576 (N_576,In_359,In_336);
nand U577 (N_577,In_245,In_182);
or U578 (N_578,In_969,In_370);
and U579 (N_579,In_205,In_410);
or U580 (N_580,In_551,In_862);
or U581 (N_581,In_833,In_876);
xor U582 (N_582,In_312,In_157);
nand U583 (N_583,In_656,In_855);
nand U584 (N_584,In_493,In_384);
and U585 (N_585,In_178,In_653);
or U586 (N_586,In_749,In_425);
and U587 (N_587,In_355,In_923);
xnor U588 (N_588,In_315,In_79);
nand U589 (N_589,In_463,In_745);
nand U590 (N_590,In_291,In_306);
or U591 (N_591,In_700,In_863);
and U592 (N_592,In_158,In_722);
and U593 (N_593,In_665,In_704);
nor U594 (N_594,In_840,In_198);
nand U595 (N_595,In_340,In_946);
nor U596 (N_596,In_318,In_489);
nand U597 (N_597,In_255,In_819);
and U598 (N_598,In_9,In_678);
and U599 (N_599,In_753,In_711);
nor U600 (N_600,In_977,In_944);
nor U601 (N_601,In_703,In_239);
nand U602 (N_602,In_255,In_672);
nand U603 (N_603,In_78,In_242);
or U604 (N_604,In_992,In_139);
nand U605 (N_605,In_679,In_604);
nor U606 (N_606,In_107,In_130);
nand U607 (N_607,In_983,In_955);
or U608 (N_608,In_323,In_708);
nand U609 (N_609,In_18,In_137);
nand U610 (N_610,In_506,In_687);
nand U611 (N_611,In_863,In_466);
nor U612 (N_612,In_550,In_528);
nand U613 (N_613,In_473,In_175);
nand U614 (N_614,In_737,In_663);
xnor U615 (N_615,In_61,In_441);
nand U616 (N_616,In_359,In_198);
or U617 (N_617,In_980,In_961);
or U618 (N_618,In_632,In_365);
or U619 (N_619,In_123,In_793);
or U620 (N_620,In_470,In_267);
and U621 (N_621,In_579,In_516);
nor U622 (N_622,In_770,In_847);
and U623 (N_623,In_44,In_947);
or U624 (N_624,In_893,In_518);
nand U625 (N_625,In_869,In_24);
nor U626 (N_626,In_136,In_31);
or U627 (N_627,In_948,In_277);
nand U628 (N_628,In_482,In_354);
or U629 (N_629,In_227,In_167);
nor U630 (N_630,In_580,In_824);
or U631 (N_631,In_927,In_287);
nor U632 (N_632,In_703,In_105);
or U633 (N_633,In_793,In_624);
xnor U634 (N_634,In_104,In_426);
and U635 (N_635,In_939,In_628);
nor U636 (N_636,In_397,In_743);
and U637 (N_637,In_202,In_533);
and U638 (N_638,In_849,In_616);
nor U639 (N_639,In_619,In_705);
and U640 (N_640,In_444,In_402);
nor U641 (N_641,In_684,In_170);
nand U642 (N_642,In_956,In_611);
nand U643 (N_643,In_994,In_978);
nor U644 (N_644,In_728,In_961);
nand U645 (N_645,In_958,In_86);
nor U646 (N_646,In_160,In_140);
and U647 (N_647,In_832,In_612);
or U648 (N_648,In_806,In_841);
or U649 (N_649,In_644,In_404);
or U650 (N_650,In_485,In_969);
or U651 (N_651,In_668,In_15);
or U652 (N_652,In_924,In_729);
and U653 (N_653,In_901,In_159);
nor U654 (N_654,In_971,In_12);
nand U655 (N_655,In_724,In_955);
nor U656 (N_656,In_377,In_849);
nand U657 (N_657,In_529,In_177);
nor U658 (N_658,In_974,In_577);
nor U659 (N_659,In_393,In_673);
nand U660 (N_660,In_191,In_581);
nand U661 (N_661,In_494,In_73);
or U662 (N_662,In_909,In_986);
or U663 (N_663,In_549,In_427);
nor U664 (N_664,In_930,In_239);
and U665 (N_665,In_393,In_433);
or U666 (N_666,In_219,In_203);
xnor U667 (N_667,In_359,In_347);
and U668 (N_668,In_225,In_488);
or U669 (N_669,In_695,In_561);
nor U670 (N_670,In_409,In_655);
and U671 (N_671,In_466,In_854);
xnor U672 (N_672,In_819,In_127);
and U673 (N_673,In_302,In_681);
nor U674 (N_674,In_719,In_131);
or U675 (N_675,In_577,In_338);
nand U676 (N_676,In_821,In_542);
and U677 (N_677,In_730,In_435);
and U678 (N_678,In_196,In_732);
or U679 (N_679,In_356,In_91);
and U680 (N_680,In_978,In_276);
nand U681 (N_681,In_274,In_839);
and U682 (N_682,In_934,In_755);
and U683 (N_683,In_897,In_838);
nand U684 (N_684,In_210,In_152);
nand U685 (N_685,In_294,In_966);
nand U686 (N_686,In_934,In_639);
and U687 (N_687,In_904,In_893);
nor U688 (N_688,In_751,In_858);
nor U689 (N_689,In_762,In_920);
nor U690 (N_690,In_370,In_477);
nor U691 (N_691,In_580,In_688);
nand U692 (N_692,In_75,In_937);
nor U693 (N_693,In_416,In_474);
and U694 (N_694,In_928,In_453);
nand U695 (N_695,In_955,In_329);
nor U696 (N_696,In_279,In_654);
nand U697 (N_697,In_39,In_584);
nand U698 (N_698,In_203,In_727);
or U699 (N_699,In_644,In_269);
nor U700 (N_700,In_786,In_634);
nor U701 (N_701,In_666,In_305);
and U702 (N_702,In_101,In_566);
and U703 (N_703,In_203,In_516);
nand U704 (N_704,In_777,In_615);
and U705 (N_705,In_76,In_439);
and U706 (N_706,In_335,In_501);
nor U707 (N_707,In_747,In_443);
nand U708 (N_708,In_959,In_481);
or U709 (N_709,In_499,In_880);
or U710 (N_710,In_856,In_530);
nor U711 (N_711,In_766,In_950);
nor U712 (N_712,In_272,In_381);
nor U713 (N_713,In_350,In_659);
xnor U714 (N_714,In_764,In_700);
and U715 (N_715,In_836,In_513);
and U716 (N_716,In_107,In_138);
nand U717 (N_717,In_451,In_802);
or U718 (N_718,In_322,In_723);
or U719 (N_719,In_729,In_363);
and U720 (N_720,In_30,In_192);
nor U721 (N_721,In_591,In_977);
nor U722 (N_722,In_983,In_589);
nand U723 (N_723,In_677,In_991);
nor U724 (N_724,In_337,In_197);
and U725 (N_725,In_160,In_646);
nor U726 (N_726,In_624,In_42);
and U727 (N_727,In_246,In_588);
nand U728 (N_728,In_770,In_166);
and U729 (N_729,In_603,In_561);
nor U730 (N_730,In_667,In_526);
nand U731 (N_731,In_729,In_482);
xnor U732 (N_732,In_41,In_537);
or U733 (N_733,In_268,In_371);
nor U734 (N_734,In_356,In_938);
nand U735 (N_735,In_408,In_390);
nor U736 (N_736,In_647,In_673);
nand U737 (N_737,In_660,In_433);
nand U738 (N_738,In_147,In_268);
or U739 (N_739,In_940,In_90);
and U740 (N_740,In_201,In_912);
nand U741 (N_741,In_379,In_822);
and U742 (N_742,In_221,In_752);
and U743 (N_743,In_875,In_264);
and U744 (N_744,In_670,In_657);
or U745 (N_745,In_414,In_500);
or U746 (N_746,In_291,In_152);
or U747 (N_747,In_153,In_786);
and U748 (N_748,In_852,In_958);
or U749 (N_749,In_546,In_658);
nor U750 (N_750,In_339,In_600);
and U751 (N_751,In_522,In_175);
nor U752 (N_752,In_224,In_890);
nor U753 (N_753,In_467,In_642);
and U754 (N_754,In_596,In_241);
or U755 (N_755,In_332,In_752);
nor U756 (N_756,In_887,In_788);
or U757 (N_757,In_599,In_191);
nand U758 (N_758,In_508,In_989);
nor U759 (N_759,In_299,In_313);
nand U760 (N_760,In_726,In_55);
or U761 (N_761,In_900,In_604);
and U762 (N_762,In_610,In_281);
nor U763 (N_763,In_449,In_190);
or U764 (N_764,In_702,In_623);
nor U765 (N_765,In_795,In_911);
nand U766 (N_766,In_743,In_686);
nor U767 (N_767,In_793,In_509);
and U768 (N_768,In_160,In_684);
nand U769 (N_769,In_386,In_535);
nand U770 (N_770,In_242,In_304);
and U771 (N_771,In_394,In_676);
nor U772 (N_772,In_968,In_42);
and U773 (N_773,In_439,In_990);
nor U774 (N_774,In_687,In_663);
nor U775 (N_775,In_657,In_601);
and U776 (N_776,In_970,In_867);
nor U777 (N_777,In_543,In_404);
and U778 (N_778,In_847,In_364);
and U779 (N_779,In_961,In_104);
and U780 (N_780,In_593,In_505);
nand U781 (N_781,In_572,In_266);
and U782 (N_782,In_683,In_365);
or U783 (N_783,In_336,In_681);
or U784 (N_784,In_103,In_27);
or U785 (N_785,In_610,In_551);
nor U786 (N_786,In_385,In_522);
and U787 (N_787,In_142,In_737);
nand U788 (N_788,In_674,In_182);
or U789 (N_789,In_19,In_804);
nor U790 (N_790,In_534,In_504);
nand U791 (N_791,In_569,In_238);
nor U792 (N_792,In_84,In_59);
nand U793 (N_793,In_344,In_345);
nor U794 (N_794,In_426,In_619);
or U795 (N_795,In_535,In_505);
or U796 (N_796,In_665,In_373);
nor U797 (N_797,In_207,In_567);
nor U798 (N_798,In_585,In_317);
and U799 (N_799,In_284,In_72);
nand U800 (N_800,In_554,In_289);
or U801 (N_801,In_931,In_317);
nand U802 (N_802,In_74,In_283);
nor U803 (N_803,In_242,In_669);
nand U804 (N_804,In_560,In_521);
or U805 (N_805,In_911,In_269);
or U806 (N_806,In_328,In_781);
nor U807 (N_807,In_6,In_45);
nand U808 (N_808,In_539,In_975);
and U809 (N_809,In_947,In_98);
nand U810 (N_810,In_740,In_211);
and U811 (N_811,In_675,In_808);
nor U812 (N_812,In_462,In_1);
and U813 (N_813,In_35,In_158);
nand U814 (N_814,In_711,In_624);
nor U815 (N_815,In_730,In_676);
or U816 (N_816,In_741,In_461);
nor U817 (N_817,In_125,In_565);
xor U818 (N_818,In_704,In_241);
or U819 (N_819,In_748,In_284);
or U820 (N_820,In_784,In_928);
or U821 (N_821,In_825,In_455);
nor U822 (N_822,In_786,In_497);
or U823 (N_823,In_575,In_85);
nand U824 (N_824,In_746,In_886);
and U825 (N_825,In_570,In_757);
or U826 (N_826,In_661,In_505);
or U827 (N_827,In_283,In_209);
nor U828 (N_828,In_723,In_9);
and U829 (N_829,In_602,In_424);
xnor U830 (N_830,In_981,In_149);
nand U831 (N_831,In_791,In_557);
nor U832 (N_832,In_990,In_574);
nor U833 (N_833,In_312,In_370);
nand U834 (N_834,In_648,In_728);
nand U835 (N_835,In_689,In_426);
nor U836 (N_836,In_861,In_163);
nor U837 (N_837,In_438,In_40);
or U838 (N_838,In_139,In_315);
xnor U839 (N_839,In_831,In_827);
nand U840 (N_840,In_105,In_15);
and U841 (N_841,In_576,In_792);
nand U842 (N_842,In_714,In_279);
nand U843 (N_843,In_427,In_307);
and U844 (N_844,In_28,In_876);
nor U845 (N_845,In_561,In_612);
and U846 (N_846,In_453,In_628);
and U847 (N_847,In_328,In_347);
and U848 (N_848,In_557,In_276);
nand U849 (N_849,In_777,In_680);
nand U850 (N_850,In_426,In_205);
nor U851 (N_851,In_991,In_803);
or U852 (N_852,In_571,In_521);
xor U853 (N_853,In_259,In_529);
and U854 (N_854,In_727,In_604);
or U855 (N_855,In_695,In_31);
nand U856 (N_856,In_978,In_750);
and U857 (N_857,In_345,In_376);
or U858 (N_858,In_54,In_884);
nand U859 (N_859,In_633,In_904);
and U860 (N_860,In_923,In_723);
or U861 (N_861,In_872,In_679);
nor U862 (N_862,In_763,In_256);
and U863 (N_863,In_191,In_697);
nor U864 (N_864,In_425,In_671);
nand U865 (N_865,In_848,In_63);
and U866 (N_866,In_428,In_157);
and U867 (N_867,In_339,In_521);
or U868 (N_868,In_62,In_720);
or U869 (N_869,In_387,In_805);
nand U870 (N_870,In_390,In_702);
nor U871 (N_871,In_443,In_797);
or U872 (N_872,In_802,In_62);
nand U873 (N_873,In_272,In_546);
and U874 (N_874,In_899,In_785);
or U875 (N_875,In_56,In_540);
nand U876 (N_876,In_820,In_872);
or U877 (N_877,In_389,In_679);
and U878 (N_878,In_701,In_72);
and U879 (N_879,In_465,In_729);
and U880 (N_880,In_709,In_470);
xor U881 (N_881,In_787,In_190);
and U882 (N_882,In_533,In_627);
nand U883 (N_883,In_896,In_25);
and U884 (N_884,In_355,In_597);
nand U885 (N_885,In_140,In_206);
and U886 (N_886,In_452,In_868);
nand U887 (N_887,In_783,In_426);
or U888 (N_888,In_749,In_785);
nor U889 (N_889,In_417,In_480);
and U890 (N_890,In_854,In_444);
and U891 (N_891,In_463,In_746);
nand U892 (N_892,In_297,In_586);
nand U893 (N_893,In_14,In_692);
nor U894 (N_894,In_574,In_625);
nor U895 (N_895,In_364,In_130);
nor U896 (N_896,In_906,In_149);
and U897 (N_897,In_212,In_558);
nor U898 (N_898,In_706,In_685);
or U899 (N_899,In_32,In_884);
and U900 (N_900,In_0,In_79);
or U901 (N_901,In_401,In_474);
and U902 (N_902,In_562,In_366);
or U903 (N_903,In_379,In_603);
and U904 (N_904,In_568,In_777);
and U905 (N_905,In_256,In_63);
xor U906 (N_906,In_269,In_149);
and U907 (N_907,In_186,In_825);
or U908 (N_908,In_955,In_665);
nor U909 (N_909,In_646,In_412);
nand U910 (N_910,In_487,In_513);
nand U911 (N_911,In_993,In_143);
nand U912 (N_912,In_697,In_822);
and U913 (N_913,In_555,In_720);
and U914 (N_914,In_117,In_549);
nor U915 (N_915,In_8,In_679);
nand U916 (N_916,In_854,In_188);
nor U917 (N_917,In_403,In_81);
nand U918 (N_918,In_344,In_465);
nand U919 (N_919,In_666,In_8);
nor U920 (N_920,In_36,In_38);
nand U921 (N_921,In_401,In_683);
or U922 (N_922,In_358,In_815);
nor U923 (N_923,In_916,In_663);
nor U924 (N_924,In_730,In_509);
nand U925 (N_925,In_510,In_791);
nor U926 (N_926,In_256,In_338);
nor U927 (N_927,In_634,In_979);
nor U928 (N_928,In_164,In_610);
or U929 (N_929,In_443,In_557);
nor U930 (N_930,In_96,In_67);
or U931 (N_931,In_585,In_423);
nand U932 (N_932,In_919,In_933);
nor U933 (N_933,In_871,In_156);
and U934 (N_934,In_178,In_552);
nand U935 (N_935,In_328,In_767);
nand U936 (N_936,In_695,In_250);
nor U937 (N_937,In_403,In_486);
or U938 (N_938,In_492,In_689);
or U939 (N_939,In_39,In_549);
nand U940 (N_940,In_760,In_436);
nand U941 (N_941,In_0,In_246);
and U942 (N_942,In_122,In_2);
nor U943 (N_943,In_622,In_915);
nand U944 (N_944,In_737,In_326);
nand U945 (N_945,In_984,In_23);
and U946 (N_946,In_390,In_763);
nor U947 (N_947,In_680,In_566);
and U948 (N_948,In_771,In_167);
nand U949 (N_949,In_402,In_690);
or U950 (N_950,In_635,In_412);
nor U951 (N_951,In_559,In_114);
xnor U952 (N_952,In_176,In_290);
and U953 (N_953,In_616,In_701);
nand U954 (N_954,In_228,In_415);
or U955 (N_955,In_993,In_612);
nor U956 (N_956,In_213,In_0);
nor U957 (N_957,In_816,In_296);
nand U958 (N_958,In_152,In_525);
xnor U959 (N_959,In_658,In_592);
nand U960 (N_960,In_312,In_736);
and U961 (N_961,In_352,In_305);
or U962 (N_962,In_636,In_534);
or U963 (N_963,In_115,In_302);
nand U964 (N_964,In_846,In_171);
or U965 (N_965,In_269,In_73);
and U966 (N_966,In_246,In_802);
and U967 (N_967,In_651,In_947);
xor U968 (N_968,In_176,In_77);
nor U969 (N_969,In_735,In_260);
nand U970 (N_970,In_337,In_73);
nand U971 (N_971,In_541,In_492);
nor U972 (N_972,In_876,In_515);
nand U973 (N_973,In_555,In_900);
and U974 (N_974,In_81,In_520);
nor U975 (N_975,In_843,In_779);
nor U976 (N_976,In_60,In_114);
and U977 (N_977,In_87,In_325);
or U978 (N_978,In_743,In_370);
and U979 (N_979,In_382,In_157);
and U980 (N_980,In_739,In_346);
nor U981 (N_981,In_925,In_773);
nand U982 (N_982,In_813,In_389);
and U983 (N_983,In_833,In_655);
nor U984 (N_984,In_752,In_689);
nor U985 (N_985,In_216,In_56);
nor U986 (N_986,In_371,In_367);
and U987 (N_987,In_459,In_695);
nor U988 (N_988,In_380,In_531);
nor U989 (N_989,In_220,In_353);
or U990 (N_990,In_457,In_447);
and U991 (N_991,In_541,In_224);
nor U992 (N_992,In_167,In_442);
nor U993 (N_993,In_71,In_751);
nor U994 (N_994,In_762,In_928);
or U995 (N_995,In_616,In_994);
nor U996 (N_996,In_132,In_633);
nor U997 (N_997,In_958,In_308);
nor U998 (N_998,In_705,In_134);
and U999 (N_999,In_35,In_541);
nand U1000 (N_1000,In_24,In_327);
or U1001 (N_1001,In_689,In_815);
nor U1002 (N_1002,In_814,In_316);
or U1003 (N_1003,In_853,In_688);
nand U1004 (N_1004,In_332,In_949);
nor U1005 (N_1005,In_81,In_951);
and U1006 (N_1006,In_553,In_396);
and U1007 (N_1007,In_267,In_713);
and U1008 (N_1008,In_3,In_753);
or U1009 (N_1009,In_114,In_975);
nand U1010 (N_1010,In_808,In_74);
and U1011 (N_1011,In_292,In_759);
or U1012 (N_1012,In_471,In_911);
nand U1013 (N_1013,In_944,In_9);
nand U1014 (N_1014,In_394,In_668);
or U1015 (N_1015,In_451,In_280);
nand U1016 (N_1016,In_76,In_701);
and U1017 (N_1017,In_459,In_680);
nor U1018 (N_1018,In_610,In_950);
nor U1019 (N_1019,In_835,In_200);
and U1020 (N_1020,In_9,In_396);
and U1021 (N_1021,In_837,In_43);
or U1022 (N_1022,In_734,In_548);
or U1023 (N_1023,In_609,In_583);
nand U1024 (N_1024,In_959,In_767);
or U1025 (N_1025,In_261,In_414);
and U1026 (N_1026,In_747,In_639);
and U1027 (N_1027,In_453,In_621);
nor U1028 (N_1028,In_415,In_705);
nor U1029 (N_1029,In_162,In_226);
nor U1030 (N_1030,In_717,In_229);
or U1031 (N_1031,In_594,In_151);
nor U1032 (N_1032,In_862,In_761);
and U1033 (N_1033,In_900,In_754);
and U1034 (N_1034,In_841,In_191);
nor U1035 (N_1035,In_959,In_542);
and U1036 (N_1036,In_419,In_396);
nor U1037 (N_1037,In_484,In_754);
nor U1038 (N_1038,In_961,In_167);
nand U1039 (N_1039,In_639,In_77);
nor U1040 (N_1040,In_783,In_208);
or U1041 (N_1041,In_744,In_72);
nor U1042 (N_1042,In_619,In_425);
nand U1043 (N_1043,In_693,In_735);
nand U1044 (N_1044,In_648,In_619);
and U1045 (N_1045,In_219,In_211);
nor U1046 (N_1046,In_57,In_954);
xor U1047 (N_1047,In_573,In_261);
and U1048 (N_1048,In_505,In_791);
or U1049 (N_1049,In_961,In_895);
nand U1050 (N_1050,In_959,In_75);
or U1051 (N_1051,In_107,In_690);
and U1052 (N_1052,In_255,In_273);
and U1053 (N_1053,In_979,In_860);
or U1054 (N_1054,In_33,In_135);
or U1055 (N_1055,In_795,In_267);
and U1056 (N_1056,In_783,In_814);
and U1057 (N_1057,In_549,In_713);
nand U1058 (N_1058,In_223,In_33);
or U1059 (N_1059,In_657,In_638);
nand U1060 (N_1060,In_362,In_281);
or U1061 (N_1061,In_106,In_55);
nand U1062 (N_1062,In_199,In_94);
nor U1063 (N_1063,In_867,In_490);
or U1064 (N_1064,In_897,In_730);
or U1065 (N_1065,In_64,In_25);
and U1066 (N_1066,In_85,In_219);
and U1067 (N_1067,In_703,In_798);
and U1068 (N_1068,In_928,In_76);
nor U1069 (N_1069,In_857,In_552);
nand U1070 (N_1070,In_524,In_492);
nand U1071 (N_1071,In_904,In_775);
and U1072 (N_1072,In_57,In_271);
and U1073 (N_1073,In_747,In_877);
or U1074 (N_1074,In_453,In_634);
nor U1075 (N_1075,In_313,In_771);
nand U1076 (N_1076,In_828,In_878);
and U1077 (N_1077,In_462,In_319);
and U1078 (N_1078,In_118,In_137);
nand U1079 (N_1079,In_967,In_285);
and U1080 (N_1080,In_554,In_338);
and U1081 (N_1081,In_277,In_858);
and U1082 (N_1082,In_72,In_896);
and U1083 (N_1083,In_493,In_86);
and U1084 (N_1084,In_422,In_540);
nor U1085 (N_1085,In_292,In_717);
and U1086 (N_1086,In_1,In_616);
or U1087 (N_1087,In_638,In_869);
and U1088 (N_1088,In_524,In_945);
or U1089 (N_1089,In_383,In_821);
nand U1090 (N_1090,In_405,In_852);
nand U1091 (N_1091,In_33,In_596);
nand U1092 (N_1092,In_256,In_260);
or U1093 (N_1093,In_863,In_423);
and U1094 (N_1094,In_591,In_156);
or U1095 (N_1095,In_655,In_283);
or U1096 (N_1096,In_880,In_340);
or U1097 (N_1097,In_897,In_573);
and U1098 (N_1098,In_62,In_217);
nor U1099 (N_1099,In_38,In_808);
and U1100 (N_1100,In_590,In_585);
nand U1101 (N_1101,In_278,In_320);
nor U1102 (N_1102,In_48,In_348);
nor U1103 (N_1103,In_724,In_83);
and U1104 (N_1104,In_961,In_869);
and U1105 (N_1105,In_95,In_794);
nor U1106 (N_1106,In_617,In_248);
nor U1107 (N_1107,In_162,In_930);
and U1108 (N_1108,In_647,In_134);
or U1109 (N_1109,In_772,In_630);
or U1110 (N_1110,In_546,In_182);
and U1111 (N_1111,In_123,In_432);
or U1112 (N_1112,In_864,In_687);
and U1113 (N_1113,In_405,In_842);
and U1114 (N_1114,In_435,In_581);
nor U1115 (N_1115,In_896,In_557);
and U1116 (N_1116,In_770,In_389);
nor U1117 (N_1117,In_322,In_33);
nand U1118 (N_1118,In_468,In_643);
and U1119 (N_1119,In_995,In_902);
nor U1120 (N_1120,In_902,In_118);
or U1121 (N_1121,In_899,In_913);
nand U1122 (N_1122,In_561,In_43);
nor U1123 (N_1123,In_411,In_56);
nand U1124 (N_1124,In_497,In_212);
and U1125 (N_1125,In_67,In_101);
and U1126 (N_1126,In_655,In_684);
and U1127 (N_1127,In_548,In_956);
and U1128 (N_1128,In_667,In_820);
nor U1129 (N_1129,In_971,In_317);
nand U1130 (N_1130,In_214,In_713);
and U1131 (N_1131,In_593,In_483);
nor U1132 (N_1132,In_646,In_505);
and U1133 (N_1133,In_711,In_778);
nor U1134 (N_1134,In_201,In_578);
or U1135 (N_1135,In_74,In_560);
nand U1136 (N_1136,In_43,In_824);
nand U1137 (N_1137,In_100,In_422);
nand U1138 (N_1138,In_327,In_217);
nor U1139 (N_1139,In_546,In_860);
nor U1140 (N_1140,In_829,In_414);
nor U1141 (N_1141,In_748,In_339);
or U1142 (N_1142,In_565,In_71);
and U1143 (N_1143,In_795,In_401);
nor U1144 (N_1144,In_999,In_253);
or U1145 (N_1145,In_421,In_499);
nand U1146 (N_1146,In_626,In_258);
nor U1147 (N_1147,In_271,In_84);
and U1148 (N_1148,In_946,In_456);
nand U1149 (N_1149,In_599,In_533);
and U1150 (N_1150,In_197,In_515);
or U1151 (N_1151,In_258,In_585);
nand U1152 (N_1152,In_347,In_265);
and U1153 (N_1153,In_452,In_458);
or U1154 (N_1154,In_183,In_753);
and U1155 (N_1155,In_46,In_435);
or U1156 (N_1156,In_678,In_412);
and U1157 (N_1157,In_783,In_74);
nand U1158 (N_1158,In_929,In_760);
or U1159 (N_1159,In_290,In_750);
nor U1160 (N_1160,In_535,In_82);
and U1161 (N_1161,In_326,In_834);
nand U1162 (N_1162,In_469,In_956);
or U1163 (N_1163,In_427,In_182);
nor U1164 (N_1164,In_890,In_153);
or U1165 (N_1165,In_584,In_425);
nand U1166 (N_1166,In_604,In_501);
or U1167 (N_1167,In_836,In_170);
and U1168 (N_1168,In_646,In_661);
nor U1169 (N_1169,In_961,In_313);
nor U1170 (N_1170,In_761,In_683);
and U1171 (N_1171,In_235,In_646);
nor U1172 (N_1172,In_560,In_962);
or U1173 (N_1173,In_876,In_25);
nor U1174 (N_1174,In_241,In_315);
or U1175 (N_1175,In_803,In_567);
nand U1176 (N_1176,In_595,In_454);
and U1177 (N_1177,In_504,In_759);
nand U1178 (N_1178,In_965,In_896);
nor U1179 (N_1179,In_932,In_983);
and U1180 (N_1180,In_645,In_758);
nor U1181 (N_1181,In_837,In_581);
xnor U1182 (N_1182,In_258,In_575);
or U1183 (N_1183,In_411,In_971);
and U1184 (N_1184,In_182,In_628);
nor U1185 (N_1185,In_858,In_338);
nand U1186 (N_1186,In_291,In_761);
nand U1187 (N_1187,In_241,In_559);
nor U1188 (N_1188,In_333,In_940);
and U1189 (N_1189,In_188,In_517);
or U1190 (N_1190,In_265,In_120);
nand U1191 (N_1191,In_403,In_430);
and U1192 (N_1192,In_249,In_898);
nand U1193 (N_1193,In_695,In_662);
or U1194 (N_1194,In_447,In_602);
or U1195 (N_1195,In_297,In_868);
or U1196 (N_1196,In_330,In_706);
nor U1197 (N_1197,In_453,In_663);
nand U1198 (N_1198,In_576,In_535);
and U1199 (N_1199,In_686,In_210);
nor U1200 (N_1200,In_244,In_100);
or U1201 (N_1201,In_360,In_321);
nor U1202 (N_1202,In_820,In_273);
nor U1203 (N_1203,In_460,In_498);
and U1204 (N_1204,In_357,In_325);
xor U1205 (N_1205,In_990,In_3);
nand U1206 (N_1206,In_65,In_274);
nor U1207 (N_1207,In_804,In_214);
or U1208 (N_1208,In_979,In_568);
nor U1209 (N_1209,In_35,In_322);
nand U1210 (N_1210,In_261,In_932);
and U1211 (N_1211,In_211,In_797);
or U1212 (N_1212,In_345,In_742);
nor U1213 (N_1213,In_501,In_512);
nor U1214 (N_1214,In_156,In_268);
xnor U1215 (N_1215,In_212,In_177);
and U1216 (N_1216,In_118,In_949);
nand U1217 (N_1217,In_739,In_73);
or U1218 (N_1218,In_792,In_321);
nand U1219 (N_1219,In_943,In_476);
nor U1220 (N_1220,In_672,In_226);
or U1221 (N_1221,In_778,In_424);
or U1222 (N_1222,In_810,In_59);
nor U1223 (N_1223,In_956,In_631);
or U1224 (N_1224,In_899,In_586);
or U1225 (N_1225,In_103,In_322);
nor U1226 (N_1226,In_663,In_652);
nand U1227 (N_1227,In_851,In_490);
nand U1228 (N_1228,In_358,In_452);
or U1229 (N_1229,In_930,In_5);
or U1230 (N_1230,In_697,In_977);
nor U1231 (N_1231,In_717,In_592);
and U1232 (N_1232,In_948,In_679);
xor U1233 (N_1233,In_28,In_781);
or U1234 (N_1234,In_801,In_505);
and U1235 (N_1235,In_667,In_771);
nand U1236 (N_1236,In_791,In_63);
nor U1237 (N_1237,In_548,In_782);
nand U1238 (N_1238,In_224,In_720);
xnor U1239 (N_1239,In_154,In_934);
and U1240 (N_1240,In_362,In_923);
xnor U1241 (N_1241,In_411,In_958);
xnor U1242 (N_1242,In_845,In_921);
or U1243 (N_1243,In_42,In_909);
and U1244 (N_1244,In_382,In_313);
nand U1245 (N_1245,In_425,In_305);
nand U1246 (N_1246,In_166,In_204);
nand U1247 (N_1247,In_930,In_392);
nor U1248 (N_1248,In_481,In_722);
or U1249 (N_1249,In_111,In_426);
or U1250 (N_1250,In_771,In_373);
or U1251 (N_1251,In_531,In_146);
nand U1252 (N_1252,In_363,In_456);
nand U1253 (N_1253,In_766,In_504);
xnor U1254 (N_1254,In_374,In_246);
and U1255 (N_1255,In_101,In_949);
nand U1256 (N_1256,In_94,In_315);
or U1257 (N_1257,In_857,In_890);
nor U1258 (N_1258,In_601,In_185);
nor U1259 (N_1259,In_459,In_931);
nor U1260 (N_1260,In_758,In_200);
and U1261 (N_1261,In_904,In_507);
or U1262 (N_1262,In_65,In_935);
nand U1263 (N_1263,In_902,In_633);
or U1264 (N_1264,In_807,In_477);
or U1265 (N_1265,In_958,In_963);
or U1266 (N_1266,In_726,In_512);
and U1267 (N_1267,In_689,In_956);
and U1268 (N_1268,In_278,In_506);
and U1269 (N_1269,In_866,In_690);
nor U1270 (N_1270,In_826,In_53);
nor U1271 (N_1271,In_80,In_234);
nor U1272 (N_1272,In_219,In_590);
nor U1273 (N_1273,In_42,In_402);
nand U1274 (N_1274,In_919,In_124);
nor U1275 (N_1275,In_42,In_27);
and U1276 (N_1276,In_238,In_679);
nand U1277 (N_1277,In_923,In_64);
and U1278 (N_1278,In_977,In_716);
nor U1279 (N_1279,In_102,In_64);
nor U1280 (N_1280,In_285,In_81);
and U1281 (N_1281,In_435,In_619);
xor U1282 (N_1282,In_811,In_183);
and U1283 (N_1283,In_946,In_739);
nand U1284 (N_1284,In_813,In_409);
or U1285 (N_1285,In_150,In_254);
nor U1286 (N_1286,In_174,In_150);
xnor U1287 (N_1287,In_559,In_946);
and U1288 (N_1288,In_229,In_324);
and U1289 (N_1289,In_844,In_506);
or U1290 (N_1290,In_844,In_78);
or U1291 (N_1291,In_14,In_828);
nand U1292 (N_1292,In_565,In_131);
nand U1293 (N_1293,In_444,In_241);
nor U1294 (N_1294,In_432,In_520);
and U1295 (N_1295,In_210,In_655);
nand U1296 (N_1296,In_716,In_785);
or U1297 (N_1297,In_55,In_991);
and U1298 (N_1298,In_245,In_931);
and U1299 (N_1299,In_536,In_227);
and U1300 (N_1300,In_216,In_3);
and U1301 (N_1301,In_370,In_468);
nor U1302 (N_1302,In_495,In_928);
xor U1303 (N_1303,In_338,In_406);
nand U1304 (N_1304,In_267,In_837);
nor U1305 (N_1305,In_477,In_3);
or U1306 (N_1306,In_976,In_968);
nand U1307 (N_1307,In_491,In_837);
xor U1308 (N_1308,In_814,In_230);
nor U1309 (N_1309,In_666,In_696);
nor U1310 (N_1310,In_158,In_461);
nand U1311 (N_1311,In_896,In_307);
or U1312 (N_1312,In_660,In_669);
nor U1313 (N_1313,In_300,In_996);
nor U1314 (N_1314,In_883,In_217);
and U1315 (N_1315,In_637,In_236);
nor U1316 (N_1316,In_607,In_514);
and U1317 (N_1317,In_239,In_584);
or U1318 (N_1318,In_135,In_56);
or U1319 (N_1319,In_599,In_700);
and U1320 (N_1320,In_240,In_677);
nand U1321 (N_1321,In_101,In_521);
nor U1322 (N_1322,In_807,In_705);
or U1323 (N_1323,In_821,In_473);
nor U1324 (N_1324,In_124,In_992);
and U1325 (N_1325,In_950,In_282);
and U1326 (N_1326,In_186,In_267);
nand U1327 (N_1327,In_349,In_510);
and U1328 (N_1328,In_293,In_738);
and U1329 (N_1329,In_566,In_949);
nand U1330 (N_1330,In_143,In_687);
or U1331 (N_1331,In_576,In_721);
nand U1332 (N_1332,In_941,In_277);
nand U1333 (N_1333,In_630,In_200);
and U1334 (N_1334,In_985,In_664);
and U1335 (N_1335,In_874,In_755);
xnor U1336 (N_1336,In_257,In_143);
nand U1337 (N_1337,In_797,In_322);
nand U1338 (N_1338,In_893,In_240);
and U1339 (N_1339,In_543,In_558);
nor U1340 (N_1340,In_61,In_43);
nor U1341 (N_1341,In_185,In_939);
or U1342 (N_1342,In_913,In_903);
nand U1343 (N_1343,In_446,In_752);
nor U1344 (N_1344,In_639,In_179);
and U1345 (N_1345,In_524,In_114);
nor U1346 (N_1346,In_548,In_680);
and U1347 (N_1347,In_140,In_285);
nor U1348 (N_1348,In_917,In_244);
nor U1349 (N_1349,In_310,In_331);
or U1350 (N_1350,In_270,In_876);
nor U1351 (N_1351,In_272,In_574);
and U1352 (N_1352,In_776,In_988);
nor U1353 (N_1353,In_280,In_120);
nand U1354 (N_1354,In_505,In_820);
nor U1355 (N_1355,In_926,In_862);
nor U1356 (N_1356,In_470,In_833);
nand U1357 (N_1357,In_595,In_19);
and U1358 (N_1358,In_716,In_619);
nand U1359 (N_1359,In_29,In_576);
nand U1360 (N_1360,In_140,In_802);
nand U1361 (N_1361,In_394,In_60);
and U1362 (N_1362,In_296,In_98);
nand U1363 (N_1363,In_391,In_196);
or U1364 (N_1364,In_12,In_118);
nor U1365 (N_1365,In_626,In_701);
or U1366 (N_1366,In_398,In_854);
nand U1367 (N_1367,In_8,In_782);
nand U1368 (N_1368,In_647,In_773);
nor U1369 (N_1369,In_930,In_884);
nor U1370 (N_1370,In_842,In_433);
or U1371 (N_1371,In_665,In_943);
nor U1372 (N_1372,In_454,In_990);
or U1373 (N_1373,In_266,In_280);
and U1374 (N_1374,In_125,In_253);
or U1375 (N_1375,In_290,In_605);
and U1376 (N_1376,In_775,In_583);
and U1377 (N_1377,In_644,In_756);
and U1378 (N_1378,In_146,In_360);
and U1379 (N_1379,In_293,In_9);
or U1380 (N_1380,In_461,In_923);
and U1381 (N_1381,In_541,In_89);
nand U1382 (N_1382,In_254,In_79);
nand U1383 (N_1383,In_623,In_35);
and U1384 (N_1384,In_960,In_605);
nand U1385 (N_1385,In_25,In_651);
nor U1386 (N_1386,In_165,In_76);
or U1387 (N_1387,In_419,In_238);
nor U1388 (N_1388,In_434,In_485);
or U1389 (N_1389,In_751,In_168);
or U1390 (N_1390,In_228,In_117);
nor U1391 (N_1391,In_227,In_454);
and U1392 (N_1392,In_993,In_5);
nor U1393 (N_1393,In_534,In_40);
nand U1394 (N_1394,In_987,In_887);
or U1395 (N_1395,In_612,In_694);
nor U1396 (N_1396,In_203,In_577);
nor U1397 (N_1397,In_78,In_721);
nor U1398 (N_1398,In_467,In_753);
nor U1399 (N_1399,In_493,In_60);
nor U1400 (N_1400,In_329,In_899);
or U1401 (N_1401,In_258,In_94);
nand U1402 (N_1402,In_594,In_414);
or U1403 (N_1403,In_674,In_105);
or U1404 (N_1404,In_896,In_905);
and U1405 (N_1405,In_13,In_39);
nand U1406 (N_1406,In_661,In_517);
or U1407 (N_1407,In_979,In_605);
or U1408 (N_1408,In_435,In_749);
and U1409 (N_1409,In_722,In_252);
nor U1410 (N_1410,In_578,In_481);
or U1411 (N_1411,In_356,In_892);
or U1412 (N_1412,In_921,In_645);
or U1413 (N_1413,In_547,In_474);
or U1414 (N_1414,In_285,In_48);
nor U1415 (N_1415,In_61,In_497);
or U1416 (N_1416,In_660,In_772);
or U1417 (N_1417,In_769,In_524);
nand U1418 (N_1418,In_311,In_107);
and U1419 (N_1419,In_358,In_55);
or U1420 (N_1420,In_536,In_946);
or U1421 (N_1421,In_289,In_869);
nand U1422 (N_1422,In_81,In_741);
or U1423 (N_1423,In_65,In_718);
nand U1424 (N_1424,In_305,In_57);
xnor U1425 (N_1425,In_414,In_539);
and U1426 (N_1426,In_308,In_750);
or U1427 (N_1427,In_549,In_159);
or U1428 (N_1428,In_80,In_405);
or U1429 (N_1429,In_290,In_708);
or U1430 (N_1430,In_293,In_546);
xor U1431 (N_1431,In_253,In_457);
and U1432 (N_1432,In_599,In_204);
and U1433 (N_1433,In_266,In_230);
and U1434 (N_1434,In_41,In_165);
and U1435 (N_1435,In_334,In_684);
or U1436 (N_1436,In_355,In_445);
nor U1437 (N_1437,In_321,In_598);
or U1438 (N_1438,In_535,In_107);
and U1439 (N_1439,In_686,In_706);
and U1440 (N_1440,In_698,In_204);
or U1441 (N_1441,In_789,In_287);
and U1442 (N_1442,In_434,In_832);
or U1443 (N_1443,In_700,In_196);
or U1444 (N_1444,In_182,In_526);
or U1445 (N_1445,In_778,In_180);
or U1446 (N_1446,In_86,In_115);
nor U1447 (N_1447,In_486,In_431);
or U1448 (N_1448,In_941,In_49);
nand U1449 (N_1449,In_479,In_528);
or U1450 (N_1450,In_983,In_484);
nand U1451 (N_1451,In_90,In_200);
or U1452 (N_1452,In_532,In_309);
or U1453 (N_1453,In_846,In_906);
or U1454 (N_1454,In_139,In_128);
and U1455 (N_1455,In_195,In_936);
and U1456 (N_1456,In_894,In_989);
or U1457 (N_1457,In_67,In_334);
nand U1458 (N_1458,In_56,In_585);
or U1459 (N_1459,In_241,In_332);
nor U1460 (N_1460,In_656,In_60);
or U1461 (N_1461,In_275,In_398);
and U1462 (N_1462,In_32,In_288);
nor U1463 (N_1463,In_847,In_713);
and U1464 (N_1464,In_63,In_718);
nand U1465 (N_1465,In_477,In_568);
or U1466 (N_1466,In_443,In_21);
nor U1467 (N_1467,In_59,In_841);
nand U1468 (N_1468,In_831,In_340);
nand U1469 (N_1469,In_525,In_997);
nor U1470 (N_1470,In_494,In_460);
or U1471 (N_1471,In_756,In_340);
nor U1472 (N_1472,In_6,In_12);
nand U1473 (N_1473,In_937,In_685);
and U1474 (N_1474,In_734,In_898);
nor U1475 (N_1475,In_32,In_157);
or U1476 (N_1476,In_177,In_781);
and U1477 (N_1477,In_668,In_637);
nor U1478 (N_1478,In_288,In_667);
or U1479 (N_1479,In_609,In_963);
nor U1480 (N_1480,In_864,In_248);
or U1481 (N_1481,In_193,In_716);
nor U1482 (N_1482,In_580,In_875);
nor U1483 (N_1483,In_605,In_425);
and U1484 (N_1484,In_557,In_337);
nand U1485 (N_1485,In_282,In_584);
nor U1486 (N_1486,In_715,In_467);
and U1487 (N_1487,In_632,In_771);
nor U1488 (N_1488,In_48,In_683);
or U1489 (N_1489,In_898,In_766);
and U1490 (N_1490,In_453,In_172);
or U1491 (N_1491,In_514,In_432);
nor U1492 (N_1492,In_996,In_976);
xor U1493 (N_1493,In_846,In_429);
or U1494 (N_1494,In_367,In_309);
and U1495 (N_1495,In_459,In_660);
nand U1496 (N_1496,In_813,In_767);
or U1497 (N_1497,In_118,In_440);
and U1498 (N_1498,In_166,In_463);
nand U1499 (N_1499,In_721,In_260);
and U1500 (N_1500,In_704,In_255);
and U1501 (N_1501,In_210,In_944);
and U1502 (N_1502,In_796,In_769);
or U1503 (N_1503,In_406,In_782);
nand U1504 (N_1504,In_934,In_195);
nand U1505 (N_1505,In_150,In_506);
and U1506 (N_1506,In_922,In_591);
xor U1507 (N_1507,In_145,In_442);
nand U1508 (N_1508,In_727,In_463);
nand U1509 (N_1509,In_379,In_128);
nand U1510 (N_1510,In_916,In_113);
nor U1511 (N_1511,In_431,In_91);
nand U1512 (N_1512,In_290,In_312);
or U1513 (N_1513,In_836,In_396);
nand U1514 (N_1514,In_674,In_476);
and U1515 (N_1515,In_354,In_909);
nor U1516 (N_1516,In_373,In_65);
nor U1517 (N_1517,In_937,In_117);
nor U1518 (N_1518,In_870,In_957);
and U1519 (N_1519,In_787,In_427);
nand U1520 (N_1520,In_731,In_375);
and U1521 (N_1521,In_831,In_295);
or U1522 (N_1522,In_721,In_235);
nand U1523 (N_1523,In_890,In_751);
or U1524 (N_1524,In_443,In_253);
nand U1525 (N_1525,In_928,In_260);
nor U1526 (N_1526,In_45,In_541);
or U1527 (N_1527,In_870,In_997);
nand U1528 (N_1528,In_982,In_667);
nor U1529 (N_1529,In_775,In_319);
nor U1530 (N_1530,In_140,In_376);
and U1531 (N_1531,In_302,In_259);
nor U1532 (N_1532,In_495,In_318);
and U1533 (N_1533,In_179,In_944);
nand U1534 (N_1534,In_771,In_997);
nand U1535 (N_1535,In_637,In_455);
xnor U1536 (N_1536,In_81,In_727);
nor U1537 (N_1537,In_417,In_634);
nor U1538 (N_1538,In_870,In_263);
nand U1539 (N_1539,In_629,In_964);
xnor U1540 (N_1540,In_239,In_806);
nor U1541 (N_1541,In_748,In_767);
nor U1542 (N_1542,In_296,In_717);
or U1543 (N_1543,In_878,In_610);
and U1544 (N_1544,In_831,In_742);
nand U1545 (N_1545,In_358,In_53);
and U1546 (N_1546,In_152,In_562);
nor U1547 (N_1547,In_34,In_902);
nor U1548 (N_1548,In_875,In_125);
or U1549 (N_1549,In_859,In_197);
or U1550 (N_1550,In_68,In_324);
nand U1551 (N_1551,In_267,In_823);
nand U1552 (N_1552,In_111,In_787);
nor U1553 (N_1553,In_775,In_23);
nor U1554 (N_1554,In_815,In_859);
nand U1555 (N_1555,In_565,In_56);
nand U1556 (N_1556,In_128,In_27);
nand U1557 (N_1557,In_487,In_247);
nand U1558 (N_1558,In_364,In_535);
nor U1559 (N_1559,In_656,In_716);
nor U1560 (N_1560,In_205,In_660);
or U1561 (N_1561,In_952,In_895);
and U1562 (N_1562,In_594,In_31);
nor U1563 (N_1563,In_474,In_459);
nand U1564 (N_1564,In_272,In_826);
nor U1565 (N_1565,In_501,In_411);
nor U1566 (N_1566,In_301,In_104);
or U1567 (N_1567,In_11,In_618);
nor U1568 (N_1568,In_199,In_611);
or U1569 (N_1569,In_116,In_315);
nor U1570 (N_1570,In_295,In_810);
and U1571 (N_1571,In_611,In_105);
and U1572 (N_1572,In_377,In_888);
nand U1573 (N_1573,In_401,In_830);
nand U1574 (N_1574,In_803,In_702);
and U1575 (N_1575,In_314,In_523);
and U1576 (N_1576,In_65,In_521);
nor U1577 (N_1577,In_185,In_607);
or U1578 (N_1578,In_642,In_817);
or U1579 (N_1579,In_549,In_65);
or U1580 (N_1580,In_505,In_24);
and U1581 (N_1581,In_605,In_574);
nor U1582 (N_1582,In_656,In_268);
nand U1583 (N_1583,In_338,In_414);
nor U1584 (N_1584,In_791,In_437);
and U1585 (N_1585,In_805,In_184);
nand U1586 (N_1586,In_890,In_605);
nand U1587 (N_1587,In_476,In_689);
nor U1588 (N_1588,In_6,In_722);
or U1589 (N_1589,In_830,In_856);
nand U1590 (N_1590,In_355,In_955);
and U1591 (N_1591,In_447,In_634);
or U1592 (N_1592,In_493,In_5);
nor U1593 (N_1593,In_744,In_360);
nor U1594 (N_1594,In_748,In_544);
nand U1595 (N_1595,In_517,In_722);
and U1596 (N_1596,In_884,In_812);
or U1597 (N_1597,In_549,In_66);
or U1598 (N_1598,In_985,In_55);
or U1599 (N_1599,In_738,In_176);
or U1600 (N_1600,In_899,In_715);
nor U1601 (N_1601,In_695,In_572);
or U1602 (N_1602,In_616,In_938);
and U1603 (N_1603,In_423,In_427);
nor U1604 (N_1604,In_383,In_769);
and U1605 (N_1605,In_279,In_597);
xor U1606 (N_1606,In_281,In_214);
and U1607 (N_1607,In_323,In_104);
xnor U1608 (N_1608,In_594,In_386);
or U1609 (N_1609,In_421,In_814);
nor U1610 (N_1610,In_624,In_73);
nand U1611 (N_1611,In_316,In_639);
and U1612 (N_1612,In_914,In_817);
nand U1613 (N_1613,In_537,In_264);
nor U1614 (N_1614,In_166,In_257);
xor U1615 (N_1615,In_326,In_237);
nand U1616 (N_1616,In_699,In_998);
nand U1617 (N_1617,In_490,In_961);
and U1618 (N_1618,In_922,In_704);
nand U1619 (N_1619,In_33,In_86);
or U1620 (N_1620,In_951,In_202);
nand U1621 (N_1621,In_137,In_201);
and U1622 (N_1622,In_796,In_738);
or U1623 (N_1623,In_379,In_989);
and U1624 (N_1624,In_798,In_985);
and U1625 (N_1625,In_66,In_101);
nand U1626 (N_1626,In_743,In_224);
xnor U1627 (N_1627,In_455,In_591);
and U1628 (N_1628,In_289,In_848);
nand U1629 (N_1629,In_916,In_73);
and U1630 (N_1630,In_861,In_19);
or U1631 (N_1631,In_496,In_29);
and U1632 (N_1632,In_428,In_617);
xor U1633 (N_1633,In_410,In_214);
nor U1634 (N_1634,In_415,In_531);
and U1635 (N_1635,In_659,In_562);
xor U1636 (N_1636,In_621,In_255);
or U1637 (N_1637,In_763,In_326);
or U1638 (N_1638,In_164,In_42);
and U1639 (N_1639,In_671,In_109);
nor U1640 (N_1640,In_535,In_640);
and U1641 (N_1641,In_594,In_856);
and U1642 (N_1642,In_410,In_649);
or U1643 (N_1643,In_580,In_138);
or U1644 (N_1644,In_884,In_644);
and U1645 (N_1645,In_936,In_11);
nor U1646 (N_1646,In_380,In_553);
nand U1647 (N_1647,In_483,In_150);
nor U1648 (N_1648,In_363,In_88);
and U1649 (N_1649,In_202,In_838);
nor U1650 (N_1650,In_244,In_895);
or U1651 (N_1651,In_799,In_307);
xor U1652 (N_1652,In_267,In_525);
and U1653 (N_1653,In_185,In_17);
and U1654 (N_1654,In_740,In_689);
nor U1655 (N_1655,In_341,In_901);
nor U1656 (N_1656,In_574,In_382);
nand U1657 (N_1657,In_881,In_992);
and U1658 (N_1658,In_155,In_523);
nand U1659 (N_1659,In_77,In_217);
nor U1660 (N_1660,In_822,In_418);
and U1661 (N_1661,In_442,In_341);
nand U1662 (N_1662,In_285,In_957);
or U1663 (N_1663,In_883,In_511);
nand U1664 (N_1664,In_702,In_131);
or U1665 (N_1665,In_406,In_553);
and U1666 (N_1666,In_87,In_597);
and U1667 (N_1667,In_778,In_283);
or U1668 (N_1668,In_912,In_423);
nor U1669 (N_1669,In_127,In_738);
xor U1670 (N_1670,In_502,In_160);
or U1671 (N_1671,In_318,In_189);
nor U1672 (N_1672,In_545,In_42);
nor U1673 (N_1673,In_285,In_689);
or U1674 (N_1674,In_854,In_547);
or U1675 (N_1675,In_21,In_101);
nor U1676 (N_1676,In_117,In_136);
xnor U1677 (N_1677,In_284,In_897);
nor U1678 (N_1678,In_680,In_76);
nand U1679 (N_1679,In_934,In_383);
or U1680 (N_1680,In_54,In_295);
and U1681 (N_1681,In_547,In_732);
and U1682 (N_1682,In_491,In_731);
nand U1683 (N_1683,In_472,In_958);
nor U1684 (N_1684,In_865,In_588);
nor U1685 (N_1685,In_113,In_735);
or U1686 (N_1686,In_870,In_516);
nand U1687 (N_1687,In_630,In_603);
or U1688 (N_1688,In_828,In_591);
or U1689 (N_1689,In_25,In_713);
or U1690 (N_1690,In_920,In_432);
or U1691 (N_1691,In_898,In_269);
nand U1692 (N_1692,In_629,In_844);
or U1693 (N_1693,In_566,In_14);
and U1694 (N_1694,In_434,In_35);
or U1695 (N_1695,In_111,In_55);
nor U1696 (N_1696,In_536,In_820);
and U1697 (N_1697,In_311,In_812);
nor U1698 (N_1698,In_127,In_673);
xnor U1699 (N_1699,In_647,In_679);
or U1700 (N_1700,In_982,In_651);
nor U1701 (N_1701,In_634,In_134);
or U1702 (N_1702,In_979,In_331);
nand U1703 (N_1703,In_548,In_621);
nor U1704 (N_1704,In_346,In_543);
or U1705 (N_1705,In_614,In_816);
nor U1706 (N_1706,In_593,In_663);
and U1707 (N_1707,In_822,In_61);
or U1708 (N_1708,In_330,In_54);
and U1709 (N_1709,In_494,In_777);
and U1710 (N_1710,In_406,In_349);
or U1711 (N_1711,In_307,In_649);
or U1712 (N_1712,In_806,In_837);
and U1713 (N_1713,In_595,In_389);
or U1714 (N_1714,In_123,In_404);
or U1715 (N_1715,In_691,In_612);
or U1716 (N_1716,In_118,In_551);
nor U1717 (N_1717,In_75,In_332);
or U1718 (N_1718,In_238,In_61);
and U1719 (N_1719,In_792,In_595);
or U1720 (N_1720,In_155,In_338);
and U1721 (N_1721,In_675,In_315);
and U1722 (N_1722,In_861,In_75);
or U1723 (N_1723,In_139,In_425);
or U1724 (N_1724,In_283,In_402);
or U1725 (N_1725,In_109,In_594);
nor U1726 (N_1726,In_664,In_485);
nor U1727 (N_1727,In_667,In_664);
nand U1728 (N_1728,In_616,In_901);
and U1729 (N_1729,In_477,In_744);
nor U1730 (N_1730,In_752,In_674);
or U1731 (N_1731,In_502,In_607);
nor U1732 (N_1732,In_949,In_457);
or U1733 (N_1733,In_716,In_514);
and U1734 (N_1734,In_177,In_883);
or U1735 (N_1735,In_989,In_67);
nand U1736 (N_1736,In_473,In_428);
and U1737 (N_1737,In_4,In_955);
nor U1738 (N_1738,In_810,In_221);
or U1739 (N_1739,In_747,In_58);
or U1740 (N_1740,In_842,In_259);
nand U1741 (N_1741,In_188,In_799);
and U1742 (N_1742,In_804,In_682);
and U1743 (N_1743,In_358,In_442);
or U1744 (N_1744,In_238,In_695);
nor U1745 (N_1745,In_960,In_301);
and U1746 (N_1746,In_382,In_134);
nand U1747 (N_1747,In_725,In_195);
xnor U1748 (N_1748,In_886,In_809);
nand U1749 (N_1749,In_679,In_127);
or U1750 (N_1750,In_696,In_136);
nor U1751 (N_1751,In_998,In_394);
nor U1752 (N_1752,In_861,In_914);
nand U1753 (N_1753,In_326,In_824);
or U1754 (N_1754,In_418,In_947);
and U1755 (N_1755,In_275,In_690);
nor U1756 (N_1756,In_984,In_291);
or U1757 (N_1757,In_266,In_646);
xor U1758 (N_1758,In_949,In_116);
and U1759 (N_1759,In_418,In_45);
and U1760 (N_1760,In_509,In_216);
and U1761 (N_1761,In_433,In_284);
nand U1762 (N_1762,In_920,In_606);
nand U1763 (N_1763,In_630,In_371);
or U1764 (N_1764,In_897,In_115);
or U1765 (N_1765,In_459,In_297);
nor U1766 (N_1766,In_540,In_783);
nand U1767 (N_1767,In_756,In_513);
nand U1768 (N_1768,In_640,In_224);
nand U1769 (N_1769,In_854,In_113);
or U1770 (N_1770,In_899,In_195);
nor U1771 (N_1771,In_446,In_516);
nand U1772 (N_1772,In_75,In_448);
and U1773 (N_1773,In_910,In_834);
nor U1774 (N_1774,In_623,In_104);
nor U1775 (N_1775,In_898,In_714);
nor U1776 (N_1776,In_327,In_868);
nand U1777 (N_1777,In_502,In_846);
and U1778 (N_1778,In_476,In_681);
nand U1779 (N_1779,In_68,In_125);
and U1780 (N_1780,In_849,In_783);
xnor U1781 (N_1781,In_819,In_96);
or U1782 (N_1782,In_103,In_40);
and U1783 (N_1783,In_292,In_510);
xnor U1784 (N_1784,In_869,In_653);
or U1785 (N_1785,In_484,In_369);
and U1786 (N_1786,In_853,In_176);
or U1787 (N_1787,In_571,In_92);
or U1788 (N_1788,In_663,In_860);
and U1789 (N_1789,In_850,In_597);
and U1790 (N_1790,In_792,In_146);
nor U1791 (N_1791,In_902,In_405);
or U1792 (N_1792,In_919,In_268);
and U1793 (N_1793,In_348,In_165);
or U1794 (N_1794,In_90,In_40);
or U1795 (N_1795,In_643,In_80);
nor U1796 (N_1796,In_561,In_428);
or U1797 (N_1797,In_746,In_64);
or U1798 (N_1798,In_782,In_199);
xnor U1799 (N_1799,In_743,In_415);
or U1800 (N_1800,In_697,In_359);
or U1801 (N_1801,In_234,In_264);
or U1802 (N_1802,In_878,In_832);
nand U1803 (N_1803,In_228,In_872);
nor U1804 (N_1804,In_97,In_139);
and U1805 (N_1805,In_510,In_303);
nand U1806 (N_1806,In_697,In_583);
or U1807 (N_1807,In_807,In_911);
nor U1808 (N_1808,In_86,In_522);
nor U1809 (N_1809,In_354,In_151);
nor U1810 (N_1810,In_859,In_377);
xnor U1811 (N_1811,In_870,In_602);
or U1812 (N_1812,In_840,In_941);
nand U1813 (N_1813,In_754,In_100);
or U1814 (N_1814,In_602,In_230);
nor U1815 (N_1815,In_229,In_419);
nor U1816 (N_1816,In_604,In_528);
xor U1817 (N_1817,In_666,In_132);
nor U1818 (N_1818,In_39,In_80);
nor U1819 (N_1819,In_839,In_43);
nand U1820 (N_1820,In_10,In_883);
nand U1821 (N_1821,In_917,In_712);
and U1822 (N_1822,In_926,In_573);
or U1823 (N_1823,In_381,In_223);
and U1824 (N_1824,In_319,In_658);
and U1825 (N_1825,In_436,In_248);
and U1826 (N_1826,In_130,In_764);
nor U1827 (N_1827,In_769,In_247);
nor U1828 (N_1828,In_469,In_109);
or U1829 (N_1829,In_356,In_498);
or U1830 (N_1830,In_25,In_257);
or U1831 (N_1831,In_848,In_177);
or U1832 (N_1832,In_654,In_635);
nand U1833 (N_1833,In_325,In_246);
and U1834 (N_1834,In_483,In_193);
nor U1835 (N_1835,In_217,In_507);
nand U1836 (N_1836,In_468,In_265);
nor U1837 (N_1837,In_785,In_587);
and U1838 (N_1838,In_747,In_69);
and U1839 (N_1839,In_341,In_960);
and U1840 (N_1840,In_394,In_54);
nand U1841 (N_1841,In_682,In_352);
or U1842 (N_1842,In_271,In_401);
nand U1843 (N_1843,In_224,In_444);
or U1844 (N_1844,In_85,In_112);
or U1845 (N_1845,In_141,In_299);
or U1846 (N_1846,In_131,In_613);
nand U1847 (N_1847,In_399,In_250);
nand U1848 (N_1848,In_170,In_249);
nor U1849 (N_1849,In_795,In_115);
nor U1850 (N_1850,In_518,In_293);
or U1851 (N_1851,In_507,In_420);
nor U1852 (N_1852,In_227,In_364);
nand U1853 (N_1853,In_349,In_691);
nand U1854 (N_1854,In_804,In_211);
or U1855 (N_1855,In_722,In_602);
nand U1856 (N_1856,In_835,In_933);
nand U1857 (N_1857,In_222,In_931);
nand U1858 (N_1858,In_376,In_280);
or U1859 (N_1859,In_679,In_540);
nor U1860 (N_1860,In_213,In_457);
and U1861 (N_1861,In_306,In_942);
or U1862 (N_1862,In_152,In_224);
xnor U1863 (N_1863,In_652,In_239);
nor U1864 (N_1864,In_2,In_180);
and U1865 (N_1865,In_910,In_687);
nor U1866 (N_1866,In_411,In_300);
or U1867 (N_1867,In_177,In_460);
or U1868 (N_1868,In_518,In_152);
xnor U1869 (N_1869,In_886,In_837);
and U1870 (N_1870,In_568,In_5);
nor U1871 (N_1871,In_218,In_988);
nand U1872 (N_1872,In_336,In_783);
nand U1873 (N_1873,In_740,In_871);
nand U1874 (N_1874,In_706,In_268);
nor U1875 (N_1875,In_630,In_777);
nor U1876 (N_1876,In_599,In_125);
or U1877 (N_1877,In_34,In_912);
and U1878 (N_1878,In_996,In_61);
and U1879 (N_1879,In_445,In_760);
or U1880 (N_1880,In_886,In_844);
nor U1881 (N_1881,In_791,In_540);
nor U1882 (N_1882,In_26,In_474);
and U1883 (N_1883,In_453,In_305);
nor U1884 (N_1884,In_894,In_978);
nor U1885 (N_1885,In_246,In_94);
and U1886 (N_1886,In_229,In_753);
xor U1887 (N_1887,In_262,In_951);
and U1888 (N_1888,In_189,In_737);
and U1889 (N_1889,In_385,In_162);
nand U1890 (N_1890,In_488,In_604);
nand U1891 (N_1891,In_551,In_11);
nor U1892 (N_1892,In_862,In_843);
xnor U1893 (N_1893,In_656,In_606);
xor U1894 (N_1894,In_620,In_594);
or U1895 (N_1895,In_50,In_310);
or U1896 (N_1896,In_942,In_673);
and U1897 (N_1897,In_750,In_898);
or U1898 (N_1898,In_127,In_488);
or U1899 (N_1899,In_370,In_366);
nor U1900 (N_1900,In_805,In_881);
nand U1901 (N_1901,In_703,In_138);
nand U1902 (N_1902,In_572,In_793);
and U1903 (N_1903,In_239,In_152);
or U1904 (N_1904,In_306,In_701);
and U1905 (N_1905,In_28,In_289);
xnor U1906 (N_1906,In_271,In_201);
and U1907 (N_1907,In_573,In_586);
or U1908 (N_1908,In_157,In_343);
and U1909 (N_1909,In_10,In_546);
nand U1910 (N_1910,In_153,In_827);
xor U1911 (N_1911,In_888,In_625);
xnor U1912 (N_1912,In_676,In_349);
nand U1913 (N_1913,In_760,In_948);
nor U1914 (N_1914,In_586,In_747);
nor U1915 (N_1915,In_638,In_432);
or U1916 (N_1916,In_797,In_751);
nand U1917 (N_1917,In_302,In_623);
and U1918 (N_1918,In_428,In_235);
and U1919 (N_1919,In_917,In_963);
nand U1920 (N_1920,In_137,In_71);
and U1921 (N_1921,In_570,In_353);
nand U1922 (N_1922,In_217,In_461);
nor U1923 (N_1923,In_894,In_903);
or U1924 (N_1924,In_661,In_466);
nor U1925 (N_1925,In_999,In_151);
and U1926 (N_1926,In_858,In_153);
or U1927 (N_1927,In_693,In_92);
and U1928 (N_1928,In_554,In_7);
nand U1929 (N_1929,In_267,In_899);
and U1930 (N_1930,In_631,In_113);
nor U1931 (N_1931,In_518,In_95);
nand U1932 (N_1932,In_328,In_795);
nor U1933 (N_1933,In_269,In_119);
and U1934 (N_1934,In_82,In_968);
nand U1935 (N_1935,In_503,In_977);
or U1936 (N_1936,In_333,In_645);
nor U1937 (N_1937,In_195,In_895);
nor U1938 (N_1938,In_987,In_259);
or U1939 (N_1939,In_123,In_361);
nand U1940 (N_1940,In_883,In_427);
or U1941 (N_1941,In_679,In_363);
and U1942 (N_1942,In_789,In_556);
and U1943 (N_1943,In_779,In_5);
nor U1944 (N_1944,In_89,In_854);
nand U1945 (N_1945,In_956,In_437);
nor U1946 (N_1946,In_893,In_53);
and U1947 (N_1947,In_95,In_93);
and U1948 (N_1948,In_343,In_841);
and U1949 (N_1949,In_278,In_72);
or U1950 (N_1950,In_917,In_101);
and U1951 (N_1951,In_804,In_731);
nor U1952 (N_1952,In_657,In_18);
and U1953 (N_1953,In_605,In_140);
and U1954 (N_1954,In_174,In_776);
nand U1955 (N_1955,In_655,In_133);
and U1956 (N_1956,In_873,In_772);
or U1957 (N_1957,In_577,In_101);
and U1958 (N_1958,In_214,In_886);
nor U1959 (N_1959,In_398,In_515);
and U1960 (N_1960,In_111,In_650);
nor U1961 (N_1961,In_570,In_748);
nor U1962 (N_1962,In_240,In_861);
nor U1963 (N_1963,In_651,In_272);
nand U1964 (N_1964,In_297,In_707);
and U1965 (N_1965,In_470,In_651);
and U1966 (N_1966,In_739,In_458);
nor U1967 (N_1967,In_738,In_356);
and U1968 (N_1968,In_199,In_151);
and U1969 (N_1969,In_918,In_988);
or U1970 (N_1970,In_369,In_762);
nor U1971 (N_1971,In_110,In_764);
or U1972 (N_1972,In_587,In_230);
or U1973 (N_1973,In_683,In_408);
nand U1974 (N_1974,In_415,In_246);
and U1975 (N_1975,In_110,In_178);
nand U1976 (N_1976,In_707,In_460);
nand U1977 (N_1977,In_498,In_100);
or U1978 (N_1978,In_152,In_890);
and U1979 (N_1979,In_159,In_67);
nor U1980 (N_1980,In_212,In_314);
nor U1981 (N_1981,In_777,In_905);
and U1982 (N_1982,In_96,In_380);
or U1983 (N_1983,In_395,In_99);
nor U1984 (N_1984,In_537,In_675);
and U1985 (N_1985,In_798,In_501);
and U1986 (N_1986,In_553,In_561);
and U1987 (N_1987,In_720,In_987);
nand U1988 (N_1988,In_237,In_426);
nor U1989 (N_1989,In_522,In_109);
and U1990 (N_1990,In_231,In_372);
or U1991 (N_1991,In_12,In_21);
nand U1992 (N_1992,In_807,In_436);
and U1993 (N_1993,In_552,In_927);
nand U1994 (N_1994,In_740,In_614);
or U1995 (N_1995,In_906,In_874);
or U1996 (N_1996,In_640,In_135);
or U1997 (N_1997,In_324,In_979);
nand U1998 (N_1998,In_539,In_878);
and U1999 (N_1999,In_762,In_422);
nor U2000 (N_2000,In_414,In_87);
xnor U2001 (N_2001,In_856,In_969);
or U2002 (N_2002,In_165,In_997);
nand U2003 (N_2003,In_380,In_567);
and U2004 (N_2004,In_295,In_951);
and U2005 (N_2005,In_630,In_503);
and U2006 (N_2006,In_569,In_800);
nand U2007 (N_2007,In_141,In_743);
nand U2008 (N_2008,In_334,In_635);
nor U2009 (N_2009,In_925,In_213);
and U2010 (N_2010,In_451,In_396);
or U2011 (N_2011,In_496,In_635);
or U2012 (N_2012,In_785,In_681);
nand U2013 (N_2013,In_367,In_228);
and U2014 (N_2014,In_983,In_677);
or U2015 (N_2015,In_190,In_189);
nor U2016 (N_2016,In_728,In_472);
nand U2017 (N_2017,In_194,In_206);
and U2018 (N_2018,In_209,In_888);
and U2019 (N_2019,In_747,In_504);
nand U2020 (N_2020,In_788,In_276);
or U2021 (N_2021,In_974,In_855);
nand U2022 (N_2022,In_90,In_494);
nor U2023 (N_2023,In_209,In_517);
nor U2024 (N_2024,In_606,In_235);
nand U2025 (N_2025,In_438,In_167);
nand U2026 (N_2026,In_178,In_754);
nor U2027 (N_2027,In_949,In_178);
or U2028 (N_2028,In_262,In_500);
nor U2029 (N_2029,In_215,In_506);
or U2030 (N_2030,In_174,In_302);
nor U2031 (N_2031,In_799,In_851);
and U2032 (N_2032,In_837,In_318);
nor U2033 (N_2033,In_87,In_177);
nand U2034 (N_2034,In_331,In_516);
and U2035 (N_2035,In_329,In_75);
nor U2036 (N_2036,In_999,In_655);
or U2037 (N_2037,In_305,In_130);
nor U2038 (N_2038,In_772,In_53);
or U2039 (N_2039,In_843,In_230);
or U2040 (N_2040,In_658,In_200);
and U2041 (N_2041,In_368,In_658);
nor U2042 (N_2042,In_779,In_215);
xor U2043 (N_2043,In_721,In_479);
or U2044 (N_2044,In_378,In_414);
and U2045 (N_2045,In_510,In_587);
nand U2046 (N_2046,In_676,In_273);
nand U2047 (N_2047,In_257,In_779);
nor U2048 (N_2048,In_617,In_198);
nand U2049 (N_2049,In_240,In_836);
or U2050 (N_2050,In_651,In_418);
nor U2051 (N_2051,In_407,In_402);
nor U2052 (N_2052,In_234,In_508);
nand U2053 (N_2053,In_799,In_199);
or U2054 (N_2054,In_40,In_246);
or U2055 (N_2055,In_313,In_640);
or U2056 (N_2056,In_628,In_608);
or U2057 (N_2057,In_36,In_377);
nand U2058 (N_2058,In_976,In_249);
and U2059 (N_2059,In_57,In_833);
nand U2060 (N_2060,In_882,In_17);
nand U2061 (N_2061,In_822,In_263);
nor U2062 (N_2062,In_25,In_559);
or U2063 (N_2063,In_672,In_110);
or U2064 (N_2064,In_333,In_287);
nand U2065 (N_2065,In_581,In_42);
and U2066 (N_2066,In_235,In_472);
and U2067 (N_2067,In_338,In_834);
and U2068 (N_2068,In_411,In_838);
and U2069 (N_2069,In_237,In_647);
nand U2070 (N_2070,In_591,In_304);
and U2071 (N_2071,In_49,In_166);
nor U2072 (N_2072,In_842,In_644);
xnor U2073 (N_2073,In_891,In_499);
or U2074 (N_2074,In_751,In_732);
and U2075 (N_2075,In_402,In_103);
or U2076 (N_2076,In_984,In_550);
nand U2077 (N_2077,In_229,In_890);
and U2078 (N_2078,In_679,In_488);
or U2079 (N_2079,In_697,In_133);
or U2080 (N_2080,In_818,In_896);
and U2081 (N_2081,In_433,In_788);
nand U2082 (N_2082,In_338,In_60);
and U2083 (N_2083,In_663,In_76);
nor U2084 (N_2084,In_432,In_473);
nor U2085 (N_2085,In_680,In_198);
xnor U2086 (N_2086,In_371,In_678);
and U2087 (N_2087,In_183,In_81);
nand U2088 (N_2088,In_249,In_887);
and U2089 (N_2089,In_212,In_271);
and U2090 (N_2090,In_316,In_277);
nand U2091 (N_2091,In_40,In_953);
nand U2092 (N_2092,In_434,In_538);
or U2093 (N_2093,In_171,In_933);
nand U2094 (N_2094,In_891,In_276);
or U2095 (N_2095,In_935,In_699);
and U2096 (N_2096,In_632,In_296);
and U2097 (N_2097,In_69,In_858);
or U2098 (N_2098,In_475,In_851);
nand U2099 (N_2099,In_604,In_331);
nand U2100 (N_2100,In_824,In_234);
and U2101 (N_2101,In_481,In_76);
nand U2102 (N_2102,In_539,In_151);
nand U2103 (N_2103,In_515,In_374);
or U2104 (N_2104,In_858,In_815);
or U2105 (N_2105,In_985,In_927);
or U2106 (N_2106,In_9,In_276);
or U2107 (N_2107,In_579,In_265);
nand U2108 (N_2108,In_20,In_788);
and U2109 (N_2109,In_933,In_887);
nand U2110 (N_2110,In_627,In_65);
and U2111 (N_2111,In_59,In_152);
nand U2112 (N_2112,In_124,In_132);
and U2113 (N_2113,In_118,In_317);
nand U2114 (N_2114,In_840,In_596);
or U2115 (N_2115,In_649,In_173);
nand U2116 (N_2116,In_434,In_99);
nand U2117 (N_2117,In_667,In_183);
xnor U2118 (N_2118,In_880,In_611);
and U2119 (N_2119,In_647,In_387);
nand U2120 (N_2120,In_100,In_4);
nor U2121 (N_2121,In_148,In_441);
nor U2122 (N_2122,In_372,In_929);
and U2123 (N_2123,In_15,In_51);
and U2124 (N_2124,In_554,In_949);
and U2125 (N_2125,In_658,In_988);
nor U2126 (N_2126,In_370,In_70);
nor U2127 (N_2127,In_783,In_743);
nor U2128 (N_2128,In_915,In_703);
and U2129 (N_2129,In_217,In_924);
nor U2130 (N_2130,In_596,In_875);
or U2131 (N_2131,In_382,In_190);
nand U2132 (N_2132,In_396,In_780);
nor U2133 (N_2133,In_623,In_826);
nand U2134 (N_2134,In_565,In_540);
nor U2135 (N_2135,In_626,In_623);
and U2136 (N_2136,In_282,In_88);
nand U2137 (N_2137,In_478,In_365);
and U2138 (N_2138,In_277,In_752);
xnor U2139 (N_2139,In_53,In_17);
nor U2140 (N_2140,In_671,In_765);
nor U2141 (N_2141,In_820,In_694);
nor U2142 (N_2142,In_85,In_555);
or U2143 (N_2143,In_481,In_661);
and U2144 (N_2144,In_629,In_59);
nor U2145 (N_2145,In_843,In_783);
nand U2146 (N_2146,In_551,In_485);
nand U2147 (N_2147,In_293,In_332);
nand U2148 (N_2148,In_762,In_586);
nor U2149 (N_2149,In_296,In_4);
and U2150 (N_2150,In_79,In_118);
nor U2151 (N_2151,In_984,In_935);
or U2152 (N_2152,In_651,In_404);
or U2153 (N_2153,In_828,In_712);
nand U2154 (N_2154,In_779,In_929);
and U2155 (N_2155,In_838,In_465);
nor U2156 (N_2156,In_548,In_566);
nor U2157 (N_2157,In_993,In_784);
nand U2158 (N_2158,In_782,In_498);
or U2159 (N_2159,In_443,In_786);
and U2160 (N_2160,In_716,In_337);
or U2161 (N_2161,In_167,In_266);
and U2162 (N_2162,In_196,In_946);
or U2163 (N_2163,In_864,In_585);
nor U2164 (N_2164,In_432,In_242);
nand U2165 (N_2165,In_199,In_881);
nand U2166 (N_2166,In_296,In_836);
and U2167 (N_2167,In_61,In_293);
or U2168 (N_2168,In_745,In_94);
and U2169 (N_2169,In_104,In_766);
xor U2170 (N_2170,In_120,In_666);
nand U2171 (N_2171,In_237,In_383);
nand U2172 (N_2172,In_771,In_232);
nand U2173 (N_2173,In_123,In_952);
nor U2174 (N_2174,In_339,In_186);
nand U2175 (N_2175,In_829,In_451);
or U2176 (N_2176,In_45,In_10);
nor U2177 (N_2177,In_4,In_722);
nor U2178 (N_2178,In_796,In_403);
or U2179 (N_2179,In_947,In_984);
or U2180 (N_2180,In_664,In_986);
and U2181 (N_2181,In_182,In_44);
or U2182 (N_2182,In_755,In_255);
or U2183 (N_2183,In_417,In_149);
or U2184 (N_2184,In_260,In_40);
and U2185 (N_2185,In_404,In_197);
or U2186 (N_2186,In_830,In_525);
or U2187 (N_2187,In_690,In_542);
and U2188 (N_2188,In_717,In_382);
nor U2189 (N_2189,In_770,In_198);
nor U2190 (N_2190,In_757,In_868);
nor U2191 (N_2191,In_579,In_497);
or U2192 (N_2192,In_82,In_172);
nand U2193 (N_2193,In_837,In_846);
nor U2194 (N_2194,In_420,In_681);
or U2195 (N_2195,In_97,In_119);
nand U2196 (N_2196,In_472,In_685);
and U2197 (N_2197,In_954,In_809);
xnor U2198 (N_2198,In_720,In_457);
and U2199 (N_2199,In_44,In_250);
nor U2200 (N_2200,In_459,In_217);
nand U2201 (N_2201,In_142,In_484);
nand U2202 (N_2202,In_955,In_952);
or U2203 (N_2203,In_550,In_989);
and U2204 (N_2204,In_407,In_698);
or U2205 (N_2205,In_998,In_182);
or U2206 (N_2206,In_136,In_204);
nand U2207 (N_2207,In_27,In_269);
nand U2208 (N_2208,In_873,In_922);
nand U2209 (N_2209,In_829,In_713);
nand U2210 (N_2210,In_812,In_96);
or U2211 (N_2211,In_272,In_188);
nor U2212 (N_2212,In_57,In_377);
or U2213 (N_2213,In_117,In_602);
and U2214 (N_2214,In_117,In_206);
nor U2215 (N_2215,In_671,In_758);
and U2216 (N_2216,In_736,In_500);
nand U2217 (N_2217,In_963,In_517);
or U2218 (N_2218,In_664,In_529);
nor U2219 (N_2219,In_502,In_114);
and U2220 (N_2220,In_658,In_925);
or U2221 (N_2221,In_255,In_426);
nand U2222 (N_2222,In_947,In_329);
and U2223 (N_2223,In_269,In_147);
or U2224 (N_2224,In_502,In_460);
or U2225 (N_2225,In_444,In_834);
nor U2226 (N_2226,In_894,In_615);
and U2227 (N_2227,In_71,In_518);
or U2228 (N_2228,In_206,In_815);
or U2229 (N_2229,In_219,In_348);
and U2230 (N_2230,In_972,In_658);
nand U2231 (N_2231,In_3,In_4);
and U2232 (N_2232,In_851,In_987);
nor U2233 (N_2233,In_890,In_121);
and U2234 (N_2234,In_55,In_757);
or U2235 (N_2235,In_225,In_338);
and U2236 (N_2236,In_789,In_62);
and U2237 (N_2237,In_701,In_345);
or U2238 (N_2238,In_303,In_590);
and U2239 (N_2239,In_123,In_154);
nand U2240 (N_2240,In_638,In_333);
or U2241 (N_2241,In_273,In_18);
and U2242 (N_2242,In_124,In_224);
nor U2243 (N_2243,In_156,In_436);
or U2244 (N_2244,In_742,In_629);
xnor U2245 (N_2245,In_157,In_10);
nor U2246 (N_2246,In_102,In_366);
or U2247 (N_2247,In_384,In_316);
nor U2248 (N_2248,In_972,In_374);
nand U2249 (N_2249,In_693,In_256);
or U2250 (N_2250,In_999,In_666);
nand U2251 (N_2251,In_96,In_160);
or U2252 (N_2252,In_190,In_514);
xnor U2253 (N_2253,In_969,In_15);
and U2254 (N_2254,In_118,In_660);
or U2255 (N_2255,In_206,In_798);
nor U2256 (N_2256,In_411,In_709);
or U2257 (N_2257,In_343,In_740);
nor U2258 (N_2258,In_162,In_520);
or U2259 (N_2259,In_690,In_964);
and U2260 (N_2260,In_390,In_940);
and U2261 (N_2261,In_23,In_179);
nand U2262 (N_2262,In_939,In_518);
nand U2263 (N_2263,In_839,In_392);
nand U2264 (N_2264,In_47,In_529);
xor U2265 (N_2265,In_242,In_256);
and U2266 (N_2266,In_885,In_600);
or U2267 (N_2267,In_816,In_46);
nor U2268 (N_2268,In_228,In_82);
and U2269 (N_2269,In_19,In_701);
nor U2270 (N_2270,In_610,In_929);
nand U2271 (N_2271,In_615,In_528);
or U2272 (N_2272,In_883,In_363);
and U2273 (N_2273,In_359,In_117);
nor U2274 (N_2274,In_281,In_775);
and U2275 (N_2275,In_602,In_838);
and U2276 (N_2276,In_3,In_723);
nand U2277 (N_2277,In_349,In_272);
or U2278 (N_2278,In_831,In_323);
nor U2279 (N_2279,In_11,In_835);
nor U2280 (N_2280,In_824,In_883);
and U2281 (N_2281,In_548,In_688);
and U2282 (N_2282,In_24,In_264);
or U2283 (N_2283,In_135,In_453);
or U2284 (N_2284,In_760,In_471);
and U2285 (N_2285,In_219,In_387);
nand U2286 (N_2286,In_120,In_545);
and U2287 (N_2287,In_12,In_527);
and U2288 (N_2288,In_15,In_109);
nand U2289 (N_2289,In_813,In_612);
and U2290 (N_2290,In_269,In_637);
nor U2291 (N_2291,In_761,In_63);
and U2292 (N_2292,In_562,In_838);
or U2293 (N_2293,In_681,In_491);
nand U2294 (N_2294,In_261,In_714);
or U2295 (N_2295,In_850,In_13);
nor U2296 (N_2296,In_837,In_831);
or U2297 (N_2297,In_346,In_231);
and U2298 (N_2298,In_933,In_814);
nor U2299 (N_2299,In_647,In_193);
and U2300 (N_2300,In_370,In_535);
nor U2301 (N_2301,In_318,In_659);
nand U2302 (N_2302,In_973,In_244);
nand U2303 (N_2303,In_950,In_557);
nor U2304 (N_2304,In_450,In_180);
xor U2305 (N_2305,In_56,In_686);
nor U2306 (N_2306,In_435,In_606);
nand U2307 (N_2307,In_450,In_440);
or U2308 (N_2308,In_753,In_52);
nand U2309 (N_2309,In_172,In_850);
xor U2310 (N_2310,In_567,In_917);
nor U2311 (N_2311,In_774,In_188);
nor U2312 (N_2312,In_904,In_330);
and U2313 (N_2313,In_141,In_410);
nand U2314 (N_2314,In_437,In_335);
or U2315 (N_2315,In_47,In_998);
and U2316 (N_2316,In_622,In_243);
nor U2317 (N_2317,In_502,In_43);
nor U2318 (N_2318,In_316,In_938);
or U2319 (N_2319,In_566,In_561);
or U2320 (N_2320,In_576,In_570);
nor U2321 (N_2321,In_240,In_234);
or U2322 (N_2322,In_28,In_851);
and U2323 (N_2323,In_393,In_516);
and U2324 (N_2324,In_424,In_323);
or U2325 (N_2325,In_859,In_608);
nand U2326 (N_2326,In_97,In_472);
nor U2327 (N_2327,In_902,In_604);
or U2328 (N_2328,In_883,In_658);
nor U2329 (N_2329,In_17,In_623);
and U2330 (N_2330,In_823,In_674);
xnor U2331 (N_2331,In_897,In_645);
or U2332 (N_2332,In_127,In_725);
nor U2333 (N_2333,In_289,In_198);
nor U2334 (N_2334,In_742,In_530);
nor U2335 (N_2335,In_505,In_460);
nand U2336 (N_2336,In_370,In_271);
nand U2337 (N_2337,In_538,In_803);
or U2338 (N_2338,In_327,In_325);
nand U2339 (N_2339,In_554,In_826);
and U2340 (N_2340,In_83,In_986);
nand U2341 (N_2341,In_392,In_568);
nand U2342 (N_2342,In_466,In_668);
and U2343 (N_2343,In_489,In_561);
and U2344 (N_2344,In_512,In_287);
xor U2345 (N_2345,In_843,In_188);
nand U2346 (N_2346,In_821,In_521);
nand U2347 (N_2347,In_87,In_741);
or U2348 (N_2348,In_552,In_815);
nand U2349 (N_2349,In_659,In_580);
or U2350 (N_2350,In_568,In_169);
or U2351 (N_2351,In_377,In_817);
or U2352 (N_2352,In_870,In_537);
or U2353 (N_2353,In_762,In_710);
nand U2354 (N_2354,In_259,In_442);
nand U2355 (N_2355,In_252,In_487);
nor U2356 (N_2356,In_216,In_4);
nor U2357 (N_2357,In_238,In_984);
or U2358 (N_2358,In_755,In_699);
nand U2359 (N_2359,In_983,In_439);
nor U2360 (N_2360,In_140,In_372);
nand U2361 (N_2361,In_946,In_941);
or U2362 (N_2362,In_600,In_713);
or U2363 (N_2363,In_309,In_42);
nor U2364 (N_2364,In_741,In_898);
and U2365 (N_2365,In_8,In_620);
nand U2366 (N_2366,In_977,In_830);
and U2367 (N_2367,In_901,In_508);
nand U2368 (N_2368,In_319,In_653);
nor U2369 (N_2369,In_547,In_758);
or U2370 (N_2370,In_97,In_373);
or U2371 (N_2371,In_562,In_684);
nand U2372 (N_2372,In_443,In_804);
nor U2373 (N_2373,In_737,In_215);
nand U2374 (N_2374,In_83,In_292);
nand U2375 (N_2375,In_697,In_428);
nand U2376 (N_2376,In_577,In_98);
nand U2377 (N_2377,In_318,In_692);
and U2378 (N_2378,In_984,In_87);
nor U2379 (N_2379,In_400,In_701);
nor U2380 (N_2380,In_913,In_54);
and U2381 (N_2381,In_645,In_713);
and U2382 (N_2382,In_69,In_8);
and U2383 (N_2383,In_829,In_15);
nand U2384 (N_2384,In_521,In_979);
or U2385 (N_2385,In_874,In_111);
and U2386 (N_2386,In_797,In_561);
and U2387 (N_2387,In_478,In_111);
or U2388 (N_2388,In_66,In_968);
nand U2389 (N_2389,In_591,In_48);
nor U2390 (N_2390,In_749,In_656);
or U2391 (N_2391,In_362,In_620);
and U2392 (N_2392,In_764,In_375);
or U2393 (N_2393,In_314,In_352);
or U2394 (N_2394,In_90,In_39);
or U2395 (N_2395,In_347,In_660);
nand U2396 (N_2396,In_163,In_219);
or U2397 (N_2397,In_180,In_592);
nand U2398 (N_2398,In_807,In_482);
nor U2399 (N_2399,In_104,In_711);
or U2400 (N_2400,In_183,In_401);
nor U2401 (N_2401,In_792,In_567);
and U2402 (N_2402,In_80,In_213);
or U2403 (N_2403,In_422,In_174);
or U2404 (N_2404,In_985,In_821);
or U2405 (N_2405,In_17,In_470);
nand U2406 (N_2406,In_478,In_728);
nor U2407 (N_2407,In_426,In_563);
and U2408 (N_2408,In_844,In_576);
and U2409 (N_2409,In_848,In_153);
and U2410 (N_2410,In_660,In_998);
nor U2411 (N_2411,In_637,In_897);
or U2412 (N_2412,In_511,In_343);
and U2413 (N_2413,In_44,In_994);
nand U2414 (N_2414,In_173,In_851);
or U2415 (N_2415,In_390,In_708);
and U2416 (N_2416,In_488,In_640);
and U2417 (N_2417,In_762,In_927);
nand U2418 (N_2418,In_201,In_923);
nor U2419 (N_2419,In_251,In_981);
nand U2420 (N_2420,In_75,In_754);
nor U2421 (N_2421,In_174,In_386);
and U2422 (N_2422,In_729,In_193);
nand U2423 (N_2423,In_461,In_538);
or U2424 (N_2424,In_528,In_734);
and U2425 (N_2425,In_647,In_320);
nor U2426 (N_2426,In_837,In_104);
or U2427 (N_2427,In_10,In_913);
nor U2428 (N_2428,In_309,In_873);
nor U2429 (N_2429,In_226,In_642);
and U2430 (N_2430,In_263,In_264);
and U2431 (N_2431,In_939,In_475);
nand U2432 (N_2432,In_801,In_530);
nand U2433 (N_2433,In_948,In_397);
or U2434 (N_2434,In_51,In_396);
nand U2435 (N_2435,In_656,In_199);
nand U2436 (N_2436,In_920,In_700);
nand U2437 (N_2437,In_730,In_960);
and U2438 (N_2438,In_558,In_329);
nor U2439 (N_2439,In_610,In_871);
or U2440 (N_2440,In_991,In_570);
nor U2441 (N_2441,In_132,In_342);
and U2442 (N_2442,In_76,In_758);
and U2443 (N_2443,In_995,In_256);
or U2444 (N_2444,In_183,In_275);
nor U2445 (N_2445,In_870,In_79);
or U2446 (N_2446,In_549,In_354);
nor U2447 (N_2447,In_737,In_54);
xnor U2448 (N_2448,In_605,In_909);
and U2449 (N_2449,In_295,In_846);
nor U2450 (N_2450,In_860,In_710);
nor U2451 (N_2451,In_104,In_817);
or U2452 (N_2452,In_827,In_519);
or U2453 (N_2453,In_528,In_211);
nand U2454 (N_2454,In_214,In_721);
nor U2455 (N_2455,In_553,In_895);
and U2456 (N_2456,In_934,In_161);
nor U2457 (N_2457,In_849,In_559);
nand U2458 (N_2458,In_352,In_997);
nor U2459 (N_2459,In_218,In_201);
or U2460 (N_2460,In_718,In_117);
and U2461 (N_2461,In_89,In_123);
and U2462 (N_2462,In_224,In_731);
and U2463 (N_2463,In_867,In_17);
and U2464 (N_2464,In_297,In_637);
nor U2465 (N_2465,In_322,In_630);
and U2466 (N_2466,In_317,In_2);
xor U2467 (N_2467,In_435,In_928);
and U2468 (N_2468,In_384,In_561);
nand U2469 (N_2469,In_627,In_502);
xor U2470 (N_2470,In_810,In_897);
or U2471 (N_2471,In_123,In_739);
nand U2472 (N_2472,In_214,In_268);
or U2473 (N_2473,In_257,In_576);
or U2474 (N_2474,In_567,In_923);
nand U2475 (N_2475,In_937,In_273);
nor U2476 (N_2476,In_924,In_743);
and U2477 (N_2477,In_739,In_448);
nand U2478 (N_2478,In_971,In_705);
nand U2479 (N_2479,In_96,In_895);
nand U2480 (N_2480,In_263,In_217);
nand U2481 (N_2481,In_728,In_667);
nand U2482 (N_2482,In_67,In_303);
or U2483 (N_2483,In_727,In_720);
and U2484 (N_2484,In_758,In_185);
nor U2485 (N_2485,In_352,In_595);
and U2486 (N_2486,In_157,In_717);
nand U2487 (N_2487,In_463,In_276);
nor U2488 (N_2488,In_682,In_491);
nand U2489 (N_2489,In_559,In_339);
and U2490 (N_2490,In_324,In_477);
nand U2491 (N_2491,In_714,In_629);
and U2492 (N_2492,In_496,In_930);
or U2493 (N_2493,In_804,In_23);
nand U2494 (N_2494,In_114,In_468);
and U2495 (N_2495,In_759,In_850);
or U2496 (N_2496,In_308,In_554);
and U2497 (N_2497,In_801,In_715);
and U2498 (N_2498,In_532,In_322);
nand U2499 (N_2499,In_172,In_987);
or U2500 (N_2500,N_2469,N_1506);
nor U2501 (N_2501,N_439,N_442);
nand U2502 (N_2502,N_974,N_1073);
or U2503 (N_2503,N_1740,N_609);
nor U2504 (N_2504,N_1937,N_600);
nand U2505 (N_2505,N_1882,N_2032);
nor U2506 (N_2506,N_913,N_186);
nor U2507 (N_2507,N_177,N_2062);
or U2508 (N_2508,N_677,N_0);
nor U2509 (N_2509,N_2128,N_1888);
or U2510 (N_2510,N_11,N_565);
and U2511 (N_2511,N_1765,N_2080);
and U2512 (N_2512,N_1735,N_1807);
nand U2513 (N_2513,N_384,N_1087);
or U2514 (N_2514,N_1804,N_1507);
nor U2515 (N_2515,N_1725,N_2244);
or U2516 (N_2516,N_194,N_1139);
or U2517 (N_2517,N_589,N_1137);
nor U2518 (N_2518,N_2069,N_316);
or U2519 (N_2519,N_717,N_1384);
xnor U2520 (N_2520,N_225,N_1926);
nand U2521 (N_2521,N_2137,N_584);
nand U2522 (N_2522,N_614,N_1272);
nor U2523 (N_2523,N_860,N_727);
nand U2524 (N_2524,N_1336,N_520);
or U2525 (N_2525,N_998,N_2364);
nor U2526 (N_2526,N_1809,N_994);
or U2527 (N_2527,N_988,N_1203);
nand U2528 (N_2528,N_2278,N_1075);
nor U2529 (N_2529,N_2479,N_363);
or U2530 (N_2530,N_2210,N_2083);
or U2531 (N_2531,N_756,N_282);
nor U2532 (N_2532,N_536,N_392);
nor U2533 (N_2533,N_1520,N_104);
or U2534 (N_2534,N_1974,N_212);
nor U2535 (N_2535,N_2207,N_1291);
nor U2536 (N_2536,N_2464,N_2280);
nand U2537 (N_2537,N_2021,N_1025);
and U2538 (N_2538,N_2357,N_339);
or U2539 (N_2539,N_783,N_676);
and U2540 (N_2540,N_527,N_465);
nand U2541 (N_2541,N_823,N_160);
or U2542 (N_2542,N_619,N_2142);
and U2543 (N_2543,N_35,N_427);
and U2544 (N_2544,N_488,N_2043);
or U2545 (N_2545,N_2466,N_2475);
nor U2546 (N_2546,N_1300,N_2138);
nor U2547 (N_2547,N_1692,N_345);
nor U2548 (N_2548,N_2489,N_1685);
and U2549 (N_2549,N_134,N_256);
nor U2550 (N_2550,N_30,N_2484);
and U2551 (N_2551,N_798,N_2406);
nand U2552 (N_2552,N_963,N_406);
nor U2553 (N_2553,N_1457,N_986);
nor U2554 (N_2554,N_389,N_858);
or U2555 (N_2555,N_1340,N_458);
or U2556 (N_2556,N_2425,N_1487);
nor U2557 (N_2557,N_105,N_2426);
nor U2558 (N_2558,N_1597,N_1298);
nor U2559 (N_2559,N_1845,N_255);
nor U2560 (N_2560,N_893,N_151);
nand U2561 (N_2561,N_1800,N_976);
or U2562 (N_2562,N_71,N_461);
nor U2563 (N_2563,N_1391,N_220);
or U2564 (N_2564,N_375,N_2378);
and U2565 (N_2565,N_423,N_1026);
nand U2566 (N_2566,N_417,N_598);
or U2567 (N_2567,N_1651,N_2433);
nand U2568 (N_2568,N_208,N_1458);
and U2569 (N_2569,N_1331,N_2294);
and U2570 (N_2570,N_901,N_22);
nor U2571 (N_2571,N_94,N_1246);
and U2572 (N_2572,N_1953,N_2423);
or U2573 (N_2573,N_621,N_1895);
nor U2574 (N_2574,N_2305,N_1706);
nor U2575 (N_2575,N_2199,N_1125);
nor U2576 (N_2576,N_1642,N_254);
or U2577 (N_2577,N_1247,N_649);
or U2578 (N_2578,N_592,N_390);
nor U2579 (N_2579,N_1252,N_2350);
nand U2580 (N_2580,N_1511,N_1761);
or U2581 (N_2581,N_2122,N_4);
nand U2582 (N_2582,N_1043,N_1949);
or U2583 (N_2583,N_1283,N_2452);
and U2584 (N_2584,N_2090,N_1583);
or U2585 (N_2585,N_1635,N_814);
and U2586 (N_2586,N_2189,N_729);
nand U2587 (N_2587,N_534,N_1606);
or U2588 (N_2588,N_305,N_1756);
nor U2589 (N_2589,N_758,N_1011);
nand U2590 (N_2590,N_1158,N_968);
or U2591 (N_2591,N_583,N_1629);
nand U2592 (N_2592,N_50,N_1307);
nand U2593 (N_2593,N_1513,N_1646);
or U2594 (N_2594,N_1449,N_1748);
or U2595 (N_2595,N_1920,N_40);
nor U2596 (N_2596,N_1015,N_608);
and U2597 (N_2597,N_65,N_1205);
or U2598 (N_2598,N_663,N_1311);
nor U2599 (N_2599,N_815,N_1899);
nand U2600 (N_2600,N_2188,N_2068);
nand U2601 (N_2601,N_294,N_685);
nand U2602 (N_2602,N_492,N_1021);
and U2603 (N_2603,N_1214,N_1971);
nand U2604 (N_2604,N_856,N_2404);
and U2605 (N_2605,N_1643,N_1035);
and U2606 (N_2606,N_499,N_689);
or U2607 (N_2607,N_2456,N_1193);
and U2608 (N_2608,N_1235,N_1820);
or U2609 (N_2609,N_1058,N_1063);
nand U2610 (N_2610,N_2013,N_1950);
nand U2611 (N_2611,N_795,N_72);
xor U2612 (N_2612,N_1145,N_1489);
and U2613 (N_2613,N_890,N_1620);
or U2614 (N_2614,N_1715,N_892);
or U2615 (N_2615,N_1463,N_2389);
nor U2616 (N_2616,N_2282,N_2323);
nand U2617 (N_2617,N_914,N_2007);
nand U2618 (N_2618,N_2162,N_725);
or U2619 (N_2619,N_1051,N_484);
or U2620 (N_2620,N_1415,N_158);
or U2621 (N_2621,N_450,N_1830);
or U2622 (N_2622,N_1481,N_1818);
or U2623 (N_2623,N_191,N_1759);
and U2624 (N_2624,N_1134,N_1044);
and U2625 (N_2625,N_673,N_182);
and U2626 (N_2626,N_355,N_632);
or U2627 (N_2627,N_2024,N_1419);
nand U2628 (N_2628,N_463,N_2299);
nor U2629 (N_2629,N_928,N_1088);
nand U2630 (N_2630,N_409,N_1680);
nand U2631 (N_2631,N_2126,N_907);
and U2632 (N_2632,N_286,N_37);
and U2633 (N_2633,N_1464,N_932);
nor U2634 (N_2634,N_1929,N_1755);
or U2635 (N_2635,N_1060,N_1541);
and U2636 (N_2636,N_1873,N_195);
nor U2637 (N_2637,N_604,N_1666);
nor U2638 (N_2638,N_1209,N_1197);
and U2639 (N_2639,N_724,N_1172);
or U2640 (N_2640,N_1922,N_537);
nand U2641 (N_2641,N_2314,N_1726);
and U2642 (N_2642,N_2018,N_2451);
nor U2643 (N_2643,N_468,N_1454);
or U2644 (N_2644,N_1738,N_558);
and U2645 (N_2645,N_1448,N_1294);
or U2646 (N_2646,N_438,N_2494);
or U2647 (N_2647,N_297,N_366);
nand U2648 (N_2648,N_1285,N_425);
nor U2649 (N_2649,N_666,N_622);
nor U2650 (N_2650,N_1282,N_1713);
nor U2651 (N_2651,N_73,N_138);
and U2652 (N_2652,N_1502,N_627);
xor U2653 (N_2653,N_1909,N_1575);
or U2654 (N_2654,N_1836,N_509);
nand U2655 (N_2655,N_588,N_732);
and U2656 (N_2656,N_2407,N_760);
and U2657 (N_2657,N_1808,N_1093);
and U2658 (N_2658,N_1693,N_772);
and U2659 (N_2659,N_1844,N_1554);
nand U2660 (N_2660,N_980,N_1274);
or U2661 (N_2661,N_1912,N_1111);
or U2662 (N_2662,N_497,N_2042);
or U2663 (N_2663,N_2267,N_2316);
nor U2664 (N_2664,N_1776,N_546);
or U2665 (N_2665,N_2224,N_1020);
nor U2666 (N_2666,N_1906,N_2220);
or U2667 (N_2667,N_644,N_1592);
and U2668 (N_2668,N_1911,N_1339);
nand U2669 (N_2669,N_276,N_1704);
nand U2670 (N_2670,N_865,N_1296);
nor U2671 (N_2671,N_1128,N_1067);
or U2672 (N_2672,N_1184,N_766);
and U2673 (N_2673,N_358,N_545);
nand U2674 (N_2674,N_2387,N_1362);
nor U2675 (N_2675,N_2156,N_1112);
nand U2676 (N_2676,N_2328,N_21);
or U2677 (N_2677,N_2020,N_1736);
or U2678 (N_2678,N_629,N_623);
nor U2679 (N_2679,N_2393,N_2059);
nand U2680 (N_2680,N_213,N_187);
or U2681 (N_2681,N_2186,N_693);
and U2682 (N_2682,N_837,N_1482);
and U2683 (N_2683,N_157,N_2442);
xor U2684 (N_2684,N_557,N_999);
nor U2685 (N_2685,N_1886,N_136);
or U2686 (N_2686,N_616,N_1933);
nor U2687 (N_2687,N_1555,N_1261);
nand U2688 (N_2688,N_1517,N_2089);
and U2689 (N_2689,N_2276,N_802);
nand U2690 (N_2690,N_1013,N_242);
or U2691 (N_2691,N_926,N_1963);
nand U2692 (N_2692,N_217,N_1443);
and U2693 (N_2693,N_1492,N_209);
or U2694 (N_2694,N_1143,N_1714);
and U2695 (N_2695,N_956,N_655);
and U2696 (N_2696,N_1954,N_684);
or U2697 (N_2697,N_422,N_658);
nor U2698 (N_2698,N_934,N_2144);
or U2699 (N_2699,N_522,N_295);
nand U2700 (N_2700,N_2440,N_664);
and U2701 (N_2701,N_2394,N_1945);
and U2702 (N_2702,N_1783,N_93);
nand U2703 (N_2703,N_2490,N_1167);
nand U2704 (N_2704,N_1613,N_686);
or U2705 (N_2705,N_1497,N_2482);
nand U2706 (N_2706,N_2372,N_1418);
nand U2707 (N_2707,N_1696,N_1303);
nand U2708 (N_2708,N_768,N_743);
or U2709 (N_2709,N_1280,N_1273);
nor U2710 (N_2710,N_2071,N_1657);
and U2711 (N_2711,N_269,N_1355);
nor U2712 (N_2712,N_1897,N_357);
and U2713 (N_2713,N_1070,N_2419);
or U2714 (N_2714,N_1802,N_188);
nor U2715 (N_2715,N_749,N_1985);
or U2716 (N_2716,N_919,N_1010);
nand U2717 (N_2717,N_2367,N_1534);
nand U2718 (N_2718,N_1412,N_307);
nand U2719 (N_2719,N_1154,N_374);
or U2720 (N_2720,N_1754,N_164);
and U2721 (N_2721,N_774,N_1263);
nor U2722 (N_2722,N_778,N_1958);
nor U2723 (N_2723,N_1286,N_691);
xor U2724 (N_2724,N_1106,N_2093);
and U2725 (N_2725,N_1966,N_1442);
nand U2726 (N_2726,N_1652,N_939);
and U2727 (N_2727,N_1540,N_1728);
nor U2728 (N_2728,N_2204,N_2289);
nor U2729 (N_2729,N_739,N_1723);
or U2730 (N_2730,N_377,N_289);
or U2731 (N_2731,N_381,N_1147);
nand U2732 (N_2732,N_1784,N_1129);
nand U2733 (N_2733,N_474,N_155);
nand U2734 (N_2734,N_82,N_2315);
or U2735 (N_2735,N_2461,N_1871);
or U2736 (N_2736,N_793,N_123);
nor U2737 (N_2737,N_74,N_1787);
nand U2738 (N_2738,N_937,N_784);
or U2739 (N_2739,N_291,N_1191);
nor U2740 (N_2740,N_400,N_1762);
or U2741 (N_2741,N_311,N_76);
nor U2742 (N_2742,N_1852,N_1893);
nand U2743 (N_2743,N_1364,N_1187);
or U2744 (N_2744,N_1901,N_1894);
or U2745 (N_2745,N_1535,N_1105);
and U2746 (N_2746,N_2121,N_1424);
nor U2747 (N_2747,N_1878,N_2130);
xor U2748 (N_2748,N_957,N_1370);
nand U2749 (N_2749,N_33,N_447);
nor U2750 (N_2750,N_292,N_429);
nand U2751 (N_2751,N_183,N_1222);
and U2752 (N_2752,N_1244,N_257);
or U2753 (N_2753,N_1925,N_841);
or U2754 (N_2754,N_1121,N_962);
nand U2755 (N_2755,N_624,N_818);
and U2756 (N_2756,N_1764,N_341);
or U2757 (N_2757,N_347,N_472);
and U2758 (N_2758,N_719,N_800);
and U2759 (N_2759,N_17,N_2217);
or U2760 (N_2760,N_654,N_1265);
nand U2761 (N_2761,N_309,N_1827);
nor U2762 (N_2762,N_2408,N_748);
or U2763 (N_2763,N_2017,N_947);
nor U2764 (N_2764,N_2055,N_129);
nand U2765 (N_2765,N_1103,N_2216);
nor U2766 (N_2766,N_45,N_801);
or U2767 (N_2767,N_745,N_2439);
or U2768 (N_2768,N_1622,N_470);
or U2769 (N_2769,N_207,N_1163);
nor U2770 (N_2770,N_1039,N_809);
nand U2771 (N_2771,N_1174,N_643);
nor U2772 (N_2772,N_523,N_1310);
nor U2773 (N_2773,N_106,N_1326);
and U2774 (N_2774,N_1459,N_2281);
or U2775 (N_2775,N_834,N_933);
or U2776 (N_2776,N_1824,N_2195);
or U2777 (N_2777,N_2159,N_2275);
or U2778 (N_2778,N_2229,N_1108);
and U2779 (N_2779,N_2322,N_1014);
nor U2780 (N_2780,N_110,N_1947);
and U2781 (N_2781,N_827,N_281);
or U2782 (N_2782,N_1667,N_700);
or U2783 (N_2783,N_2252,N_1570);
nor U2784 (N_2784,N_2061,N_69);
xnor U2785 (N_2785,N_1964,N_2264);
nand U2786 (N_2786,N_1934,N_1752);
nor U2787 (N_2787,N_1055,N_1100);
nor U2788 (N_2788,N_1289,N_741);
nand U2789 (N_2789,N_1169,N_1981);
or U2790 (N_2790,N_41,N_487);
nor U2791 (N_2791,N_179,N_2338);
or U2792 (N_2792,N_2343,N_861);
or U2793 (N_2793,N_1938,N_839);
and U2794 (N_2794,N_2127,N_1879);
nand U2795 (N_2795,N_296,N_706);
nand U2796 (N_2796,N_181,N_1584);
nand U2797 (N_2797,N_787,N_174);
and U2798 (N_2798,N_993,N_1445);
nand U2799 (N_2799,N_386,N_2286);
or U2800 (N_2800,N_2180,N_451);
or U2801 (N_2801,N_280,N_2167);
and U2802 (N_2802,N_1290,N_326);
or U2803 (N_2803,N_163,N_109);
or U2804 (N_2804,N_368,N_825);
and U2805 (N_2805,N_440,N_917);
or U2806 (N_2806,N_273,N_1777);
and U2807 (N_2807,N_1078,N_385);
nor U2808 (N_2808,N_1250,N_2087);
and U2809 (N_2809,N_210,N_1375);
nor U2810 (N_2810,N_1505,N_353);
and U2811 (N_2811,N_1686,N_555);
xnor U2812 (N_2812,N_551,N_1624);
and U2813 (N_2813,N_633,N_2421);
nand U2814 (N_2814,N_1630,N_369);
nand U2815 (N_2815,N_1324,N_554);
or U2816 (N_2816,N_2164,N_1379);
nand U2817 (N_2817,N_1677,N_2014);
nor U2818 (N_2818,N_1860,N_308);
or U2819 (N_2819,N_599,N_1188);
nor U2820 (N_2820,N_1304,N_464);
nand U2821 (N_2821,N_2391,N_2073);
or U2822 (N_2822,N_1219,N_1493);
or U2823 (N_2823,N_66,N_435);
nor U2824 (N_2824,N_2066,N_2115);
nor U2825 (N_2825,N_2105,N_1293);
or U2826 (N_2826,N_1376,N_241);
nor U2827 (N_2827,N_1429,N_2190);
nor U2828 (N_2828,N_1416,N_1631);
or U2829 (N_2829,N_1413,N_2169);
and U2830 (N_2830,N_2301,N_180);
nand U2831 (N_2831,N_874,N_737);
nand U2832 (N_2832,N_1135,N_1889);
or U2833 (N_2833,N_169,N_330);
and U2834 (N_2834,N_2483,N_620);
or U2835 (N_2835,N_1936,N_2459);
nor U2836 (N_2836,N_1645,N_1159);
nor U2837 (N_2837,N_2279,N_99);
or U2838 (N_2838,N_662,N_1305);
nand U2839 (N_2839,N_2410,N_1612);
and U2840 (N_2840,N_2455,N_651);
nand U2841 (N_2841,N_279,N_984);
nand U2842 (N_2842,N_757,N_1269);
and U2843 (N_2843,N_1831,N_1395);
nand U2844 (N_2844,N_1287,N_580);
or U2845 (N_2845,N_2086,N_1607);
or U2846 (N_2846,N_652,N_1399);
nor U2847 (N_2847,N_510,N_2400);
and U2848 (N_2848,N_119,N_1773);
and U2849 (N_2849,N_2444,N_306);
and U2850 (N_2850,N_1637,N_1315);
or U2851 (N_2851,N_1733,N_694);
or U2852 (N_2852,N_596,N_1455);
nand U2853 (N_2853,N_569,N_753);
and U2854 (N_2854,N_514,N_1092);
and U2855 (N_2855,N_1072,N_1530);
or U2856 (N_2856,N_2203,N_539);
nor U2857 (N_2857,N_2385,N_637);
nor U2858 (N_2858,N_2476,N_263);
or U2859 (N_2859,N_2182,N_2390);
and U2860 (N_2860,N_2249,N_108);
and U2861 (N_2861,N_2392,N_638);
and U2862 (N_2862,N_1790,N_819);
nand U2863 (N_2863,N_246,N_981);
nor U2864 (N_2864,N_2245,N_462);
nand U2865 (N_2865,N_1373,N_2472);
and U2866 (N_2866,N_713,N_1732);
nor U2867 (N_2867,N_971,N_1967);
nor U2868 (N_2868,N_1385,N_805);
nor U2869 (N_2869,N_1335,N_2260);
xor U2870 (N_2870,N_1970,N_1718);
nor U2871 (N_2871,N_1891,N_228);
and U2872 (N_2872,N_343,N_1392);
nand U2873 (N_2873,N_1245,N_1120);
nand U2874 (N_2874,N_990,N_2006);
or U2875 (N_2875,N_457,N_211);
nand U2876 (N_2876,N_2165,N_1450);
nand U2877 (N_2877,N_587,N_2099);
nor U2878 (N_2878,N_722,N_875);
and U2879 (N_2879,N_404,N_873);
nand U2880 (N_2880,N_2430,N_421);
nor U2881 (N_2881,N_2349,N_236);
nor U2882 (N_2882,N_121,N_1348);
nor U2883 (N_2883,N_333,N_53);
nand U2884 (N_2884,N_2376,N_1545);
and U2885 (N_2885,N_262,N_921);
or U2886 (N_2886,N_361,N_1593);
nand U2887 (N_2887,N_1533,N_991);
or U2888 (N_2888,N_475,N_1835);
nor U2889 (N_2889,N_1608,N_2236);
and U2890 (N_2890,N_2211,N_786);
or U2891 (N_2891,N_1959,N_92);
xor U2892 (N_2892,N_2306,N_1037);
and U2893 (N_2893,N_641,N_1354);
nand U2894 (N_2894,N_1236,N_2037);
and U2895 (N_2895,N_416,N_192);
and U2896 (N_2896,N_1708,N_172);
and U2897 (N_2897,N_1192,N_2);
nand U2898 (N_2898,N_578,N_635);
nor U2899 (N_2899,N_1647,N_1898);
and U2900 (N_2900,N_2074,N_2172);
nand U2901 (N_2901,N_1536,N_266);
nor U2902 (N_2902,N_2434,N_915);
nor U2903 (N_2903,N_2424,N_2302);
nor U2904 (N_2904,N_1052,N_251);
and U2905 (N_2905,N_1504,N_518);
or U2906 (N_2906,N_1080,N_1655);
and U2907 (N_2907,N_1869,N_1863);
or U2908 (N_2908,N_1007,N_55);
xor U2909 (N_2909,N_657,N_525);
or U2910 (N_2910,N_460,N_1832);
nor U2911 (N_2911,N_2076,N_1915);
or U2912 (N_2912,N_1525,N_1550);
and U2913 (N_2913,N_1817,N_86);
nand U2914 (N_2914,N_1356,N_2320);
xor U2915 (N_2915,N_1242,N_1956);
and U2916 (N_2916,N_1737,N_36);
nor U2917 (N_2917,N_1665,N_153);
nand U2918 (N_2918,N_543,N_1903);
or U2919 (N_2919,N_43,N_313);
nor U2920 (N_2920,N_2183,N_1485);
nor U2921 (N_2921,N_2317,N_770);
nor U2922 (N_2922,N_1478,N_653);
nand U2923 (N_2923,N_2191,N_337);
nand U2924 (N_2924,N_1779,N_77);
nor U2925 (N_2925,N_852,N_2246);
nand U2926 (N_2926,N_1019,N_101);
and U2927 (N_2927,N_989,N_965);
nand U2928 (N_2928,N_1609,N_2341);
nand U2929 (N_2929,N_1578,N_1634);
or U2930 (N_2930,N_720,N_348);
nand U2931 (N_2931,N_942,N_293);
nand U2932 (N_2932,N_38,N_883);
xnor U2933 (N_2933,N_2096,N_1381);
nand U2934 (N_2934,N_849,N_1008);
and U2935 (N_2935,N_1856,N_1476);
or U2936 (N_2936,N_1678,N_2187);
or U2937 (N_2937,N_1268,N_1644);
or U2938 (N_2938,N_2432,N_1576);
and U2939 (N_2939,N_2497,N_1202);
or U2940 (N_2940,N_1460,N_1695);
nor U2941 (N_2941,N_1679,N_319);
nor U2942 (N_2942,N_453,N_755);
nor U2943 (N_2943,N_2227,N_1372);
nor U2944 (N_2944,N_1386,N_1004);
nand U2945 (N_2945,N_1470,N_1102);
and U2946 (N_2946,N_2103,N_1997);
nor U2947 (N_2947,N_1230,N_196);
or U2948 (N_2948,N_1965,N_324);
or U2949 (N_2949,N_200,N_2234);
nor U2950 (N_2950,N_1743,N_1491);
and U2951 (N_2951,N_2292,N_1700);
nand U2952 (N_2952,N_647,N_762);
or U2953 (N_2953,N_120,N_707);
nor U2954 (N_2954,N_709,N_1683);
nand U2955 (N_2955,N_561,N_1232);
xor U2956 (N_2956,N_1278,N_1890);
nand U2957 (N_2957,N_603,N_1027);
xor U2958 (N_2958,N_1982,N_1430);
nand U2959 (N_2959,N_2222,N_173);
or U2960 (N_2960,N_205,N_935);
or U2961 (N_2961,N_740,N_137);
nand U2962 (N_2962,N_1472,N_167);
nand U2963 (N_2963,N_714,N_1900);
xor U2964 (N_2964,N_1420,N_227);
nor U2965 (N_2965,N_322,N_265);
xor U2966 (N_2966,N_233,N_350);
and U2967 (N_2967,N_1594,N_1603);
or U2968 (N_2968,N_1212,N_1018);
and U2969 (N_2969,N_1640,N_2088);
or U2970 (N_2970,N_1774,N_864);
nand U2971 (N_2971,N_1249,N_1140);
nor U2972 (N_2972,N_1320,N_821);
nor U2973 (N_2973,N_408,N_2051);
nor U2974 (N_2974,N_1164,N_1234);
nor U2975 (N_2975,N_2303,N_244);
nor U2976 (N_2976,N_1876,N_734);
nor U2977 (N_2977,N_391,N_1739);
nand U2978 (N_2978,N_1514,N_2208);
and U2979 (N_2979,N_27,N_2300);
or U2980 (N_2980,N_1330,N_387);
nand U2981 (N_2981,N_202,N_9);
and U2982 (N_2982,N_738,N_176);
and U2983 (N_2983,N_1266,N_781);
nand U2984 (N_2984,N_2354,N_1864);
or U2985 (N_2985,N_832,N_1149);
nor U2986 (N_2986,N_2241,N_171);
nor U2987 (N_2987,N_2257,N_1819);
nor U2988 (N_2988,N_2492,N_2272);
or U2989 (N_2989,N_1763,N_746);
nand U2990 (N_2990,N_446,N_2369);
or U2991 (N_2991,N_334,N_1799);
or U2992 (N_2992,N_1377,N_1941);
or U2993 (N_2993,N_2250,N_1849);
or U2994 (N_2994,N_143,N_2095);
nand U2995 (N_2995,N_1874,N_2049);
and U2996 (N_2996,N_1024,N_576);
nand U2997 (N_2997,N_1091,N_2136);
nor U2998 (N_2998,N_1892,N_672);
nand U2999 (N_2999,N_742,N_1798);
nor U3000 (N_3000,N_28,N_2005);
and U3001 (N_3001,N_1224,N_1671);
nand U3002 (N_3002,N_1099,N_969);
or U3003 (N_3003,N_512,N_49);
nand U3004 (N_3004,N_1940,N_564);
nand U3005 (N_3005,N_1569,N_631);
and U3006 (N_3006,N_659,N_1337);
and U3007 (N_3007,N_2064,N_1617);
nor U3008 (N_3008,N_904,N_1987);
nand U3009 (N_3009,N_103,N_2102);
nand U3010 (N_3010,N_591,N_1730);
xor U3011 (N_3011,N_1760,N_2200);
or U3012 (N_3012,N_1257,N_977);
xor U3013 (N_3013,N_1838,N_1387);
and U3014 (N_3014,N_2101,N_1626);
or U3015 (N_3015,N_1297,N_2397);
nor U3016 (N_3016,N_2336,N_1851);
or U3017 (N_3017,N_1368,N_661);
or U3018 (N_3018,N_1907,N_145);
and U3019 (N_3019,N_2319,N_411);
nor U3020 (N_3020,N_1117,N_2048);
nor U3021 (N_3021,N_154,N_2325);
nand U3022 (N_3022,N_8,N_2462);
and U3023 (N_3023,N_848,N_2449);
or U3024 (N_3024,N_2015,N_1213);
nor U3025 (N_3025,N_733,N_3);
or U3026 (N_3026,N_776,N_1623);
and U3027 (N_3027,N_2332,N_586);
nand U3028 (N_3028,N_2375,N_701);
and U3029 (N_3029,N_2358,N_648);
nor U3030 (N_3030,N_2178,N_547);
nor U3031 (N_3031,N_476,N_1902);
or U3032 (N_3032,N_790,N_765);
nor U3033 (N_3033,N_2181,N_70);
or U3034 (N_3034,N_1281,N_1488);
or U3035 (N_3035,N_1582,N_581);
nor U3036 (N_3036,N_204,N_95);
nand U3037 (N_3037,N_1532,N_48);
nor U3038 (N_3038,N_16,N_113);
and U3039 (N_3039,N_290,N_1896);
or U3040 (N_3040,N_2114,N_185);
and U3041 (N_3041,N_975,N_1208);
nand U3042 (N_3042,N_668,N_2185);
nand U3043 (N_3043,N_1223,N_301);
nor U3044 (N_3044,N_607,N_2333);
or U3045 (N_3045,N_2431,N_13);
or U3046 (N_3046,N_1215,N_1432);
or U3047 (N_3047,N_304,N_1453);
xor U3048 (N_3048,N_57,N_2238);
nand U3049 (N_3049,N_215,N_1986);
nor U3050 (N_3050,N_885,N_529);
and U3051 (N_3051,N_1309,N_606);
nor U3052 (N_3052,N_230,N_1618);
nor U3053 (N_3053,N_2176,N_826);
nor U3054 (N_3054,N_1401,N_2395);
and U3055 (N_3055,N_615,N_354);
or U3056 (N_3056,N_1133,N_1277);
or U3057 (N_3057,N_1833,N_797);
nor U3058 (N_3058,N_247,N_2386);
nor U3059 (N_3059,N_2356,N_221);
nand U3060 (N_3060,N_2453,N_1227);
nor U3061 (N_3061,N_81,N_1961);
or U3062 (N_3062,N_199,N_133);
nand U3063 (N_3063,N_1029,N_2151);
and U3064 (N_3064,N_436,N_1341);
or U3065 (N_3065,N_415,N_1322);
and U3066 (N_3066,N_495,N_853);
nand U3067 (N_3067,N_549,N_1423);
nor U3068 (N_3068,N_494,N_2415);
or U3069 (N_3069,N_1116,N_2065);
nor U3070 (N_3070,N_443,N_1753);
or U3071 (N_3071,N_1402,N_336);
nand U3072 (N_3072,N_1983,N_47);
or U3073 (N_3073,N_822,N_1688);
or U3074 (N_3074,N_894,N_862);
or U3075 (N_3075,N_918,N_32);
and U3076 (N_3076,N_1181,N_1495);
xnor U3077 (N_3077,N_1621,N_502);
or U3078 (N_3078,N_521,N_2310);
nor U3079 (N_3079,N_261,N_107);
and U3080 (N_3080,N_1255,N_329);
or U3081 (N_3081,N_1825,N_1334);
and U3082 (N_3082,N_1927,N_1744);
nor U3083 (N_3083,N_1747,N_1012);
nand U3084 (N_3084,N_2119,N_2417);
nor U3085 (N_3085,N_857,N_538);
xor U3086 (N_3086,N_20,N_640);
or U3087 (N_3087,N_639,N_238);
nand U3088 (N_3088,N_1564,N_1132);
nand U3089 (N_3089,N_871,N_2486);
or U3090 (N_3090,N_838,N_115);
and U3091 (N_3091,N_506,N_466);
nor U3092 (N_3092,N_2171,N_1600);
and U3093 (N_3093,N_2324,N_1095);
nand U3094 (N_3094,N_1467,N_2437);
nand U3095 (N_3095,N_1829,N_660);
or U3096 (N_3096,N_1358,N_2329);
or U3097 (N_3097,N_1360,N_730);
or U3098 (N_3098,N_708,N_886);
nand U3099 (N_3099,N_2379,N_367);
and U3100 (N_3100,N_1332,N_2077);
and U3101 (N_3101,N_2111,N_595);
or U3102 (N_3102,N_277,N_1796);
nor U3103 (N_3103,N_1789,N_2174);
nand U3104 (N_3104,N_2226,N_1653);
nor U3105 (N_3105,N_1975,N_1840);
or U3106 (N_3106,N_2152,N_1539);
nor U3107 (N_3107,N_1699,N_1639);
or U3108 (N_3108,N_597,N_2031);
or U3109 (N_3109,N_877,N_1812);
and U3110 (N_3110,N_2420,N_1049);
or U3111 (N_3111,N_1544,N_83);
or U3112 (N_3112,N_131,N_2100);
nor U3113 (N_3113,N_424,N_1867);
and U3114 (N_3114,N_274,N_2063);
nor U3115 (N_3115,N_1681,N_1703);
and U3116 (N_3116,N_785,N_895);
and U3117 (N_3117,N_1248,N_2273);
nor U3118 (N_3118,N_2034,N_419);
and U3119 (N_3119,N_2135,N_1880);
and U3120 (N_3120,N_1302,N_548);
nor U3121 (N_3121,N_1705,N_1742);
or U3122 (N_3122,N_252,N_1500);
or U3123 (N_3123,N_150,N_1923);
or U3124 (N_3124,N_80,N_754);
nor U3125 (N_3125,N_2265,N_1910);
nand U3126 (N_3126,N_26,N_1451);
or U3127 (N_3127,N_165,N_888);
nand U3128 (N_3128,N_29,N_1085);
or U3129 (N_3129,N_1847,N_1691);
or U3130 (N_3130,N_1628,N_1727);
or U3131 (N_3131,N_1148,N_1673);
nand U3132 (N_3132,N_1225,N_590);
and U3133 (N_3133,N_1846,N_490);
nor U3134 (N_3134,N_444,N_2163);
or U3135 (N_3135,N_1171,N_328);
or U3136 (N_3136,N_489,N_1096);
nor U3137 (N_3137,N_2277,N_2027);
nand U3138 (N_3138,N_949,N_2344);
nand U3139 (N_3139,N_690,N_1960);
or U3140 (N_3140,N_1082,N_2283);
nand U3141 (N_3141,N_231,N_2262);
or U3142 (N_3142,N_63,N_2327);
nor U3143 (N_3143,N_1327,N_1206);
or U3144 (N_3144,N_2471,N_91);
or U3145 (N_3145,N_2029,N_567);
xor U3146 (N_3146,N_764,N_454);
nand U3147 (N_3147,N_2113,N_2012);
nand U3148 (N_3148,N_1510,N_382);
nand U3149 (N_3149,N_51,N_1397);
or U3150 (N_3150,N_842,N_1862);
nand U3151 (N_3151,N_61,N_432);
or U3152 (N_3152,N_1059,N_1389);
nand U3153 (N_3153,N_1587,N_310);
nor U3154 (N_3154,N_2384,N_594);
or U3155 (N_3155,N_950,N_922);
nand U3156 (N_3156,N_613,N_1857);
nor U3157 (N_3157,N_298,N_248);
nor U3158 (N_3158,N_1267,N_500);
and U3159 (N_3159,N_346,N_605);
nor U3160 (N_3160,N_1750,N_2374);
or U3161 (N_3161,N_1408,N_1547);
nand U3162 (N_3162,N_831,N_1130);
nand U3163 (N_3163,N_2269,N_2457);
or U3164 (N_3164,N_397,N_1674);
nor U3165 (N_3165,N_718,N_1444);
and U3166 (N_3166,N_1041,N_1183);
and U3167 (N_3167,N_2271,N_433);
xnor U3168 (N_3168,N_528,N_1233);
nor U3169 (N_3169,N_201,N_1076);
and U3170 (N_3170,N_2003,N_1690);
nor U3171 (N_3171,N_1904,N_1426);
nand U3172 (N_3172,N_315,N_1745);
nor U3173 (N_3173,N_1259,N_370);
nand U3174 (N_3174,N_2498,N_1660);
or U3175 (N_3175,N_127,N_2296);
and U3176 (N_3176,N_1791,N_2118);
nand U3177 (N_3177,N_1196,N_278);
nand U3178 (N_3178,N_1042,N_721);
nor U3179 (N_3179,N_373,N_1931);
nand U3180 (N_3180,N_1394,N_1988);
nor U3181 (N_3181,N_2362,N_1369);
nand U3182 (N_3182,N_1056,N_2155);
nand U3183 (N_3183,N_2078,N_847);
or U3184 (N_3184,N_1995,N_1839);
or U3185 (N_3185,N_559,N_7);
and U3186 (N_3186,N_2075,N_2041);
and U3187 (N_3187,N_1345,N_1684);
or U3188 (N_3188,N_2237,N_1383);
or U3189 (N_3189,N_1552,N_1317);
or U3190 (N_3190,N_1425,N_945);
or U3191 (N_3191,N_1295,N_898);
xor U3192 (N_3192,N_2402,N_232);
or U3193 (N_3193,N_1538,N_486);
xor U3194 (N_3194,N_1207,N_840);
nor U3195 (N_3195,N_1329,N_1074);
or U3196 (N_3196,N_1546,N_2291);
nor U3197 (N_3197,N_1712,N_2295);
and U3198 (N_3198,N_1741,N_953);
nand U3199 (N_3199,N_1016,N_1284);
and U3200 (N_3200,N_2033,N_130);
or U3201 (N_3201,N_1301,N_941);
nand U3202 (N_3202,N_2438,N_6);
and U3203 (N_3203,N_1841,N_1185);
or U3204 (N_3204,N_1580,N_1720);
and U3205 (N_3205,N_2468,N_688);
or U3206 (N_3206,N_1328,N_190);
or U3207 (N_3207,N_479,N_1405);
nand U3208 (N_3208,N_2487,N_1722);
nor U3209 (N_3209,N_1153,N_2219);
nand U3210 (N_3210,N_2057,N_2359);
nand U3211 (N_3211,N_2470,N_1537);
and U3212 (N_3212,N_156,N_2184);
nor U3213 (N_3213,N_936,N_1664);
nand U3214 (N_3214,N_1241,N_1932);
and U3215 (N_3215,N_2107,N_900);
and U3216 (N_3216,N_517,N_1853);
nand U3217 (N_3217,N_1469,N_1176);
and U3218 (N_3218,N_2092,N_1319);
nand U3219 (N_3219,N_1884,N_2266);
or U3220 (N_3220,N_1471,N_206);
and U3221 (N_3221,N_1151,N_891);
nor U3222 (N_3222,N_1930,N_759);
nor U3223 (N_3223,N_1406,N_1299);
or U3224 (N_3224,N_2478,N_1556);
nand U3225 (N_3225,N_1687,N_1486);
xor U3226 (N_3226,N_2230,N_1553);
and U3227 (N_3227,N_752,N_1437);
and U3228 (N_3228,N_1479,N_1905);
nor U3229 (N_3229,N_2290,N_723);
nor U3230 (N_3230,N_650,N_1589);
or U3231 (N_3231,N_493,N_909);
and U3232 (N_3232,N_910,N_882);
or U3233 (N_3233,N_1611,N_866);
or U3234 (N_3234,N_1670,N_747);
and U3235 (N_3235,N_237,N_698);
nor U3236 (N_3236,N_782,N_2496);
nor U3237 (N_3237,N_1939,N_1211);
nand U3238 (N_3238,N_2120,N_2082);
or U3239 (N_3239,N_380,N_2212);
and U3240 (N_3240,N_1136,N_2435);
nor U3241 (N_3241,N_2416,N_132);
and U3242 (N_3242,N_1000,N_1398);
and U3243 (N_3243,N_1990,N_1661);
nor U3244 (N_3244,N_869,N_412);
and U3245 (N_3245,N_2148,N_2366);
nand U3246 (N_3246,N_2373,N_1276);
and U3247 (N_3247,N_1483,N_360);
nor U3248 (N_3248,N_1872,N_1079);
or U3249 (N_3249,N_1976,N_828);
and U3250 (N_3250,N_1568,N_2331);
and U3251 (N_3251,N_418,N_2345);
nand U3252 (N_3252,N_1101,N_830);
and U3253 (N_3253,N_259,N_964);
nand U3254 (N_3254,N_62,N_1821);
and U3255 (N_3255,N_601,N_1758);
nand U3256 (N_3256,N_1175,N_2150);
or U3257 (N_3257,N_511,N_1549);
nor U3258 (N_3258,N_1676,N_2412);
nand U3259 (N_3259,N_2427,N_703);
nand U3260 (N_3260,N_229,N_2117);
nand U3261 (N_3261,N_98,N_162);
and U3262 (N_3262,N_626,N_944);
or U3263 (N_3263,N_321,N_1516);
or U3264 (N_3264,N_1484,N_14);
and U3265 (N_3265,N_1313,N_1162);
or U3266 (N_3266,N_2428,N_1349);
and U3267 (N_3267,N_25,N_340);
nor U3268 (N_3268,N_1731,N_807);
nor U3269 (N_3269,N_630,N_887);
or U3270 (N_3270,N_2110,N_572);
or U3271 (N_3271,N_2084,N_2218);
nor U3272 (N_3272,N_2247,N_498);
nor U3273 (N_3273,N_1751,N_1573);
nand U3274 (N_3274,N_1746,N_2312);
or U3275 (N_3275,N_515,N_2193);
and U3276 (N_3276,N_112,N_1881);
nand U3277 (N_3277,N_1127,N_923);
nand U3278 (N_3278,N_1770,N_264);
nand U3279 (N_3279,N_2170,N_2154);
and U3280 (N_3280,N_1672,N_351);
and U3281 (N_3281,N_19,N_2382);
and U3282 (N_3282,N_970,N_966);
nand U3283 (N_3283,N_1475,N_929);
and U3284 (N_3284,N_2153,N_982);
nor U3285 (N_3285,N_1201,N_780);
and U3286 (N_3286,N_2044,N_480);
or U3287 (N_3287,N_2477,N_1709);
or U3288 (N_3288,N_1599,N_1757);
nor U3289 (N_3289,N_1081,N_1619);
nor U3290 (N_3290,N_1574,N_302);
nor U3291 (N_3291,N_2481,N_2405);
nand U3292 (N_3292,N_1456,N_34);
and U3293 (N_3293,N_855,N_1396);
xor U3294 (N_3294,N_2141,N_1438);
or U3295 (N_3295,N_1256,N_716);
and U3296 (N_3296,N_562,N_2008);
and U3297 (N_3297,N_2243,N_2206);
nor U3298 (N_3298,N_312,N_532);
or U3299 (N_3299,N_912,N_833);
or U3300 (N_3300,N_1501,N_2258);
nor U3301 (N_3301,N_2140,N_526);
nor U3302 (N_3302,N_1957,N_1523);
and U3303 (N_3303,N_1795,N_2287);
nor U3304 (N_3304,N_1654,N_2388);
nor U3305 (N_3305,N_87,N_2240);
nor U3306 (N_3306,N_1031,N_1338);
nand U3307 (N_3307,N_193,N_152);
nand U3308 (N_3308,N_2205,N_1778);
nor U3309 (N_3309,N_1615,N_471);
nor U3310 (N_3310,N_2371,N_2360);
or U3311 (N_3311,N_1916,N_288);
and U3312 (N_3312,N_1682,N_1969);
nand U3313 (N_3313,N_2039,N_1913);
and U3314 (N_3314,N_1165,N_2253);
or U3315 (N_3315,N_67,N_1788);
nor U3316 (N_3316,N_2129,N_253);
and U3317 (N_3317,N_1144,N_820);
or U3318 (N_3318,N_249,N_574);
nand U3319 (N_3319,N_1367,N_985);
and U3320 (N_3320,N_473,N_835);
or U3321 (N_3321,N_449,N_140);
nand U3322 (N_3322,N_1865,N_1104);
or U3323 (N_3323,N_2132,N_582);
or U3324 (N_3324,N_1382,N_958);
nand U3325 (N_3325,N_602,N_2177);
or U3326 (N_3326,N_338,N_1919);
or U3327 (N_3327,N_44,N_593);
or U3328 (N_3328,N_2403,N_680);
or U3329 (N_3329,N_751,N_1566);
or U3330 (N_3330,N_961,N_1194);
nor U3331 (N_3331,N_379,N_478);
or U3332 (N_3332,N_2436,N_1033);
and U3333 (N_3333,N_712,N_349);
or U3334 (N_3334,N_2368,N_2488);
nor U3335 (N_3335,N_1887,N_1400);
nand U3336 (N_3336,N_359,N_2318);
nand U3337 (N_3337,N_2004,N_2175);
nand U3338 (N_3338,N_2214,N_284);
and U3339 (N_3339,N_642,N_1989);
nor U3340 (N_3340,N_799,N_184);
or U3341 (N_3341,N_2108,N_222);
and U3342 (N_3342,N_198,N_362);
nor U3343 (N_3343,N_75,N_1602);
nor U3344 (N_3344,N_906,N_166);
nand U3345 (N_3345,N_2070,N_2396);
nor U3346 (N_3346,N_2256,N_482);
and U3347 (N_3347,N_836,N_667);
and U3348 (N_3348,N_2019,N_553);
nand U3349 (N_3349,N_1526,N_1077);
nand U3350 (N_3350,N_2288,N_1388);
or U3351 (N_3351,N_1859,N_58);
and U3352 (N_3352,N_2067,N_1199);
nor U3353 (N_3353,N_791,N_1001);
and U3354 (N_3354,N_88,N_1694);
nand U3355 (N_3355,N_1498,N_144);
nand U3356 (N_3356,N_1883,N_983);
and U3357 (N_3357,N_711,N_1123);
or U3358 (N_3358,N_1404,N_2337);
and U3359 (N_3359,N_1823,N_1480);
or U3360 (N_3360,N_459,N_2228);
and U3361 (N_3361,N_1801,N_1002);
nand U3362 (N_3362,N_1238,N_2016);
nand U3363 (N_3363,N_1633,N_203);
or U3364 (N_3364,N_808,N_496);
and U3365 (N_3365,N_2146,N_2198);
or U3366 (N_3366,N_1993,N_1198);
or U3367 (N_3367,N_2401,N_804);
nand U3368 (N_3368,N_430,N_491);
and U3369 (N_3369,N_1239,N_1858);
and U3370 (N_3370,N_2454,N_1581);
or U3371 (N_3371,N_736,N_1527);
or U3372 (N_3372,N_611,N_1979);
nand U3373 (N_3373,N_1614,N_1048);
or U3374 (N_3374,N_775,N_1109);
or U3375 (N_3375,N_2270,N_441);
and U3376 (N_3376,N_2157,N_2334);
and U3377 (N_3377,N_1107,N_1343);
or U3378 (N_3378,N_2010,N_1772);
nor U3379 (N_3379,N_656,N_2340);
and U3380 (N_3380,N_135,N_2284);
or U3381 (N_3381,N_1084,N_1962);
or U3382 (N_3382,N_1781,N_2352);
or U3383 (N_3383,N_1040,N_1279);
or U3384 (N_3384,N_1407,N_960);
nand U3385 (N_3385,N_335,N_102);
and U3386 (N_3386,N_452,N_1032);
nand U3387 (N_3387,N_530,N_2197);
nor U3388 (N_3388,N_1689,N_1275);
nand U3389 (N_3389,N_388,N_1022);
nand U3390 (N_3390,N_1638,N_1353);
nor U3391 (N_3391,N_1854,N_1697);
nor U3392 (N_3392,N_533,N_556);
and U3393 (N_3393,N_2465,N_318);
or U3394 (N_3394,N_1509,N_2035);
nor U3395 (N_3395,N_2473,N_2098);
nand U3396 (N_3396,N_1089,N_1782);
or U3397 (N_3397,N_1441,N_1503);
or U3398 (N_3398,N_1822,N_851);
nor U3399 (N_3399,N_405,N_704);
nor U3400 (N_3400,N_979,N_695);
or U3401 (N_3401,N_1610,N_2339);
nand U3402 (N_3402,N_1944,N_448);
nand U3403 (N_3403,N_1494,N_2480);
and U3404 (N_3404,N_1216,N_1598);
or U3405 (N_3405,N_407,N_414);
nor U3406 (N_3406,N_1034,N_868);
and U3407 (N_3407,N_159,N_967);
or U3408 (N_3408,N_1605,N_1561);
nand U3409 (N_3409,N_2124,N_125);
xnor U3410 (N_3410,N_1409,N_846);
nand U3411 (N_3411,N_897,N_1724);
nor U3412 (N_3412,N_816,N_2399);
nand U3413 (N_3413,N_1585,N_1124);
nand U3414 (N_3414,N_1625,N_744);
and U3415 (N_3415,N_2450,N_372);
and U3416 (N_3416,N_467,N_2125);
and U3417 (N_3417,N_1071,N_97);
and U3418 (N_3418,N_258,N_1814);
nor U3419 (N_3419,N_122,N_796);
nand U3420 (N_3420,N_1766,N_1528);
nand U3421 (N_3421,N_2202,N_1806);
nor U3422 (N_3422,N_610,N_2409);
nor U3423 (N_3423,N_1179,N_323);
and U3424 (N_3424,N_1427,N_617);
nor U3425 (N_3425,N_485,N_1924);
nand U3426 (N_3426,N_788,N_1411);
or U3427 (N_3427,N_1943,N_1359);
nor U3428 (N_3428,N_930,N_2297);
nand U3429 (N_3429,N_1543,N_12);
nor U3430 (N_3430,N_46,N_39);
and U3431 (N_3431,N_1204,N_342);
nand U3432 (N_3432,N_1237,N_2248);
or U3433 (N_3433,N_902,N_1146);
or U3434 (N_3434,N_767,N_117);
and U3435 (N_3435,N_434,N_1057);
or U3436 (N_3436,N_997,N_1542);
nor U3437 (N_3437,N_1551,N_1436);
nor U3438 (N_3438,N_750,N_1734);
nor U3439 (N_3439,N_1499,N_1308);
nand U3440 (N_3440,N_168,N_2441);
nor U3441 (N_3441,N_1361,N_1521);
or U3442 (N_3442,N_777,N_899);
nand U3443 (N_3443,N_2221,N_1115);
or U3444 (N_3444,N_1254,N_817);
nor U3445 (N_3445,N_1050,N_1166);
or U3446 (N_3446,N_2139,N_1371);
nor U3447 (N_3447,N_1565,N_728);
and U3448 (N_3448,N_671,N_1984);
nor U3449 (N_3449,N_1721,N_1999);
or U3450 (N_3450,N_469,N_995);
nand U3451 (N_3451,N_1160,N_761);
or U3452 (N_3452,N_2255,N_2028);
nand U3453 (N_3453,N_1529,N_1870);
nor U3454 (N_3454,N_1170,N_715);
nor U3455 (N_3455,N_1342,N_1908);
nor U3456 (N_3456,N_1119,N_1918);
nand U3457 (N_3457,N_669,N_2046);
nand U3458 (N_3458,N_1632,N_1951);
and U3459 (N_3459,N_1098,N_2231);
and U3460 (N_3460,N_175,N_1769);
nor U3461 (N_3461,N_1921,N_271);
nor U3462 (N_3462,N_2443,N_2307);
and U3463 (N_3463,N_1243,N_1186);
nand U3464 (N_3464,N_161,N_519);
and U3465 (N_3465,N_15,N_1054);
and U3466 (N_3466,N_779,N_911);
nand U3467 (N_3467,N_878,N_1251);
nor U3468 (N_3468,N_1531,N_1793);
or U3469 (N_3469,N_331,N_697);
and U3470 (N_3470,N_2000,N_1113);
or U3471 (N_3471,N_566,N_18);
nand U3472 (N_3472,N_1161,N_2149);
and U3473 (N_3473,N_2050,N_2448);
and U3474 (N_3474,N_1837,N_954);
nor U3475 (N_3475,N_952,N_332);
and U3476 (N_3476,N_674,N_2134);
and U3477 (N_3477,N_1352,N_612);
nor U3478 (N_3478,N_1710,N_1262);
nand U3479 (N_3479,N_844,N_1935);
nand U3480 (N_3480,N_428,N_2104);
nor U3481 (N_3481,N_735,N_2009);
nand U3482 (N_3482,N_2145,N_2311);
nand U3483 (N_3483,N_535,N_938);
nor U3484 (N_3484,N_223,N_1562);
and U3485 (N_3485,N_1711,N_905);
nor U3486 (N_3486,N_560,N_1228);
and U3487 (N_3487,N_24,N_769);
or U3488 (N_3488,N_111,N_1118);
nor U3489 (N_3489,N_2085,N_996);
nor U3490 (N_3490,N_2225,N_1805);
nor U3491 (N_3491,N_1811,N_683);
or U3492 (N_3492,N_2213,N_5);
and U3493 (N_3493,N_682,N_1131);
nand U3494 (N_3494,N_675,N_1955);
and U3495 (N_3495,N_56,N_1595);
nor U3496 (N_3496,N_2274,N_903);
nor U3497 (N_3497,N_889,N_299);
and U3498 (N_3498,N_1195,N_1659);
or U3499 (N_3499,N_678,N_563);
and U3500 (N_3500,N_1767,N_1466);
nor U3501 (N_3501,N_1452,N_1948);
nor U3502 (N_3502,N_410,N_413);
and U3503 (N_3503,N_1972,N_763);
nor U3504 (N_3504,N_2094,N_1240);
or U3505 (N_3505,N_726,N_2351);
nor U3506 (N_3506,N_1157,N_1351);
or U3507 (N_3507,N_1428,N_1434);
nand U3508 (N_3508,N_1519,N_1559);
and U3509 (N_3509,N_189,N_1828);
nor U3510 (N_3510,N_925,N_1698);
and U3511 (N_3511,N_1596,N_1097);
nand U3512 (N_3512,N_1473,N_1771);
and U3513 (N_3513,N_2251,N_1604);
nor U3514 (N_3514,N_1142,N_1810);
and U3515 (N_3515,N_812,N_420);
and U3516 (N_3516,N_1843,N_2235);
or U3517 (N_3517,N_52,N_2383);
or U3518 (N_3518,N_287,N_1270);
or U3519 (N_3519,N_1155,N_702);
or U3520 (N_3520,N_645,N_2414);
and U3521 (N_3521,N_2091,N_2147);
or U3522 (N_3522,N_1522,N_1992);
nand U3523 (N_3523,N_356,N_829);
and U3524 (N_3524,N_2022,N_618);
or U3525 (N_3525,N_2458,N_170);
nor U3526 (N_3526,N_1462,N_1446);
nand U3527 (N_3527,N_573,N_139);
or U3528 (N_3528,N_940,N_68);
and U3529 (N_3529,N_1220,N_2040);
or U3530 (N_3530,N_1226,N_224);
nor U3531 (N_3531,N_503,N_1928);
nand U3532 (N_3532,N_78,N_2268);
and U3533 (N_3533,N_2418,N_31);
nor U3534 (N_3534,N_2030,N_1586);
nand U3535 (N_3535,N_1422,N_2036);
nor U3536 (N_3536,N_1816,N_916);
or U3537 (N_3537,N_2321,N_1558);
nand U3538 (N_3538,N_64,N_1288);
nand U3539 (N_3539,N_142,N_399);
nor U3540 (N_3540,N_2348,N_2168);
and U3541 (N_3541,N_426,N_810);
nor U3542 (N_3542,N_1946,N_1333);
nand U3543 (N_3543,N_285,N_1068);
and U3544 (N_3544,N_505,N_1065);
and U3545 (N_3545,N_1182,N_1156);
or U3546 (N_3546,N_1390,N_696);
nand U3547 (N_3547,N_456,N_710);
or U3548 (N_3548,N_1729,N_872);
and U3549 (N_3549,N_1180,N_1114);
or U3550 (N_3550,N_1508,N_1563);
and U3551 (N_3551,N_395,N_1572);
nor U3552 (N_3552,N_585,N_1260);
and U3553 (N_3553,N_275,N_1577);
and U3554 (N_3554,N_1998,N_845);
and U3555 (N_3555,N_1036,N_501);
xnor U3556 (N_3556,N_1421,N_1649);
nor U3557 (N_3557,N_84,N_1658);
nand U3558 (N_3558,N_1346,N_2232);
nor U3559 (N_3559,N_141,N_2411);
and U3560 (N_3560,N_2056,N_2233);
or U3561 (N_3561,N_1431,N_243);
xor U3562 (N_3562,N_881,N_1591);
and U3563 (N_3563,N_524,N_1834);
nor U3564 (N_3564,N_2365,N_114);
nand U3565 (N_3565,N_234,N_2097);
nand U3566 (N_3566,N_402,N_1749);
and U3567 (N_3567,N_1440,N_2353);
or U3568 (N_3568,N_531,N_625);
xor U3569 (N_3569,N_2161,N_2377);
nand U3570 (N_3570,N_2370,N_867);
or U3571 (N_3571,N_1023,N_1177);
nor U3572 (N_3572,N_1548,N_1090);
or U3573 (N_3573,N_2047,N_575);
or U3574 (N_3574,N_1062,N_2446);
and U3575 (N_3575,N_544,N_2326);
nor U3576 (N_3576,N_1868,N_1557);
or U3577 (N_3577,N_1006,N_687);
nand U3578 (N_3578,N_1496,N_1465);
nand U3579 (N_3579,N_2143,N_1061);
and U3580 (N_3580,N_214,N_283);
nor U3581 (N_3581,N_568,N_541);
nor U3582 (N_3582,N_1028,N_2467);
xor U3583 (N_3583,N_863,N_1588);
nor U3584 (N_3584,N_2447,N_2158);
nor U3585 (N_3585,N_1866,N_1579);
and U3586 (N_3586,N_383,N_2261);
or U3587 (N_3587,N_550,N_2045);
nand U3588 (N_3588,N_116,N_2079);
or U3589 (N_3589,N_1848,N_972);
nor U3590 (N_3590,N_1217,N_1785);
or U3591 (N_3591,N_245,N_219);
and U3592 (N_3592,N_178,N_1264);
and U3593 (N_3593,N_1813,N_705);
or U3594 (N_3594,N_477,N_1797);
or U3595 (N_3595,N_268,N_218);
nor U3596 (N_3596,N_1292,N_226);
nor U3597 (N_3597,N_1417,N_1768);
or U3598 (N_3598,N_128,N_42);
and U3599 (N_3599,N_1656,N_2485);
or U3600 (N_3600,N_1258,N_2499);
nor U3601 (N_3601,N_1786,N_260);
and U3602 (N_3602,N_992,N_670);
nor U3603 (N_3603,N_973,N_1590);
nor U3604 (N_3604,N_118,N_1323);
nor U3605 (N_3605,N_146,N_1347);
or U3606 (N_3606,N_2285,N_1150);
or U3607 (N_3607,N_327,N_2106);
and U3608 (N_3608,N_1627,N_2001);
or U3609 (N_3609,N_79,N_1173);
and U3610 (N_3610,N_1447,N_1168);
nor U3611 (N_3611,N_314,N_1318);
nor U3612 (N_3612,N_2363,N_1403);
nor U3613 (N_3613,N_959,N_955);
and U3614 (N_3614,N_636,N_2112);
xnor U3615 (N_3615,N_1378,N_59);
and U3616 (N_3616,N_393,N_2422);
nor U3617 (N_3617,N_1468,N_1086);
nand U3618 (N_3618,N_850,N_571);
nand U3619 (N_3619,N_927,N_2002);
and U3620 (N_3620,N_2026,N_1321);
and U3621 (N_3621,N_1005,N_811);
or U3622 (N_3622,N_2474,N_508);
nand U3623 (N_3623,N_646,N_1325);
nor U3624 (N_3624,N_876,N_1662);
or U3625 (N_3625,N_1792,N_792);
nand U3626 (N_3626,N_1474,N_2330);
or U3627 (N_3627,N_1190,N_481);
nor U3628 (N_3628,N_1009,N_250);
and U3629 (N_3629,N_437,N_1775);
or U3630 (N_3630,N_2166,N_2025);
nand U3631 (N_3631,N_681,N_1312);
nand U3632 (N_3632,N_124,N_1122);
or U3633 (N_3633,N_378,N_445);
nor U3634 (N_3634,N_924,N_1571);
nor U3635 (N_3635,N_2131,N_2058);
or U3636 (N_3636,N_2060,N_731);
xnor U3637 (N_3637,N_665,N_1363);
and U3638 (N_3638,N_325,N_2160);
and U3639 (N_3639,N_90,N_1877);
or U3640 (N_3640,N_2081,N_1030);
nand U3641 (N_3641,N_2298,N_978);
or U3642 (N_3642,N_1366,N_240);
nor U3643 (N_3643,N_946,N_1842);
nand U3644 (N_3644,N_1229,N_579);
and U3645 (N_3645,N_2335,N_1701);
xnor U3646 (N_3646,N_96,N_1719);
or U3647 (N_3647,N_1410,N_854);
nor U3648 (N_3648,N_1875,N_1231);
and U3649 (N_3649,N_1046,N_272);
or U3650 (N_3650,N_2192,N_806);
nand U3651 (N_3651,N_2346,N_1973);
xor U3652 (N_3652,N_2038,N_364);
and U3653 (N_3653,N_1861,N_1914);
nand U3654 (N_3654,N_1414,N_2123);
nand U3655 (N_3655,N_2309,N_1126);
xnor U3656 (N_3656,N_2313,N_147);
nand U3657 (N_3657,N_2133,N_1942);
nor U3658 (N_3658,N_239,N_824);
and U3659 (N_3659,N_2116,N_2429);
and U3660 (N_3660,N_54,N_376);
or U3661 (N_3661,N_1567,N_896);
xor U3662 (N_3662,N_1094,N_1641);
or U3663 (N_3663,N_1616,N_1306);
nand U3664 (N_3664,N_1991,N_344);
or U3665 (N_3665,N_1707,N_789);
and U3666 (N_3666,N_2381,N_2380);
or U3667 (N_3667,N_2242,N_1053);
nor U3668 (N_3668,N_2052,N_2263);
nand U3669 (N_3669,N_843,N_1668);
and U3670 (N_3670,N_1850,N_126);
nor U3671 (N_3671,N_2011,N_403);
nor U3672 (N_3672,N_431,N_2398);
and U3673 (N_3673,N_2413,N_1200);
nor U3674 (N_3674,N_1780,N_1045);
or U3675 (N_3675,N_197,N_1461);
nand U3676 (N_3676,N_516,N_60);
nand U3677 (N_3677,N_1917,N_773);
and U3678 (N_3678,N_1271,N_1210);
nor U3679 (N_3679,N_692,N_1003);
and U3680 (N_3680,N_1433,N_813);
nand U3681 (N_3681,N_2259,N_1110);
nor U3682 (N_3682,N_1996,N_1515);
or U3683 (N_3683,N_483,N_1968);
or U3684 (N_3684,N_1980,N_1017);
nor U3685 (N_3685,N_948,N_2355);
or U3686 (N_3686,N_1350,N_2053);
nand U3687 (N_3687,N_23,N_1702);
nand U3688 (N_3688,N_699,N_317);
nand U3689 (N_3689,N_148,N_1675);
nand U3690 (N_3690,N_1994,N_1189);
nor U3691 (N_3691,N_1344,N_879);
nor U3692 (N_3692,N_1038,N_1435);
and U3693 (N_3693,N_85,N_552);
and U3694 (N_3694,N_859,N_2308);
nand U3695 (N_3695,N_1512,N_2493);
nor U3696 (N_3696,N_1141,N_870);
or U3697 (N_3697,N_2491,N_2179);
nand U3698 (N_3698,N_1663,N_1393);
nand U3699 (N_3699,N_794,N_398);
nand U3700 (N_3700,N_2342,N_1138);
or U3701 (N_3701,N_2347,N_507);
or U3702 (N_3702,N_2361,N_908);
or U3703 (N_3703,N_1316,N_10);
nand U3704 (N_3704,N_2196,N_1650);
and U3705 (N_3705,N_270,N_1490);
or U3706 (N_3706,N_396,N_1855);
nor U3707 (N_3707,N_1978,N_1439);
nor U3708 (N_3708,N_1066,N_1815);
nor U3709 (N_3709,N_2215,N_300);
and U3710 (N_3710,N_1826,N_1560);
nor U3711 (N_3711,N_1069,N_634);
nor U3712 (N_3712,N_371,N_540);
nor U3713 (N_3713,N_1152,N_880);
nand U3714 (N_3714,N_1977,N_1357);
and U3715 (N_3715,N_1221,N_267);
nor U3716 (N_3716,N_2445,N_504);
and U3717 (N_3717,N_2239,N_2460);
or U3718 (N_3718,N_394,N_577);
xor U3719 (N_3719,N_1601,N_2173);
or U3720 (N_3720,N_1794,N_931);
and U3721 (N_3721,N_1374,N_1477);
or U3722 (N_3722,N_943,N_1047);
nor U3723 (N_3723,N_1178,N_1218);
nor U3724 (N_3724,N_803,N_216);
nand U3725 (N_3725,N_1365,N_1380);
nor U3726 (N_3726,N_1064,N_570);
or U3727 (N_3727,N_2463,N_89);
and U3728 (N_3728,N_1648,N_1);
nor U3729 (N_3729,N_2254,N_149);
xnor U3730 (N_3730,N_1518,N_352);
or U3731 (N_3731,N_513,N_920);
or U3732 (N_3732,N_2072,N_2201);
nor U3733 (N_3733,N_2054,N_303);
and U3734 (N_3734,N_1669,N_2109);
and U3735 (N_3735,N_1636,N_1083);
nand U3736 (N_3736,N_2304,N_1314);
or U3737 (N_3737,N_1803,N_951);
or U3738 (N_3738,N_235,N_542);
or U3739 (N_3739,N_320,N_771);
nand U3740 (N_3740,N_455,N_1717);
and U3741 (N_3741,N_2495,N_987);
nor U3742 (N_3742,N_1716,N_2023);
or U3743 (N_3743,N_679,N_2209);
and U3744 (N_3744,N_100,N_628);
and U3745 (N_3745,N_365,N_2194);
nand U3746 (N_3746,N_401,N_1524);
nand U3747 (N_3747,N_1952,N_2293);
xor U3748 (N_3748,N_884,N_2223);
and U3749 (N_3749,N_1885,N_1253);
nor U3750 (N_3750,N_1642,N_1037);
xnor U3751 (N_3751,N_2287,N_2259);
and U3752 (N_3752,N_2240,N_1420);
nor U3753 (N_3753,N_1955,N_382);
nand U3754 (N_3754,N_848,N_1655);
or U3755 (N_3755,N_1814,N_2063);
nand U3756 (N_3756,N_132,N_115);
and U3757 (N_3757,N_1451,N_927);
or U3758 (N_3758,N_1841,N_2030);
nand U3759 (N_3759,N_837,N_1262);
and U3760 (N_3760,N_1639,N_1338);
nor U3761 (N_3761,N_499,N_922);
or U3762 (N_3762,N_1256,N_719);
and U3763 (N_3763,N_2499,N_1728);
nor U3764 (N_3764,N_1937,N_190);
nand U3765 (N_3765,N_1747,N_641);
or U3766 (N_3766,N_1512,N_55);
or U3767 (N_3767,N_1208,N_1918);
and U3768 (N_3768,N_516,N_173);
nor U3769 (N_3769,N_1227,N_2429);
nand U3770 (N_3770,N_1743,N_2401);
nor U3771 (N_3771,N_2040,N_318);
and U3772 (N_3772,N_619,N_1630);
nand U3773 (N_3773,N_1797,N_2183);
nand U3774 (N_3774,N_25,N_247);
or U3775 (N_3775,N_306,N_723);
nand U3776 (N_3776,N_2022,N_1321);
nor U3777 (N_3777,N_1426,N_706);
nor U3778 (N_3778,N_203,N_1032);
and U3779 (N_3779,N_1546,N_1477);
or U3780 (N_3780,N_762,N_1763);
nand U3781 (N_3781,N_1714,N_381);
nor U3782 (N_3782,N_655,N_241);
nand U3783 (N_3783,N_273,N_2388);
and U3784 (N_3784,N_2343,N_849);
and U3785 (N_3785,N_1889,N_1044);
and U3786 (N_3786,N_1427,N_1765);
nand U3787 (N_3787,N_815,N_2206);
nor U3788 (N_3788,N_1969,N_115);
or U3789 (N_3789,N_462,N_2100);
and U3790 (N_3790,N_2278,N_107);
nand U3791 (N_3791,N_618,N_1379);
xnor U3792 (N_3792,N_1026,N_1528);
and U3793 (N_3793,N_1136,N_2451);
nand U3794 (N_3794,N_886,N_1206);
nor U3795 (N_3795,N_676,N_1290);
or U3796 (N_3796,N_107,N_639);
or U3797 (N_3797,N_746,N_904);
or U3798 (N_3798,N_1678,N_91);
and U3799 (N_3799,N_2208,N_2284);
nor U3800 (N_3800,N_1616,N_2387);
and U3801 (N_3801,N_1414,N_912);
and U3802 (N_3802,N_2167,N_2194);
or U3803 (N_3803,N_363,N_760);
and U3804 (N_3804,N_1534,N_799);
nor U3805 (N_3805,N_215,N_945);
or U3806 (N_3806,N_590,N_791);
nand U3807 (N_3807,N_192,N_374);
nand U3808 (N_3808,N_787,N_1454);
nor U3809 (N_3809,N_1075,N_157);
or U3810 (N_3810,N_1334,N_856);
and U3811 (N_3811,N_345,N_388);
nor U3812 (N_3812,N_2433,N_627);
nand U3813 (N_3813,N_2259,N_1340);
nor U3814 (N_3814,N_2032,N_1533);
nand U3815 (N_3815,N_964,N_1372);
nor U3816 (N_3816,N_929,N_1024);
nand U3817 (N_3817,N_1478,N_2274);
nor U3818 (N_3818,N_19,N_1749);
nor U3819 (N_3819,N_59,N_1068);
and U3820 (N_3820,N_2407,N_2321);
and U3821 (N_3821,N_1583,N_1099);
nor U3822 (N_3822,N_1190,N_2490);
nor U3823 (N_3823,N_1236,N_2490);
or U3824 (N_3824,N_400,N_2288);
and U3825 (N_3825,N_1447,N_508);
or U3826 (N_3826,N_361,N_427);
or U3827 (N_3827,N_359,N_492);
nor U3828 (N_3828,N_271,N_1688);
nor U3829 (N_3829,N_613,N_1869);
or U3830 (N_3830,N_967,N_2084);
or U3831 (N_3831,N_2451,N_17);
and U3832 (N_3832,N_732,N_2160);
nand U3833 (N_3833,N_328,N_2354);
or U3834 (N_3834,N_1708,N_391);
or U3835 (N_3835,N_203,N_391);
or U3836 (N_3836,N_763,N_984);
nor U3837 (N_3837,N_2314,N_2102);
nor U3838 (N_3838,N_903,N_1323);
or U3839 (N_3839,N_2387,N_1507);
or U3840 (N_3840,N_529,N_332);
nand U3841 (N_3841,N_1687,N_452);
or U3842 (N_3842,N_1003,N_844);
and U3843 (N_3843,N_654,N_353);
nand U3844 (N_3844,N_1995,N_2093);
nand U3845 (N_3845,N_1501,N_505);
or U3846 (N_3846,N_2216,N_2207);
nand U3847 (N_3847,N_1206,N_807);
or U3848 (N_3848,N_1341,N_1683);
nor U3849 (N_3849,N_113,N_1931);
or U3850 (N_3850,N_1037,N_1127);
or U3851 (N_3851,N_1419,N_2202);
or U3852 (N_3852,N_1449,N_439);
or U3853 (N_3853,N_1447,N_206);
nand U3854 (N_3854,N_815,N_1673);
nor U3855 (N_3855,N_1789,N_1560);
or U3856 (N_3856,N_445,N_1407);
nand U3857 (N_3857,N_1784,N_1326);
nor U3858 (N_3858,N_668,N_1038);
and U3859 (N_3859,N_1599,N_596);
and U3860 (N_3860,N_1736,N_738);
and U3861 (N_3861,N_103,N_886);
or U3862 (N_3862,N_1575,N_943);
nor U3863 (N_3863,N_2397,N_1205);
nand U3864 (N_3864,N_1447,N_1846);
nand U3865 (N_3865,N_1838,N_556);
nand U3866 (N_3866,N_982,N_551);
and U3867 (N_3867,N_1238,N_2044);
or U3868 (N_3868,N_332,N_51);
or U3869 (N_3869,N_118,N_1135);
nand U3870 (N_3870,N_2365,N_692);
and U3871 (N_3871,N_860,N_1679);
nand U3872 (N_3872,N_963,N_890);
nor U3873 (N_3873,N_306,N_207);
and U3874 (N_3874,N_375,N_1356);
nor U3875 (N_3875,N_681,N_1237);
nor U3876 (N_3876,N_1220,N_1531);
nor U3877 (N_3877,N_1399,N_2375);
nand U3878 (N_3878,N_301,N_809);
or U3879 (N_3879,N_2218,N_1153);
nor U3880 (N_3880,N_287,N_926);
or U3881 (N_3881,N_623,N_648);
nor U3882 (N_3882,N_2073,N_455);
and U3883 (N_3883,N_1397,N_757);
or U3884 (N_3884,N_1314,N_2380);
nand U3885 (N_3885,N_102,N_62);
or U3886 (N_3886,N_738,N_599);
and U3887 (N_3887,N_468,N_2351);
or U3888 (N_3888,N_476,N_1377);
and U3889 (N_3889,N_1539,N_2201);
nor U3890 (N_3890,N_342,N_2395);
nor U3891 (N_3891,N_2261,N_54);
nor U3892 (N_3892,N_1557,N_2447);
nor U3893 (N_3893,N_702,N_1632);
and U3894 (N_3894,N_2452,N_2071);
nand U3895 (N_3895,N_2266,N_671);
nand U3896 (N_3896,N_1428,N_1785);
nor U3897 (N_3897,N_832,N_2368);
nand U3898 (N_3898,N_1097,N_2445);
nor U3899 (N_3899,N_41,N_8);
or U3900 (N_3900,N_701,N_196);
and U3901 (N_3901,N_1665,N_1702);
nand U3902 (N_3902,N_1828,N_755);
nand U3903 (N_3903,N_1823,N_378);
nor U3904 (N_3904,N_2128,N_2116);
nor U3905 (N_3905,N_23,N_157);
nand U3906 (N_3906,N_634,N_882);
and U3907 (N_3907,N_1853,N_2228);
and U3908 (N_3908,N_885,N_1198);
and U3909 (N_3909,N_802,N_1440);
and U3910 (N_3910,N_184,N_2426);
nand U3911 (N_3911,N_2043,N_593);
nor U3912 (N_3912,N_2375,N_636);
nand U3913 (N_3913,N_2405,N_162);
nand U3914 (N_3914,N_195,N_964);
or U3915 (N_3915,N_206,N_1830);
or U3916 (N_3916,N_1854,N_277);
or U3917 (N_3917,N_855,N_1016);
and U3918 (N_3918,N_1332,N_1255);
xor U3919 (N_3919,N_1103,N_1353);
nand U3920 (N_3920,N_301,N_721);
and U3921 (N_3921,N_2444,N_1033);
nand U3922 (N_3922,N_1146,N_194);
nand U3923 (N_3923,N_2031,N_1000);
and U3924 (N_3924,N_906,N_1171);
and U3925 (N_3925,N_2235,N_111);
or U3926 (N_3926,N_1069,N_1330);
xnor U3927 (N_3927,N_696,N_2150);
nor U3928 (N_3928,N_1348,N_1365);
xnor U3929 (N_3929,N_847,N_1966);
nand U3930 (N_3930,N_1166,N_703);
xor U3931 (N_3931,N_2082,N_915);
nand U3932 (N_3932,N_1121,N_1020);
nor U3933 (N_3933,N_680,N_1499);
nand U3934 (N_3934,N_1688,N_937);
nand U3935 (N_3935,N_2021,N_2108);
or U3936 (N_3936,N_2498,N_1411);
nand U3937 (N_3937,N_383,N_247);
nand U3938 (N_3938,N_1878,N_1639);
or U3939 (N_3939,N_1045,N_1957);
nand U3940 (N_3940,N_577,N_1907);
nand U3941 (N_3941,N_943,N_1541);
xor U3942 (N_3942,N_2231,N_1243);
nand U3943 (N_3943,N_2,N_870);
or U3944 (N_3944,N_2022,N_1450);
nand U3945 (N_3945,N_1123,N_1483);
or U3946 (N_3946,N_509,N_2439);
nor U3947 (N_3947,N_276,N_357);
nand U3948 (N_3948,N_582,N_235);
and U3949 (N_3949,N_4,N_468);
and U3950 (N_3950,N_12,N_1407);
xor U3951 (N_3951,N_1430,N_2297);
or U3952 (N_3952,N_327,N_602);
nand U3953 (N_3953,N_1846,N_1990);
and U3954 (N_3954,N_104,N_2210);
nand U3955 (N_3955,N_1107,N_2303);
nand U3956 (N_3956,N_939,N_1233);
or U3957 (N_3957,N_140,N_872);
xor U3958 (N_3958,N_2337,N_1918);
or U3959 (N_3959,N_1566,N_428);
and U3960 (N_3960,N_2428,N_2185);
or U3961 (N_3961,N_765,N_221);
or U3962 (N_3962,N_90,N_1817);
or U3963 (N_3963,N_1051,N_2466);
nand U3964 (N_3964,N_864,N_2111);
nand U3965 (N_3965,N_109,N_1172);
nand U3966 (N_3966,N_468,N_1307);
and U3967 (N_3967,N_741,N_2123);
xnor U3968 (N_3968,N_1338,N_855);
and U3969 (N_3969,N_2092,N_1102);
or U3970 (N_3970,N_1689,N_1647);
or U3971 (N_3971,N_149,N_586);
nand U3972 (N_3972,N_2246,N_1580);
and U3973 (N_3973,N_2350,N_663);
and U3974 (N_3974,N_163,N_1547);
and U3975 (N_3975,N_1425,N_1828);
or U3976 (N_3976,N_1972,N_601);
and U3977 (N_3977,N_1266,N_529);
nor U3978 (N_3978,N_1731,N_1626);
and U3979 (N_3979,N_1561,N_2120);
or U3980 (N_3980,N_1018,N_1635);
or U3981 (N_3981,N_601,N_1447);
nor U3982 (N_3982,N_1304,N_156);
nor U3983 (N_3983,N_2310,N_1398);
nor U3984 (N_3984,N_133,N_1662);
nand U3985 (N_3985,N_2417,N_344);
nor U3986 (N_3986,N_1227,N_943);
nor U3987 (N_3987,N_1996,N_590);
or U3988 (N_3988,N_408,N_1802);
nand U3989 (N_3989,N_333,N_1197);
nand U3990 (N_3990,N_241,N_1913);
or U3991 (N_3991,N_1579,N_1465);
nand U3992 (N_3992,N_1286,N_48);
or U3993 (N_3993,N_354,N_1597);
nor U3994 (N_3994,N_506,N_1595);
nor U3995 (N_3995,N_351,N_52);
and U3996 (N_3996,N_2420,N_738);
or U3997 (N_3997,N_1226,N_114);
nand U3998 (N_3998,N_1253,N_1093);
and U3999 (N_3999,N_411,N_1814);
and U4000 (N_4000,N_2036,N_194);
xor U4001 (N_4001,N_2433,N_565);
and U4002 (N_4002,N_1595,N_1653);
nor U4003 (N_4003,N_2173,N_1855);
and U4004 (N_4004,N_1132,N_227);
nor U4005 (N_4005,N_81,N_876);
or U4006 (N_4006,N_1484,N_2102);
nor U4007 (N_4007,N_1009,N_494);
and U4008 (N_4008,N_435,N_2010);
nor U4009 (N_4009,N_1039,N_1563);
and U4010 (N_4010,N_498,N_1645);
nor U4011 (N_4011,N_274,N_1453);
nand U4012 (N_4012,N_1379,N_476);
nor U4013 (N_4013,N_1160,N_1514);
nand U4014 (N_4014,N_449,N_1279);
or U4015 (N_4015,N_389,N_146);
and U4016 (N_4016,N_815,N_1184);
nand U4017 (N_4017,N_1101,N_2274);
and U4018 (N_4018,N_134,N_1153);
nor U4019 (N_4019,N_2491,N_1284);
and U4020 (N_4020,N_2119,N_412);
or U4021 (N_4021,N_1905,N_795);
nand U4022 (N_4022,N_1539,N_9);
and U4023 (N_4023,N_1090,N_945);
nand U4024 (N_4024,N_965,N_793);
or U4025 (N_4025,N_2293,N_1263);
nand U4026 (N_4026,N_36,N_927);
xor U4027 (N_4027,N_817,N_158);
or U4028 (N_4028,N_2368,N_1722);
or U4029 (N_4029,N_1247,N_104);
or U4030 (N_4030,N_2356,N_2065);
and U4031 (N_4031,N_252,N_1668);
or U4032 (N_4032,N_1639,N_623);
nor U4033 (N_4033,N_1797,N_108);
and U4034 (N_4034,N_2379,N_567);
nor U4035 (N_4035,N_394,N_850);
nand U4036 (N_4036,N_860,N_2413);
nand U4037 (N_4037,N_2406,N_260);
nand U4038 (N_4038,N_1981,N_279);
and U4039 (N_4039,N_273,N_210);
nand U4040 (N_4040,N_187,N_147);
and U4041 (N_4041,N_1885,N_2219);
and U4042 (N_4042,N_1898,N_310);
nand U4043 (N_4043,N_1788,N_1498);
nand U4044 (N_4044,N_1422,N_1931);
nor U4045 (N_4045,N_1789,N_1276);
nor U4046 (N_4046,N_464,N_1798);
or U4047 (N_4047,N_743,N_2459);
or U4048 (N_4048,N_1191,N_300);
and U4049 (N_4049,N_1536,N_497);
and U4050 (N_4050,N_1057,N_24);
nand U4051 (N_4051,N_1573,N_8);
or U4052 (N_4052,N_917,N_955);
nand U4053 (N_4053,N_349,N_847);
nor U4054 (N_4054,N_1994,N_2130);
nor U4055 (N_4055,N_1388,N_1162);
nand U4056 (N_4056,N_200,N_1639);
nand U4057 (N_4057,N_2445,N_1457);
nor U4058 (N_4058,N_1772,N_1452);
or U4059 (N_4059,N_1291,N_677);
or U4060 (N_4060,N_681,N_814);
or U4061 (N_4061,N_834,N_774);
nor U4062 (N_4062,N_61,N_2172);
or U4063 (N_4063,N_129,N_760);
and U4064 (N_4064,N_181,N_1044);
nand U4065 (N_4065,N_2355,N_1256);
or U4066 (N_4066,N_1313,N_1967);
and U4067 (N_4067,N_2129,N_2400);
nand U4068 (N_4068,N_817,N_1067);
or U4069 (N_4069,N_1360,N_1983);
and U4070 (N_4070,N_1504,N_1973);
and U4071 (N_4071,N_1391,N_786);
nand U4072 (N_4072,N_449,N_213);
nand U4073 (N_4073,N_2046,N_540);
nand U4074 (N_4074,N_198,N_1908);
nor U4075 (N_4075,N_1561,N_1484);
or U4076 (N_4076,N_2174,N_1200);
nand U4077 (N_4077,N_1048,N_1490);
or U4078 (N_4078,N_270,N_207);
xnor U4079 (N_4079,N_728,N_1426);
or U4080 (N_4080,N_251,N_850);
and U4081 (N_4081,N_1579,N_474);
and U4082 (N_4082,N_1040,N_2068);
nor U4083 (N_4083,N_1669,N_910);
or U4084 (N_4084,N_119,N_123);
nor U4085 (N_4085,N_962,N_1600);
and U4086 (N_4086,N_2204,N_1842);
and U4087 (N_4087,N_1405,N_1511);
or U4088 (N_4088,N_19,N_1559);
nor U4089 (N_4089,N_1714,N_1505);
nor U4090 (N_4090,N_1774,N_800);
or U4091 (N_4091,N_366,N_607);
nand U4092 (N_4092,N_209,N_2192);
and U4093 (N_4093,N_607,N_1729);
nor U4094 (N_4094,N_684,N_80);
nand U4095 (N_4095,N_929,N_151);
or U4096 (N_4096,N_170,N_47);
or U4097 (N_4097,N_1941,N_185);
and U4098 (N_4098,N_727,N_2152);
and U4099 (N_4099,N_1532,N_2119);
nand U4100 (N_4100,N_228,N_366);
nand U4101 (N_4101,N_2183,N_790);
nor U4102 (N_4102,N_1246,N_1335);
and U4103 (N_4103,N_2056,N_709);
nand U4104 (N_4104,N_1997,N_1467);
or U4105 (N_4105,N_97,N_2181);
nor U4106 (N_4106,N_2330,N_902);
or U4107 (N_4107,N_205,N_1462);
nor U4108 (N_4108,N_1002,N_1191);
and U4109 (N_4109,N_1870,N_1211);
nor U4110 (N_4110,N_2459,N_2441);
nor U4111 (N_4111,N_1563,N_2080);
and U4112 (N_4112,N_1905,N_697);
or U4113 (N_4113,N_1620,N_1680);
and U4114 (N_4114,N_1504,N_1726);
xnor U4115 (N_4115,N_1884,N_1106);
nand U4116 (N_4116,N_764,N_930);
nor U4117 (N_4117,N_2362,N_850);
nor U4118 (N_4118,N_1739,N_294);
nor U4119 (N_4119,N_1220,N_635);
or U4120 (N_4120,N_2473,N_1145);
nand U4121 (N_4121,N_1052,N_1503);
and U4122 (N_4122,N_1025,N_2418);
and U4123 (N_4123,N_686,N_1433);
and U4124 (N_4124,N_758,N_1393);
nand U4125 (N_4125,N_561,N_213);
and U4126 (N_4126,N_1763,N_1499);
nor U4127 (N_4127,N_518,N_965);
or U4128 (N_4128,N_1570,N_35);
or U4129 (N_4129,N_1951,N_2310);
nand U4130 (N_4130,N_1460,N_983);
nand U4131 (N_4131,N_1158,N_1771);
nand U4132 (N_4132,N_1917,N_470);
or U4133 (N_4133,N_2081,N_1037);
nor U4134 (N_4134,N_312,N_153);
nand U4135 (N_4135,N_592,N_1000);
xor U4136 (N_4136,N_505,N_2488);
xor U4137 (N_4137,N_87,N_999);
nor U4138 (N_4138,N_582,N_689);
or U4139 (N_4139,N_299,N_2311);
nor U4140 (N_4140,N_283,N_1256);
and U4141 (N_4141,N_1170,N_843);
or U4142 (N_4142,N_1490,N_930);
nor U4143 (N_4143,N_926,N_1353);
nand U4144 (N_4144,N_1542,N_623);
nand U4145 (N_4145,N_1591,N_1382);
or U4146 (N_4146,N_2239,N_1017);
nor U4147 (N_4147,N_1571,N_971);
and U4148 (N_4148,N_663,N_1679);
and U4149 (N_4149,N_2263,N_1168);
nand U4150 (N_4150,N_1122,N_1451);
xor U4151 (N_4151,N_2360,N_474);
nand U4152 (N_4152,N_1903,N_2098);
nand U4153 (N_4153,N_2234,N_1366);
and U4154 (N_4154,N_1317,N_1923);
nand U4155 (N_4155,N_1489,N_1572);
nor U4156 (N_4156,N_2371,N_967);
nand U4157 (N_4157,N_1081,N_1030);
nand U4158 (N_4158,N_2300,N_900);
nand U4159 (N_4159,N_1796,N_1386);
nor U4160 (N_4160,N_2239,N_1789);
and U4161 (N_4161,N_597,N_1420);
or U4162 (N_4162,N_1379,N_219);
and U4163 (N_4163,N_2176,N_201);
or U4164 (N_4164,N_790,N_170);
or U4165 (N_4165,N_69,N_575);
nand U4166 (N_4166,N_419,N_1838);
or U4167 (N_4167,N_2238,N_581);
nand U4168 (N_4168,N_2033,N_1233);
nand U4169 (N_4169,N_2416,N_1607);
nor U4170 (N_4170,N_364,N_1991);
or U4171 (N_4171,N_1288,N_1920);
and U4172 (N_4172,N_2178,N_332);
nand U4173 (N_4173,N_733,N_1494);
nor U4174 (N_4174,N_999,N_1854);
nand U4175 (N_4175,N_1201,N_1818);
nand U4176 (N_4176,N_1035,N_173);
and U4177 (N_4177,N_425,N_1372);
or U4178 (N_4178,N_1755,N_853);
and U4179 (N_4179,N_1865,N_2242);
nand U4180 (N_4180,N_2495,N_260);
nor U4181 (N_4181,N_2335,N_638);
nand U4182 (N_4182,N_95,N_2124);
nor U4183 (N_4183,N_1830,N_2380);
and U4184 (N_4184,N_2168,N_58);
nand U4185 (N_4185,N_1664,N_2016);
or U4186 (N_4186,N_1171,N_1134);
or U4187 (N_4187,N_1514,N_2465);
or U4188 (N_4188,N_2186,N_1837);
and U4189 (N_4189,N_781,N_1290);
and U4190 (N_4190,N_2489,N_885);
and U4191 (N_4191,N_1737,N_1776);
or U4192 (N_4192,N_1035,N_2085);
nor U4193 (N_4193,N_2079,N_1894);
and U4194 (N_4194,N_1455,N_537);
or U4195 (N_4195,N_945,N_508);
or U4196 (N_4196,N_1019,N_2381);
and U4197 (N_4197,N_446,N_2235);
nor U4198 (N_4198,N_1734,N_1179);
and U4199 (N_4199,N_1226,N_1509);
and U4200 (N_4200,N_1543,N_2211);
or U4201 (N_4201,N_2071,N_1025);
nand U4202 (N_4202,N_887,N_1965);
and U4203 (N_4203,N_1865,N_845);
nor U4204 (N_4204,N_1997,N_166);
and U4205 (N_4205,N_781,N_980);
or U4206 (N_4206,N_1224,N_972);
and U4207 (N_4207,N_316,N_1889);
nand U4208 (N_4208,N_689,N_276);
nand U4209 (N_4209,N_295,N_1860);
nor U4210 (N_4210,N_354,N_629);
xor U4211 (N_4211,N_1247,N_1653);
or U4212 (N_4212,N_1963,N_1341);
or U4213 (N_4213,N_1452,N_1296);
nor U4214 (N_4214,N_340,N_23);
nand U4215 (N_4215,N_1158,N_920);
nand U4216 (N_4216,N_1283,N_1899);
or U4217 (N_4217,N_162,N_2449);
and U4218 (N_4218,N_186,N_205);
and U4219 (N_4219,N_1938,N_542);
or U4220 (N_4220,N_120,N_2185);
nand U4221 (N_4221,N_1269,N_2478);
or U4222 (N_4222,N_1867,N_191);
or U4223 (N_4223,N_1841,N_1578);
nor U4224 (N_4224,N_1609,N_1151);
and U4225 (N_4225,N_720,N_773);
and U4226 (N_4226,N_2314,N_1418);
nor U4227 (N_4227,N_848,N_393);
nand U4228 (N_4228,N_671,N_56);
or U4229 (N_4229,N_1892,N_893);
and U4230 (N_4230,N_2170,N_177);
or U4231 (N_4231,N_2035,N_734);
nand U4232 (N_4232,N_1468,N_466);
and U4233 (N_4233,N_2360,N_1288);
nand U4234 (N_4234,N_1267,N_1442);
or U4235 (N_4235,N_1548,N_467);
nand U4236 (N_4236,N_500,N_879);
or U4237 (N_4237,N_1212,N_1238);
or U4238 (N_4238,N_1391,N_2365);
nor U4239 (N_4239,N_2059,N_2101);
and U4240 (N_4240,N_1075,N_1986);
or U4241 (N_4241,N_578,N_1831);
nor U4242 (N_4242,N_56,N_1097);
and U4243 (N_4243,N_706,N_1269);
nand U4244 (N_4244,N_1197,N_503);
nand U4245 (N_4245,N_698,N_2084);
nor U4246 (N_4246,N_2384,N_2377);
nand U4247 (N_4247,N_1910,N_2280);
and U4248 (N_4248,N_1590,N_1123);
nand U4249 (N_4249,N_310,N_1736);
xnor U4250 (N_4250,N_630,N_2400);
or U4251 (N_4251,N_1499,N_1007);
nand U4252 (N_4252,N_414,N_1050);
nor U4253 (N_4253,N_82,N_887);
and U4254 (N_4254,N_1810,N_1606);
or U4255 (N_4255,N_2437,N_994);
nor U4256 (N_4256,N_252,N_411);
or U4257 (N_4257,N_2379,N_2208);
nor U4258 (N_4258,N_1159,N_1898);
nand U4259 (N_4259,N_2008,N_2137);
xnor U4260 (N_4260,N_1100,N_2407);
and U4261 (N_4261,N_2184,N_1284);
or U4262 (N_4262,N_1477,N_1957);
nor U4263 (N_4263,N_1087,N_1224);
or U4264 (N_4264,N_761,N_551);
nand U4265 (N_4265,N_2408,N_803);
nand U4266 (N_4266,N_585,N_400);
and U4267 (N_4267,N_1665,N_1574);
or U4268 (N_4268,N_1128,N_448);
and U4269 (N_4269,N_1154,N_656);
xor U4270 (N_4270,N_1693,N_2217);
and U4271 (N_4271,N_440,N_2173);
or U4272 (N_4272,N_1636,N_1211);
nor U4273 (N_4273,N_1823,N_1315);
or U4274 (N_4274,N_1163,N_2483);
and U4275 (N_4275,N_1104,N_1138);
nand U4276 (N_4276,N_2341,N_1122);
nand U4277 (N_4277,N_1221,N_99);
nor U4278 (N_4278,N_667,N_512);
or U4279 (N_4279,N_741,N_1020);
or U4280 (N_4280,N_2089,N_403);
nand U4281 (N_4281,N_1167,N_2450);
or U4282 (N_4282,N_1931,N_2019);
xnor U4283 (N_4283,N_1969,N_256);
nor U4284 (N_4284,N_541,N_2091);
nand U4285 (N_4285,N_526,N_747);
nor U4286 (N_4286,N_2349,N_1815);
or U4287 (N_4287,N_1927,N_857);
nand U4288 (N_4288,N_61,N_2278);
nand U4289 (N_4289,N_253,N_2267);
and U4290 (N_4290,N_1306,N_1766);
nor U4291 (N_4291,N_298,N_594);
nor U4292 (N_4292,N_1659,N_366);
xnor U4293 (N_4293,N_2440,N_709);
nand U4294 (N_4294,N_1352,N_114);
and U4295 (N_4295,N_1140,N_743);
and U4296 (N_4296,N_2339,N_890);
nor U4297 (N_4297,N_1381,N_1578);
or U4298 (N_4298,N_2150,N_895);
nor U4299 (N_4299,N_1600,N_2280);
nand U4300 (N_4300,N_486,N_268);
or U4301 (N_4301,N_1741,N_645);
nand U4302 (N_4302,N_2086,N_2324);
or U4303 (N_4303,N_0,N_747);
nand U4304 (N_4304,N_2157,N_2169);
or U4305 (N_4305,N_2098,N_965);
or U4306 (N_4306,N_1737,N_1295);
nand U4307 (N_4307,N_1985,N_2439);
nor U4308 (N_4308,N_1818,N_966);
and U4309 (N_4309,N_2224,N_180);
or U4310 (N_4310,N_2278,N_789);
or U4311 (N_4311,N_2032,N_794);
nand U4312 (N_4312,N_194,N_1837);
nor U4313 (N_4313,N_2003,N_29);
or U4314 (N_4314,N_194,N_651);
and U4315 (N_4315,N_969,N_1170);
nor U4316 (N_4316,N_1164,N_2456);
nand U4317 (N_4317,N_2435,N_1587);
nor U4318 (N_4318,N_453,N_664);
or U4319 (N_4319,N_402,N_1304);
nand U4320 (N_4320,N_1865,N_698);
nand U4321 (N_4321,N_509,N_231);
or U4322 (N_4322,N_460,N_2009);
nand U4323 (N_4323,N_342,N_400);
xor U4324 (N_4324,N_2349,N_12);
and U4325 (N_4325,N_346,N_2435);
and U4326 (N_4326,N_1040,N_1219);
or U4327 (N_4327,N_1012,N_1349);
and U4328 (N_4328,N_1815,N_2157);
and U4329 (N_4329,N_1644,N_644);
and U4330 (N_4330,N_1843,N_2375);
nand U4331 (N_4331,N_1984,N_1946);
nand U4332 (N_4332,N_917,N_1088);
nor U4333 (N_4333,N_2431,N_326);
or U4334 (N_4334,N_703,N_1309);
and U4335 (N_4335,N_789,N_2173);
nor U4336 (N_4336,N_2417,N_1684);
nor U4337 (N_4337,N_582,N_1464);
nand U4338 (N_4338,N_335,N_1299);
or U4339 (N_4339,N_2381,N_1002);
or U4340 (N_4340,N_2108,N_2232);
or U4341 (N_4341,N_122,N_765);
nor U4342 (N_4342,N_421,N_1917);
and U4343 (N_4343,N_1398,N_2436);
or U4344 (N_4344,N_274,N_2449);
nand U4345 (N_4345,N_791,N_2258);
nand U4346 (N_4346,N_1701,N_728);
xnor U4347 (N_4347,N_2142,N_854);
or U4348 (N_4348,N_2316,N_1102);
or U4349 (N_4349,N_2166,N_2137);
and U4350 (N_4350,N_1499,N_1211);
and U4351 (N_4351,N_1209,N_1431);
nor U4352 (N_4352,N_2430,N_1520);
and U4353 (N_4353,N_1359,N_729);
or U4354 (N_4354,N_2296,N_26);
nor U4355 (N_4355,N_208,N_1776);
or U4356 (N_4356,N_2188,N_1913);
and U4357 (N_4357,N_1401,N_1542);
nand U4358 (N_4358,N_117,N_150);
xor U4359 (N_4359,N_724,N_173);
nand U4360 (N_4360,N_267,N_1865);
and U4361 (N_4361,N_294,N_811);
nor U4362 (N_4362,N_2351,N_638);
nor U4363 (N_4363,N_2215,N_1464);
nor U4364 (N_4364,N_226,N_143);
or U4365 (N_4365,N_477,N_622);
and U4366 (N_4366,N_917,N_1844);
or U4367 (N_4367,N_1060,N_200);
and U4368 (N_4368,N_652,N_12);
and U4369 (N_4369,N_497,N_1682);
and U4370 (N_4370,N_2232,N_243);
nand U4371 (N_4371,N_8,N_1341);
and U4372 (N_4372,N_386,N_1173);
and U4373 (N_4373,N_1295,N_949);
nor U4374 (N_4374,N_34,N_2111);
xor U4375 (N_4375,N_435,N_965);
nand U4376 (N_4376,N_2404,N_1221);
or U4377 (N_4377,N_2358,N_536);
nor U4378 (N_4378,N_1896,N_1634);
and U4379 (N_4379,N_1756,N_1406);
nor U4380 (N_4380,N_2424,N_1446);
nand U4381 (N_4381,N_2330,N_591);
or U4382 (N_4382,N_1947,N_399);
and U4383 (N_4383,N_749,N_185);
nor U4384 (N_4384,N_742,N_2184);
nand U4385 (N_4385,N_2494,N_1859);
and U4386 (N_4386,N_1597,N_967);
or U4387 (N_4387,N_1415,N_1419);
nor U4388 (N_4388,N_233,N_1503);
nor U4389 (N_4389,N_547,N_1314);
nor U4390 (N_4390,N_353,N_416);
nand U4391 (N_4391,N_1471,N_2049);
or U4392 (N_4392,N_1264,N_1400);
nand U4393 (N_4393,N_324,N_1341);
nand U4394 (N_4394,N_2177,N_1262);
nor U4395 (N_4395,N_624,N_1851);
xnor U4396 (N_4396,N_993,N_2268);
nor U4397 (N_4397,N_1333,N_1356);
and U4398 (N_4398,N_2064,N_1991);
and U4399 (N_4399,N_1381,N_2049);
or U4400 (N_4400,N_1626,N_2026);
nor U4401 (N_4401,N_469,N_325);
nand U4402 (N_4402,N_1430,N_2134);
nand U4403 (N_4403,N_539,N_1569);
and U4404 (N_4404,N_2300,N_1298);
and U4405 (N_4405,N_1788,N_2259);
or U4406 (N_4406,N_370,N_1936);
and U4407 (N_4407,N_1765,N_892);
nand U4408 (N_4408,N_703,N_416);
and U4409 (N_4409,N_234,N_1209);
nor U4410 (N_4410,N_2219,N_8);
or U4411 (N_4411,N_2351,N_1052);
or U4412 (N_4412,N_912,N_2283);
xor U4413 (N_4413,N_1530,N_415);
and U4414 (N_4414,N_2263,N_1322);
nand U4415 (N_4415,N_1287,N_1886);
nand U4416 (N_4416,N_1922,N_2473);
nor U4417 (N_4417,N_123,N_603);
xor U4418 (N_4418,N_621,N_1734);
nand U4419 (N_4419,N_916,N_735);
nand U4420 (N_4420,N_988,N_2212);
nand U4421 (N_4421,N_57,N_1444);
and U4422 (N_4422,N_1033,N_585);
and U4423 (N_4423,N_1215,N_2034);
or U4424 (N_4424,N_40,N_1769);
nor U4425 (N_4425,N_1296,N_860);
and U4426 (N_4426,N_2194,N_584);
nand U4427 (N_4427,N_1535,N_93);
and U4428 (N_4428,N_1424,N_152);
nor U4429 (N_4429,N_988,N_213);
or U4430 (N_4430,N_17,N_1802);
or U4431 (N_4431,N_2460,N_360);
or U4432 (N_4432,N_2418,N_186);
or U4433 (N_4433,N_180,N_2445);
nand U4434 (N_4434,N_1267,N_967);
or U4435 (N_4435,N_600,N_1050);
nor U4436 (N_4436,N_2439,N_836);
or U4437 (N_4437,N_1293,N_789);
nor U4438 (N_4438,N_1899,N_905);
nand U4439 (N_4439,N_887,N_1669);
nor U4440 (N_4440,N_2389,N_2247);
nor U4441 (N_4441,N_1293,N_1883);
or U4442 (N_4442,N_1104,N_877);
xor U4443 (N_4443,N_671,N_1850);
nor U4444 (N_4444,N_1985,N_2223);
nand U4445 (N_4445,N_880,N_2260);
nand U4446 (N_4446,N_23,N_880);
nand U4447 (N_4447,N_1934,N_99);
nor U4448 (N_4448,N_1367,N_1201);
xor U4449 (N_4449,N_190,N_1528);
or U4450 (N_4450,N_1274,N_885);
and U4451 (N_4451,N_1007,N_181);
nor U4452 (N_4452,N_2492,N_2458);
or U4453 (N_4453,N_2459,N_307);
and U4454 (N_4454,N_1345,N_720);
nand U4455 (N_4455,N_1698,N_1922);
nor U4456 (N_4456,N_1523,N_1506);
or U4457 (N_4457,N_1967,N_1137);
and U4458 (N_4458,N_1215,N_2167);
and U4459 (N_4459,N_1650,N_127);
nor U4460 (N_4460,N_961,N_1062);
and U4461 (N_4461,N_322,N_1796);
nand U4462 (N_4462,N_1832,N_566);
nor U4463 (N_4463,N_1637,N_903);
and U4464 (N_4464,N_1023,N_604);
and U4465 (N_4465,N_863,N_2184);
nand U4466 (N_4466,N_272,N_2361);
and U4467 (N_4467,N_79,N_1019);
and U4468 (N_4468,N_94,N_1373);
xnor U4469 (N_4469,N_1600,N_666);
or U4470 (N_4470,N_196,N_2392);
nor U4471 (N_4471,N_1923,N_2468);
nand U4472 (N_4472,N_1904,N_108);
or U4473 (N_4473,N_1176,N_1798);
nand U4474 (N_4474,N_1227,N_1552);
or U4475 (N_4475,N_2015,N_2308);
or U4476 (N_4476,N_901,N_1749);
and U4477 (N_4477,N_1459,N_348);
nand U4478 (N_4478,N_1408,N_972);
and U4479 (N_4479,N_165,N_63);
nand U4480 (N_4480,N_299,N_2364);
or U4481 (N_4481,N_1936,N_1517);
nand U4482 (N_4482,N_2141,N_1970);
nand U4483 (N_4483,N_1829,N_1639);
and U4484 (N_4484,N_2027,N_871);
nand U4485 (N_4485,N_813,N_1021);
nand U4486 (N_4486,N_1971,N_992);
and U4487 (N_4487,N_1282,N_1312);
or U4488 (N_4488,N_962,N_2214);
and U4489 (N_4489,N_131,N_731);
and U4490 (N_4490,N_2094,N_1232);
nand U4491 (N_4491,N_815,N_2074);
or U4492 (N_4492,N_353,N_1990);
or U4493 (N_4493,N_2310,N_694);
and U4494 (N_4494,N_2448,N_1654);
nor U4495 (N_4495,N_1064,N_466);
nor U4496 (N_4496,N_1577,N_77);
nand U4497 (N_4497,N_783,N_1507);
xor U4498 (N_4498,N_1577,N_1065);
and U4499 (N_4499,N_2259,N_590);
nor U4500 (N_4500,N_648,N_1293);
nand U4501 (N_4501,N_816,N_1996);
and U4502 (N_4502,N_619,N_2447);
nand U4503 (N_4503,N_628,N_990);
nor U4504 (N_4504,N_8,N_950);
nor U4505 (N_4505,N_722,N_1515);
nor U4506 (N_4506,N_2153,N_82);
or U4507 (N_4507,N_955,N_163);
nand U4508 (N_4508,N_1185,N_2323);
nand U4509 (N_4509,N_1517,N_1044);
and U4510 (N_4510,N_299,N_1003);
nor U4511 (N_4511,N_1131,N_1741);
or U4512 (N_4512,N_2278,N_554);
and U4513 (N_4513,N_1352,N_2100);
or U4514 (N_4514,N_836,N_1506);
nand U4515 (N_4515,N_793,N_460);
and U4516 (N_4516,N_678,N_160);
or U4517 (N_4517,N_1718,N_1895);
nand U4518 (N_4518,N_1483,N_138);
or U4519 (N_4519,N_897,N_1916);
or U4520 (N_4520,N_1339,N_514);
nand U4521 (N_4521,N_875,N_1141);
nor U4522 (N_4522,N_1865,N_473);
nand U4523 (N_4523,N_2256,N_416);
nand U4524 (N_4524,N_1316,N_2251);
and U4525 (N_4525,N_1589,N_1293);
or U4526 (N_4526,N_1436,N_141);
and U4527 (N_4527,N_1444,N_1159);
nor U4528 (N_4528,N_1782,N_2298);
and U4529 (N_4529,N_950,N_158);
and U4530 (N_4530,N_698,N_1238);
nor U4531 (N_4531,N_1138,N_345);
and U4532 (N_4532,N_166,N_263);
or U4533 (N_4533,N_2497,N_169);
and U4534 (N_4534,N_1794,N_434);
and U4535 (N_4535,N_2147,N_949);
nand U4536 (N_4536,N_546,N_1471);
nand U4537 (N_4537,N_797,N_1328);
xnor U4538 (N_4538,N_1716,N_1524);
and U4539 (N_4539,N_2360,N_2094);
nand U4540 (N_4540,N_300,N_635);
and U4541 (N_4541,N_1261,N_2277);
nand U4542 (N_4542,N_496,N_2035);
nand U4543 (N_4543,N_2195,N_2350);
or U4544 (N_4544,N_1749,N_1483);
or U4545 (N_4545,N_791,N_5);
nor U4546 (N_4546,N_106,N_1057);
and U4547 (N_4547,N_822,N_1813);
nand U4548 (N_4548,N_1695,N_276);
nand U4549 (N_4549,N_109,N_2485);
nand U4550 (N_4550,N_1017,N_2064);
or U4551 (N_4551,N_1726,N_2028);
nor U4552 (N_4552,N_1083,N_467);
and U4553 (N_4553,N_493,N_2008);
or U4554 (N_4554,N_1688,N_302);
or U4555 (N_4555,N_1318,N_2105);
nand U4556 (N_4556,N_1957,N_1634);
nand U4557 (N_4557,N_2346,N_626);
and U4558 (N_4558,N_307,N_741);
and U4559 (N_4559,N_2270,N_2177);
nor U4560 (N_4560,N_373,N_736);
nand U4561 (N_4561,N_2117,N_1973);
nand U4562 (N_4562,N_1005,N_2115);
nor U4563 (N_4563,N_943,N_1715);
or U4564 (N_4564,N_1872,N_1405);
xnor U4565 (N_4565,N_568,N_1365);
nor U4566 (N_4566,N_1649,N_818);
nand U4567 (N_4567,N_359,N_1313);
nor U4568 (N_4568,N_1761,N_2076);
or U4569 (N_4569,N_2041,N_1839);
and U4570 (N_4570,N_25,N_1012);
nor U4571 (N_4571,N_1553,N_2127);
or U4572 (N_4572,N_1477,N_1473);
xnor U4573 (N_4573,N_2462,N_1178);
or U4574 (N_4574,N_1836,N_238);
nand U4575 (N_4575,N_1031,N_121);
nor U4576 (N_4576,N_1508,N_1952);
and U4577 (N_4577,N_277,N_476);
nor U4578 (N_4578,N_1736,N_2484);
or U4579 (N_4579,N_4,N_2424);
nand U4580 (N_4580,N_2347,N_1228);
nor U4581 (N_4581,N_770,N_1015);
and U4582 (N_4582,N_1139,N_1540);
nor U4583 (N_4583,N_18,N_1497);
and U4584 (N_4584,N_2360,N_2042);
nand U4585 (N_4585,N_939,N_1624);
and U4586 (N_4586,N_996,N_2359);
or U4587 (N_4587,N_784,N_1297);
nand U4588 (N_4588,N_2468,N_476);
or U4589 (N_4589,N_298,N_1463);
nand U4590 (N_4590,N_1191,N_1983);
or U4591 (N_4591,N_222,N_1676);
nand U4592 (N_4592,N_2167,N_1899);
or U4593 (N_4593,N_1558,N_2102);
or U4594 (N_4594,N_394,N_1147);
nand U4595 (N_4595,N_1182,N_748);
or U4596 (N_4596,N_1902,N_2335);
and U4597 (N_4597,N_1348,N_1666);
or U4598 (N_4598,N_1776,N_122);
nand U4599 (N_4599,N_2492,N_1704);
or U4600 (N_4600,N_729,N_711);
nand U4601 (N_4601,N_2384,N_468);
and U4602 (N_4602,N_1495,N_1994);
or U4603 (N_4603,N_630,N_1030);
nand U4604 (N_4604,N_1322,N_1472);
nor U4605 (N_4605,N_749,N_967);
nor U4606 (N_4606,N_688,N_2411);
and U4607 (N_4607,N_741,N_2206);
and U4608 (N_4608,N_1353,N_334);
nor U4609 (N_4609,N_141,N_2056);
nand U4610 (N_4610,N_2203,N_1764);
nor U4611 (N_4611,N_446,N_2156);
nor U4612 (N_4612,N_2112,N_2220);
nand U4613 (N_4613,N_1603,N_2294);
or U4614 (N_4614,N_762,N_1957);
and U4615 (N_4615,N_203,N_835);
or U4616 (N_4616,N_139,N_1862);
nor U4617 (N_4617,N_440,N_179);
nand U4618 (N_4618,N_63,N_1488);
or U4619 (N_4619,N_832,N_770);
or U4620 (N_4620,N_1742,N_785);
and U4621 (N_4621,N_2389,N_1752);
nand U4622 (N_4622,N_1196,N_1760);
nor U4623 (N_4623,N_956,N_885);
or U4624 (N_4624,N_1304,N_708);
or U4625 (N_4625,N_2339,N_1396);
nand U4626 (N_4626,N_442,N_306);
or U4627 (N_4627,N_2209,N_2387);
and U4628 (N_4628,N_2389,N_912);
nand U4629 (N_4629,N_2197,N_815);
and U4630 (N_4630,N_1607,N_1832);
nand U4631 (N_4631,N_1999,N_1964);
and U4632 (N_4632,N_2157,N_2056);
nor U4633 (N_4633,N_2204,N_1174);
or U4634 (N_4634,N_1063,N_617);
and U4635 (N_4635,N_893,N_1337);
nor U4636 (N_4636,N_2149,N_2224);
nor U4637 (N_4637,N_1569,N_1363);
or U4638 (N_4638,N_2051,N_2261);
nor U4639 (N_4639,N_2346,N_2248);
nor U4640 (N_4640,N_2011,N_967);
and U4641 (N_4641,N_1102,N_908);
or U4642 (N_4642,N_1515,N_447);
and U4643 (N_4643,N_2150,N_2175);
nand U4644 (N_4644,N_2177,N_2268);
nor U4645 (N_4645,N_2289,N_430);
or U4646 (N_4646,N_777,N_569);
or U4647 (N_4647,N_1575,N_2384);
nor U4648 (N_4648,N_2124,N_1190);
or U4649 (N_4649,N_522,N_997);
or U4650 (N_4650,N_1006,N_797);
and U4651 (N_4651,N_286,N_860);
and U4652 (N_4652,N_954,N_1223);
or U4653 (N_4653,N_832,N_835);
nor U4654 (N_4654,N_2436,N_869);
nand U4655 (N_4655,N_1649,N_27);
or U4656 (N_4656,N_2363,N_572);
nor U4657 (N_4657,N_64,N_1872);
and U4658 (N_4658,N_1090,N_1118);
or U4659 (N_4659,N_647,N_552);
nand U4660 (N_4660,N_1294,N_1503);
nor U4661 (N_4661,N_1998,N_1993);
nor U4662 (N_4662,N_1005,N_939);
nand U4663 (N_4663,N_2197,N_215);
or U4664 (N_4664,N_2223,N_1619);
nor U4665 (N_4665,N_243,N_1603);
nor U4666 (N_4666,N_1052,N_634);
or U4667 (N_4667,N_981,N_2110);
nor U4668 (N_4668,N_2159,N_713);
or U4669 (N_4669,N_1129,N_612);
nor U4670 (N_4670,N_730,N_2435);
and U4671 (N_4671,N_1867,N_1510);
nor U4672 (N_4672,N_66,N_939);
or U4673 (N_4673,N_1689,N_1481);
nor U4674 (N_4674,N_931,N_1953);
and U4675 (N_4675,N_762,N_1899);
nand U4676 (N_4676,N_1549,N_908);
nor U4677 (N_4677,N_1471,N_241);
nor U4678 (N_4678,N_1699,N_1240);
nor U4679 (N_4679,N_321,N_743);
nand U4680 (N_4680,N_1194,N_2058);
and U4681 (N_4681,N_1548,N_1479);
nor U4682 (N_4682,N_149,N_2107);
nand U4683 (N_4683,N_819,N_1315);
or U4684 (N_4684,N_2443,N_816);
and U4685 (N_4685,N_1594,N_1259);
nor U4686 (N_4686,N_528,N_1526);
and U4687 (N_4687,N_1923,N_1152);
nor U4688 (N_4688,N_1424,N_1947);
nand U4689 (N_4689,N_418,N_313);
nor U4690 (N_4690,N_2271,N_600);
or U4691 (N_4691,N_461,N_1222);
nor U4692 (N_4692,N_1178,N_1633);
and U4693 (N_4693,N_641,N_1043);
and U4694 (N_4694,N_994,N_389);
and U4695 (N_4695,N_624,N_2019);
and U4696 (N_4696,N_405,N_1198);
nor U4697 (N_4697,N_2192,N_1301);
and U4698 (N_4698,N_1674,N_1861);
and U4699 (N_4699,N_1922,N_1529);
or U4700 (N_4700,N_1888,N_125);
nor U4701 (N_4701,N_334,N_741);
nand U4702 (N_4702,N_1601,N_1076);
nor U4703 (N_4703,N_2356,N_2064);
and U4704 (N_4704,N_1596,N_1590);
nor U4705 (N_4705,N_1590,N_760);
and U4706 (N_4706,N_58,N_1818);
and U4707 (N_4707,N_1854,N_504);
nand U4708 (N_4708,N_465,N_1836);
nor U4709 (N_4709,N_1553,N_1747);
nor U4710 (N_4710,N_2483,N_2354);
nor U4711 (N_4711,N_1966,N_260);
nor U4712 (N_4712,N_1739,N_1636);
nor U4713 (N_4713,N_1753,N_907);
nor U4714 (N_4714,N_1758,N_663);
or U4715 (N_4715,N_1850,N_892);
nand U4716 (N_4716,N_1861,N_967);
nor U4717 (N_4717,N_1974,N_2440);
nor U4718 (N_4718,N_2115,N_1354);
nand U4719 (N_4719,N_120,N_1299);
nor U4720 (N_4720,N_2033,N_1274);
nor U4721 (N_4721,N_613,N_2347);
or U4722 (N_4722,N_1113,N_1997);
nor U4723 (N_4723,N_1448,N_933);
nor U4724 (N_4724,N_300,N_41);
or U4725 (N_4725,N_765,N_1695);
nor U4726 (N_4726,N_1852,N_1644);
nand U4727 (N_4727,N_2246,N_2231);
nand U4728 (N_4728,N_658,N_2299);
or U4729 (N_4729,N_2093,N_2166);
or U4730 (N_4730,N_2281,N_1907);
nor U4731 (N_4731,N_967,N_1664);
or U4732 (N_4732,N_1541,N_745);
xnor U4733 (N_4733,N_1625,N_1410);
and U4734 (N_4734,N_1666,N_30);
or U4735 (N_4735,N_1190,N_1901);
nor U4736 (N_4736,N_102,N_1800);
nor U4737 (N_4737,N_899,N_1106);
nor U4738 (N_4738,N_491,N_676);
nand U4739 (N_4739,N_512,N_1037);
or U4740 (N_4740,N_467,N_900);
nand U4741 (N_4741,N_1307,N_2296);
or U4742 (N_4742,N_2428,N_2380);
nand U4743 (N_4743,N_2207,N_1397);
and U4744 (N_4744,N_1239,N_596);
and U4745 (N_4745,N_265,N_707);
nor U4746 (N_4746,N_970,N_2444);
nand U4747 (N_4747,N_1678,N_1277);
and U4748 (N_4748,N_1621,N_332);
nor U4749 (N_4749,N_2089,N_407);
and U4750 (N_4750,N_1965,N_1114);
and U4751 (N_4751,N_362,N_382);
and U4752 (N_4752,N_1640,N_1260);
or U4753 (N_4753,N_1899,N_1255);
nand U4754 (N_4754,N_331,N_2429);
nand U4755 (N_4755,N_900,N_1647);
nand U4756 (N_4756,N_1900,N_1873);
or U4757 (N_4757,N_1705,N_1429);
nand U4758 (N_4758,N_1337,N_1076);
and U4759 (N_4759,N_1845,N_1254);
nor U4760 (N_4760,N_1661,N_1958);
or U4761 (N_4761,N_586,N_50);
nand U4762 (N_4762,N_1678,N_1410);
and U4763 (N_4763,N_2099,N_2213);
nor U4764 (N_4764,N_324,N_2249);
and U4765 (N_4765,N_283,N_2371);
or U4766 (N_4766,N_2201,N_1008);
xnor U4767 (N_4767,N_1371,N_572);
nor U4768 (N_4768,N_2495,N_28);
and U4769 (N_4769,N_1562,N_810);
nor U4770 (N_4770,N_1718,N_62);
xor U4771 (N_4771,N_1492,N_615);
nor U4772 (N_4772,N_1215,N_298);
or U4773 (N_4773,N_1403,N_646);
nand U4774 (N_4774,N_666,N_2059);
or U4775 (N_4775,N_1962,N_2249);
nand U4776 (N_4776,N_2154,N_2267);
and U4777 (N_4777,N_2269,N_1833);
nor U4778 (N_4778,N_1162,N_1057);
nand U4779 (N_4779,N_2054,N_1728);
and U4780 (N_4780,N_1296,N_572);
or U4781 (N_4781,N_1597,N_278);
or U4782 (N_4782,N_919,N_1791);
nand U4783 (N_4783,N_1033,N_884);
or U4784 (N_4784,N_712,N_1050);
nand U4785 (N_4785,N_68,N_1748);
nand U4786 (N_4786,N_1588,N_1317);
or U4787 (N_4787,N_1184,N_2464);
nor U4788 (N_4788,N_2145,N_579);
nand U4789 (N_4789,N_1024,N_1510);
nor U4790 (N_4790,N_2301,N_2069);
nor U4791 (N_4791,N_2439,N_1073);
nor U4792 (N_4792,N_346,N_1723);
and U4793 (N_4793,N_1081,N_585);
nor U4794 (N_4794,N_122,N_2479);
nor U4795 (N_4795,N_291,N_683);
nor U4796 (N_4796,N_1648,N_2351);
nor U4797 (N_4797,N_1243,N_2128);
nor U4798 (N_4798,N_313,N_1807);
nor U4799 (N_4799,N_596,N_1134);
nor U4800 (N_4800,N_2242,N_2404);
and U4801 (N_4801,N_38,N_127);
nor U4802 (N_4802,N_1824,N_806);
nand U4803 (N_4803,N_109,N_2478);
nand U4804 (N_4804,N_722,N_801);
nor U4805 (N_4805,N_1346,N_2423);
and U4806 (N_4806,N_996,N_1571);
nand U4807 (N_4807,N_1413,N_1470);
and U4808 (N_4808,N_1611,N_2350);
and U4809 (N_4809,N_2130,N_203);
nand U4810 (N_4810,N_73,N_1151);
nor U4811 (N_4811,N_2474,N_1057);
xnor U4812 (N_4812,N_2184,N_1933);
nand U4813 (N_4813,N_1463,N_1190);
or U4814 (N_4814,N_1008,N_330);
nor U4815 (N_4815,N_1334,N_2052);
nand U4816 (N_4816,N_1733,N_1318);
nand U4817 (N_4817,N_1854,N_1876);
nand U4818 (N_4818,N_64,N_1794);
nor U4819 (N_4819,N_227,N_2013);
nor U4820 (N_4820,N_808,N_1628);
nand U4821 (N_4821,N_1640,N_294);
nand U4822 (N_4822,N_2441,N_2440);
or U4823 (N_4823,N_1498,N_210);
or U4824 (N_4824,N_1131,N_937);
and U4825 (N_4825,N_1758,N_933);
or U4826 (N_4826,N_1418,N_1209);
nand U4827 (N_4827,N_1062,N_2364);
and U4828 (N_4828,N_2090,N_800);
nor U4829 (N_4829,N_1602,N_1416);
or U4830 (N_4830,N_1036,N_1592);
nor U4831 (N_4831,N_1036,N_458);
and U4832 (N_4832,N_1142,N_2434);
and U4833 (N_4833,N_373,N_583);
nand U4834 (N_4834,N_2125,N_873);
nand U4835 (N_4835,N_2180,N_1537);
or U4836 (N_4836,N_1188,N_1954);
and U4837 (N_4837,N_1911,N_2000);
nand U4838 (N_4838,N_1451,N_1820);
and U4839 (N_4839,N_594,N_717);
and U4840 (N_4840,N_478,N_2385);
nor U4841 (N_4841,N_1633,N_2279);
and U4842 (N_4842,N_608,N_641);
or U4843 (N_4843,N_31,N_1173);
or U4844 (N_4844,N_896,N_174);
nand U4845 (N_4845,N_2061,N_1143);
nand U4846 (N_4846,N_1880,N_844);
nor U4847 (N_4847,N_384,N_160);
and U4848 (N_4848,N_970,N_975);
and U4849 (N_4849,N_689,N_567);
nor U4850 (N_4850,N_1888,N_1345);
nand U4851 (N_4851,N_1364,N_15);
and U4852 (N_4852,N_1499,N_435);
nand U4853 (N_4853,N_1693,N_416);
and U4854 (N_4854,N_1858,N_511);
nand U4855 (N_4855,N_803,N_2466);
or U4856 (N_4856,N_1568,N_446);
nand U4857 (N_4857,N_555,N_1062);
nand U4858 (N_4858,N_1884,N_1256);
nand U4859 (N_4859,N_40,N_764);
nand U4860 (N_4860,N_1582,N_2483);
nor U4861 (N_4861,N_653,N_202);
xnor U4862 (N_4862,N_275,N_436);
nand U4863 (N_4863,N_85,N_268);
or U4864 (N_4864,N_1058,N_1637);
or U4865 (N_4865,N_1655,N_894);
and U4866 (N_4866,N_1944,N_263);
and U4867 (N_4867,N_2363,N_2123);
nand U4868 (N_4868,N_975,N_790);
and U4869 (N_4869,N_2415,N_130);
and U4870 (N_4870,N_703,N_134);
nor U4871 (N_4871,N_1542,N_1592);
and U4872 (N_4872,N_1764,N_2032);
nor U4873 (N_4873,N_1199,N_1961);
nand U4874 (N_4874,N_1703,N_1658);
nor U4875 (N_4875,N_716,N_619);
nand U4876 (N_4876,N_2115,N_1849);
nand U4877 (N_4877,N_531,N_2095);
or U4878 (N_4878,N_231,N_605);
nor U4879 (N_4879,N_86,N_188);
nand U4880 (N_4880,N_1224,N_753);
or U4881 (N_4881,N_699,N_2406);
or U4882 (N_4882,N_1700,N_1807);
and U4883 (N_4883,N_2166,N_1214);
or U4884 (N_4884,N_1783,N_801);
nor U4885 (N_4885,N_832,N_1413);
nor U4886 (N_4886,N_1209,N_1857);
and U4887 (N_4887,N_1441,N_1530);
and U4888 (N_4888,N_1130,N_76);
and U4889 (N_4889,N_680,N_1624);
nand U4890 (N_4890,N_2244,N_103);
or U4891 (N_4891,N_2456,N_1129);
and U4892 (N_4892,N_1971,N_2123);
and U4893 (N_4893,N_2097,N_2481);
and U4894 (N_4894,N_2234,N_1035);
and U4895 (N_4895,N_2043,N_383);
and U4896 (N_4896,N_1427,N_893);
nor U4897 (N_4897,N_1123,N_1268);
nor U4898 (N_4898,N_1074,N_2479);
or U4899 (N_4899,N_2169,N_1500);
nor U4900 (N_4900,N_847,N_504);
or U4901 (N_4901,N_644,N_1125);
or U4902 (N_4902,N_1479,N_158);
and U4903 (N_4903,N_2225,N_2306);
nand U4904 (N_4904,N_372,N_714);
nor U4905 (N_4905,N_385,N_528);
nor U4906 (N_4906,N_1252,N_2128);
and U4907 (N_4907,N_908,N_2239);
and U4908 (N_4908,N_191,N_3);
nor U4909 (N_4909,N_1878,N_1946);
or U4910 (N_4910,N_1866,N_832);
or U4911 (N_4911,N_2425,N_2206);
nor U4912 (N_4912,N_64,N_1446);
or U4913 (N_4913,N_2153,N_2063);
and U4914 (N_4914,N_1525,N_422);
nand U4915 (N_4915,N_2011,N_407);
and U4916 (N_4916,N_2128,N_1739);
or U4917 (N_4917,N_1071,N_1237);
and U4918 (N_4918,N_904,N_1731);
nor U4919 (N_4919,N_1380,N_1149);
and U4920 (N_4920,N_233,N_163);
nor U4921 (N_4921,N_681,N_2087);
nor U4922 (N_4922,N_636,N_766);
nor U4923 (N_4923,N_1681,N_1571);
and U4924 (N_4924,N_577,N_187);
nand U4925 (N_4925,N_587,N_704);
nand U4926 (N_4926,N_2225,N_2017);
or U4927 (N_4927,N_1584,N_2116);
xor U4928 (N_4928,N_125,N_291);
nor U4929 (N_4929,N_2152,N_148);
and U4930 (N_4930,N_1497,N_645);
nand U4931 (N_4931,N_2427,N_1297);
or U4932 (N_4932,N_459,N_1201);
and U4933 (N_4933,N_1767,N_873);
nand U4934 (N_4934,N_991,N_427);
nor U4935 (N_4935,N_1356,N_1283);
nand U4936 (N_4936,N_1316,N_2231);
or U4937 (N_4937,N_1037,N_2358);
and U4938 (N_4938,N_1997,N_2381);
and U4939 (N_4939,N_626,N_2227);
nand U4940 (N_4940,N_2422,N_1922);
or U4941 (N_4941,N_1200,N_401);
or U4942 (N_4942,N_1957,N_2259);
nand U4943 (N_4943,N_91,N_2135);
and U4944 (N_4944,N_1542,N_246);
and U4945 (N_4945,N_49,N_669);
nand U4946 (N_4946,N_1564,N_1227);
or U4947 (N_4947,N_1317,N_1540);
nor U4948 (N_4948,N_2362,N_492);
or U4949 (N_4949,N_1552,N_480);
nand U4950 (N_4950,N_272,N_1163);
nand U4951 (N_4951,N_2486,N_665);
nand U4952 (N_4952,N_1812,N_2309);
and U4953 (N_4953,N_1755,N_2108);
nand U4954 (N_4954,N_583,N_974);
and U4955 (N_4955,N_1414,N_1283);
xnor U4956 (N_4956,N_1910,N_297);
xor U4957 (N_4957,N_1334,N_626);
nor U4958 (N_4958,N_2039,N_53);
or U4959 (N_4959,N_1663,N_2049);
and U4960 (N_4960,N_1200,N_479);
and U4961 (N_4961,N_1856,N_816);
or U4962 (N_4962,N_1036,N_2346);
nor U4963 (N_4963,N_1344,N_178);
and U4964 (N_4964,N_85,N_2036);
nor U4965 (N_4965,N_1003,N_1894);
or U4966 (N_4966,N_1881,N_1395);
nor U4967 (N_4967,N_373,N_342);
and U4968 (N_4968,N_1095,N_2408);
nor U4969 (N_4969,N_732,N_2410);
and U4970 (N_4970,N_952,N_2129);
nand U4971 (N_4971,N_1573,N_1106);
nand U4972 (N_4972,N_1528,N_924);
nand U4973 (N_4973,N_1306,N_2295);
nand U4974 (N_4974,N_96,N_1990);
nand U4975 (N_4975,N_2024,N_886);
nor U4976 (N_4976,N_2032,N_80);
and U4977 (N_4977,N_178,N_2196);
and U4978 (N_4978,N_1497,N_659);
and U4979 (N_4979,N_939,N_2248);
and U4980 (N_4980,N_2358,N_1690);
nor U4981 (N_4981,N_1667,N_1236);
nand U4982 (N_4982,N_1200,N_31);
nor U4983 (N_4983,N_364,N_1275);
nor U4984 (N_4984,N_1151,N_185);
or U4985 (N_4985,N_1061,N_1729);
nand U4986 (N_4986,N_1732,N_1877);
or U4987 (N_4987,N_502,N_1186);
nand U4988 (N_4988,N_606,N_2242);
or U4989 (N_4989,N_1799,N_170);
nor U4990 (N_4990,N_97,N_1857);
nor U4991 (N_4991,N_631,N_2173);
nor U4992 (N_4992,N_1586,N_250);
and U4993 (N_4993,N_308,N_2043);
and U4994 (N_4994,N_2224,N_1520);
nor U4995 (N_4995,N_1461,N_1399);
or U4996 (N_4996,N_169,N_2260);
and U4997 (N_4997,N_362,N_2373);
xor U4998 (N_4998,N_1664,N_2017);
and U4999 (N_4999,N_1773,N_668);
or U5000 (N_5000,N_2810,N_3799);
or U5001 (N_5001,N_4138,N_3696);
nand U5002 (N_5002,N_3135,N_4588);
and U5003 (N_5003,N_4617,N_3435);
and U5004 (N_5004,N_4486,N_4529);
and U5005 (N_5005,N_2767,N_3713);
or U5006 (N_5006,N_3840,N_3862);
and U5007 (N_5007,N_4370,N_2728);
nand U5008 (N_5008,N_2758,N_2833);
or U5009 (N_5009,N_2535,N_4911);
nor U5010 (N_5010,N_2698,N_3918);
and U5011 (N_5011,N_4531,N_3309);
nand U5012 (N_5012,N_3284,N_4608);
and U5013 (N_5013,N_2913,N_3186);
nand U5014 (N_5014,N_3084,N_3831);
and U5015 (N_5015,N_3397,N_4979);
nor U5016 (N_5016,N_4291,N_3410);
nand U5017 (N_5017,N_3211,N_3905);
nor U5018 (N_5018,N_3063,N_3562);
nand U5019 (N_5019,N_2583,N_3537);
nor U5020 (N_5020,N_3990,N_2511);
nor U5021 (N_5021,N_4191,N_3520);
nor U5022 (N_5022,N_4441,N_2628);
and U5023 (N_5023,N_3471,N_4935);
nand U5024 (N_5024,N_3803,N_2696);
or U5025 (N_5025,N_3867,N_3480);
or U5026 (N_5026,N_3173,N_2902);
or U5027 (N_5027,N_3658,N_4671);
or U5028 (N_5028,N_4254,N_3829);
and U5029 (N_5029,N_4577,N_3743);
nand U5030 (N_5030,N_3947,N_4073);
nor U5031 (N_5031,N_4903,N_4110);
xor U5032 (N_5032,N_3639,N_2757);
or U5033 (N_5033,N_4941,N_4201);
nor U5034 (N_5034,N_4996,N_3275);
and U5035 (N_5035,N_3155,N_3832);
nand U5036 (N_5036,N_4691,N_4228);
nand U5037 (N_5037,N_2620,N_4366);
or U5038 (N_5038,N_3444,N_4490);
nor U5039 (N_5039,N_3857,N_3041);
nand U5040 (N_5040,N_3351,N_3834);
nand U5041 (N_5041,N_3254,N_2800);
nor U5042 (N_5042,N_4263,N_2789);
and U5043 (N_5043,N_3280,N_3675);
and U5044 (N_5044,N_4783,N_2540);
nand U5045 (N_5045,N_3133,N_4510);
nor U5046 (N_5046,N_4333,N_4025);
nand U5047 (N_5047,N_3912,N_2675);
and U5048 (N_5048,N_3736,N_4233);
nand U5049 (N_5049,N_4837,N_2704);
xnor U5050 (N_5050,N_3023,N_4625);
nand U5051 (N_5051,N_4086,N_4369);
nand U5052 (N_5052,N_2639,N_4285);
nand U5053 (N_5053,N_3367,N_2822);
nand U5054 (N_5054,N_3965,N_2917);
nand U5055 (N_5055,N_3866,N_4148);
and U5056 (N_5056,N_4600,N_2992);
and U5057 (N_5057,N_3755,N_4683);
or U5058 (N_5058,N_4178,N_3113);
nand U5059 (N_5059,N_4975,N_4619);
and U5060 (N_5060,N_3466,N_3092);
nor U5061 (N_5061,N_3493,N_2731);
nor U5062 (N_5062,N_3190,N_3760);
nor U5063 (N_5063,N_4117,N_4288);
or U5064 (N_5064,N_2989,N_3256);
or U5065 (N_5065,N_3595,N_3338);
and U5066 (N_5066,N_3602,N_4232);
nand U5067 (N_5067,N_2910,N_3777);
nor U5068 (N_5068,N_2874,N_3532);
and U5069 (N_5069,N_4072,N_3085);
and U5070 (N_5070,N_2997,N_4825);
nand U5071 (N_5071,N_4978,N_4303);
or U5072 (N_5072,N_4259,N_3228);
nand U5073 (N_5073,N_3530,N_4475);
and U5074 (N_5074,N_2750,N_3315);
and U5075 (N_5075,N_2570,N_2574);
and U5076 (N_5076,N_4289,N_4764);
xnor U5077 (N_5077,N_4275,N_4000);
or U5078 (N_5078,N_2705,N_4169);
and U5079 (N_5079,N_3408,N_3292);
nor U5080 (N_5080,N_3141,N_3664);
nand U5081 (N_5081,N_4828,N_4896);
nor U5082 (N_5082,N_4419,N_3618);
or U5083 (N_5083,N_3222,N_4244);
nor U5084 (N_5084,N_4981,N_4964);
and U5085 (N_5085,N_4061,N_4195);
nand U5086 (N_5086,N_3195,N_4253);
nand U5087 (N_5087,N_3772,N_4400);
nand U5088 (N_5088,N_2761,N_2632);
or U5089 (N_5089,N_2848,N_4090);
and U5090 (N_5090,N_4884,N_3100);
nand U5091 (N_5091,N_4874,N_3843);
nand U5092 (N_5092,N_2857,N_4105);
or U5093 (N_5093,N_3541,N_4066);
nor U5094 (N_5094,N_2618,N_4394);
or U5095 (N_5095,N_3654,N_3514);
nand U5096 (N_5096,N_2873,N_4858);
or U5097 (N_5097,N_2607,N_4237);
xor U5098 (N_5098,N_3767,N_3603);
or U5099 (N_5099,N_2746,N_2572);
or U5100 (N_5100,N_4031,N_4349);
or U5101 (N_5101,N_4524,N_3503);
or U5102 (N_5102,N_3216,N_4326);
or U5103 (N_5103,N_4920,N_3392);
nand U5104 (N_5104,N_4950,N_3705);
and U5105 (N_5105,N_3691,N_4823);
nor U5106 (N_5106,N_2772,N_4800);
nor U5107 (N_5107,N_4423,N_4666);
and U5108 (N_5108,N_2871,N_4980);
nor U5109 (N_5109,N_4043,N_3168);
nand U5110 (N_5110,N_3235,N_4261);
nand U5111 (N_5111,N_4406,N_3332);
and U5112 (N_5112,N_4750,N_3849);
nand U5113 (N_5113,N_2596,N_4306);
nor U5114 (N_5114,N_3915,N_4271);
and U5115 (N_5115,N_4035,N_4779);
nand U5116 (N_5116,N_3628,N_3679);
nor U5117 (N_5117,N_3874,N_3106);
and U5118 (N_5118,N_2724,N_2613);
nor U5119 (N_5119,N_4984,N_4093);
and U5120 (N_5120,N_4824,N_3764);
xnor U5121 (N_5121,N_3950,N_2877);
xnor U5122 (N_5122,N_3634,N_3110);
and U5123 (N_5123,N_3643,N_4116);
and U5124 (N_5124,N_2663,N_2697);
nor U5125 (N_5125,N_2561,N_4012);
nand U5126 (N_5126,N_4310,N_2633);
or U5127 (N_5127,N_2905,N_4305);
nor U5128 (N_5128,N_4765,N_4409);
or U5129 (N_5129,N_3335,N_3241);
or U5130 (N_5130,N_3425,N_3393);
xor U5131 (N_5131,N_3566,N_2550);
nand U5132 (N_5132,N_4209,N_2911);
and U5133 (N_5133,N_4538,N_4468);
or U5134 (N_5134,N_3180,N_4746);
and U5135 (N_5135,N_3420,N_4397);
or U5136 (N_5136,N_4471,N_3613);
and U5137 (N_5137,N_4982,N_2876);
nor U5138 (N_5138,N_2991,N_4702);
nand U5139 (N_5139,N_2771,N_4346);
or U5140 (N_5140,N_2666,N_4578);
or U5141 (N_5141,N_2653,N_4211);
nand U5142 (N_5142,N_4021,N_4899);
and U5143 (N_5143,N_4141,N_2891);
or U5144 (N_5144,N_3997,N_3976);
nand U5145 (N_5145,N_4572,N_3515);
or U5146 (N_5146,N_4342,N_4567);
nand U5147 (N_5147,N_4785,N_3593);
nor U5148 (N_5148,N_3459,N_3975);
nor U5149 (N_5149,N_4241,N_3258);
nor U5150 (N_5150,N_4362,N_4304);
nand U5151 (N_5151,N_3517,N_2740);
xnor U5152 (N_5152,N_4912,N_2687);
nand U5153 (N_5153,N_3886,N_4831);
and U5154 (N_5154,N_4249,N_3183);
or U5155 (N_5155,N_4904,N_3497);
and U5156 (N_5156,N_4123,N_3477);
and U5157 (N_5157,N_4482,N_3242);
or U5158 (N_5158,N_4755,N_2853);
nor U5159 (N_5159,N_3481,N_2667);
or U5160 (N_5160,N_4604,N_4995);
or U5161 (N_5161,N_3249,N_3060);
and U5162 (N_5162,N_4041,N_3261);
xor U5163 (N_5163,N_2519,N_4242);
nor U5164 (N_5164,N_3651,N_3430);
nor U5165 (N_5165,N_3895,N_4563);
nand U5166 (N_5166,N_4284,N_4870);
nand U5167 (N_5167,N_4564,N_3227);
or U5168 (N_5168,N_4348,N_3236);
nand U5169 (N_5169,N_4794,N_4484);
nor U5170 (N_5170,N_2962,N_4157);
nand U5171 (N_5171,N_4393,N_3287);
nand U5172 (N_5172,N_3052,N_3766);
nor U5173 (N_5173,N_3270,N_3265);
or U5174 (N_5174,N_4640,N_2586);
or U5175 (N_5175,N_4094,N_4959);
and U5176 (N_5176,N_3327,N_4469);
and U5177 (N_5177,N_2975,N_4380);
or U5178 (N_5178,N_4388,N_4915);
and U5179 (N_5179,N_3939,N_3166);
or U5180 (N_5180,N_3962,N_4493);
nand U5181 (N_5181,N_3179,N_4880);
nand U5182 (N_5182,N_2787,N_2644);
and U5183 (N_5183,N_3836,N_3479);
nor U5184 (N_5184,N_2851,N_3729);
nand U5185 (N_5185,N_4379,N_4257);
and U5186 (N_5186,N_2907,N_4585);
and U5187 (N_5187,N_3115,N_2528);
or U5188 (N_5188,N_4042,N_4082);
and U5189 (N_5189,N_2834,N_4177);
or U5190 (N_5190,N_2845,N_4933);
or U5191 (N_5191,N_3358,N_4451);
and U5192 (N_5192,N_3429,N_4733);
and U5193 (N_5193,N_4940,N_3486);
or U5194 (N_5194,N_3900,N_3967);
or U5195 (N_5195,N_2875,N_3108);
nand U5196 (N_5196,N_2756,N_3207);
nand U5197 (N_5197,N_4894,N_2706);
nand U5198 (N_5198,N_4756,N_2568);
nor U5199 (N_5199,N_4653,N_3293);
and U5200 (N_5200,N_3333,N_3310);
nand U5201 (N_5201,N_2709,N_3066);
and U5202 (N_5202,N_3376,N_4491);
or U5203 (N_5203,N_2737,N_3601);
or U5204 (N_5204,N_4329,N_4848);
nor U5205 (N_5205,N_4056,N_2624);
and U5206 (N_5206,N_4422,N_3586);
and U5207 (N_5207,N_4147,N_4286);
or U5208 (N_5208,N_2591,N_3462);
or U5209 (N_5209,N_3090,N_2929);
xnor U5210 (N_5210,N_3272,N_2608);
nand U5211 (N_5211,N_4410,N_4768);
nand U5212 (N_5212,N_4331,N_4944);
or U5213 (N_5213,N_4556,N_2951);
nand U5214 (N_5214,N_3695,N_3762);
nor U5215 (N_5215,N_4555,N_3123);
and U5216 (N_5216,N_4074,N_2749);
xnor U5217 (N_5217,N_3257,N_2641);
nor U5218 (N_5218,N_4532,N_4902);
and U5219 (N_5219,N_3276,N_4862);
nand U5220 (N_5220,N_2931,N_3660);
nor U5221 (N_5221,N_4692,N_4954);
nor U5222 (N_5222,N_2721,N_4158);
nand U5223 (N_5223,N_4196,N_3336);
nor U5224 (N_5224,N_2522,N_4763);
and U5225 (N_5225,N_4961,N_3058);
or U5226 (N_5226,N_3055,N_4221);
nor U5227 (N_5227,N_4676,N_3542);
or U5228 (N_5228,N_4416,N_2534);
nor U5229 (N_5229,N_4445,N_3298);
and U5230 (N_5230,N_4735,N_3700);
or U5231 (N_5231,N_2819,N_3107);
nand U5232 (N_5232,N_4392,N_3094);
nor U5233 (N_5233,N_4091,N_3154);
nand U5234 (N_5234,N_3534,N_4223);
nand U5235 (N_5235,N_3329,N_2577);
nand U5236 (N_5236,N_4027,N_3391);
or U5237 (N_5237,N_3765,N_3926);
nand U5238 (N_5238,N_4877,N_2744);
or U5239 (N_5239,N_3458,N_3259);
nand U5240 (N_5240,N_2802,N_2868);
and U5241 (N_5241,N_2604,N_3856);
nor U5242 (N_5242,N_3209,N_3378);
nand U5243 (N_5243,N_2942,N_4186);
or U5244 (N_5244,N_4973,N_2571);
nand U5245 (N_5245,N_3991,N_4450);
and U5246 (N_5246,N_4236,N_2673);
nand U5247 (N_5247,N_2773,N_4001);
nand U5248 (N_5248,N_4222,N_3850);
nor U5249 (N_5249,N_2580,N_2879);
nor U5250 (N_5250,N_3632,N_4173);
and U5251 (N_5251,N_2759,N_3956);
nand U5252 (N_5252,N_3509,N_4871);
nor U5253 (N_5253,N_2841,N_4923);
and U5254 (N_5254,N_4953,N_4396);
or U5255 (N_5255,N_4558,N_4723);
nor U5256 (N_5256,N_4553,N_3746);
or U5257 (N_5257,N_2774,N_4741);
and U5258 (N_5258,N_4174,N_2747);
or U5259 (N_5259,N_3657,N_3314);
nor U5260 (N_5260,N_3971,N_3267);
or U5261 (N_5261,N_2982,N_3897);
and U5262 (N_5262,N_2768,N_3600);
or U5263 (N_5263,N_2974,N_3042);
or U5264 (N_5264,N_4946,N_3182);
and U5265 (N_5265,N_4994,N_3868);
and U5266 (N_5266,N_2584,N_4598);
nand U5267 (N_5267,N_4167,N_2979);
nand U5268 (N_5268,N_3604,N_4266);
or U5269 (N_5269,N_3551,N_2963);
nor U5270 (N_5270,N_3513,N_2617);
and U5271 (N_5271,N_3587,N_4562);
and U5272 (N_5272,N_4227,N_2516);
nor U5273 (N_5273,N_4151,N_3716);
nand U5274 (N_5274,N_3288,N_4264);
nor U5275 (N_5275,N_3768,N_3590);
and U5276 (N_5276,N_2743,N_2593);
or U5277 (N_5277,N_3201,N_3086);
nand U5278 (N_5278,N_3942,N_3330);
nor U5279 (N_5279,N_3592,N_3262);
and U5280 (N_5280,N_4963,N_3553);
nand U5281 (N_5281,N_2898,N_4854);
and U5282 (N_5282,N_4998,N_3873);
or U5283 (N_5283,N_4296,N_4402);
and U5284 (N_5284,N_4155,N_3781);
or U5285 (N_5285,N_2527,N_3467);
nand U5286 (N_5286,N_3159,N_3363);
nand U5287 (N_5287,N_3098,N_2543);
nor U5288 (N_5288,N_4515,N_3820);
xnor U5289 (N_5289,N_3104,N_4150);
nand U5290 (N_5290,N_2569,N_4465);
and U5291 (N_5291,N_3732,N_3611);
nor U5292 (N_5292,N_4710,N_3099);
and U5293 (N_5293,N_2738,N_2692);
nor U5294 (N_5294,N_3011,N_3698);
nor U5295 (N_5295,N_3492,N_2852);
nor U5296 (N_5296,N_4922,N_3783);
nand U5297 (N_5297,N_3434,N_4417);
nor U5298 (N_5298,N_4686,N_4489);
or U5299 (N_5299,N_3761,N_3788);
and U5300 (N_5300,N_3854,N_4891);
or U5301 (N_5301,N_2887,N_2914);
or U5302 (N_5302,N_4190,N_3305);
and U5303 (N_5303,N_2884,N_2627);
nand U5304 (N_5304,N_3878,N_3318);
nor U5305 (N_5305,N_4717,N_4347);
or U5306 (N_5306,N_3271,N_3723);
nor U5307 (N_5307,N_3730,N_3161);
and U5308 (N_5308,N_4309,N_3581);
nand U5309 (N_5309,N_4808,N_2986);
or U5310 (N_5310,N_2642,N_3510);
nand U5311 (N_5311,N_2560,N_4725);
and U5312 (N_5312,N_4002,N_4013);
nor U5313 (N_5313,N_2683,N_2549);
or U5314 (N_5314,N_4139,N_3296);
or U5315 (N_5315,N_4520,N_3822);
nor U5316 (N_5316,N_2507,N_2861);
nor U5317 (N_5317,N_3715,N_4294);
and U5318 (N_5318,N_4140,N_2995);
xor U5319 (N_5319,N_2700,N_4218);
or U5320 (N_5320,N_4925,N_4714);
nand U5321 (N_5321,N_2803,N_3291);
nand U5322 (N_5322,N_3811,N_4054);
nand U5323 (N_5323,N_3582,N_4868);
nor U5324 (N_5324,N_2866,N_4519);
and U5325 (N_5325,N_3518,N_4582);
or U5326 (N_5326,N_4844,N_3782);
or U5327 (N_5327,N_4560,N_3511);
nand U5328 (N_5328,N_4525,N_2969);
and U5329 (N_5329,N_3004,N_2736);
and U5330 (N_5330,N_2732,N_4052);
nand U5331 (N_5331,N_3012,N_4951);
or U5332 (N_5332,N_2764,N_2563);
nand U5333 (N_5333,N_4752,N_3891);
and U5334 (N_5334,N_3349,N_3787);
and U5335 (N_5335,N_4770,N_3118);
or U5336 (N_5336,N_2918,N_3577);
or U5337 (N_5337,N_3313,N_3718);
nand U5338 (N_5338,N_2518,N_3116);
nor U5339 (N_5339,N_2623,N_3077);
or U5340 (N_5340,N_4599,N_4480);
or U5341 (N_5341,N_4740,N_3753);
nand U5342 (N_5342,N_3724,N_3337);
and U5343 (N_5343,N_2582,N_3250);
nor U5344 (N_5344,N_3072,N_2948);
xnor U5345 (N_5345,N_2643,N_3655);
and U5346 (N_5346,N_3331,N_3026);
and U5347 (N_5347,N_3974,N_4193);
nand U5348 (N_5348,N_4145,N_3504);
and U5349 (N_5349,N_4727,N_4918);
and U5350 (N_5350,N_4373,N_3682);
nand U5351 (N_5351,N_2984,N_3162);
nand U5352 (N_5352,N_3957,N_4220);
nand U5353 (N_5353,N_3031,N_4098);
and U5354 (N_5354,N_4660,N_3500);
nor U5355 (N_5355,N_4597,N_4488);
and U5356 (N_5356,N_4730,N_3101);
nand U5357 (N_5357,N_2946,N_2509);
or U5358 (N_5358,N_3020,N_4936);
xnor U5359 (N_5359,N_2878,N_2512);
nor U5360 (N_5360,N_3252,N_4064);
or U5361 (N_5361,N_4202,N_4118);
nor U5362 (N_5362,N_2869,N_4212);
and U5363 (N_5363,N_4019,N_3346);
or U5364 (N_5364,N_3584,N_3144);
and U5365 (N_5365,N_4112,N_3818);
and U5366 (N_5366,N_4969,N_4413);
and U5367 (N_5367,N_2558,N_4914);
nand U5368 (N_5368,N_4645,N_3837);
nand U5369 (N_5369,N_3627,N_4811);
and U5370 (N_5370,N_2978,N_3759);
nand U5371 (N_5371,N_3969,N_4804);
or U5372 (N_5372,N_2688,N_3153);
nand U5373 (N_5373,N_3689,N_4507);
or U5374 (N_5374,N_3299,N_4059);
and U5375 (N_5375,N_4967,N_2909);
nor U5376 (N_5376,N_2966,N_4203);
or U5377 (N_5377,N_3779,N_4452);
or U5378 (N_5378,N_2777,N_4955);
or U5379 (N_5379,N_4464,N_3411);
nor U5380 (N_5380,N_4295,N_3127);
or U5381 (N_5381,N_4569,N_3398);
and U5382 (N_5382,N_4467,N_4210);
nor U5383 (N_5383,N_4198,N_3588);
and U5384 (N_5384,N_3049,N_3741);
xor U5385 (N_5385,N_2842,N_3936);
and U5386 (N_5386,N_4917,N_3533);
nor U5387 (N_5387,N_3953,N_3921);
and U5388 (N_5388,N_4606,N_4711);
and U5389 (N_5389,N_3455,N_2635);
and U5390 (N_5390,N_4162,N_3778);
and U5391 (N_5391,N_4044,N_2953);
nand U5392 (N_5392,N_3062,N_4972);
nor U5393 (N_5393,N_3290,N_3297);
nand U5394 (N_5394,N_2537,N_2923);
nand U5395 (N_5395,N_3079,N_4592);
and U5396 (N_5396,N_4743,N_3087);
nand U5397 (N_5397,N_3374,N_3285);
or U5398 (N_5398,N_3263,N_4229);
nor U5399 (N_5399,N_3268,N_4016);
nand U5400 (N_5400,N_4483,N_3559);
or U5401 (N_5401,N_3930,N_2716);
and U5402 (N_5402,N_2835,N_4070);
nor U5403 (N_5403,N_3366,N_3217);
or U5404 (N_5404,N_4080,N_3403);
nand U5405 (N_5405,N_4749,N_4930);
nand U5406 (N_5406,N_3641,N_4866);
nor U5407 (N_5407,N_2755,N_2536);
xnor U5408 (N_5408,N_4620,N_3708);
nand U5409 (N_5409,N_4197,N_4820);
or U5410 (N_5410,N_3171,N_3334);
nor U5411 (N_5411,N_3576,N_4670);
nor U5412 (N_5412,N_4712,N_3648);
xnor U5413 (N_5413,N_2788,N_2664);
and U5414 (N_5414,N_3640,N_3899);
or U5415 (N_5415,N_4631,N_2694);
or U5416 (N_5416,N_2562,N_3388);
nor U5417 (N_5417,N_2718,N_4938);
nand U5418 (N_5418,N_3952,N_3827);
nor U5419 (N_5419,N_4580,N_3609);
and U5420 (N_5420,N_4504,N_4842);
and U5421 (N_5421,N_3359,N_4337);
nor U5422 (N_5422,N_3984,N_3785);
nor U5423 (N_5423,N_3360,N_4360);
or U5424 (N_5424,N_3826,N_4732);
or U5425 (N_5425,N_4602,N_3951);
or U5426 (N_5426,N_4830,N_3733);
or U5427 (N_5427,N_2708,N_3687);
nand U5428 (N_5428,N_2850,N_3901);
nand U5429 (N_5429,N_2936,N_3633);
and U5430 (N_5430,N_4230,N_3894);
nand U5431 (N_5431,N_4103,N_4087);
nor U5432 (N_5432,N_4986,N_2640);
nand U5433 (N_5433,N_4571,N_2922);
nor U5434 (N_5434,N_3968,N_2542);
and U5435 (N_5435,N_4956,N_3860);
nand U5436 (N_5436,N_3567,N_3699);
xor U5437 (N_5437,N_4603,N_4976);
nor U5438 (N_5438,N_3663,N_3131);
and U5439 (N_5439,N_4900,N_3876);
or U5440 (N_5440,N_4199,N_3711);
nor U5441 (N_5441,N_3786,N_3616);
and U5442 (N_5442,N_3771,N_3050);
and U5443 (N_5443,N_2904,N_2657);
nand U5444 (N_5444,N_4125,N_4458);
and U5445 (N_5445,N_4270,N_4506);
or U5446 (N_5446,N_3357,N_4340);
nand U5447 (N_5447,N_3117,N_3463);
nor U5448 (N_5448,N_4869,N_4274);
nor U5449 (N_5449,N_2606,N_2860);
and U5450 (N_5450,N_3917,N_4414);
nand U5451 (N_5451,N_4134,N_3549);
nand U5452 (N_5452,N_3321,N_4026);
and U5453 (N_5453,N_4239,N_2846);
and U5454 (N_5454,N_3128,N_2605);
nand U5455 (N_5455,N_3656,N_3206);
nand U5456 (N_5456,N_3596,N_4096);
and U5457 (N_5457,N_4361,N_3018);
or U5458 (N_5458,N_4790,N_4100);
or U5459 (N_5459,N_4772,N_4937);
nor U5460 (N_5460,N_3034,N_4624);
nor U5461 (N_5461,N_4101,N_4355);
and U5462 (N_5462,N_4840,N_3088);
nor U5463 (N_5463,N_2901,N_2713);
nand U5464 (N_5464,N_4443,N_3476);
nand U5465 (N_5465,N_4526,N_3306);
and U5466 (N_5466,N_3855,N_4308);
nand U5467 (N_5467,N_4822,N_4888);
nor U5468 (N_5468,N_4573,N_2968);
or U5469 (N_5469,N_3863,N_4364);
nand U5470 (N_5470,N_2616,N_3989);
nand U5471 (N_5471,N_3224,N_4251);
nor U5472 (N_5472,N_4238,N_3935);
nand U5473 (N_5473,N_2592,N_4024);
or U5474 (N_5474,N_3607,N_4613);
and U5475 (N_5475,N_3669,N_2615);
nor U5476 (N_5476,N_4133,N_3987);
and U5477 (N_5477,N_3067,N_3013);
nand U5478 (N_5478,N_3234,N_2798);
or U5479 (N_5479,N_2714,N_4492);
nor U5480 (N_5480,N_3585,N_3629);
nand U5481 (N_5481,N_3053,N_4709);
nand U5482 (N_5482,N_3483,N_4479);
nor U5483 (N_5483,N_3409,N_4508);
xor U5484 (N_5484,N_4857,N_3519);
or U5485 (N_5485,N_3036,N_2515);
or U5486 (N_5486,N_4539,N_4543);
nand U5487 (N_5487,N_3692,N_2818);
and U5488 (N_5488,N_3342,N_3960);
nor U5489 (N_5489,N_3494,N_4985);
nor U5490 (N_5490,N_2813,N_4183);
nand U5491 (N_5491,N_4172,N_2811);
xnor U5492 (N_5492,N_2647,N_2677);
nor U5493 (N_5493,N_3693,N_2958);
nor U5494 (N_5494,N_3615,N_4418);
and U5495 (N_5495,N_4076,N_3554);
and U5496 (N_5496,N_4618,N_4590);
nand U5497 (N_5497,N_2899,N_3137);
and U5498 (N_5498,N_4966,N_2839);
nand U5499 (N_5499,N_4144,N_4260);
nor U5500 (N_5500,N_4062,N_3880);
nand U5501 (N_5501,N_2973,N_2600);
nor U5502 (N_5502,N_4643,N_4459);
nor U5503 (N_5503,N_3931,N_4371);
xnor U5504 (N_5504,N_4166,N_4566);
or U5505 (N_5505,N_2530,N_2648);
and U5506 (N_5506,N_4814,N_2685);
and U5507 (N_5507,N_4656,N_3636);
nor U5508 (N_5508,N_2524,N_4909);
and U5509 (N_5509,N_4622,N_4281);
nand U5510 (N_5510,N_4832,N_3218);
or U5511 (N_5511,N_4007,N_4104);
xor U5512 (N_5512,N_2935,N_4313);
and U5513 (N_5513,N_4766,N_2676);
nor U5514 (N_5514,N_2682,N_4290);
and U5515 (N_5515,N_3598,N_4338);
or U5516 (N_5516,N_2883,N_3683);
nand U5517 (N_5517,N_4107,N_4328);
or U5518 (N_5518,N_3972,N_3805);
and U5519 (N_5519,N_2939,N_4781);
nand U5520 (N_5520,N_4159,N_3769);
nor U5521 (N_5521,N_2533,N_3830);
nand U5522 (N_5522,N_3903,N_4171);
or U5523 (N_5523,N_4330,N_3808);
and U5524 (N_5524,N_2609,N_3312);
xor U5525 (N_5525,N_3564,N_3028);
and U5526 (N_5526,N_4987,N_4385);
or U5527 (N_5527,N_3379,N_2735);
nand U5528 (N_5528,N_3919,N_4252);
or U5529 (N_5529,N_2556,N_4427);
nand U5530 (N_5530,N_3896,N_3122);
nor U5531 (N_5531,N_2662,N_3383);
nand U5532 (N_5532,N_3447,N_4415);
or U5533 (N_5533,N_4185,N_3670);
nand U5534 (N_5534,N_4399,N_3422);
or U5535 (N_5535,N_2622,N_3454);
xor U5536 (N_5536,N_4168,N_4028);
or U5537 (N_5537,N_3726,N_3922);
or U5538 (N_5538,N_3273,N_3734);
and U5539 (N_5539,N_4687,N_4272);
nor U5540 (N_5540,N_3302,N_2824);
nand U5541 (N_5541,N_2988,N_4404);
and U5542 (N_5542,N_4462,N_3631);
and U5543 (N_5543,N_4224,N_4817);
and U5544 (N_5544,N_4570,N_3416);
nand U5545 (N_5545,N_4292,N_3341);
and U5546 (N_5546,N_2987,N_3526);
nand U5547 (N_5547,N_3111,N_4789);
nand U5548 (N_5548,N_2741,N_3943);
nor U5549 (N_5549,N_2652,N_3097);
and U5550 (N_5550,N_3756,N_4847);
nor U5551 (N_5551,N_3213,N_3239);
or U5552 (N_5552,N_3591,N_3966);
or U5553 (N_5553,N_2927,N_3823);
and U5554 (N_5554,N_3438,N_3907);
nor U5555 (N_5555,N_3134,N_4293);
and U5556 (N_5556,N_3286,N_2684);
nor U5557 (N_5557,N_4511,N_4641);
and U5558 (N_5558,N_4276,N_2691);
or U5559 (N_5559,N_3124,N_4039);
xor U5560 (N_5560,N_4428,N_2924);
nor U5561 (N_5561,N_4075,N_4432);
and U5562 (N_5562,N_3372,N_4352);
and U5563 (N_5563,N_3704,N_4835);
and U5564 (N_5564,N_3869,N_4088);
or U5565 (N_5565,N_3599,N_3248);
xor U5566 (N_5566,N_4113,N_3149);
nand U5567 (N_5567,N_3375,N_2589);
nand U5568 (N_5568,N_3000,N_4705);
or U5569 (N_5569,N_3074,N_4225);
nand U5570 (N_5570,N_4748,N_4403);
and U5571 (N_5571,N_3070,N_4111);
and U5572 (N_5572,N_3441,N_3040);
or U5573 (N_5573,N_4895,N_3326);
or U5574 (N_5574,N_3697,N_4217);
nand U5575 (N_5575,N_3612,N_4420);
or U5576 (N_5576,N_4128,N_4401);
and U5577 (N_5577,N_3946,N_2894);
and U5578 (N_5578,N_2654,N_4838);
nand U5579 (N_5579,N_3246,N_2855);
nand U5580 (N_5580,N_3694,N_3839);
and U5581 (N_5581,N_2538,N_4881);
or U5582 (N_5582,N_4661,N_3913);
and U5583 (N_5583,N_3238,N_3350);
and U5584 (N_5584,N_4787,N_2546);
nand U5585 (N_5585,N_3221,N_3064);
nand U5586 (N_5586,N_4067,N_4009);
nor U5587 (N_5587,N_2906,N_2679);
and U5588 (N_5588,N_4312,N_4367);
nor U5589 (N_5589,N_2885,N_3061);
nand U5590 (N_5590,N_4689,N_2889);
and U5591 (N_5591,N_3057,N_4109);
and U5592 (N_5592,N_4188,N_3266);
nor U5593 (N_5593,N_4208,N_4815);
and U5594 (N_5594,N_3630,N_2693);
and U5595 (N_5595,N_3745,N_4023);
or U5596 (N_5596,N_4463,N_2890);
and U5597 (N_5597,N_3784,N_2897);
nand U5598 (N_5598,N_3798,N_3009);
nor U5599 (N_5599,N_3146,N_4161);
nor U5600 (N_5600,N_3789,N_3638);
and U5601 (N_5601,N_2864,N_3245);
or U5602 (N_5602,N_3156,N_2928);
nand U5603 (N_5603,N_3521,N_2965);
nand U5604 (N_5604,N_3973,N_4788);
or U5605 (N_5605,N_3776,N_3215);
nor U5606 (N_5606,N_4127,N_2595);
or U5607 (N_5607,N_3451,N_3401);
nor U5608 (N_5608,N_3738,N_2996);
and U5609 (N_5609,N_4892,N_4063);
or U5610 (N_5610,N_4997,N_3080);
and U5611 (N_5611,N_4568,N_3706);
or U5612 (N_5612,N_4398,N_3399);
nand U5613 (N_5613,N_4797,N_2545);
nand U5614 (N_5614,N_3608,N_4928);
nor U5615 (N_5615,N_4623,N_4136);
nor U5616 (N_5616,N_2808,N_4747);
nor U5617 (N_5617,N_2967,N_2983);
nand U5618 (N_5618,N_3390,N_3138);
or U5619 (N_5619,N_3712,N_4267);
and U5620 (N_5620,N_2838,N_4957);
nand U5621 (N_5621,N_4099,N_4389);
xor U5622 (N_5622,N_3446,N_4301);
nor U5623 (N_5623,N_4678,N_3384);
or U5624 (N_5624,N_3037,N_4548);
or U5625 (N_5625,N_3821,N_3557);
nand U5626 (N_5626,N_2815,N_3439);
and U5627 (N_5627,N_3714,N_2597);
or U5628 (N_5628,N_3690,N_4949);
xnor U5629 (N_5629,N_2668,N_4176);
and U5630 (N_5630,N_3255,N_4821);
or U5631 (N_5631,N_4846,N_4774);
nand U5632 (N_5632,N_3828,N_4541);
and U5633 (N_5633,N_3484,N_4910);
nor U5634 (N_5634,N_3996,N_4472);
or U5635 (N_5635,N_4051,N_2778);
nand U5636 (N_5636,N_3980,N_4048);
or U5637 (N_5637,N_3871,N_3556);
and U5638 (N_5638,N_4341,N_4703);
nor U5639 (N_5639,N_4908,N_4132);
or U5640 (N_5640,N_4863,N_3121);
and U5641 (N_5641,N_3202,N_3852);
nand U5642 (N_5642,N_4943,N_2601);
and U5643 (N_5643,N_3538,N_4707);
nand U5644 (N_5644,N_4268,N_2829);
or U5645 (N_5645,N_3370,N_2722);
nand U5646 (N_5646,N_3610,N_4855);
and U5647 (N_5647,N_3095,N_3181);
nand U5648 (N_5648,N_2598,N_4298);
and U5649 (N_5649,N_3560,N_4078);
or U5650 (N_5650,N_4890,N_3642);
nor U5651 (N_5651,N_3021,N_3910);
nor U5652 (N_5652,N_3864,N_2831);
nand U5653 (N_5653,N_4461,N_2517);
and U5654 (N_5654,N_4307,N_2754);
or U5655 (N_5655,N_2720,N_4213);
and U5656 (N_5656,N_3456,N_4235);
nor U5657 (N_5657,N_4374,N_3301);
nand U5658 (N_5658,N_4786,N_2990);
nand U5659 (N_5659,N_2867,N_2804);
nand U5660 (N_5660,N_4047,N_3279);
or U5661 (N_5661,N_4247,N_3177);
nand U5662 (N_5662,N_4170,N_4681);
nor U5663 (N_5663,N_3428,N_4574);
nor U5664 (N_5664,N_3014,N_2825);
nor U5665 (N_5665,N_4906,N_2920);
nand U5666 (N_5666,N_4089,N_3352);
nand U5667 (N_5667,N_2590,N_3949);
or U5668 (N_5668,N_3877,N_4215);
and U5669 (N_5669,N_3237,N_2726);
or U5670 (N_5670,N_2947,N_4905);
nand U5671 (N_5671,N_2753,N_2651);
nor U5672 (N_5672,N_4758,N_4505);
nand U5673 (N_5673,N_4595,N_3316);
or U5674 (N_5674,N_3594,N_3614);
nand U5675 (N_5675,N_3119,N_2817);
nor U5676 (N_5676,N_3999,N_3906);
or U5677 (N_5677,N_4030,N_3964);
and U5678 (N_5678,N_2814,N_4836);
nor U5679 (N_5679,N_2500,N_3103);
and U5680 (N_5680,N_3424,N_4079);
and U5681 (N_5681,N_4189,N_4376);
and U5682 (N_5682,N_3210,N_4856);
or U5683 (N_5683,N_4485,N_2539);
or U5684 (N_5684,N_3096,N_3016);
nor U5685 (N_5685,N_4744,N_3528);
nor U5686 (N_5686,N_4421,N_3470);
and U5687 (N_5687,N_3810,N_4356);
nor U5688 (N_5688,N_4336,N_3196);
nand U5689 (N_5689,N_3308,N_4680);
nor U5690 (N_5690,N_4165,N_4665);
and U5691 (N_5691,N_2847,N_4607);
and U5692 (N_5692,N_4350,N_3568);
and U5693 (N_5693,N_3019,N_4153);
nor U5694 (N_5694,N_3727,N_3737);
or U5695 (N_5695,N_4501,N_4557);
or U5696 (N_5696,N_2502,N_2896);
or U5697 (N_5697,N_2870,N_4206);
nand U5698 (N_5698,N_3892,N_4882);
or U5699 (N_5699,N_3703,N_4243);
nand U5700 (N_5700,N_3569,N_3686);
and U5701 (N_5701,N_3325,N_3547);
and U5702 (N_5702,N_3158,N_3003);
or U5703 (N_5703,N_4672,N_3883);
nand U5704 (N_5704,N_4444,N_2566);
nand U5705 (N_5705,N_4200,N_4497);
or U5706 (N_5706,N_4283,N_3885);
and U5707 (N_5707,N_3791,N_3774);
nor U5708 (N_5708,N_4833,N_3389);
nor U5709 (N_5709,N_3381,N_3637);
and U5710 (N_5710,N_4583,N_3445);
and U5711 (N_5711,N_4160,N_3005);
and U5712 (N_5712,N_3231,N_4500);
nand U5713 (N_5713,N_4791,N_2837);
nor U5714 (N_5714,N_3015,N_4311);
nor U5715 (N_5715,N_2506,N_4965);
and U5716 (N_5716,N_4514,N_3548);
nor U5717 (N_5717,N_3512,N_2710);
nor U5718 (N_5718,N_2999,N_3469);
nor U5719 (N_5719,N_3571,N_4591);
and U5720 (N_5720,N_2636,N_2949);
and U5721 (N_5721,N_3208,N_4934);
nor U5722 (N_5722,N_2832,N_4586);
nand U5723 (N_5723,N_2793,N_3865);
nand U5724 (N_5724,N_3954,N_2564);
and U5725 (N_5725,N_3790,N_3251);
nand U5726 (N_5726,N_3311,N_2826);
or U5727 (N_5727,N_3544,N_4332);
or U5728 (N_5728,N_3606,N_2933);
nor U5729 (N_5729,N_4826,N_4509);
and U5730 (N_5730,N_2573,N_3688);
and U5731 (N_5731,N_2541,N_3859);
nand U5732 (N_5732,N_4429,N_3324);
and U5733 (N_5733,N_3659,N_3728);
and U5734 (N_5734,N_3780,N_3552);
or U5735 (N_5735,N_3188,N_4697);
or U5736 (N_5736,N_3433,N_2611);
nor U5737 (N_5737,N_3491,N_3522);
nor U5738 (N_5738,N_4316,N_4659);
and U5739 (N_5739,N_3945,N_3888);
nand U5740 (N_5740,N_2678,N_3496);
or U5741 (N_5741,N_3032,N_3735);
and U5742 (N_5742,N_3498,N_3143);
and U5743 (N_5743,N_3872,N_3205);
nand U5744 (N_5744,N_4003,N_3775);
and U5745 (N_5745,N_4688,N_4050);
nor U5746 (N_5746,N_3406,N_4273);
or U5747 (N_5747,N_4518,N_3531);
and U5748 (N_5748,N_2950,N_4095);
nand U5749 (N_5749,N_2863,N_3934);
or U5750 (N_5750,N_2915,N_4129);
or U5751 (N_5751,N_3998,N_4040);
or U5752 (N_5752,N_3535,N_3875);
nand U5753 (N_5753,N_3666,N_2908);
nand U5754 (N_5754,N_2581,N_3758);
nor U5755 (N_5755,N_3619,N_3043);
and U5756 (N_5756,N_4551,N_3450);
nand U5757 (N_5757,N_3506,N_4187);
or U5758 (N_5758,N_2782,N_3744);
or U5759 (N_5759,N_4447,N_3147);
or U5760 (N_5760,N_4642,N_3176);
or U5761 (N_5761,N_4055,N_4547);
nand U5762 (N_5762,N_4049,N_4083);
nor U5763 (N_5763,N_3881,N_3045);
nor U5764 (N_5764,N_3817,N_3322);
nand U5765 (N_5765,N_3804,N_3833);
nor U5766 (N_5766,N_2729,N_2960);
and U5767 (N_5767,N_4754,N_4742);
or U5768 (N_5768,N_4611,N_3081);
nor U5769 (N_5769,N_3460,N_3847);
nand U5770 (N_5770,N_3536,N_4999);
or U5771 (N_5771,N_4375,N_4684);
and U5772 (N_5772,N_2742,N_4771);
and U5773 (N_5773,N_2531,N_3625);
and U5774 (N_5774,N_4581,N_3033);
nor U5775 (N_5775,N_3561,N_2760);
and U5776 (N_5776,N_3165,N_2715);
nor U5777 (N_5777,N_2791,N_4460);
and U5778 (N_5778,N_3073,N_3887);
and U5779 (N_5779,N_2961,N_2579);
and U5780 (N_5780,N_3340,N_3345);
or U5781 (N_5781,N_2766,N_3412);
nand U5782 (N_5782,N_3740,N_4860);
and U5783 (N_5783,N_2660,N_4038);
nand U5784 (N_5784,N_3039,N_4887);
nor U5785 (N_5785,N_4926,N_4231);
and U5786 (N_5786,N_3685,N_3923);
or U5787 (N_5787,N_3405,N_4793);
or U5788 (N_5788,N_2707,N_4455);
xor U5789 (N_5789,N_2576,N_4384);
nand U5790 (N_5790,N_3136,N_3395);
and U5791 (N_5791,N_3807,N_3986);
nor U5792 (N_5792,N_3944,N_4248);
xnor U5793 (N_5793,N_2783,N_4942);
nor U5794 (N_5794,N_4782,N_2769);
nor U5795 (N_5795,N_2836,N_3212);
nand U5796 (N_5796,N_3382,N_2938);
nand U5797 (N_5797,N_2565,N_2944);
nor U5798 (N_5798,N_3908,N_4279);
and U5799 (N_5799,N_4875,N_4020);
nand U5800 (N_5800,N_4246,N_2505);
and U5801 (N_5801,N_3731,N_4207);
nand U5802 (N_5802,N_4446,N_4164);
and U5803 (N_5803,N_4799,N_2523);
or U5804 (N_5804,N_3197,N_4803);
or U5805 (N_5805,N_2526,N_3125);
nor U5806 (N_5806,N_2893,N_3579);
nor U5807 (N_5807,N_4004,N_3001);
and U5808 (N_5808,N_4699,N_4287);
nor U5809 (N_5809,N_3684,N_2637);
or U5810 (N_5810,N_4865,N_4628);
nor U5811 (N_5811,N_2998,N_2723);
nand U5812 (N_5812,N_4876,N_4700);
or U5813 (N_5813,N_3461,N_3489);
or U5814 (N_5814,N_2785,N_4124);
nand U5815 (N_5815,N_3150,N_4878);
and U5816 (N_5816,N_3139,N_2959);
nand U5817 (N_5817,N_2925,N_3354);
nand U5818 (N_5818,N_4277,N_3431);
or U5819 (N_5819,N_3059,N_3889);
nor U5820 (N_5820,N_4992,N_3861);
nor U5821 (N_5821,N_3985,N_4149);
or U5822 (N_5822,N_4381,N_4931);
and U5823 (N_5823,N_3508,N_4767);
nor U5824 (N_5824,N_2752,N_4022);
or U5825 (N_5825,N_3501,N_4269);
or U5826 (N_5826,N_4448,N_3160);
nand U5827 (N_5827,N_4037,N_2882);
nor U5828 (N_5828,N_3157,N_3750);
xnor U5829 (N_5829,N_4180,N_2781);
nor U5830 (N_5830,N_4005,N_4841);
nand U5831 (N_5831,N_2681,N_3898);
nor U5832 (N_5832,N_4439,N_2547);
and U5833 (N_5833,N_3701,N_3364);
or U5834 (N_5834,N_4255,N_4728);
nor U5835 (N_5835,N_2994,N_4314);
nor U5836 (N_5836,N_2659,N_2521);
nand U5837 (N_5837,N_3233,N_3848);
and U5838 (N_5838,N_4302,N_3488);
nor U5839 (N_5839,N_2603,N_2790);
nor U5840 (N_5840,N_3665,N_3992);
nand U5841 (N_5841,N_4849,N_3002);
and U5842 (N_5842,N_3432,N_4523);
nand U5843 (N_5843,N_4609,N_4544);
nor U5844 (N_5844,N_2544,N_3427);
or U5845 (N_5845,N_4664,N_4806);
nor U5846 (N_5846,N_4114,N_3148);
and U5847 (N_5847,N_2779,N_3343);
nor U5848 (N_5848,N_3749,N_4395);
nand U5849 (N_5849,N_3419,N_3644);
or U5850 (N_5850,N_4258,N_2612);
and U5851 (N_5851,N_3068,N_4873);
and U5852 (N_5852,N_4893,N_3893);
or U5853 (N_5853,N_3482,N_2625);
or U5854 (N_5854,N_3824,N_4792);
nor U5855 (N_5855,N_3008,N_4412);
nand U5856 (N_5856,N_2823,N_3928);
or U5857 (N_5857,N_4784,N_4426);
nand U5858 (N_5858,N_3371,N_4593);
nand U5859 (N_5859,N_4530,N_4634);
and U5860 (N_5860,N_4655,N_3024);
or U5861 (N_5861,N_4575,N_4674);
nand U5862 (N_5862,N_3796,N_2776);
or U5863 (N_5863,N_4565,N_4646);
nor U5864 (N_5864,N_2730,N_3924);
and U5865 (N_5865,N_4751,N_4801);
and U5866 (N_5866,N_4718,N_2780);
nand U5867 (N_5867,N_3605,N_2599);
nand U5868 (N_5868,N_3938,N_3082);
nand U5869 (N_5869,N_3543,N_4142);
xnor U5870 (N_5870,N_4068,N_3940);
nor U5871 (N_5871,N_4760,N_4885);
and U5872 (N_5872,N_2554,N_3283);
nand U5873 (N_5873,N_3048,N_4677);
xnor U5874 (N_5874,N_4550,N_3816);
and U5875 (N_5875,N_3890,N_3870);
and U5876 (N_5876,N_2702,N_3170);
xnor U5877 (N_5877,N_3961,N_3677);
nor U5878 (N_5878,N_2680,N_2849);
nand U5879 (N_5879,N_3635,N_3193);
or U5880 (N_5880,N_3941,N_4119);
nor U5881 (N_5881,N_4032,N_2508);
or U5882 (N_5882,N_4610,N_4194);
or U5883 (N_5883,N_4425,N_3578);
nand U5884 (N_5884,N_3184,N_2650);
and U5885 (N_5885,N_3289,N_2809);
nand U5886 (N_5886,N_4204,N_4146);
nor U5887 (N_5887,N_4060,N_3958);
nand U5888 (N_5888,N_3858,N_2903);
nor U5889 (N_5889,N_4382,N_3814);
nor U5890 (N_5890,N_4179,N_3140);
xnor U5891 (N_5891,N_4839,N_4616);
xor U5892 (N_5892,N_2945,N_4993);
nor U5893 (N_5893,N_3678,N_2830);
nor U5894 (N_5894,N_3617,N_3414);
and U5895 (N_5895,N_3105,N_3415);
xor U5896 (N_5896,N_3189,N_3244);
and U5897 (N_5897,N_4813,N_4053);
or U5898 (N_5898,N_3361,N_3933);
and U5899 (N_5899,N_2649,N_2733);
and U5900 (N_5900,N_4719,N_4156);
and U5901 (N_5901,N_3046,N_2557);
nor U5902 (N_5902,N_4321,N_4708);
and U5903 (N_5903,N_3356,N_4921);
nor U5904 (N_5904,N_4737,N_3214);
and U5905 (N_5905,N_4383,N_2919);
nor U5906 (N_5906,N_2690,N_4605);
xnor U5907 (N_5907,N_3240,N_3253);
and U5908 (N_5908,N_3927,N_4736);
or U5909 (N_5909,N_2739,N_3192);
and U5910 (N_5910,N_4115,N_3194);
or U5911 (N_5911,N_4802,N_3129);
nor U5912 (N_5912,N_3126,N_3668);
nor U5913 (N_5913,N_4454,N_3373);
or U5914 (N_5914,N_4913,N_3558);
nand U5915 (N_5915,N_3440,N_2689);
or U5916 (N_5916,N_4927,N_4351);
and U5917 (N_5917,N_3710,N_2795);
or U5918 (N_5918,N_2671,N_3851);
and U5919 (N_5919,N_3529,N_4759);
nor U5920 (N_5920,N_2844,N_2725);
xnor U5921 (N_5921,N_3763,N_3575);
xnor U5922 (N_5922,N_4205,N_2786);
xor U5923 (N_5923,N_3963,N_4108);
and U5924 (N_5924,N_3646,N_2912);
nand U5925 (N_5925,N_4405,N_2672);
or U5926 (N_5926,N_4651,N_3845);
or U5927 (N_5927,N_4407,N_2638);
nand U5928 (N_5928,N_4516,N_3988);
nor U5929 (N_5929,N_3320,N_2971);
nand U5930 (N_5930,N_2658,N_4470);
and U5931 (N_5931,N_3109,N_3387);
or U5932 (N_5932,N_4635,N_2964);
or U5933 (N_5933,N_3465,N_3672);
or U5934 (N_5934,N_2807,N_3673);
and U5935 (N_5935,N_2712,N_4968);
or U5936 (N_5936,N_4630,N_4829);
and U5937 (N_5937,N_3007,N_4853);
or U5938 (N_5938,N_2794,N_3436);
and U5939 (N_5939,N_3220,N_4970);
and U5940 (N_5940,N_3502,N_2858);
nor U5941 (N_5941,N_2548,N_3932);
or U5942 (N_5942,N_4435,N_3344);
nand U5943 (N_5943,N_4796,N_4102);
xnor U5944 (N_5944,N_3574,N_4652);
nor U5945 (N_5945,N_4528,N_3219);
nand U5946 (N_5946,N_3819,N_3167);
or U5947 (N_5947,N_2529,N_4131);
and U5948 (N_5948,N_4390,N_2792);
nor U5949 (N_5949,N_2745,N_4775);
nand U5950 (N_5950,N_4667,N_3792);
nand U5951 (N_5951,N_3006,N_3929);
and U5952 (N_5952,N_4436,N_3802);
or U5953 (N_5953,N_4627,N_3597);
and U5954 (N_5954,N_4721,N_4126);
or U5955 (N_5955,N_3421,N_2575);
or U5956 (N_5956,N_3717,N_3539);
xor U5957 (N_5957,N_3555,N_3487);
nor U5958 (N_5958,N_3457,N_3368);
nor U5959 (N_5959,N_4549,N_3038);
and U5960 (N_5960,N_2943,N_4120);
nand U5961 (N_5961,N_4442,N_2840);
or U5962 (N_5962,N_3621,N_4245);
nor U5963 (N_5963,N_4654,N_4503);
or U5964 (N_5964,N_3151,N_4536);
nor U5965 (N_5965,N_4773,N_2559);
and U5966 (N_5966,N_4325,N_4932);
and U5967 (N_5967,N_2872,N_3093);
nor U5968 (N_5968,N_2567,N_3065);
nor U5969 (N_5969,N_4434,N_4029);
and U5970 (N_5970,N_4805,N_4474);
nand U5971 (N_5971,N_3937,N_4335);
or U5972 (N_5972,N_4345,N_4521);
nand U5973 (N_5973,N_2748,N_2552);
and U5974 (N_5974,N_3979,N_3920);
and U5975 (N_5975,N_4487,N_4477);
nand U5976 (N_5976,N_3112,N_3164);
and U5977 (N_5977,N_4889,N_4014);
and U5978 (N_5978,N_4476,N_3620);
or U5979 (N_5979,N_3959,N_2940);
nand U5980 (N_5980,N_3948,N_4377);
or U5981 (N_5981,N_4738,N_3914);
nand U5982 (N_5982,N_3770,N_4069);
and U5983 (N_5983,N_3468,N_4731);
and U5984 (N_5984,N_2957,N_3995);
nor U5985 (N_5985,N_4265,N_4262);
or U5986 (N_5986,N_3223,N_4638);
or U5987 (N_5987,N_3809,N_3773);
nand U5988 (N_5988,N_4685,N_3443);
nor U5989 (N_5989,N_4872,N_4698);
and U5990 (N_5990,N_4092,N_3505);
or U5991 (N_5991,N_3583,N_3978);
and U5992 (N_5992,N_4280,N_3747);
and U5993 (N_5993,N_3623,N_2588);
and U5994 (N_5994,N_3328,N_2551);
or U5995 (N_5995,N_3754,N_4675);
nor U5996 (N_5996,N_3709,N_4008);
nand U5997 (N_5997,N_4673,N_4859);
nand U5998 (N_5998,N_4701,N_2614);
and U5999 (N_5999,N_2775,N_3200);
nor U6000 (N_6000,N_4216,N_4319);
nand U6001 (N_6001,N_4576,N_3172);
and U6002 (N_6002,N_3174,N_4391);
and U6003 (N_6003,N_4299,N_2796);
and U6004 (N_6004,N_2520,N_4639);
nand U6005 (N_6005,N_3071,N_4378);
nand U6006 (N_6006,N_3982,N_2629);
nor U6007 (N_6007,N_2665,N_2525);
nor U6008 (N_6008,N_2670,N_2734);
or U6009 (N_6009,N_3573,N_3247);
and U6010 (N_6010,N_3229,N_4163);
nand U6011 (N_6011,N_4135,N_2926);
or U6012 (N_6012,N_4916,N_4184);
nor U6013 (N_6013,N_4081,N_4363);
nor U6014 (N_6014,N_2952,N_4430);
nand U6015 (N_6015,N_4977,N_2820);
or U6016 (N_6016,N_4658,N_3981);
nor U6017 (N_6017,N_4502,N_3295);
and U6018 (N_6018,N_3386,N_2504);
or U6019 (N_6019,N_2656,N_2762);
and U6020 (N_6020,N_4851,N_4561);
xnor U6021 (N_6021,N_3132,N_4776);
or U6022 (N_6022,N_3353,N_4991);
nor U6023 (N_6023,N_2806,N_2892);
and U6024 (N_6024,N_4353,N_4234);
or U6025 (N_6025,N_4358,N_3017);
nor U6026 (N_6026,N_2621,N_4512);
nand U6027 (N_6027,N_4724,N_4240);
nand U6028 (N_6028,N_2886,N_3203);
and U6029 (N_6029,N_4522,N_3076);
nand U6030 (N_6030,N_4084,N_4478);
and U6031 (N_6031,N_3707,N_3452);
or U6032 (N_6032,N_2645,N_2514);
nand U6033 (N_6033,N_4834,N_3524);
or U6034 (N_6034,N_4449,N_3626);
nand U6035 (N_6035,N_3369,N_4143);
and U6036 (N_6036,N_3916,N_4372);
nand U6037 (N_6037,N_3453,N_3317);
nor U6038 (N_6038,N_3563,N_4850);
nor U6039 (N_6039,N_4121,N_4344);
nor U6040 (N_6040,N_4974,N_4812);
nand U6041 (N_6041,N_3442,N_3163);
nor U6042 (N_6042,N_4011,N_2661);
nor U6043 (N_6043,N_2630,N_2976);
nand U6044 (N_6044,N_3879,N_4122);
nand U6045 (N_6045,N_3377,N_3970);
or U6046 (N_6046,N_3977,N_4534);
and U6047 (N_6047,N_4540,N_4695);
or U6048 (N_6048,N_3035,N_2717);
or U6049 (N_6049,N_4780,N_4679);
xnor U6050 (N_6050,N_2553,N_4761);
nor U6051 (N_6051,N_4322,N_4753);
nor U6052 (N_6052,N_3475,N_3294);
and U6053 (N_6053,N_4424,N_4365);
nor U6054 (N_6054,N_3993,N_4867);
nand U6055 (N_6055,N_3720,N_3243);
and U6056 (N_6056,N_4722,N_4990);
nor U6057 (N_6057,N_3813,N_3825);
nand U6058 (N_6058,N_3365,N_4589);
and U6059 (N_6059,N_4387,N_4919);
and U6060 (N_6060,N_2921,N_2669);
nor U6061 (N_6061,N_4045,N_4006);
or U6062 (N_6062,N_3650,N_4453);
nor U6063 (N_6063,N_3348,N_4769);
nand U6064 (N_6064,N_4696,N_4219);
nor U6065 (N_6065,N_4408,N_3054);
or U6066 (N_6066,N_3725,N_3281);
or U6067 (N_6067,N_3647,N_4669);
nor U6068 (N_6068,N_3955,N_4952);
nor U6069 (N_6069,N_4594,N_4734);
and U6070 (N_6070,N_4250,N_2930);
and U6071 (N_6071,N_4852,N_4033);
and U6072 (N_6072,N_3794,N_4626);
nand U6073 (N_6073,N_4632,N_3089);
nor U6074 (N_6074,N_3417,N_4034);
nor U6075 (N_6075,N_3187,N_4300);
or U6076 (N_6076,N_4542,N_4354);
nor U6077 (N_6077,N_2993,N_2816);
nor U6078 (N_6078,N_3846,N_3402);
nand U6079 (N_6079,N_2900,N_3925);
xor U6080 (N_6080,N_3835,N_4843);
nor U6081 (N_6081,N_3495,N_3550);
nand U6082 (N_6082,N_4816,N_2763);
nor U6083 (N_6083,N_3274,N_3674);
and U6084 (N_6084,N_4810,N_3815);
nand U6085 (N_6085,N_3499,N_4945);
or U6086 (N_6086,N_4898,N_4989);
nor U6087 (N_6087,N_3800,N_4682);
and U6088 (N_6088,N_3680,N_3842);
nor U6089 (N_6089,N_3667,N_4879);
xor U6090 (N_6090,N_2578,N_4948);
nand U6091 (N_6091,N_3178,N_4897);
or U6092 (N_6092,N_3304,N_2854);
nand U6093 (N_6093,N_3490,N_4827);
nand U6094 (N_6094,N_2503,N_4411);
or U6095 (N_6095,N_4960,N_4494);
and U6096 (N_6096,N_4729,N_4318);
and U6097 (N_6097,N_2827,N_2510);
or U6098 (N_6098,N_4621,N_3676);
nand U6099 (N_6099,N_4317,N_4473);
or U6100 (N_6100,N_4085,N_4662);
nor U6101 (N_6101,N_3022,N_3806);
and U6102 (N_6102,N_4152,N_4552);
xnor U6103 (N_6103,N_3473,N_2646);
or U6104 (N_6104,N_4323,N_4579);
nor U6105 (N_6105,N_4537,N_4130);
and U6106 (N_6106,N_3102,N_4648);
nor U6107 (N_6107,N_4587,N_2937);
nor U6108 (N_6108,N_2859,N_3622);
nor U6109 (N_6109,N_3185,N_2856);
nor U6110 (N_6110,N_4601,N_3904);
nor U6111 (N_6111,N_4057,N_4546);
nand U6112 (N_6112,N_4690,N_2619);
or U6113 (N_6113,N_4663,N_3225);
nand U6114 (N_6114,N_3478,N_2956);
nor U6115 (N_6115,N_4017,N_4693);
and U6116 (N_6116,N_4739,N_2888);
and U6117 (N_6117,N_4065,N_3844);
or U6118 (N_6118,N_2634,N_4282);
nor U6119 (N_6119,N_3722,N_3339);
nand U6120 (N_6120,N_4559,N_3719);
nand U6121 (N_6121,N_4650,N_4357);
or U6122 (N_6122,N_4636,N_3323);
and U6123 (N_6123,N_4334,N_4614);
nor U6124 (N_6124,N_3449,N_4495);
and U6125 (N_6125,N_2610,N_4818);
nor U6126 (N_6126,N_3662,N_2916);
nand U6127 (N_6127,N_4757,N_3472);
nand U6128 (N_6128,N_3029,N_2977);
or U6129 (N_6129,N_2701,N_2880);
and U6130 (N_6130,N_4181,N_3751);
or U6131 (N_6131,N_3516,N_2703);
or U6132 (N_6132,N_4809,N_2895);
nand U6133 (N_6133,N_2765,N_2594);
nand U6134 (N_6134,N_4629,N_4720);
nand U6135 (N_6135,N_4046,N_2862);
or U6136 (N_6136,N_3114,N_4864);
or U6137 (N_6137,N_2501,N_4545);
or U6138 (N_6138,N_4745,N_3507);
nor U6139 (N_6139,N_2865,N_4431);
nand U6140 (N_6140,N_3437,N_3671);
nor U6141 (N_6141,N_3909,N_3230);
nand U6142 (N_6142,N_3030,N_4036);
nand U6143 (N_6143,N_3565,N_3277);
or U6144 (N_6144,N_3380,N_4513);
xnor U6145 (N_6145,N_4010,N_2955);
nand U6146 (N_6146,N_3801,N_2513);
xor U6147 (N_6147,N_3418,N_2805);
nand U6148 (N_6148,N_3523,N_2828);
and U6149 (N_6149,N_4535,N_3527);
nor U6150 (N_6150,N_3362,N_4386);
nor U6151 (N_6151,N_2585,N_4924);
nor U6152 (N_6152,N_4988,N_4777);
nor U6153 (N_6153,N_4694,N_4554);
and U6154 (N_6154,N_3407,N_3757);
nand U6155 (N_6155,N_3570,N_3282);
nand U6156 (N_6156,N_3198,N_4798);
nand U6157 (N_6157,N_2602,N_4704);
and U6158 (N_6158,N_2801,N_3797);
nand U6159 (N_6159,N_3091,N_3044);
or U6160 (N_6160,N_2821,N_3423);
and U6161 (N_6161,N_4637,N_3152);
or U6162 (N_6162,N_3540,N_4154);
and U6163 (N_6163,N_4324,N_3911);
nand U6164 (N_6164,N_3653,N_4726);
nor U6165 (N_6165,N_3580,N_3300);
or U6166 (N_6166,N_4339,N_4861);
xnor U6167 (N_6167,N_3589,N_3075);
xor U6168 (N_6168,N_3025,N_2980);
nand U6169 (N_6169,N_4359,N_2674);
nor U6170 (N_6170,N_4437,N_3347);
or U6171 (N_6171,N_4715,N_3199);
and U6172 (N_6172,N_4907,N_2695);
or U6173 (N_6173,N_2799,N_4983);
nor U6174 (N_6174,N_4962,N_3394);
and U6175 (N_6175,N_4106,N_2626);
xnor U6176 (N_6176,N_3681,N_2932);
nor U6177 (N_6177,N_3130,N_2719);
nor U6178 (N_6178,N_4533,N_4716);
or U6179 (N_6179,N_4649,N_4327);
and U6180 (N_6180,N_3385,N_4320);
and U6181 (N_6181,N_4343,N_2631);
nand U6182 (N_6182,N_2686,N_4498);
nor U6183 (N_6183,N_4192,N_2711);
nand U6184 (N_6184,N_3232,N_3191);
nand U6185 (N_6185,N_3742,N_3884);
nand U6186 (N_6186,N_4795,N_3525);
nor U6187 (N_6187,N_4807,N_3795);
nor U6188 (N_6188,N_4315,N_4368);
nand U6189 (N_6189,N_4778,N_4644);
nor U6190 (N_6190,N_3739,N_3078);
nand U6191 (N_6191,N_4929,N_2784);
and U6192 (N_6192,N_3545,N_2532);
nand U6193 (N_6193,N_4015,N_2985);
and U6194 (N_6194,N_3010,N_2555);
nand U6195 (N_6195,N_3142,N_4527);
nand U6196 (N_6196,N_3264,N_3355);
or U6197 (N_6197,N_3396,N_3169);
nand U6198 (N_6198,N_4297,N_4819);
or U6199 (N_6199,N_3120,N_3260);
or U6200 (N_6200,N_4182,N_4706);
nand U6201 (N_6201,N_4175,N_4517);
and U6202 (N_6202,N_3047,N_3413);
nor U6203 (N_6203,N_3645,N_4657);
or U6204 (N_6204,N_4496,N_2655);
nand U6205 (N_6205,N_3464,N_2981);
nand U6206 (N_6206,N_3838,N_2941);
and U6207 (N_6207,N_4071,N_4947);
xnor U6208 (N_6208,N_4433,N_4971);
nor U6209 (N_6209,N_4584,N_3624);
or U6210 (N_6210,N_3572,N_3069);
and U6211 (N_6211,N_3841,N_3983);
or U6212 (N_6212,N_3226,N_4633);
or U6213 (N_6213,N_3303,N_4883);
nand U6214 (N_6214,N_2843,N_3702);
nor U6215 (N_6215,N_4596,N_4226);
nand U6216 (N_6216,N_4762,N_4939);
nand U6217 (N_6217,N_4438,N_3204);
and U6218 (N_6218,N_3882,N_3307);
and U6219 (N_6219,N_3400,N_4612);
nand U6220 (N_6220,N_3721,N_3793);
nand U6221 (N_6221,N_4440,N_4466);
nand U6222 (N_6222,N_3278,N_3853);
or U6223 (N_6223,N_2797,N_2970);
or U6224 (N_6224,N_4886,N_3994);
or U6225 (N_6225,N_4901,N_3175);
nand U6226 (N_6226,N_2881,N_3485);
or U6227 (N_6227,N_4058,N_4499);
nor U6228 (N_6228,N_2812,N_4137);
nand U6229 (N_6229,N_4958,N_3649);
nand U6230 (N_6230,N_4615,N_3474);
and U6231 (N_6231,N_4647,N_2727);
nand U6232 (N_6232,N_3661,N_3056);
or U6233 (N_6233,N_2587,N_4018);
and U6234 (N_6234,N_2954,N_4214);
or U6235 (N_6235,N_4457,N_3269);
or U6236 (N_6236,N_4256,N_3752);
and U6237 (N_6237,N_2934,N_2751);
nor U6238 (N_6238,N_2770,N_3546);
and U6239 (N_6239,N_3319,N_3652);
nor U6240 (N_6240,N_3426,N_3404);
nand U6241 (N_6241,N_3748,N_4668);
or U6242 (N_6242,N_3051,N_3448);
or U6243 (N_6243,N_4845,N_4097);
nand U6244 (N_6244,N_4713,N_4481);
or U6245 (N_6245,N_2972,N_4456);
nand U6246 (N_6246,N_4278,N_3902);
and U6247 (N_6247,N_3083,N_4077);
nor U6248 (N_6248,N_3145,N_2699);
nor U6249 (N_6249,N_3027,N_3812);
and U6250 (N_6250,N_4572,N_4634);
nor U6251 (N_6251,N_4028,N_2916);
nand U6252 (N_6252,N_3535,N_4177);
or U6253 (N_6253,N_4985,N_3574);
and U6254 (N_6254,N_3381,N_3040);
nand U6255 (N_6255,N_4010,N_4400);
xor U6256 (N_6256,N_3035,N_3102);
nor U6257 (N_6257,N_4981,N_2895);
nand U6258 (N_6258,N_4299,N_3686);
and U6259 (N_6259,N_3613,N_3761);
and U6260 (N_6260,N_3375,N_4996);
and U6261 (N_6261,N_3363,N_4604);
nor U6262 (N_6262,N_3345,N_3080);
or U6263 (N_6263,N_4665,N_4896);
and U6264 (N_6264,N_2814,N_2740);
and U6265 (N_6265,N_2956,N_3554);
nand U6266 (N_6266,N_3829,N_2670);
nor U6267 (N_6267,N_2949,N_2529);
nand U6268 (N_6268,N_4386,N_3371);
or U6269 (N_6269,N_4704,N_2657);
nor U6270 (N_6270,N_4575,N_2572);
or U6271 (N_6271,N_3872,N_4746);
nand U6272 (N_6272,N_3793,N_2846);
nor U6273 (N_6273,N_2572,N_3007);
nand U6274 (N_6274,N_4841,N_3696);
nand U6275 (N_6275,N_3345,N_3195);
nor U6276 (N_6276,N_4084,N_4881);
or U6277 (N_6277,N_3904,N_2956);
nand U6278 (N_6278,N_3025,N_3305);
and U6279 (N_6279,N_3771,N_2649);
nand U6280 (N_6280,N_4511,N_3214);
nor U6281 (N_6281,N_2853,N_3649);
nand U6282 (N_6282,N_3321,N_2870);
or U6283 (N_6283,N_4561,N_2991);
or U6284 (N_6284,N_3141,N_4121);
or U6285 (N_6285,N_4984,N_4778);
or U6286 (N_6286,N_3633,N_2709);
nand U6287 (N_6287,N_3716,N_4662);
nor U6288 (N_6288,N_4745,N_3018);
nor U6289 (N_6289,N_4655,N_3962);
nor U6290 (N_6290,N_4555,N_4594);
nand U6291 (N_6291,N_4898,N_2812);
and U6292 (N_6292,N_4457,N_3088);
nand U6293 (N_6293,N_4736,N_4152);
and U6294 (N_6294,N_4256,N_2734);
xor U6295 (N_6295,N_3516,N_2829);
and U6296 (N_6296,N_2869,N_4339);
nand U6297 (N_6297,N_3278,N_3022);
xnor U6298 (N_6298,N_4986,N_3668);
nor U6299 (N_6299,N_2896,N_3652);
nand U6300 (N_6300,N_4726,N_3132);
and U6301 (N_6301,N_2813,N_2715);
and U6302 (N_6302,N_4466,N_2865);
or U6303 (N_6303,N_2967,N_4907);
nand U6304 (N_6304,N_2516,N_4925);
nor U6305 (N_6305,N_3455,N_4398);
nor U6306 (N_6306,N_4994,N_3707);
nand U6307 (N_6307,N_3832,N_4050);
nand U6308 (N_6308,N_4006,N_3326);
nand U6309 (N_6309,N_2506,N_4810);
or U6310 (N_6310,N_3014,N_4962);
nand U6311 (N_6311,N_4571,N_3410);
and U6312 (N_6312,N_3499,N_3074);
nand U6313 (N_6313,N_2507,N_3732);
nor U6314 (N_6314,N_4898,N_3150);
nand U6315 (N_6315,N_4357,N_3004);
or U6316 (N_6316,N_2924,N_4112);
nor U6317 (N_6317,N_3963,N_4351);
or U6318 (N_6318,N_2526,N_3412);
nor U6319 (N_6319,N_3722,N_3525);
nand U6320 (N_6320,N_2656,N_4653);
nor U6321 (N_6321,N_4638,N_3189);
and U6322 (N_6322,N_2517,N_3564);
and U6323 (N_6323,N_2561,N_4111);
or U6324 (N_6324,N_2521,N_2554);
and U6325 (N_6325,N_2869,N_4221);
and U6326 (N_6326,N_2885,N_4872);
nand U6327 (N_6327,N_2501,N_4866);
nand U6328 (N_6328,N_4408,N_4076);
and U6329 (N_6329,N_4307,N_2935);
and U6330 (N_6330,N_3562,N_3519);
or U6331 (N_6331,N_4210,N_4538);
or U6332 (N_6332,N_2974,N_4481);
or U6333 (N_6333,N_4689,N_3667);
and U6334 (N_6334,N_2788,N_4873);
and U6335 (N_6335,N_4995,N_4780);
nor U6336 (N_6336,N_2984,N_3224);
or U6337 (N_6337,N_4126,N_3900);
and U6338 (N_6338,N_3969,N_4437);
nor U6339 (N_6339,N_4860,N_3188);
or U6340 (N_6340,N_3702,N_3428);
and U6341 (N_6341,N_4503,N_3996);
nand U6342 (N_6342,N_3678,N_3255);
nand U6343 (N_6343,N_2767,N_4258);
xor U6344 (N_6344,N_4984,N_2778);
and U6345 (N_6345,N_3324,N_2891);
nor U6346 (N_6346,N_4988,N_3304);
nor U6347 (N_6347,N_4855,N_4881);
nand U6348 (N_6348,N_3503,N_3924);
xor U6349 (N_6349,N_4934,N_2775);
nand U6350 (N_6350,N_4098,N_4825);
or U6351 (N_6351,N_3809,N_4933);
and U6352 (N_6352,N_3145,N_4508);
xor U6353 (N_6353,N_2658,N_3611);
nor U6354 (N_6354,N_2608,N_4723);
and U6355 (N_6355,N_3768,N_3623);
or U6356 (N_6356,N_4846,N_2902);
and U6357 (N_6357,N_2871,N_3507);
nand U6358 (N_6358,N_4160,N_2889);
nor U6359 (N_6359,N_3195,N_3788);
and U6360 (N_6360,N_4909,N_4992);
nor U6361 (N_6361,N_2923,N_2969);
or U6362 (N_6362,N_2963,N_3987);
or U6363 (N_6363,N_3011,N_2812);
nand U6364 (N_6364,N_3446,N_2749);
and U6365 (N_6365,N_3117,N_3121);
or U6366 (N_6366,N_3670,N_2535);
nand U6367 (N_6367,N_4331,N_2594);
and U6368 (N_6368,N_3822,N_3935);
nor U6369 (N_6369,N_3276,N_3129);
and U6370 (N_6370,N_4436,N_4887);
xor U6371 (N_6371,N_3673,N_4333);
xor U6372 (N_6372,N_2639,N_2597);
nor U6373 (N_6373,N_3683,N_2719);
or U6374 (N_6374,N_4576,N_4949);
xor U6375 (N_6375,N_3625,N_3412);
nor U6376 (N_6376,N_2980,N_2844);
nor U6377 (N_6377,N_4670,N_3125);
or U6378 (N_6378,N_2762,N_2820);
nor U6379 (N_6379,N_4535,N_3186);
or U6380 (N_6380,N_4628,N_3522);
and U6381 (N_6381,N_2575,N_4864);
nor U6382 (N_6382,N_2894,N_3227);
or U6383 (N_6383,N_3536,N_3050);
and U6384 (N_6384,N_2511,N_4488);
xnor U6385 (N_6385,N_4288,N_4637);
nand U6386 (N_6386,N_2838,N_4966);
nor U6387 (N_6387,N_4852,N_2935);
and U6388 (N_6388,N_4344,N_4305);
nor U6389 (N_6389,N_2526,N_2569);
or U6390 (N_6390,N_4818,N_4776);
or U6391 (N_6391,N_3161,N_3558);
and U6392 (N_6392,N_2866,N_4784);
nor U6393 (N_6393,N_3943,N_3518);
and U6394 (N_6394,N_4102,N_4237);
nor U6395 (N_6395,N_3564,N_3464);
nor U6396 (N_6396,N_3285,N_4598);
or U6397 (N_6397,N_3804,N_4167);
nand U6398 (N_6398,N_4255,N_3672);
or U6399 (N_6399,N_3885,N_3592);
or U6400 (N_6400,N_4660,N_3864);
and U6401 (N_6401,N_4401,N_2521);
or U6402 (N_6402,N_4365,N_2996);
nor U6403 (N_6403,N_2595,N_3195);
or U6404 (N_6404,N_3740,N_3785);
nor U6405 (N_6405,N_3339,N_2871);
and U6406 (N_6406,N_4952,N_2640);
or U6407 (N_6407,N_3920,N_2738);
nand U6408 (N_6408,N_3626,N_2553);
nand U6409 (N_6409,N_4081,N_3199);
nor U6410 (N_6410,N_3241,N_3921);
nand U6411 (N_6411,N_3626,N_3373);
or U6412 (N_6412,N_2758,N_4394);
and U6413 (N_6413,N_3231,N_4176);
and U6414 (N_6414,N_4925,N_3039);
nand U6415 (N_6415,N_3620,N_4614);
and U6416 (N_6416,N_3583,N_2791);
or U6417 (N_6417,N_4359,N_4569);
nand U6418 (N_6418,N_3124,N_2645);
and U6419 (N_6419,N_2926,N_3048);
nand U6420 (N_6420,N_4872,N_4827);
or U6421 (N_6421,N_2701,N_2636);
nand U6422 (N_6422,N_2854,N_3026);
or U6423 (N_6423,N_3794,N_4544);
or U6424 (N_6424,N_3382,N_4052);
and U6425 (N_6425,N_3942,N_3731);
nand U6426 (N_6426,N_4806,N_4437);
nor U6427 (N_6427,N_4798,N_4684);
and U6428 (N_6428,N_3005,N_4535);
and U6429 (N_6429,N_3553,N_4949);
and U6430 (N_6430,N_4095,N_3605);
nand U6431 (N_6431,N_4790,N_4389);
or U6432 (N_6432,N_2879,N_4281);
nor U6433 (N_6433,N_4243,N_3523);
or U6434 (N_6434,N_4566,N_4663);
nor U6435 (N_6435,N_3556,N_2813);
nand U6436 (N_6436,N_3407,N_2974);
xnor U6437 (N_6437,N_2534,N_3309);
or U6438 (N_6438,N_4505,N_4194);
and U6439 (N_6439,N_2639,N_3612);
nand U6440 (N_6440,N_2955,N_3795);
nor U6441 (N_6441,N_4914,N_4777);
nor U6442 (N_6442,N_3773,N_2658);
nor U6443 (N_6443,N_4037,N_4818);
nand U6444 (N_6444,N_3068,N_3724);
nor U6445 (N_6445,N_2976,N_3029);
nor U6446 (N_6446,N_3955,N_3405);
and U6447 (N_6447,N_3963,N_3787);
nor U6448 (N_6448,N_2695,N_2795);
and U6449 (N_6449,N_3716,N_3024);
nand U6450 (N_6450,N_3247,N_3555);
or U6451 (N_6451,N_4360,N_3760);
nor U6452 (N_6452,N_4960,N_4622);
xnor U6453 (N_6453,N_3750,N_3560);
or U6454 (N_6454,N_3307,N_4507);
and U6455 (N_6455,N_4727,N_3733);
nand U6456 (N_6456,N_3482,N_3298);
or U6457 (N_6457,N_3616,N_4032);
or U6458 (N_6458,N_2836,N_2940);
nor U6459 (N_6459,N_3418,N_4194);
nand U6460 (N_6460,N_4055,N_2594);
nand U6461 (N_6461,N_3819,N_4975);
and U6462 (N_6462,N_4850,N_4822);
nor U6463 (N_6463,N_3985,N_4327);
nand U6464 (N_6464,N_3135,N_4058);
and U6465 (N_6465,N_2585,N_4451);
nor U6466 (N_6466,N_4796,N_4078);
nand U6467 (N_6467,N_4859,N_4371);
nand U6468 (N_6468,N_3216,N_2733);
nand U6469 (N_6469,N_3416,N_4196);
or U6470 (N_6470,N_2811,N_4792);
and U6471 (N_6471,N_3624,N_3153);
nand U6472 (N_6472,N_4646,N_3088);
or U6473 (N_6473,N_4813,N_4309);
nor U6474 (N_6474,N_2600,N_3695);
nand U6475 (N_6475,N_4318,N_4074);
nor U6476 (N_6476,N_4808,N_3150);
and U6477 (N_6477,N_3643,N_3207);
nand U6478 (N_6478,N_4226,N_2699);
nand U6479 (N_6479,N_3338,N_4959);
nor U6480 (N_6480,N_4894,N_3408);
nand U6481 (N_6481,N_3820,N_3988);
nand U6482 (N_6482,N_3270,N_4444);
or U6483 (N_6483,N_4069,N_3280);
and U6484 (N_6484,N_2695,N_4011);
and U6485 (N_6485,N_4645,N_2800);
nand U6486 (N_6486,N_3567,N_3178);
and U6487 (N_6487,N_3306,N_4812);
and U6488 (N_6488,N_4478,N_4884);
or U6489 (N_6489,N_4563,N_3503);
nor U6490 (N_6490,N_2595,N_2826);
and U6491 (N_6491,N_4990,N_2666);
nor U6492 (N_6492,N_4181,N_4515);
or U6493 (N_6493,N_4927,N_2655);
nor U6494 (N_6494,N_4672,N_3050);
or U6495 (N_6495,N_2516,N_3340);
and U6496 (N_6496,N_4702,N_3087);
or U6497 (N_6497,N_3765,N_3144);
and U6498 (N_6498,N_3942,N_3564);
xnor U6499 (N_6499,N_3074,N_2803);
and U6500 (N_6500,N_3880,N_3239);
or U6501 (N_6501,N_3922,N_4177);
or U6502 (N_6502,N_2740,N_4432);
or U6503 (N_6503,N_4161,N_4259);
and U6504 (N_6504,N_3878,N_3373);
xor U6505 (N_6505,N_4598,N_3737);
nor U6506 (N_6506,N_3904,N_2741);
and U6507 (N_6507,N_2593,N_4626);
or U6508 (N_6508,N_2812,N_4418);
nor U6509 (N_6509,N_4118,N_3982);
or U6510 (N_6510,N_4909,N_4603);
and U6511 (N_6511,N_4069,N_3580);
and U6512 (N_6512,N_3598,N_3984);
nand U6513 (N_6513,N_2670,N_3313);
and U6514 (N_6514,N_2888,N_3802);
or U6515 (N_6515,N_4732,N_3865);
nand U6516 (N_6516,N_4850,N_2914);
or U6517 (N_6517,N_4585,N_3181);
and U6518 (N_6518,N_2892,N_4823);
or U6519 (N_6519,N_4182,N_4684);
or U6520 (N_6520,N_2605,N_2813);
xor U6521 (N_6521,N_4185,N_4701);
and U6522 (N_6522,N_3589,N_4247);
and U6523 (N_6523,N_3800,N_3488);
nor U6524 (N_6524,N_2964,N_3167);
nand U6525 (N_6525,N_4610,N_3254);
nand U6526 (N_6526,N_3906,N_3287);
or U6527 (N_6527,N_4812,N_4242);
nor U6528 (N_6528,N_3225,N_4735);
or U6529 (N_6529,N_4049,N_2799);
and U6530 (N_6530,N_4883,N_2523);
or U6531 (N_6531,N_4294,N_3198);
or U6532 (N_6532,N_3841,N_4138);
nand U6533 (N_6533,N_4806,N_3180);
and U6534 (N_6534,N_3118,N_3560);
nor U6535 (N_6535,N_3528,N_3376);
nor U6536 (N_6536,N_2589,N_4569);
nor U6537 (N_6537,N_3365,N_3192);
and U6538 (N_6538,N_3616,N_4384);
nand U6539 (N_6539,N_3807,N_4403);
or U6540 (N_6540,N_3930,N_4599);
and U6541 (N_6541,N_2785,N_3333);
nor U6542 (N_6542,N_4107,N_3812);
and U6543 (N_6543,N_3367,N_3438);
xor U6544 (N_6544,N_3730,N_3853);
xor U6545 (N_6545,N_3391,N_3395);
or U6546 (N_6546,N_4352,N_3277);
or U6547 (N_6547,N_3644,N_2928);
nor U6548 (N_6548,N_3543,N_3560);
xnor U6549 (N_6549,N_4437,N_3353);
or U6550 (N_6550,N_4590,N_3768);
nand U6551 (N_6551,N_4886,N_4363);
or U6552 (N_6552,N_4002,N_4909);
and U6553 (N_6553,N_2932,N_2939);
nor U6554 (N_6554,N_3822,N_4465);
or U6555 (N_6555,N_4178,N_4682);
or U6556 (N_6556,N_2685,N_2916);
and U6557 (N_6557,N_2775,N_2906);
xnor U6558 (N_6558,N_4282,N_3265);
and U6559 (N_6559,N_2841,N_3538);
nor U6560 (N_6560,N_3348,N_3559);
or U6561 (N_6561,N_4454,N_2703);
nor U6562 (N_6562,N_3157,N_4492);
and U6563 (N_6563,N_4158,N_3896);
nor U6564 (N_6564,N_2566,N_4166);
or U6565 (N_6565,N_3877,N_3287);
or U6566 (N_6566,N_3562,N_3864);
or U6567 (N_6567,N_3433,N_4827);
and U6568 (N_6568,N_4233,N_4449);
nor U6569 (N_6569,N_3372,N_2854);
nand U6570 (N_6570,N_3811,N_3609);
or U6571 (N_6571,N_3939,N_4784);
nor U6572 (N_6572,N_2774,N_2562);
nand U6573 (N_6573,N_3974,N_3890);
nand U6574 (N_6574,N_4409,N_3742);
or U6575 (N_6575,N_2760,N_4131);
nand U6576 (N_6576,N_3708,N_4718);
nor U6577 (N_6577,N_3396,N_2837);
and U6578 (N_6578,N_3582,N_3450);
nand U6579 (N_6579,N_4300,N_4464);
nor U6580 (N_6580,N_2663,N_4388);
or U6581 (N_6581,N_3063,N_4338);
nand U6582 (N_6582,N_4519,N_3673);
nand U6583 (N_6583,N_4239,N_3773);
nor U6584 (N_6584,N_4067,N_3358);
or U6585 (N_6585,N_2876,N_4566);
nor U6586 (N_6586,N_3541,N_4888);
nor U6587 (N_6587,N_3797,N_3923);
nor U6588 (N_6588,N_4927,N_3226);
nor U6589 (N_6589,N_3031,N_3048);
nand U6590 (N_6590,N_3391,N_3875);
nor U6591 (N_6591,N_3269,N_3863);
nor U6592 (N_6592,N_4094,N_3783);
or U6593 (N_6593,N_4618,N_4042);
or U6594 (N_6594,N_3544,N_3216);
or U6595 (N_6595,N_4231,N_4467);
nand U6596 (N_6596,N_2568,N_2640);
nor U6597 (N_6597,N_4258,N_4516);
nand U6598 (N_6598,N_3576,N_3790);
nand U6599 (N_6599,N_4179,N_2715);
nor U6600 (N_6600,N_3605,N_4538);
or U6601 (N_6601,N_2975,N_4952);
and U6602 (N_6602,N_3872,N_2809);
nand U6603 (N_6603,N_4184,N_4629);
or U6604 (N_6604,N_4153,N_3454);
nand U6605 (N_6605,N_3369,N_3654);
nor U6606 (N_6606,N_3614,N_2909);
nor U6607 (N_6607,N_3538,N_2791);
and U6608 (N_6608,N_3670,N_4783);
nor U6609 (N_6609,N_4081,N_3662);
nand U6610 (N_6610,N_4095,N_2836);
nand U6611 (N_6611,N_3438,N_3959);
nand U6612 (N_6612,N_4440,N_3073);
nor U6613 (N_6613,N_3290,N_2669);
or U6614 (N_6614,N_3689,N_3077);
or U6615 (N_6615,N_4460,N_4626);
or U6616 (N_6616,N_3618,N_3596);
nor U6617 (N_6617,N_4967,N_2746);
and U6618 (N_6618,N_3949,N_2614);
nor U6619 (N_6619,N_3239,N_3931);
nand U6620 (N_6620,N_3458,N_3982);
and U6621 (N_6621,N_3058,N_3925);
nand U6622 (N_6622,N_4214,N_3867);
and U6623 (N_6623,N_3672,N_3396);
nand U6624 (N_6624,N_3328,N_3081);
nand U6625 (N_6625,N_2872,N_2801);
or U6626 (N_6626,N_3725,N_2959);
and U6627 (N_6627,N_4676,N_4370);
xnor U6628 (N_6628,N_4923,N_3825);
nand U6629 (N_6629,N_3272,N_2692);
or U6630 (N_6630,N_2535,N_4275);
nor U6631 (N_6631,N_2734,N_4203);
or U6632 (N_6632,N_3072,N_4550);
and U6633 (N_6633,N_4334,N_4033);
and U6634 (N_6634,N_4601,N_4854);
and U6635 (N_6635,N_2823,N_4019);
xor U6636 (N_6636,N_4645,N_3632);
nor U6637 (N_6637,N_4371,N_3316);
nor U6638 (N_6638,N_3463,N_4589);
xor U6639 (N_6639,N_2924,N_3041);
and U6640 (N_6640,N_3353,N_3019);
or U6641 (N_6641,N_3678,N_2621);
nand U6642 (N_6642,N_3000,N_4279);
nor U6643 (N_6643,N_4937,N_3235);
or U6644 (N_6644,N_3576,N_3411);
nor U6645 (N_6645,N_3925,N_4432);
and U6646 (N_6646,N_4695,N_2776);
nor U6647 (N_6647,N_2508,N_2570);
or U6648 (N_6648,N_3306,N_4614);
nor U6649 (N_6649,N_2507,N_2852);
nor U6650 (N_6650,N_4809,N_4674);
nor U6651 (N_6651,N_4809,N_3363);
or U6652 (N_6652,N_4076,N_4928);
nor U6653 (N_6653,N_3567,N_2757);
or U6654 (N_6654,N_2943,N_4253);
or U6655 (N_6655,N_3489,N_2611);
nand U6656 (N_6656,N_4092,N_3866);
or U6657 (N_6657,N_3234,N_3421);
and U6658 (N_6658,N_3051,N_3208);
nor U6659 (N_6659,N_4165,N_2967);
or U6660 (N_6660,N_3562,N_2561);
nor U6661 (N_6661,N_3295,N_3559);
nor U6662 (N_6662,N_4700,N_4435);
nand U6663 (N_6663,N_4502,N_2697);
nor U6664 (N_6664,N_4553,N_3627);
nor U6665 (N_6665,N_3899,N_4490);
and U6666 (N_6666,N_4618,N_3341);
nor U6667 (N_6667,N_4908,N_2907);
and U6668 (N_6668,N_4046,N_3864);
or U6669 (N_6669,N_2681,N_4012);
xor U6670 (N_6670,N_4034,N_4531);
nand U6671 (N_6671,N_3548,N_4165);
nand U6672 (N_6672,N_3437,N_4146);
and U6673 (N_6673,N_3058,N_3240);
nor U6674 (N_6674,N_3383,N_4441);
nor U6675 (N_6675,N_4129,N_3935);
nand U6676 (N_6676,N_3277,N_4877);
and U6677 (N_6677,N_4458,N_3051);
and U6678 (N_6678,N_3148,N_3782);
nor U6679 (N_6679,N_3265,N_4725);
nand U6680 (N_6680,N_2724,N_3616);
nor U6681 (N_6681,N_2525,N_3026);
nor U6682 (N_6682,N_3573,N_4198);
nor U6683 (N_6683,N_4788,N_4010);
nor U6684 (N_6684,N_4260,N_4175);
or U6685 (N_6685,N_3857,N_3614);
nand U6686 (N_6686,N_3796,N_3867);
nor U6687 (N_6687,N_4118,N_3972);
nand U6688 (N_6688,N_4862,N_2511);
or U6689 (N_6689,N_3415,N_4154);
nor U6690 (N_6690,N_3782,N_4895);
or U6691 (N_6691,N_4203,N_3649);
or U6692 (N_6692,N_3753,N_3381);
or U6693 (N_6693,N_2569,N_4545);
nor U6694 (N_6694,N_2849,N_3762);
or U6695 (N_6695,N_2955,N_4124);
nor U6696 (N_6696,N_2937,N_3508);
and U6697 (N_6697,N_3552,N_4734);
and U6698 (N_6698,N_4201,N_3774);
or U6699 (N_6699,N_2740,N_3640);
xor U6700 (N_6700,N_4619,N_3080);
or U6701 (N_6701,N_4825,N_3059);
nand U6702 (N_6702,N_2943,N_4974);
nor U6703 (N_6703,N_2625,N_3780);
and U6704 (N_6704,N_2739,N_4537);
nand U6705 (N_6705,N_4914,N_3051);
nand U6706 (N_6706,N_4047,N_4574);
or U6707 (N_6707,N_4307,N_4536);
nand U6708 (N_6708,N_4861,N_4624);
nand U6709 (N_6709,N_4305,N_4179);
xnor U6710 (N_6710,N_4714,N_2875);
xor U6711 (N_6711,N_2904,N_3581);
nor U6712 (N_6712,N_4897,N_3923);
nor U6713 (N_6713,N_4808,N_3930);
xnor U6714 (N_6714,N_2960,N_3263);
nand U6715 (N_6715,N_3827,N_3872);
nor U6716 (N_6716,N_4007,N_4429);
nor U6717 (N_6717,N_4012,N_3264);
nor U6718 (N_6718,N_2514,N_3369);
nor U6719 (N_6719,N_2771,N_4734);
nand U6720 (N_6720,N_3655,N_4041);
nand U6721 (N_6721,N_4010,N_3247);
or U6722 (N_6722,N_4841,N_3996);
nor U6723 (N_6723,N_4269,N_3443);
xor U6724 (N_6724,N_3650,N_3732);
nand U6725 (N_6725,N_4869,N_3791);
and U6726 (N_6726,N_4472,N_2575);
and U6727 (N_6727,N_3324,N_4550);
nand U6728 (N_6728,N_3727,N_2562);
or U6729 (N_6729,N_3196,N_3423);
nor U6730 (N_6730,N_2515,N_4186);
nand U6731 (N_6731,N_4833,N_4479);
nand U6732 (N_6732,N_3929,N_4865);
or U6733 (N_6733,N_3117,N_2660);
nor U6734 (N_6734,N_4535,N_3034);
or U6735 (N_6735,N_4298,N_2579);
and U6736 (N_6736,N_4887,N_4575);
nor U6737 (N_6737,N_3585,N_2769);
nand U6738 (N_6738,N_4829,N_4485);
nor U6739 (N_6739,N_4842,N_3667);
and U6740 (N_6740,N_3784,N_4045);
nor U6741 (N_6741,N_4986,N_3956);
xnor U6742 (N_6742,N_2691,N_4550);
nor U6743 (N_6743,N_2763,N_3125);
nor U6744 (N_6744,N_3368,N_2950);
nand U6745 (N_6745,N_4160,N_2909);
nor U6746 (N_6746,N_3330,N_4773);
xor U6747 (N_6747,N_4621,N_2983);
or U6748 (N_6748,N_4024,N_3903);
and U6749 (N_6749,N_3989,N_4568);
or U6750 (N_6750,N_3726,N_3698);
nor U6751 (N_6751,N_3948,N_2689);
nand U6752 (N_6752,N_3876,N_4222);
nand U6753 (N_6753,N_3569,N_3654);
or U6754 (N_6754,N_3950,N_4393);
and U6755 (N_6755,N_3571,N_4081);
and U6756 (N_6756,N_4014,N_4377);
and U6757 (N_6757,N_4862,N_4805);
nor U6758 (N_6758,N_2611,N_3670);
nand U6759 (N_6759,N_4801,N_4273);
nor U6760 (N_6760,N_4727,N_3499);
nor U6761 (N_6761,N_2942,N_4264);
or U6762 (N_6762,N_3752,N_4322);
and U6763 (N_6763,N_3434,N_4953);
nor U6764 (N_6764,N_3018,N_2902);
nand U6765 (N_6765,N_3914,N_2521);
or U6766 (N_6766,N_4610,N_3690);
and U6767 (N_6767,N_4251,N_3471);
and U6768 (N_6768,N_4411,N_2904);
and U6769 (N_6769,N_4388,N_4788);
or U6770 (N_6770,N_3244,N_4955);
nor U6771 (N_6771,N_3089,N_3075);
or U6772 (N_6772,N_3044,N_4586);
nand U6773 (N_6773,N_4891,N_3677);
and U6774 (N_6774,N_3498,N_3944);
xor U6775 (N_6775,N_4888,N_4938);
and U6776 (N_6776,N_2772,N_3363);
nor U6777 (N_6777,N_3847,N_3130);
or U6778 (N_6778,N_4710,N_2647);
nand U6779 (N_6779,N_3161,N_4706);
nand U6780 (N_6780,N_4694,N_3691);
nor U6781 (N_6781,N_4141,N_4826);
or U6782 (N_6782,N_3752,N_4919);
or U6783 (N_6783,N_4974,N_4534);
and U6784 (N_6784,N_4647,N_2730);
nand U6785 (N_6785,N_2693,N_2932);
nor U6786 (N_6786,N_2832,N_4322);
or U6787 (N_6787,N_3735,N_3210);
or U6788 (N_6788,N_4775,N_3593);
nand U6789 (N_6789,N_2958,N_2562);
nor U6790 (N_6790,N_3001,N_3075);
and U6791 (N_6791,N_4623,N_3971);
and U6792 (N_6792,N_2592,N_4104);
or U6793 (N_6793,N_2608,N_2626);
nor U6794 (N_6794,N_4387,N_2754);
or U6795 (N_6795,N_2895,N_4053);
nor U6796 (N_6796,N_2751,N_2866);
or U6797 (N_6797,N_3142,N_4897);
and U6798 (N_6798,N_4057,N_2959);
and U6799 (N_6799,N_4715,N_3985);
or U6800 (N_6800,N_4451,N_3549);
nor U6801 (N_6801,N_2977,N_4861);
nor U6802 (N_6802,N_4705,N_4637);
nor U6803 (N_6803,N_4986,N_3570);
nor U6804 (N_6804,N_2612,N_3035);
nand U6805 (N_6805,N_3727,N_3259);
nor U6806 (N_6806,N_4170,N_2710);
nor U6807 (N_6807,N_3100,N_2953);
or U6808 (N_6808,N_4651,N_3815);
and U6809 (N_6809,N_4976,N_4808);
nor U6810 (N_6810,N_4038,N_3176);
nor U6811 (N_6811,N_3824,N_4445);
and U6812 (N_6812,N_4977,N_2910);
and U6813 (N_6813,N_4256,N_4645);
nand U6814 (N_6814,N_4175,N_3343);
or U6815 (N_6815,N_4193,N_3056);
and U6816 (N_6816,N_2923,N_2996);
or U6817 (N_6817,N_3518,N_4251);
and U6818 (N_6818,N_2547,N_2662);
or U6819 (N_6819,N_4814,N_3818);
or U6820 (N_6820,N_4276,N_3376);
or U6821 (N_6821,N_2725,N_4600);
nand U6822 (N_6822,N_4679,N_2961);
or U6823 (N_6823,N_3195,N_2931);
nand U6824 (N_6824,N_3402,N_2534);
or U6825 (N_6825,N_4877,N_4746);
nor U6826 (N_6826,N_4581,N_4997);
nor U6827 (N_6827,N_3493,N_4455);
nor U6828 (N_6828,N_4816,N_4637);
or U6829 (N_6829,N_2669,N_3160);
and U6830 (N_6830,N_3756,N_3711);
nand U6831 (N_6831,N_2635,N_3773);
or U6832 (N_6832,N_4903,N_2963);
or U6833 (N_6833,N_4232,N_4682);
nand U6834 (N_6834,N_3099,N_3912);
or U6835 (N_6835,N_3640,N_4882);
nor U6836 (N_6836,N_3408,N_2506);
or U6837 (N_6837,N_2744,N_4631);
nand U6838 (N_6838,N_4454,N_4167);
nand U6839 (N_6839,N_3230,N_4970);
or U6840 (N_6840,N_3348,N_3164);
nor U6841 (N_6841,N_2523,N_4145);
nor U6842 (N_6842,N_4002,N_4582);
nand U6843 (N_6843,N_2983,N_3594);
nand U6844 (N_6844,N_4016,N_2546);
nand U6845 (N_6845,N_4588,N_3701);
nand U6846 (N_6846,N_4307,N_4202);
and U6847 (N_6847,N_4127,N_2939);
nand U6848 (N_6848,N_3131,N_4488);
nor U6849 (N_6849,N_3501,N_2729);
and U6850 (N_6850,N_4356,N_3921);
nand U6851 (N_6851,N_2641,N_4756);
nand U6852 (N_6852,N_3689,N_4626);
nor U6853 (N_6853,N_2910,N_4922);
nor U6854 (N_6854,N_3522,N_4499);
and U6855 (N_6855,N_3067,N_3225);
nand U6856 (N_6856,N_2939,N_4245);
and U6857 (N_6857,N_3895,N_4295);
or U6858 (N_6858,N_4745,N_3761);
and U6859 (N_6859,N_4283,N_2969);
and U6860 (N_6860,N_4094,N_4824);
nor U6861 (N_6861,N_4079,N_3616);
or U6862 (N_6862,N_4122,N_4709);
nand U6863 (N_6863,N_2622,N_4503);
or U6864 (N_6864,N_4417,N_3417);
and U6865 (N_6865,N_2538,N_4407);
nand U6866 (N_6866,N_3922,N_3448);
xnor U6867 (N_6867,N_2806,N_3394);
nor U6868 (N_6868,N_4665,N_4505);
and U6869 (N_6869,N_3407,N_3072);
nor U6870 (N_6870,N_4067,N_2598);
nand U6871 (N_6871,N_3285,N_4935);
nand U6872 (N_6872,N_2560,N_2840);
nor U6873 (N_6873,N_4384,N_4108);
or U6874 (N_6874,N_2958,N_3708);
nor U6875 (N_6875,N_3916,N_3993);
nor U6876 (N_6876,N_3399,N_3718);
nor U6877 (N_6877,N_3194,N_4437);
nor U6878 (N_6878,N_4052,N_2751);
nand U6879 (N_6879,N_4668,N_4693);
or U6880 (N_6880,N_4538,N_2724);
and U6881 (N_6881,N_4198,N_2845);
nand U6882 (N_6882,N_2993,N_3574);
or U6883 (N_6883,N_3553,N_4082);
and U6884 (N_6884,N_4756,N_3689);
and U6885 (N_6885,N_3982,N_2917);
nand U6886 (N_6886,N_2600,N_3956);
and U6887 (N_6887,N_2984,N_4035);
nor U6888 (N_6888,N_3215,N_3309);
or U6889 (N_6889,N_4713,N_2764);
nor U6890 (N_6890,N_3781,N_3986);
nand U6891 (N_6891,N_3958,N_3047);
and U6892 (N_6892,N_2967,N_4211);
or U6893 (N_6893,N_2531,N_4592);
nand U6894 (N_6894,N_4131,N_2725);
xor U6895 (N_6895,N_2586,N_2728);
and U6896 (N_6896,N_4235,N_2640);
or U6897 (N_6897,N_4054,N_3080);
or U6898 (N_6898,N_4871,N_4804);
nand U6899 (N_6899,N_3380,N_2596);
nor U6900 (N_6900,N_4302,N_4256);
nand U6901 (N_6901,N_2981,N_3615);
xor U6902 (N_6902,N_3615,N_4506);
nand U6903 (N_6903,N_4507,N_3345);
and U6904 (N_6904,N_2685,N_4772);
and U6905 (N_6905,N_3603,N_2941);
nor U6906 (N_6906,N_2597,N_2675);
nand U6907 (N_6907,N_2974,N_2908);
nand U6908 (N_6908,N_3972,N_2717);
nand U6909 (N_6909,N_4554,N_2895);
and U6910 (N_6910,N_3184,N_4527);
xor U6911 (N_6911,N_2682,N_4127);
nand U6912 (N_6912,N_4738,N_4993);
nor U6913 (N_6913,N_2609,N_3229);
or U6914 (N_6914,N_3679,N_4916);
nand U6915 (N_6915,N_2839,N_2520);
nand U6916 (N_6916,N_4210,N_4258);
and U6917 (N_6917,N_4778,N_2828);
or U6918 (N_6918,N_2626,N_3216);
and U6919 (N_6919,N_2522,N_3479);
nor U6920 (N_6920,N_4121,N_3704);
or U6921 (N_6921,N_3107,N_3987);
nand U6922 (N_6922,N_2700,N_3155);
and U6923 (N_6923,N_4986,N_3263);
nor U6924 (N_6924,N_3326,N_4113);
and U6925 (N_6925,N_2598,N_4232);
nor U6926 (N_6926,N_3497,N_3347);
nor U6927 (N_6927,N_3315,N_3492);
and U6928 (N_6928,N_2506,N_4165);
nand U6929 (N_6929,N_4271,N_4567);
nor U6930 (N_6930,N_4755,N_3261);
nand U6931 (N_6931,N_4959,N_2925);
nor U6932 (N_6932,N_4779,N_3033);
nand U6933 (N_6933,N_4682,N_4778);
or U6934 (N_6934,N_2623,N_4766);
or U6935 (N_6935,N_4746,N_3094);
or U6936 (N_6936,N_4819,N_4383);
nand U6937 (N_6937,N_3644,N_2561);
or U6938 (N_6938,N_3115,N_3072);
nor U6939 (N_6939,N_3488,N_3975);
nor U6940 (N_6940,N_4062,N_2728);
nand U6941 (N_6941,N_4213,N_3733);
and U6942 (N_6942,N_3968,N_4754);
and U6943 (N_6943,N_3751,N_4011);
nor U6944 (N_6944,N_2566,N_4705);
or U6945 (N_6945,N_3905,N_3595);
and U6946 (N_6946,N_3315,N_3251);
nor U6947 (N_6947,N_3794,N_4159);
and U6948 (N_6948,N_4112,N_3440);
and U6949 (N_6949,N_3067,N_4288);
nand U6950 (N_6950,N_3400,N_2879);
or U6951 (N_6951,N_4550,N_4128);
nand U6952 (N_6952,N_4564,N_4512);
nor U6953 (N_6953,N_2724,N_4605);
nor U6954 (N_6954,N_4724,N_3870);
nor U6955 (N_6955,N_3291,N_4429);
and U6956 (N_6956,N_3272,N_2720);
nand U6957 (N_6957,N_3771,N_4389);
nor U6958 (N_6958,N_4876,N_3504);
and U6959 (N_6959,N_3409,N_2770);
nor U6960 (N_6960,N_2696,N_4347);
nand U6961 (N_6961,N_3311,N_2958);
nand U6962 (N_6962,N_3771,N_3475);
and U6963 (N_6963,N_4147,N_3688);
xor U6964 (N_6964,N_4433,N_4192);
and U6965 (N_6965,N_4652,N_2850);
or U6966 (N_6966,N_4343,N_3934);
nand U6967 (N_6967,N_3918,N_3478);
nor U6968 (N_6968,N_2911,N_3412);
nor U6969 (N_6969,N_4908,N_2903);
nand U6970 (N_6970,N_2746,N_3945);
nor U6971 (N_6971,N_4769,N_2926);
or U6972 (N_6972,N_4448,N_3905);
and U6973 (N_6973,N_4779,N_3680);
and U6974 (N_6974,N_4364,N_3226);
nor U6975 (N_6975,N_2746,N_3780);
or U6976 (N_6976,N_4402,N_2870);
nand U6977 (N_6977,N_3643,N_3911);
and U6978 (N_6978,N_4826,N_2605);
and U6979 (N_6979,N_3511,N_4942);
or U6980 (N_6980,N_3787,N_3688);
or U6981 (N_6981,N_4562,N_3589);
nand U6982 (N_6982,N_4002,N_4786);
and U6983 (N_6983,N_2519,N_3145);
and U6984 (N_6984,N_3405,N_4495);
and U6985 (N_6985,N_4733,N_2699);
and U6986 (N_6986,N_2548,N_2503);
nor U6987 (N_6987,N_2601,N_4054);
and U6988 (N_6988,N_3175,N_3394);
or U6989 (N_6989,N_4863,N_2877);
nand U6990 (N_6990,N_4615,N_3421);
nand U6991 (N_6991,N_4036,N_3224);
or U6992 (N_6992,N_3981,N_4579);
nor U6993 (N_6993,N_4470,N_3014);
or U6994 (N_6994,N_3350,N_3277);
and U6995 (N_6995,N_3411,N_4911);
or U6996 (N_6996,N_3603,N_3819);
nand U6997 (N_6997,N_4202,N_4982);
or U6998 (N_6998,N_4094,N_3611);
nand U6999 (N_6999,N_4578,N_4520);
nor U7000 (N_7000,N_2826,N_4549);
nor U7001 (N_7001,N_4133,N_4464);
nand U7002 (N_7002,N_3532,N_3765);
nor U7003 (N_7003,N_4472,N_3513);
or U7004 (N_7004,N_3883,N_4885);
nor U7005 (N_7005,N_4320,N_4729);
nand U7006 (N_7006,N_4731,N_4536);
or U7007 (N_7007,N_3168,N_2578);
nor U7008 (N_7008,N_4310,N_4342);
nor U7009 (N_7009,N_4415,N_4162);
and U7010 (N_7010,N_3897,N_4075);
nor U7011 (N_7011,N_2819,N_4142);
and U7012 (N_7012,N_3332,N_2872);
nor U7013 (N_7013,N_4339,N_3754);
or U7014 (N_7014,N_4177,N_4943);
and U7015 (N_7015,N_3341,N_3998);
xnor U7016 (N_7016,N_3522,N_2708);
nor U7017 (N_7017,N_4837,N_4670);
or U7018 (N_7018,N_3425,N_3320);
and U7019 (N_7019,N_4109,N_4488);
nor U7020 (N_7020,N_2818,N_3099);
or U7021 (N_7021,N_4360,N_3430);
nand U7022 (N_7022,N_3583,N_4125);
nor U7023 (N_7023,N_3267,N_4050);
nor U7024 (N_7024,N_4522,N_4515);
or U7025 (N_7025,N_4258,N_4266);
or U7026 (N_7026,N_4401,N_3579);
nor U7027 (N_7027,N_3743,N_4789);
and U7028 (N_7028,N_2889,N_2677);
and U7029 (N_7029,N_3925,N_3994);
and U7030 (N_7030,N_3987,N_4372);
or U7031 (N_7031,N_4924,N_3924);
and U7032 (N_7032,N_4031,N_3690);
nand U7033 (N_7033,N_2518,N_2788);
nor U7034 (N_7034,N_4057,N_3429);
or U7035 (N_7035,N_4127,N_4143);
nand U7036 (N_7036,N_3041,N_2808);
or U7037 (N_7037,N_3993,N_4997);
nand U7038 (N_7038,N_4825,N_2502);
nand U7039 (N_7039,N_4294,N_4125);
nand U7040 (N_7040,N_4954,N_3369);
and U7041 (N_7041,N_3548,N_3943);
or U7042 (N_7042,N_4229,N_4334);
nor U7043 (N_7043,N_4706,N_4328);
or U7044 (N_7044,N_3637,N_4052);
nand U7045 (N_7045,N_4055,N_4924);
and U7046 (N_7046,N_4766,N_3604);
or U7047 (N_7047,N_3375,N_2665);
xnor U7048 (N_7048,N_2506,N_3283);
nand U7049 (N_7049,N_4217,N_3792);
nor U7050 (N_7050,N_3270,N_4924);
nor U7051 (N_7051,N_4548,N_2612);
and U7052 (N_7052,N_2669,N_4584);
or U7053 (N_7053,N_4231,N_3490);
and U7054 (N_7054,N_4663,N_3496);
or U7055 (N_7055,N_3438,N_3583);
or U7056 (N_7056,N_4329,N_3538);
nand U7057 (N_7057,N_4951,N_4629);
or U7058 (N_7058,N_4377,N_4185);
and U7059 (N_7059,N_3697,N_3250);
xnor U7060 (N_7060,N_4206,N_4963);
and U7061 (N_7061,N_3043,N_3388);
nor U7062 (N_7062,N_3362,N_2835);
nor U7063 (N_7063,N_4403,N_4617);
or U7064 (N_7064,N_4942,N_3699);
or U7065 (N_7065,N_3229,N_3935);
nor U7066 (N_7066,N_3191,N_4771);
nand U7067 (N_7067,N_3952,N_4760);
nand U7068 (N_7068,N_3597,N_3815);
and U7069 (N_7069,N_3440,N_3213);
and U7070 (N_7070,N_3486,N_3347);
and U7071 (N_7071,N_3177,N_4248);
nand U7072 (N_7072,N_3051,N_4122);
or U7073 (N_7073,N_3987,N_4787);
nand U7074 (N_7074,N_2923,N_4831);
xor U7075 (N_7075,N_2685,N_3646);
and U7076 (N_7076,N_4126,N_4093);
nand U7077 (N_7077,N_3846,N_4371);
and U7078 (N_7078,N_4628,N_3628);
and U7079 (N_7079,N_3152,N_3410);
or U7080 (N_7080,N_3476,N_3601);
or U7081 (N_7081,N_3658,N_3574);
nor U7082 (N_7082,N_3022,N_3645);
nor U7083 (N_7083,N_3230,N_3518);
and U7084 (N_7084,N_4899,N_4193);
nand U7085 (N_7085,N_2811,N_4468);
nor U7086 (N_7086,N_3681,N_3743);
nand U7087 (N_7087,N_2565,N_3669);
nand U7088 (N_7088,N_3807,N_2902);
or U7089 (N_7089,N_2905,N_3839);
or U7090 (N_7090,N_4689,N_4597);
nor U7091 (N_7091,N_3244,N_3342);
nor U7092 (N_7092,N_4231,N_4472);
and U7093 (N_7093,N_4626,N_2950);
nor U7094 (N_7094,N_3395,N_2719);
and U7095 (N_7095,N_2873,N_4221);
and U7096 (N_7096,N_3269,N_2517);
nand U7097 (N_7097,N_3909,N_2537);
or U7098 (N_7098,N_4942,N_4445);
nand U7099 (N_7099,N_3052,N_3979);
nand U7100 (N_7100,N_4638,N_4905);
nand U7101 (N_7101,N_3018,N_4374);
and U7102 (N_7102,N_4289,N_2879);
and U7103 (N_7103,N_2664,N_4257);
and U7104 (N_7104,N_4816,N_4165);
and U7105 (N_7105,N_3482,N_3780);
or U7106 (N_7106,N_4663,N_4060);
or U7107 (N_7107,N_4107,N_3266);
nor U7108 (N_7108,N_3971,N_4983);
nand U7109 (N_7109,N_4000,N_3243);
xor U7110 (N_7110,N_4450,N_3078);
xnor U7111 (N_7111,N_2752,N_3585);
xnor U7112 (N_7112,N_3136,N_2731);
nor U7113 (N_7113,N_4608,N_3267);
nor U7114 (N_7114,N_4783,N_4546);
nor U7115 (N_7115,N_4601,N_3250);
or U7116 (N_7116,N_2884,N_3361);
or U7117 (N_7117,N_4033,N_4624);
nor U7118 (N_7118,N_3262,N_4974);
nor U7119 (N_7119,N_4468,N_4173);
and U7120 (N_7120,N_2668,N_3937);
or U7121 (N_7121,N_4562,N_4001);
nand U7122 (N_7122,N_3672,N_3708);
nand U7123 (N_7123,N_3969,N_3158);
xnor U7124 (N_7124,N_2930,N_3927);
nand U7125 (N_7125,N_2841,N_3086);
and U7126 (N_7126,N_3624,N_2551);
nor U7127 (N_7127,N_4530,N_4734);
nor U7128 (N_7128,N_4048,N_4950);
and U7129 (N_7129,N_4146,N_4857);
and U7130 (N_7130,N_3980,N_3979);
and U7131 (N_7131,N_2763,N_4000);
nor U7132 (N_7132,N_2570,N_3155);
and U7133 (N_7133,N_3041,N_4001);
or U7134 (N_7134,N_2675,N_4736);
and U7135 (N_7135,N_3338,N_4149);
or U7136 (N_7136,N_3824,N_3163);
nor U7137 (N_7137,N_2716,N_4420);
and U7138 (N_7138,N_4399,N_2591);
nor U7139 (N_7139,N_3420,N_3769);
and U7140 (N_7140,N_3404,N_3468);
nor U7141 (N_7141,N_4570,N_4384);
or U7142 (N_7142,N_4145,N_3541);
and U7143 (N_7143,N_4144,N_3488);
and U7144 (N_7144,N_3414,N_2885);
and U7145 (N_7145,N_2560,N_4897);
nand U7146 (N_7146,N_4574,N_4251);
and U7147 (N_7147,N_3082,N_3565);
nand U7148 (N_7148,N_3953,N_3763);
and U7149 (N_7149,N_4622,N_4012);
or U7150 (N_7150,N_3135,N_2769);
nor U7151 (N_7151,N_3529,N_4070);
or U7152 (N_7152,N_2640,N_4669);
nand U7153 (N_7153,N_3142,N_3108);
xnor U7154 (N_7154,N_4814,N_2953);
and U7155 (N_7155,N_4845,N_4969);
and U7156 (N_7156,N_4651,N_4622);
or U7157 (N_7157,N_4139,N_4817);
and U7158 (N_7158,N_2669,N_2748);
and U7159 (N_7159,N_3404,N_4579);
or U7160 (N_7160,N_3147,N_4602);
nor U7161 (N_7161,N_4530,N_4009);
and U7162 (N_7162,N_3031,N_3225);
nor U7163 (N_7163,N_3147,N_4771);
nand U7164 (N_7164,N_4878,N_2576);
and U7165 (N_7165,N_4481,N_4610);
xnor U7166 (N_7166,N_4055,N_3517);
nand U7167 (N_7167,N_3537,N_2918);
and U7168 (N_7168,N_4419,N_4477);
nor U7169 (N_7169,N_3886,N_2770);
or U7170 (N_7170,N_3584,N_4070);
and U7171 (N_7171,N_2906,N_2666);
nand U7172 (N_7172,N_3643,N_4087);
or U7173 (N_7173,N_4877,N_4119);
nand U7174 (N_7174,N_4586,N_3771);
or U7175 (N_7175,N_4582,N_3355);
nand U7176 (N_7176,N_4690,N_4197);
and U7177 (N_7177,N_3307,N_3770);
and U7178 (N_7178,N_2640,N_4563);
or U7179 (N_7179,N_4034,N_4851);
or U7180 (N_7180,N_2938,N_4662);
or U7181 (N_7181,N_3451,N_4141);
and U7182 (N_7182,N_4029,N_3622);
xor U7183 (N_7183,N_4837,N_3668);
and U7184 (N_7184,N_4236,N_3103);
nor U7185 (N_7185,N_4400,N_4744);
or U7186 (N_7186,N_4485,N_4691);
nor U7187 (N_7187,N_3969,N_4874);
and U7188 (N_7188,N_3348,N_3249);
nand U7189 (N_7189,N_2975,N_2632);
nor U7190 (N_7190,N_3538,N_3636);
or U7191 (N_7191,N_3118,N_4055);
xor U7192 (N_7192,N_3981,N_4637);
nor U7193 (N_7193,N_4889,N_3182);
nor U7194 (N_7194,N_4693,N_4375);
nor U7195 (N_7195,N_4108,N_4240);
nand U7196 (N_7196,N_3232,N_2632);
or U7197 (N_7197,N_4562,N_2519);
nand U7198 (N_7198,N_4866,N_3300);
and U7199 (N_7199,N_3393,N_3095);
and U7200 (N_7200,N_4175,N_3165);
nor U7201 (N_7201,N_4985,N_4567);
nor U7202 (N_7202,N_2906,N_2994);
nand U7203 (N_7203,N_4438,N_4598);
or U7204 (N_7204,N_4640,N_3630);
nor U7205 (N_7205,N_2939,N_2570);
nor U7206 (N_7206,N_3707,N_3224);
and U7207 (N_7207,N_4805,N_3819);
nand U7208 (N_7208,N_3553,N_2739);
and U7209 (N_7209,N_4099,N_3690);
or U7210 (N_7210,N_2899,N_4409);
or U7211 (N_7211,N_3631,N_3032);
nor U7212 (N_7212,N_4545,N_2510);
nand U7213 (N_7213,N_4917,N_4811);
and U7214 (N_7214,N_4900,N_2811);
and U7215 (N_7215,N_4841,N_3121);
xor U7216 (N_7216,N_4162,N_2799);
xor U7217 (N_7217,N_2941,N_2638);
nor U7218 (N_7218,N_4296,N_2569);
nand U7219 (N_7219,N_3760,N_4322);
nor U7220 (N_7220,N_4114,N_2712);
nor U7221 (N_7221,N_3994,N_3571);
and U7222 (N_7222,N_3202,N_4477);
or U7223 (N_7223,N_2786,N_2899);
nor U7224 (N_7224,N_2585,N_2804);
nor U7225 (N_7225,N_2578,N_3120);
and U7226 (N_7226,N_4181,N_2935);
and U7227 (N_7227,N_3685,N_4642);
nand U7228 (N_7228,N_4653,N_4401);
nand U7229 (N_7229,N_2790,N_3095);
nor U7230 (N_7230,N_3682,N_3644);
nand U7231 (N_7231,N_3303,N_4943);
or U7232 (N_7232,N_3433,N_4711);
or U7233 (N_7233,N_3008,N_4177);
and U7234 (N_7234,N_4883,N_2872);
or U7235 (N_7235,N_3486,N_3500);
and U7236 (N_7236,N_4182,N_4513);
or U7237 (N_7237,N_3719,N_3215);
or U7238 (N_7238,N_3074,N_3067);
or U7239 (N_7239,N_4758,N_4421);
or U7240 (N_7240,N_3404,N_3198);
or U7241 (N_7241,N_2725,N_4134);
or U7242 (N_7242,N_4442,N_3205);
xnor U7243 (N_7243,N_4790,N_3477);
and U7244 (N_7244,N_3739,N_3090);
or U7245 (N_7245,N_4748,N_3153);
nand U7246 (N_7246,N_2793,N_3628);
nor U7247 (N_7247,N_4917,N_3526);
or U7248 (N_7248,N_3521,N_4279);
and U7249 (N_7249,N_3873,N_2817);
or U7250 (N_7250,N_2681,N_3968);
or U7251 (N_7251,N_3562,N_4506);
or U7252 (N_7252,N_4546,N_4753);
and U7253 (N_7253,N_3023,N_3517);
nand U7254 (N_7254,N_4040,N_4161);
nor U7255 (N_7255,N_4386,N_2960);
nand U7256 (N_7256,N_3254,N_4169);
and U7257 (N_7257,N_4772,N_4071);
or U7258 (N_7258,N_3479,N_3853);
or U7259 (N_7259,N_4411,N_4869);
or U7260 (N_7260,N_4734,N_3133);
nand U7261 (N_7261,N_3007,N_3326);
and U7262 (N_7262,N_3801,N_3418);
nand U7263 (N_7263,N_3302,N_3211);
or U7264 (N_7264,N_4803,N_3064);
nor U7265 (N_7265,N_3938,N_3191);
nand U7266 (N_7266,N_4722,N_2969);
nand U7267 (N_7267,N_4682,N_4295);
nor U7268 (N_7268,N_2972,N_2796);
nor U7269 (N_7269,N_4565,N_2970);
and U7270 (N_7270,N_2539,N_4522);
nor U7271 (N_7271,N_4823,N_3922);
and U7272 (N_7272,N_4760,N_2593);
and U7273 (N_7273,N_4385,N_3119);
or U7274 (N_7274,N_4402,N_4880);
nand U7275 (N_7275,N_3093,N_2573);
nand U7276 (N_7276,N_4281,N_3280);
nor U7277 (N_7277,N_4963,N_2934);
and U7278 (N_7278,N_4558,N_3843);
nor U7279 (N_7279,N_3012,N_3546);
nand U7280 (N_7280,N_4114,N_3552);
nor U7281 (N_7281,N_3735,N_2954);
xnor U7282 (N_7282,N_2978,N_3627);
and U7283 (N_7283,N_4410,N_4570);
and U7284 (N_7284,N_3758,N_2843);
or U7285 (N_7285,N_2620,N_4882);
or U7286 (N_7286,N_4448,N_3356);
nor U7287 (N_7287,N_4635,N_4243);
and U7288 (N_7288,N_3281,N_4539);
or U7289 (N_7289,N_3466,N_3639);
nand U7290 (N_7290,N_3425,N_4937);
and U7291 (N_7291,N_3634,N_4137);
nor U7292 (N_7292,N_3096,N_4154);
nand U7293 (N_7293,N_4206,N_3354);
and U7294 (N_7294,N_3890,N_3262);
nor U7295 (N_7295,N_4155,N_4504);
and U7296 (N_7296,N_3279,N_4444);
nand U7297 (N_7297,N_3144,N_3500);
and U7298 (N_7298,N_3204,N_2792);
nand U7299 (N_7299,N_3506,N_4865);
or U7300 (N_7300,N_4905,N_2785);
nand U7301 (N_7301,N_3348,N_2867);
nor U7302 (N_7302,N_4823,N_3899);
and U7303 (N_7303,N_4918,N_4175);
nand U7304 (N_7304,N_3833,N_4428);
or U7305 (N_7305,N_4784,N_3682);
nand U7306 (N_7306,N_3376,N_2577);
nor U7307 (N_7307,N_4176,N_4429);
nand U7308 (N_7308,N_3423,N_2547);
and U7309 (N_7309,N_3637,N_4496);
and U7310 (N_7310,N_3381,N_3391);
nand U7311 (N_7311,N_3316,N_4370);
and U7312 (N_7312,N_4386,N_3788);
and U7313 (N_7313,N_4124,N_3834);
or U7314 (N_7314,N_2738,N_4028);
nor U7315 (N_7315,N_4843,N_3478);
nor U7316 (N_7316,N_2856,N_3586);
and U7317 (N_7317,N_4728,N_3696);
and U7318 (N_7318,N_2736,N_3744);
nor U7319 (N_7319,N_3268,N_4692);
and U7320 (N_7320,N_4991,N_3053);
or U7321 (N_7321,N_4502,N_4932);
and U7322 (N_7322,N_3396,N_3816);
nor U7323 (N_7323,N_3281,N_4700);
nand U7324 (N_7324,N_3962,N_3572);
nor U7325 (N_7325,N_3501,N_4888);
and U7326 (N_7326,N_3406,N_3177);
or U7327 (N_7327,N_4617,N_4847);
nor U7328 (N_7328,N_3163,N_4980);
or U7329 (N_7329,N_3816,N_3040);
and U7330 (N_7330,N_4319,N_3052);
nor U7331 (N_7331,N_2660,N_3702);
and U7332 (N_7332,N_2798,N_3476);
and U7333 (N_7333,N_4212,N_3170);
nand U7334 (N_7334,N_2683,N_4292);
nand U7335 (N_7335,N_4493,N_3748);
and U7336 (N_7336,N_3848,N_2507);
nor U7337 (N_7337,N_3099,N_4466);
and U7338 (N_7338,N_4722,N_2504);
and U7339 (N_7339,N_4546,N_3557);
nand U7340 (N_7340,N_2757,N_4539);
or U7341 (N_7341,N_4628,N_3234);
or U7342 (N_7342,N_3199,N_2960);
or U7343 (N_7343,N_2782,N_4488);
and U7344 (N_7344,N_3753,N_2817);
nor U7345 (N_7345,N_3773,N_4480);
xnor U7346 (N_7346,N_3953,N_2904);
or U7347 (N_7347,N_3911,N_4266);
or U7348 (N_7348,N_2827,N_4017);
or U7349 (N_7349,N_2825,N_2857);
nand U7350 (N_7350,N_3214,N_3062);
xor U7351 (N_7351,N_3844,N_4005);
or U7352 (N_7352,N_4106,N_2937);
nor U7353 (N_7353,N_2562,N_4024);
nand U7354 (N_7354,N_4846,N_2505);
nor U7355 (N_7355,N_4088,N_4276);
nand U7356 (N_7356,N_4971,N_3716);
nor U7357 (N_7357,N_4240,N_4720);
nor U7358 (N_7358,N_3845,N_4936);
or U7359 (N_7359,N_3830,N_2797);
nand U7360 (N_7360,N_3525,N_3111);
nand U7361 (N_7361,N_4859,N_3952);
or U7362 (N_7362,N_3622,N_3229);
nand U7363 (N_7363,N_4858,N_2578);
or U7364 (N_7364,N_4202,N_2573);
nand U7365 (N_7365,N_3626,N_2659);
and U7366 (N_7366,N_4875,N_4189);
or U7367 (N_7367,N_4471,N_3437);
nand U7368 (N_7368,N_4573,N_3849);
nor U7369 (N_7369,N_3221,N_2717);
and U7370 (N_7370,N_4743,N_3468);
nor U7371 (N_7371,N_3244,N_3812);
and U7372 (N_7372,N_4244,N_3211);
or U7373 (N_7373,N_2617,N_2583);
and U7374 (N_7374,N_3668,N_3634);
and U7375 (N_7375,N_3409,N_3191);
or U7376 (N_7376,N_4438,N_4541);
and U7377 (N_7377,N_4829,N_3244);
nor U7378 (N_7378,N_3030,N_4799);
xor U7379 (N_7379,N_3245,N_4204);
and U7380 (N_7380,N_4458,N_3565);
or U7381 (N_7381,N_4916,N_4534);
and U7382 (N_7382,N_4366,N_3716);
nand U7383 (N_7383,N_2635,N_2573);
and U7384 (N_7384,N_3156,N_2666);
nor U7385 (N_7385,N_2962,N_3752);
nor U7386 (N_7386,N_4370,N_3993);
and U7387 (N_7387,N_2925,N_3217);
or U7388 (N_7388,N_4262,N_3288);
nor U7389 (N_7389,N_4274,N_3363);
or U7390 (N_7390,N_4614,N_3516);
and U7391 (N_7391,N_3031,N_3756);
nand U7392 (N_7392,N_4686,N_3698);
nor U7393 (N_7393,N_3895,N_2992);
nand U7394 (N_7394,N_2613,N_3196);
or U7395 (N_7395,N_2690,N_2920);
and U7396 (N_7396,N_2618,N_4382);
and U7397 (N_7397,N_2631,N_4816);
or U7398 (N_7398,N_3538,N_4746);
nor U7399 (N_7399,N_3043,N_4266);
nor U7400 (N_7400,N_3879,N_3232);
nand U7401 (N_7401,N_3681,N_2986);
nand U7402 (N_7402,N_2579,N_4953);
or U7403 (N_7403,N_4151,N_3603);
nand U7404 (N_7404,N_3747,N_3926);
or U7405 (N_7405,N_3846,N_4512);
and U7406 (N_7406,N_3487,N_3210);
or U7407 (N_7407,N_3803,N_3199);
nand U7408 (N_7408,N_3776,N_2983);
nand U7409 (N_7409,N_4101,N_3231);
or U7410 (N_7410,N_4321,N_3572);
nand U7411 (N_7411,N_4576,N_3362);
nor U7412 (N_7412,N_4805,N_4085);
and U7413 (N_7413,N_4992,N_4445);
or U7414 (N_7414,N_4731,N_4076);
or U7415 (N_7415,N_3462,N_3698);
or U7416 (N_7416,N_4655,N_4093);
xor U7417 (N_7417,N_4230,N_3882);
nor U7418 (N_7418,N_2980,N_2971);
and U7419 (N_7419,N_2671,N_3128);
or U7420 (N_7420,N_4585,N_2730);
nand U7421 (N_7421,N_4824,N_4234);
nor U7422 (N_7422,N_3542,N_3813);
nor U7423 (N_7423,N_2520,N_3114);
nor U7424 (N_7424,N_3327,N_4999);
xor U7425 (N_7425,N_3968,N_4815);
and U7426 (N_7426,N_2549,N_2779);
and U7427 (N_7427,N_3999,N_3207);
nand U7428 (N_7428,N_4016,N_4298);
nor U7429 (N_7429,N_3262,N_2993);
nand U7430 (N_7430,N_2839,N_4784);
nand U7431 (N_7431,N_3347,N_4667);
or U7432 (N_7432,N_4865,N_2718);
or U7433 (N_7433,N_2614,N_3673);
or U7434 (N_7434,N_2979,N_4782);
and U7435 (N_7435,N_4509,N_2672);
nor U7436 (N_7436,N_4683,N_3034);
or U7437 (N_7437,N_3701,N_4637);
and U7438 (N_7438,N_3887,N_4312);
and U7439 (N_7439,N_3340,N_4452);
and U7440 (N_7440,N_4271,N_3091);
nor U7441 (N_7441,N_4233,N_3861);
nor U7442 (N_7442,N_4090,N_2502);
nor U7443 (N_7443,N_4280,N_4855);
nand U7444 (N_7444,N_4123,N_2517);
or U7445 (N_7445,N_4382,N_2631);
nand U7446 (N_7446,N_2962,N_2543);
nand U7447 (N_7447,N_4063,N_2707);
or U7448 (N_7448,N_3910,N_4253);
nand U7449 (N_7449,N_4677,N_4513);
nand U7450 (N_7450,N_2604,N_4265);
and U7451 (N_7451,N_4371,N_3610);
nor U7452 (N_7452,N_4294,N_3972);
nand U7453 (N_7453,N_3097,N_3104);
nand U7454 (N_7454,N_4643,N_3554);
nor U7455 (N_7455,N_3274,N_4667);
or U7456 (N_7456,N_2711,N_3570);
xor U7457 (N_7457,N_2843,N_4817);
nor U7458 (N_7458,N_2855,N_3357);
nand U7459 (N_7459,N_3273,N_3126);
and U7460 (N_7460,N_2960,N_4184);
or U7461 (N_7461,N_2773,N_4733);
nor U7462 (N_7462,N_4556,N_4309);
nand U7463 (N_7463,N_2815,N_3796);
or U7464 (N_7464,N_4608,N_4127);
or U7465 (N_7465,N_3658,N_3576);
nand U7466 (N_7466,N_4028,N_4680);
nand U7467 (N_7467,N_3617,N_3721);
nand U7468 (N_7468,N_2883,N_4376);
and U7469 (N_7469,N_3736,N_3115);
or U7470 (N_7470,N_4966,N_3049);
nor U7471 (N_7471,N_2662,N_4261);
xnor U7472 (N_7472,N_2623,N_3225);
or U7473 (N_7473,N_2845,N_3944);
nand U7474 (N_7474,N_3740,N_3975);
nand U7475 (N_7475,N_4886,N_3128);
nand U7476 (N_7476,N_2980,N_3460);
and U7477 (N_7477,N_2756,N_3643);
nand U7478 (N_7478,N_3383,N_3456);
nand U7479 (N_7479,N_4897,N_2538);
nor U7480 (N_7480,N_4662,N_4425);
and U7481 (N_7481,N_4674,N_3961);
nor U7482 (N_7482,N_4995,N_4884);
or U7483 (N_7483,N_4263,N_3855);
nor U7484 (N_7484,N_3381,N_4870);
or U7485 (N_7485,N_4408,N_3451);
nand U7486 (N_7486,N_4036,N_4120);
nor U7487 (N_7487,N_3398,N_3282);
nand U7488 (N_7488,N_3141,N_4946);
nor U7489 (N_7489,N_3197,N_4404);
or U7490 (N_7490,N_4548,N_3044);
and U7491 (N_7491,N_3046,N_2678);
nand U7492 (N_7492,N_3550,N_2897);
and U7493 (N_7493,N_3526,N_4670);
and U7494 (N_7494,N_3972,N_2614);
and U7495 (N_7495,N_3251,N_3547);
nor U7496 (N_7496,N_2664,N_3341);
and U7497 (N_7497,N_4856,N_3554);
nor U7498 (N_7498,N_4250,N_2534);
or U7499 (N_7499,N_4731,N_3041);
and U7500 (N_7500,N_5386,N_5942);
nor U7501 (N_7501,N_5605,N_5065);
and U7502 (N_7502,N_5253,N_7021);
nand U7503 (N_7503,N_6368,N_5374);
nor U7504 (N_7504,N_6819,N_7215);
nand U7505 (N_7505,N_6832,N_5892);
nor U7506 (N_7506,N_6130,N_7230);
nor U7507 (N_7507,N_7101,N_6144);
nand U7508 (N_7508,N_6867,N_6806);
nand U7509 (N_7509,N_6479,N_6741);
nor U7510 (N_7510,N_6054,N_6831);
nor U7511 (N_7511,N_7104,N_5122);
nor U7512 (N_7512,N_7367,N_5393);
nor U7513 (N_7513,N_5720,N_7190);
xnor U7514 (N_7514,N_6138,N_6692);
nor U7515 (N_7515,N_7071,N_6122);
and U7516 (N_7516,N_6030,N_5927);
nor U7517 (N_7517,N_5263,N_5724);
and U7518 (N_7518,N_7066,N_5516);
or U7519 (N_7519,N_6757,N_7084);
or U7520 (N_7520,N_5482,N_6855);
nand U7521 (N_7521,N_5604,N_5014);
and U7522 (N_7522,N_7034,N_6481);
nand U7523 (N_7523,N_5112,N_7060);
or U7524 (N_7524,N_5385,N_6955);
and U7525 (N_7525,N_5662,N_6927);
nor U7526 (N_7526,N_5049,N_7002);
nor U7527 (N_7527,N_6857,N_5952);
nand U7528 (N_7528,N_5555,N_5660);
nor U7529 (N_7529,N_5856,N_5025);
nand U7530 (N_7530,N_6794,N_5843);
or U7531 (N_7531,N_5209,N_6235);
xor U7532 (N_7532,N_6667,N_5291);
or U7533 (N_7533,N_5827,N_5855);
nand U7534 (N_7534,N_7323,N_6502);
and U7535 (N_7535,N_6427,N_5506);
and U7536 (N_7536,N_7380,N_6319);
nor U7537 (N_7537,N_6388,N_7290);
and U7538 (N_7538,N_6615,N_6928);
or U7539 (N_7539,N_5747,N_5916);
or U7540 (N_7540,N_7417,N_6082);
nor U7541 (N_7541,N_5896,N_7177);
and U7542 (N_7542,N_6643,N_5858);
and U7543 (N_7543,N_7315,N_5676);
or U7544 (N_7544,N_6554,N_6820);
xnor U7545 (N_7545,N_7109,N_6445);
or U7546 (N_7546,N_6317,N_5473);
and U7547 (N_7547,N_6715,N_5093);
or U7548 (N_7548,N_6576,N_6705);
and U7549 (N_7549,N_6188,N_7379);
and U7550 (N_7550,N_5109,N_7468);
nand U7551 (N_7551,N_6733,N_6258);
and U7552 (N_7552,N_5568,N_5762);
and U7553 (N_7553,N_6273,N_6934);
or U7554 (N_7554,N_5459,N_7339);
nor U7555 (N_7555,N_6509,N_7309);
nor U7556 (N_7556,N_5074,N_5594);
nor U7557 (N_7557,N_5941,N_6204);
nor U7558 (N_7558,N_7075,N_5307);
or U7559 (N_7559,N_5343,N_5082);
and U7560 (N_7560,N_6147,N_5134);
nand U7561 (N_7561,N_5123,N_6395);
nand U7562 (N_7562,N_5749,N_6918);
or U7563 (N_7563,N_7486,N_6069);
or U7564 (N_7564,N_5174,N_5582);
or U7565 (N_7565,N_6078,N_5371);
nor U7566 (N_7566,N_6354,N_5641);
nand U7567 (N_7567,N_5384,N_5237);
or U7568 (N_7568,N_5692,N_5854);
or U7569 (N_7569,N_6942,N_6558);
nand U7570 (N_7570,N_7059,N_5187);
nand U7571 (N_7571,N_5153,N_5330);
nor U7572 (N_7572,N_6662,N_5850);
nor U7573 (N_7573,N_6250,N_5729);
nor U7574 (N_7574,N_5390,N_7457);
or U7575 (N_7575,N_6207,N_6193);
nor U7576 (N_7576,N_6598,N_7181);
or U7577 (N_7577,N_6646,N_6364);
nand U7578 (N_7578,N_6683,N_7436);
and U7579 (N_7579,N_6039,N_7319);
nand U7580 (N_7580,N_6212,N_7204);
and U7581 (N_7581,N_5005,N_5230);
nor U7582 (N_7582,N_5813,N_5550);
and U7583 (N_7583,N_5966,N_5759);
and U7584 (N_7584,N_5267,N_6062);
or U7585 (N_7585,N_6665,N_5133);
nand U7586 (N_7586,N_6717,N_6604);
or U7587 (N_7587,N_6448,N_6392);
nor U7588 (N_7588,N_6756,N_5935);
nand U7589 (N_7589,N_7439,N_5932);
or U7590 (N_7590,N_6600,N_6327);
nand U7591 (N_7591,N_6626,N_6792);
and U7592 (N_7592,N_5549,N_5987);
and U7593 (N_7593,N_7119,N_5336);
xor U7594 (N_7594,N_5258,N_5271);
or U7595 (N_7595,N_5541,N_5751);
nand U7596 (N_7596,N_5592,N_6522);
or U7597 (N_7597,N_5272,N_6027);
and U7598 (N_7598,N_5488,N_6902);
nor U7599 (N_7599,N_6861,N_5113);
nand U7600 (N_7600,N_5306,N_5644);
nor U7601 (N_7601,N_7283,N_5965);
nand U7602 (N_7602,N_6377,N_7227);
and U7603 (N_7603,N_6999,N_6883);
nand U7604 (N_7604,N_6888,N_5106);
or U7605 (N_7605,N_5764,N_5163);
or U7606 (N_7606,N_7316,N_5578);
xor U7607 (N_7607,N_6812,N_6483);
or U7608 (N_7608,N_5763,N_6609);
nand U7609 (N_7609,N_6386,N_5453);
nor U7610 (N_7610,N_7078,N_5557);
or U7611 (N_7611,N_5417,N_5790);
and U7612 (N_7612,N_6680,N_7171);
and U7613 (N_7613,N_7240,N_5047);
nand U7614 (N_7614,N_5733,N_6492);
nand U7615 (N_7615,N_7001,N_5873);
nand U7616 (N_7616,N_6149,N_5494);
nand U7617 (N_7617,N_7278,N_6310);
nor U7618 (N_7618,N_6898,N_7173);
nor U7619 (N_7619,N_5536,N_6910);
nor U7620 (N_7620,N_5670,N_5580);
nand U7621 (N_7621,N_7079,N_6749);
nor U7622 (N_7622,N_6220,N_5534);
nor U7623 (N_7623,N_6526,N_5003);
or U7624 (N_7624,N_5125,N_5831);
nor U7625 (N_7625,N_5440,N_6419);
or U7626 (N_7626,N_5444,N_6309);
nand U7627 (N_7627,N_7389,N_6011);
and U7628 (N_7628,N_5829,N_6961);
or U7629 (N_7629,N_6924,N_5428);
and U7630 (N_7630,N_7451,N_5776);
and U7631 (N_7631,N_7462,N_5804);
or U7632 (N_7632,N_6244,N_6067);
nor U7633 (N_7633,N_6729,N_6734);
or U7634 (N_7634,N_5523,N_5658);
nand U7635 (N_7635,N_7282,N_6561);
nor U7636 (N_7636,N_6889,N_5796);
nor U7637 (N_7637,N_6352,N_6628);
nor U7638 (N_7638,N_5333,N_5496);
or U7639 (N_7639,N_6495,N_6557);
xor U7640 (N_7640,N_6029,N_6323);
xnor U7641 (N_7641,N_6892,N_5070);
or U7642 (N_7642,N_5436,N_6346);
nor U7643 (N_7643,N_5566,N_6257);
nor U7644 (N_7644,N_5392,N_6496);
and U7645 (N_7645,N_5197,N_6994);
nor U7646 (N_7646,N_5849,N_5499);
or U7647 (N_7647,N_6172,N_5182);
and U7648 (N_7648,N_7040,N_5632);
and U7649 (N_7649,N_6470,N_6420);
nand U7650 (N_7650,N_6535,N_5475);
and U7651 (N_7651,N_7147,N_5190);
or U7652 (N_7652,N_5063,N_5705);
nand U7653 (N_7653,N_5521,N_7183);
nand U7654 (N_7654,N_6219,N_5840);
and U7655 (N_7655,N_6002,N_6754);
nor U7656 (N_7656,N_6485,N_6666);
or U7657 (N_7657,N_6223,N_7141);
or U7658 (N_7658,N_7428,N_7268);
or U7659 (N_7659,N_5640,N_5503);
nor U7660 (N_7660,N_5379,N_5391);
and U7661 (N_7661,N_6610,N_7005);
or U7662 (N_7662,N_5789,N_5338);
nor U7663 (N_7663,N_6624,N_6896);
nor U7664 (N_7664,N_5205,N_5443);
or U7665 (N_7665,N_6956,N_7284);
nand U7666 (N_7666,N_6539,N_5681);
and U7667 (N_7667,N_6958,N_6949);
nand U7668 (N_7668,N_7242,N_6348);
nand U7669 (N_7669,N_6374,N_5151);
nor U7670 (N_7670,N_6176,N_6232);
or U7671 (N_7671,N_5377,N_5526);
or U7672 (N_7672,N_6043,N_5707);
or U7673 (N_7673,N_5077,N_5527);
nor U7674 (N_7674,N_6866,N_6673);
nor U7675 (N_7675,N_5667,N_7427);
or U7676 (N_7676,N_6467,N_5259);
or U7677 (N_7677,N_7429,N_7238);
and U7678 (N_7678,N_6688,N_6684);
and U7679 (N_7679,N_6096,N_5016);
nor U7680 (N_7680,N_7178,N_5409);
and U7681 (N_7681,N_6822,N_7411);
and U7682 (N_7682,N_7343,N_5609);
and U7683 (N_7683,N_5685,N_5294);
nor U7684 (N_7684,N_5874,N_5738);
and U7685 (N_7685,N_6728,N_5997);
nor U7686 (N_7686,N_6196,N_7351);
and U7687 (N_7687,N_5027,N_5994);
or U7688 (N_7688,N_7218,N_7495);
or U7689 (N_7689,N_7117,N_5906);
or U7690 (N_7690,N_6727,N_6966);
and U7691 (N_7691,N_6974,N_5572);
or U7692 (N_7692,N_5086,N_5465);
nor U7693 (N_7693,N_7294,N_5778);
or U7694 (N_7694,N_7346,N_5522);
nand U7695 (N_7695,N_7364,N_5606);
nor U7696 (N_7696,N_6387,N_6167);
nor U7697 (N_7697,N_5570,N_5815);
nand U7698 (N_7698,N_6530,N_7382);
nand U7699 (N_7699,N_5710,N_6523);
nand U7700 (N_7700,N_5870,N_6917);
and U7701 (N_7701,N_5618,N_6066);
or U7702 (N_7702,N_5899,N_6446);
nor U7703 (N_7703,N_6519,N_7063);
nor U7704 (N_7704,N_7482,N_7026);
nand U7705 (N_7705,N_5629,N_7267);
nor U7706 (N_7706,N_5171,N_5262);
or U7707 (N_7707,N_6511,N_5381);
nor U7708 (N_7708,N_7111,N_5974);
or U7709 (N_7709,N_5576,N_6114);
nor U7710 (N_7710,N_5767,N_6246);
or U7711 (N_7711,N_7031,N_6085);
nand U7712 (N_7712,N_6629,N_6834);
and U7713 (N_7713,N_6976,N_5004);
or U7714 (N_7714,N_6887,N_5655);
and U7715 (N_7715,N_7206,N_6622);
or U7716 (N_7716,N_5007,N_5554);
or U7717 (N_7717,N_6058,N_6660);
xnor U7718 (N_7718,N_6544,N_6120);
and U7719 (N_7719,N_5281,N_5953);
nand U7720 (N_7720,N_5754,N_6764);
nand U7721 (N_7721,N_6647,N_6700);
nand U7722 (N_7722,N_6914,N_7237);
or U7723 (N_7723,N_5525,N_7179);
nor U7724 (N_7724,N_6516,N_5904);
nand U7725 (N_7725,N_5311,N_7122);
and U7726 (N_7726,N_5193,N_5117);
nand U7727 (N_7727,N_5244,N_6126);
and U7728 (N_7728,N_7326,N_5735);
and U7729 (N_7729,N_6788,N_5823);
xnor U7730 (N_7730,N_5455,N_6200);
nand U7731 (N_7731,N_5001,N_5567);
and U7732 (N_7732,N_5400,N_5556);
nand U7733 (N_7733,N_7003,N_5945);
and U7734 (N_7734,N_5663,N_5518);
and U7735 (N_7735,N_6453,N_5860);
nand U7736 (N_7736,N_6159,N_5411);
nand U7737 (N_7737,N_5329,N_6814);
nand U7738 (N_7738,N_6322,N_5220);
and U7739 (N_7739,N_7293,N_5884);
nor U7740 (N_7740,N_6251,N_6150);
nor U7741 (N_7741,N_5347,N_5235);
nor U7742 (N_7742,N_5427,N_6477);
nor U7743 (N_7743,N_5588,N_7055);
nor U7744 (N_7744,N_5889,N_7246);
nor U7745 (N_7745,N_6844,N_5674);
nand U7746 (N_7746,N_6044,N_5806);
nor U7747 (N_7747,N_6846,N_6585);
nand U7748 (N_7748,N_6426,N_5466);
nor U7749 (N_7749,N_5985,N_5880);
nand U7750 (N_7750,N_6803,N_6165);
or U7751 (N_7751,N_6641,N_5183);
nand U7752 (N_7752,N_5430,N_5591);
and U7753 (N_7753,N_7113,N_5888);
or U7754 (N_7754,N_6074,N_5920);
or U7755 (N_7755,N_6407,N_6525);
and U7756 (N_7756,N_5223,N_5625);
nor U7757 (N_7757,N_5717,N_5741);
and U7758 (N_7758,N_5489,N_6294);
and U7759 (N_7759,N_7187,N_6260);
nand U7760 (N_7760,N_7211,N_6638);
and U7761 (N_7761,N_6290,N_5130);
nor U7762 (N_7762,N_6378,N_7488);
and U7763 (N_7763,N_7249,N_6627);
or U7764 (N_7764,N_6022,N_5801);
and U7765 (N_7765,N_6103,N_6802);
nand U7766 (N_7766,N_7160,N_6656);
nor U7767 (N_7767,N_5703,N_6882);
nand U7768 (N_7768,N_5671,N_6451);
nand U7769 (N_7769,N_6972,N_6343);
or U7770 (N_7770,N_6277,N_5178);
or U7771 (N_7771,N_6422,N_7285);
nand U7772 (N_7772,N_7363,N_6156);
nor U7773 (N_7773,N_5711,N_5201);
or U7774 (N_7774,N_7289,N_7329);
nor U7775 (N_7775,N_5479,N_5579);
nor U7776 (N_7776,N_6636,N_6623);
or U7777 (N_7777,N_5161,N_7112);
and U7778 (N_7778,N_6102,N_6381);
and U7779 (N_7779,N_6904,N_5115);
nor U7780 (N_7780,N_6342,N_7466);
nor U7781 (N_7781,N_5288,N_7234);
or U7782 (N_7782,N_6770,N_6115);
or U7783 (N_7783,N_7094,N_6474);
xor U7784 (N_7784,N_6135,N_6036);
nor U7785 (N_7785,N_6498,N_5487);
nor U7786 (N_7786,N_7229,N_5104);
and U7787 (N_7787,N_6650,N_6107);
nor U7788 (N_7788,N_6977,N_6552);
and U7789 (N_7789,N_5470,N_6895);
nor U7790 (N_7790,N_6563,N_7261);
and U7791 (N_7791,N_5124,N_5395);
or U7792 (N_7792,N_6175,N_6051);
or U7793 (N_7793,N_5561,N_5947);
and U7794 (N_7794,N_5697,N_6905);
or U7795 (N_7795,N_5375,N_7394);
and U7796 (N_7796,N_7402,N_5457);
or U7797 (N_7797,N_6166,N_7196);
nor U7798 (N_7798,N_6264,N_6815);
and U7799 (N_7799,N_5114,N_5434);
nand U7800 (N_7800,N_7362,N_6452);
nor U7801 (N_7801,N_6852,N_6210);
nor U7802 (N_7802,N_6296,N_5745);
xor U7803 (N_7803,N_7180,N_6588);
nand U7804 (N_7804,N_5872,N_6383);
and U7805 (N_7805,N_6567,N_6726);
nor U7806 (N_7806,N_6435,N_5492);
or U7807 (N_7807,N_7263,N_6618);
or U7808 (N_7808,N_6291,N_5398);
and U7809 (N_7809,N_6858,N_7375);
nand U7810 (N_7810,N_7009,N_5407);
nor U7811 (N_7811,N_6874,N_5156);
or U7812 (N_7812,N_5540,N_6265);
nor U7813 (N_7813,N_5836,N_6288);
nand U7814 (N_7814,N_6925,N_5689);
and U7815 (N_7815,N_6920,N_5603);
nor U7816 (N_7816,N_6414,N_5647);
and U7817 (N_7817,N_7469,N_5092);
or U7818 (N_7818,N_5295,N_7232);
or U7819 (N_7819,N_7374,N_5486);
and U7820 (N_7820,N_6468,N_5933);
and U7821 (N_7821,N_5563,N_6391);
nand U7822 (N_7822,N_6841,N_6649);
nor U7823 (N_7823,N_6578,N_5073);
nand U7824 (N_7824,N_6347,N_6982);
nand U7825 (N_7825,N_5274,N_6123);
or U7826 (N_7826,N_7200,N_5046);
nand U7827 (N_7827,N_7461,N_5078);
nand U7828 (N_7828,N_5537,N_5925);
nand U7829 (N_7829,N_5367,N_7090);
xor U7830 (N_7830,N_6514,N_7061);
or U7831 (N_7831,N_6004,N_6399);
nand U7832 (N_7832,N_7203,N_5838);
nor U7833 (N_7833,N_7460,N_7483);
nand U7834 (N_7834,N_5943,N_5290);
nand U7835 (N_7835,N_5217,N_6911);
and U7836 (N_7836,N_7220,N_5988);
nor U7837 (N_7837,N_6341,N_6952);
and U7838 (N_7838,N_5844,N_6358);
and U7839 (N_7839,N_6041,N_7129);
nand U7840 (N_7840,N_6878,N_5203);
and U7841 (N_7841,N_7022,N_5296);
nor U7842 (N_7842,N_5520,N_6143);
and U7843 (N_7843,N_5321,N_6686);
or U7844 (N_7844,N_7372,N_6571);
nor U7845 (N_7845,N_7033,N_5902);
nand U7846 (N_7846,N_6935,N_5100);
and U7847 (N_7847,N_5155,N_6055);
nand U7848 (N_7848,N_7091,N_7320);
nand U7849 (N_7849,N_5071,N_5204);
and U7850 (N_7850,N_5481,N_5224);
nand U7851 (N_7851,N_5501,N_5015);
and U7852 (N_7852,N_6682,N_5653);
nor U7853 (N_7853,N_6735,N_6782);
or U7854 (N_7854,N_6304,N_6712);
nand U7855 (N_7855,N_6589,N_7041);
nand U7856 (N_7856,N_6053,N_7485);
or U7857 (N_7857,N_5261,N_6367);
or U7858 (N_7858,N_6139,N_6423);
or U7859 (N_7859,N_7365,N_7214);
or U7860 (N_7860,N_5981,N_5227);
and U7861 (N_7861,N_5613,N_5195);
nor U7862 (N_7862,N_6353,N_7287);
nand U7863 (N_7863,N_5243,N_7455);
nand U7864 (N_7864,N_7395,N_6997);
xor U7865 (N_7865,N_7440,N_5731);
or U7866 (N_7866,N_6384,N_6351);
nor U7867 (N_7867,N_5175,N_5743);
or U7868 (N_7868,N_5539,N_6020);
nor U7869 (N_7869,N_5266,N_5739);
or U7870 (N_7870,N_7192,N_7271);
and U7871 (N_7871,N_7404,N_5062);
nand U7872 (N_7872,N_6325,N_5273);
xor U7873 (N_7873,N_7105,N_5786);
or U7874 (N_7874,N_5999,N_5706);
or U7875 (N_7875,N_5661,N_5146);
nand U7876 (N_7876,N_6625,N_5975);
and U7877 (N_7877,N_6269,N_7303);
and U7878 (N_7878,N_5694,N_7070);
nand U7879 (N_7879,N_5450,N_5158);
and U7880 (N_7880,N_6124,N_6117);
or U7881 (N_7881,N_5478,N_6293);
xnor U7882 (N_7882,N_5010,N_5638);
nand U7883 (N_7883,N_6722,N_5532);
and U7884 (N_7884,N_6213,N_6690);
nand U7885 (N_7885,N_5508,N_7262);
nor U7886 (N_7886,N_6978,N_5043);
xnor U7887 (N_7887,N_6181,N_6940);
and U7888 (N_7888,N_5405,N_7068);
xor U7889 (N_7889,N_6289,N_7370);
nor U7890 (N_7890,N_5748,N_7381);
nor U7891 (N_7891,N_5725,N_5191);
and U7892 (N_7892,N_6695,N_6698);
nor U7893 (N_7893,N_6259,N_5363);
nor U7894 (N_7894,N_6936,N_7023);
nand U7895 (N_7895,N_6602,N_5257);
and U7896 (N_7896,N_6462,N_6410);
or U7897 (N_7897,N_5651,N_5634);
nor U7898 (N_7898,N_6752,N_7472);
nor U7899 (N_7899,N_5126,N_5402);
or U7900 (N_7900,N_6237,N_7304);
nor U7901 (N_7901,N_6416,N_6009);
nor U7902 (N_7902,N_5432,N_5324);
nor U7903 (N_7903,N_5437,N_7291);
nand U7904 (N_7904,N_5924,N_7277);
and U7905 (N_7905,N_6573,N_5959);
nor U7906 (N_7906,N_5898,N_7130);
or U7907 (N_7907,N_6340,N_6789);
and U7908 (N_7908,N_5538,N_6872);
nand U7909 (N_7909,N_5067,N_7473);
or U7910 (N_7910,N_6026,N_5657);
nor U7911 (N_7911,N_7449,N_6829);
nand U7912 (N_7912,N_5373,N_5420);
nand U7913 (N_7913,N_6438,N_5853);
nand U7914 (N_7914,N_5793,N_5809);
nand U7915 (N_7915,N_5037,N_7115);
and U7916 (N_7916,N_6891,N_7114);
or U7917 (N_7917,N_6086,N_6371);
nor U7918 (N_7918,N_7347,N_5814);
or U7919 (N_7919,N_6405,N_6357);
nand U7920 (N_7920,N_6981,N_5602);
nor U7921 (N_7921,N_6548,N_6517);
nor U7922 (N_7922,N_5326,N_7341);
nand U7923 (N_7923,N_5977,N_6187);
and U7924 (N_7924,N_6033,N_5246);
nor U7925 (N_7925,N_7244,N_7385);
nand U7926 (N_7926,N_5847,N_5700);
and U7927 (N_7927,N_5654,N_6651);
or U7928 (N_7928,N_6654,N_5008);
or U7929 (N_7929,N_5510,N_5505);
nor U7930 (N_7930,N_6224,N_7138);
xor U7931 (N_7931,N_6710,N_6580);
or U7932 (N_7932,N_6531,N_5646);
xnor U7933 (N_7933,N_7313,N_7366);
and U7934 (N_7934,N_6818,N_6180);
or U7935 (N_7935,N_6308,N_5963);
or U7936 (N_7936,N_7074,N_5919);
nor U7937 (N_7937,N_5552,N_5728);
nor U7938 (N_7938,N_5967,N_6694);
and U7939 (N_7939,N_5573,N_6214);
or U7940 (N_7940,N_6153,N_5968);
nor U7941 (N_7941,N_6222,N_5713);
and U7942 (N_7942,N_6747,N_7116);
or U7943 (N_7943,N_7133,N_6233);
and U7944 (N_7944,N_5595,N_6179);
and U7945 (N_7945,N_6007,N_6094);
nand U7946 (N_7946,N_5930,N_5531);
or U7947 (N_7947,N_5797,N_5325);
nand U7948 (N_7948,N_5439,N_6313);
and U7949 (N_7949,N_6990,N_6635);
nor U7950 (N_7950,N_5144,N_7151);
nand U7951 (N_7951,N_6969,N_7008);
nor U7952 (N_7952,N_5617,N_7208);
xor U7953 (N_7953,N_7197,N_7088);
nor U7954 (N_7954,N_7489,N_6973);
nand U7955 (N_7955,N_5252,N_5524);
xor U7956 (N_7956,N_5339,N_7156);
and U7957 (N_7957,N_6015,N_5396);
nor U7958 (N_7958,N_6106,N_7118);
and U7959 (N_7959,N_6856,N_5996);
or U7960 (N_7960,N_7281,N_6853);
nand U7961 (N_7961,N_6606,N_5835);
and U7962 (N_7962,N_5159,N_7231);
or U7963 (N_7963,N_6778,N_5045);
or U7964 (N_7964,N_7383,N_6801);
and U7965 (N_7965,N_7340,N_6595);
and U7966 (N_7966,N_5784,N_7490);
nand U7967 (N_7967,N_6398,N_7435);
nand U7968 (N_7968,N_6285,N_5758);
nor U7969 (N_7969,N_5560,N_6837);
and U7970 (N_7970,N_7175,N_7085);
and U7971 (N_7971,N_6760,N_6776);
and U7972 (N_7972,N_5756,N_5472);
xor U7973 (N_7973,N_6965,N_5234);
nor U7974 (N_7974,N_5098,N_6537);
or U7975 (N_7975,N_5317,N_6489);
nand U7976 (N_7976,N_5308,N_6810);
xnor U7977 (N_7977,N_6068,N_6605);
xnor U7978 (N_7978,N_7210,N_7251);
nor U7979 (N_7979,N_6879,N_6010);
nand U7980 (N_7980,N_6948,N_6267);
nor U7981 (N_7981,N_5345,N_5712);
and U7982 (N_7982,N_7241,N_6711);
and U7983 (N_7983,N_5226,N_6389);
nand U7984 (N_7984,N_5931,N_5485);
or U7985 (N_7985,N_7017,N_6425);
nor U7986 (N_7986,N_6132,N_6963);
or U7987 (N_7987,N_5620,N_5683);
or U7988 (N_7988,N_5140,N_5009);
nor U7989 (N_7989,N_7006,N_5213);
or U7990 (N_7990,N_5264,N_7297);
and U7991 (N_7991,N_5571,N_5359);
or U7992 (N_7992,N_5229,N_6243);
nor U7993 (N_7993,N_6283,N_6017);
nand U7994 (N_7994,N_5513,N_5160);
nor U7995 (N_7995,N_6297,N_5719);
xor U7996 (N_7996,N_5066,N_5038);
and U7997 (N_7997,N_5715,N_6234);
nor U7998 (N_7998,N_5989,N_5905);
xor U7999 (N_7999,N_5322,N_6478);
and U8000 (N_8000,N_7235,N_6061);
or U8001 (N_8001,N_5079,N_6324);
nor U8002 (N_8002,N_6930,N_6476);
nand U8003 (N_8003,N_5631,N_6230);
and U8004 (N_8004,N_5212,N_5154);
and U8005 (N_8005,N_5955,N_6075);
nand U8006 (N_8006,N_6746,N_5075);
or U8007 (N_8007,N_6461,N_5280);
nor U8008 (N_8008,N_7328,N_7288);
nand U8009 (N_8009,N_6797,N_6140);
and U8010 (N_8010,N_5490,N_6953);
and U8011 (N_8011,N_6944,N_5839);
and U8012 (N_8012,N_7095,N_6490);
or U8013 (N_8013,N_5169,N_7012);
nand U8014 (N_8014,N_5279,N_6284);
xnor U8015 (N_8015,N_5141,N_7015);
and U8016 (N_8016,N_6753,N_6499);
nor U8017 (N_8017,N_5438,N_5315);
and U8018 (N_8018,N_5971,N_7414);
and U8019 (N_8019,N_6817,N_5519);
nor U8020 (N_8020,N_5184,N_5127);
nor U8021 (N_8021,N_6256,N_6447);
and U8022 (N_8022,N_5131,N_6975);
nor U8023 (N_8023,N_6873,N_6830);
and U8024 (N_8024,N_6781,N_5755);
or U8025 (N_8025,N_5334,N_5084);
or U8026 (N_8026,N_5956,N_6549);
and U8027 (N_8027,N_6145,N_6208);
nand U8028 (N_8028,N_6744,N_7207);
nand U8029 (N_8029,N_6767,N_5688);
nor U8030 (N_8030,N_6229,N_6921);
or U8031 (N_8031,N_7202,N_6545);
and U8032 (N_8032,N_6550,N_6677);
nor U8033 (N_8033,N_7030,N_6894);
nor U8034 (N_8034,N_6370,N_6050);
or U8035 (N_8035,N_6708,N_5799);
nand U8036 (N_8036,N_7058,N_5085);
and U8037 (N_8037,N_6697,N_7226);
and U8038 (N_8038,N_6513,N_6473);
nand U8039 (N_8039,N_5709,N_5533);
nand U8040 (N_8040,N_5447,N_6311);
and U8041 (N_8041,N_6360,N_6136);
and U8042 (N_8042,N_6076,N_6245);
and U8043 (N_8043,N_5547,N_7188);
and U8044 (N_8044,N_7421,N_7123);
and U8045 (N_8045,N_6460,N_5771);
and U8046 (N_8046,N_6562,N_5911);
nand U8047 (N_8047,N_6266,N_7047);
nand U8048 (N_8048,N_6217,N_5869);
or U8049 (N_8049,N_5669,N_6111);
nand U8050 (N_8050,N_5456,N_6424);
nand U8051 (N_8051,N_5451,N_5744);
nor U8052 (N_8052,N_5864,N_5000);
and U8053 (N_8053,N_6964,N_5668);
nand U8054 (N_8054,N_7193,N_5636);
nand U8055 (N_8055,N_7336,N_6724);
nand U8056 (N_8056,N_5833,N_7325);
nand U8057 (N_8057,N_6572,N_6648);
nor U8058 (N_8058,N_5172,N_5462);
nand U8059 (N_8059,N_6546,N_7280);
and U8060 (N_8060,N_5480,N_7317);
and U8061 (N_8061,N_6751,N_7121);
nor U8062 (N_8062,N_5382,N_7463);
nor U8063 (N_8063,N_7185,N_5355);
and U8064 (N_8064,N_5121,N_5507);
nor U8065 (N_8065,N_5626,N_6031);
or U8066 (N_8066,N_6864,N_5410);
xnor U8067 (N_8067,N_6119,N_7205);
nand U8068 (N_8068,N_6931,N_5736);
or U8069 (N_8069,N_5292,N_5242);
nand U8070 (N_8070,N_5587,N_6334);
or U8071 (N_8071,N_5546,N_5337);
or U8072 (N_8072,N_6216,N_6769);
nor U8073 (N_8073,N_7494,N_7139);
nand U8074 (N_8074,N_5166,N_5342);
nand U8075 (N_8075,N_6540,N_6696);
and U8076 (N_8076,N_6174,N_5331);
nor U8077 (N_8077,N_6359,N_5630);
and U8078 (N_8078,N_5150,N_5320);
nor U8079 (N_8079,N_5575,N_6507);
or U8080 (N_8080,N_5984,N_6890);
or U8081 (N_8081,N_5599,N_5773);
and U8082 (N_8082,N_6743,N_6701);
and U8083 (N_8083,N_6632,N_6592);
and U8084 (N_8084,N_6253,N_6827);
and U8085 (N_8085,N_6303,N_5842);
and U8086 (N_8086,N_5774,N_7170);
or U8087 (N_8087,N_7330,N_6899);
nand U8088 (N_8088,N_5319,N_6908);
nand U8089 (N_8089,N_7191,N_5388);
nor U8090 (N_8090,N_5699,N_7219);
nand U8091 (N_8091,N_6871,N_5690);
nor U8092 (N_8092,N_6774,N_7425);
and U8093 (N_8093,N_6035,N_7128);
or U8094 (N_8094,N_6434,N_7132);
nor U8095 (N_8095,N_5593,N_7442);
and U8096 (N_8096,N_5791,N_5530);
nand U8097 (N_8097,N_5615,N_5287);
nand U8098 (N_8098,N_5300,N_5800);
and U8099 (N_8099,N_6912,N_5394);
nand U8100 (N_8100,N_6807,N_7174);
nand U8101 (N_8101,N_5723,N_5059);
nor U8102 (N_8102,N_7166,N_6658);
and U8103 (N_8103,N_6236,N_5118);
and U8104 (N_8104,N_6152,N_6272);
and U8105 (N_8105,N_5951,N_5677);
and U8106 (N_8106,N_7252,N_6279);
nand U8107 (N_8107,N_7499,N_5471);
nor U8108 (N_8108,N_6318,N_6090);
and U8109 (N_8109,N_5794,N_6183);
and U8110 (N_8110,N_7043,N_5845);
or U8111 (N_8111,N_5529,N_5035);
and U8112 (N_8112,N_5349,N_6418);
nand U8113 (N_8113,N_6611,N_7163);
and U8114 (N_8114,N_6003,N_6345);
nand U8115 (N_8115,N_5061,N_6455);
and U8116 (N_8116,N_5129,N_5957);
nor U8117 (N_8117,N_5152,N_7308);
nand U8118 (N_8118,N_6791,N_6761);
nor U8119 (N_8119,N_7433,N_7186);
nor U8120 (N_8120,N_5727,N_7477);
and U8121 (N_8121,N_6702,N_5649);
nor U8122 (N_8122,N_5737,N_6671);
or U8123 (N_8123,N_6186,N_5251);
and U8124 (N_8124,N_5039,N_5199);
nor U8125 (N_8125,N_6951,N_6241);
nand U8126 (N_8126,N_5019,N_6730);
nor U8127 (N_8127,N_6185,N_7048);
nand U8128 (N_8128,N_5348,N_5344);
nand U8129 (N_8129,N_6206,N_6286);
or U8130 (N_8130,N_6762,N_7137);
nor U8131 (N_8131,N_5050,N_7087);
nand U8132 (N_8132,N_5021,N_6019);
and U8133 (N_8133,N_6335,N_6777);
or U8134 (N_8134,N_6038,N_5176);
and U8135 (N_8135,N_5760,N_5650);
and U8136 (N_8136,N_7158,N_5165);
and U8137 (N_8137,N_6597,N_6986);
nand U8138 (N_8138,N_6162,N_6566);
nor U8139 (N_8139,N_5431,N_6500);
nor U8140 (N_8140,N_5897,N_7239);
and U8141 (N_8141,N_6057,N_6333);
or U8142 (N_8142,N_7360,N_6528);
nand U8143 (N_8143,N_6028,N_7353);
nor U8144 (N_8144,N_5586,N_5148);
or U8145 (N_8145,N_5376,N_6869);
nand U8146 (N_8146,N_5900,N_6463);
nor U8147 (N_8147,N_6991,N_5275);
nor U8148 (N_8148,N_7161,N_5309);
nor U8149 (N_8149,N_6521,N_6110);
nor U8150 (N_8150,N_5332,N_5639);
nand U8151 (N_8151,N_5335,N_5214);
nand U8152 (N_8152,N_5364,N_6491);
or U8153 (N_8153,N_6529,N_6177);
nor U8154 (N_8154,N_5598,N_5107);
nand U8155 (N_8155,N_6191,N_7453);
nor U8156 (N_8156,N_5024,N_7286);
nor U8157 (N_8157,N_7276,N_6475);
and U8158 (N_8158,N_5248,N_6980);
or U8159 (N_8159,N_6630,N_7103);
and U8160 (N_8160,N_7126,N_5569);
nor U8161 (N_8161,N_6608,N_5366);
or U8162 (N_8162,N_7247,N_6863);
nand U8163 (N_8163,N_6569,N_5441);
nor U8164 (N_8164,N_5859,N_5832);
and U8165 (N_8165,N_6691,N_7089);
nor U8166 (N_8166,N_5080,N_7037);
and U8167 (N_8167,N_7481,N_6025);
nand U8168 (N_8168,N_7076,N_6329);
nand U8169 (N_8169,N_7419,N_6466);
and U8170 (N_8170,N_5553,N_5323);
or U8171 (N_8171,N_6240,N_6765);
nor U8172 (N_8172,N_7377,N_6201);
nor U8173 (N_8173,N_6954,N_6169);
or U8174 (N_8174,N_6785,N_5596);
or U8175 (N_8175,N_6886,N_5426);
and U8176 (N_8176,N_6616,N_5610);
nand U8177 (N_8177,N_6915,N_6763);
nor U8178 (N_8178,N_6639,N_7256);
and U8179 (N_8179,N_5369,N_5006);
and U8180 (N_8180,N_7408,N_6060);
nor U8181 (N_8181,N_6064,N_5318);
nand U8182 (N_8182,N_7097,N_6657);
nor U8183 (N_8183,N_6645,N_6709);
nand U8184 (N_8184,N_5356,N_5691);
nand U8185 (N_8185,N_6811,N_5881);
or U8186 (N_8186,N_5585,N_5044);
or U8187 (N_8187,N_6992,N_7406);
nand U8188 (N_8188,N_6821,N_6520);
nor U8189 (N_8189,N_5215,N_5659);
and U8190 (N_8190,N_5581,N_5054);
or U8191 (N_8191,N_5623,N_7467);
nand U8192 (N_8192,N_6979,N_6089);
nand U8193 (N_8193,N_6676,N_6836);
or U8194 (N_8194,N_5678,N_5142);
nor U8195 (N_8195,N_7348,N_6436);
nand U8196 (N_8196,N_6238,N_5820);
nor U8197 (N_8197,N_5535,N_5218);
nor U8198 (N_8198,N_5002,N_5087);
and U8199 (N_8199,N_6255,N_6155);
nand U8200 (N_8200,N_5788,N_5013);
nor U8201 (N_8201,N_6583,N_7318);
nand U8202 (N_8202,N_5198,N_7416);
xnor U8203 (N_8203,N_5088,N_6534);
and U8204 (N_8204,N_7306,N_5415);
or U8205 (N_8205,N_6298,N_5232);
nor U8206 (N_8206,N_6154,N_5514);
nor U8207 (N_8207,N_7127,N_5435);
nor U8208 (N_8208,N_5656,N_6518);
and U8209 (N_8209,N_6305,N_5511);
nand U8210 (N_8210,N_6664,N_6946);
or U8211 (N_8211,N_5876,N_5819);
or U8212 (N_8212,N_5372,N_6369);
or U8213 (N_8213,N_6704,N_5895);
nor U8214 (N_8214,N_6163,N_6738);
or U8215 (N_8215,N_7136,N_7057);
and U8216 (N_8216,N_5608,N_7011);
nand U8217 (N_8217,N_5196,N_6996);
or U8218 (N_8218,N_6449,N_6759);
or U8219 (N_8219,N_7184,N_5944);
nand U8220 (N_8220,N_7258,N_7493);
nand U8221 (N_8221,N_5991,N_6900);
or U8222 (N_8222,N_5029,N_7456);
nand U8223 (N_8223,N_5069,N_6194);
nor U8224 (N_8224,N_7195,N_5095);
nand U8225 (N_8225,N_7447,N_6221);
nand U8226 (N_8226,N_6430,N_5105);
nand U8227 (N_8227,N_7373,N_5493);
nand U8228 (N_8228,N_7140,N_6320);
nor U8229 (N_8229,N_7260,N_6338);
xor U8230 (N_8230,N_6116,N_6556);
or U8231 (N_8231,N_5811,N_6706);
and U8232 (N_8232,N_5111,N_6292);
nor U8233 (N_8233,N_6839,N_5289);
and U8234 (N_8234,N_6349,N_7444);
or U8235 (N_8235,N_7036,N_6040);
or U8236 (N_8236,N_7045,N_5939);
nor U8237 (N_8237,N_7430,N_5882);
nand U8238 (N_8238,N_5718,N_6745);
or U8239 (N_8239,N_5387,N_7393);
nand U8240 (N_8240,N_5887,N_7352);
nor U8241 (N_8241,N_6168,N_5885);
nand U8242 (N_8242,N_7299,N_6137);
nor U8243 (N_8243,N_7431,N_6501);
and U8244 (N_8244,N_5316,N_6252);
nand U8245 (N_8245,N_7273,N_5285);
and U8246 (N_8246,N_5469,N_7038);
or U8247 (N_8247,N_6849,N_6672);
or U8248 (N_8248,N_6939,N_5137);
or U8249 (N_8249,N_5500,N_5361);
nand U8250 (N_8250,N_7209,N_7243);
nand U8251 (N_8251,N_5732,N_6736);
or U8252 (N_8252,N_5162,N_5277);
or U8253 (N_8253,N_5299,N_7253);
or U8254 (N_8254,N_7479,N_5350);
and U8255 (N_8255,N_5216,N_5722);
and U8256 (N_8256,N_6884,N_5675);
nand U8257 (N_8257,N_6287,N_7024);
nand U8258 (N_8258,N_5401,N_6417);
nor U8259 (N_8259,N_6112,N_5775);
or U8260 (N_8260,N_7018,N_5852);
and U8261 (N_8261,N_5483,N_5240);
nor U8262 (N_8262,N_7342,N_7400);
and U8263 (N_8263,N_6787,N_5408);
nand U8264 (N_8264,N_7110,N_6988);
nand U8265 (N_8265,N_6613,N_6034);
or U8266 (N_8266,N_6714,N_7446);
and U8267 (N_8267,N_6415,N_6393);
and U8268 (N_8268,N_6877,N_6458);
or U8269 (N_8269,N_7475,N_6907);
nand U8270 (N_8270,N_5934,N_7052);
and U8271 (N_8271,N_6541,N_6109);
nor U8272 (N_8272,N_6570,N_7484);
nor U8273 (N_8273,N_6375,N_7331);
nand U8274 (N_8274,N_5202,N_5558);
or U8275 (N_8275,N_7107,N_6784);
or U8276 (N_8276,N_7275,N_6321);
xnor U8277 (N_8277,N_6129,N_5180);
and U8278 (N_8278,N_5765,N_6750);
or U8279 (N_8279,N_5721,N_6823);
and U8280 (N_8280,N_6780,N_5284);
nor U8281 (N_8281,N_6494,N_6881);
nand U8282 (N_8282,N_6052,N_6689);
and U8283 (N_8283,N_7491,N_5474);
or U8284 (N_8284,N_6725,N_6118);
nand U8285 (N_8285,N_7423,N_6073);
nand U8286 (N_8286,N_7324,N_6740);
or U8287 (N_8287,N_6970,N_5921);
or U8288 (N_8288,N_5103,N_6312);
or U8289 (N_8289,N_6845,N_7014);
nor U8290 (N_8290,N_6012,N_5422);
nand U8291 (N_8291,N_5803,N_7387);
nor U8292 (N_8292,N_6164,N_6198);
and U8293 (N_8293,N_6184,N_5979);
nor U8294 (N_8294,N_7474,N_5821);
nand U8295 (N_8295,N_5628,N_6527);
and U8296 (N_8296,N_5302,N_5042);
and U8297 (N_8297,N_6299,N_5110);
nor U8298 (N_8298,N_7392,N_5056);
and U8299 (N_8299,N_5517,N_6248);
or U8300 (N_8300,N_5851,N_5051);
and U8301 (N_8301,N_5149,N_6401);
nor U8302 (N_8302,N_6016,N_7257);
or U8303 (N_8303,N_5468,N_5303);
and U8304 (N_8304,N_5250,N_6331);
nor U8305 (N_8305,N_5389,N_5032);
or U8306 (N_8306,N_6773,N_5868);
nor U8307 (N_8307,N_6719,N_5917);
nand U8308 (N_8308,N_5026,N_6631);
nor U8309 (N_8309,N_6771,N_6772);
and U8310 (N_8310,N_6433,N_5207);
and U8311 (N_8311,N_6488,N_6362);
or U8312 (N_8312,N_5826,N_7213);
nor U8313 (N_8313,N_6301,N_6097);
nand U8314 (N_8314,N_6486,N_5076);
or U8315 (N_8315,N_6300,N_6687);
and U8316 (N_8316,N_7259,N_6805);
and U8317 (N_8317,N_6865,N_7314);
and U8318 (N_8318,N_5779,N_6077);
xnor U8319 (N_8319,N_7201,N_6508);
and U8320 (N_8320,N_5053,N_6307);
xnor U8321 (N_8321,N_7027,N_5574);
and U8322 (N_8322,N_6013,N_5020);
and U8323 (N_8323,N_5484,N_5972);
nor U8324 (N_8324,N_6203,N_5269);
nor U8325 (N_8325,N_5816,N_5805);
or U8326 (N_8326,N_5825,N_7358);
or U8327 (N_8327,N_7388,N_7054);
nor U8328 (N_8328,N_5397,N_5753);
nor U8329 (N_8329,N_6737,N_5992);
nor U8330 (N_8330,N_6633,N_5730);
and U8331 (N_8331,N_5068,N_5590);
and U8332 (N_8332,N_6049,N_5477);
and U8333 (N_8333,N_5664,N_6380);
and U8334 (N_8334,N_6828,N_5017);
nand U8335 (N_8335,N_5562,N_5241);
or U8336 (N_8336,N_5861,N_5188);
nor U8337 (N_8337,N_5340,N_7487);
and U8338 (N_8338,N_7099,N_6095);
nand U8339 (N_8339,N_7295,N_6409);
nor U8340 (N_8340,N_5559,N_5040);
and U8341 (N_8341,N_5512,N_7056);
and U8342 (N_8342,N_6947,N_6215);
or U8343 (N_8343,N_5648,N_6731);
and U8344 (N_8344,N_6938,N_6707);
or U8345 (N_8345,N_6024,N_5990);
nor U8346 (N_8346,N_7134,N_5022);
nand U8347 (N_8347,N_6985,N_6431);
or U8348 (N_8348,N_6723,N_7264);
and U8349 (N_8349,N_7361,N_6497);
nor U8350 (N_8350,N_5497,N_5362);
or U8351 (N_8351,N_7216,N_5119);
nand U8352 (N_8352,N_5268,N_5726);
or U8353 (N_8353,N_5177,N_6239);
nand U8354 (N_8354,N_6906,N_5179);
nor U8355 (N_8355,N_7221,N_5544);
nand U8356 (N_8356,N_6553,N_5282);
and U8357 (N_8357,N_6356,N_6859);
and U8358 (N_8358,N_5249,N_5312);
nor U8359 (N_8359,N_7357,N_6441);
and U8360 (N_8360,N_7154,N_6350);
and U8361 (N_8361,N_5425,N_7149);
nor U8362 (N_8362,N_5102,N_7356);
nand U8363 (N_8363,N_5052,N_5089);
or U8364 (N_8364,N_6023,N_5239);
nand U8365 (N_8365,N_5616,N_5708);
nor U8366 (N_8366,N_5878,N_6275);
or U8367 (N_8367,N_6783,N_5909);
and U8368 (N_8368,N_6903,N_5018);
or U8369 (N_8369,N_6046,N_6071);
nand U8370 (N_8370,N_7443,N_5766);
nand U8371 (N_8371,N_6848,N_6480);
nand U8372 (N_8372,N_7310,N_7042);
or U8373 (N_8373,N_5260,N_6000);
or U8374 (N_8374,N_5890,N_7450);
nand U8375 (N_8375,N_5564,N_5783);
and U8376 (N_8376,N_6796,N_5034);
xnor U8377 (N_8377,N_6775,N_5170);
nand U8378 (N_8378,N_6444,N_6242);
nor U8379 (N_8379,N_6679,N_6601);
nand U8380 (N_8380,N_5695,N_7403);
or U8381 (N_8381,N_6402,N_6400);
xnor U8382 (N_8382,N_6316,N_5841);
nor U8383 (N_8383,N_5090,N_5652);
and U8384 (N_8384,N_5096,N_5360);
nand U8385 (N_8385,N_7172,N_5993);
and U8386 (N_8386,N_5383,N_6505);
and U8387 (N_8387,N_7153,N_5116);
nor U8388 (N_8388,N_5802,N_7300);
nand U8389 (N_8389,N_5830,N_7386);
nand U8390 (N_8390,N_5624,N_6226);
and U8391 (N_8391,N_6555,N_5740);
and U8392 (N_8392,N_6582,N_7333);
or U8393 (N_8393,N_6560,N_5908);
or U8394 (N_8394,N_5752,N_6365);
nand U8395 (N_8395,N_5445,N_5938);
nor U8396 (N_8396,N_7236,N_7407);
or U8397 (N_8397,N_6231,N_5192);
or U8398 (N_8398,N_5686,N_7124);
xnor U8399 (N_8399,N_5293,N_5621);
and U8400 (N_8400,N_5954,N_5378);
or U8401 (N_8401,N_6413,N_6533);
nor U8402 (N_8402,N_5173,N_5031);
and U8403 (N_8403,N_6021,N_7093);
nor U8404 (N_8404,N_5922,N_5354);
nor U8405 (N_8405,N_7167,N_6396);
or U8406 (N_8406,N_5138,N_6950);
and U8407 (N_8407,N_5509,N_6579);
nor U8408 (N_8408,N_5635,N_5464);
or U8409 (N_8409,N_5687,N_7080);
nor U8410 (N_8410,N_6121,N_6984);
or U8411 (N_8411,N_6825,N_6993);
nor U8412 (N_8412,N_5028,N_7415);
or U8413 (N_8413,N_5057,N_6941);
nand U8414 (N_8414,N_7053,N_6809);
nor U8415 (N_8415,N_5637,N_7100);
nand U8416 (N_8416,N_6620,N_5128);
and U8417 (N_8417,N_6048,N_7422);
nand U8418 (N_8418,N_5101,N_6681);
and U8419 (N_8419,N_6758,N_7098);
or U8420 (N_8420,N_6428,N_6919);
or U8421 (N_8421,N_6072,N_5147);
or U8422 (N_8422,N_6596,N_5498);
or U8423 (N_8423,N_7399,N_5433);
and U8424 (N_8424,N_7029,N_6943);
nand U8425 (N_8425,N_6644,N_5701);
and U8426 (N_8426,N_5341,N_5418);
and U8427 (N_8427,N_5696,N_7194);
and U8428 (N_8428,N_7250,N_6412);
or U8429 (N_8429,N_6617,N_5879);
nand U8430 (N_8430,N_6178,N_5301);
nor U8431 (N_8431,N_5219,N_7035);
or U8432 (N_8432,N_5970,N_6464);
or U8433 (N_8433,N_5780,N_6125);
and U8434 (N_8434,N_6456,N_7051);
and U8435 (N_8435,N_6440,N_7398);
nand U8436 (N_8436,N_5785,N_5454);
nor U8437 (N_8437,N_6840,N_5421);
and U8438 (N_8438,N_7438,N_6826);
or U8439 (N_8439,N_5837,N_7471);
and U8440 (N_8440,N_6742,N_7418);
nor U8441 (N_8441,N_6280,N_5419);
and U8442 (N_8442,N_7305,N_5449);
nor U8443 (N_8443,N_5238,N_6768);
nor U8444 (N_8444,N_5750,N_6157);
or U8445 (N_8445,N_5871,N_5682);
nand U8446 (N_8446,N_5867,N_5283);
and U8447 (N_8447,N_6218,N_6404);
nor U8448 (N_8448,N_5463,N_5915);
nand U8449 (N_8449,N_6510,N_5886);
xor U8450 (N_8450,N_5351,N_5937);
nor U8451 (N_8451,N_7065,N_7050);
nand U8452 (N_8452,N_6800,N_7498);
or U8453 (N_8453,N_5467,N_5787);
nand U8454 (N_8454,N_6748,N_5929);
and U8455 (N_8455,N_5055,N_7322);
nor U8456 (N_8456,N_5704,N_6059);
or U8457 (N_8457,N_5742,N_6363);
nor U8458 (N_8458,N_7198,N_6372);
or U8459 (N_8459,N_6083,N_6146);
nor U8460 (N_8460,N_7102,N_5448);
or U8461 (N_8461,N_6101,N_6442);
nor U8462 (N_8462,N_7384,N_7269);
nand U8463 (N_8463,N_5099,N_5946);
or U8464 (N_8464,N_5060,N_6599);
nor U8465 (N_8465,N_7405,N_6084);
and U8466 (N_8466,N_7199,N_6199);
or U8467 (N_8467,N_5012,N_5304);
and U8468 (N_8468,N_7150,N_5297);
nor U8469 (N_8469,N_7233,N_5633);
nor U8470 (N_8470,N_6674,N_6808);
or U8471 (N_8471,N_5094,N_6142);
or U8472 (N_8472,N_6591,N_5181);
nor U8473 (N_8473,N_7073,N_5875);
nand U8474 (N_8474,N_7369,N_5757);
and U8475 (N_8475,N_6995,N_6568);
or U8476 (N_8476,N_7162,N_6989);
and U8477 (N_8477,N_7020,N_5761);
xnor U8478 (N_8478,N_7049,N_5627);
nor U8479 (N_8479,N_6282,N_5962);
and U8480 (N_8480,N_7312,N_7376);
nor U8481 (N_8481,N_5452,N_5157);
and U8482 (N_8482,N_6099,N_6278);
nor U8483 (N_8483,N_5792,N_5423);
nand U8484 (N_8484,N_6661,N_5940);
nor U8485 (N_8485,N_5914,N_6161);
nand U8486 (N_8486,N_7298,N_5097);
nand U8487 (N_8487,N_6971,N_6472);
nand U8488 (N_8488,N_5327,N_5948);
and U8489 (N_8489,N_6432,N_6659);
nand U8490 (N_8490,N_5406,N_6295);
nand U8491 (N_8491,N_7165,N_5168);
and U8492 (N_8492,N_5357,N_7189);
or U8493 (N_8493,N_5314,N_7355);
nand U8494 (N_8494,N_7145,N_6361);
or U8495 (N_8495,N_6968,N_6851);
nand U8496 (N_8496,N_5973,N_6652);
and U8497 (N_8497,N_6699,N_6983);
nor U8498 (N_8498,N_7224,N_5584);
and U8499 (N_8499,N_6885,N_5011);
and U8500 (N_8500,N_7000,N_5980);
nand U8501 (N_8501,N_7390,N_7445);
nand U8502 (N_8502,N_5672,N_6998);
or U8503 (N_8503,N_5772,N_7410);
and U8504 (N_8504,N_5298,N_6854);
and U8505 (N_8505,N_7152,N_5036);
and U8506 (N_8506,N_6835,N_5145);
nor U8507 (N_8507,N_6394,N_6766);
nor U8508 (N_8508,N_6330,N_6227);
and U8509 (N_8509,N_6503,N_6614);
and U8510 (N_8510,N_6875,N_5961);
xor U8511 (N_8511,N_5824,N_5958);
nor U8512 (N_8512,N_5714,N_7492);
or U8513 (N_8513,N_6087,N_7092);
nor U8514 (N_8514,N_7142,N_5781);
nand U8515 (N_8515,N_6131,N_6713);
nand U8516 (N_8516,N_6482,N_7274);
or U8517 (N_8517,N_6314,N_7086);
or U8518 (N_8518,N_7228,N_6876);
nand U8519 (N_8519,N_6205,N_7108);
nand U8520 (N_8520,N_6070,N_6913);
nor U8521 (N_8521,N_7321,N_6575);
nand U8522 (N_8522,N_5186,N_6141);
nand U8523 (N_8523,N_6247,N_7144);
and U8524 (N_8524,N_6559,N_6397);
nor U8525 (N_8525,N_6668,N_6344);
or U8526 (N_8526,N_5270,N_6929);
nand U8527 (N_8527,N_5404,N_6670);
nor U8528 (N_8528,N_6270,N_6005);
nor U8529 (N_8529,N_6842,N_6092);
nor U8530 (N_8530,N_7081,N_5891);
and U8531 (N_8531,N_5208,N_6133);
or U8532 (N_8532,N_5041,N_5461);
and U8533 (N_8533,N_5583,N_7157);
nor U8534 (N_8534,N_6716,N_7378);
and U8535 (N_8535,N_6262,N_5206);
nand U8536 (N_8536,N_7135,N_5200);
and U8537 (N_8537,N_5189,N_5368);
nand U8538 (N_8538,N_7125,N_5132);
and U8539 (N_8539,N_6276,N_5358);
nor U8540 (N_8540,N_7349,N_7470);
nor U8541 (N_8541,N_5865,N_5998);
nor U8542 (N_8542,N_7225,N_6406);
or U8543 (N_8543,N_5846,N_5446);
nand U8544 (N_8544,N_6880,N_6437);
nand U8545 (N_8545,N_7441,N_6228);
and U8546 (N_8546,N_5666,N_5565);
xnor U8547 (N_8547,N_5982,N_6901);
xnor U8548 (N_8548,N_5255,N_5622);
and U8549 (N_8549,N_6653,N_5458);
nand U8550 (N_8550,N_5542,N_5476);
nor U8551 (N_8551,N_6261,N_5866);
nand U8552 (N_8552,N_7413,N_5528);
nand U8553 (N_8553,N_5673,N_5548);
or U8554 (N_8554,N_7062,N_6487);
and U8555 (N_8555,N_6584,N_6373);
and U8556 (N_8556,N_6862,N_6813);
or U8557 (N_8557,N_6326,N_5964);
and U8558 (N_8558,N_5139,N_6209);
or U8559 (N_8559,N_5679,N_6274);
and U8560 (N_8560,N_6577,N_6047);
nor U8561 (N_8561,N_6640,N_5352);
xnor U8562 (N_8562,N_6006,N_7272);
nand U8563 (N_8563,N_6543,N_6594);
or U8564 (N_8564,N_5995,N_5949);
nand U8565 (N_8565,N_6634,N_5907);
nor U8566 (N_8566,N_6798,N_5614);
and U8567 (N_8567,N_5912,N_6459);
xor U8568 (N_8568,N_7350,N_5491);
or U8569 (N_8569,N_6148,N_6916);
or U8570 (N_8570,N_6192,N_6158);
and U8571 (N_8571,N_5680,N_5828);
and U8572 (N_8572,N_6268,N_6926);
nand U8573 (N_8573,N_7223,N_6302);
nand U8574 (N_8574,N_5817,N_6108);
nand U8575 (N_8575,N_5416,N_5228);
and U8576 (N_8576,N_6408,N_6045);
nor U8577 (N_8577,N_6457,N_7296);
xnor U8578 (N_8578,N_7391,N_6824);
and U8579 (N_8579,N_7164,N_7311);
and U8580 (N_8580,N_5834,N_5429);
xnor U8581 (N_8581,N_5716,N_5612);
nand U8582 (N_8582,N_6281,N_6306);
nor U8583 (N_8583,N_5983,N_5848);
nand U8584 (N_8584,N_6128,N_5143);
nor U8585 (N_8585,N_6962,N_5822);
and U8586 (N_8586,N_6512,N_6590);
nand U8587 (N_8587,N_6524,N_5918);
xor U8588 (N_8588,N_6190,N_5286);
nand U8589 (N_8589,N_5619,N_6443);
or U8590 (N_8590,N_7337,N_6542);
nand U8591 (N_8591,N_6868,N_7335);
nand U8592 (N_8592,N_6484,N_6833);
nor U8593 (N_8593,N_7046,N_7143);
nand U8594 (N_8594,N_7354,N_6933);
nor U8595 (N_8595,N_5265,N_6454);
xnor U8596 (N_8596,N_5233,N_6538);
or U8597 (N_8597,N_6065,N_5928);
nand U8598 (N_8598,N_5808,N_5515);
or U8599 (N_8599,N_5403,N_6337);
or U8600 (N_8600,N_5231,N_5135);
or U8601 (N_8601,N_5734,N_6655);
nor U8602 (N_8602,N_6850,N_5412);
and U8603 (N_8603,N_5807,N_5589);
or U8604 (N_8604,N_5030,N_5926);
nand U8605 (N_8605,N_7437,N_6739);
or U8606 (N_8606,N_7010,N_7412);
and U8607 (N_8607,N_6593,N_7013);
nand U8608 (N_8608,N_6088,N_6637);
or U8609 (N_8609,N_5072,N_6465);
and U8610 (N_8610,N_5545,N_6870);
nor U8611 (N_8611,N_6339,N_6450);
nand U8612 (N_8612,N_5863,N_6581);
nand U8613 (N_8613,N_6779,N_6171);
nand U8614 (N_8614,N_7039,N_7497);
nor U8615 (N_8615,N_7025,N_5611);
or U8616 (N_8616,N_5064,N_7072);
nor U8617 (N_8617,N_6603,N_6063);
or U8618 (N_8618,N_7397,N_6959);
nor U8619 (N_8619,N_7265,N_5960);
and U8620 (N_8620,N_6037,N_6001);
and U8621 (N_8621,N_6564,N_5768);
nand U8622 (N_8622,N_6790,N_7255);
and U8623 (N_8623,N_7266,N_6376);
nor U8624 (N_8624,N_7032,N_7007);
nand U8625 (N_8625,N_7345,N_6008);
or U8626 (N_8626,N_5597,N_6195);
or U8627 (N_8627,N_6091,N_6675);
and U8628 (N_8628,N_5081,N_6421);
nor U8629 (N_8629,N_5913,N_5399);
xnor U8630 (N_8630,N_5665,N_7448);
nor U8631 (N_8631,N_7401,N_6860);
and U8632 (N_8632,N_7434,N_6100);
nand U8633 (N_8633,N_5645,N_5310);
and U8634 (N_8634,N_5221,N_6718);
and U8635 (N_8635,N_7064,N_7432);
nand U8636 (N_8636,N_5353,N_5167);
nand U8637 (N_8637,N_6263,N_7222);
nor U8638 (N_8638,N_7067,N_7426);
or U8639 (N_8639,N_5413,N_5033);
or U8640 (N_8640,N_5194,N_7176);
or U8641 (N_8641,N_7465,N_6189);
or U8642 (N_8642,N_7480,N_6151);
or U8643 (N_8643,N_6182,N_7458);
xor U8644 (N_8644,N_6170,N_6469);
nor U8645 (N_8645,N_6439,N_6685);
or U8646 (N_8646,N_7159,N_6032);
nor U8647 (N_8647,N_6804,N_5812);
and U8648 (N_8648,N_5380,N_7359);
nand U8649 (N_8649,N_7409,N_7254);
xnor U8650 (N_8650,N_5254,N_7279);
nor U8651 (N_8651,N_6693,N_5607);
or U8652 (N_8652,N_5903,N_6669);
nor U8653 (N_8653,N_5795,N_7301);
nor U8654 (N_8654,N_7155,N_6897);
or U8655 (N_8655,N_7019,N_7245);
or U8656 (N_8656,N_6847,N_5236);
nor U8657 (N_8657,N_5023,N_6080);
or U8658 (N_8658,N_6471,N_5460);
or U8659 (N_8659,N_7004,N_5698);
nand U8660 (N_8660,N_6134,N_5978);
or U8661 (N_8661,N_7334,N_6574);
nand U8662 (N_8662,N_6547,N_7452);
or U8663 (N_8663,N_6249,N_6987);
or U8664 (N_8664,N_6838,N_5442);
nand U8665 (N_8665,N_7182,N_6551);
or U8666 (N_8666,N_7420,N_5862);
nand U8667 (N_8667,N_7169,N_7454);
or U8668 (N_8668,N_5769,N_6042);
or U8669 (N_8669,N_7424,N_7478);
nor U8670 (N_8670,N_5782,N_5684);
nand U8671 (N_8671,N_7302,N_6957);
and U8672 (N_8672,N_6382,N_5256);
nand U8673 (N_8673,N_6703,N_6893);
nor U8674 (N_8674,N_5083,N_6127);
or U8675 (N_8675,N_6922,N_6909);
and U8676 (N_8676,N_5225,N_7168);
and U8677 (N_8677,N_6587,N_5901);
or U8678 (N_8678,N_6721,N_7083);
or U8679 (N_8679,N_5222,N_7270);
or U8680 (N_8680,N_5936,N_6923);
or U8681 (N_8681,N_6786,N_6104);
and U8682 (N_8682,N_5883,N_6211);
or U8683 (N_8683,N_7459,N_5857);
nand U8684 (N_8684,N_7106,N_6536);
nand U8685 (N_8685,N_7464,N_6202);
or U8686 (N_8686,N_7338,N_5877);
and U8687 (N_8687,N_6379,N_5245);
and U8688 (N_8688,N_5365,N_5328);
or U8689 (N_8689,N_6336,N_5950);
or U8690 (N_8690,N_7217,N_6937);
nand U8691 (N_8691,N_5551,N_5642);
and U8692 (N_8692,N_6271,N_6225);
or U8693 (N_8693,N_6795,N_6018);
and U8694 (N_8694,N_7344,N_6098);
xor U8695 (N_8695,N_6366,N_5210);
or U8696 (N_8696,N_7371,N_7396);
nand U8697 (N_8697,N_6532,N_6720);
and U8698 (N_8698,N_5893,N_6355);
or U8699 (N_8699,N_7044,N_6621);
nor U8700 (N_8700,N_6793,N_5986);
or U8701 (N_8701,N_6586,N_5091);
nor U8702 (N_8702,N_6506,N_5211);
nand U8703 (N_8703,N_5346,N_5894);
or U8704 (N_8704,N_6843,N_5185);
nor U8705 (N_8705,N_7069,N_6607);
or U8706 (N_8706,N_7332,N_6197);
or U8707 (N_8707,N_6565,N_5313);
or U8708 (N_8708,N_6932,N_5502);
and U8709 (N_8709,N_6332,N_5370);
or U8710 (N_8710,N_6612,N_7248);
and U8711 (N_8711,N_7212,N_5108);
or U8712 (N_8712,N_6390,N_5048);
nor U8713 (N_8713,N_6642,N_5120);
or U8714 (N_8714,N_6678,N_6732);
nor U8715 (N_8715,N_5136,N_6254);
nor U8716 (N_8716,N_7292,N_5818);
or U8717 (N_8717,N_7307,N_6328);
or U8718 (N_8718,N_5601,N_6493);
nand U8719 (N_8719,N_7146,N_5693);
and U8720 (N_8720,N_7148,N_6411);
and U8721 (N_8721,N_5923,N_5976);
and U8722 (N_8722,N_6515,N_7082);
nand U8723 (N_8723,N_5770,N_5164);
nor U8724 (N_8724,N_6403,N_6816);
and U8725 (N_8725,N_6093,N_6663);
xnor U8726 (N_8726,N_5746,N_5577);
nand U8727 (N_8727,N_6945,N_6113);
nand U8728 (N_8728,N_5777,N_5910);
nand U8729 (N_8729,N_6105,N_5543);
and U8730 (N_8730,N_5702,N_6429);
or U8731 (N_8731,N_5969,N_6755);
or U8732 (N_8732,N_7496,N_5600);
or U8733 (N_8733,N_5810,N_6960);
nand U8734 (N_8734,N_6056,N_6967);
or U8735 (N_8735,N_6079,N_5424);
nor U8736 (N_8736,N_7131,N_7096);
nand U8737 (N_8737,N_6160,N_5643);
and U8738 (N_8738,N_5305,N_5276);
and U8739 (N_8739,N_6799,N_5414);
nor U8740 (N_8740,N_5504,N_7327);
nand U8741 (N_8741,N_7476,N_6014);
or U8742 (N_8742,N_6315,N_7120);
nor U8743 (N_8743,N_7077,N_7368);
or U8744 (N_8744,N_6385,N_6619);
nand U8745 (N_8745,N_6081,N_5278);
nor U8746 (N_8746,N_7028,N_7016);
nor U8747 (N_8747,N_6504,N_5058);
nand U8748 (N_8748,N_5495,N_5798);
nand U8749 (N_8749,N_6173,N_5247);
nor U8750 (N_8750,N_5512,N_7376);
nor U8751 (N_8751,N_5474,N_7279);
and U8752 (N_8752,N_5688,N_5496);
nor U8753 (N_8753,N_5774,N_6113);
nand U8754 (N_8754,N_6288,N_7380);
nand U8755 (N_8755,N_7327,N_6068);
nand U8756 (N_8756,N_5853,N_6887);
or U8757 (N_8757,N_5350,N_5662);
nor U8758 (N_8758,N_6598,N_5105);
or U8759 (N_8759,N_7049,N_5280);
nor U8760 (N_8760,N_7466,N_5373);
and U8761 (N_8761,N_7260,N_5652);
nor U8762 (N_8762,N_5151,N_6897);
nand U8763 (N_8763,N_7086,N_6948);
and U8764 (N_8764,N_6770,N_5427);
nor U8765 (N_8765,N_6469,N_6027);
and U8766 (N_8766,N_5686,N_5351);
nor U8767 (N_8767,N_5239,N_6450);
nor U8768 (N_8768,N_5909,N_7260);
and U8769 (N_8769,N_5491,N_5957);
nor U8770 (N_8770,N_7071,N_5317);
and U8771 (N_8771,N_7024,N_6092);
nand U8772 (N_8772,N_5292,N_6902);
or U8773 (N_8773,N_5528,N_5086);
and U8774 (N_8774,N_7193,N_6715);
or U8775 (N_8775,N_6943,N_6433);
and U8776 (N_8776,N_6864,N_7085);
nand U8777 (N_8777,N_6313,N_6072);
nor U8778 (N_8778,N_7009,N_7208);
or U8779 (N_8779,N_5200,N_7028);
and U8780 (N_8780,N_7477,N_6619);
nand U8781 (N_8781,N_6988,N_6831);
and U8782 (N_8782,N_7094,N_5306);
or U8783 (N_8783,N_7461,N_5348);
and U8784 (N_8784,N_6478,N_5955);
nor U8785 (N_8785,N_5116,N_6579);
nand U8786 (N_8786,N_6684,N_5674);
nand U8787 (N_8787,N_5718,N_6067);
or U8788 (N_8788,N_6823,N_7295);
and U8789 (N_8789,N_7237,N_5972);
nand U8790 (N_8790,N_5693,N_5343);
or U8791 (N_8791,N_5251,N_7424);
nand U8792 (N_8792,N_7275,N_6662);
nand U8793 (N_8793,N_6224,N_5856);
or U8794 (N_8794,N_7102,N_5498);
and U8795 (N_8795,N_7479,N_7308);
nand U8796 (N_8796,N_7120,N_6208);
nand U8797 (N_8797,N_7293,N_7068);
and U8798 (N_8798,N_5726,N_7282);
nor U8799 (N_8799,N_7470,N_6281);
nor U8800 (N_8800,N_5984,N_5596);
or U8801 (N_8801,N_6135,N_6989);
and U8802 (N_8802,N_5444,N_5650);
nor U8803 (N_8803,N_5782,N_6954);
nor U8804 (N_8804,N_5941,N_5994);
and U8805 (N_8805,N_5671,N_5608);
xor U8806 (N_8806,N_6398,N_5393);
nor U8807 (N_8807,N_5979,N_7279);
nor U8808 (N_8808,N_5065,N_5889);
and U8809 (N_8809,N_5304,N_5244);
or U8810 (N_8810,N_6007,N_6261);
and U8811 (N_8811,N_6507,N_7097);
nor U8812 (N_8812,N_6935,N_5179);
or U8813 (N_8813,N_6621,N_5391);
nand U8814 (N_8814,N_5947,N_6470);
nor U8815 (N_8815,N_6928,N_5679);
xor U8816 (N_8816,N_5632,N_6110);
or U8817 (N_8817,N_6919,N_7432);
and U8818 (N_8818,N_5779,N_6757);
and U8819 (N_8819,N_5937,N_5099);
and U8820 (N_8820,N_5152,N_6607);
nor U8821 (N_8821,N_7226,N_5485);
and U8822 (N_8822,N_7488,N_6754);
xor U8823 (N_8823,N_6581,N_7102);
nand U8824 (N_8824,N_6238,N_5090);
xor U8825 (N_8825,N_7038,N_6200);
nand U8826 (N_8826,N_5048,N_6329);
and U8827 (N_8827,N_5672,N_6519);
or U8828 (N_8828,N_7031,N_6242);
nor U8829 (N_8829,N_6017,N_5861);
and U8830 (N_8830,N_6482,N_5091);
nand U8831 (N_8831,N_6580,N_6456);
nand U8832 (N_8832,N_6969,N_5500);
nor U8833 (N_8833,N_6538,N_6899);
or U8834 (N_8834,N_7098,N_5655);
nand U8835 (N_8835,N_5292,N_5890);
or U8836 (N_8836,N_6773,N_5078);
or U8837 (N_8837,N_7355,N_7424);
nor U8838 (N_8838,N_7339,N_6539);
or U8839 (N_8839,N_5546,N_5259);
or U8840 (N_8840,N_6140,N_6687);
nor U8841 (N_8841,N_6368,N_6249);
and U8842 (N_8842,N_5202,N_5768);
or U8843 (N_8843,N_6789,N_5081);
nand U8844 (N_8844,N_7309,N_6112);
nand U8845 (N_8845,N_7212,N_5139);
nand U8846 (N_8846,N_5834,N_5490);
and U8847 (N_8847,N_5663,N_5003);
nand U8848 (N_8848,N_6502,N_6049);
or U8849 (N_8849,N_6697,N_5983);
and U8850 (N_8850,N_6265,N_6533);
nand U8851 (N_8851,N_7271,N_6987);
nand U8852 (N_8852,N_6760,N_5935);
and U8853 (N_8853,N_7208,N_6947);
and U8854 (N_8854,N_7218,N_6454);
or U8855 (N_8855,N_6266,N_5659);
nor U8856 (N_8856,N_6110,N_6372);
and U8857 (N_8857,N_6357,N_7258);
or U8858 (N_8858,N_6669,N_5029);
nor U8859 (N_8859,N_5356,N_6058);
nand U8860 (N_8860,N_6175,N_5177);
nand U8861 (N_8861,N_5770,N_6103);
nand U8862 (N_8862,N_6772,N_7085);
or U8863 (N_8863,N_6461,N_5127);
or U8864 (N_8864,N_6998,N_5262);
and U8865 (N_8865,N_5848,N_5502);
nand U8866 (N_8866,N_6596,N_6732);
or U8867 (N_8867,N_5598,N_5145);
nor U8868 (N_8868,N_5702,N_6397);
or U8869 (N_8869,N_7073,N_5318);
nor U8870 (N_8870,N_5640,N_5248);
nand U8871 (N_8871,N_5089,N_5084);
nand U8872 (N_8872,N_6757,N_6745);
or U8873 (N_8873,N_5309,N_6484);
and U8874 (N_8874,N_5910,N_6193);
and U8875 (N_8875,N_5746,N_7466);
and U8876 (N_8876,N_5410,N_6154);
or U8877 (N_8877,N_5232,N_5118);
and U8878 (N_8878,N_5391,N_7120);
or U8879 (N_8879,N_5745,N_6153);
or U8880 (N_8880,N_6120,N_5034);
or U8881 (N_8881,N_5952,N_5591);
or U8882 (N_8882,N_6600,N_5031);
or U8883 (N_8883,N_6013,N_6939);
or U8884 (N_8884,N_7095,N_6114);
nor U8885 (N_8885,N_5287,N_5186);
nand U8886 (N_8886,N_5318,N_7148);
or U8887 (N_8887,N_5073,N_6377);
nand U8888 (N_8888,N_6808,N_6067);
nand U8889 (N_8889,N_6830,N_7067);
nand U8890 (N_8890,N_6683,N_5830);
nor U8891 (N_8891,N_5796,N_5181);
nor U8892 (N_8892,N_6110,N_6748);
or U8893 (N_8893,N_6051,N_5047);
nor U8894 (N_8894,N_5999,N_5568);
and U8895 (N_8895,N_6795,N_7102);
and U8896 (N_8896,N_5050,N_5379);
and U8897 (N_8897,N_5573,N_6748);
nand U8898 (N_8898,N_6252,N_5996);
nor U8899 (N_8899,N_7441,N_7254);
or U8900 (N_8900,N_6829,N_5027);
or U8901 (N_8901,N_6314,N_6966);
nor U8902 (N_8902,N_7051,N_6900);
nor U8903 (N_8903,N_5395,N_5165);
and U8904 (N_8904,N_6263,N_7015);
and U8905 (N_8905,N_6826,N_5844);
nor U8906 (N_8906,N_6775,N_6565);
nand U8907 (N_8907,N_6791,N_6114);
nor U8908 (N_8908,N_7260,N_5869);
or U8909 (N_8909,N_7267,N_5866);
nor U8910 (N_8910,N_6062,N_6467);
or U8911 (N_8911,N_5267,N_5139);
and U8912 (N_8912,N_7272,N_5483);
nand U8913 (N_8913,N_6759,N_6703);
nor U8914 (N_8914,N_6412,N_6189);
nand U8915 (N_8915,N_7196,N_5379);
or U8916 (N_8916,N_7347,N_5190);
nand U8917 (N_8917,N_7098,N_5632);
nand U8918 (N_8918,N_7421,N_6240);
and U8919 (N_8919,N_6663,N_5191);
and U8920 (N_8920,N_6737,N_5335);
or U8921 (N_8921,N_5899,N_5369);
nand U8922 (N_8922,N_5097,N_7146);
nand U8923 (N_8923,N_7061,N_6736);
xor U8924 (N_8924,N_7335,N_7081);
nand U8925 (N_8925,N_6931,N_6365);
and U8926 (N_8926,N_5496,N_6487);
or U8927 (N_8927,N_7209,N_5759);
nand U8928 (N_8928,N_6331,N_5936);
nor U8929 (N_8929,N_5040,N_7120);
or U8930 (N_8930,N_5973,N_6487);
nand U8931 (N_8931,N_6224,N_5493);
nand U8932 (N_8932,N_7278,N_6784);
nor U8933 (N_8933,N_5315,N_7115);
or U8934 (N_8934,N_5980,N_6044);
nand U8935 (N_8935,N_7416,N_7448);
xor U8936 (N_8936,N_7054,N_5220);
nor U8937 (N_8937,N_6753,N_7357);
nor U8938 (N_8938,N_6959,N_5326);
or U8939 (N_8939,N_6978,N_5325);
or U8940 (N_8940,N_6381,N_5601);
nand U8941 (N_8941,N_6785,N_6658);
and U8942 (N_8942,N_5202,N_5818);
xnor U8943 (N_8943,N_7128,N_5825);
nor U8944 (N_8944,N_7149,N_5974);
nor U8945 (N_8945,N_5048,N_5356);
and U8946 (N_8946,N_7413,N_5320);
and U8947 (N_8947,N_5795,N_6892);
nand U8948 (N_8948,N_6757,N_5055);
nand U8949 (N_8949,N_7159,N_6162);
nand U8950 (N_8950,N_5662,N_5009);
or U8951 (N_8951,N_6611,N_5083);
or U8952 (N_8952,N_6605,N_6531);
and U8953 (N_8953,N_5705,N_6063);
or U8954 (N_8954,N_5390,N_5278);
and U8955 (N_8955,N_5854,N_6616);
or U8956 (N_8956,N_5890,N_6173);
nor U8957 (N_8957,N_5644,N_5064);
nand U8958 (N_8958,N_7065,N_5314);
and U8959 (N_8959,N_6735,N_6508);
or U8960 (N_8960,N_7331,N_7445);
nand U8961 (N_8961,N_6696,N_6569);
and U8962 (N_8962,N_5411,N_5585);
nor U8963 (N_8963,N_5123,N_7145);
and U8964 (N_8964,N_5628,N_5157);
and U8965 (N_8965,N_6520,N_6315);
nand U8966 (N_8966,N_5820,N_7316);
nor U8967 (N_8967,N_6076,N_6567);
nor U8968 (N_8968,N_6912,N_5789);
nand U8969 (N_8969,N_6159,N_5087);
or U8970 (N_8970,N_6915,N_5440);
nor U8971 (N_8971,N_5242,N_6540);
and U8972 (N_8972,N_6935,N_6029);
or U8973 (N_8973,N_5350,N_7127);
xnor U8974 (N_8974,N_6296,N_5517);
or U8975 (N_8975,N_7433,N_5914);
nand U8976 (N_8976,N_5624,N_7211);
nor U8977 (N_8977,N_6166,N_5399);
and U8978 (N_8978,N_7026,N_6040);
or U8979 (N_8979,N_6896,N_5658);
and U8980 (N_8980,N_7372,N_7098);
and U8981 (N_8981,N_6880,N_5706);
or U8982 (N_8982,N_7121,N_5417);
nor U8983 (N_8983,N_6595,N_7404);
or U8984 (N_8984,N_5516,N_5805);
nand U8985 (N_8985,N_7030,N_5163);
nor U8986 (N_8986,N_7480,N_5870);
nand U8987 (N_8987,N_5605,N_5443);
nand U8988 (N_8988,N_7099,N_6610);
nand U8989 (N_8989,N_6765,N_5293);
nand U8990 (N_8990,N_7220,N_5457);
and U8991 (N_8991,N_5996,N_6031);
and U8992 (N_8992,N_5125,N_6131);
and U8993 (N_8993,N_5310,N_5313);
nor U8994 (N_8994,N_6127,N_5293);
and U8995 (N_8995,N_5421,N_6567);
nand U8996 (N_8996,N_5603,N_5260);
nand U8997 (N_8997,N_5765,N_5805);
and U8998 (N_8998,N_5383,N_6077);
nand U8999 (N_8999,N_6950,N_5750);
or U9000 (N_9000,N_6160,N_6897);
nor U9001 (N_9001,N_5125,N_6635);
and U9002 (N_9002,N_6971,N_6297);
nor U9003 (N_9003,N_5030,N_7107);
nor U9004 (N_9004,N_5357,N_5365);
nor U9005 (N_9005,N_6091,N_5621);
nand U9006 (N_9006,N_7092,N_6635);
and U9007 (N_9007,N_5712,N_5733);
and U9008 (N_9008,N_5462,N_6006);
nor U9009 (N_9009,N_6616,N_5594);
nor U9010 (N_9010,N_5454,N_5948);
or U9011 (N_9011,N_5688,N_7382);
nand U9012 (N_9012,N_5403,N_7373);
nor U9013 (N_9013,N_7214,N_6089);
or U9014 (N_9014,N_5151,N_6097);
and U9015 (N_9015,N_6079,N_7046);
and U9016 (N_9016,N_6184,N_6344);
and U9017 (N_9017,N_5044,N_6722);
nor U9018 (N_9018,N_7182,N_6165);
nand U9019 (N_9019,N_7141,N_5055);
nor U9020 (N_9020,N_6623,N_5268);
and U9021 (N_9021,N_5431,N_5297);
nor U9022 (N_9022,N_5537,N_6496);
and U9023 (N_9023,N_5174,N_5883);
and U9024 (N_9024,N_6180,N_5782);
and U9025 (N_9025,N_7456,N_6923);
nand U9026 (N_9026,N_5165,N_7451);
or U9027 (N_9027,N_5954,N_5579);
nand U9028 (N_9028,N_5484,N_5481);
and U9029 (N_9029,N_6415,N_7168);
nor U9030 (N_9030,N_6239,N_5955);
nor U9031 (N_9031,N_7217,N_5646);
and U9032 (N_9032,N_6132,N_7427);
nor U9033 (N_9033,N_5153,N_6166);
nand U9034 (N_9034,N_5769,N_7081);
or U9035 (N_9035,N_7379,N_7232);
nor U9036 (N_9036,N_6997,N_6805);
nand U9037 (N_9037,N_5454,N_6034);
or U9038 (N_9038,N_5934,N_7013);
or U9039 (N_9039,N_6915,N_5191);
and U9040 (N_9040,N_5419,N_5473);
and U9041 (N_9041,N_6913,N_6666);
nor U9042 (N_9042,N_5402,N_5548);
nand U9043 (N_9043,N_6557,N_7083);
or U9044 (N_9044,N_5058,N_6451);
nor U9045 (N_9045,N_5998,N_5575);
and U9046 (N_9046,N_7029,N_6934);
nor U9047 (N_9047,N_6671,N_5830);
nor U9048 (N_9048,N_5292,N_5490);
nand U9049 (N_9049,N_5753,N_5447);
or U9050 (N_9050,N_7293,N_7330);
or U9051 (N_9051,N_5716,N_7089);
and U9052 (N_9052,N_6696,N_5004);
and U9053 (N_9053,N_5342,N_6215);
nor U9054 (N_9054,N_6346,N_7034);
nand U9055 (N_9055,N_5671,N_6080);
nor U9056 (N_9056,N_6095,N_6977);
nor U9057 (N_9057,N_6872,N_6322);
nor U9058 (N_9058,N_6619,N_7401);
or U9059 (N_9059,N_6129,N_5289);
and U9060 (N_9060,N_5356,N_6832);
and U9061 (N_9061,N_6992,N_6058);
and U9062 (N_9062,N_7009,N_5259);
nor U9063 (N_9063,N_7097,N_6136);
xor U9064 (N_9064,N_7350,N_6389);
nand U9065 (N_9065,N_6949,N_6426);
nand U9066 (N_9066,N_6586,N_5735);
nand U9067 (N_9067,N_6753,N_6553);
nor U9068 (N_9068,N_6821,N_5365);
nor U9069 (N_9069,N_5046,N_6654);
and U9070 (N_9070,N_6241,N_6514);
and U9071 (N_9071,N_5965,N_5598);
nand U9072 (N_9072,N_5933,N_6093);
and U9073 (N_9073,N_6706,N_7097);
nor U9074 (N_9074,N_6352,N_6073);
nor U9075 (N_9075,N_5368,N_6077);
or U9076 (N_9076,N_7145,N_6321);
nand U9077 (N_9077,N_6011,N_6300);
nor U9078 (N_9078,N_5330,N_6108);
nand U9079 (N_9079,N_6900,N_6452);
and U9080 (N_9080,N_7118,N_7243);
nor U9081 (N_9081,N_5355,N_7215);
and U9082 (N_9082,N_6928,N_5174);
nor U9083 (N_9083,N_5071,N_6154);
or U9084 (N_9084,N_7415,N_6080);
nor U9085 (N_9085,N_5995,N_7422);
nand U9086 (N_9086,N_7129,N_6518);
and U9087 (N_9087,N_5648,N_6429);
or U9088 (N_9088,N_6332,N_5342);
or U9089 (N_9089,N_5476,N_6671);
and U9090 (N_9090,N_5169,N_5362);
or U9091 (N_9091,N_6583,N_6866);
or U9092 (N_9092,N_5638,N_7483);
or U9093 (N_9093,N_5154,N_5765);
nor U9094 (N_9094,N_5430,N_7103);
nand U9095 (N_9095,N_6785,N_7121);
nor U9096 (N_9096,N_5186,N_5884);
nand U9097 (N_9097,N_6470,N_6586);
nor U9098 (N_9098,N_6241,N_5501);
or U9099 (N_9099,N_6056,N_5115);
nand U9100 (N_9100,N_5397,N_6292);
or U9101 (N_9101,N_6152,N_7232);
nand U9102 (N_9102,N_6658,N_6609);
or U9103 (N_9103,N_5439,N_6078);
or U9104 (N_9104,N_5175,N_5404);
nand U9105 (N_9105,N_5231,N_5818);
nand U9106 (N_9106,N_7304,N_6189);
or U9107 (N_9107,N_5323,N_6001);
and U9108 (N_9108,N_6462,N_6661);
nor U9109 (N_9109,N_7279,N_6931);
and U9110 (N_9110,N_5640,N_5666);
xnor U9111 (N_9111,N_5561,N_5320);
nor U9112 (N_9112,N_6167,N_5042);
and U9113 (N_9113,N_6401,N_6917);
nor U9114 (N_9114,N_5590,N_5617);
nand U9115 (N_9115,N_5971,N_6986);
nor U9116 (N_9116,N_6199,N_6240);
nand U9117 (N_9117,N_7487,N_5687);
or U9118 (N_9118,N_5337,N_6584);
nor U9119 (N_9119,N_5939,N_5699);
or U9120 (N_9120,N_7072,N_6060);
nor U9121 (N_9121,N_6587,N_6000);
and U9122 (N_9122,N_6066,N_7353);
and U9123 (N_9123,N_5227,N_7446);
and U9124 (N_9124,N_5938,N_5515);
nand U9125 (N_9125,N_6597,N_6361);
nor U9126 (N_9126,N_7440,N_7487);
or U9127 (N_9127,N_7327,N_6461);
or U9128 (N_9128,N_5890,N_5214);
nor U9129 (N_9129,N_6094,N_6853);
nor U9130 (N_9130,N_6904,N_6628);
and U9131 (N_9131,N_6942,N_7339);
nor U9132 (N_9132,N_7085,N_7409);
or U9133 (N_9133,N_6645,N_6392);
or U9134 (N_9134,N_5241,N_7158);
nor U9135 (N_9135,N_7239,N_6468);
nand U9136 (N_9136,N_5925,N_6433);
or U9137 (N_9137,N_6778,N_7282);
and U9138 (N_9138,N_7436,N_6912);
or U9139 (N_9139,N_7365,N_7060);
and U9140 (N_9140,N_6861,N_7206);
xnor U9141 (N_9141,N_5839,N_6186);
nor U9142 (N_9142,N_5837,N_5801);
nor U9143 (N_9143,N_6195,N_7218);
nor U9144 (N_9144,N_7128,N_5110);
nor U9145 (N_9145,N_7401,N_6550);
nand U9146 (N_9146,N_5007,N_6177);
xnor U9147 (N_9147,N_6678,N_6306);
nor U9148 (N_9148,N_6059,N_6153);
or U9149 (N_9149,N_7301,N_5431);
and U9150 (N_9150,N_5208,N_5747);
or U9151 (N_9151,N_5644,N_6531);
or U9152 (N_9152,N_7086,N_5534);
nand U9153 (N_9153,N_7298,N_6296);
nor U9154 (N_9154,N_5362,N_6516);
or U9155 (N_9155,N_6943,N_5595);
and U9156 (N_9156,N_5540,N_5765);
and U9157 (N_9157,N_6234,N_5762);
and U9158 (N_9158,N_6876,N_6506);
nand U9159 (N_9159,N_5994,N_6105);
xnor U9160 (N_9160,N_6797,N_7203);
nor U9161 (N_9161,N_5599,N_5675);
and U9162 (N_9162,N_5577,N_7435);
nand U9163 (N_9163,N_5744,N_5825);
and U9164 (N_9164,N_6413,N_6828);
or U9165 (N_9165,N_6951,N_6428);
or U9166 (N_9166,N_5955,N_6360);
and U9167 (N_9167,N_6299,N_6409);
and U9168 (N_9168,N_7226,N_5814);
nand U9169 (N_9169,N_7206,N_5035);
and U9170 (N_9170,N_6133,N_6706);
nand U9171 (N_9171,N_5746,N_5683);
nor U9172 (N_9172,N_7094,N_6083);
and U9173 (N_9173,N_6959,N_7375);
and U9174 (N_9174,N_5035,N_7328);
and U9175 (N_9175,N_6865,N_5853);
and U9176 (N_9176,N_5764,N_6682);
nand U9177 (N_9177,N_5254,N_6100);
and U9178 (N_9178,N_6348,N_5858);
nand U9179 (N_9179,N_5950,N_6111);
xnor U9180 (N_9180,N_5344,N_5497);
nand U9181 (N_9181,N_5194,N_7062);
or U9182 (N_9182,N_6352,N_6790);
and U9183 (N_9183,N_7056,N_6549);
nor U9184 (N_9184,N_7314,N_5221);
or U9185 (N_9185,N_6327,N_5348);
nor U9186 (N_9186,N_7149,N_6500);
nor U9187 (N_9187,N_5071,N_7216);
nor U9188 (N_9188,N_6905,N_7331);
nand U9189 (N_9189,N_5585,N_5311);
and U9190 (N_9190,N_5336,N_6840);
or U9191 (N_9191,N_6167,N_5153);
and U9192 (N_9192,N_7134,N_5294);
or U9193 (N_9193,N_7415,N_6815);
nor U9194 (N_9194,N_6771,N_5086);
or U9195 (N_9195,N_6511,N_7268);
and U9196 (N_9196,N_6503,N_6898);
nand U9197 (N_9197,N_5077,N_7340);
nor U9198 (N_9198,N_6519,N_6848);
nand U9199 (N_9199,N_5145,N_5848);
nand U9200 (N_9200,N_6430,N_5886);
nor U9201 (N_9201,N_6164,N_5935);
xnor U9202 (N_9202,N_5672,N_6191);
nor U9203 (N_9203,N_7080,N_6257);
nor U9204 (N_9204,N_7287,N_5913);
nor U9205 (N_9205,N_5411,N_6058);
nor U9206 (N_9206,N_5584,N_6307);
or U9207 (N_9207,N_5386,N_6267);
or U9208 (N_9208,N_5164,N_5174);
nand U9209 (N_9209,N_6504,N_5180);
or U9210 (N_9210,N_6061,N_5687);
and U9211 (N_9211,N_7370,N_7268);
or U9212 (N_9212,N_7056,N_6678);
nand U9213 (N_9213,N_6859,N_6963);
nor U9214 (N_9214,N_5923,N_6633);
nor U9215 (N_9215,N_7162,N_7361);
and U9216 (N_9216,N_6673,N_7048);
nor U9217 (N_9217,N_6440,N_6427);
or U9218 (N_9218,N_6387,N_6493);
or U9219 (N_9219,N_6450,N_5449);
and U9220 (N_9220,N_5534,N_5640);
or U9221 (N_9221,N_6515,N_7415);
and U9222 (N_9222,N_6065,N_5268);
nand U9223 (N_9223,N_7195,N_5265);
nor U9224 (N_9224,N_6354,N_5908);
and U9225 (N_9225,N_5793,N_7350);
nor U9226 (N_9226,N_5571,N_6282);
or U9227 (N_9227,N_5327,N_5174);
nor U9228 (N_9228,N_5575,N_6626);
nand U9229 (N_9229,N_7209,N_6381);
nor U9230 (N_9230,N_6536,N_6998);
nor U9231 (N_9231,N_6008,N_6377);
and U9232 (N_9232,N_5756,N_6441);
nor U9233 (N_9233,N_6787,N_6884);
and U9234 (N_9234,N_6898,N_6980);
nor U9235 (N_9235,N_6339,N_5549);
nand U9236 (N_9236,N_5626,N_6680);
and U9237 (N_9237,N_6190,N_5295);
nand U9238 (N_9238,N_5813,N_7242);
xnor U9239 (N_9239,N_6698,N_5109);
or U9240 (N_9240,N_5704,N_6828);
or U9241 (N_9241,N_6636,N_6016);
nand U9242 (N_9242,N_6856,N_5707);
nand U9243 (N_9243,N_6203,N_5211);
nor U9244 (N_9244,N_5852,N_6173);
nand U9245 (N_9245,N_6125,N_7286);
nand U9246 (N_9246,N_5394,N_5587);
and U9247 (N_9247,N_6199,N_5135);
nor U9248 (N_9248,N_6787,N_5643);
nor U9249 (N_9249,N_6053,N_5680);
nor U9250 (N_9250,N_5814,N_5790);
or U9251 (N_9251,N_7407,N_5814);
and U9252 (N_9252,N_5075,N_6565);
and U9253 (N_9253,N_5140,N_7199);
and U9254 (N_9254,N_6950,N_5148);
nand U9255 (N_9255,N_6269,N_7276);
and U9256 (N_9256,N_5996,N_6796);
and U9257 (N_9257,N_5010,N_5315);
and U9258 (N_9258,N_6716,N_7107);
nand U9259 (N_9259,N_5795,N_7492);
nor U9260 (N_9260,N_5265,N_7090);
and U9261 (N_9261,N_5376,N_6577);
and U9262 (N_9262,N_6715,N_5709);
nand U9263 (N_9263,N_6373,N_7421);
nand U9264 (N_9264,N_6811,N_7332);
and U9265 (N_9265,N_6182,N_7494);
and U9266 (N_9266,N_6641,N_5442);
and U9267 (N_9267,N_6478,N_7463);
or U9268 (N_9268,N_7350,N_5795);
and U9269 (N_9269,N_6021,N_6805);
xor U9270 (N_9270,N_7059,N_5409);
or U9271 (N_9271,N_5259,N_7046);
and U9272 (N_9272,N_7078,N_7327);
nor U9273 (N_9273,N_6774,N_6320);
nand U9274 (N_9274,N_5527,N_7466);
or U9275 (N_9275,N_5919,N_7468);
nand U9276 (N_9276,N_5757,N_5831);
and U9277 (N_9277,N_5219,N_7409);
nand U9278 (N_9278,N_6905,N_6509);
nor U9279 (N_9279,N_7328,N_5387);
nand U9280 (N_9280,N_6986,N_6874);
nand U9281 (N_9281,N_6140,N_6693);
nand U9282 (N_9282,N_5051,N_5789);
nand U9283 (N_9283,N_5129,N_7317);
or U9284 (N_9284,N_5170,N_7433);
nand U9285 (N_9285,N_6673,N_5585);
nand U9286 (N_9286,N_5167,N_6460);
nand U9287 (N_9287,N_5293,N_6803);
nor U9288 (N_9288,N_6377,N_5062);
and U9289 (N_9289,N_5718,N_6859);
nand U9290 (N_9290,N_6641,N_6330);
nor U9291 (N_9291,N_5785,N_6244);
nand U9292 (N_9292,N_5102,N_6840);
nor U9293 (N_9293,N_6848,N_5938);
nand U9294 (N_9294,N_6660,N_5390);
nor U9295 (N_9295,N_5369,N_6046);
xor U9296 (N_9296,N_5834,N_6729);
and U9297 (N_9297,N_7024,N_5361);
nand U9298 (N_9298,N_5256,N_6638);
and U9299 (N_9299,N_7036,N_7196);
and U9300 (N_9300,N_6190,N_5717);
nor U9301 (N_9301,N_7131,N_6286);
and U9302 (N_9302,N_5566,N_5034);
and U9303 (N_9303,N_6536,N_5455);
nand U9304 (N_9304,N_5189,N_5209);
and U9305 (N_9305,N_6944,N_7370);
nand U9306 (N_9306,N_6127,N_6814);
nand U9307 (N_9307,N_6514,N_5478);
or U9308 (N_9308,N_6431,N_6874);
and U9309 (N_9309,N_5388,N_6759);
and U9310 (N_9310,N_5351,N_5676);
and U9311 (N_9311,N_6075,N_6012);
and U9312 (N_9312,N_6424,N_5031);
nor U9313 (N_9313,N_7480,N_7179);
nor U9314 (N_9314,N_5978,N_7075);
nand U9315 (N_9315,N_5848,N_5914);
nor U9316 (N_9316,N_7053,N_5768);
nor U9317 (N_9317,N_6629,N_7180);
nor U9318 (N_9318,N_6645,N_6042);
or U9319 (N_9319,N_6698,N_7469);
xor U9320 (N_9320,N_6015,N_7112);
or U9321 (N_9321,N_7207,N_5687);
or U9322 (N_9322,N_6368,N_5161);
and U9323 (N_9323,N_7214,N_6861);
or U9324 (N_9324,N_5915,N_6365);
nor U9325 (N_9325,N_7234,N_7100);
nand U9326 (N_9326,N_5007,N_5436);
and U9327 (N_9327,N_6015,N_7242);
nor U9328 (N_9328,N_5809,N_6692);
nor U9329 (N_9329,N_5101,N_5261);
or U9330 (N_9330,N_5874,N_5377);
and U9331 (N_9331,N_5961,N_5823);
and U9332 (N_9332,N_6023,N_5977);
and U9333 (N_9333,N_6202,N_6204);
nor U9334 (N_9334,N_5995,N_5838);
or U9335 (N_9335,N_5625,N_6132);
and U9336 (N_9336,N_5431,N_6429);
nand U9337 (N_9337,N_5231,N_5892);
nand U9338 (N_9338,N_5758,N_5534);
nor U9339 (N_9339,N_6256,N_5662);
nor U9340 (N_9340,N_6645,N_7262);
or U9341 (N_9341,N_7442,N_5610);
or U9342 (N_9342,N_5040,N_5573);
or U9343 (N_9343,N_5449,N_7009);
nor U9344 (N_9344,N_5059,N_6932);
nor U9345 (N_9345,N_6898,N_5995);
nor U9346 (N_9346,N_7088,N_6884);
and U9347 (N_9347,N_6706,N_7080);
nand U9348 (N_9348,N_6017,N_5489);
nor U9349 (N_9349,N_6503,N_5362);
nor U9350 (N_9350,N_6723,N_7431);
nand U9351 (N_9351,N_5297,N_7450);
nor U9352 (N_9352,N_7350,N_7311);
nand U9353 (N_9353,N_6465,N_7199);
or U9354 (N_9354,N_5788,N_6768);
nand U9355 (N_9355,N_7371,N_6102);
nor U9356 (N_9356,N_6369,N_7463);
nand U9357 (N_9357,N_6502,N_6203);
nor U9358 (N_9358,N_7043,N_5785);
and U9359 (N_9359,N_6305,N_5210);
nor U9360 (N_9360,N_5462,N_6924);
nor U9361 (N_9361,N_5945,N_7364);
and U9362 (N_9362,N_7476,N_5266);
nand U9363 (N_9363,N_6991,N_6195);
and U9364 (N_9364,N_5218,N_5322);
nor U9365 (N_9365,N_5367,N_6716);
and U9366 (N_9366,N_5838,N_6720);
or U9367 (N_9367,N_5127,N_5269);
xor U9368 (N_9368,N_5885,N_6443);
or U9369 (N_9369,N_5316,N_7198);
nor U9370 (N_9370,N_5392,N_5402);
nor U9371 (N_9371,N_5250,N_6411);
and U9372 (N_9372,N_7419,N_6194);
xor U9373 (N_9373,N_6380,N_5893);
nor U9374 (N_9374,N_6847,N_7113);
xor U9375 (N_9375,N_5729,N_5184);
nor U9376 (N_9376,N_5089,N_5502);
nand U9377 (N_9377,N_5525,N_5861);
and U9378 (N_9378,N_6070,N_6703);
nor U9379 (N_9379,N_5248,N_5727);
nand U9380 (N_9380,N_7408,N_6725);
nand U9381 (N_9381,N_7322,N_7217);
nand U9382 (N_9382,N_7322,N_7081);
nor U9383 (N_9383,N_5716,N_6926);
and U9384 (N_9384,N_5404,N_5557);
nor U9385 (N_9385,N_5810,N_7418);
or U9386 (N_9386,N_5162,N_6547);
nand U9387 (N_9387,N_6393,N_5826);
nor U9388 (N_9388,N_7099,N_5108);
and U9389 (N_9389,N_6431,N_6272);
and U9390 (N_9390,N_6537,N_6134);
and U9391 (N_9391,N_6229,N_6096);
and U9392 (N_9392,N_7393,N_6836);
and U9393 (N_9393,N_5717,N_5989);
and U9394 (N_9394,N_5351,N_6757);
nand U9395 (N_9395,N_6698,N_5096);
and U9396 (N_9396,N_5824,N_6236);
or U9397 (N_9397,N_6693,N_5479);
or U9398 (N_9398,N_6603,N_5454);
and U9399 (N_9399,N_7173,N_7358);
nand U9400 (N_9400,N_7463,N_7330);
nor U9401 (N_9401,N_5235,N_7419);
nand U9402 (N_9402,N_7496,N_7250);
nand U9403 (N_9403,N_6993,N_5555);
or U9404 (N_9404,N_5257,N_6301);
xor U9405 (N_9405,N_5117,N_6343);
nand U9406 (N_9406,N_5783,N_5392);
or U9407 (N_9407,N_5201,N_7373);
or U9408 (N_9408,N_5161,N_5722);
and U9409 (N_9409,N_6136,N_7217);
nor U9410 (N_9410,N_7242,N_7482);
nor U9411 (N_9411,N_5698,N_6246);
or U9412 (N_9412,N_6446,N_5925);
nand U9413 (N_9413,N_6736,N_7494);
nand U9414 (N_9414,N_5218,N_6469);
nand U9415 (N_9415,N_5947,N_6855);
and U9416 (N_9416,N_6851,N_5808);
or U9417 (N_9417,N_7194,N_5307);
or U9418 (N_9418,N_6288,N_5983);
nand U9419 (N_9419,N_6228,N_5211);
and U9420 (N_9420,N_5522,N_7446);
or U9421 (N_9421,N_5921,N_5494);
nor U9422 (N_9422,N_7108,N_6222);
or U9423 (N_9423,N_6014,N_6651);
nand U9424 (N_9424,N_7111,N_6761);
or U9425 (N_9425,N_6136,N_6153);
and U9426 (N_9426,N_6481,N_7378);
and U9427 (N_9427,N_7000,N_5057);
or U9428 (N_9428,N_7423,N_7079);
or U9429 (N_9429,N_6710,N_5675);
nor U9430 (N_9430,N_6263,N_7347);
nor U9431 (N_9431,N_6231,N_5445);
nor U9432 (N_9432,N_6614,N_6093);
and U9433 (N_9433,N_5745,N_6783);
nand U9434 (N_9434,N_6725,N_5033);
or U9435 (N_9435,N_5025,N_5366);
or U9436 (N_9436,N_7235,N_6646);
and U9437 (N_9437,N_5878,N_6223);
and U9438 (N_9438,N_5296,N_6953);
nand U9439 (N_9439,N_6639,N_5811);
nor U9440 (N_9440,N_5253,N_5904);
nor U9441 (N_9441,N_7146,N_5049);
nand U9442 (N_9442,N_7386,N_7160);
nand U9443 (N_9443,N_6882,N_6395);
and U9444 (N_9444,N_5218,N_5389);
xnor U9445 (N_9445,N_5491,N_7376);
or U9446 (N_9446,N_5158,N_6083);
nor U9447 (N_9447,N_6063,N_5368);
nand U9448 (N_9448,N_6081,N_5490);
and U9449 (N_9449,N_7284,N_5513);
nor U9450 (N_9450,N_5425,N_6053);
nand U9451 (N_9451,N_6351,N_6856);
and U9452 (N_9452,N_5061,N_6169);
and U9453 (N_9453,N_6031,N_5892);
nand U9454 (N_9454,N_7465,N_6852);
nand U9455 (N_9455,N_5038,N_5769);
or U9456 (N_9456,N_6828,N_5242);
and U9457 (N_9457,N_6529,N_7019);
or U9458 (N_9458,N_5109,N_6257);
or U9459 (N_9459,N_5890,N_5074);
nand U9460 (N_9460,N_6156,N_5804);
nand U9461 (N_9461,N_7320,N_5064);
or U9462 (N_9462,N_6873,N_6750);
nor U9463 (N_9463,N_5766,N_7160);
or U9464 (N_9464,N_6070,N_6875);
or U9465 (N_9465,N_6398,N_6928);
or U9466 (N_9466,N_7275,N_5593);
or U9467 (N_9467,N_5663,N_5489);
and U9468 (N_9468,N_5261,N_5029);
and U9469 (N_9469,N_6071,N_5036);
nand U9470 (N_9470,N_5307,N_6423);
or U9471 (N_9471,N_7144,N_5981);
or U9472 (N_9472,N_6443,N_6649);
and U9473 (N_9473,N_6916,N_7419);
nor U9474 (N_9474,N_6237,N_5669);
xnor U9475 (N_9475,N_5862,N_5812);
nand U9476 (N_9476,N_5595,N_6007);
nor U9477 (N_9477,N_7488,N_6984);
xor U9478 (N_9478,N_5102,N_6058);
and U9479 (N_9479,N_6197,N_5786);
and U9480 (N_9480,N_6427,N_6534);
nor U9481 (N_9481,N_6543,N_6327);
or U9482 (N_9482,N_5805,N_7085);
nand U9483 (N_9483,N_5824,N_6303);
nor U9484 (N_9484,N_5721,N_6880);
and U9485 (N_9485,N_5642,N_6385);
nor U9486 (N_9486,N_5583,N_7240);
or U9487 (N_9487,N_6143,N_5936);
nand U9488 (N_9488,N_5845,N_6246);
nor U9489 (N_9489,N_6895,N_6328);
and U9490 (N_9490,N_6906,N_5791);
and U9491 (N_9491,N_6558,N_6457);
nor U9492 (N_9492,N_6733,N_7475);
and U9493 (N_9493,N_5487,N_6727);
nor U9494 (N_9494,N_6977,N_6753);
or U9495 (N_9495,N_5549,N_6556);
nand U9496 (N_9496,N_6271,N_6289);
nor U9497 (N_9497,N_6440,N_6784);
nand U9498 (N_9498,N_5075,N_6829);
or U9499 (N_9499,N_6454,N_7228);
xnor U9500 (N_9500,N_6191,N_6929);
and U9501 (N_9501,N_7084,N_5959);
nor U9502 (N_9502,N_5506,N_5388);
and U9503 (N_9503,N_6223,N_5962);
nand U9504 (N_9504,N_5923,N_6382);
and U9505 (N_9505,N_5230,N_6462);
nor U9506 (N_9506,N_5491,N_7486);
nand U9507 (N_9507,N_6862,N_6803);
or U9508 (N_9508,N_7201,N_7125);
nand U9509 (N_9509,N_6095,N_6758);
nor U9510 (N_9510,N_5400,N_5640);
nor U9511 (N_9511,N_6832,N_6417);
and U9512 (N_9512,N_6019,N_6948);
nand U9513 (N_9513,N_6762,N_5241);
nor U9514 (N_9514,N_5444,N_7489);
or U9515 (N_9515,N_6435,N_6409);
nand U9516 (N_9516,N_5971,N_6219);
xor U9517 (N_9517,N_5580,N_6948);
or U9518 (N_9518,N_6550,N_6029);
nor U9519 (N_9519,N_5019,N_5171);
nor U9520 (N_9520,N_5628,N_5622);
or U9521 (N_9521,N_5592,N_6733);
nor U9522 (N_9522,N_6846,N_5759);
nand U9523 (N_9523,N_6809,N_6228);
nand U9524 (N_9524,N_6929,N_7299);
nand U9525 (N_9525,N_6017,N_5746);
and U9526 (N_9526,N_5486,N_5849);
nand U9527 (N_9527,N_7219,N_7103);
nand U9528 (N_9528,N_5382,N_6537);
and U9529 (N_9529,N_5490,N_6678);
nand U9530 (N_9530,N_6780,N_7314);
and U9531 (N_9531,N_5659,N_5805);
and U9532 (N_9532,N_5653,N_6014);
and U9533 (N_9533,N_5316,N_7110);
or U9534 (N_9534,N_6649,N_7383);
and U9535 (N_9535,N_5551,N_7167);
nand U9536 (N_9536,N_5052,N_7191);
nor U9537 (N_9537,N_5006,N_5138);
nor U9538 (N_9538,N_7047,N_5721);
nor U9539 (N_9539,N_5121,N_5221);
nor U9540 (N_9540,N_5674,N_6601);
or U9541 (N_9541,N_7477,N_7178);
xor U9542 (N_9542,N_6676,N_6076);
nand U9543 (N_9543,N_5487,N_5819);
nor U9544 (N_9544,N_6025,N_5647);
or U9545 (N_9545,N_5441,N_6265);
nand U9546 (N_9546,N_6720,N_7191);
nor U9547 (N_9547,N_6821,N_5680);
and U9548 (N_9548,N_5632,N_6633);
or U9549 (N_9549,N_5987,N_5678);
nor U9550 (N_9550,N_5156,N_5557);
and U9551 (N_9551,N_6464,N_5980);
nor U9552 (N_9552,N_5425,N_5505);
and U9553 (N_9553,N_5099,N_6100);
xor U9554 (N_9554,N_6433,N_5930);
or U9555 (N_9555,N_5300,N_6538);
or U9556 (N_9556,N_6739,N_7397);
xnor U9557 (N_9557,N_6599,N_5274);
nand U9558 (N_9558,N_6914,N_6735);
or U9559 (N_9559,N_6471,N_6834);
or U9560 (N_9560,N_5423,N_5098);
or U9561 (N_9561,N_5043,N_5897);
or U9562 (N_9562,N_5221,N_5194);
nand U9563 (N_9563,N_6137,N_7239);
nand U9564 (N_9564,N_6919,N_5459);
nand U9565 (N_9565,N_5870,N_5375);
or U9566 (N_9566,N_5809,N_5023);
xnor U9567 (N_9567,N_6659,N_5894);
nand U9568 (N_9568,N_6280,N_5873);
nor U9569 (N_9569,N_5345,N_6339);
nor U9570 (N_9570,N_6648,N_5707);
nor U9571 (N_9571,N_5555,N_6275);
or U9572 (N_9572,N_5909,N_5853);
and U9573 (N_9573,N_6108,N_5266);
and U9574 (N_9574,N_5233,N_6363);
nor U9575 (N_9575,N_7342,N_5574);
nor U9576 (N_9576,N_5439,N_6912);
nand U9577 (N_9577,N_7337,N_5648);
nor U9578 (N_9578,N_5509,N_5757);
or U9579 (N_9579,N_5037,N_7253);
nor U9580 (N_9580,N_7465,N_6900);
and U9581 (N_9581,N_6906,N_6895);
nor U9582 (N_9582,N_7430,N_5609);
or U9583 (N_9583,N_6160,N_6751);
nor U9584 (N_9584,N_5283,N_5785);
or U9585 (N_9585,N_7056,N_6418);
and U9586 (N_9586,N_6859,N_7185);
nand U9587 (N_9587,N_5111,N_5433);
nor U9588 (N_9588,N_5446,N_5166);
nor U9589 (N_9589,N_5980,N_7181);
or U9590 (N_9590,N_7443,N_6879);
and U9591 (N_9591,N_6114,N_6492);
nor U9592 (N_9592,N_7370,N_6942);
nor U9593 (N_9593,N_6878,N_7436);
or U9594 (N_9594,N_7194,N_7073);
and U9595 (N_9595,N_5415,N_5066);
nor U9596 (N_9596,N_5277,N_7356);
nand U9597 (N_9597,N_6870,N_7280);
and U9598 (N_9598,N_6662,N_6454);
and U9599 (N_9599,N_6340,N_7009);
nand U9600 (N_9600,N_6231,N_6417);
nand U9601 (N_9601,N_5153,N_7275);
or U9602 (N_9602,N_6712,N_6055);
or U9603 (N_9603,N_6624,N_7159);
nor U9604 (N_9604,N_6771,N_5212);
nand U9605 (N_9605,N_7289,N_5676);
nor U9606 (N_9606,N_5177,N_6817);
and U9607 (N_9607,N_6563,N_6144);
and U9608 (N_9608,N_6090,N_5689);
nor U9609 (N_9609,N_6041,N_5916);
nor U9610 (N_9610,N_6180,N_5527);
nand U9611 (N_9611,N_6119,N_7243);
and U9612 (N_9612,N_5546,N_6187);
nor U9613 (N_9613,N_5109,N_6091);
and U9614 (N_9614,N_6001,N_6794);
nand U9615 (N_9615,N_5901,N_6528);
nor U9616 (N_9616,N_6373,N_5518);
and U9617 (N_9617,N_6004,N_7423);
or U9618 (N_9618,N_6837,N_7389);
xor U9619 (N_9619,N_6979,N_7453);
or U9620 (N_9620,N_6050,N_5123);
nor U9621 (N_9621,N_5945,N_5376);
xnor U9622 (N_9622,N_6902,N_5444);
nor U9623 (N_9623,N_7159,N_5606);
or U9624 (N_9624,N_6380,N_5451);
nor U9625 (N_9625,N_5456,N_6955);
nor U9626 (N_9626,N_5901,N_5298);
and U9627 (N_9627,N_6903,N_5279);
nand U9628 (N_9628,N_7189,N_6655);
and U9629 (N_9629,N_5339,N_7193);
and U9630 (N_9630,N_6074,N_5601);
or U9631 (N_9631,N_6255,N_6799);
and U9632 (N_9632,N_5262,N_5523);
and U9633 (N_9633,N_5027,N_7142);
nor U9634 (N_9634,N_6196,N_6891);
nand U9635 (N_9635,N_5999,N_7403);
and U9636 (N_9636,N_5852,N_5620);
or U9637 (N_9637,N_6625,N_5718);
and U9638 (N_9638,N_5812,N_7445);
nand U9639 (N_9639,N_6586,N_6503);
or U9640 (N_9640,N_5268,N_7189);
or U9641 (N_9641,N_5814,N_6317);
and U9642 (N_9642,N_7133,N_6089);
nand U9643 (N_9643,N_7270,N_5323);
nor U9644 (N_9644,N_6022,N_5117);
nor U9645 (N_9645,N_5772,N_5098);
or U9646 (N_9646,N_6837,N_5674);
or U9647 (N_9647,N_5159,N_5454);
nor U9648 (N_9648,N_5688,N_6619);
nor U9649 (N_9649,N_5077,N_5225);
and U9650 (N_9650,N_5993,N_6411);
nand U9651 (N_9651,N_6524,N_5851);
nand U9652 (N_9652,N_5610,N_6166);
nor U9653 (N_9653,N_5550,N_5744);
or U9654 (N_9654,N_6933,N_7173);
nor U9655 (N_9655,N_7163,N_5768);
nand U9656 (N_9656,N_5743,N_5904);
nor U9657 (N_9657,N_5954,N_6584);
and U9658 (N_9658,N_5203,N_6923);
or U9659 (N_9659,N_6712,N_5856);
and U9660 (N_9660,N_5151,N_7404);
or U9661 (N_9661,N_7002,N_6499);
and U9662 (N_9662,N_6582,N_6516);
nor U9663 (N_9663,N_7066,N_6564);
nand U9664 (N_9664,N_5219,N_5262);
nand U9665 (N_9665,N_5198,N_5420);
nand U9666 (N_9666,N_5510,N_5877);
and U9667 (N_9667,N_6882,N_6598);
nor U9668 (N_9668,N_5548,N_6824);
xor U9669 (N_9669,N_7155,N_7357);
nor U9670 (N_9670,N_7290,N_7032);
nor U9671 (N_9671,N_7288,N_6625);
nand U9672 (N_9672,N_5286,N_6750);
and U9673 (N_9673,N_7494,N_6410);
and U9674 (N_9674,N_5045,N_5289);
or U9675 (N_9675,N_7100,N_6899);
and U9676 (N_9676,N_6198,N_5977);
nand U9677 (N_9677,N_7086,N_5162);
nand U9678 (N_9678,N_6915,N_7355);
or U9679 (N_9679,N_7336,N_5291);
or U9680 (N_9680,N_6055,N_5222);
nor U9681 (N_9681,N_7021,N_6833);
and U9682 (N_9682,N_6052,N_7152);
and U9683 (N_9683,N_5105,N_5949);
or U9684 (N_9684,N_5400,N_5537);
nand U9685 (N_9685,N_6531,N_6472);
nand U9686 (N_9686,N_5745,N_5367);
and U9687 (N_9687,N_7427,N_6149);
or U9688 (N_9688,N_5920,N_6466);
or U9689 (N_9689,N_6388,N_6613);
nor U9690 (N_9690,N_5977,N_6415);
nor U9691 (N_9691,N_5665,N_7282);
nor U9692 (N_9692,N_5047,N_5799);
or U9693 (N_9693,N_6646,N_7486);
nor U9694 (N_9694,N_6574,N_6332);
or U9695 (N_9695,N_6256,N_6039);
and U9696 (N_9696,N_7127,N_6864);
nor U9697 (N_9697,N_5005,N_5364);
or U9698 (N_9698,N_7481,N_6467);
nand U9699 (N_9699,N_5511,N_5103);
nand U9700 (N_9700,N_5638,N_6432);
nor U9701 (N_9701,N_7414,N_7390);
nand U9702 (N_9702,N_6814,N_6832);
or U9703 (N_9703,N_6212,N_5643);
nor U9704 (N_9704,N_5028,N_5997);
and U9705 (N_9705,N_5192,N_6705);
and U9706 (N_9706,N_5044,N_5019);
nor U9707 (N_9707,N_6627,N_6456);
nand U9708 (N_9708,N_7316,N_7301);
nor U9709 (N_9709,N_6765,N_5832);
nand U9710 (N_9710,N_5080,N_6753);
or U9711 (N_9711,N_6274,N_7058);
or U9712 (N_9712,N_6813,N_6083);
or U9713 (N_9713,N_5429,N_5082);
nor U9714 (N_9714,N_6299,N_6839);
or U9715 (N_9715,N_5773,N_5127);
nor U9716 (N_9716,N_5505,N_5233);
and U9717 (N_9717,N_5679,N_5472);
nor U9718 (N_9718,N_7017,N_5455);
and U9719 (N_9719,N_5584,N_7209);
or U9720 (N_9720,N_7480,N_5174);
nor U9721 (N_9721,N_6491,N_7009);
nand U9722 (N_9722,N_5097,N_7342);
nor U9723 (N_9723,N_6276,N_5363);
or U9724 (N_9724,N_6361,N_5177);
nor U9725 (N_9725,N_7050,N_5191);
and U9726 (N_9726,N_6148,N_6176);
nor U9727 (N_9727,N_7335,N_7304);
nand U9728 (N_9728,N_6423,N_5065);
or U9729 (N_9729,N_7260,N_6514);
and U9730 (N_9730,N_5725,N_6472);
and U9731 (N_9731,N_5011,N_6487);
nor U9732 (N_9732,N_6982,N_7446);
nand U9733 (N_9733,N_6613,N_5041);
nor U9734 (N_9734,N_7375,N_6260);
xor U9735 (N_9735,N_6005,N_7021);
nand U9736 (N_9736,N_6749,N_6615);
or U9737 (N_9737,N_6954,N_7226);
nand U9738 (N_9738,N_5018,N_6702);
nor U9739 (N_9739,N_6002,N_7119);
and U9740 (N_9740,N_5626,N_5417);
and U9741 (N_9741,N_5291,N_7298);
or U9742 (N_9742,N_6293,N_5938);
nor U9743 (N_9743,N_7053,N_6665);
nor U9744 (N_9744,N_5862,N_7288);
nor U9745 (N_9745,N_5426,N_5515);
or U9746 (N_9746,N_7294,N_6521);
nand U9747 (N_9747,N_6326,N_6437);
or U9748 (N_9748,N_5288,N_5076);
and U9749 (N_9749,N_5630,N_5988);
nor U9750 (N_9750,N_5474,N_5653);
xor U9751 (N_9751,N_6809,N_5095);
or U9752 (N_9752,N_6443,N_6404);
nand U9753 (N_9753,N_6012,N_5670);
nand U9754 (N_9754,N_7278,N_6992);
or U9755 (N_9755,N_5344,N_6426);
and U9756 (N_9756,N_5653,N_7176);
nand U9757 (N_9757,N_7217,N_6477);
or U9758 (N_9758,N_5483,N_6011);
or U9759 (N_9759,N_7161,N_6286);
nand U9760 (N_9760,N_5345,N_5169);
nand U9761 (N_9761,N_5228,N_6570);
nor U9762 (N_9762,N_7207,N_7313);
and U9763 (N_9763,N_7323,N_6101);
xor U9764 (N_9764,N_5921,N_5428);
nor U9765 (N_9765,N_7456,N_5757);
nor U9766 (N_9766,N_6438,N_6227);
or U9767 (N_9767,N_5853,N_6874);
nor U9768 (N_9768,N_5521,N_6156);
or U9769 (N_9769,N_5084,N_6344);
nand U9770 (N_9770,N_7468,N_7008);
nand U9771 (N_9771,N_6897,N_5580);
and U9772 (N_9772,N_5891,N_6265);
nor U9773 (N_9773,N_5628,N_5635);
nor U9774 (N_9774,N_7288,N_6551);
xnor U9775 (N_9775,N_6251,N_5752);
nand U9776 (N_9776,N_7409,N_6532);
nand U9777 (N_9777,N_7116,N_7039);
and U9778 (N_9778,N_6447,N_7375);
xnor U9779 (N_9779,N_6445,N_6229);
or U9780 (N_9780,N_6859,N_5250);
nand U9781 (N_9781,N_6235,N_6156);
nand U9782 (N_9782,N_5056,N_6711);
nand U9783 (N_9783,N_5591,N_6174);
and U9784 (N_9784,N_6625,N_7033);
nand U9785 (N_9785,N_6855,N_6980);
or U9786 (N_9786,N_5417,N_6794);
nor U9787 (N_9787,N_6639,N_7285);
nand U9788 (N_9788,N_5156,N_7171);
or U9789 (N_9789,N_6210,N_6215);
and U9790 (N_9790,N_6356,N_7453);
nand U9791 (N_9791,N_7371,N_6399);
nand U9792 (N_9792,N_7011,N_5114);
xnor U9793 (N_9793,N_6576,N_7171);
nand U9794 (N_9794,N_6070,N_5548);
nor U9795 (N_9795,N_6287,N_6649);
and U9796 (N_9796,N_6825,N_6529);
nor U9797 (N_9797,N_7144,N_6674);
and U9798 (N_9798,N_7159,N_7143);
nor U9799 (N_9799,N_5540,N_5725);
nand U9800 (N_9800,N_7229,N_5852);
nor U9801 (N_9801,N_7453,N_5380);
and U9802 (N_9802,N_7218,N_6898);
nor U9803 (N_9803,N_6250,N_6644);
nand U9804 (N_9804,N_6849,N_6147);
nand U9805 (N_9805,N_7332,N_6183);
nor U9806 (N_9806,N_6551,N_5421);
or U9807 (N_9807,N_5286,N_5306);
or U9808 (N_9808,N_5404,N_6237);
or U9809 (N_9809,N_5066,N_5561);
or U9810 (N_9810,N_7443,N_6998);
nand U9811 (N_9811,N_6285,N_7380);
nand U9812 (N_9812,N_7190,N_7375);
nand U9813 (N_9813,N_7374,N_5401);
or U9814 (N_9814,N_6844,N_7118);
or U9815 (N_9815,N_5720,N_6799);
or U9816 (N_9816,N_5000,N_5498);
or U9817 (N_9817,N_5730,N_5503);
or U9818 (N_9818,N_5417,N_6210);
and U9819 (N_9819,N_6557,N_6064);
and U9820 (N_9820,N_6163,N_7191);
and U9821 (N_9821,N_6443,N_7137);
or U9822 (N_9822,N_6587,N_7001);
nor U9823 (N_9823,N_5589,N_5087);
nor U9824 (N_9824,N_6791,N_6280);
or U9825 (N_9825,N_6216,N_6588);
nor U9826 (N_9826,N_6584,N_7180);
and U9827 (N_9827,N_5785,N_6558);
nand U9828 (N_9828,N_5478,N_6839);
and U9829 (N_9829,N_6261,N_7090);
or U9830 (N_9830,N_6167,N_5635);
or U9831 (N_9831,N_7464,N_5073);
or U9832 (N_9832,N_7172,N_5420);
or U9833 (N_9833,N_6944,N_7339);
or U9834 (N_9834,N_5560,N_7233);
nand U9835 (N_9835,N_7273,N_5623);
and U9836 (N_9836,N_7445,N_6106);
or U9837 (N_9837,N_6804,N_6163);
nand U9838 (N_9838,N_6587,N_5755);
nand U9839 (N_9839,N_5903,N_5589);
xor U9840 (N_9840,N_5240,N_5587);
and U9841 (N_9841,N_5170,N_6287);
or U9842 (N_9842,N_6767,N_5140);
nand U9843 (N_9843,N_7339,N_6181);
xnor U9844 (N_9844,N_7235,N_6406);
and U9845 (N_9845,N_6277,N_5687);
and U9846 (N_9846,N_5471,N_5525);
and U9847 (N_9847,N_6766,N_7035);
xnor U9848 (N_9848,N_6937,N_6416);
and U9849 (N_9849,N_5906,N_7332);
or U9850 (N_9850,N_7403,N_5349);
nor U9851 (N_9851,N_5296,N_6198);
and U9852 (N_9852,N_5540,N_7229);
or U9853 (N_9853,N_7333,N_6165);
and U9854 (N_9854,N_5700,N_6482);
nand U9855 (N_9855,N_6736,N_5442);
nand U9856 (N_9856,N_7236,N_7234);
and U9857 (N_9857,N_6305,N_5944);
and U9858 (N_9858,N_6172,N_5224);
and U9859 (N_9859,N_7063,N_6748);
or U9860 (N_9860,N_7390,N_7327);
and U9861 (N_9861,N_7091,N_6288);
or U9862 (N_9862,N_6549,N_6997);
nand U9863 (N_9863,N_5779,N_6676);
and U9864 (N_9864,N_5210,N_6838);
nor U9865 (N_9865,N_5656,N_5133);
or U9866 (N_9866,N_7299,N_7021);
nor U9867 (N_9867,N_7052,N_6713);
nor U9868 (N_9868,N_5455,N_6574);
or U9869 (N_9869,N_5240,N_6843);
nand U9870 (N_9870,N_6563,N_6771);
nand U9871 (N_9871,N_5507,N_6575);
and U9872 (N_9872,N_6634,N_7377);
nand U9873 (N_9873,N_6157,N_6065);
and U9874 (N_9874,N_6543,N_6451);
or U9875 (N_9875,N_5764,N_7113);
nand U9876 (N_9876,N_5578,N_7373);
nor U9877 (N_9877,N_6771,N_6062);
nand U9878 (N_9878,N_5072,N_6992);
or U9879 (N_9879,N_6358,N_5071);
or U9880 (N_9880,N_7148,N_5716);
nand U9881 (N_9881,N_6294,N_7017);
nand U9882 (N_9882,N_6236,N_7405);
nor U9883 (N_9883,N_5541,N_6546);
nand U9884 (N_9884,N_7080,N_5095);
and U9885 (N_9885,N_6347,N_5966);
nand U9886 (N_9886,N_6371,N_6846);
or U9887 (N_9887,N_6535,N_6711);
nor U9888 (N_9888,N_7009,N_5124);
nor U9889 (N_9889,N_5399,N_5682);
nand U9890 (N_9890,N_5541,N_5468);
or U9891 (N_9891,N_6845,N_5651);
nand U9892 (N_9892,N_7364,N_6911);
and U9893 (N_9893,N_5934,N_6458);
nor U9894 (N_9894,N_5104,N_5213);
nor U9895 (N_9895,N_6073,N_5656);
and U9896 (N_9896,N_6268,N_5605);
or U9897 (N_9897,N_6241,N_6815);
nand U9898 (N_9898,N_6858,N_6915);
and U9899 (N_9899,N_7389,N_5244);
nor U9900 (N_9900,N_6441,N_7439);
and U9901 (N_9901,N_7158,N_6161);
or U9902 (N_9902,N_7148,N_6318);
and U9903 (N_9903,N_7345,N_7231);
nor U9904 (N_9904,N_6022,N_5643);
and U9905 (N_9905,N_5711,N_6940);
nand U9906 (N_9906,N_5672,N_7157);
and U9907 (N_9907,N_7463,N_5655);
and U9908 (N_9908,N_7144,N_5491);
nand U9909 (N_9909,N_5791,N_7453);
nand U9910 (N_9910,N_6850,N_5028);
nand U9911 (N_9911,N_5826,N_5516);
and U9912 (N_9912,N_6131,N_5864);
nand U9913 (N_9913,N_5235,N_6139);
and U9914 (N_9914,N_7344,N_6820);
or U9915 (N_9915,N_6216,N_6145);
or U9916 (N_9916,N_5470,N_5550);
nor U9917 (N_9917,N_5017,N_6294);
or U9918 (N_9918,N_7035,N_5651);
and U9919 (N_9919,N_6879,N_6255);
nand U9920 (N_9920,N_6698,N_6460);
nand U9921 (N_9921,N_6922,N_5324);
nand U9922 (N_9922,N_6247,N_7310);
and U9923 (N_9923,N_7457,N_6252);
nor U9924 (N_9924,N_5162,N_6233);
nand U9925 (N_9925,N_7197,N_7018);
nor U9926 (N_9926,N_5006,N_6788);
nand U9927 (N_9927,N_6083,N_7369);
nand U9928 (N_9928,N_5648,N_5910);
nor U9929 (N_9929,N_6885,N_5772);
and U9930 (N_9930,N_6135,N_5535);
and U9931 (N_9931,N_6872,N_5705);
nor U9932 (N_9932,N_5232,N_6072);
and U9933 (N_9933,N_5286,N_5460);
or U9934 (N_9934,N_6118,N_7030);
and U9935 (N_9935,N_5638,N_6313);
nand U9936 (N_9936,N_5321,N_7085);
and U9937 (N_9937,N_6634,N_6194);
nand U9938 (N_9938,N_5681,N_5725);
and U9939 (N_9939,N_5317,N_6395);
and U9940 (N_9940,N_7068,N_5797);
or U9941 (N_9941,N_5980,N_6054);
and U9942 (N_9942,N_6914,N_6007);
or U9943 (N_9943,N_6784,N_5286);
or U9944 (N_9944,N_6996,N_5438);
or U9945 (N_9945,N_7175,N_6772);
and U9946 (N_9946,N_6728,N_7347);
and U9947 (N_9947,N_5459,N_6851);
nor U9948 (N_9948,N_5817,N_6408);
nand U9949 (N_9949,N_5037,N_6523);
or U9950 (N_9950,N_6503,N_6111);
nand U9951 (N_9951,N_6250,N_5350);
xnor U9952 (N_9952,N_6810,N_6041);
or U9953 (N_9953,N_6762,N_6065);
nand U9954 (N_9954,N_6507,N_5809);
nor U9955 (N_9955,N_6574,N_7363);
and U9956 (N_9956,N_6195,N_6238);
nor U9957 (N_9957,N_6069,N_6349);
nand U9958 (N_9958,N_7374,N_5631);
or U9959 (N_9959,N_7008,N_5047);
and U9960 (N_9960,N_5273,N_5149);
nor U9961 (N_9961,N_5514,N_5895);
or U9962 (N_9962,N_5876,N_7037);
and U9963 (N_9963,N_5847,N_5081);
and U9964 (N_9964,N_7357,N_5439);
nand U9965 (N_9965,N_6359,N_7377);
xor U9966 (N_9966,N_6896,N_5562);
nand U9967 (N_9967,N_5846,N_6955);
or U9968 (N_9968,N_6079,N_6777);
and U9969 (N_9969,N_5080,N_6976);
or U9970 (N_9970,N_5378,N_5216);
nor U9971 (N_9971,N_6363,N_6981);
nand U9972 (N_9972,N_5852,N_5383);
nand U9973 (N_9973,N_6345,N_7100);
nor U9974 (N_9974,N_5832,N_6736);
nand U9975 (N_9975,N_7159,N_6845);
nor U9976 (N_9976,N_5344,N_7122);
and U9977 (N_9977,N_6864,N_5695);
nand U9978 (N_9978,N_7263,N_6944);
nor U9979 (N_9979,N_6376,N_6558);
nand U9980 (N_9980,N_5381,N_6067);
or U9981 (N_9981,N_5027,N_5033);
nor U9982 (N_9982,N_7162,N_6703);
nor U9983 (N_9983,N_6324,N_6773);
or U9984 (N_9984,N_6974,N_5544);
nand U9985 (N_9985,N_5176,N_7153);
nor U9986 (N_9986,N_7257,N_5905);
nand U9987 (N_9987,N_5424,N_6981);
nand U9988 (N_9988,N_6025,N_6856);
or U9989 (N_9989,N_5015,N_5953);
nor U9990 (N_9990,N_6287,N_6643);
or U9991 (N_9991,N_7464,N_5617);
nand U9992 (N_9992,N_5722,N_7488);
nor U9993 (N_9993,N_6833,N_6067);
or U9994 (N_9994,N_6875,N_7468);
or U9995 (N_9995,N_5150,N_6991);
and U9996 (N_9996,N_5805,N_5635);
nor U9997 (N_9997,N_7065,N_6254);
and U9998 (N_9998,N_6200,N_5917);
xnor U9999 (N_9999,N_6254,N_5416);
or UO_0 (O_0,N_8217,N_8359);
nand UO_1 (O_1,N_9666,N_7553);
nor UO_2 (O_2,N_8633,N_9259);
xnor UO_3 (O_3,N_8938,N_8513);
nand UO_4 (O_4,N_7888,N_7829);
nor UO_5 (O_5,N_9693,N_9633);
nand UO_6 (O_6,N_8128,N_7599);
and UO_7 (O_7,N_9062,N_9940);
nand UO_8 (O_8,N_7697,N_8953);
nand UO_9 (O_9,N_7979,N_9898);
nand UO_10 (O_10,N_7756,N_8675);
or UO_11 (O_11,N_7900,N_9987);
nor UO_12 (O_12,N_9829,N_9254);
nor UO_13 (O_13,N_7731,N_7866);
and UO_14 (O_14,N_8635,N_9539);
or UO_15 (O_15,N_9239,N_7556);
and UO_16 (O_16,N_8986,N_8244);
nor UO_17 (O_17,N_9065,N_7919);
nor UO_18 (O_18,N_7615,N_9314);
or UO_19 (O_19,N_8255,N_8700);
or UO_20 (O_20,N_9715,N_8252);
or UO_21 (O_21,N_9051,N_9282);
nand UO_22 (O_22,N_7739,N_8145);
nand UO_23 (O_23,N_8914,N_8548);
nand UO_24 (O_24,N_9344,N_9193);
or UO_25 (O_25,N_7635,N_9774);
or UO_26 (O_26,N_7534,N_7962);
nand UO_27 (O_27,N_8107,N_8231);
and UO_28 (O_28,N_8417,N_8027);
nand UO_29 (O_29,N_9077,N_8623);
nand UO_30 (O_30,N_8447,N_9567);
nor UO_31 (O_31,N_8903,N_8339);
or UO_32 (O_32,N_8710,N_7800);
xnor UO_33 (O_33,N_9104,N_8684);
and UO_34 (O_34,N_8076,N_8759);
nor UO_35 (O_35,N_9985,N_8337);
nand UO_36 (O_36,N_8280,N_9771);
or UO_37 (O_37,N_8628,N_7719);
xnor UO_38 (O_38,N_8752,N_9155);
and UO_39 (O_39,N_9569,N_8381);
and UO_40 (O_40,N_7580,N_8419);
and UO_41 (O_41,N_7746,N_7708);
and UO_42 (O_42,N_9989,N_8834);
nand UO_43 (O_43,N_7652,N_9637);
nand UO_44 (O_44,N_9682,N_9749);
nand UO_45 (O_45,N_9769,N_9802);
nand UO_46 (O_46,N_8606,N_9589);
nor UO_47 (O_47,N_9203,N_9098);
nor UO_48 (O_48,N_9632,N_8783);
or UO_49 (O_49,N_9468,N_8390);
nor UO_50 (O_50,N_7810,N_7895);
nand UO_51 (O_51,N_8894,N_9755);
or UO_52 (O_52,N_8556,N_9507);
and UO_53 (O_53,N_8453,N_7533);
and UO_54 (O_54,N_7871,N_9484);
and UO_55 (O_55,N_8492,N_9641);
and UO_56 (O_56,N_9429,N_9742);
and UO_57 (O_57,N_8038,N_7943);
nand UO_58 (O_58,N_7679,N_9007);
or UO_59 (O_59,N_8004,N_9928);
and UO_60 (O_60,N_9028,N_9426);
nor UO_61 (O_61,N_9945,N_8477);
xor UO_62 (O_62,N_7591,N_8388);
and UO_63 (O_63,N_9325,N_8857);
nor UO_64 (O_64,N_8179,N_8006);
and UO_65 (O_65,N_9927,N_9806);
nand UO_66 (O_66,N_8432,N_7993);
nor UO_67 (O_67,N_9501,N_8241);
nand UO_68 (O_68,N_9827,N_9859);
nor UO_69 (O_69,N_8075,N_9370);
nand UO_70 (O_70,N_8977,N_7820);
nand UO_71 (O_71,N_8097,N_8227);
nand UO_72 (O_72,N_8139,N_9346);
nor UO_73 (O_73,N_8655,N_7791);
nand UO_74 (O_74,N_9323,N_7862);
nor UO_75 (O_75,N_8459,N_7514);
and UO_76 (O_76,N_8020,N_8908);
or UO_77 (O_77,N_8910,N_9964);
or UO_78 (O_78,N_7890,N_8992);
nand UO_79 (O_79,N_8304,N_8287);
nand UO_80 (O_80,N_8742,N_8362);
nor UO_81 (O_81,N_9422,N_9247);
nand UO_82 (O_82,N_9610,N_8412);
nor UO_83 (O_83,N_8592,N_8303);
and UO_84 (O_84,N_7620,N_8220);
nor UO_85 (O_85,N_8768,N_7834);
or UO_86 (O_86,N_8468,N_9969);
or UO_87 (O_87,N_7964,N_8413);
or UO_88 (O_88,N_8746,N_8425);
nand UO_89 (O_89,N_9371,N_8129);
nor UO_90 (O_90,N_8519,N_7554);
nand UO_91 (O_91,N_8100,N_8801);
or UO_92 (O_92,N_9582,N_9981);
or UO_93 (O_93,N_9948,N_9008);
and UO_94 (O_94,N_9034,N_8581);
nand UO_95 (O_95,N_9384,N_8266);
or UO_96 (O_96,N_8888,N_8836);
xor UO_97 (O_97,N_7913,N_9931);
or UO_98 (O_98,N_7994,N_7680);
nand UO_99 (O_99,N_9949,N_9509);
nand UO_100 (O_100,N_8000,N_9258);
nand UO_101 (O_101,N_8593,N_8315);
and UO_102 (O_102,N_9256,N_9116);
or UO_103 (O_103,N_8011,N_9498);
or UO_104 (O_104,N_9112,N_9505);
and UO_105 (O_105,N_8921,N_8336);
nor UO_106 (O_106,N_8144,N_9456);
and UO_107 (O_107,N_8818,N_8162);
nand UO_108 (O_108,N_9230,N_8773);
nor UO_109 (O_109,N_8407,N_9257);
nand UO_110 (O_110,N_9364,N_9932);
nand UO_111 (O_111,N_9482,N_8278);
nor UO_112 (O_112,N_9452,N_7968);
or UO_113 (O_113,N_8999,N_9957);
or UO_114 (O_114,N_7836,N_8104);
nor UO_115 (O_115,N_9551,N_9673);
nand UO_116 (O_116,N_9503,N_7629);
nor UO_117 (O_117,N_8269,N_8907);
nor UO_118 (O_118,N_9188,N_8532);
nor UO_119 (O_119,N_8579,N_8415);
nor UO_120 (O_120,N_8307,N_9655);
and UO_121 (O_121,N_8658,N_8463);
or UO_122 (O_122,N_9372,N_9500);
and UO_123 (O_123,N_8512,N_7725);
and UO_124 (O_124,N_8137,N_8837);
or UO_125 (O_125,N_8561,N_9022);
nand UO_126 (O_126,N_8958,N_8219);
nor UO_127 (O_127,N_8835,N_8276);
nand UO_128 (O_128,N_9643,N_8717);
or UO_129 (O_129,N_9407,N_8366);
or UO_130 (O_130,N_8673,N_9118);
and UO_131 (O_131,N_8612,N_9374);
and UO_132 (O_132,N_7601,N_8571);
and UO_133 (O_133,N_8611,N_8887);
or UO_134 (O_134,N_9237,N_9553);
nand UO_135 (O_135,N_9638,N_9302);
nor UO_136 (O_136,N_7813,N_7526);
nand UO_137 (O_137,N_8474,N_7980);
nand UO_138 (O_138,N_7602,N_7718);
nand UO_139 (O_139,N_7654,N_7677);
or UO_140 (O_140,N_8472,N_8896);
and UO_141 (O_141,N_9812,N_8165);
and UO_142 (O_142,N_7869,N_9664);
nand UO_143 (O_143,N_8186,N_7872);
or UO_144 (O_144,N_7575,N_8657);
or UO_145 (O_145,N_9273,N_8018);
nor UO_146 (O_146,N_8654,N_8972);
and UO_147 (O_147,N_8901,N_8461);
or UO_148 (O_148,N_8349,N_9462);
nand UO_149 (O_149,N_9318,N_8214);
or UO_150 (O_150,N_9778,N_7887);
and UO_151 (O_151,N_8721,N_8886);
nand UO_152 (O_152,N_8465,N_8796);
nor UO_153 (O_153,N_8210,N_7548);
xor UO_154 (O_154,N_9326,N_9397);
or UO_155 (O_155,N_8501,N_8072);
or UO_156 (O_156,N_9005,N_9861);
xor UO_157 (O_157,N_9905,N_9951);
or UO_158 (O_158,N_9076,N_9182);
and UO_159 (O_159,N_8713,N_8950);
or UO_160 (O_160,N_8155,N_7894);
or UO_161 (O_161,N_9692,N_9950);
nand UO_162 (O_162,N_9408,N_9274);
nand UO_163 (O_163,N_9466,N_7550);
nor UO_164 (O_164,N_7990,N_9049);
or UO_165 (O_165,N_7734,N_7710);
or UO_166 (O_166,N_9853,N_7774);
nand UO_167 (O_167,N_9331,N_9296);
nand UO_168 (O_168,N_8288,N_8061);
nand UO_169 (O_169,N_8136,N_8848);
nand UO_170 (O_170,N_9440,N_7683);
and UO_171 (O_171,N_9026,N_9517);
and UO_172 (O_172,N_8709,N_9856);
nand UO_173 (O_173,N_9317,N_8181);
and UO_174 (O_174,N_8060,N_9622);
nand UO_175 (O_175,N_9211,N_8927);
nor UO_176 (O_176,N_9731,N_8828);
and UO_177 (O_177,N_9917,N_8201);
and UO_178 (O_178,N_7597,N_8542);
nor UO_179 (O_179,N_8427,N_7507);
or UO_180 (O_180,N_7547,N_7752);
nand UO_181 (O_181,N_9578,N_9094);
or UO_182 (O_182,N_9297,N_7864);
nand UO_183 (O_183,N_8987,N_8749);
nor UO_184 (O_184,N_9107,N_7584);
or UO_185 (O_185,N_8706,N_9227);
nor UO_186 (O_186,N_9588,N_9037);
and UO_187 (O_187,N_8878,N_7847);
or UO_188 (O_188,N_9139,N_8125);
nor UO_189 (O_189,N_8180,N_7692);
or UO_190 (O_190,N_8829,N_8433);
nor UO_191 (O_191,N_8567,N_7702);
nor UO_192 (O_192,N_8974,N_8583);
and UO_193 (O_193,N_7779,N_7832);
and UO_194 (O_194,N_8726,N_7647);
and UO_195 (O_195,N_8577,N_8728);
and UO_196 (O_196,N_9903,N_9916);
and UO_197 (O_197,N_9820,N_8044);
nand UO_198 (O_198,N_8729,N_7787);
or UO_199 (O_199,N_8504,N_9128);
and UO_200 (O_200,N_7541,N_8598);
nor UO_201 (O_201,N_7579,N_7600);
nand UO_202 (O_202,N_9518,N_9670);
or UO_203 (O_203,N_8329,N_8452);
or UO_204 (O_204,N_8310,N_8355);
or UO_205 (O_205,N_9956,N_9497);
nand UO_206 (O_206,N_7642,N_9123);
and UO_207 (O_207,N_7730,N_7870);
nor UO_208 (O_208,N_9773,N_9625);
nand UO_209 (O_209,N_8521,N_8631);
nor UO_210 (O_210,N_7559,N_8079);
and UO_211 (O_211,N_7846,N_9563);
nor UO_212 (O_212,N_8377,N_8617);
nand UO_213 (O_213,N_8274,N_9597);
or UO_214 (O_214,N_8694,N_7638);
or UO_215 (O_215,N_8962,N_7755);
nand UO_216 (O_216,N_9840,N_9058);
nor UO_217 (O_217,N_9975,N_9477);
and UO_218 (O_218,N_9063,N_7923);
or UO_219 (O_219,N_8699,N_9513);
or UO_220 (O_220,N_9779,N_9402);
nand UO_221 (O_221,N_9250,N_8790);
or UO_222 (O_222,N_7537,N_8402);
or UO_223 (O_223,N_9910,N_9399);
nor UO_224 (O_224,N_8607,N_8926);
or UO_225 (O_225,N_8531,N_8480);
nand UO_226 (O_226,N_8849,N_9711);
and UO_227 (O_227,N_8229,N_7812);
and UO_228 (O_228,N_8423,N_9321);
nor UO_229 (O_229,N_9675,N_8394);
and UO_230 (O_230,N_9411,N_8960);
and UO_231 (O_231,N_8846,N_9191);
nor UO_232 (O_232,N_9499,N_9612);
nand UO_233 (O_233,N_9281,N_9209);
or UO_234 (O_234,N_8822,N_8923);
nand UO_235 (O_235,N_8948,N_8015);
nand UO_236 (O_236,N_8338,N_7724);
nand UO_237 (O_237,N_7793,N_7997);
nor UO_238 (O_238,N_8246,N_8161);
or UO_239 (O_239,N_7539,N_7711);
and UO_240 (O_240,N_9704,N_9733);
and UO_241 (O_241,N_7751,N_8140);
nor UO_242 (O_242,N_8070,N_8807);
or UO_243 (O_243,N_8956,N_8373);
and UO_244 (O_244,N_9119,N_8518);
nor UO_245 (O_245,N_8971,N_8185);
and UO_246 (O_246,N_8770,N_8985);
and UO_247 (O_247,N_9432,N_9142);
nor UO_248 (O_248,N_7795,N_8391);
or UO_249 (O_249,N_8672,N_7714);
nand UO_250 (O_250,N_8664,N_9968);
and UO_251 (O_251,N_8268,N_8558);
nand UO_252 (O_252,N_7880,N_8372);
and UO_253 (O_253,N_9178,N_8871);
and UO_254 (O_254,N_7703,N_8467);
nand UO_255 (O_255,N_8363,N_7960);
nand UO_256 (O_256,N_7560,N_8582);
and UO_257 (O_257,N_9900,N_9447);
nand UO_258 (O_258,N_8641,N_7833);
and UO_259 (O_259,N_7852,N_7838);
nand UO_260 (O_260,N_7903,N_9690);
and UO_261 (O_261,N_9961,N_7590);
or UO_262 (O_262,N_9716,N_8046);
and UO_263 (O_263,N_9029,N_8755);
nand UO_264 (O_264,N_9546,N_8460);
nand UO_265 (O_265,N_8141,N_9923);
or UO_266 (O_266,N_9572,N_8080);
nand UO_267 (O_267,N_9925,N_9515);
nor UO_268 (O_268,N_9556,N_9168);
nor UO_269 (O_269,N_7940,N_9018);
or UO_270 (O_270,N_7513,N_9242);
nor UO_271 (O_271,N_7650,N_7571);
xnor UO_272 (O_272,N_8990,N_9414);
nor UO_273 (O_273,N_9004,N_9100);
nand UO_274 (O_274,N_8434,N_9952);
and UO_275 (O_275,N_7543,N_8959);
or UO_276 (O_276,N_8570,N_8902);
and UO_277 (O_277,N_8481,N_8799);
nand UO_278 (O_278,N_8979,N_7529);
nand UO_279 (O_279,N_9712,N_9640);
nor UO_280 (O_280,N_9381,N_8895);
or UO_281 (O_281,N_8753,N_9490);
and UO_282 (O_282,N_7592,N_7564);
and UO_283 (O_283,N_8462,N_8994);
and UO_284 (O_284,N_9453,N_7848);
nor UO_285 (O_285,N_9213,N_8313);
or UO_286 (O_286,N_7959,N_7639);
and UO_287 (O_287,N_8067,N_9683);
nand UO_288 (O_288,N_7565,N_9228);
nand UO_289 (O_289,N_8360,N_8970);
nor UO_290 (O_290,N_7896,N_9271);
or UO_291 (O_291,N_8915,N_8774);
and UO_292 (O_292,N_7897,N_8007);
or UO_293 (O_293,N_9521,N_9786);
or UO_294 (O_294,N_9628,N_9721);
nand UO_295 (O_295,N_9174,N_8010);
nand UO_296 (O_296,N_8376,N_9998);
nor UO_297 (O_297,N_7874,N_8560);
nand UO_298 (O_298,N_9959,N_8573);
nand UO_299 (O_299,N_7763,N_8230);
and UO_300 (O_300,N_7566,N_9870);
nor UO_301 (O_301,N_9125,N_7891);
xnor UO_302 (O_302,N_8855,N_8319);
nand UO_303 (O_303,N_7552,N_7986);
and UO_304 (O_304,N_8098,N_7821);
nor UO_305 (O_305,N_9357,N_9745);
or UO_306 (O_306,N_9815,N_8057);
nand UO_307 (O_307,N_8647,N_8646);
or UO_308 (O_308,N_9290,N_8904);
nand UO_309 (O_309,N_9377,N_7624);
and UO_310 (O_310,N_8215,N_9485);
nand UO_311 (O_311,N_8300,N_8416);
nor UO_312 (O_312,N_8357,N_9417);
or UO_313 (O_313,N_8042,N_9003);
xor UO_314 (O_314,N_7694,N_9489);
and UO_315 (O_315,N_8844,N_7925);
nand UO_316 (O_316,N_8158,N_8808);
nor UO_317 (O_317,N_7910,N_9087);
and UO_318 (O_318,N_7957,N_7531);
nor UO_319 (O_319,N_8105,N_9519);
nor UO_320 (O_320,N_7740,N_8688);
or UO_321 (O_321,N_9061,N_7562);
or UO_322 (O_322,N_7551,N_7569);
xnor UO_323 (O_323,N_7728,N_9801);
and UO_324 (O_324,N_9554,N_9423);
nand UO_325 (O_325,N_7645,N_8758);
nor UO_326 (O_326,N_9792,N_9857);
nor UO_327 (O_327,N_7656,N_8810);
or UO_328 (O_328,N_7792,N_9093);
or UO_329 (O_329,N_9043,N_8618);
nand UO_330 (O_330,N_9092,N_9210);
or UO_331 (O_331,N_9449,N_9298);
nor UO_332 (O_332,N_8594,N_7856);
or UO_333 (O_333,N_9580,N_8036);
nand UO_334 (O_334,N_9761,N_8195);
nor UO_335 (O_335,N_8533,N_8663);
nor UO_336 (O_336,N_8508,N_9783);
nor UO_337 (O_337,N_9019,N_9869);
nor UO_338 (O_338,N_9953,N_7517);
and UO_339 (O_339,N_8980,N_8937);
nor UO_340 (O_340,N_8609,N_8171);
nor UO_341 (O_341,N_8265,N_9467);
nor UO_342 (O_342,N_8760,N_8997);
and UO_343 (O_343,N_7875,N_9156);
nor UO_344 (O_344,N_8649,N_7744);
nor UO_345 (O_345,N_7664,N_8850);
nor UO_346 (O_346,N_8114,N_9260);
or UO_347 (O_347,N_8820,N_9152);
or UO_348 (O_348,N_9780,N_8949);
nand UO_349 (O_349,N_9868,N_7912);
nor UO_350 (O_350,N_8873,N_8714);
nand UO_351 (O_351,N_8976,N_8989);
or UO_352 (O_352,N_8955,N_9451);
or UO_353 (O_353,N_7860,N_9849);
nand UO_354 (O_354,N_8147,N_7884);
or UO_355 (O_355,N_7809,N_9681);
and UO_356 (O_356,N_8775,N_9656);
nor UO_357 (O_357,N_9966,N_9891);
and UO_358 (O_358,N_8111,N_8443);
and UO_359 (O_359,N_7618,N_9676);
nand UO_360 (O_360,N_9995,N_7988);
or UO_361 (O_361,N_9036,N_7532);
or UO_362 (O_362,N_9338,N_9618);
nand UO_363 (O_363,N_8900,N_9838);
nor UO_364 (O_364,N_8741,N_8778);
and UO_365 (O_365,N_9754,N_8854);
and UO_366 (O_366,N_7955,N_8207);
nand UO_367 (O_367,N_8662,N_9251);
or UO_368 (O_368,N_9115,N_9504);
and UO_369 (O_369,N_8745,N_8256);
nor UO_370 (O_370,N_9329,N_8912);
and UO_371 (O_371,N_9844,N_8942);
or UO_372 (O_372,N_8931,N_8471);
nand UO_373 (O_373,N_7608,N_8639);
and UO_374 (O_374,N_9709,N_9933);
and UO_375 (O_375,N_7742,N_9201);
or UO_376 (O_376,N_8473,N_9926);
or UO_377 (O_377,N_9304,N_9516);
or UO_378 (O_378,N_9958,N_8321);
nand UO_379 (O_379,N_8340,N_8167);
nand UO_380 (O_380,N_8037,N_9579);
nand UO_381 (O_381,N_8716,N_8557);
nand UO_382 (O_382,N_7911,N_9831);
or UO_383 (O_383,N_8211,N_7717);
and UO_384 (O_384,N_7991,N_9538);
nor UO_385 (O_385,N_8242,N_8392);
nand UO_386 (O_386,N_8206,N_9124);
nand UO_387 (O_387,N_9858,N_8762);
or UO_388 (O_388,N_8676,N_7825);
or UO_389 (O_389,N_9739,N_9396);
nand UO_390 (O_390,N_9566,N_8049);
nand UO_391 (O_391,N_8156,N_8187);
and UO_392 (O_392,N_9481,N_7572);
nand UO_393 (O_393,N_7503,N_9383);
nor UO_394 (O_394,N_9176,N_9053);
or UO_395 (O_395,N_7595,N_7768);
and UO_396 (O_396,N_7935,N_9261);
and UO_397 (O_397,N_9642,N_7563);
nor UO_398 (O_398,N_9270,N_7839);
and UO_399 (O_399,N_7506,N_9993);
nor UO_400 (O_400,N_8597,N_9021);
or UO_401 (O_401,N_9608,N_7920);
or UO_402 (O_402,N_8817,N_9624);
or UO_403 (O_403,N_9760,N_9984);
nor UO_404 (O_404,N_8034,N_8839);
nand UO_405 (O_405,N_8348,N_7762);
or UO_406 (O_406,N_8780,N_9573);
nand UO_407 (O_407,N_7523,N_8146);
or UO_408 (O_408,N_8543,N_8929);
or UO_409 (O_409,N_7589,N_8464);
nand UO_410 (O_410,N_9224,N_8798);
or UO_411 (O_411,N_8869,N_9272);
or UO_412 (O_412,N_7950,N_8189);
nor UO_413 (O_413,N_8764,N_9919);
and UO_414 (O_414,N_9292,N_9924);
nand UO_415 (O_415,N_8382,N_9699);
nand UO_416 (O_416,N_9050,N_9535);
nand UO_417 (O_417,N_9091,N_9723);
nor UO_418 (O_418,N_8719,N_8361);
nor UO_419 (O_419,N_9421,N_8346);
nand UO_420 (O_420,N_8751,N_8627);
nor UO_421 (O_421,N_8205,N_9635);
and UO_422 (O_422,N_8550,N_7732);
and UO_423 (O_423,N_9389,N_7705);
or UO_424 (O_424,N_9889,N_8791);
nand UO_425 (O_425,N_7630,N_7678);
or UO_426 (O_426,N_9141,N_8715);
and UO_427 (O_427,N_7616,N_9850);
nor UO_428 (O_428,N_7876,N_8698);
and UO_429 (O_429,N_9601,N_8736);
and UO_430 (O_430,N_7873,N_7588);
and UO_431 (O_431,N_8420,N_8648);
and UO_432 (O_432,N_9241,N_8693);
nor UO_433 (O_433,N_9287,N_8541);
nor UO_434 (O_434,N_8743,N_9121);
nand UO_435 (O_435,N_9753,N_8174);
and UO_436 (O_436,N_9027,N_9198);
and UO_437 (O_437,N_8112,N_9543);
and UO_438 (O_438,N_9986,N_7606);
xor UO_439 (O_439,N_8450,N_9054);
and UO_440 (O_440,N_7818,N_9825);
and UO_441 (O_441,N_9069,N_8784);
nand UO_442 (O_442,N_8251,N_8578);
nand UO_443 (O_443,N_8602,N_9348);
or UO_444 (O_444,N_8811,N_8476);
nand UO_445 (O_445,N_8496,N_9181);
nor UO_446 (O_446,N_7609,N_8405);
and UO_447 (O_447,N_8151,N_7961);
or UO_448 (O_448,N_8920,N_9097);
nor UO_449 (O_449,N_7555,N_9415);
or UO_450 (O_450,N_9854,N_7691);
or UO_451 (O_451,N_7977,N_7504);
nor UO_452 (O_452,N_7817,N_9584);
or UO_453 (O_453,N_8073,N_9725);
nor UO_454 (O_454,N_9390,N_9083);
and UO_455 (O_455,N_7685,N_8951);
xnor UO_456 (O_456,N_7996,N_9147);
nor UO_457 (O_457,N_8198,N_9057);
nand UO_458 (O_458,N_8192,N_9388);
or UO_459 (O_459,N_8991,N_9688);
nor UO_460 (O_460,N_8967,N_9767);
nor UO_461 (O_461,N_9560,N_7796);
nor UO_462 (O_462,N_9459,N_8881);
or UO_463 (O_463,N_9609,N_9430);
and UO_464 (O_464,N_8317,N_9263);
and UO_465 (O_465,N_9627,N_9602);
and UO_466 (O_466,N_8776,N_7826);
nand UO_467 (O_467,N_9883,N_9108);
or UO_468 (O_468,N_9526,N_8383);
nand UO_469 (O_469,N_7966,N_9531);
and UO_470 (O_470,N_9621,N_8169);
and UO_471 (O_471,N_9285,N_9896);
and UO_472 (O_472,N_9997,N_9342);
nand UO_473 (O_473,N_8142,N_8932);
nor UO_474 (O_474,N_7790,N_8071);
nor UO_475 (O_475,N_9033,N_9345);
nand UO_476 (O_476,N_8122,N_9450);
and UO_477 (O_477,N_7727,N_9536);
and UO_478 (O_478,N_9818,N_9701);
or UO_479 (O_479,N_9179,N_9730);
and UO_480 (O_480,N_9525,N_7978);
nand UO_481 (O_481,N_9394,N_7771);
or UO_482 (O_482,N_8569,N_9594);
or UO_483 (O_483,N_8106,N_7593);
nand UO_484 (O_484,N_7759,N_8968);
nor UO_485 (O_485,N_8580,N_7781);
and UO_486 (O_486,N_8860,N_8421);
nand UO_487 (O_487,N_9544,N_9267);
and UO_488 (O_488,N_9040,N_7646);
nand UO_489 (O_489,N_8704,N_8286);
nand UO_490 (O_490,N_7803,N_7509);
or UO_491 (O_491,N_8279,N_8086);
and UO_492 (O_492,N_9136,N_9249);
or UO_493 (O_493,N_9977,N_9127);
nor UO_494 (O_494,N_8094,N_7519);
nor UO_495 (O_495,N_9277,N_9074);
xnor UO_496 (O_496,N_9491,N_9316);
nand UO_497 (O_497,N_8535,N_9159);
nor UO_498 (O_498,N_7929,N_8002);
or UO_499 (O_499,N_9685,N_8576);
nand UO_500 (O_500,N_8812,N_7885);
or UO_501 (O_501,N_9145,N_8127);
nand UO_502 (O_502,N_8679,N_8389);
nand UO_503 (O_503,N_8085,N_7587);
and UO_504 (O_504,N_8124,N_9486);
nor UO_505 (O_505,N_9359,N_8964);
nor UO_506 (O_506,N_7956,N_7849);
nor UO_507 (O_507,N_7926,N_8514);
nand UO_508 (O_508,N_9436,N_7631);
and UO_509 (O_509,N_8975,N_9403);
and UO_510 (O_510,N_8291,N_9591);
nor UO_511 (O_511,N_9445,N_7879);
or UO_512 (O_512,N_9912,N_8893);
and UO_513 (O_513,N_7696,N_8188);
nand UO_514 (O_514,N_8874,N_7798);
or UO_515 (O_515,N_8879,N_8905);
and UO_516 (O_516,N_7510,N_8625);
nand UO_517 (O_517,N_9524,N_7586);
nor UO_518 (O_518,N_9080,N_7845);
nor UO_519 (O_519,N_8685,N_9428);
or UO_520 (O_520,N_9192,N_8170);
or UO_521 (O_521,N_9552,N_8194);
nor UO_522 (O_522,N_7814,N_9424);
nand UO_523 (O_523,N_8064,N_7861);
nand UO_524 (O_524,N_8538,N_9965);
or UO_525 (O_525,N_8936,N_9382);
nand UO_526 (O_526,N_8439,N_8534);
and UO_527 (O_527,N_9212,N_9023);
nand UO_528 (O_528,N_9532,N_9218);
nor UO_529 (O_529,N_9911,N_9439);
nor UO_530 (O_530,N_9163,N_8160);
nor UO_531 (O_531,N_7682,N_8610);
or UO_532 (O_532,N_8119,N_9474);
nor UO_533 (O_533,N_9565,N_8720);
or UO_534 (O_534,N_9743,N_8074);
nor UO_535 (O_535,N_8705,N_9041);
nand UO_536 (O_536,N_8549,N_9144);
or UO_537 (O_537,N_9153,N_8261);
nor UO_538 (O_538,N_7527,N_9970);
nor UO_539 (O_539,N_8485,N_8234);
and UO_540 (O_540,N_7699,N_7837);
nor UO_541 (O_541,N_9888,N_7819);
nand UO_542 (O_542,N_8586,N_8707);
and UO_543 (O_543,N_8826,N_8152);
nor UO_544 (O_544,N_9262,N_9583);
and UO_545 (O_545,N_7583,N_9180);
nor UO_546 (O_546,N_8494,N_9807);
nor UO_547 (O_547,N_9186,N_7688);
and UO_548 (O_548,N_8232,N_8297);
and UO_549 (O_549,N_9758,N_9702);
nor UO_550 (O_550,N_8025,N_8154);
and UO_551 (O_551,N_7877,N_8536);
or UO_552 (O_552,N_9885,N_8842);
or UO_553 (O_553,N_9920,N_9705);
nor UO_554 (O_554,N_8335,N_9365);
nor UO_555 (O_555,N_8877,N_9511);
nor UO_556 (O_556,N_9475,N_8506);
nor UO_557 (O_557,N_7637,N_9537);
nor UO_558 (O_558,N_7892,N_9939);
nor UO_559 (O_559,N_8540,N_9199);
nor UO_560 (O_560,N_9620,N_7749);
and UO_561 (O_561,N_8327,N_7806);
xnor UO_562 (O_562,N_8622,N_8944);
or UO_563 (O_563,N_9157,N_7614);
and UO_564 (O_564,N_7850,N_9851);
or UO_565 (O_565,N_9616,N_9719);
nand UO_566 (O_566,N_8634,N_7799);
nand UO_567 (O_567,N_8334,N_9379);
nand UO_568 (O_568,N_9626,N_8995);
nor UO_569 (O_569,N_8455,N_9710);
nor UO_570 (O_570,N_7713,N_8865);
nand UO_571 (O_571,N_8354,N_8123);
nand UO_572 (O_572,N_8233,N_9623);
nor UO_573 (O_573,N_9133,N_9915);
nand UO_574 (O_574,N_7761,N_8711);
nor UO_575 (O_575,N_8099,N_9955);
and UO_576 (O_576,N_8864,N_9406);
or UO_577 (O_577,N_9605,N_7636);
or UO_578 (O_578,N_9391,N_9322);
nor UO_579 (O_579,N_8816,N_9520);
or UO_580 (O_580,N_7835,N_9744);
and UO_581 (O_581,N_8756,N_9547);
nor UO_582 (O_582,N_8794,N_8781);
nor UO_583 (O_583,N_8225,N_8978);
nand UO_584 (O_584,N_9558,N_8619);
or UO_585 (O_585,N_9113,N_8028);
or UO_586 (O_586,N_9312,N_9284);
nor UO_587 (O_587,N_7748,N_9599);
nand UO_588 (O_588,N_7686,N_8983);
and UO_589 (O_589,N_8294,N_9410);
nor UO_590 (O_590,N_8285,N_9660);
nor UO_591 (O_591,N_8380,N_9533);
nand UO_592 (O_592,N_7842,N_7906);
nand UO_593 (O_593,N_8574,N_9967);
or UO_594 (O_594,N_8498,N_8148);
nor UO_595 (O_595,N_8862,N_8084);
nor UO_596 (O_596,N_8840,N_9648);
nor UO_597 (O_597,N_8176,N_9495);
nand UO_598 (O_598,N_9434,N_7938);
nand UO_599 (O_599,N_9587,N_8089);
or UO_600 (O_600,N_7784,N_7975);
or UO_601 (O_601,N_8030,N_8701);
or UO_602 (O_602,N_9070,N_9225);
nor UO_603 (O_603,N_8438,N_7893);
and UO_604 (O_604,N_9992,N_9740);
nand UO_605 (O_605,N_7934,N_9630);
nand UO_606 (O_606,N_8551,N_7681);
nand UO_607 (O_607,N_8870,N_8651);
nor UO_608 (O_608,N_9880,N_7741);
nor UO_609 (O_609,N_9165,N_9512);
and UO_610 (O_610,N_9300,N_8032);
nor UO_611 (O_611,N_7577,N_9472);
and UO_612 (O_612,N_8785,N_8424);
or UO_613 (O_613,N_8515,N_8973);
and UO_614 (O_614,N_7585,N_9483);
and UO_615 (O_615,N_9138,N_9607);
nor UO_616 (O_616,N_7743,N_8545);
nor UO_617 (O_617,N_9206,N_8275);
nor UO_618 (O_618,N_9708,N_9826);
nand UO_619 (O_619,N_8113,N_9066);
and UO_620 (O_620,N_8998,N_8302);
and UO_621 (O_621,N_8369,N_9487);
nor UO_622 (O_622,N_8562,N_8456);
and UO_623 (O_623,N_9109,N_9636);
nand UO_624 (O_624,N_8021,N_9461);
or UO_625 (O_625,N_9315,N_7675);
or UO_626 (O_626,N_9697,N_8223);
or UO_627 (O_627,N_7623,N_8718);
nor UO_628 (O_628,N_8118,N_9140);
nand UO_629 (O_629,N_8493,N_7914);
and UO_630 (O_630,N_7757,N_9020);
nor UO_631 (O_631,N_9283,N_9763);
nor UO_632 (O_632,N_7985,N_8322);
nor UO_633 (O_633,N_7573,N_7687);
nor UO_634 (O_634,N_8308,N_8016);
and UO_635 (O_635,N_9700,N_8740);
nor UO_636 (O_636,N_9764,N_9234);
nor UO_637 (O_637,N_8945,N_9131);
xnor UO_638 (O_638,N_9813,N_9465);
and UO_639 (O_639,N_8899,N_8517);
nand UO_640 (O_640,N_9568,N_9380);
nand UO_641 (O_641,N_8430,N_9289);
nor UO_642 (O_642,N_7859,N_9895);
xor UO_643 (O_643,N_9471,N_9324);
or UO_644 (O_644,N_7927,N_9823);
and UO_645 (O_645,N_7698,N_9613);
nor UO_646 (O_646,N_8963,N_9223);
and UO_647 (O_647,N_9677,N_8565);
nand UO_648 (O_648,N_9862,N_7651);
nor UO_649 (O_649,N_8555,N_8221);
nand UO_650 (O_650,N_9330,N_8792);
nor UO_651 (O_651,N_8744,N_8883);
nor UO_652 (O_652,N_8595,N_9375);
or UO_653 (O_653,N_9842,N_8239);
nor UO_654 (O_654,N_8727,N_9634);
nor UO_655 (O_655,N_7570,N_9530);
nand UO_656 (O_656,N_8765,N_8367);
and UO_657 (O_657,N_9446,N_9847);
and UO_658 (O_658,N_8023,N_9438);
or UO_659 (O_659,N_8414,N_7807);
and UO_660 (O_660,N_8564,N_9207);
and UO_661 (O_661,N_9863,N_7783);
nor UO_662 (O_662,N_7780,N_8273);
nor UO_663 (O_663,N_9934,N_9243);
or UO_664 (O_664,N_8454,N_9855);
nand UO_665 (O_665,N_9879,N_8356);
nand UO_666 (O_666,N_8868,N_7844);
nand UO_667 (O_667,N_8117,N_8324);
nand UO_668 (O_668,N_8428,N_8306);
and UO_669 (O_669,N_7901,N_8404);
or UO_670 (O_670,N_8109,N_9014);
nand UO_671 (O_671,N_9313,N_7581);
or UO_672 (O_672,N_7804,N_7865);
nand UO_673 (O_673,N_7811,N_9336);
and UO_674 (O_674,N_8019,N_7972);
or UO_675 (O_675,N_9071,N_8845);
nand UO_676 (O_676,N_8919,N_8445);
or UO_677 (O_677,N_8786,N_9770);
nand UO_678 (O_678,N_7788,N_8691);
or UO_679 (O_679,N_8375,N_9696);
or UO_680 (O_680,N_9834,N_8703);
nand UO_681 (O_681,N_8224,N_8831);
nor UO_682 (O_682,N_8856,N_7878);
nor UO_683 (O_683,N_9420,N_9334);
nand UO_684 (O_684,N_8632,N_9514);
or UO_685 (O_685,N_8399,N_8406);
and UO_686 (O_686,N_9154,N_8422);
or UO_687 (O_687,N_9143,N_8193);
nand UO_688 (O_688,N_9571,N_9787);
and UO_689 (O_689,N_9220,N_8292);
and UO_690 (O_690,N_8048,N_8670);
or UO_691 (O_691,N_9361,N_7574);
or UO_692 (O_692,N_9954,N_8656);
and UO_693 (O_693,N_7853,N_9280);
nand UO_694 (O_694,N_8033,N_9392);
and UO_695 (O_695,N_8134,N_8689);
or UO_696 (O_696,N_8793,N_9079);
nor UO_697 (O_697,N_9833,N_9574);
and UO_698 (O_698,N_8572,N_8458);
and UO_699 (O_699,N_7726,N_9906);
and UO_700 (O_700,N_8469,N_7603);
nand UO_701 (O_701,N_8777,N_7625);
or UO_702 (O_702,N_9734,N_8008);
and UO_703 (O_703,N_9522,N_7989);
and UO_704 (O_704,N_9320,N_8613);
or UO_705 (O_705,N_9814,N_8925);
and UO_706 (O_706,N_7954,N_7634);
and UO_707 (O_707,N_7941,N_9045);
and UO_708 (O_708,N_9691,N_9795);
nand UO_709 (O_709,N_7944,N_8328);
or UO_710 (O_710,N_9030,N_9120);
nand UO_711 (O_711,N_9351,N_9886);
nand UO_712 (O_712,N_7704,N_8299);
and UO_713 (O_713,N_9562,N_8050);
nor UO_714 (O_714,N_8325,N_9089);
nand UO_715 (O_715,N_8270,N_8667);
nor UO_716 (O_716,N_8253,N_9830);
or UO_717 (O_717,N_7775,N_8101);
nor UO_718 (O_718,N_8153,N_9367);
and UO_719 (O_719,N_8343,N_8725);
nor UO_720 (O_720,N_8088,N_8884);
and UO_721 (O_721,N_8761,N_9615);
nand UO_722 (O_722,N_8166,N_7967);
or UO_723 (O_723,N_9729,N_8708);
nor UO_724 (O_724,N_8260,N_8830);
nand UO_725 (O_725,N_7643,N_9177);
nor UO_726 (O_726,N_7521,N_8750);
nand UO_727 (O_727,N_7690,N_9614);
nor UO_728 (O_728,N_7605,N_8012);
nor UO_729 (O_729,N_7617,N_8947);
nand UO_730 (O_730,N_8608,N_8599);
nand UO_731 (O_731,N_9738,N_9170);
nand UO_732 (O_732,N_7668,N_9860);
and UO_733 (O_733,N_7701,N_9096);
xnor UO_734 (O_734,N_9835,N_7520);
nand UO_735 (O_735,N_8218,N_9090);
or UO_736 (O_736,N_9246,N_8825);
nand UO_737 (O_737,N_9189,N_8813);
or UO_738 (O_738,N_8397,N_9999);
or UO_739 (O_739,N_8082,N_8282);
or UO_740 (O_740,N_7516,N_7767);
or UO_741 (O_741,N_9035,N_9810);
and UO_742 (O_742,N_9458,N_7641);
or UO_743 (O_743,N_8961,N_7627);
and UO_744 (O_744,N_8823,N_7610);
nor UO_745 (O_745,N_9663,N_8370);
or UO_746 (O_746,N_9836,N_7736);
or UO_747 (O_747,N_8588,N_8930);
and UO_748 (O_748,N_8544,N_9718);
and UO_749 (O_749,N_7653,N_8296);
nor UO_750 (O_750,N_7709,N_9398);
xor UO_751 (O_751,N_8164,N_9943);
nand UO_752 (O_752,N_9162,N_8316);
nand UO_753 (O_753,N_7917,N_9132);
or UO_754 (O_754,N_8352,N_9843);
or UO_755 (O_755,N_8668,N_7969);
nor UO_756 (O_756,N_9356,N_9668);
nand UO_757 (O_757,N_9214,N_8630);
nor UO_758 (O_758,N_8090,N_7815);
or UO_759 (O_759,N_7666,N_9173);
nor UO_760 (O_760,N_9982,N_9158);
or UO_761 (O_761,N_7949,N_9301);
nor UO_762 (O_762,N_9837,N_7863);
nand UO_763 (O_763,N_7808,N_8563);
or UO_764 (O_764,N_9311,N_9110);
or UO_765 (O_765,N_7770,N_9674);
nor UO_766 (O_766,N_7907,N_7655);
and UO_767 (O_767,N_8384,N_8530);
or UO_768 (O_768,N_7621,N_7659);
or UO_769 (O_769,N_8680,N_8345);
nand UO_770 (O_770,N_8184,N_9160);
nor UO_771 (O_771,N_9319,N_7626);
nand UO_772 (O_772,N_9882,N_9236);
xor UO_773 (O_773,N_9724,N_9355);
nor UO_774 (O_774,N_9117,N_9473);
and UO_775 (O_775,N_8644,N_8502);
or UO_776 (O_776,N_8525,N_9476);
nand UO_777 (O_777,N_9233,N_8078);
nand UO_778 (O_778,N_8511,N_9431);
or UO_779 (O_779,N_8248,N_9349);
or UO_780 (O_780,N_7712,N_9817);
nor UO_781 (O_781,N_7764,N_8035);
nor UO_782 (O_782,N_7596,N_8451);
and UO_783 (O_783,N_9974,N_9044);
nor UO_784 (O_784,N_9413,N_9478);
nor UO_785 (O_785,N_7505,N_8723);
and UO_786 (O_786,N_9360,N_9661);
or UO_787 (O_787,N_9590,N_9873);
or UO_788 (O_788,N_9548,N_7857);
nand UO_789 (O_789,N_9679,N_9751);
or UO_790 (O_790,N_9848,N_9291);
or UO_791 (O_791,N_7715,N_9839);
nand UO_792 (O_792,N_8435,N_8130);
or UO_793 (O_793,N_9901,N_9726);
nor UO_794 (O_794,N_8358,N_9493);
nor UO_795 (O_795,N_7660,N_8505);
or UO_796 (O_796,N_9204,N_7558);
or UO_797 (O_797,N_8478,N_9068);
nand UO_798 (O_798,N_7611,N_9288);
nor UO_799 (O_799,N_7754,N_7998);
nor UO_800 (O_800,N_9653,N_9707);
or UO_801 (O_801,N_8490,N_9728);
nor UO_802 (O_802,N_8293,N_9752);
nor UO_803 (O_803,N_7662,N_7928);
and UO_804 (O_804,N_8882,N_9405);
or UO_805 (O_805,N_9766,N_7931);
nand UO_806 (O_806,N_8281,N_9400);
or UO_807 (O_807,N_7716,N_8026);
or UO_808 (O_808,N_9060,N_8748);
nand UO_809 (O_809,N_7987,N_8769);
or UO_810 (O_810,N_9373,N_9540);
or UO_811 (O_811,N_7640,N_8429);
or UO_812 (O_812,N_9278,N_7905);
nand UO_813 (O_813,N_8009,N_9866);
nor UO_814 (O_814,N_8507,N_8175);
or UO_815 (O_815,N_7918,N_9047);
nor UO_816 (O_816,N_9048,N_8398);
nand UO_817 (O_817,N_9581,N_7899);
and UO_818 (O_818,N_7965,N_8954);
and UO_819 (O_819,N_9269,N_9937);
or UO_820 (O_820,N_9376,N_9976);
or UO_821 (O_821,N_8411,N_9652);
or UO_822 (O_822,N_9443,N_9890);
nor UO_823 (O_823,N_8172,N_9695);
nor UO_824 (O_824,N_8190,N_7670);
nor UO_825 (O_825,N_9195,N_9646);
or UO_826 (O_826,N_9171,N_9941);
nand UO_827 (O_827,N_9042,N_9404);
nand UO_828 (O_828,N_7982,N_9268);
nand UO_829 (O_829,N_7772,N_8523);
and UO_830 (O_830,N_7578,N_7958);
nor UO_831 (O_831,N_9872,N_8283);
nand UO_832 (O_832,N_8066,N_9617);
nand UO_833 (O_833,N_8386,N_9464);
nand UO_834 (O_834,N_7542,N_8022);
or UO_835 (O_835,N_7689,N_8695);
nor UO_836 (O_836,N_7765,N_7745);
nor UO_837 (O_837,N_8539,N_8731);
nand UO_838 (O_838,N_9215,N_9494);
or UO_839 (O_839,N_8733,N_8482);
or UO_840 (O_840,N_7594,N_9962);
and UO_841 (O_841,N_8486,N_9226);
nor UO_842 (O_842,N_8838,N_7760);
nor UO_843 (O_843,N_9502,N_7823);
and UO_844 (O_844,N_8739,N_7797);
or UO_845 (O_845,N_8442,N_9595);
nor UO_846 (O_846,N_9253,N_9914);
nand UO_847 (O_847,N_9904,N_9146);
or UO_848 (O_848,N_9781,N_8487);
or UO_849 (O_849,N_9056,N_7776);
nand UO_850 (O_850,N_9990,N_8204);
and UO_851 (O_851,N_8788,N_8133);
nand UO_852 (O_852,N_8933,N_9276);
or UO_853 (O_853,N_9101,N_9988);
nand UO_854 (O_854,N_8516,N_8364);
nand UO_855 (O_855,N_8917,N_9776);
or UO_856 (O_856,N_7904,N_7827);
nor UO_857 (O_857,N_9216,N_9435);
or UO_858 (O_858,N_7536,N_9864);
nor UO_859 (O_859,N_8393,N_8867);
or UO_860 (O_860,N_8489,N_8081);
and UO_861 (O_861,N_8906,N_8236);
nand UO_862 (O_862,N_7729,N_8982);
nor UO_863 (O_863,N_7546,N_8062);
and UO_864 (O_864,N_9161,N_8800);
or UO_865 (O_865,N_8051,N_8787);
nand UO_866 (O_866,N_7882,N_9222);
and UO_867 (O_867,N_9684,N_8092);
nand UO_868 (O_868,N_8196,N_9286);
or UO_869 (O_869,N_8149,N_8457);
and UO_870 (O_870,N_9757,N_9735);
and UO_871 (O_871,N_8250,N_7628);
or UO_872 (O_872,N_9576,N_7632);
and UO_873 (O_873,N_9687,N_7633);
nor UO_874 (O_874,N_7501,N_9921);
xnor UO_875 (O_875,N_8885,N_8898);
nand UO_876 (O_876,N_8290,N_9819);
xor UO_877 (O_877,N_9341,N_9479);
nor UO_878 (O_878,N_7648,N_9103);
and UO_879 (O_879,N_8120,N_9877);
nor UO_880 (O_880,N_8110,N_9647);
nand UO_881 (O_881,N_9328,N_9264);
nand UO_882 (O_882,N_9549,N_9386);
or UO_883 (O_883,N_9006,N_8686);
or UO_884 (O_884,N_7721,N_7737);
and UO_885 (O_885,N_9122,N_9644);
nand UO_886 (O_886,N_8408,N_7946);
nand UO_887 (O_887,N_7855,N_9665);
nor UO_888 (O_888,N_8918,N_9463);
and UO_889 (O_889,N_9909,N_8730);
nor UO_890 (O_890,N_8584,N_8387);
nor UO_891 (O_891,N_8591,N_7528);
and UO_892 (O_892,N_9387,N_9748);
nand UO_893 (O_893,N_8529,N_8228);
and UO_894 (O_894,N_9793,N_9032);
and UO_895 (O_895,N_8289,N_7886);
nand UO_896 (O_896,N_8326,N_9130);
and UO_897 (O_897,N_9929,N_9293);
nand UO_898 (O_898,N_7693,N_8191);
and UO_899 (O_899,N_7561,N_8103);
nand UO_900 (O_900,N_8678,N_9416);
and UO_901 (O_901,N_7801,N_9790);
and UO_902 (O_902,N_7604,N_9395);
and UO_903 (O_903,N_8601,N_9564);
or UO_904 (O_904,N_8795,N_9893);
nor UO_905 (O_905,N_8712,N_9221);
and UO_906 (O_906,N_8671,N_8660);
nor UO_907 (O_907,N_7672,N_7785);
nand UO_908 (O_908,N_8069,N_9245);
nand UO_909 (O_909,N_7802,N_9184);
or UO_910 (O_910,N_8437,N_8614);
or UO_911 (O_911,N_8928,N_9662);
nand UO_912 (O_912,N_8603,N_8068);
and UO_913 (O_913,N_8131,N_9996);
or UO_914 (O_914,N_9310,N_9275);
nor UO_915 (O_915,N_8298,N_9577);
and UO_916 (O_916,N_8017,N_8858);
or UO_917 (O_917,N_8911,N_8257);
or UO_918 (O_918,N_9631,N_7948);
nand UO_919 (O_919,N_8431,N_8237);
or UO_920 (O_920,N_8889,N_8448);
or UO_921 (O_921,N_9393,N_9654);
or UO_922 (O_922,N_9265,N_9678);
nand UO_923 (O_923,N_7671,N_7598);
and UO_924 (O_924,N_9936,N_8183);
nor UO_925 (O_925,N_8566,N_9845);
nor UO_926 (O_926,N_7753,N_8258);
or UO_927 (O_927,N_8330,N_8653);
nand UO_928 (O_928,N_9052,N_7500);
or UO_929 (O_929,N_7661,N_8254);
and UO_930 (O_930,N_7930,N_8093);
xor UO_931 (O_931,N_9401,N_8396);
or UO_932 (O_932,N_9299,N_8247);
nor UO_933 (O_933,N_9200,N_7824);
nand UO_934 (O_934,N_7695,N_9194);
and UO_935 (O_935,N_8853,N_9134);
xnor UO_936 (O_936,N_8637,N_7789);
nand UO_937 (O_937,N_7773,N_7576);
and UO_938 (O_938,N_9347,N_9106);
nor UO_939 (O_939,N_8702,N_8546);
xnor UO_940 (O_940,N_8135,N_8295);
nor UO_941 (O_941,N_8333,N_7974);
or UO_942 (O_942,N_8216,N_8677);
and UO_943 (O_943,N_9078,N_8568);
xnor UO_944 (O_944,N_8491,N_8924);
or UO_945 (O_945,N_8934,N_8063);
or UO_946 (O_946,N_8984,N_9991);
or UO_947 (O_947,N_8410,N_8772);
and UO_948 (O_948,N_9196,N_8267);
nand UO_949 (O_949,N_8824,N_9480);
and UO_950 (O_950,N_9978,N_8409);
nand UO_951 (O_951,N_9913,N_9598);
nor UO_952 (O_952,N_7544,N_8890);
nand UO_953 (O_953,N_9010,N_7524);
nor UO_954 (O_954,N_8872,N_8789);
nor UO_955 (O_955,N_7854,N_8056);
or UO_956 (O_956,N_8863,N_9187);
nand UO_957 (O_957,N_8522,N_9167);
nor UO_958 (O_958,N_8054,N_8126);
or UO_959 (O_959,N_8401,N_8559);
nand UO_960 (O_960,N_9876,N_7921);
nand UO_961 (O_961,N_7992,N_9454);
and UO_962 (O_962,N_9555,N_7936);
nand UO_963 (O_963,N_9166,N_8484);
nor UO_964 (O_964,N_7841,N_9067);
nand UO_965 (O_965,N_9875,N_7502);
nand UO_966 (O_966,N_8892,N_8636);
nand UO_967 (O_967,N_8503,N_9785);
and UO_968 (O_968,N_9114,N_8587);
nor UO_969 (O_969,N_8520,N_8440);
nand UO_970 (O_970,N_8674,N_9585);
and UO_971 (O_971,N_8163,N_8859);
nor UO_972 (O_972,N_8497,N_8935);
or UO_973 (O_973,N_7843,N_8500);
or UO_974 (O_974,N_9694,N_8626);
or UO_975 (O_975,N_8108,N_9667);
and UO_976 (O_976,N_7657,N_9437);
or UO_977 (O_977,N_7981,N_7889);
or UO_978 (O_978,N_9327,N_7758);
nor UO_979 (O_979,N_9427,N_9703);
nand UO_980 (O_980,N_9689,N_8347);
and UO_981 (O_981,N_7937,N_8168);
and UO_982 (O_982,N_9305,N_7983);
and UO_983 (O_983,N_8368,N_9102);
or UO_984 (O_984,N_7667,N_9164);
nand UO_985 (O_985,N_8735,N_8262);
and UO_986 (O_986,N_7916,N_8722);
and UO_987 (O_987,N_9570,N_9255);
and UO_988 (O_988,N_9841,N_8029);
or UO_989 (O_989,N_7706,N_7805);
and UO_990 (O_990,N_8537,N_8600);
and UO_991 (O_991,N_8724,N_9492);
nand UO_992 (O_992,N_8053,N_7995);
or UO_993 (O_993,N_7540,N_8754);
nor UO_994 (O_994,N_9340,N_8590);
and UO_995 (O_995,N_8524,N_8866);
xor UO_996 (O_996,N_8263,N_7619);
nor UO_997 (O_997,N_8449,N_8638);
nor UO_998 (O_998,N_9508,N_9015);
and UO_999 (O_999,N_8897,N_8277);
or UO_1000 (O_1000,N_8996,N_9645);
nor UO_1001 (O_1001,N_8909,N_9619);
nor UO_1002 (O_1002,N_8235,N_7568);
or UO_1003 (O_1003,N_9460,N_9922);
and UO_1004 (O_1004,N_9650,N_8197);
and UO_1005 (O_1005,N_9534,N_7947);
and UO_1006 (O_1006,N_9441,N_8552);
and UO_1007 (O_1007,N_9409,N_8843);
or UO_1008 (O_1008,N_9031,N_8052);
nor UO_1009 (O_1009,N_9604,N_8797);
nand UO_1010 (O_1010,N_8077,N_9894);
or UO_1011 (O_1011,N_9747,N_9603);
nand UO_1012 (O_1012,N_9960,N_9671);
and UO_1013 (O_1013,N_8353,N_7649);
and UO_1014 (O_1014,N_7794,N_9073);
nand UO_1015 (O_1015,N_8243,N_8005);
nor UO_1016 (O_1016,N_9002,N_8138);
and UO_1017 (O_1017,N_8213,N_8876);
and UO_1018 (O_1018,N_9808,N_8734);
and UO_1019 (O_1019,N_8318,N_8470);
and UO_1020 (O_1020,N_7769,N_9629);
nor UO_1021 (O_1021,N_7700,N_7951);
nor UO_1022 (O_1022,N_8441,N_8395);
nor UO_1023 (O_1023,N_9082,N_8821);
and UO_1024 (O_1024,N_9983,N_9252);
nor UO_1025 (O_1025,N_9368,N_9129);
nor UO_1026 (O_1026,N_9659,N_8351);
nand UO_1027 (O_1027,N_9169,N_8604);
and UO_1028 (O_1028,N_9714,N_9084);
and UO_1029 (O_1029,N_9528,N_9680);
nor UO_1030 (O_1030,N_9899,N_9971);
or UO_1031 (O_1031,N_8847,N_7999);
and UO_1032 (O_1032,N_9907,N_9527);
and UO_1033 (O_1033,N_9308,N_9669);
nor UO_1034 (O_1034,N_7828,N_9803);
and UO_1035 (O_1035,N_8311,N_9000);
or UO_1036 (O_1036,N_9865,N_9930);
nor UO_1037 (O_1037,N_9828,N_8272);
and UO_1038 (O_1038,N_9219,N_8495);
nand UO_1039 (O_1039,N_9229,N_9658);
xnor UO_1040 (O_1040,N_7738,N_9205);
nand UO_1041 (O_1041,N_8596,N_9765);
nor UO_1042 (O_1042,N_8585,N_9183);
nor UO_1043 (O_1043,N_9686,N_8669);
and UO_1044 (O_1044,N_9303,N_9529);
and UO_1045 (O_1045,N_8426,N_9244);
nor UO_1046 (O_1046,N_9559,N_9782);
xor UO_1047 (O_1047,N_8605,N_9412);
or UO_1048 (O_1048,N_7549,N_9175);
or UO_1049 (O_1049,N_8965,N_8483);
nor UO_1050 (O_1050,N_8509,N_9852);
nor UO_1051 (O_1051,N_9418,N_9016);
nor UO_1052 (O_1052,N_9086,N_9231);
nor UO_1053 (O_1053,N_9720,N_9038);
nor UO_1054 (O_1054,N_7952,N_7567);
nand UO_1055 (O_1055,N_8940,N_9649);
and UO_1056 (O_1056,N_7644,N_9722);
and UO_1057 (O_1057,N_8087,N_8804);
nand UO_1058 (O_1058,N_8238,N_9994);
nor UO_1059 (O_1059,N_8757,N_7777);
nand UO_1060 (O_1060,N_8575,N_9248);
or UO_1061 (O_1061,N_8766,N_8832);
xnor UO_1062 (O_1062,N_8365,N_9150);
nor UO_1063 (O_1063,N_7669,N_9541);
or UO_1064 (O_1064,N_8814,N_8116);
and UO_1065 (O_1065,N_9510,N_9784);
and UO_1066 (O_1066,N_9240,N_7782);
and UO_1067 (O_1067,N_9172,N_9821);
nor UO_1068 (O_1068,N_8045,N_8475);
and UO_1069 (O_1069,N_7607,N_8966);
or UO_1070 (O_1070,N_7663,N_8320);
or UO_1071 (O_1071,N_9777,N_7963);
nor UO_1072 (O_1072,N_7613,N_9425);
or UO_1073 (O_1073,N_7723,N_9433);
nor UO_1074 (O_1074,N_7973,N_8091);
nor UO_1075 (O_1075,N_8916,N_9059);
or UO_1076 (O_1076,N_8661,N_8031);
nand UO_1077 (O_1077,N_7840,N_9797);
nor UO_1078 (O_1078,N_8891,N_8400);
nand UO_1079 (O_1079,N_8479,N_8157);
nand UO_1080 (O_1080,N_9775,N_8014);
nor UO_1081 (O_1081,N_9039,N_7720);
nor UO_1082 (O_1082,N_9788,N_7902);
nor UO_1083 (O_1083,N_9362,N_7622);
nor UO_1084 (O_1084,N_9072,N_7538);
or UO_1085 (O_1085,N_8013,N_9887);
and UO_1086 (O_1086,N_9542,N_9013);
nor UO_1087 (O_1087,N_8499,N_9469);
xor UO_1088 (O_1088,N_8403,N_8208);
and UO_1089 (O_1089,N_8341,N_8779);
nand UO_1090 (O_1090,N_7515,N_9266);
nand UO_1091 (O_1091,N_8643,N_9111);
nand UO_1092 (O_1092,N_8747,N_8943);
or UO_1093 (O_1093,N_9706,N_9972);
or UO_1094 (O_1094,N_9444,N_9075);
nand UO_1095 (O_1095,N_8527,N_9448);
nor UO_1096 (O_1096,N_9756,N_9055);
nor UO_1097 (O_1097,N_9746,N_8802);
or UO_1098 (O_1098,N_8102,N_9791);
and UO_1099 (O_1099,N_9081,N_7582);
nor UO_1100 (O_1100,N_9798,N_9717);
nand UO_1101 (O_1101,N_9596,N_8629);
or UO_1102 (O_1102,N_9095,N_8659);
and UO_1103 (O_1103,N_9796,N_8547);
and UO_1104 (O_1104,N_8173,N_9385);
and UO_1105 (O_1105,N_8737,N_9306);
nor UO_1106 (O_1106,N_9025,N_9750);
nor UO_1107 (O_1107,N_7665,N_9333);
xnor UO_1108 (O_1108,N_9973,N_7511);
nand UO_1109 (O_1109,N_8178,N_8696);
or UO_1110 (O_1110,N_9759,N_7750);
nand UO_1111 (O_1111,N_9938,N_9369);
nor UO_1112 (O_1112,N_9980,N_8841);
nor UO_1113 (O_1113,N_7612,N_7735);
or UO_1114 (O_1114,N_9488,N_8271);
or UO_1115 (O_1115,N_7733,N_9867);
and UO_1116 (O_1116,N_9046,N_8681);
and UO_1117 (O_1117,N_7830,N_9523);
xnor UO_1118 (O_1118,N_7535,N_7883);
nand UO_1119 (O_1119,N_7831,N_8988);
nor UO_1120 (O_1120,N_8687,N_8177);
nor UO_1121 (O_1121,N_9235,N_8350);
nand UO_1122 (O_1122,N_8305,N_8624);
nor UO_1123 (O_1123,N_9363,N_7518);
nor UO_1124 (O_1124,N_8665,N_8024);
nor UO_1125 (O_1125,N_7722,N_9611);
nand UO_1126 (O_1126,N_9639,N_8553);
xor UO_1127 (O_1127,N_9358,N_9496);
nor UO_1128 (O_1128,N_9592,N_9366);
and UO_1129 (O_1129,N_9024,N_8374);
or UO_1130 (O_1130,N_9772,N_9575);
nand UO_1131 (O_1131,N_8065,N_9586);
nor UO_1132 (O_1132,N_8809,N_8620);
and UO_1133 (O_1133,N_7881,N_8309);
or UO_1134 (O_1134,N_9001,N_9935);
nand UO_1135 (O_1135,N_8803,N_9550);
and UO_1136 (O_1136,N_9762,N_9470);
nand UO_1137 (O_1137,N_9350,N_9185);
nor UO_1138 (O_1138,N_9354,N_8616);
nor UO_1139 (O_1139,N_9963,N_8059);
or UO_1140 (O_1140,N_8993,N_9064);
nand UO_1141 (O_1141,N_7933,N_9009);
and UO_1142 (O_1142,N_8880,N_7684);
nor UO_1143 (O_1143,N_8554,N_7953);
nand UO_1144 (O_1144,N_8436,N_7530);
nor UO_1145 (O_1145,N_8058,N_8738);
nand UO_1146 (O_1146,N_7658,N_8589);
and UO_1147 (O_1147,N_8782,N_9800);
or UO_1148 (O_1148,N_9713,N_7674);
nand UO_1149 (O_1149,N_7976,N_8957);
and UO_1150 (O_1150,N_8332,N_9099);
nand UO_1151 (O_1151,N_8819,N_9732);
nand UO_1152 (O_1152,N_7545,N_8245);
nand UO_1153 (O_1153,N_8922,N_7707);
or UO_1154 (O_1154,N_9918,N_9657);
nor UO_1155 (O_1155,N_9012,N_8690);
or UO_1156 (O_1156,N_8642,N_9606);
and UO_1157 (O_1157,N_8314,N_7915);
or UO_1158 (O_1158,N_8323,N_8132);
or UO_1159 (O_1159,N_7898,N_7512);
nand UO_1160 (O_1160,N_9442,N_9419);
nor UO_1161 (O_1161,N_8418,N_9727);
nand UO_1162 (O_1162,N_9335,N_7676);
or UO_1163 (O_1163,N_8121,N_7766);
nand UO_1164 (O_1164,N_8003,N_9892);
nand UO_1165 (O_1165,N_9908,N_8939);
nand UO_1166 (O_1166,N_8083,N_9149);
or UO_1167 (O_1167,N_8645,N_9804);
and UO_1168 (O_1168,N_8941,N_7970);
nor UO_1169 (O_1169,N_8692,N_8732);
nand UO_1170 (O_1170,N_9455,N_7909);
nand UO_1171 (O_1171,N_8301,N_9884);
nor UO_1172 (O_1172,N_9457,N_8001);
nor UO_1173 (O_1173,N_9871,N_8041);
and UO_1174 (O_1174,N_9088,N_9811);
and UO_1175 (O_1175,N_8209,N_8952);
nand UO_1176 (O_1176,N_8650,N_9672);
nor UO_1177 (O_1177,N_9208,N_8652);
and UO_1178 (O_1178,N_9202,N_8805);
xor UO_1179 (O_1179,N_9343,N_7867);
or UO_1180 (O_1180,N_7922,N_8199);
or UO_1181 (O_1181,N_8040,N_9137);
nor UO_1182 (O_1182,N_8697,N_9736);
and UO_1183 (O_1183,N_7924,N_8528);
or UO_1184 (O_1184,N_8371,N_8150);
or UO_1185 (O_1185,N_7747,N_9942);
and UO_1186 (O_1186,N_8212,N_9874);
nand UO_1187 (O_1187,N_8852,N_9339);
nor UO_1188 (O_1188,N_9809,N_9561);
nand UO_1189 (O_1189,N_8861,N_9232);
and UO_1190 (O_1190,N_8875,N_8342);
nand UO_1191 (O_1191,N_8913,N_9011);
or UO_1192 (O_1192,N_8143,N_8640);
and UO_1193 (O_1193,N_8240,N_9126);
or UO_1194 (O_1194,N_8444,N_9148);
nor UO_1195 (O_1195,N_9979,N_9295);
nand UO_1196 (O_1196,N_9947,N_8806);
or UO_1197 (O_1197,N_8682,N_9135);
or UO_1198 (O_1198,N_9794,N_9651);
and UO_1199 (O_1199,N_8771,N_7945);
nor UO_1200 (O_1200,N_8202,N_7868);
and UO_1201 (O_1201,N_8115,N_9105);
or UO_1202 (O_1202,N_8615,N_8159);
or UO_1203 (O_1203,N_9294,N_9593);
and UO_1204 (O_1204,N_8200,N_7851);
nor UO_1205 (O_1205,N_9698,N_9307);
and UO_1206 (O_1206,N_7778,N_8039);
or UO_1207 (O_1207,N_8182,N_8763);
nand UO_1208 (O_1208,N_8095,N_8683);
xor UO_1209 (O_1209,N_9824,N_8047);
nor UO_1210 (O_1210,N_9944,N_8385);
or UO_1211 (O_1211,N_9545,N_8827);
xor UO_1212 (O_1212,N_8249,N_7525);
or UO_1213 (O_1213,N_7508,N_9332);
or UO_1214 (O_1214,N_8203,N_9600);
or UO_1215 (O_1215,N_8526,N_9279);
or UO_1216 (O_1216,N_9017,N_9085);
nand UO_1217 (O_1217,N_9902,N_9378);
nand UO_1218 (O_1218,N_9946,N_9805);
xor UO_1219 (O_1219,N_7557,N_8378);
nand UO_1220 (O_1220,N_8969,N_9337);
or UO_1221 (O_1221,N_9217,N_9799);
nand UO_1222 (O_1222,N_9789,N_8379);
or UO_1223 (O_1223,N_8226,N_9816);
and UO_1224 (O_1224,N_7673,N_9881);
nand UO_1225 (O_1225,N_8851,N_7939);
or UO_1226 (O_1226,N_8055,N_7984);
nor UO_1227 (O_1227,N_8666,N_9737);
nor UO_1228 (O_1228,N_8259,N_8815);
and UO_1229 (O_1229,N_8981,N_8466);
xnor UO_1230 (O_1230,N_7942,N_8767);
nand UO_1231 (O_1231,N_9832,N_7932);
or UO_1232 (O_1232,N_7822,N_8264);
nand UO_1233 (O_1233,N_9151,N_9846);
and UO_1234 (O_1234,N_9190,N_8446);
xor UO_1235 (O_1235,N_8946,N_7786);
and UO_1236 (O_1236,N_8096,N_9557);
or UO_1237 (O_1237,N_8344,N_9897);
or UO_1238 (O_1238,N_8284,N_8043);
nor UO_1239 (O_1239,N_8621,N_9309);
or UO_1240 (O_1240,N_9768,N_9352);
nand UO_1241 (O_1241,N_8312,N_8833);
nor UO_1242 (O_1242,N_8488,N_7816);
nor UO_1243 (O_1243,N_8222,N_7522);
nand UO_1244 (O_1244,N_9197,N_9506);
and UO_1245 (O_1245,N_8331,N_7971);
and UO_1246 (O_1246,N_7858,N_8510);
or UO_1247 (O_1247,N_9238,N_9822);
or UO_1248 (O_1248,N_9878,N_9353);
and UO_1249 (O_1249,N_7908,N_9741);
or UO_1250 (O_1250,N_7671,N_8787);
nand UO_1251 (O_1251,N_8188,N_8824);
or UO_1252 (O_1252,N_9802,N_9549);
and UO_1253 (O_1253,N_7760,N_8592);
nand UO_1254 (O_1254,N_8476,N_9753);
and UO_1255 (O_1255,N_8131,N_7756);
and UO_1256 (O_1256,N_9321,N_8351);
nor UO_1257 (O_1257,N_9575,N_8095);
and UO_1258 (O_1258,N_7565,N_8865);
or UO_1259 (O_1259,N_8533,N_7655);
nor UO_1260 (O_1260,N_9951,N_9807);
nor UO_1261 (O_1261,N_9213,N_8537);
nand UO_1262 (O_1262,N_9855,N_8923);
or UO_1263 (O_1263,N_9881,N_9641);
nor UO_1264 (O_1264,N_8947,N_7930);
nand UO_1265 (O_1265,N_9608,N_9342);
nor UO_1266 (O_1266,N_7607,N_7810);
and UO_1267 (O_1267,N_8949,N_8736);
and UO_1268 (O_1268,N_7810,N_9168);
nor UO_1269 (O_1269,N_8099,N_9161);
and UO_1270 (O_1270,N_7732,N_7703);
or UO_1271 (O_1271,N_8116,N_8148);
or UO_1272 (O_1272,N_9570,N_8478);
and UO_1273 (O_1273,N_7958,N_9015);
xnor UO_1274 (O_1274,N_9986,N_9877);
and UO_1275 (O_1275,N_8143,N_7859);
or UO_1276 (O_1276,N_9954,N_8093);
and UO_1277 (O_1277,N_9004,N_9732);
and UO_1278 (O_1278,N_9417,N_8371);
or UO_1279 (O_1279,N_7972,N_9654);
nand UO_1280 (O_1280,N_7963,N_7745);
nor UO_1281 (O_1281,N_8132,N_7727);
nand UO_1282 (O_1282,N_7585,N_8324);
and UO_1283 (O_1283,N_9218,N_7854);
or UO_1284 (O_1284,N_8590,N_8712);
and UO_1285 (O_1285,N_8431,N_8317);
or UO_1286 (O_1286,N_9831,N_9527);
nor UO_1287 (O_1287,N_8020,N_9455);
or UO_1288 (O_1288,N_9794,N_8456);
nand UO_1289 (O_1289,N_7586,N_7650);
nor UO_1290 (O_1290,N_8970,N_8179);
or UO_1291 (O_1291,N_9325,N_9736);
nand UO_1292 (O_1292,N_8168,N_9747);
and UO_1293 (O_1293,N_9271,N_8638);
xnor UO_1294 (O_1294,N_9369,N_9407);
or UO_1295 (O_1295,N_9335,N_7580);
and UO_1296 (O_1296,N_7539,N_8928);
nand UO_1297 (O_1297,N_7579,N_9845);
nor UO_1298 (O_1298,N_9603,N_9889);
xor UO_1299 (O_1299,N_8514,N_7507);
nor UO_1300 (O_1300,N_9423,N_8211);
nand UO_1301 (O_1301,N_8550,N_9178);
nor UO_1302 (O_1302,N_9960,N_9183);
nor UO_1303 (O_1303,N_7993,N_9268);
nor UO_1304 (O_1304,N_7851,N_7996);
or UO_1305 (O_1305,N_7847,N_8649);
and UO_1306 (O_1306,N_8452,N_9799);
nor UO_1307 (O_1307,N_8981,N_8117);
and UO_1308 (O_1308,N_8462,N_9598);
nand UO_1309 (O_1309,N_8691,N_8593);
nand UO_1310 (O_1310,N_9835,N_9790);
and UO_1311 (O_1311,N_8633,N_9915);
nor UO_1312 (O_1312,N_8611,N_8674);
and UO_1313 (O_1313,N_9163,N_8067);
nand UO_1314 (O_1314,N_9350,N_9956);
nor UO_1315 (O_1315,N_9518,N_9547);
nand UO_1316 (O_1316,N_9848,N_9909);
xnor UO_1317 (O_1317,N_9511,N_7903);
nor UO_1318 (O_1318,N_9640,N_9980);
nand UO_1319 (O_1319,N_8596,N_8116);
and UO_1320 (O_1320,N_8108,N_7671);
nand UO_1321 (O_1321,N_7737,N_8936);
and UO_1322 (O_1322,N_8029,N_7585);
or UO_1323 (O_1323,N_9026,N_8049);
or UO_1324 (O_1324,N_8367,N_8060);
nor UO_1325 (O_1325,N_8460,N_9456);
or UO_1326 (O_1326,N_9940,N_9840);
nand UO_1327 (O_1327,N_9372,N_7850);
nor UO_1328 (O_1328,N_9319,N_8040);
nor UO_1329 (O_1329,N_8976,N_8119);
and UO_1330 (O_1330,N_7669,N_8507);
nor UO_1331 (O_1331,N_8393,N_8134);
nand UO_1332 (O_1332,N_9422,N_7868);
or UO_1333 (O_1333,N_8999,N_8942);
or UO_1334 (O_1334,N_8274,N_9630);
nand UO_1335 (O_1335,N_9352,N_7565);
nand UO_1336 (O_1336,N_7532,N_8110);
and UO_1337 (O_1337,N_9030,N_9602);
nand UO_1338 (O_1338,N_7726,N_8915);
or UO_1339 (O_1339,N_8955,N_9476);
nand UO_1340 (O_1340,N_7891,N_8664);
nor UO_1341 (O_1341,N_8707,N_8532);
and UO_1342 (O_1342,N_8694,N_8216);
nor UO_1343 (O_1343,N_9511,N_9036);
and UO_1344 (O_1344,N_9164,N_8403);
and UO_1345 (O_1345,N_9897,N_8326);
nand UO_1346 (O_1346,N_9462,N_9051);
nor UO_1347 (O_1347,N_8559,N_7721);
or UO_1348 (O_1348,N_8886,N_7920);
or UO_1349 (O_1349,N_8609,N_9245);
nor UO_1350 (O_1350,N_9720,N_8515);
nand UO_1351 (O_1351,N_8167,N_8760);
nor UO_1352 (O_1352,N_8330,N_8089);
nand UO_1353 (O_1353,N_9323,N_9147);
and UO_1354 (O_1354,N_9082,N_9182);
or UO_1355 (O_1355,N_8484,N_9540);
and UO_1356 (O_1356,N_8003,N_7753);
xnor UO_1357 (O_1357,N_9425,N_8845);
nand UO_1358 (O_1358,N_8357,N_8978);
and UO_1359 (O_1359,N_8789,N_8251);
nand UO_1360 (O_1360,N_9553,N_8854);
nand UO_1361 (O_1361,N_9333,N_8445);
and UO_1362 (O_1362,N_9769,N_9433);
nand UO_1363 (O_1363,N_8074,N_8715);
nand UO_1364 (O_1364,N_9547,N_9673);
and UO_1365 (O_1365,N_8865,N_9709);
or UO_1366 (O_1366,N_7969,N_8951);
or UO_1367 (O_1367,N_9919,N_9810);
nor UO_1368 (O_1368,N_8233,N_8129);
nor UO_1369 (O_1369,N_7602,N_9131);
or UO_1370 (O_1370,N_9744,N_9933);
nand UO_1371 (O_1371,N_8322,N_8426);
or UO_1372 (O_1372,N_8252,N_8060);
or UO_1373 (O_1373,N_8905,N_9996);
nand UO_1374 (O_1374,N_8780,N_8776);
nand UO_1375 (O_1375,N_8883,N_7999);
or UO_1376 (O_1376,N_7650,N_9291);
nor UO_1377 (O_1377,N_9542,N_9436);
nand UO_1378 (O_1378,N_9374,N_8593);
nand UO_1379 (O_1379,N_9387,N_8326);
and UO_1380 (O_1380,N_8916,N_8128);
nor UO_1381 (O_1381,N_8494,N_7945);
or UO_1382 (O_1382,N_9321,N_9281);
nand UO_1383 (O_1383,N_8370,N_9848);
nand UO_1384 (O_1384,N_7614,N_9442);
nor UO_1385 (O_1385,N_7866,N_9905);
and UO_1386 (O_1386,N_7781,N_9951);
or UO_1387 (O_1387,N_8057,N_8527);
or UO_1388 (O_1388,N_8517,N_7903);
and UO_1389 (O_1389,N_8935,N_8113);
nor UO_1390 (O_1390,N_7533,N_9080);
and UO_1391 (O_1391,N_8093,N_8860);
nand UO_1392 (O_1392,N_7788,N_9972);
nand UO_1393 (O_1393,N_8458,N_8580);
nor UO_1394 (O_1394,N_9910,N_9007);
nor UO_1395 (O_1395,N_9365,N_8875);
or UO_1396 (O_1396,N_9848,N_8831);
nand UO_1397 (O_1397,N_7701,N_9734);
or UO_1398 (O_1398,N_9405,N_9087);
nand UO_1399 (O_1399,N_9069,N_7565);
nor UO_1400 (O_1400,N_9586,N_8377);
and UO_1401 (O_1401,N_8455,N_8180);
nor UO_1402 (O_1402,N_8581,N_9686);
and UO_1403 (O_1403,N_8576,N_8535);
nor UO_1404 (O_1404,N_9445,N_9328);
xor UO_1405 (O_1405,N_9407,N_8842);
xor UO_1406 (O_1406,N_8604,N_8236);
and UO_1407 (O_1407,N_8065,N_8890);
nand UO_1408 (O_1408,N_8696,N_9686);
or UO_1409 (O_1409,N_7667,N_9117);
and UO_1410 (O_1410,N_7652,N_9737);
xnor UO_1411 (O_1411,N_8506,N_9769);
and UO_1412 (O_1412,N_8119,N_7667);
or UO_1413 (O_1413,N_9219,N_7800);
and UO_1414 (O_1414,N_9226,N_9662);
or UO_1415 (O_1415,N_7618,N_8405);
xnor UO_1416 (O_1416,N_7966,N_7538);
and UO_1417 (O_1417,N_8416,N_9977);
nand UO_1418 (O_1418,N_8658,N_9415);
nand UO_1419 (O_1419,N_9897,N_7742);
nor UO_1420 (O_1420,N_7612,N_8773);
nor UO_1421 (O_1421,N_9428,N_8264);
nor UO_1422 (O_1422,N_8711,N_8109);
nor UO_1423 (O_1423,N_9892,N_9107);
nor UO_1424 (O_1424,N_9497,N_7605);
and UO_1425 (O_1425,N_9715,N_8395);
and UO_1426 (O_1426,N_9636,N_8802);
and UO_1427 (O_1427,N_9383,N_9838);
or UO_1428 (O_1428,N_8409,N_8635);
nand UO_1429 (O_1429,N_9866,N_9912);
and UO_1430 (O_1430,N_8557,N_8154);
or UO_1431 (O_1431,N_9040,N_7841);
nand UO_1432 (O_1432,N_8244,N_8511);
nand UO_1433 (O_1433,N_9693,N_8035);
and UO_1434 (O_1434,N_8562,N_9405);
nand UO_1435 (O_1435,N_8509,N_8057);
or UO_1436 (O_1436,N_7536,N_7797);
or UO_1437 (O_1437,N_9573,N_9112);
xor UO_1438 (O_1438,N_8432,N_7820);
nor UO_1439 (O_1439,N_7937,N_7975);
or UO_1440 (O_1440,N_8705,N_7739);
nand UO_1441 (O_1441,N_8089,N_9970);
nand UO_1442 (O_1442,N_9017,N_8153);
and UO_1443 (O_1443,N_9968,N_8791);
nand UO_1444 (O_1444,N_8405,N_9633);
nand UO_1445 (O_1445,N_8572,N_9364);
nand UO_1446 (O_1446,N_8758,N_8010);
nand UO_1447 (O_1447,N_9804,N_9871);
nand UO_1448 (O_1448,N_8145,N_8392);
nor UO_1449 (O_1449,N_9449,N_8731);
nand UO_1450 (O_1450,N_9485,N_8210);
or UO_1451 (O_1451,N_9301,N_9745);
nand UO_1452 (O_1452,N_8940,N_7729);
or UO_1453 (O_1453,N_7749,N_8579);
nor UO_1454 (O_1454,N_7630,N_9160);
and UO_1455 (O_1455,N_9228,N_8132);
nor UO_1456 (O_1456,N_9413,N_9461);
and UO_1457 (O_1457,N_8478,N_7897);
and UO_1458 (O_1458,N_7520,N_8633);
nand UO_1459 (O_1459,N_9804,N_9823);
nor UO_1460 (O_1460,N_8574,N_7715);
xnor UO_1461 (O_1461,N_8078,N_9977);
xnor UO_1462 (O_1462,N_7880,N_8741);
nand UO_1463 (O_1463,N_8212,N_8148);
nand UO_1464 (O_1464,N_7521,N_7878);
nand UO_1465 (O_1465,N_8592,N_9776);
nand UO_1466 (O_1466,N_9445,N_8001);
nand UO_1467 (O_1467,N_7770,N_9871);
nand UO_1468 (O_1468,N_8823,N_9294);
nand UO_1469 (O_1469,N_9723,N_7773);
and UO_1470 (O_1470,N_9063,N_8478);
and UO_1471 (O_1471,N_7873,N_8204);
nand UO_1472 (O_1472,N_7535,N_8826);
nand UO_1473 (O_1473,N_9360,N_9060);
xnor UO_1474 (O_1474,N_8701,N_9785);
nand UO_1475 (O_1475,N_7858,N_8640);
xnor UO_1476 (O_1476,N_9323,N_9666);
or UO_1477 (O_1477,N_8315,N_8738);
nor UO_1478 (O_1478,N_8679,N_9485);
and UO_1479 (O_1479,N_9643,N_9889);
or UO_1480 (O_1480,N_9920,N_7882);
nand UO_1481 (O_1481,N_9819,N_7899);
nand UO_1482 (O_1482,N_9680,N_9892);
and UO_1483 (O_1483,N_9134,N_8777);
and UO_1484 (O_1484,N_8319,N_8072);
nor UO_1485 (O_1485,N_9628,N_9177);
or UO_1486 (O_1486,N_8675,N_8116);
nand UO_1487 (O_1487,N_8333,N_8962);
or UO_1488 (O_1488,N_8270,N_8616);
nor UO_1489 (O_1489,N_8632,N_9259);
and UO_1490 (O_1490,N_7696,N_9084);
or UO_1491 (O_1491,N_8732,N_9998);
nor UO_1492 (O_1492,N_7633,N_8689);
and UO_1493 (O_1493,N_9764,N_8502);
or UO_1494 (O_1494,N_9557,N_9346);
or UO_1495 (O_1495,N_8784,N_9518);
and UO_1496 (O_1496,N_9220,N_9290);
nor UO_1497 (O_1497,N_8512,N_8856);
or UO_1498 (O_1498,N_8078,N_8877);
or UO_1499 (O_1499,N_8466,N_8586);
endmodule