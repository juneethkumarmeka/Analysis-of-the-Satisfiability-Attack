module basic_2000_20000_2500_10_levels_1xor_7(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999;
and U0 (N_0,In_1249,In_1470);
nor U1 (N_1,In_292,In_17);
or U2 (N_2,In_0,In_1481);
and U3 (N_3,In_318,In_1520);
and U4 (N_4,In_1033,In_1706);
nor U5 (N_5,In_1143,In_1908);
nor U6 (N_6,In_1058,In_791);
nand U7 (N_7,In_1190,In_521);
and U8 (N_8,In_271,In_336);
nand U9 (N_9,In_1675,In_1133);
and U10 (N_10,In_1756,In_1251);
and U11 (N_11,In_1105,In_342);
or U12 (N_12,In_1808,In_26);
or U13 (N_13,In_658,In_619);
and U14 (N_14,In_847,In_1055);
nor U15 (N_15,In_1552,In_437);
or U16 (N_16,In_1676,In_747);
nand U17 (N_17,In_1708,In_43);
or U18 (N_18,In_535,In_741);
nand U19 (N_19,In_345,In_1902);
or U20 (N_20,In_740,In_1715);
or U21 (N_21,In_327,In_1483);
nor U22 (N_22,In_766,In_1303);
nor U23 (N_23,In_1726,In_131);
nor U24 (N_24,In_659,In_1496);
or U25 (N_25,In_93,In_1005);
and U26 (N_26,In_146,In_1168);
nand U27 (N_27,In_963,In_715);
and U28 (N_28,In_1090,In_1984);
nand U29 (N_29,In_1876,In_514);
or U30 (N_30,In_1311,In_1751);
and U31 (N_31,In_729,In_679);
and U32 (N_32,In_153,In_636);
or U33 (N_33,In_1772,In_133);
or U34 (N_34,In_98,In_485);
and U35 (N_35,In_1639,In_995);
and U36 (N_36,In_260,In_800);
and U37 (N_37,In_1500,In_630);
and U38 (N_38,In_194,In_1445);
xnor U39 (N_39,In_114,In_230);
nor U40 (N_40,In_1009,In_383);
xor U41 (N_41,In_868,In_382);
xor U42 (N_42,In_1854,In_991);
nor U43 (N_43,In_386,In_1697);
nor U44 (N_44,In_1926,In_1887);
xor U45 (N_45,In_1124,In_655);
nor U46 (N_46,In_421,In_1084);
or U47 (N_47,In_662,In_145);
nand U48 (N_48,In_419,In_539);
nand U49 (N_49,In_1664,In_1636);
nor U50 (N_50,In_712,In_1172);
nor U51 (N_51,In_1346,In_478);
and U52 (N_52,In_723,In_1853);
nor U53 (N_53,In_1580,In_1779);
or U54 (N_54,In_1948,In_126);
nor U55 (N_55,In_241,In_646);
nand U56 (N_56,In_393,In_798);
or U57 (N_57,In_1237,In_1645);
nand U58 (N_58,In_304,In_1831);
nand U59 (N_59,In_1391,In_900);
nor U60 (N_60,In_1007,In_1243);
and U61 (N_61,In_1551,In_795);
and U62 (N_62,In_918,In_1129);
and U63 (N_63,In_276,In_1492);
nand U64 (N_64,In_545,In_610);
nor U65 (N_65,In_772,In_1582);
or U66 (N_66,In_1620,In_15);
nor U67 (N_67,In_1031,In_1755);
and U68 (N_68,In_1915,In_310);
nor U69 (N_69,In_1283,In_598);
nor U70 (N_70,In_1192,In_1765);
nand U71 (N_71,In_838,In_1263);
or U72 (N_72,In_1858,In_1712);
nor U73 (N_73,In_41,In_1187);
nor U74 (N_74,In_87,In_1486);
and U75 (N_75,In_623,In_816);
nand U76 (N_76,In_4,In_1231);
nand U77 (N_77,In_986,In_1424);
and U78 (N_78,In_138,In_1724);
nand U79 (N_79,In_1956,In_1619);
nand U80 (N_80,In_496,In_877);
nand U81 (N_81,In_261,In_1438);
nor U82 (N_82,In_1489,In_1701);
nand U83 (N_83,In_89,In_568);
and U84 (N_84,In_884,In_1986);
and U85 (N_85,In_1484,In_61);
xor U86 (N_86,In_1562,In_1678);
and U87 (N_87,In_1611,In_746);
nand U88 (N_88,In_82,In_1316);
or U89 (N_89,In_675,In_811);
nand U90 (N_90,In_760,In_1434);
nand U91 (N_91,In_66,In_1212);
and U92 (N_92,In_890,In_563);
nor U93 (N_93,In_1314,In_391);
nand U94 (N_94,In_1906,In_1721);
or U95 (N_95,In_1768,In_1790);
or U96 (N_96,In_924,In_657);
and U97 (N_97,In_1688,In_1178);
nand U98 (N_98,In_628,In_745);
and U99 (N_99,In_885,In_1602);
and U100 (N_100,In_70,In_1803);
and U101 (N_101,In_992,In_287);
or U102 (N_102,In_1725,In_1837);
or U103 (N_103,In_463,In_286);
and U104 (N_104,In_1279,In_1974);
and U105 (N_105,In_916,In_865);
and U106 (N_106,In_111,In_953);
nand U107 (N_107,In_1487,In_1420);
nor U108 (N_108,In_631,In_1397);
nand U109 (N_109,In_987,In_852);
and U110 (N_110,In_1820,In_1878);
or U111 (N_111,In_569,In_961);
or U112 (N_112,In_1817,In_1430);
and U113 (N_113,In_688,In_1855);
nand U114 (N_114,In_1656,In_719);
or U115 (N_115,In_403,In_605);
and U116 (N_116,In_1449,In_2);
and U117 (N_117,In_1441,In_633);
or U118 (N_118,In_978,In_667);
nor U119 (N_119,In_1624,In_578);
or U120 (N_120,In_673,In_141);
or U121 (N_121,In_860,In_209);
nand U122 (N_122,In_1082,In_224);
nand U123 (N_123,In_459,In_1793);
xnor U124 (N_124,In_246,In_1250);
nand U125 (N_125,In_759,In_405);
or U126 (N_126,In_509,In_1258);
or U127 (N_127,In_58,In_594);
and U128 (N_128,In_820,In_222);
nor U129 (N_129,In_892,In_532);
and U130 (N_130,In_1961,In_653);
or U131 (N_131,In_743,In_1147);
or U132 (N_132,In_210,In_1788);
nor U133 (N_133,In_39,In_505);
and U134 (N_134,In_1839,In_72);
and U135 (N_135,In_666,In_238);
and U136 (N_136,In_1248,In_1600);
or U137 (N_137,In_878,In_122);
or U138 (N_138,In_1658,In_1633);
and U139 (N_139,In_1215,In_758);
nor U140 (N_140,In_1392,In_748);
and U141 (N_141,In_221,In_526);
and U142 (N_142,In_768,In_474);
or U143 (N_143,In_25,In_600);
and U144 (N_144,In_1920,In_1293);
nand U145 (N_145,In_508,In_450);
nor U146 (N_146,In_709,In_1732);
and U147 (N_147,In_45,In_1262);
and U148 (N_148,In_552,In_1466);
and U149 (N_149,In_48,In_1395);
and U150 (N_150,In_399,In_1744);
nor U151 (N_151,In_449,In_239);
or U152 (N_152,In_889,In_179);
nor U153 (N_153,In_972,In_1485);
or U154 (N_154,In_35,In_1269);
nand U155 (N_155,In_1205,In_1347);
and U156 (N_156,In_529,In_27);
nand U157 (N_157,In_1669,In_1569);
and U158 (N_158,In_173,In_412);
or U159 (N_159,In_803,In_447);
nor U160 (N_160,In_429,In_911);
nand U161 (N_161,In_118,In_189);
nand U162 (N_162,In_1535,In_1474);
nand U163 (N_163,In_997,In_394);
or U164 (N_164,In_988,In_81);
nor U165 (N_165,In_951,In_1581);
or U166 (N_166,In_1657,In_190);
nand U167 (N_167,In_1864,In_651);
nor U168 (N_168,In_67,In_1812);
nand U169 (N_169,In_1370,In_1412);
nand U170 (N_170,In_197,In_1561);
nand U171 (N_171,In_1219,In_255);
nand U172 (N_172,In_1478,In_540);
and U173 (N_173,In_1904,In_895);
nand U174 (N_174,In_1153,In_841);
and U175 (N_175,In_1067,In_786);
and U176 (N_176,In_710,In_302);
nor U177 (N_177,In_1975,In_320);
nand U178 (N_178,In_1748,In_379);
and U179 (N_179,In_845,In_192);
or U180 (N_180,In_732,In_827);
and U181 (N_181,In_548,In_999);
or U182 (N_182,In_1696,In_781);
or U183 (N_183,In_418,In_368);
or U184 (N_184,In_1140,In_19);
nor U185 (N_185,In_1197,In_400);
and U186 (N_186,In_49,In_1044);
nand U187 (N_187,In_1185,In_641);
nand U188 (N_188,In_595,In_677);
and U189 (N_189,In_549,In_1589);
or U190 (N_190,In_182,In_1849);
or U191 (N_191,In_125,In_1013);
nand U192 (N_192,In_909,In_780);
nor U193 (N_193,In_1368,In_1157);
nand U194 (N_194,In_1637,In_1548);
and U195 (N_195,In_519,In_353);
nor U196 (N_196,In_1266,In_1415);
or U197 (N_197,In_120,In_958);
or U198 (N_198,In_1149,In_1861);
nand U199 (N_199,In_971,In_269);
or U200 (N_200,In_1665,In_152);
and U201 (N_201,In_1587,In_1931);
nor U202 (N_202,In_1951,In_1081);
or U203 (N_203,In_1816,In_1450);
nand U204 (N_204,In_714,In_477);
or U205 (N_205,In_778,In_763);
and U206 (N_206,In_177,In_1737);
or U207 (N_207,In_1881,In_1355);
xor U208 (N_208,In_1608,In_861);
nor U209 (N_209,In_728,In_1138);
or U210 (N_210,In_476,In_1700);
nand U211 (N_211,In_1893,In_172);
nor U212 (N_212,In_1076,In_590);
nor U213 (N_213,In_356,In_1718);
nor U214 (N_214,In_409,In_425);
nor U215 (N_215,In_830,In_1462);
and U216 (N_216,In_1448,In_1834);
and U217 (N_217,In_465,In_661);
and U218 (N_218,In_471,In_178);
or U219 (N_219,In_1773,In_1301);
nand U220 (N_220,In_1331,In_939);
nand U221 (N_221,In_231,In_1417);
nor U222 (N_222,In_490,In_1338);
and U223 (N_223,In_1505,In_585);
nand U224 (N_224,In_637,In_165);
xnor U225 (N_225,In_1814,In_649);
nand U226 (N_226,In_1091,In_1358);
and U227 (N_227,In_1194,In_775);
nor U228 (N_228,In_357,In_245);
and U229 (N_229,In_1384,In_910);
nand U230 (N_230,In_829,In_1119);
nand U231 (N_231,In_375,In_366);
nor U232 (N_232,In_1195,In_160);
nor U233 (N_233,In_1169,In_305);
or U234 (N_234,In_1042,In_322);
nor U235 (N_235,In_1239,In_851);
nor U236 (N_236,In_12,In_46);
nor U237 (N_237,In_1959,In_1443);
nor U238 (N_238,In_794,In_3);
and U239 (N_239,In_60,In_301);
nor U240 (N_240,In_1928,In_614);
or U241 (N_241,In_325,In_1776);
nor U242 (N_242,In_882,In_1813);
nor U243 (N_243,In_640,In_1380);
nand U244 (N_244,In_1795,In_1519);
or U245 (N_245,In_55,In_134);
and U246 (N_246,In_581,In_1026);
nand U247 (N_247,In_1317,In_94);
nand U248 (N_248,In_557,In_524);
and U249 (N_249,In_1378,In_592);
nor U250 (N_250,In_749,In_950);
and U251 (N_251,In_371,In_1404);
or U252 (N_252,In_1334,In_634);
or U253 (N_253,In_135,In_831);
nor U254 (N_254,In_776,In_14);
and U255 (N_255,In_1739,In_1039);
nor U256 (N_256,In_439,In_248);
or U257 (N_257,In_792,In_112);
nor U258 (N_258,In_299,In_456);
nand U259 (N_259,In_343,In_110);
and U260 (N_260,In_683,In_905);
nand U261 (N_261,In_159,In_1764);
nor U262 (N_262,In_180,In_9);
or U263 (N_263,In_1894,In_249);
or U264 (N_264,In_123,In_1660);
nor U265 (N_265,In_589,In_1597);
nor U266 (N_266,In_1429,In_1282);
nand U267 (N_267,In_788,In_1092);
nand U268 (N_268,In_888,In_1782);
nand U269 (N_269,In_1069,In_870);
and U270 (N_270,In_1668,In_989);
nand U271 (N_271,In_1118,In_1040);
and U272 (N_272,In_1122,In_1145);
nand U273 (N_273,In_1944,In_143);
nor U274 (N_274,In_452,In_654);
nor U275 (N_275,In_1369,In_523);
xor U276 (N_276,In_1333,In_18);
nor U277 (N_277,In_1048,In_385);
or U278 (N_278,In_1563,In_565);
and U279 (N_279,In_1440,In_1230);
nor U280 (N_280,In_1032,In_1228);
nand U281 (N_281,In_983,In_351);
and U282 (N_282,In_1006,In_556);
nor U283 (N_283,In_1494,In_919);
or U284 (N_284,In_1842,In_1418);
nand U285 (N_285,In_1968,In_1681);
and U286 (N_286,In_1240,In_1770);
nor U287 (N_287,In_86,In_697);
or U288 (N_288,In_1888,In_1227);
nand U289 (N_289,In_212,In_53);
and U290 (N_290,In_285,In_416);
nand U291 (N_291,In_448,In_220);
nor U292 (N_292,In_1917,In_1160);
nand U293 (N_293,In_534,In_1838);
or U294 (N_294,In_1024,In_1162);
and U295 (N_295,In_1967,In_1818);
and U296 (N_296,In_671,In_374);
nand U297 (N_297,In_1151,In_1324);
xor U298 (N_298,In_1905,In_1361);
and U299 (N_299,In_648,In_367);
or U300 (N_300,In_378,In_1588);
nor U301 (N_301,In_1463,In_186);
nor U302 (N_302,In_1936,In_959);
nor U303 (N_303,In_1875,In_1146);
nor U304 (N_304,In_1177,In_213);
and U305 (N_305,In_730,In_1390);
and U306 (N_306,In_499,In_1617);
nor U307 (N_307,In_672,In_468);
and U308 (N_308,In_1873,In_1037);
nor U309 (N_309,In_1342,In_1419);
and U310 (N_310,In_381,In_1281);
or U311 (N_311,In_1274,In_1043);
or U312 (N_312,In_1183,In_1738);
xnor U313 (N_313,In_596,In_101);
nor U314 (N_314,In_836,In_1503);
nand U315 (N_315,In_445,In_1318);
nor U316 (N_316,In_1305,In_1934);
nand U317 (N_317,In_591,In_1155);
nor U318 (N_318,In_949,In_137);
nor U319 (N_319,In_433,In_282);
nor U320 (N_320,In_91,In_1543);
or U321 (N_321,In_1689,In_1822);
and U322 (N_322,In_517,In_1570);
nor U323 (N_323,In_1259,In_1654);
nand U324 (N_324,In_1472,In_461);
or U325 (N_325,In_1014,In_365);
and U326 (N_326,In_1422,In_864);
nand U327 (N_327,In_1425,In_1444);
and U328 (N_328,In_702,In_1692);
and U329 (N_329,In_1973,In_1607);
nand U330 (N_330,In_977,In_11);
and U331 (N_331,In_942,In_1459);
or U332 (N_332,In_1389,In_886);
and U333 (N_333,In_196,In_891);
or U334 (N_334,In_721,In_616);
nor U335 (N_335,In_843,In_1965);
nand U336 (N_336,In_1528,In_162);
or U337 (N_337,In_370,In_1203);
nand U338 (N_338,In_1727,In_1041);
nand U339 (N_339,In_139,In_1957);
nor U340 (N_340,In_756,In_819);
or U341 (N_341,In_65,In_1760);
nand U342 (N_342,In_1056,In_290);
and U343 (N_343,In_1476,In_946);
nor U344 (N_344,In_266,In_1942);
nand U345 (N_345,In_344,In_1717);
nand U346 (N_346,In_388,In_1539);
nor U347 (N_347,In_510,In_1232);
or U348 (N_348,In_1652,In_1402);
nor U349 (N_349,In_1698,In_1966);
nand U350 (N_350,In_1290,In_1271);
nor U351 (N_351,In_1901,In_1513);
or U352 (N_352,In_823,In_970);
and U353 (N_353,In_150,In_1769);
nand U354 (N_354,In_1542,In_1340);
nor U355 (N_355,In_157,In_542);
and U356 (N_356,In_701,In_1287);
or U357 (N_357,In_774,In_1720);
or U358 (N_358,In_1534,In_1008);
or U359 (N_359,In_1156,In_1387);
nor U360 (N_360,In_572,In_583);
nand U361 (N_361,In_752,In_680);
or U362 (N_362,In_938,In_1300);
nor U363 (N_363,In_1353,In_373);
and U364 (N_364,In_1999,In_346);
or U365 (N_365,In_1112,In_559);
and U366 (N_366,In_296,In_44);
or U367 (N_367,In_1778,In_980);
or U368 (N_368,In_813,In_789);
nand U369 (N_369,In_458,In_1547);
and U370 (N_370,In_779,In_1386);
and U371 (N_371,In_364,In_1110);
nand U372 (N_372,In_1188,In_940);
and U373 (N_373,In_117,In_1763);
and U374 (N_374,In_129,In_1436);
or U375 (N_375,In_1964,In_1867);
and U376 (N_376,In_1360,In_976);
or U377 (N_377,In_417,In_799);
nor U378 (N_378,In_1846,In_155);
nand U379 (N_379,In_809,In_805);
and U380 (N_380,In_1377,In_1932);
or U381 (N_381,In_764,In_1252);
or U382 (N_382,In_446,In_175);
or U383 (N_383,In_1735,In_430);
or U384 (N_384,In_812,In_1328);
nand U385 (N_385,In_1821,In_1108);
and U386 (N_386,In_1586,In_1452);
nor U387 (N_387,In_42,In_692);
and U388 (N_388,In_1711,In_79);
nor U389 (N_389,In_1128,In_1601);
nand U390 (N_390,In_975,In_883);
nor U391 (N_391,In_151,In_1029);
or U392 (N_392,In_1116,In_1127);
nand U393 (N_393,In_470,In_564);
and U394 (N_394,In_1348,In_926);
nor U395 (N_395,In_1860,In_1703);
or U396 (N_396,In_229,In_1512);
nand U397 (N_397,In_887,In_1865);
and U398 (N_398,In_384,In_1545);
nor U399 (N_399,In_1167,In_1107);
nor U400 (N_400,In_682,In_908);
nor U401 (N_401,In_1265,In_291);
nand U402 (N_402,In_254,In_954);
nor U403 (N_403,In_1913,In_1480);
or U404 (N_404,In_828,In_853);
nor U405 (N_405,In_1015,In_903);
and U406 (N_406,In_1729,In_1207);
or U407 (N_407,In_863,In_1549);
xnor U408 (N_408,In_1848,In_599);
and U409 (N_409,In_1068,In_331);
nor U410 (N_410,In_361,In_1253);
nand U411 (N_411,In_1622,In_473);
and U412 (N_412,In_664,In_1217);
nand U413 (N_413,In_934,In_1992);
xor U414 (N_414,In_223,In_1501);
nand U415 (N_415,In_1863,In_1245);
or U416 (N_416,In_871,In_738);
and U417 (N_417,In_395,In_1914);
xor U418 (N_418,In_1201,In_1113);
or U419 (N_419,In_1457,In_38);
or U420 (N_420,In_339,In_1065);
nor U421 (N_421,In_1437,In_74);
nand U422 (N_422,In_376,In_1687);
and U423 (N_423,In_531,In_103);
or U424 (N_424,In_1104,In_1955);
or U425 (N_425,In_842,In_867);
and U426 (N_426,In_1019,In_1332);
nand U427 (N_427,In_575,In_337);
and U428 (N_428,In_1504,In_1604);
nor U429 (N_429,In_1879,In_551);
nor U430 (N_430,In_1310,In_584);
or U431 (N_431,In_753,In_288);
and U432 (N_432,In_250,In_1979);
and U433 (N_433,In_1388,In_964);
and U434 (N_434,In_1912,In_1704);
nand U435 (N_435,In_736,In_263);
and U436 (N_436,In_132,In_1161);
or U437 (N_437,In_544,In_1246);
or U438 (N_438,In_1456,In_1969);
and U439 (N_439,In_1135,In_817);
and U440 (N_440,In_1750,In_1066);
and U441 (N_441,In_1923,In_1070);
nand U442 (N_442,In_307,In_1088);
nand U443 (N_443,In_1101,In_475);
and U444 (N_444,In_1576,In_927);
nor U445 (N_445,In_1947,In_898);
and U446 (N_446,In_148,In_232);
nand U447 (N_447,In_879,In_1139);
nor U448 (N_448,In_199,In_1074);
and U449 (N_449,In_698,In_1121);
nand U450 (N_450,In_1978,In_411);
or U451 (N_451,In_1175,In_1001);
or U452 (N_452,In_850,In_428);
nor U453 (N_453,In_1798,In_1130);
nand U454 (N_454,In_52,In_1981);
nor U455 (N_455,In_611,In_629);
and U456 (N_456,In_1653,In_284);
and U457 (N_457,In_1164,In_1983);
nand U458 (N_458,In_1736,In_538);
or U459 (N_459,In_1125,In_912);
and U460 (N_460,In_1034,In_1646);
or U461 (N_461,In_1850,In_414);
nor U462 (N_462,In_167,In_265);
and U463 (N_463,In_420,In_1921);
nand U464 (N_464,In_1359,In_562);
nand U465 (N_465,In_77,In_1158);
and U466 (N_466,In_1538,In_225);
and U467 (N_467,In_1012,In_492);
and U468 (N_468,In_1394,In_553);
nor U469 (N_469,In_1722,In_1784);
and U470 (N_470,In_996,In_665);
or U471 (N_471,In_90,In_1841);
and U472 (N_472,In_1383,In_1002);
nand U473 (N_473,In_1767,In_1943);
nand U474 (N_474,In_205,In_489);
or U475 (N_475,In_525,In_1609);
or U476 (N_476,In_1408,In_783);
and U477 (N_477,In_1544,In_1379);
or U478 (N_478,In_1911,In_586);
and U479 (N_479,In_313,In_495);
nor U480 (N_480,In_1963,In_1728);
nand U481 (N_481,In_280,In_1367);
or U482 (N_482,In_685,In_68);
and U483 (N_483,In_1527,In_1997);
nor U484 (N_484,In_142,In_237);
and U485 (N_485,In_1907,In_85);
and U486 (N_486,In_1635,In_158);
or U487 (N_487,In_1264,In_1524);
nand U488 (N_488,In_506,In_1442);
or U489 (N_489,In_1550,In_670);
nor U490 (N_490,In_434,In_453);
xnor U491 (N_491,In_435,In_432);
or U492 (N_492,In_1847,In_99);
nor U493 (N_493,In_627,In_1810);
nand U494 (N_494,In_1323,In_703);
and U495 (N_495,In_537,In_1017);
or U496 (N_496,In_1060,In_1777);
or U497 (N_497,In_494,In_566);
or U498 (N_498,In_603,In_1381);
or U499 (N_499,In_979,In_604);
nand U500 (N_500,In_929,In_1200);
or U501 (N_501,In_1482,In_1210);
or U502 (N_502,In_1774,In_1330);
nand U503 (N_503,In_501,In_389);
xor U504 (N_504,In_576,In_423);
nor U505 (N_505,In_875,In_1345);
nor U506 (N_506,In_1366,In_1691);
and U507 (N_507,In_451,In_1522);
nand U508 (N_508,In_952,In_1087);
nand U509 (N_509,In_1234,In_848);
and U510 (N_510,In_696,In_233);
or U511 (N_511,In_407,In_1890);
and U512 (N_512,In_873,In_256);
nand U513 (N_513,In_293,In_1758);
nand U514 (N_514,In_1018,In_571);
or U515 (N_515,In_725,In_967);
or U516 (N_516,In_274,In_1506);
xnor U517 (N_517,In_1439,In_1510);
or U518 (N_518,In_1372,In_486);
or U519 (N_519,In_1674,In_771);
nor U520 (N_520,In_300,In_1642);
or U521 (N_521,In_1743,In_1325);
nand U522 (N_522,In_854,In_1591);
and U523 (N_523,In_1661,In_597);
or U524 (N_524,In_1291,In_1294);
nand U525 (N_525,In_500,In_309);
nand U526 (N_526,In_656,In_1114);
nand U527 (N_527,In_1357,In_1536);
or U528 (N_528,In_208,In_856);
or U529 (N_529,In_1181,In_406);
and U530 (N_530,In_482,In_621);
and U531 (N_531,In_1971,In_1794);
nand U532 (N_532,In_1579,In_1613);
nand U533 (N_533,In_1643,In_1312);
and U534 (N_534,In_1254,In_1214);
and U535 (N_535,In_113,In_1994);
nor U536 (N_536,In_47,In_904);
nor U537 (N_537,In_1927,In_1830);
or U538 (N_538,In_574,In_104);
nor U539 (N_539,In_1629,In_1889);
nand U540 (N_540,In_1455,In_840);
or U541 (N_541,In_1080,In_1733);
or U542 (N_542,In_1242,In_240);
nor U543 (N_543,In_1453,In_396);
or U544 (N_544,In_1786,In_1693);
nand U545 (N_545,In_1421,In_319);
nor U546 (N_546,In_298,In_62);
nor U547 (N_547,In_694,In_1625);
and U548 (N_548,In_1883,In_1828);
or U549 (N_549,In_1100,In_358);
and U550 (N_550,In_1209,In_1761);
nand U551 (N_551,In_1451,In_769);
or U552 (N_552,In_1224,In_957);
nand U553 (N_553,In_427,In_1663);
nor U554 (N_554,In_855,In_1071);
and U555 (N_555,In_608,In_207);
nor U556 (N_556,In_1713,In_198);
nand U557 (N_557,In_1924,In_1671);
and U558 (N_558,In_1020,In_1475);
nor U559 (N_559,In_1222,In_844);
or U560 (N_560,In_247,In_1937);
nand U561 (N_561,In_1174,In_876);
nand U562 (N_562,In_773,In_1196);
and U563 (N_563,In_140,In_1953);
nand U564 (N_564,In_1364,In_1393);
or U565 (N_565,In_899,In_777);
nor U566 (N_566,In_1411,In_917);
nor U567 (N_567,In_1980,In_279);
nor U568 (N_568,In_1583,In_1471);
nand U569 (N_569,In_607,In_1835);
and U570 (N_570,In_1556,In_206);
nor U571 (N_571,In_1446,In_40);
xor U572 (N_572,In_639,In_1626);
and U573 (N_573,In_56,In_1028);
nor U574 (N_574,In_8,In_1584);
nand U575 (N_575,In_814,In_355);
nand U576 (N_576,In_1035,In_1433);
or U577 (N_577,In_1952,In_724);
nor U578 (N_578,In_253,In_1376);
nand U579 (N_579,In_1996,In_1374);
nand U580 (N_580,In_1131,In_708);
and U581 (N_581,In_297,In_415);
or U582 (N_582,In_826,In_1062);
and U583 (N_583,In_37,In_1897);
nand U584 (N_584,In_602,In_1598);
nand U585 (N_585,In_1106,In_734);
nor U586 (N_586,In_914,In_1603);
nand U587 (N_587,In_457,In_716);
nor U588 (N_588,In_1811,In_1123);
nand U589 (N_589,In_1049,In_275);
and U590 (N_590,In_1918,In_1061);
nand U591 (N_591,In_21,In_985);
nand U592 (N_592,In_982,In_1593);
and U593 (N_593,In_1780,In_154);
nor U594 (N_594,In_947,In_762);
or U595 (N_595,In_488,In_965);
nand U596 (N_596,In_770,In_71);
nor U597 (N_597,In_398,In_59);
and U598 (N_598,In_930,In_1191);
or U599 (N_599,In_483,In_413);
nand U600 (N_600,In_20,In_1339);
and U601 (N_601,In_1218,In_442);
nor U602 (N_602,In_1805,In_426);
and U603 (N_603,In_1270,In_1710);
and U604 (N_604,In_97,In_1874);
nand U605 (N_605,In_765,In_354);
and U606 (N_606,In_1428,In_1050);
and U607 (N_607,In_422,In_1179);
nor U608 (N_608,In_1740,In_1085);
or U609 (N_609,In_431,In_1000);
nor U610 (N_610,In_1523,In_219);
and U611 (N_611,In_1186,In_1723);
nor U612 (N_612,In_349,In_1165);
nand U613 (N_613,In_441,In_1575);
nor U614 (N_614,In_184,In_1343);
or U615 (N_615,In_156,In_202);
and U616 (N_616,In_377,In_1565);
nor U617 (N_617,In_1126,In_1115);
nor U618 (N_618,In_824,In_1079);
nand U619 (N_619,In_1714,In_668);
nand U620 (N_620,In_1843,In_1925);
xnor U621 (N_621,In_176,In_1574);
or U622 (N_622,In_1949,In_1958);
nor U623 (N_623,In_928,In_944);
and U624 (N_624,In_502,In_1871);
nand U625 (N_625,In_533,In_387);
nand U626 (N_626,In_1416,In_168);
and U627 (N_627,In_1337,In_684);
or U628 (N_628,In_1309,In_1465);
or U629 (N_629,In_711,In_1159);
or U630 (N_630,In_1238,In_193);
nor U631 (N_631,In_102,In_144);
nand U632 (N_632,In_128,In_936);
or U633 (N_633,In_1344,In_981);
nand U634 (N_634,In_1257,In_1078);
nand U635 (N_635,In_464,In_935);
or U636 (N_636,In_1315,In_1326);
and U637 (N_637,In_579,In_1063);
and U638 (N_638,In_64,In_897);
and U639 (N_639,In_541,In_1351);
nand U640 (N_640,In_1819,In_1809);
or U641 (N_641,In_1117,In_226);
and U642 (N_642,In_1644,In_1884);
and U643 (N_643,In_1526,In_1572);
nor U644 (N_644,In_314,In_1286);
nand U645 (N_645,In_1199,In_1403);
nor U646 (N_646,In_968,In_570);
or U647 (N_647,In_1086,In_340);
or U648 (N_648,In_1235,In_960);
nor U649 (N_649,In_1244,In_802);
nor U650 (N_650,In_1277,In_1023);
or U651 (N_651,In_1320,In_1170);
nor U652 (N_652,In_1566,In_846);
nor U653 (N_653,In_1615,In_1605);
nor U654 (N_654,In_948,In_323);
or U655 (N_655,In_1016,In_438);
or U656 (N_656,In_622,In_1783);
nand U657 (N_657,In_1295,In_181);
nand U658 (N_658,In_858,In_1946);
nor U659 (N_659,In_530,In_1414);
nand U660 (N_660,In_166,In_606);
nor U661 (N_661,In_955,In_401);
and U662 (N_662,In_1336,In_1898);
nand U663 (N_663,In_1749,In_504);
xor U664 (N_664,In_1686,In_700);
and U665 (N_665,In_1531,In_1089);
nor U666 (N_666,In_707,In_234);
or U667 (N_667,In_1616,In_1546);
or U668 (N_668,In_1939,In_402);
or U669 (N_669,In_513,In_1432);
and U670 (N_670,In_1435,In_1753);
or U671 (N_671,In_1892,In_1690);
and U672 (N_672,In_907,In_834);
nor U673 (N_673,In_880,In_1073);
and U674 (N_674,In_647,In_303);
or U675 (N_675,In_515,In_217);
or U676 (N_676,In_1498,In_1189);
nor U677 (N_677,In_1298,In_1288);
nand U678 (N_678,In_1801,In_1594);
nor U679 (N_679,In_1426,In_1695);
nand U680 (N_680,In_1350,In_1382);
nand U681 (N_681,In_1038,In_1826);
and U682 (N_682,In_1988,In_1659);
nor U683 (N_683,In_105,In_315);
and U684 (N_684,In_869,In_615);
nor U685 (N_685,In_1166,In_1998);
nor U686 (N_686,In_1667,In_1606);
or U687 (N_687,In_1954,In_822);
and U688 (N_688,In_1304,In_1857);
nand U689 (N_689,In_161,In_787);
and U690 (N_690,In_106,In_554);
nor U691 (N_691,In_1094,In_1491);
or U692 (N_692,In_941,In_34);
nor U693 (N_693,In_1694,In_1137);
nor U694 (N_694,In_1991,In_837);
or U695 (N_695,In_1844,In_797);
nor U696 (N_696,In_1899,In_436);
nand U697 (N_697,In_1734,In_742);
and U698 (N_698,In_1627,In_687);
nand U699 (N_699,In_283,In_1972);
and U700 (N_700,In_1521,In_1910);
and U701 (N_701,In_1184,In_1509);
nor U702 (N_702,In_1699,In_1313);
nor U703 (N_703,In_1278,In_1719);
or U704 (N_704,In_1585,In_107);
or U705 (N_705,In_1802,In_218);
nor U706 (N_706,In_278,In_1);
and U707 (N_707,In_1533,In_1540);
and U708 (N_708,In_462,In_1297);
nand U709 (N_709,In_1950,In_268);
or U710 (N_710,In_1064,In_1638);
or U711 (N_711,In_1880,In_16);
nand U712 (N_712,In_1059,In_922);
or U713 (N_713,In_874,In_832);
or U714 (N_714,In_663,In_1634);
or U715 (N_715,In_1869,In_1595);
nor U716 (N_716,In_652,In_1375);
or U717 (N_717,In_1511,In_1111);
nor U718 (N_718,In_392,In_624);
nor U719 (N_719,In_332,In_1508);
and U720 (N_720,In_1684,In_1276);
or U721 (N_721,In_1651,In_187);
or U722 (N_722,In_1025,In_1047);
and U723 (N_723,In_130,In_550);
xor U724 (N_724,In_258,In_1938);
and U725 (N_725,In_121,In_1216);
and U726 (N_726,In_720,In_1321);
or U727 (N_727,In_1977,In_1208);
or U728 (N_728,In_1083,In_335);
nand U729 (N_729,In_1054,In_460);
nand U730 (N_730,In_956,In_348);
and U731 (N_731,In_28,In_1682);
and U732 (N_732,In_119,In_1284);
and U733 (N_733,In_469,In_109);
or U734 (N_734,In_1306,In_536);
nor U735 (N_735,In_1976,In_1507);
and U736 (N_736,In_915,In_404);
xnor U737 (N_737,In_1202,In_511);
nand U738 (N_738,In_1142,In_334);
or U739 (N_739,In_609,In_1406);
or U740 (N_740,In_1102,In_527);
nor U741 (N_741,In_1895,In_306);
nand U742 (N_742,In_259,In_1672);
nand U743 (N_743,In_1413,In_149);
nor U744 (N_744,In_1027,In_1670);
and U745 (N_745,In_1985,In_635);
nor U746 (N_746,In_216,In_1922);
nand U747 (N_747,In_1488,In_312);
or U748 (N_748,In_943,In_1903);
and U749 (N_749,In_601,In_674);
nor U750 (N_750,In_1578,In_1648);
or U751 (N_751,In_835,In_1220);
and U752 (N_752,In_507,In_1401);
nand U753 (N_753,In_1827,In_1929);
or U754 (N_754,In_1612,In_1398);
or U755 (N_755,In_78,In_1799);
and U756 (N_756,In_455,In_705);
xor U757 (N_757,In_1785,In_1962);
nor U758 (N_758,In_862,In_1352);
nor U759 (N_759,In_1075,In_750);
nand U760 (N_760,In_1098,In_1564);
and U761 (N_761,In_397,In_295);
or U762 (N_762,In_1173,In_1077);
nand U763 (N_763,In_211,In_1356);
nor U764 (N_764,In_1807,In_1499);
nand U765 (N_765,In_1529,In_839);
or U766 (N_766,In_1132,In_487);
nand U767 (N_767,In_516,In_580);
and U768 (N_768,In_1396,In_1308);
nand U769 (N_769,In_1256,In_214);
and U770 (N_770,In_793,In_625);
and U771 (N_771,In_1502,In_691);
or U772 (N_772,In_1053,In_1933);
or U773 (N_773,In_1730,In_1557);
and U774 (N_774,In_88,In_1716);
or U775 (N_775,In_311,In_699);
and U776 (N_776,In_408,In_108);
nand U777 (N_777,In_1163,In_984);
nand U778 (N_778,In_1677,In_1577);
nand U779 (N_779,In_235,In_493);
nand U780 (N_780,In_92,In_277);
and U781 (N_781,In_818,In_262);
nand U782 (N_782,In_472,In_363);
and U783 (N_783,In_10,In_1516);
and U784 (N_784,In_1647,In_1862);
nor U785 (N_785,In_191,In_1493);
nor U786 (N_786,In_528,In_1630);
or U787 (N_787,In_1285,In_543);
nor U788 (N_788,In_1791,In_1872);
and U789 (N_789,In_1845,In_116);
nor U790 (N_790,In_587,In_645);
or U791 (N_791,In_969,In_785);
nand U792 (N_792,In_815,In_1307);
and U793 (N_793,In_632,In_1916);
or U794 (N_794,In_1833,In_1649);
nand U795 (N_795,In_1182,In_906);
nand U796 (N_796,In_1640,In_1354);
nor U797 (N_797,In_1211,In_1628);
nand U798 (N_798,In_96,In_1832);
or U799 (N_799,In_1225,In_1815);
nor U800 (N_800,In_227,In_642);
or U801 (N_801,In_1517,In_22);
nor U802 (N_802,In_369,In_1447);
or U803 (N_803,In_350,In_1945);
and U804 (N_804,In_727,In_326);
or U805 (N_805,In_1405,In_893);
and U806 (N_806,In_1468,In_1399);
nor U807 (N_807,In_1096,In_1747);
nand U808 (N_808,In_1571,In_1775);
nor U809 (N_809,In_228,In_754);
nor U810 (N_810,In_681,In_454);
nand U811 (N_811,In_801,In_1093);
or U812 (N_812,In_1103,In_1229);
and U813 (N_813,In_1226,In_80);
or U814 (N_814,In_1144,In_95);
nor U815 (N_815,In_796,In_410);
or U816 (N_816,In_5,In_1891);
and U817 (N_817,In_1400,In_1655);
or U818 (N_818,In_1267,In_821);
or U819 (N_819,In_1233,In_170);
and U820 (N_820,In_1851,In_1460);
or U821 (N_821,In_1003,In_717);
nor U822 (N_822,In_512,In_347);
and U823 (N_823,In_1004,In_1707);
nand U824 (N_824,In_329,In_1859);
xnor U825 (N_825,In_731,In_810);
and U826 (N_826,In_1057,In_1632);
and U827 (N_827,In_1097,In_1618);
nand U828 (N_828,In_1631,In_1458);
nand U829 (N_829,In_1731,In_693);
nand U830 (N_830,In_1995,In_466);
nand U831 (N_831,In_1590,In_1662);
nor U832 (N_832,In_236,In_1427);
nor U833 (N_833,In_1781,In_1641);
or U834 (N_834,In_480,In_270);
and U835 (N_835,In_560,In_638);
nand U836 (N_836,In_1806,In_1614);
nand U837 (N_837,In_620,In_63);
nand U838 (N_838,In_761,In_1477);
nand U839 (N_839,In_567,In_726);
nor U840 (N_840,In_75,In_147);
and U841 (N_841,In_923,In_1423);
or U842 (N_842,In_273,In_333);
and U843 (N_843,In_440,In_1680);
or U844 (N_844,In_1204,In_518);
and U845 (N_845,In_1373,In_29);
nand U846 (N_846,In_966,In_522);
and U847 (N_847,In_1567,In_660);
nand U848 (N_848,In_896,In_866);
nor U849 (N_849,In_136,In_998);
or U850 (N_850,In_1010,In_24);
and U851 (N_851,In_1247,In_744);
and U852 (N_852,In_859,In_443);
nand U853 (N_853,In_808,In_1150);
nand U854 (N_854,In_308,In_1941);
and U855 (N_855,In_1789,In_784);
nor U856 (N_856,In_1148,In_1322);
nand U857 (N_857,In_1407,In_973);
nand U858 (N_858,In_1555,In_1198);
and U859 (N_859,In_913,In_1341);
nor U860 (N_860,In_933,In_1823);
and U861 (N_861,In_1762,In_689);
and U862 (N_862,In_618,In_901);
and U863 (N_863,In_1515,In_1479);
nand U864 (N_864,In_920,In_7);
or U865 (N_865,In_881,In_1840);
nor U866 (N_866,In_690,In_1152);
nor U867 (N_867,In_1241,In_1771);
and U868 (N_868,In_215,In_825);
or U869 (N_869,In_1072,In_1683);
nor U870 (N_870,In_790,In_1919);
and U871 (N_871,In_644,In_243);
nand U872 (N_872,In_1454,In_200);
or U873 (N_873,In_124,In_735);
nor U874 (N_874,In_1464,In_330);
and U875 (N_875,In_1490,In_163);
nand U876 (N_876,In_1742,In_1206);
nor U877 (N_877,In_974,In_1261);
nor U878 (N_878,In_1221,In_484);
nor U879 (N_879,In_317,In_722);
or U880 (N_880,In_424,In_612);
and U881 (N_881,In_1989,In_737);
or U882 (N_882,In_1558,In_1319);
nor U883 (N_883,In_1530,In_1745);
and U884 (N_884,In_686,In_1560);
and U885 (N_885,In_1268,In_1800);
and U886 (N_886,In_1970,In_1363);
nand U887 (N_887,In_1896,In_362);
nand U888 (N_888,In_1856,In_36);
xor U889 (N_889,In_546,In_1011);
or U890 (N_890,In_164,In_338);
nor U891 (N_891,In_704,In_782);
nor U892 (N_892,In_359,In_294);
and U893 (N_893,In_1882,In_1852);
and U894 (N_894,In_23,In_1099);
nor U895 (N_895,In_1514,In_573);
and U896 (N_896,In_1596,In_1495);
and U897 (N_897,In_990,In_1021);
nand U898 (N_898,In_360,In_1825);
nand U899 (N_899,In_1746,In_1829);
nand U900 (N_900,In_1797,In_1327);
nand U901 (N_901,In_582,In_1051);
or U902 (N_902,In_324,In_444);
xnor U903 (N_903,In_757,In_1537);
nand U904 (N_904,In_1052,In_321);
nor U905 (N_905,In_547,In_1236);
and U906 (N_906,In_577,In_1296);
nor U907 (N_907,In_1154,In_872);
nand U908 (N_908,In_706,In_185);
and U909 (N_909,In_1302,In_1702);
or U910 (N_910,In_1223,In_1193);
and U911 (N_911,In_1568,In_171);
nor U912 (N_912,In_902,In_57);
nor U913 (N_913,In_33,In_804);
and U914 (N_914,In_1705,In_1095);
or U915 (N_915,In_1046,In_1673);
xor U916 (N_916,In_1599,In_1532);
or U917 (N_917,In_1935,In_1752);
and U918 (N_918,In_520,In_1836);
nand U919 (N_919,In_479,In_1409);
or U920 (N_920,In_169,In_50);
nand U921 (N_921,In_1610,In_894);
nand U922 (N_922,In_1679,In_1909);
nor U923 (N_923,In_1541,In_69);
nand U924 (N_924,In_1371,In_1497);
nand U925 (N_925,In_1993,In_588);
or U926 (N_926,In_257,In_1554);
and U927 (N_927,In_1741,In_1868);
and U928 (N_928,In_561,In_244);
and U929 (N_929,In_352,In_1553);
and U930 (N_930,In_497,In_1885);
nor U931 (N_931,In_264,In_1141);
nand U932 (N_932,In_857,In_115);
and U933 (N_933,In_1045,In_1134);
and U934 (N_934,In_558,In_1030);
and U935 (N_935,In_1759,In_733);
or U936 (N_936,In_1299,In_1518);
or U937 (N_937,In_1866,In_76);
nor U938 (N_938,In_739,In_251);
nor U939 (N_939,In_195,In_203);
nor U940 (N_940,In_1559,In_678);
or U941 (N_941,In_1990,In_1787);
nor U942 (N_942,In_1685,In_849);
or U943 (N_943,In_1473,In_281);
nor U944 (N_944,In_6,In_1292);
nand U945 (N_945,In_1275,In_481);
and U946 (N_946,In_1573,In_626);
and U947 (N_947,In_1877,In_1940);
nand U948 (N_948,In_669,In_1982);
nand U949 (N_949,In_242,In_613);
or U950 (N_950,In_713,In_1036);
and U951 (N_951,In_84,In_31);
nand U952 (N_952,In_617,In_643);
nand U953 (N_953,In_945,In_188);
nor U954 (N_954,In_1525,In_1431);
and U955 (N_955,In_1272,In_1792);
or U956 (N_956,In_328,In_755);
or U957 (N_957,In_1766,In_390);
or U958 (N_958,In_1176,In_1824);
nor U959 (N_959,In_498,In_937);
and U960 (N_960,In_1757,In_252);
nand U961 (N_961,In_807,In_1349);
or U962 (N_962,In_289,In_1410);
nor U963 (N_963,In_676,In_1365);
and U964 (N_964,In_1329,In_83);
nand U965 (N_965,In_380,In_1109);
nand U966 (N_966,In_925,In_932);
or U967 (N_967,In_1120,In_1796);
and U968 (N_968,In_1930,In_1213);
nand U969 (N_969,In_316,In_201);
nand U970 (N_970,In_1870,In_100);
nand U971 (N_971,In_174,In_833);
or U972 (N_972,In_1960,In_806);
and U973 (N_973,In_1335,In_1469);
nand U974 (N_974,In_54,In_1592);
and U975 (N_975,In_1280,In_13);
nand U976 (N_976,In_1886,In_1362);
or U977 (N_977,In_921,In_491);
nor U978 (N_978,In_767,In_1255);
or U979 (N_979,In_1461,In_555);
nor U980 (N_980,In_204,In_503);
nor U981 (N_981,In_1709,In_1754);
and U982 (N_982,In_372,In_962);
and U983 (N_983,In_267,In_30);
nor U984 (N_984,In_1273,In_32);
and U985 (N_985,In_1467,In_593);
nor U986 (N_986,In_1650,In_1260);
and U987 (N_987,In_1666,In_127);
or U988 (N_988,In_1171,In_73);
nand U989 (N_989,In_1621,In_718);
nor U990 (N_990,In_1987,In_272);
nor U991 (N_991,In_1804,In_1180);
nor U992 (N_992,In_751,In_1623);
or U993 (N_993,In_1289,In_994);
or U994 (N_994,In_183,In_993);
nor U995 (N_995,In_695,In_1385);
nand U996 (N_996,In_341,In_1022);
nand U997 (N_997,In_467,In_931);
or U998 (N_998,In_51,In_650);
nand U999 (N_999,In_1136,In_1900);
or U1000 (N_1000,In_861,In_1935);
and U1001 (N_1001,In_1787,In_1601);
or U1002 (N_1002,In_52,In_489);
nand U1003 (N_1003,In_714,In_1265);
nand U1004 (N_1004,In_1161,In_1716);
or U1005 (N_1005,In_1404,In_1148);
nor U1006 (N_1006,In_625,In_456);
or U1007 (N_1007,In_1442,In_1009);
nand U1008 (N_1008,In_161,In_1325);
nand U1009 (N_1009,In_19,In_982);
and U1010 (N_1010,In_1007,In_526);
or U1011 (N_1011,In_69,In_1533);
and U1012 (N_1012,In_1775,In_32);
nor U1013 (N_1013,In_1537,In_1440);
or U1014 (N_1014,In_1696,In_1561);
and U1015 (N_1015,In_456,In_1425);
nor U1016 (N_1016,In_1510,In_553);
nor U1017 (N_1017,In_1128,In_17);
or U1018 (N_1018,In_1314,In_694);
or U1019 (N_1019,In_711,In_1813);
nand U1020 (N_1020,In_625,In_833);
and U1021 (N_1021,In_1108,In_584);
and U1022 (N_1022,In_829,In_554);
nor U1023 (N_1023,In_1320,In_190);
and U1024 (N_1024,In_1412,In_1603);
and U1025 (N_1025,In_1388,In_1686);
nand U1026 (N_1026,In_69,In_630);
nor U1027 (N_1027,In_1273,In_1557);
nor U1028 (N_1028,In_843,In_1981);
nand U1029 (N_1029,In_1942,In_649);
and U1030 (N_1030,In_645,In_357);
or U1031 (N_1031,In_1453,In_1934);
and U1032 (N_1032,In_1541,In_1250);
or U1033 (N_1033,In_1254,In_1912);
or U1034 (N_1034,In_1341,In_578);
or U1035 (N_1035,In_296,In_204);
nand U1036 (N_1036,In_1390,In_1447);
or U1037 (N_1037,In_1572,In_508);
or U1038 (N_1038,In_735,In_1666);
and U1039 (N_1039,In_280,In_1071);
nand U1040 (N_1040,In_737,In_22);
nor U1041 (N_1041,In_225,In_610);
and U1042 (N_1042,In_932,In_799);
or U1043 (N_1043,In_1577,In_412);
and U1044 (N_1044,In_1045,In_979);
or U1045 (N_1045,In_1910,In_1508);
and U1046 (N_1046,In_1828,In_824);
and U1047 (N_1047,In_1296,In_424);
and U1048 (N_1048,In_1379,In_98);
nor U1049 (N_1049,In_371,In_368);
or U1050 (N_1050,In_1467,In_187);
nand U1051 (N_1051,In_697,In_1055);
xnor U1052 (N_1052,In_892,In_1550);
nor U1053 (N_1053,In_1633,In_111);
nand U1054 (N_1054,In_1104,In_849);
nor U1055 (N_1055,In_930,In_695);
or U1056 (N_1056,In_1794,In_1657);
nand U1057 (N_1057,In_1924,In_464);
and U1058 (N_1058,In_400,In_1899);
and U1059 (N_1059,In_547,In_607);
nor U1060 (N_1060,In_617,In_1529);
nand U1061 (N_1061,In_1009,In_346);
nand U1062 (N_1062,In_1919,In_1337);
nor U1063 (N_1063,In_1168,In_1427);
nor U1064 (N_1064,In_1575,In_930);
and U1065 (N_1065,In_697,In_1688);
and U1066 (N_1066,In_1047,In_1998);
nand U1067 (N_1067,In_1313,In_1196);
nand U1068 (N_1068,In_1150,In_1827);
and U1069 (N_1069,In_878,In_1016);
or U1070 (N_1070,In_1276,In_1556);
nor U1071 (N_1071,In_1776,In_1591);
nor U1072 (N_1072,In_1166,In_1205);
nor U1073 (N_1073,In_962,In_907);
nor U1074 (N_1074,In_437,In_552);
and U1075 (N_1075,In_240,In_39);
and U1076 (N_1076,In_454,In_1877);
or U1077 (N_1077,In_237,In_1580);
nor U1078 (N_1078,In_1132,In_1514);
nand U1079 (N_1079,In_1525,In_79);
and U1080 (N_1080,In_1122,In_1428);
nand U1081 (N_1081,In_950,In_549);
nor U1082 (N_1082,In_1135,In_1698);
nand U1083 (N_1083,In_1163,In_905);
or U1084 (N_1084,In_906,In_283);
nand U1085 (N_1085,In_1388,In_1158);
nor U1086 (N_1086,In_119,In_1750);
or U1087 (N_1087,In_1427,In_1770);
or U1088 (N_1088,In_235,In_672);
nand U1089 (N_1089,In_1416,In_784);
and U1090 (N_1090,In_870,In_862);
nand U1091 (N_1091,In_453,In_1101);
nand U1092 (N_1092,In_452,In_1008);
or U1093 (N_1093,In_20,In_41);
or U1094 (N_1094,In_1548,In_1340);
or U1095 (N_1095,In_1857,In_576);
or U1096 (N_1096,In_145,In_1307);
nor U1097 (N_1097,In_920,In_730);
or U1098 (N_1098,In_1142,In_169);
or U1099 (N_1099,In_798,In_749);
nor U1100 (N_1100,In_1962,In_194);
nand U1101 (N_1101,In_599,In_596);
nand U1102 (N_1102,In_1793,In_1296);
nand U1103 (N_1103,In_1594,In_1785);
or U1104 (N_1104,In_767,In_951);
or U1105 (N_1105,In_981,In_1327);
and U1106 (N_1106,In_1659,In_448);
xnor U1107 (N_1107,In_1646,In_1178);
and U1108 (N_1108,In_1260,In_117);
or U1109 (N_1109,In_586,In_152);
and U1110 (N_1110,In_1318,In_893);
nand U1111 (N_1111,In_169,In_803);
and U1112 (N_1112,In_837,In_1250);
nand U1113 (N_1113,In_1380,In_85);
or U1114 (N_1114,In_934,In_101);
nor U1115 (N_1115,In_37,In_1782);
nand U1116 (N_1116,In_1501,In_1351);
nor U1117 (N_1117,In_5,In_928);
and U1118 (N_1118,In_1820,In_787);
or U1119 (N_1119,In_604,In_36);
and U1120 (N_1120,In_1885,In_663);
nand U1121 (N_1121,In_1609,In_1423);
nand U1122 (N_1122,In_1910,In_225);
and U1123 (N_1123,In_499,In_166);
nor U1124 (N_1124,In_1549,In_92);
and U1125 (N_1125,In_368,In_795);
nand U1126 (N_1126,In_907,In_1411);
and U1127 (N_1127,In_1218,In_742);
nand U1128 (N_1128,In_552,In_643);
nor U1129 (N_1129,In_558,In_1024);
nor U1130 (N_1130,In_947,In_607);
and U1131 (N_1131,In_816,In_1431);
nand U1132 (N_1132,In_491,In_164);
and U1133 (N_1133,In_831,In_256);
nor U1134 (N_1134,In_1570,In_665);
nor U1135 (N_1135,In_810,In_1827);
nand U1136 (N_1136,In_419,In_1491);
or U1137 (N_1137,In_1998,In_1196);
and U1138 (N_1138,In_1703,In_1505);
nand U1139 (N_1139,In_212,In_1405);
nand U1140 (N_1140,In_135,In_1499);
nand U1141 (N_1141,In_786,In_984);
xor U1142 (N_1142,In_354,In_732);
nand U1143 (N_1143,In_492,In_376);
nor U1144 (N_1144,In_1097,In_510);
nand U1145 (N_1145,In_1845,In_1814);
or U1146 (N_1146,In_862,In_86);
nand U1147 (N_1147,In_459,In_941);
nor U1148 (N_1148,In_551,In_1212);
nand U1149 (N_1149,In_196,In_1519);
and U1150 (N_1150,In_203,In_1601);
nand U1151 (N_1151,In_78,In_810);
nor U1152 (N_1152,In_808,In_643);
or U1153 (N_1153,In_823,In_68);
or U1154 (N_1154,In_1128,In_319);
and U1155 (N_1155,In_435,In_209);
nand U1156 (N_1156,In_1562,In_347);
nor U1157 (N_1157,In_1365,In_276);
or U1158 (N_1158,In_507,In_1651);
nor U1159 (N_1159,In_1944,In_1459);
nor U1160 (N_1160,In_1845,In_1435);
or U1161 (N_1161,In_1991,In_1068);
nor U1162 (N_1162,In_77,In_1712);
nand U1163 (N_1163,In_1354,In_1253);
nand U1164 (N_1164,In_1026,In_260);
nor U1165 (N_1165,In_846,In_1918);
nor U1166 (N_1166,In_286,In_363);
and U1167 (N_1167,In_1212,In_565);
or U1168 (N_1168,In_1625,In_775);
and U1169 (N_1169,In_641,In_1848);
nand U1170 (N_1170,In_574,In_1788);
or U1171 (N_1171,In_1586,In_604);
nor U1172 (N_1172,In_416,In_655);
nor U1173 (N_1173,In_269,In_430);
nand U1174 (N_1174,In_1467,In_1563);
nand U1175 (N_1175,In_566,In_475);
or U1176 (N_1176,In_481,In_550);
or U1177 (N_1177,In_1620,In_1933);
nor U1178 (N_1178,In_1132,In_7);
and U1179 (N_1179,In_385,In_1156);
and U1180 (N_1180,In_617,In_1582);
nor U1181 (N_1181,In_1988,In_657);
or U1182 (N_1182,In_1952,In_604);
nor U1183 (N_1183,In_1630,In_909);
and U1184 (N_1184,In_1723,In_1779);
and U1185 (N_1185,In_906,In_269);
or U1186 (N_1186,In_922,In_909);
nand U1187 (N_1187,In_92,In_760);
and U1188 (N_1188,In_1111,In_26);
nand U1189 (N_1189,In_1094,In_1890);
and U1190 (N_1190,In_212,In_1187);
and U1191 (N_1191,In_1140,In_1861);
nand U1192 (N_1192,In_822,In_1864);
nor U1193 (N_1193,In_1818,In_868);
nor U1194 (N_1194,In_748,In_1436);
or U1195 (N_1195,In_1453,In_1043);
and U1196 (N_1196,In_1102,In_312);
and U1197 (N_1197,In_881,In_323);
and U1198 (N_1198,In_494,In_1499);
nor U1199 (N_1199,In_1328,In_1381);
and U1200 (N_1200,In_924,In_1464);
and U1201 (N_1201,In_622,In_610);
nand U1202 (N_1202,In_611,In_1734);
or U1203 (N_1203,In_815,In_550);
and U1204 (N_1204,In_1817,In_1503);
nand U1205 (N_1205,In_947,In_299);
nand U1206 (N_1206,In_88,In_810);
and U1207 (N_1207,In_958,In_898);
or U1208 (N_1208,In_622,In_869);
nand U1209 (N_1209,In_246,In_755);
nor U1210 (N_1210,In_575,In_51);
nand U1211 (N_1211,In_1282,In_576);
nor U1212 (N_1212,In_1058,In_1602);
nand U1213 (N_1213,In_1747,In_1451);
nor U1214 (N_1214,In_367,In_669);
and U1215 (N_1215,In_1092,In_1963);
and U1216 (N_1216,In_1215,In_1685);
and U1217 (N_1217,In_1118,In_1855);
nand U1218 (N_1218,In_1169,In_571);
xor U1219 (N_1219,In_250,In_899);
or U1220 (N_1220,In_384,In_963);
nor U1221 (N_1221,In_1851,In_1916);
nor U1222 (N_1222,In_715,In_1714);
and U1223 (N_1223,In_1550,In_631);
nor U1224 (N_1224,In_936,In_851);
xnor U1225 (N_1225,In_138,In_218);
and U1226 (N_1226,In_1693,In_369);
nor U1227 (N_1227,In_970,In_1804);
and U1228 (N_1228,In_1366,In_1598);
and U1229 (N_1229,In_679,In_749);
or U1230 (N_1230,In_699,In_1954);
nand U1231 (N_1231,In_1704,In_1791);
or U1232 (N_1232,In_1508,In_1941);
or U1233 (N_1233,In_1483,In_314);
and U1234 (N_1234,In_1765,In_123);
and U1235 (N_1235,In_252,In_560);
or U1236 (N_1236,In_741,In_638);
nor U1237 (N_1237,In_679,In_858);
or U1238 (N_1238,In_1615,In_1773);
nor U1239 (N_1239,In_1256,In_1754);
and U1240 (N_1240,In_634,In_951);
nand U1241 (N_1241,In_545,In_1234);
or U1242 (N_1242,In_222,In_307);
nor U1243 (N_1243,In_1129,In_1352);
nand U1244 (N_1244,In_1154,In_875);
or U1245 (N_1245,In_1197,In_82);
nor U1246 (N_1246,In_1505,In_33);
and U1247 (N_1247,In_337,In_506);
or U1248 (N_1248,In_1683,In_492);
or U1249 (N_1249,In_329,In_1156);
nor U1250 (N_1250,In_1280,In_173);
nor U1251 (N_1251,In_388,In_915);
and U1252 (N_1252,In_812,In_1857);
nor U1253 (N_1253,In_1823,In_1485);
xnor U1254 (N_1254,In_1403,In_1879);
or U1255 (N_1255,In_1428,In_1166);
nor U1256 (N_1256,In_282,In_379);
and U1257 (N_1257,In_1492,In_871);
or U1258 (N_1258,In_435,In_949);
nand U1259 (N_1259,In_649,In_1128);
and U1260 (N_1260,In_260,In_438);
nand U1261 (N_1261,In_708,In_1481);
or U1262 (N_1262,In_1139,In_1674);
nand U1263 (N_1263,In_1627,In_130);
and U1264 (N_1264,In_173,In_946);
nor U1265 (N_1265,In_444,In_437);
nor U1266 (N_1266,In_1973,In_377);
or U1267 (N_1267,In_1988,In_1460);
nand U1268 (N_1268,In_975,In_361);
and U1269 (N_1269,In_1,In_297);
or U1270 (N_1270,In_719,In_1095);
nand U1271 (N_1271,In_1931,In_1340);
or U1272 (N_1272,In_1815,In_112);
and U1273 (N_1273,In_1221,In_19);
nor U1274 (N_1274,In_182,In_1899);
nand U1275 (N_1275,In_157,In_624);
nor U1276 (N_1276,In_201,In_461);
and U1277 (N_1277,In_1979,In_362);
and U1278 (N_1278,In_368,In_1193);
nor U1279 (N_1279,In_898,In_170);
nand U1280 (N_1280,In_1419,In_1040);
or U1281 (N_1281,In_1555,In_1674);
nand U1282 (N_1282,In_1068,In_1495);
nor U1283 (N_1283,In_1330,In_519);
nor U1284 (N_1284,In_1785,In_1452);
or U1285 (N_1285,In_921,In_330);
nand U1286 (N_1286,In_689,In_543);
nor U1287 (N_1287,In_117,In_780);
and U1288 (N_1288,In_1972,In_816);
or U1289 (N_1289,In_744,In_1434);
nor U1290 (N_1290,In_1929,In_1196);
nand U1291 (N_1291,In_222,In_917);
and U1292 (N_1292,In_543,In_1864);
nand U1293 (N_1293,In_1182,In_1918);
nand U1294 (N_1294,In_483,In_463);
nor U1295 (N_1295,In_419,In_1001);
nand U1296 (N_1296,In_692,In_1090);
and U1297 (N_1297,In_644,In_875);
or U1298 (N_1298,In_1296,In_1465);
and U1299 (N_1299,In_457,In_470);
nor U1300 (N_1300,In_485,In_524);
and U1301 (N_1301,In_458,In_905);
nor U1302 (N_1302,In_463,In_1119);
and U1303 (N_1303,In_97,In_454);
nand U1304 (N_1304,In_1366,In_1775);
and U1305 (N_1305,In_994,In_713);
nand U1306 (N_1306,In_1984,In_354);
nand U1307 (N_1307,In_1865,In_420);
nor U1308 (N_1308,In_1749,In_1961);
and U1309 (N_1309,In_1038,In_756);
nand U1310 (N_1310,In_1522,In_497);
and U1311 (N_1311,In_52,In_1777);
nor U1312 (N_1312,In_1569,In_288);
or U1313 (N_1313,In_1330,In_1434);
and U1314 (N_1314,In_1315,In_981);
nand U1315 (N_1315,In_544,In_1524);
and U1316 (N_1316,In_1457,In_78);
nor U1317 (N_1317,In_1591,In_118);
and U1318 (N_1318,In_1868,In_486);
nand U1319 (N_1319,In_722,In_1151);
nand U1320 (N_1320,In_729,In_124);
nand U1321 (N_1321,In_1564,In_1663);
nor U1322 (N_1322,In_1450,In_1258);
or U1323 (N_1323,In_362,In_1305);
and U1324 (N_1324,In_878,In_187);
and U1325 (N_1325,In_717,In_318);
nor U1326 (N_1326,In_948,In_1932);
nor U1327 (N_1327,In_1761,In_525);
nor U1328 (N_1328,In_1373,In_1487);
and U1329 (N_1329,In_1349,In_1441);
nor U1330 (N_1330,In_934,In_1039);
nand U1331 (N_1331,In_419,In_593);
and U1332 (N_1332,In_1927,In_1619);
nor U1333 (N_1333,In_426,In_435);
and U1334 (N_1334,In_107,In_348);
and U1335 (N_1335,In_1052,In_868);
nand U1336 (N_1336,In_824,In_777);
and U1337 (N_1337,In_526,In_399);
and U1338 (N_1338,In_1868,In_433);
nor U1339 (N_1339,In_1651,In_1628);
or U1340 (N_1340,In_62,In_1566);
nand U1341 (N_1341,In_1838,In_1725);
and U1342 (N_1342,In_1574,In_1118);
nor U1343 (N_1343,In_875,In_1844);
nand U1344 (N_1344,In_389,In_1802);
or U1345 (N_1345,In_828,In_898);
nor U1346 (N_1346,In_439,In_1481);
and U1347 (N_1347,In_1315,In_1701);
and U1348 (N_1348,In_207,In_934);
nor U1349 (N_1349,In_174,In_1115);
nand U1350 (N_1350,In_255,In_633);
or U1351 (N_1351,In_45,In_1744);
and U1352 (N_1352,In_1993,In_282);
nor U1353 (N_1353,In_1060,In_676);
nor U1354 (N_1354,In_1848,In_0);
nor U1355 (N_1355,In_722,In_935);
nor U1356 (N_1356,In_1292,In_415);
and U1357 (N_1357,In_658,In_976);
nor U1358 (N_1358,In_1137,In_1086);
nand U1359 (N_1359,In_809,In_241);
or U1360 (N_1360,In_745,In_287);
nor U1361 (N_1361,In_526,In_1927);
or U1362 (N_1362,In_1582,In_892);
nor U1363 (N_1363,In_26,In_83);
and U1364 (N_1364,In_587,In_101);
and U1365 (N_1365,In_1540,In_543);
and U1366 (N_1366,In_719,In_1306);
or U1367 (N_1367,In_1012,In_390);
and U1368 (N_1368,In_404,In_894);
nand U1369 (N_1369,In_559,In_1536);
nand U1370 (N_1370,In_965,In_769);
nor U1371 (N_1371,In_286,In_1478);
or U1372 (N_1372,In_1638,In_1910);
nand U1373 (N_1373,In_793,In_561);
nor U1374 (N_1374,In_195,In_1517);
nand U1375 (N_1375,In_789,In_149);
and U1376 (N_1376,In_905,In_1720);
and U1377 (N_1377,In_1020,In_295);
nand U1378 (N_1378,In_1969,In_973);
and U1379 (N_1379,In_1151,In_1823);
and U1380 (N_1380,In_677,In_223);
or U1381 (N_1381,In_749,In_1143);
or U1382 (N_1382,In_733,In_1043);
and U1383 (N_1383,In_510,In_1827);
nor U1384 (N_1384,In_557,In_818);
and U1385 (N_1385,In_170,In_1743);
nor U1386 (N_1386,In_1696,In_1611);
and U1387 (N_1387,In_1144,In_1290);
and U1388 (N_1388,In_850,In_756);
nor U1389 (N_1389,In_796,In_321);
nor U1390 (N_1390,In_374,In_214);
or U1391 (N_1391,In_19,In_870);
nand U1392 (N_1392,In_211,In_1273);
nand U1393 (N_1393,In_1605,In_399);
nand U1394 (N_1394,In_1816,In_1073);
nor U1395 (N_1395,In_688,In_1823);
nand U1396 (N_1396,In_568,In_455);
or U1397 (N_1397,In_1587,In_1901);
or U1398 (N_1398,In_758,In_1153);
nor U1399 (N_1399,In_1461,In_242);
and U1400 (N_1400,In_1444,In_872);
or U1401 (N_1401,In_427,In_1475);
or U1402 (N_1402,In_1259,In_1712);
or U1403 (N_1403,In_663,In_439);
nand U1404 (N_1404,In_999,In_1201);
or U1405 (N_1405,In_405,In_441);
nor U1406 (N_1406,In_563,In_543);
or U1407 (N_1407,In_216,In_458);
nor U1408 (N_1408,In_1610,In_266);
xor U1409 (N_1409,In_239,In_1057);
or U1410 (N_1410,In_972,In_1657);
or U1411 (N_1411,In_250,In_1802);
nor U1412 (N_1412,In_1060,In_944);
nand U1413 (N_1413,In_1182,In_176);
nor U1414 (N_1414,In_93,In_323);
nor U1415 (N_1415,In_1857,In_1342);
nand U1416 (N_1416,In_251,In_520);
nor U1417 (N_1417,In_1604,In_364);
or U1418 (N_1418,In_472,In_881);
or U1419 (N_1419,In_1212,In_489);
or U1420 (N_1420,In_1289,In_757);
and U1421 (N_1421,In_1619,In_1405);
and U1422 (N_1422,In_233,In_120);
nor U1423 (N_1423,In_727,In_1271);
or U1424 (N_1424,In_1170,In_688);
or U1425 (N_1425,In_381,In_1211);
nor U1426 (N_1426,In_726,In_882);
nor U1427 (N_1427,In_1287,In_73);
or U1428 (N_1428,In_59,In_1598);
nand U1429 (N_1429,In_223,In_389);
nand U1430 (N_1430,In_1133,In_670);
and U1431 (N_1431,In_1914,In_934);
and U1432 (N_1432,In_933,In_1241);
nand U1433 (N_1433,In_216,In_921);
and U1434 (N_1434,In_1797,In_1828);
and U1435 (N_1435,In_958,In_341);
nor U1436 (N_1436,In_1148,In_1182);
nor U1437 (N_1437,In_1521,In_1250);
or U1438 (N_1438,In_789,In_1288);
or U1439 (N_1439,In_874,In_1135);
nor U1440 (N_1440,In_1890,In_516);
and U1441 (N_1441,In_1618,In_1314);
or U1442 (N_1442,In_487,In_979);
nand U1443 (N_1443,In_746,In_1927);
or U1444 (N_1444,In_1400,In_1778);
and U1445 (N_1445,In_1581,In_375);
nand U1446 (N_1446,In_1133,In_1760);
nand U1447 (N_1447,In_30,In_1252);
nand U1448 (N_1448,In_421,In_1778);
and U1449 (N_1449,In_372,In_46);
nand U1450 (N_1450,In_179,In_1181);
nand U1451 (N_1451,In_1768,In_1957);
nand U1452 (N_1452,In_6,In_750);
or U1453 (N_1453,In_102,In_1569);
or U1454 (N_1454,In_1114,In_1390);
and U1455 (N_1455,In_1080,In_720);
nor U1456 (N_1456,In_438,In_838);
and U1457 (N_1457,In_566,In_396);
or U1458 (N_1458,In_808,In_1298);
nand U1459 (N_1459,In_424,In_625);
or U1460 (N_1460,In_554,In_1676);
and U1461 (N_1461,In_1509,In_1688);
nor U1462 (N_1462,In_1899,In_1056);
and U1463 (N_1463,In_392,In_632);
nand U1464 (N_1464,In_785,In_1913);
nand U1465 (N_1465,In_662,In_1906);
or U1466 (N_1466,In_1791,In_508);
or U1467 (N_1467,In_625,In_1548);
and U1468 (N_1468,In_717,In_1655);
or U1469 (N_1469,In_1338,In_1179);
and U1470 (N_1470,In_1111,In_687);
nor U1471 (N_1471,In_984,In_1158);
nand U1472 (N_1472,In_894,In_1173);
nand U1473 (N_1473,In_1140,In_1279);
and U1474 (N_1474,In_1116,In_252);
and U1475 (N_1475,In_1619,In_1767);
nor U1476 (N_1476,In_14,In_941);
or U1477 (N_1477,In_1402,In_17);
nor U1478 (N_1478,In_1989,In_1403);
and U1479 (N_1479,In_420,In_1082);
nand U1480 (N_1480,In_973,In_1009);
nor U1481 (N_1481,In_1141,In_1625);
nand U1482 (N_1482,In_1957,In_501);
and U1483 (N_1483,In_1488,In_20);
nor U1484 (N_1484,In_773,In_1897);
and U1485 (N_1485,In_532,In_453);
nand U1486 (N_1486,In_1886,In_1090);
and U1487 (N_1487,In_564,In_1284);
and U1488 (N_1488,In_169,In_1589);
nand U1489 (N_1489,In_1040,In_1660);
and U1490 (N_1490,In_1971,In_59);
nor U1491 (N_1491,In_1510,In_784);
and U1492 (N_1492,In_1689,In_1098);
and U1493 (N_1493,In_183,In_1103);
or U1494 (N_1494,In_1698,In_24);
or U1495 (N_1495,In_1867,In_192);
or U1496 (N_1496,In_1512,In_1759);
and U1497 (N_1497,In_1307,In_1846);
and U1498 (N_1498,In_1269,In_445);
and U1499 (N_1499,In_1810,In_644);
nand U1500 (N_1500,In_1544,In_1052);
nor U1501 (N_1501,In_1890,In_63);
nor U1502 (N_1502,In_811,In_1367);
nor U1503 (N_1503,In_1818,In_1819);
and U1504 (N_1504,In_1991,In_983);
nor U1505 (N_1505,In_68,In_896);
nor U1506 (N_1506,In_190,In_1588);
nor U1507 (N_1507,In_1677,In_1076);
nor U1508 (N_1508,In_735,In_882);
and U1509 (N_1509,In_1713,In_353);
nand U1510 (N_1510,In_1657,In_1762);
or U1511 (N_1511,In_1469,In_240);
nor U1512 (N_1512,In_488,In_1098);
nand U1513 (N_1513,In_677,In_238);
or U1514 (N_1514,In_939,In_647);
and U1515 (N_1515,In_1434,In_1205);
or U1516 (N_1516,In_891,In_480);
or U1517 (N_1517,In_1683,In_1607);
or U1518 (N_1518,In_1338,In_896);
and U1519 (N_1519,In_530,In_986);
nand U1520 (N_1520,In_278,In_1524);
and U1521 (N_1521,In_416,In_1057);
or U1522 (N_1522,In_650,In_767);
or U1523 (N_1523,In_711,In_84);
or U1524 (N_1524,In_1309,In_1714);
or U1525 (N_1525,In_2,In_1497);
or U1526 (N_1526,In_545,In_1810);
or U1527 (N_1527,In_222,In_1897);
nor U1528 (N_1528,In_1722,In_504);
nand U1529 (N_1529,In_71,In_20);
nor U1530 (N_1530,In_1671,In_727);
nor U1531 (N_1531,In_1659,In_524);
or U1532 (N_1532,In_1445,In_1662);
and U1533 (N_1533,In_1725,In_947);
or U1534 (N_1534,In_1352,In_1391);
nor U1535 (N_1535,In_472,In_1428);
and U1536 (N_1536,In_797,In_744);
nor U1537 (N_1537,In_776,In_71);
and U1538 (N_1538,In_233,In_802);
nor U1539 (N_1539,In_9,In_712);
or U1540 (N_1540,In_104,In_1211);
or U1541 (N_1541,In_1657,In_1363);
nor U1542 (N_1542,In_689,In_643);
and U1543 (N_1543,In_86,In_1403);
and U1544 (N_1544,In_1529,In_1065);
or U1545 (N_1545,In_643,In_1239);
and U1546 (N_1546,In_918,In_258);
nand U1547 (N_1547,In_203,In_1348);
and U1548 (N_1548,In_275,In_1292);
nand U1549 (N_1549,In_327,In_519);
and U1550 (N_1550,In_1191,In_1094);
xor U1551 (N_1551,In_1430,In_1777);
and U1552 (N_1552,In_520,In_1205);
and U1553 (N_1553,In_358,In_208);
nand U1554 (N_1554,In_149,In_225);
nand U1555 (N_1555,In_1636,In_329);
or U1556 (N_1556,In_887,In_86);
nand U1557 (N_1557,In_1183,In_1905);
nand U1558 (N_1558,In_1938,In_1018);
nor U1559 (N_1559,In_1087,In_1310);
and U1560 (N_1560,In_298,In_1535);
and U1561 (N_1561,In_685,In_458);
nor U1562 (N_1562,In_1283,In_1233);
nand U1563 (N_1563,In_1330,In_1693);
and U1564 (N_1564,In_979,In_129);
xor U1565 (N_1565,In_1377,In_994);
nand U1566 (N_1566,In_1843,In_478);
and U1567 (N_1567,In_1231,In_1693);
or U1568 (N_1568,In_489,In_1566);
or U1569 (N_1569,In_1941,In_680);
nand U1570 (N_1570,In_1679,In_348);
nand U1571 (N_1571,In_268,In_151);
or U1572 (N_1572,In_513,In_1620);
or U1573 (N_1573,In_1495,In_1541);
or U1574 (N_1574,In_677,In_1004);
and U1575 (N_1575,In_1875,In_1180);
or U1576 (N_1576,In_676,In_195);
nor U1577 (N_1577,In_188,In_1142);
nor U1578 (N_1578,In_108,In_191);
nand U1579 (N_1579,In_1062,In_1600);
and U1580 (N_1580,In_1009,In_1356);
or U1581 (N_1581,In_1271,In_1532);
and U1582 (N_1582,In_1010,In_1223);
and U1583 (N_1583,In_670,In_1922);
nand U1584 (N_1584,In_1008,In_1525);
nor U1585 (N_1585,In_27,In_84);
nand U1586 (N_1586,In_1759,In_1706);
or U1587 (N_1587,In_376,In_1676);
or U1588 (N_1588,In_685,In_1165);
or U1589 (N_1589,In_1742,In_394);
or U1590 (N_1590,In_282,In_1879);
nand U1591 (N_1591,In_1989,In_1668);
nor U1592 (N_1592,In_1790,In_1097);
and U1593 (N_1593,In_1426,In_823);
or U1594 (N_1594,In_1524,In_1910);
or U1595 (N_1595,In_666,In_1184);
nand U1596 (N_1596,In_514,In_1287);
nor U1597 (N_1597,In_962,In_289);
nand U1598 (N_1598,In_249,In_1515);
or U1599 (N_1599,In_436,In_476);
nor U1600 (N_1600,In_1605,In_1817);
and U1601 (N_1601,In_1672,In_547);
or U1602 (N_1602,In_560,In_1049);
and U1603 (N_1603,In_28,In_189);
or U1604 (N_1604,In_344,In_1558);
nand U1605 (N_1605,In_729,In_1587);
or U1606 (N_1606,In_1816,In_1149);
and U1607 (N_1607,In_567,In_1119);
or U1608 (N_1608,In_1249,In_1469);
nand U1609 (N_1609,In_1736,In_1924);
nand U1610 (N_1610,In_1168,In_1326);
nand U1611 (N_1611,In_29,In_159);
or U1612 (N_1612,In_335,In_626);
or U1613 (N_1613,In_438,In_1378);
and U1614 (N_1614,In_822,In_1779);
and U1615 (N_1615,In_1718,In_89);
and U1616 (N_1616,In_1224,In_51);
and U1617 (N_1617,In_794,In_1126);
and U1618 (N_1618,In_180,In_525);
nor U1619 (N_1619,In_893,In_1322);
nand U1620 (N_1620,In_1162,In_638);
and U1621 (N_1621,In_316,In_1294);
and U1622 (N_1622,In_1036,In_401);
nand U1623 (N_1623,In_1528,In_1214);
nand U1624 (N_1624,In_1954,In_1999);
and U1625 (N_1625,In_853,In_1593);
nand U1626 (N_1626,In_1791,In_1196);
and U1627 (N_1627,In_1601,In_1652);
nor U1628 (N_1628,In_428,In_1975);
or U1629 (N_1629,In_1004,In_1870);
and U1630 (N_1630,In_781,In_201);
and U1631 (N_1631,In_1601,In_367);
or U1632 (N_1632,In_1836,In_1299);
nand U1633 (N_1633,In_1864,In_1655);
and U1634 (N_1634,In_131,In_962);
nand U1635 (N_1635,In_716,In_1516);
nor U1636 (N_1636,In_1329,In_160);
nor U1637 (N_1637,In_732,In_753);
nor U1638 (N_1638,In_844,In_1825);
nand U1639 (N_1639,In_1287,In_719);
or U1640 (N_1640,In_643,In_38);
nor U1641 (N_1641,In_1867,In_591);
nand U1642 (N_1642,In_1646,In_86);
or U1643 (N_1643,In_129,In_686);
or U1644 (N_1644,In_933,In_1507);
or U1645 (N_1645,In_1085,In_646);
nor U1646 (N_1646,In_1698,In_492);
nand U1647 (N_1647,In_1239,In_331);
nand U1648 (N_1648,In_936,In_1643);
or U1649 (N_1649,In_467,In_1245);
nand U1650 (N_1650,In_1828,In_485);
nand U1651 (N_1651,In_1536,In_624);
nor U1652 (N_1652,In_44,In_29);
and U1653 (N_1653,In_205,In_707);
nand U1654 (N_1654,In_1223,In_1699);
or U1655 (N_1655,In_1776,In_350);
nand U1656 (N_1656,In_1052,In_1983);
and U1657 (N_1657,In_208,In_928);
nor U1658 (N_1658,In_748,In_1215);
or U1659 (N_1659,In_330,In_1743);
and U1660 (N_1660,In_1476,In_1870);
or U1661 (N_1661,In_1262,In_864);
or U1662 (N_1662,In_496,In_1181);
or U1663 (N_1663,In_1386,In_1975);
or U1664 (N_1664,In_1045,In_1853);
and U1665 (N_1665,In_944,In_1875);
nand U1666 (N_1666,In_381,In_1602);
nor U1667 (N_1667,In_900,In_1785);
or U1668 (N_1668,In_891,In_1311);
nand U1669 (N_1669,In_1057,In_1510);
or U1670 (N_1670,In_1277,In_600);
nor U1671 (N_1671,In_743,In_748);
nor U1672 (N_1672,In_1618,In_1946);
nor U1673 (N_1673,In_1821,In_499);
and U1674 (N_1674,In_638,In_1976);
and U1675 (N_1675,In_1342,In_861);
nand U1676 (N_1676,In_600,In_1667);
nand U1677 (N_1677,In_924,In_1988);
nand U1678 (N_1678,In_586,In_939);
or U1679 (N_1679,In_345,In_1557);
and U1680 (N_1680,In_1436,In_363);
nor U1681 (N_1681,In_461,In_1292);
and U1682 (N_1682,In_191,In_786);
nand U1683 (N_1683,In_1888,In_1844);
or U1684 (N_1684,In_1761,In_1187);
or U1685 (N_1685,In_1269,In_108);
nor U1686 (N_1686,In_621,In_1329);
or U1687 (N_1687,In_383,In_1486);
and U1688 (N_1688,In_1005,In_1645);
or U1689 (N_1689,In_705,In_1606);
nor U1690 (N_1690,In_1592,In_177);
nand U1691 (N_1691,In_592,In_714);
and U1692 (N_1692,In_25,In_738);
nor U1693 (N_1693,In_1769,In_483);
nor U1694 (N_1694,In_456,In_1385);
nor U1695 (N_1695,In_952,In_920);
and U1696 (N_1696,In_608,In_870);
and U1697 (N_1697,In_1629,In_735);
or U1698 (N_1698,In_130,In_292);
and U1699 (N_1699,In_1987,In_1778);
nor U1700 (N_1700,In_137,In_1547);
and U1701 (N_1701,In_714,In_1862);
nor U1702 (N_1702,In_796,In_1724);
nor U1703 (N_1703,In_1800,In_161);
or U1704 (N_1704,In_850,In_1765);
nand U1705 (N_1705,In_190,In_1385);
nand U1706 (N_1706,In_1235,In_1625);
nor U1707 (N_1707,In_1614,In_1374);
nor U1708 (N_1708,In_1307,In_150);
nand U1709 (N_1709,In_457,In_1658);
nand U1710 (N_1710,In_1065,In_721);
or U1711 (N_1711,In_1469,In_1667);
nor U1712 (N_1712,In_1762,In_1921);
or U1713 (N_1713,In_422,In_397);
or U1714 (N_1714,In_1997,In_514);
or U1715 (N_1715,In_710,In_1382);
nor U1716 (N_1716,In_1531,In_1127);
or U1717 (N_1717,In_1108,In_631);
and U1718 (N_1718,In_466,In_1881);
nand U1719 (N_1719,In_340,In_1999);
nor U1720 (N_1720,In_772,In_1534);
nor U1721 (N_1721,In_698,In_1035);
and U1722 (N_1722,In_1403,In_1093);
or U1723 (N_1723,In_194,In_645);
nand U1724 (N_1724,In_205,In_1543);
or U1725 (N_1725,In_29,In_72);
and U1726 (N_1726,In_718,In_353);
nand U1727 (N_1727,In_1912,In_1686);
nand U1728 (N_1728,In_552,In_1683);
nand U1729 (N_1729,In_1803,In_1530);
and U1730 (N_1730,In_118,In_95);
nand U1731 (N_1731,In_609,In_16);
or U1732 (N_1732,In_1622,In_958);
nand U1733 (N_1733,In_1254,In_418);
nand U1734 (N_1734,In_524,In_1013);
or U1735 (N_1735,In_1423,In_333);
and U1736 (N_1736,In_1794,In_1106);
nand U1737 (N_1737,In_1036,In_930);
or U1738 (N_1738,In_1394,In_1708);
or U1739 (N_1739,In_559,In_308);
or U1740 (N_1740,In_18,In_214);
nor U1741 (N_1741,In_1860,In_254);
nand U1742 (N_1742,In_397,In_624);
and U1743 (N_1743,In_1602,In_93);
nor U1744 (N_1744,In_1671,In_1609);
and U1745 (N_1745,In_1153,In_371);
and U1746 (N_1746,In_1383,In_130);
nand U1747 (N_1747,In_1755,In_39);
and U1748 (N_1748,In_1403,In_1884);
nor U1749 (N_1749,In_251,In_776);
nand U1750 (N_1750,In_1188,In_287);
nor U1751 (N_1751,In_755,In_1269);
or U1752 (N_1752,In_88,In_367);
nor U1753 (N_1753,In_1869,In_1350);
nand U1754 (N_1754,In_772,In_1993);
or U1755 (N_1755,In_490,In_320);
or U1756 (N_1756,In_1690,In_1023);
and U1757 (N_1757,In_1,In_53);
and U1758 (N_1758,In_96,In_293);
or U1759 (N_1759,In_1799,In_151);
nand U1760 (N_1760,In_161,In_383);
nor U1761 (N_1761,In_235,In_1063);
nand U1762 (N_1762,In_747,In_204);
nand U1763 (N_1763,In_1371,In_684);
or U1764 (N_1764,In_1777,In_270);
nand U1765 (N_1765,In_1960,In_1846);
nand U1766 (N_1766,In_921,In_259);
nor U1767 (N_1767,In_612,In_1898);
nor U1768 (N_1768,In_1267,In_1547);
nand U1769 (N_1769,In_1697,In_1328);
and U1770 (N_1770,In_156,In_551);
nand U1771 (N_1771,In_359,In_393);
nand U1772 (N_1772,In_446,In_1935);
nor U1773 (N_1773,In_626,In_1632);
nand U1774 (N_1774,In_1393,In_1099);
nand U1775 (N_1775,In_907,In_1838);
or U1776 (N_1776,In_129,In_687);
nor U1777 (N_1777,In_296,In_1981);
nand U1778 (N_1778,In_167,In_541);
or U1779 (N_1779,In_660,In_186);
nor U1780 (N_1780,In_154,In_941);
or U1781 (N_1781,In_719,In_861);
or U1782 (N_1782,In_475,In_1668);
nor U1783 (N_1783,In_829,In_1865);
and U1784 (N_1784,In_1209,In_1944);
or U1785 (N_1785,In_1214,In_1534);
nand U1786 (N_1786,In_1437,In_509);
nand U1787 (N_1787,In_1558,In_472);
xnor U1788 (N_1788,In_543,In_1399);
and U1789 (N_1789,In_479,In_1653);
and U1790 (N_1790,In_755,In_1625);
nor U1791 (N_1791,In_1913,In_134);
and U1792 (N_1792,In_1168,In_917);
or U1793 (N_1793,In_1722,In_873);
xor U1794 (N_1794,In_540,In_911);
and U1795 (N_1795,In_200,In_347);
and U1796 (N_1796,In_915,In_764);
nand U1797 (N_1797,In_488,In_1116);
and U1798 (N_1798,In_1750,In_1274);
and U1799 (N_1799,In_1893,In_69);
nor U1800 (N_1800,In_1803,In_1772);
or U1801 (N_1801,In_439,In_648);
nand U1802 (N_1802,In_745,In_1104);
and U1803 (N_1803,In_511,In_1683);
nand U1804 (N_1804,In_1574,In_121);
nand U1805 (N_1805,In_58,In_1653);
and U1806 (N_1806,In_758,In_1384);
nor U1807 (N_1807,In_725,In_1885);
or U1808 (N_1808,In_1977,In_1893);
nand U1809 (N_1809,In_1801,In_1449);
and U1810 (N_1810,In_1230,In_110);
or U1811 (N_1811,In_288,In_439);
nand U1812 (N_1812,In_129,In_210);
or U1813 (N_1813,In_1852,In_1165);
and U1814 (N_1814,In_855,In_798);
nor U1815 (N_1815,In_652,In_1607);
nor U1816 (N_1816,In_1888,In_1630);
or U1817 (N_1817,In_1333,In_178);
or U1818 (N_1818,In_1275,In_911);
nand U1819 (N_1819,In_313,In_531);
nand U1820 (N_1820,In_1163,In_1374);
nand U1821 (N_1821,In_1207,In_1617);
and U1822 (N_1822,In_1654,In_1721);
or U1823 (N_1823,In_1244,In_1400);
or U1824 (N_1824,In_1124,In_1226);
nand U1825 (N_1825,In_1029,In_1548);
nor U1826 (N_1826,In_653,In_304);
nand U1827 (N_1827,In_1195,In_106);
nand U1828 (N_1828,In_1358,In_1414);
nor U1829 (N_1829,In_1245,In_523);
nand U1830 (N_1830,In_914,In_606);
and U1831 (N_1831,In_1274,In_1911);
nor U1832 (N_1832,In_1529,In_1456);
or U1833 (N_1833,In_1873,In_249);
and U1834 (N_1834,In_1484,In_1609);
and U1835 (N_1835,In_333,In_1379);
nand U1836 (N_1836,In_427,In_1420);
or U1837 (N_1837,In_1578,In_366);
nand U1838 (N_1838,In_1849,In_1547);
and U1839 (N_1839,In_792,In_1849);
and U1840 (N_1840,In_672,In_1129);
or U1841 (N_1841,In_769,In_369);
nor U1842 (N_1842,In_1399,In_537);
nand U1843 (N_1843,In_240,In_366);
and U1844 (N_1844,In_980,In_1372);
and U1845 (N_1845,In_737,In_1728);
nor U1846 (N_1846,In_946,In_635);
or U1847 (N_1847,In_1384,In_279);
nor U1848 (N_1848,In_1892,In_325);
and U1849 (N_1849,In_935,In_46);
or U1850 (N_1850,In_331,In_505);
nor U1851 (N_1851,In_1452,In_1488);
and U1852 (N_1852,In_503,In_1063);
or U1853 (N_1853,In_1455,In_1649);
and U1854 (N_1854,In_345,In_1839);
and U1855 (N_1855,In_1585,In_892);
nand U1856 (N_1856,In_805,In_1872);
or U1857 (N_1857,In_3,In_691);
nand U1858 (N_1858,In_1091,In_1131);
nand U1859 (N_1859,In_281,In_86);
nor U1860 (N_1860,In_290,In_1757);
and U1861 (N_1861,In_1548,In_334);
nand U1862 (N_1862,In_450,In_1952);
nand U1863 (N_1863,In_1282,In_1616);
xnor U1864 (N_1864,In_1508,In_1051);
nand U1865 (N_1865,In_1297,In_1735);
and U1866 (N_1866,In_1250,In_1108);
or U1867 (N_1867,In_1083,In_41);
nand U1868 (N_1868,In_1154,In_100);
xnor U1869 (N_1869,In_862,In_1295);
nor U1870 (N_1870,In_1962,In_228);
and U1871 (N_1871,In_797,In_808);
nor U1872 (N_1872,In_828,In_581);
nand U1873 (N_1873,In_476,In_1835);
and U1874 (N_1874,In_707,In_1781);
xor U1875 (N_1875,In_551,In_1514);
and U1876 (N_1876,In_1776,In_1957);
and U1877 (N_1877,In_1889,In_288);
nor U1878 (N_1878,In_1853,In_644);
nor U1879 (N_1879,In_1441,In_353);
or U1880 (N_1880,In_1398,In_1864);
or U1881 (N_1881,In_1477,In_783);
and U1882 (N_1882,In_996,In_410);
nand U1883 (N_1883,In_1611,In_1409);
or U1884 (N_1884,In_1265,In_1003);
nor U1885 (N_1885,In_604,In_1641);
and U1886 (N_1886,In_726,In_39);
or U1887 (N_1887,In_291,In_1363);
nand U1888 (N_1888,In_1480,In_71);
nand U1889 (N_1889,In_805,In_261);
nand U1890 (N_1890,In_1313,In_261);
nor U1891 (N_1891,In_719,In_1357);
and U1892 (N_1892,In_614,In_1999);
and U1893 (N_1893,In_667,In_1063);
nand U1894 (N_1894,In_106,In_765);
nor U1895 (N_1895,In_469,In_432);
or U1896 (N_1896,In_716,In_1407);
or U1897 (N_1897,In_1825,In_199);
or U1898 (N_1898,In_558,In_1504);
or U1899 (N_1899,In_1724,In_51);
nor U1900 (N_1900,In_872,In_154);
nand U1901 (N_1901,In_732,In_1231);
nand U1902 (N_1902,In_550,In_772);
nor U1903 (N_1903,In_1775,In_901);
and U1904 (N_1904,In_607,In_800);
and U1905 (N_1905,In_823,In_1110);
nor U1906 (N_1906,In_1596,In_516);
and U1907 (N_1907,In_523,In_309);
nor U1908 (N_1908,In_639,In_1624);
nor U1909 (N_1909,In_450,In_1165);
nand U1910 (N_1910,In_168,In_446);
nand U1911 (N_1911,In_1345,In_1919);
nand U1912 (N_1912,In_1151,In_1406);
nand U1913 (N_1913,In_1402,In_788);
and U1914 (N_1914,In_353,In_1213);
nand U1915 (N_1915,In_489,In_1646);
nor U1916 (N_1916,In_194,In_1276);
nand U1917 (N_1917,In_993,In_1806);
and U1918 (N_1918,In_1712,In_1540);
nand U1919 (N_1919,In_729,In_1011);
or U1920 (N_1920,In_1935,In_1276);
or U1921 (N_1921,In_69,In_966);
nor U1922 (N_1922,In_704,In_1989);
and U1923 (N_1923,In_560,In_1641);
or U1924 (N_1924,In_1910,In_720);
and U1925 (N_1925,In_1733,In_1555);
and U1926 (N_1926,In_487,In_1702);
and U1927 (N_1927,In_516,In_1416);
and U1928 (N_1928,In_1880,In_945);
nor U1929 (N_1929,In_138,In_45);
or U1930 (N_1930,In_698,In_302);
nor U1931 (N_1931,In_1048,In_1883);
or U1932 (N_1932,In_1782,In_1929);
nor U1933 (N_1933,In_611,In_1789);
nand U1934 (N_1934,In_1676,In_547);
or U1935 (N_1935,In_1749,In_1245);
or U1936 (N_1936,In_1258,In_388);
or U1937 (N_1937,In_1910,In_169);
nor U1938 (N_1938,In_517,In_978);
and U1939 (N_1939,In_1034,In_1862);
nand U1940 (N_1940,In_1177,In_1771);
and U1941 (N_1941,In_1656,In_770);
nor U1942 (N_1942,In_1983,In_1450);
and U1943 (N_1943,In_616,In_1751);
nor U1944 (N_1944,In_275,In_458);
nand U1945 (N_1945,In_11,In_303);
or U1946 (N_1946,In_1637,In_328);
nor U1947 (N_1947,In_164,In_262);
nand U1948 (N_1948,In_1054,In_1372);
nand U1949 (N_1949,In_916,In_1984);
nand U1950 (N_1950,In_306,In_1827);
or U1951 (N_1951,In_1281,In_1337);
nor U1952 (N_1952,In_327,In_1967);
and U1953 (N_1953,In_717,In_762);
nor U1954 (N_1954,In_936,In_1543);
nor U1955 (N_1955,In_1137,In_5);
or U1956 (N_1956,In_649,In_107);
nor U1957 (N_1957,In_836,In_216);
nor U1958 (N_1958,In_1623,In_1594);
or U1959 (N_1959,In_1841,In_384);
nand U1960 (N_1960,In_530,In_261);
nand U1961 (N_1961,In_528,In_1086);
nand U1962 (N_1962,In_1602,In_176);
nand U1963 (N_1963,In_58,In_457);
nand U1964 (N_1964,In_101,In_1835);
nand U1965 (N_1965,In_1870,In_1212);
nor U1966 (N_1966,In_1135,In_206);
or U1967 (N_1967,In_745,In_850);
nor U1968 (N_1968,In_922,In_1781);
nor U1969 (N_1969,In_957,In_1647);
and U1970 (N_1970,In_492,In_450);
or U1971 (N_1971,In_1291,In_120);
or U1972 (N_1972,In_1981,In_317);
xnor U1973 (N_1973,In_1182,In_551);
nand U1974 (N_1974,In_1319,In_391);
xor U1975 (N_1975,In_937,In_156);
nor U1976 (N_1976,In_443,In_1650);
and U1977 (N_1977,In_641,In_1827);
nand U1978 (N_1978,In_631,In_1216);
nor U1979 (N_1979,In_1909,In_1132);
and U1980 (N_1980,In_1245,In_405);
and U1981 (N_1981,In_1772,In_1499);
nor U1982 (N_1982,In_361,In_257);
xnor U1983 (N_1983,In_864,In_290);
nand U1984 (N_1984,In_921,In_638);
and U1985 (N_1985,In_1625,In_1691);
and U1986 (N_1986,In_1986,In_957);
or U1987 (N_1987,In_680,In_131);
nor U1988 (N_1988,In_1364,In_473);
nand U1989 (N_1989,In_1,In_117);
or U1990 (N_1990,In_1634,In_1894);
nor U1991 (N_1991,In_423,In_851);
nor U1992 (N_1992,In_1372,In_1718);
or U1993 (N_1993,In_1450,In_1028);
nand U1994 (N_1994,In_1418,In_546);
nand U1995 (N_1995,In_720,In_1488);
nand U1996 (N_1996,In_272,In_1671);
and U1997 (N_1997,In_1638,In_1089);
or U1998 (N_1998,In_567,In_724);
and U1999 (N_1999,In_142,In_525);
or U2000 (N_2000,N_1654,N_930);
nand U2001 (N_2001,N_1475,N_1775);
and U2002 (N_2002,N_1983,N_716);
nand U2003 (N_2003,N_1341,N_537);
nand U2004 (N_2004,N_1295,N_1995);
nand U2005 (N_2005,N_1910,N_1687);
nand U2006 (N_2006,N_558,N_953);
nor U2007 (N_2007,N_1957,N_71);
and U2008 (N_2008,N_1879,N_162);
nor U2009 (N_2009,N_161,N_11);
and U2010 (N_2010,N_977,N_330);
nand U2011 (N_2011,N_90,N_324);
or U2012 (N_2012,N_925,N_1579);
and U2013 (N_2013,N_163,N_1316);
or U2014 (N_2014,N_383,N_1195);
nand U2015 (N_2015,N_1999,N_1671);
or U2016 (N_2016,N_1478,N_1078);
nand U2017 (N_2017,N_580,N_1784);
and U2018 (N_2018,N_1126,N_531);
nor U2019 (N_2019,N_1806,N_1206);
xor U2020 (N_2020,N_1972,N_1681);
or U2021 (N_2021,N_1889,N_1301);
nand U2022 (N_2022,N_1779,N_1915);
or U2023 (N_2023,N_434,N_1383);
or U2024 (N_2024,N_1019,N_1607);
and U2025 (N_2025,N_181,N_1457);
and U2026 (N_2026,N_250,N_44);
nor U2027 (N_2027,N_515,N_209);
nor U2028 (N_2028,N_217,N_145);
or U2029 (N_2029,N_129,N_1861);
or U2030 (N_2030,N_282,N_13);
nand U2031 (N_2031,N_1192,N_1270);
nand U2032 (N_2032,N_1535,N_1296);
and U2033 (N_2033,N_684,N_584);
nand U2034 (N_2034,N_205,N_271);
and U2035 (N_2035,N_1197,N_1893);
nand U2036 (N_2036,N_1808,N_751);
nand U2037 (N_2037,N_933,N_1146);
and U2038 (N_2038,N_306,N_1318);
or U2039 (N_2039,N_1143,N_1596);
and U2040 (N_2040,N_171,N_1015);
or U2041 (N_2041,N_960,N_1070);
nor U2042 (N_2042,N_1561,N_381);
nand U2043 (N_2043,N_298,N_64);
nor U2044 (N_2044,N_34,N_1500);
nand U2045 (N_2045,N_302,N_1660);
or U2046 (N_2046,N_1831,N_1502);
or U2047 (N_2047,N_22,N_854);
or U2048 (N_2048,N_93,N_1066);
or U2049 (N_2049,N_834,N_848);
or U2050 (N_2050,N_241,N_42);
or U2051 (N_2051,N_313,N_506);
xnor U2052 (N_2052,N_1486,N_1555);
and U2053 (N_2053,N_1191,N_1073);
xnor U2054 (N_2054,N_1700,N_1683);
and U2055 (N_2055,N_1127,N_1437);
nor U2056 (N_2056,N_1274,N_1372);
or U2057 (N_2057,N_206,N_1046);
and U2058 (N_2058,N_1042,N_1719);
or U2059 (N_2059,N_1794,N_1242);
or U2060 (N_2060,N_299,N_1175);
and U2061 (N_2061,N_51,N_1501);
and U2062 (N_2062,N_375,N_144);
or U2063 (N_2063,N_649,N_802);
nand U2064 (N_2064,N_1346,N_1853);
nor U2065 (N_2065,N_1967,N_1287);
nor U2066 (N_2066,N_1503,N_1940);
nand U2067 (N_2067,N_1132,N_365);
or U2068 (N_2068,N_267,N_653);
or U2069 (N_2069,N_1523,N_1416);
or U2070 (N_2070,N_53,N_208);
or U2071 (N_2071,N_619,N_1674);
nor U2072 (N_2072,N_692,N_19);
nand U2073 (N_2073,N_1487,N_1053);
or U2074 (N_2074,N_1268,N_1842);
nand U2075 (N_2075,N_12,N_1543);
and U2076 (N_2076,N_165,N_147);
and U2077 (N_2077,N_1797,N_1067);
or U2078 (N_2078,N_588,N_1215);
nand U2079 (N_2079,N_429,N_1360);
and U2080 (N_2080,N_1944,N_800);
or U2081 (N_2081,N_103,N_456);
or U2082 (N_2082,N_743,N_1116);
and U2083 (N_2083,N_52,N_362);
nand U2084 (N_2084,N_1311,N_808);
xor U2085 (N_2085,N_762,N_1920);
nand U2086 (N_2086,N_155,N_469);
nor U2087 (N_2087,N_244,N_1337);
and U2088 (N_2088,N_1027,N_352);
or U2089 (N_2089,N_1599,N_693);
or U2090 (N_2090,N_308,N_650);
nor U2091 (N_2091,N_1955,N_715);
nand U2092 (N_2092,N_221,N_571);
and U2093 (N_2093,N_1905,N_1895);
nand U2094 (N_2094,N_1964,N_310);
or U2095 (N_2095,N_113,N_307);
nand U2096 (N_2096,N_1716,N_47);
or U2097 (N_2097,N_1682,N_1664);
and U2098 (N_2098,N_1379,N_242);
and U2099 (N_2099,N_104,N_1025);
nand U2100 (N_2100,N_461,N_1385);
and U2101 (N_2101,N_1836,N_1460);
nand U2102 (N_2102,N_245,N_1426);
and U2103 (N_2103,N_1373,N_1355);
and U2104 (N_2104,N_1581,N_1858);
nand U2105 (N_2105,N_1627,N_1584);
nor U2106 (N_2106,N_397,N_1239);
nor U2107 (N_2107,N_1470,N_1041);
nor U2108 (N_2108,N_927,N_1894);
nor U2109 (N_2109,N_1252,N_570);
and U2110 (N_2110,N_1878,N_1254);
and U2111 (N_2111,N_86,N_230);
nor U2112 (N_2112,N_1589,N_1171);
or U2113 (N_2113,N_201,N_884);
or U2114 (N_2114,N_822,N_1266);
and U2115 (N_2115,N_380,N_5);
or U2116 (N_2116,N_1233,N_756);
or U2117 (N_2117,N_1058,N_29);
nand U2118 (N_2118,N_855,N_475);
or U2119 (N_2119,N_1100,N_688);
nand U2120 (N_2120,N_1077,N_556);
and U2121 (N_2121,N_830,N_1272);
xnor U2122 (N_2122,N_439,N_1404);
nor U2123 (N_2123,N_1976,N_1873);
or U2124 (N_2124,N_581,N_615);
nor U2125 (N_2125,N_1782,N_1286);
and U2126 (N_2126,N_1044,N_143);
nor U2127 (N_2127,N_745,N_33);
or U2128 (N_2128,N_175,N_341);
and U2129 (N_2129,N_266,N_1697);
and U2130 (N_2130,N_664,N_281);
or U2131 (N_2131,N_1986,N_26);
or U2132 (N_2132,N_1557,N_1668);
or U2133 (N_2133,N_1803,N_1098);
nor U2134 (N_2134,N_1055,N_1248);
and U2135 (N_2135,N_1706,N_316);
nor U2136 (N_2136,N_1819,N_782);
and U2137 (N_2137,N_1780,N_1510);
nand U2138 (N_2138,N_699,N_1768);
nor U2139 (N_2139,N_1689,N_852);
and U2140 (N_2140,N_1332,N_1409);
nor U2141 (N_2141,N_998,N_1860);
or U2142 (N_2142,N_734,N_1635);
nor U2143 (N_2143,N_376,N_1834);
or U2144 (N_2144,N_1956,N_1425);
nor U2145 (N_2145,N_82,N_1913);
and U2146 (N_2146,N_17,N_797);
nor U2147 (N_2147,N_74,N_1473);
nor U2148 (N_2148,N_1419,N_771);
and U2149 (N_2149,N_864,N_717);
nor U2150 (N_2150,N_679,N_671);
and U2151 (N_2151,N_120,N_228);
and U2152 (N_2152,N_1317,N_421);
or U2153 (N_2153,N_520,N_983);
nand U2154 (N_2154,N_1892,N_1507);
nor U2155 (N_2155,N_958,N_1748);
nor U2156 (N_2156,N_1315,N_1488);
or U2157 (N_2157,N_15,N_423);
or U2158 (N_2158,N_632,N_1408);
and U2159 (N_2159,N_334,N_1139);
nor U2160 (N_2160,N_1929,N_1764);
and U2161 (N_2161,N_1129,N_1928);
and U2162 (N_2162,N_567,N_411);
and U2163 (N_2163,N_1282,N_1628);
nor U2164 (N_2164,N_1908,N_1050);
nor U2165 (N_2165,N_1189,N_873);
nor U2166 (N_2166,N_1556,N_246);
nor U2167 (N_2167,N_318,N_465);
and U2168 (N_2168,N_262,N_1812);
and U2169 (N_2169,N_658,N_433);
nor U2170 (N_2170,N_1199,N_1006);
or U2171 (N_2171,N_1981,N_151);
and U2172 (N_2172,N_521,N_1529);
and U2173 (N_2173,N_50,N_1303);
and U2174 (N_2174,N_623,N_753);
and U2175 (N_2175,N_417,N_1875);
and U2176 (N_2176,N_1839,N_735);
or U2177 (N_2177,N_160,N_1182);
and U2178 (N_2178,N_1977,N_1791);
or U2179 (N_2179,N_1212,N_1902);
nor U2180 (N_2180,N_133,N_900);
nand U2181 (N_2181,N_1644,N_911);
nand U2182 (N_2182,N_709,N_754);
nor U2183 (N_2183,N_1708,N_1134);
nor U2184 (N_2184,N_661,N_270);
or U2185 (N_2185,N_1594,N_593);
nor U2186 (N_2186,N_849,N_952);
or U2187 (N_2187,N_283,N_744);
nand U2188 (N_2188,N_1749,N_583);
nand U2189 (N_2189,N_861,N_440);
nor U2190 (N_2190,N_1676,N_1474);
nor U2191 (N_2191,N_339,N_264);
nand U2192 (N_2192,N_1484,N_1265);
nand U2193 (N_2193,N_1445,N_257);
nand U2194 (N_2194,N_1970,N_1769);
or U2195 (N_2195,N_895,N_824);
and U2196 (N_2196,N_1813,N_1651);
nor U2197 (N_2197,N_1863,N_1397);
nor U2198 (N_2198,N_342,N_94);
nor U2199 (N_2199,N_1653,N_1969);
nor U2200 (N_2200,N_712,N_956);
nand U2201 (N_2201,N_872,N_424);
or U2202 (N_2202,N_81,N_1342);
nand U2203 (N_2203,N_89,N_111);
or U2204 (N_2204,N_1188,N_1792);
and U2205 (N_2205,N_1824,N_1950);
nand U2206 (N_2206,N_792,N_1637);
or U2207 (N_2207,N_741,N_415);
and U2208 (N_2208,N_123,N_356);
or U2209 (N_2209,N_1766,N_1264);
nor U2210 (N_2210,N_1776,N_1020);
and U2211 (N_2211,N_490,N_533);
nor U2212 (N_2212,N_839,N_182);
or U2213 (N_2213,N_609,N_249);
nand U2214 (N_2214,N_1176,N_156);
nand U2215 (N_2215,N_1851,N_1026);
or U2216 (N_2216,N_586,N_368);
nand U2217 (N_2217,N_1288,N_1525);
nand U2218 (N_2218,N_1711,N_951);
nor U2219 (N_2219,N_1917,N_1490);
or U2220 (N_2220,N_1434,N_1647);
nor U2221 (N_2221,N_562,N_1057);
nand U2222 (N_2222,N_829,N_1843);
and U2223 (N_2223,N_638,N_1211);
and U2224 (N_2224,N_1773,N_1045);
nor U2225 (N_2225,N_1411,N_1008);
or U2226 (N_2226,N_1805,N_1850);
and U2227 (N_2227,N_1076,N_237);
or U2228 (N_2228,N_494,N_1430);
nand U2229 (N_2229,N_174,N_678);
or U2230 (N_2230,N_560,N_1688);
xor U2231 (N_2231,N_1323,N_578);
nor U2232 (N_2232,N_179,N_1418);
nor U2233 (N_2233,N_636,N_385);
nor U2234 (N_2234,N_323,N_932);
and U2235 (N_2235,N_1033,N_1241);
nor U2236 (N_2236,N_1174,N_991);
and U2237 (N_2237,N_1110,N_523);
or U2238 (N_2238,N_351,N_301);
nor U2239 (N_2239,N_1690,N_1225);
nand U2240 (N_2240,N_577,N_1335);
nor U2241 (N_2241,N_1573,N_1344);
nor U2242 (N_2242,N_1312,N_974);
and U2243 (N_2243,N_305,N_1043);
nand U2244 (N_2244,N_1642,N_997);
nor U2245 (N_2245,N_1975,N_367);
and U2246 (N_2246,N_1403,N_1996);
and U2247 (N_2247,N_37,N_1240);
or U2248 (N_2248,N_1338,N_1722);
nor U2249 (N_2249,N_1289,N_360);
nand U2250 (N_2250,N_812,N_467);
or U2251 (N_2251,N_818,N_168);
xor U2252 (N_2252,N_1513,N_134);
nand U2253 (N_2253,N_1809,N_651);
and U2254 (N_2254,N_277,N_1083);
or U2255 (N_2255,N_1105,N_1923);
or U2256 (N_2256,N_730,N_532);
nor U2257 (N_2257,N_1941,N_1800);
and U2258 (N_2258,N_216,N_1151);
and U2259 (N_2259,N_396,N_1250);
or U2260 (N_2260,N_1514,N_1984);
nor U2261 (N_2261,N_1997,N_41);
nand U2262 (N_2262,N_1161,N_784);
nand U2263 (N_2263,N_187,N_729);
nand U2264 (N_2264,N_1082,N_70);
and U2265 (N_2265,N_1302,N_297);
and U2266 (N_2266,N_964,N_61);
nor U2267 (N_2267,N_1547,N_1833);
nor U2268 (N_2268,N_659,N_164);
and U2269 (N_2269,N_1063,N_137);
nand U2270 (N_2270,N_377,N_1278);
nor U2271 (N_2271,N_1872,N_826);
nor U2272 (N_2272,N_1592,N_763);
and U2273 (N_2273,N_1612,N_700);
nand U2274 (N_2274,N_1115,N_1621);
nor U2275 (N_2275,N_1365,N_1680);
or U2276 (N_2276,N_665,N_1150);
nand U2277 (N_2277,N_1770,N_1414);
and U2278 (N_2278,N_1217,N_1125);
nor U2279 (N_2279,N_1155,N_99);
and U2280 (N_2280,N_592,N_1060);
and U2281 (N_2281,N_598,N_1994);
and U2282 (N_2282,N_1595,N_1079);
nor U2283 (N_2283,N_259,N_176);
nor U2284 (N_2284,N_1458,N_315);
and U2285 (N_2285,N_1085,N_1597);
nor U2286 (N_2286,N_1630,N_1691);
nor U2287 (N_2287,N_810,N_149);
and U2288 (N_2288,N_1269,N_519);
nand U2289 (N_2289,N_867,N_1799);
nand U2290 (N_2290,N_1421,N_290);
or U2291 (N_2291,N_138,N_1754);
nand U2292 (N_2292,N_1821,N_1904);
nand U2293 (N_2293,N_685,N_1971);
nor U2294 (N_2294,N_1389,N_1712);
nand U2295 (N_2295,N_1101,N_1329);
nand U2296 (N_2296,N_1614,N_1030);
or U2297 (N_2297,N_1260,N_1652);
nor U2298 (N_2298,N_476,N_68);
or U2299 (N_2299,N_1147,N_1334);
and U2300 (N_2300,N_642,N_496);
nor U2301 (N_2301,N_210,N_1013);
nand U2302 (N_2302,N_1855,N_1731);
nand U2303 (N_2303,N_1222,N_1795);
nor U2304 (N_2304,N_202,N_935);
nand U2305 (N_2305,N_1159,N_1307);
or U2306 (N_2306,N_1750,N_1518);
nor U2307 (N_2307,N_1559,N_1485);
and U2308 (N_2308,N_1505,N_887);
nand U2309 (N_2309,N_1005,N_1292);
nor U2310 (N_2310,N_764,N_117);
nor U2311 (N_2311,N_1393,N_1281);
and U2312 (N_2312,N_321,N_488);
or U2313 (N_2313,N_1112,N_1720);
nor U2314 (N_2314,N_1565,N_1531);
and U2315 (N_2315,N_1131,N_255);
nand U2316 (N_2316,N_454,N_527);
and U2317 (N_2317,N_414,N_406);
nor U2318 (N_2318,N_837,N_84);
or U2319 (N_2319,N_1616,N_1570);
and U2320 (N_2320,N_916,N_1152);
or U2321 (N_2321,N_1351,N_1890);
and U2322 (N_2322,N_166,N_723);
and U2323 (N_2323,N_1162,N_992);
or U2324 (N_2324,N_1608,N_364);
or U2325 (N_2325,N_881,N_680);
xor U2326 (N_2326,N_3,N_1932);
nor U2327 (N_2327,N_1183,N_379);
and U2328 (N_2328,N_1789,N_758);
or U2329 (N_2329,N_1745,N_1758);
and U2330 (N_2330,N_668,N_1601);
or U2331 (N_2331,N_1477,N_934);
and U2332 (N_2332,N_590,N_211);
and U2333 (N_2333,N_1440,N_938);
nor U2334 (N_2334,N_1386,N_1390);
nand U2335 (N_2335,N_1636,N_1925);
nand U2336 (N_2336,N_1919,N_1947);
or U2337 (N_2337,N_254,N_616);
and U2338 (N_2338,N_1609,N_1056);
nand U2339 (N_2339,N_1548,N_789);
and U2340 (N_2340,N_1065,N_919);
or U2341 (N_2341,N_199,N_1086);
or U2342 (N_2342,N_407,N_1811);
and U2343 (N_2343,N_564,N_1271);
and U2344 (N_2344,N_1516,N_981);
nor U2345 (N_2345,N_1898,N_691);
nand U2346 (N_2346,N_1023,N_273);
nand U2347 (N_2347,N_1255,N_1364);
nor U2348 (N_2348,N_197,N_1590);
or U2349 (N_2349,N_338,N_1762);
nor U2350 (N_2350,N_1366,N_814);
nor U2351 (N_2351,N_1347,N_1450);
nor U2352 (N_2352,N_336,N_189);
or U2353 (N_2353,N_1359,N_1499);
or U2354 (N_2354,N_428,N_234);
nand U2355 (N_2355,N_832,N_885);
nor U2356 (N_2356,N_1498,N_1140);
nor U2357 (N_2357,N_198,N_1737);
or U2358 (N_2358,N_652,N_1244);
or U2359 (N_2359,N_1992,N_1857);
or U2360 (N_2360,N_77,N_759);
or U2361 (N_2361,N_512,N_1822);
nor U2362 (N_2362,N_431,N_403);
nor U2363 (N_2363,N_1088,N_1071);
and U2364 (N_2364,N_122,N_393);
or U2365 (N_2365,N_1021,N_227);
or U2366 (N_2366,N_1294,N_1771);
nor U2367 (N_2367,N_1228,N_224);
and U2368 (N_2368,N_1208,N_1884);
nand U2369 (N_2369,N_1184,N_1675);
nand U2370 (N_2370,N_453,N_1849);
and U2371 (N_2371,N_576,N_942);
or U2372 (N_2372,N_517,N_472);
or U2373 (N_2373,N_1847,N_1009);
or U2374 (N_2374,N_999,N_425);
nand U2375 (N_2375,N_158,N_1862);
nand U2376 (N_2376,N_621,N_435);
nand U2377 (N_2377,N_474,N_223);
nand U2378 (N_2378,N_1693,N_98);
and U2379 (N_2379,N_1090,N_1136);
or U2380 (N_2380,N_1550,N_1968);
nor U2381 (N_2381,N_728,N_449);
nand U2382 (N_2382,N_720,N_1883);
nand U2383 (N_2383,N_550,N_889);
and U2384 (N_2384,N_838,N_1449);
nand U2385 (N_2385,N_420,N_194);
and U2386 (N_2386,N_528,N_833);
or U2387 (N_2387,N_1464,N_1452);
and U2388 (N_2388,N_464,N_1456);
or U2389 (N_2389,N_1804,N_513);
nor U2390 (N_2390,N_1528,N_1432);
or U2391 (N_2391,N_1137,N_1541);
nand U2392 (N_2392,N_278,N_967);
or U2393 (N_2393,N_1837,N_275);
or U2394 (N_2394,N_1939,N_480);
nor U2395 (N_2395,N_1887,N_54);
nor U2396 (N_2396,N_401,N_767);
and U2397 (N_2397,N_1280,N_49);
nor U2398 (N_2398,N_561,N_1870);
or U2399 (N_2399,N_1761,N_252);
nor U2400 (N_2400,N_1966,N_1562);
and U2401 (N_2401,N_755,N_121);
nand U2402 (N_2402,N_1661,N_1190);
or U2403 (N_2403,N_1276,N_647);
or U2404 (N_2404,N_1869,N_689);
nor U2405 (N_2405,N_25,N_45);
nor U2406 (N_2406,N_1459,N_618);
and U2407 (N_2407,N_1061,N_59);
or U2408 (N_2408,N_775,N_1882);
nand U2409 (N_2409,N_914,N_1102);
nor U2410 (N_2410,N_777,N_1625);
and U2411 (N_2411,N_1508,N_768);
or U2412 (N_2412,N_1376,N_1059);
or U2413 (N_2413,N_1428,N_1168);
and U2414 (N_2414,N_43,N_157);
nor U2415 (N_2415,N_1527,N_1238);
nand U2416 (N_2416,N_460,N_863);
and U2417 (N_2417,N_1031,N_293);
nor U2418 (N_2418,N_845,N_805);
and U2419 (N_2419,N_870,N_1924);
nand U2420 (N_2420,N_1236,N_769);
and U2421 (N_2421,N_1521,N_1325);
and U2422 (N_2422,N_1454,N_14);
and U2423 (N_2423,N_1845,N_1838);
and U2424 (N_2424,N_1173,N_303);
or U2425 (N_2425,N_1656,N_1374);
or U2426 (N_2426,N_272,N_886);
nand U2427 (N_2427,N_1909,N_154);
nor U2428 (N_2428,N_1624,N_312);
and U2429 (N_2429,N_1167,N_1558);
nand U2430 (N_2430,N_1308,N_28);
nand U2431 (N_2431,N_1504,N_1622);
nor U2432 (N_2432,N_627,N_1667);
nand U2433 (N_2433,N_146,N_950);
and U2434 (N_2434,N_436,N_1153);
or U2435 (N_2435,N_795,N_633);
nor U2436 (N_2436,N_1468,N_1638);
or U2437 (N_2437,N_124,N_1388);
nand U2438 (N_2438,N_787,N_733);
nor U2439 (N_2439,N_686,N_1089);
or U2440 (N_2440,N_109,N_91);
or U2441 (N_2441,N_1551,N_1728);
nor U2442 (N_2442,N_505,N_1802);
nand U2443 (N_2443,N_1600,N_441);
and U2444 (N_2444,N_100,N_604);
nand U2445 (N_2445,N_1576,N_46);
or U2446 (N_2446,N_178,N_1854);
or U2447 (N_2447,N_322,N_625);
or U2448 (N_2448,N_116,N_416);
or U2449 (N_2449,N_937,N_1074);
nor U2450 (N_2450,N_1778,N_1165);
nor U2451 (N_2451,N_1001,N_430);
or U2452 (N_2452,N_1736,N_1117);
nand U2453 (N_2453,N_856,N_947);
nand U2454 (N_2454,N_335,N_32);
or U2455 (N_2455,N_1520,N_1896);
and U2456 (N_2456,N_1170,N_865);
nand U2457 (N_2457,N_631,N_746);
and U2458 (N_2458,N_1942,N_188);
nor U2459 (N_2459,N_1180,N_719);
nand U2460 (N_2460,N_648,N_1451);
or U2461 (N_2461,N_690,N_1582);
and U2462 (N_2462,N_1205,N_1899);
nor U2463 (N_2463,N_1113,N_400);
or U2464 (N_2464,N_1623,N_1943);
nand U2465 (N_2465,N_1011,N_1705);
or U2466 (N_2466,N_1517,N_939);
and U2467 (N_2467,N_366,N_518);
nor U2468 (N_2468,N_545,N_1832);
nor U2469 (N_2469,N_1032,N_1727);
nor U2470 (N_2470,N_1954,N_582);
and U2471 (N_2471,N_1793,N_159);
nand U2472 (N_2472,N_612,N_1072);
nor U2473 (N_2473,N_220,N_896);
nand U2474 (N_2474,N_1497,N_1111);
nand U2475 (N_2475,N_1413,N_819);
or U2476 (N_2476,N_4,N_1692);
nand U2477 (N_2477,N_1099,N_1039);
nor U2478 (N_2478,N_1874,N_391);
nor U2479 (N_2479,N_479,N_959);
nand U2480 (N_2480,N_1370,N_57);
or U2481 (N_2481,N_1398,N_1107);
nor U2482 (N_2482,N_345,N_905);
or U2483 (N_2483,N_748,N_697);
nand U2484 (N_2484,N_1330,N_477);
or U2485 (N_2485,N_183,N_1069);
nor U2486 (N_2486,N_635,N_1114);
nand U2487 (N_2487,N_135,N_1827);
or U2488 (N_2488,N_1801,N_78);
nand U2489 (N_2489,N_522,N_304);
or U2490 (N_2490,N_1038,N_1577);
nand U2491 (N_2491,N_128,N_1880);
xor U2492 (N_2492,N_1,N_793);
or U2493 (N_2493,N_1480,N_404);
and U2494 (N_2494,N_1256,N_901);
nand U2495 (N_2495,N_1544,N_243);
or U2496 (N_2496,N_1953,N_1258);
or U2497 (N_2497,N_546,N_509);
and U2498 (N_2498,N_655,N_1305);
nand U2499 (N_2499,N_1319,N_1820);
and U2500 (N_2500,N_1017,N_1620);
and U2501 (N_2501,N_1665,N_126);
nand U2502 (N_2502,N_125,N_529);
or U2503 (N_2503,N_1328,N_831);
and U2504 (N_2504,N_1912,N_761);
nor U2505 (N_2505,N_713,N_139);
or U2506 (N_2506,N_1493,N_548);
nor U2507 (N_2507,N_820,N_127);
nor U2508 (N_2508,N_778,N_1934);
nor U2509 (N_2509,N_1427,N_1369);
nand U2510 (N_2510,N_300,N_248);
or U2511 (N_2511,N_56,N_1049);
and U2512 (N_2512,N_888,N_276);
nor U2513 (N_2513,N_614,N_1724);
and U2514 (N_2514,N_1304,N_1387);
or U2515 (N_2515,N_996,N_1429);
or U2516 (N_2516,N_470,N_909);
nor U2517 (N_2517,N_35,N_1759);
and U2518 (N_2518,N_329,N_1533);
or U2519 (N_2519,N_1816,N_97);
and U2520 (N_2520,N_1564,N_554);
and U2521 (N_2521,N_1817,N_115);
nand U2522 (N_2522,N_192,N_1396);
xnor U2523 (N_2523,N_811,N_346);
or U2524 (N_2524,N_1657,N_501);
or U2525 (N_2525,N_253,N_1193);
and U2526 (N_2526,N_1530,N_1361);
nor U2527 (N_2527,N_801,N_1141);
and U2528 (N_2528,N_269,N_940);
xnor U2529 (N_2529,N_130,N_1410);
and U2530 (N_2530,N_817,N_1560);
or U2531 (N_2531,N_1704,N_288);
nor U2532 (N_2532,N_413,N_287);
nor U2533 (N_2533,N_514,N_478);
nand U2534 (N_2534,N_102,N_40);
nand U2535 (N_2535,N_1243,N_540);
nor U2536 (N_2536,N_1699,N_1982);
and U2537 (N_2537,N_114,N_840);
and U2538 (N_2538,N_790,N_1695);
and U2539 (N_2539,N_1763,N_450);
nand U2540 (N_2540,N_140,N_1283);
and U2541 (N_2541,N_1990,N_542);
and U2542 (N_2542,N_1848,N_402);
or U2543 (N_2543,N_1443,N_1713);
or U2544 (N_2544,N_1751,N_995);
or U2545 (N_2545,N_1650,N_1048);
and U2546 (N_2546,N_55,N_1187);
and U2547 (N_2547,N_1670,N_459);
nor U2548 (N_2548,N_1399,N_1207);
nor U2549 (N_2549,N_1718,N_662);
nor U2550 (N_2550,N_634,N_485);
and U2551 (N_2551,N_1204,N_1588);
or U2552 (N_2552,N_231,N_1198);
and U2553 (N_2553,N_1911,N_853);
xnor U2554 (N_2554,N_484,N_1569);
or U2555 (N_2555,N_1160,N_268);
xnor U2556 (N_2556,N_711,N_898);
or U2557 (N_2557,N_170,N_1733);
or U2558 (N_2558,N_1918,N_382);
or U2559 (N_2559,N_357,N_1133);
and U2560 (N_2560,N_1512,N_58);
nor U2561 (N_2561,N_1807,N_1231);
nand U2562 (N_2562,N_468,N_1586);
nor U2563 (N_2563,N_1602,N_1273);
nand U2564 (N_2564,N_695,N_1299);
or U2565 (N_2565,N_60,N_426);
nor U2566 (N_2566,N_328,N_314);
or U2567 (N_2567,N_1743,N_447);
or U2568 (N_2568,N_0,N_1262);
and U2569 (N_2569,N_731,N_261);
nor U2570 (N_2570,N_343,N_492);
and U2571 (N_2571,N_674,N_585);
and U2572 (N_2572,N_1277,N_437);
and U2573 (N_2573,N_1774,N_1864);
nor U2574 (N_2574,N_710,N_1865);
or U2575 (N_2575,N_804,N_1016);
or U2576 (N_2576,N_669,N_279);
and U2577 (N_2577,N_108,N_395);
and U2578 (N_2578,N_1717,N_1352);
or U2579 (N_2579,N_1353,N_1868);
or U2580 (N_2580,N_1752,N_24);
nor U2581 (N_2581,N_706,N_1406);
or U2582 (N_2582,N_1223,N_384);
or U2583 (N_2583,N_1343,N_549);
nand U2584 (N_2584,N_226,N_1613);
or U2585 (N_2585,N_1679,N_552);
and U2586 (N_2586,N_446,N_1358);
or U2587 (N_2587,N_594,N_1639);
or U2588 (N_2588,N_796,N_31);
or U2589 (N_2589,N_106,N_880);
nor U2590 (N_2590,N_603,N_1815);
nor U2591 (N_2591,N_1010,N_725);
and U2592 (N_2592,N_663,N_707);
or U2593 (N_2593,N_906,N_1991);
nor U2594 (N_2594,N_1400,N_1309);
or U2595 (N_2595,N_772,N_1542);
nor U2596 (N_2596,N_274,N_1298);
and U2597 (N_2597,N_563,N_412);
nand U2598 (N_2598,N_841,N_354);
or U2599 (N_2599,N_788,N_258);
nor U2600 (N_2600,N_132,N_1574);
and U2601 (N_2601,N_1442,N_681);
or U2602 (N_2602,N_457,N_260);
and U2603 (N_2603,N_859,N_1135);
or U2604 (N_2604,N_656,N_1097);
nor U2605 (N_2605,N_587,N_1221);
and U2606 (N_2606,N_605,N_1081);
or U2607 (N_2607,N_1962,N_791);
and U2608 (N_2608,N_1979,N_372);
or U2609 (N_2609,N_1022,N_214);
nor U2610 (N_2610,N_703,N_455);
and U2611 (N_2611,N_1448,N_36);
nor U2612 (N_2612,N_1961,N_676);
nand U2613 (N_2613,N_781,N_295);
or U2614 (N_2614,N_191,N_1035);
or U2615 (N_2615,N_1438,N_982);
or U2616 (N_2616,N_1471,N_890);
or U2617 (N_2617,N_868,N_432);
and U2618 (N_2618,N_1783,N_1785);
or U2619 (N_2619,N_979,N_541);
or U2620 (N_2620,N_110,N_1634);
nor U2621 (N_2621,N_72,N_500);
or U2622 (N_2622,N_1757,N_617);
nand U2623 (N_2623,N_371,N_816);
nand U2624 (N_2624,N_1818,N_511);
nor U2625 (N_2625,N_1554,N_891);
and U2626 (N_2626,N_1906,N_215);
and U2627 (N_2627,N_1522,N_390);
or U2628 (N_2628,N_1538,N_1447);
or U2629 (N_2629,N_18,N_1756);
or U2630 (N_2630,N_1327,N_1157);
or U2631 (N_2631,N_1885,N_629);
nor U2632 (N_2632,N_1466,N_1084);
nand U2633 (N_2633,N_608,N_683);
nand U2634 (N_2634,N_1106,N_1877);
nand U2635 (N_2635,N_773,N_1900);
nand U2636 (N_2636,N_1201,N_6);
and U2637 (N_2637,N_1825,N_628);
and U2638 (N_2638,N_1333,N_1746);
or U2639 (N_2639,N_1788,N_1279);
and U2640 (N_2640,N_153,N_600);
nand U2641 (N_2641,N_378,N_332);
nor U2642 (N_2642,N_495,N_1075);
nand U2643 (N_2643,N_361,N_325);
or U2644 (N_2644,N_1128,N_835);
nor U2645 (N_2645,N_1753,N_320);
or U2646 (N_2646,N_1598,N_1666);
nor U2647 (N_2647,N_196,N_1730);
nor U2648 (N_2648,N_1246,N_212);
or U2649 (N_2649,N_1796,N_622);
and U2650 (N_2650,N_851,N_1441);
and U2651 (N_2651,N_1213,N_957);
nor U2652 (N_2652,N_1203,N_553);
nor U2653 (N_2653,N_539,N_606);
or U2654 (N_2654,N_213,N_10);
and U2655 (N_2655,N_798,N_892);
nand U2656 (N_2656,N_487,N_1958);
or U2657 (N_2657,N_1871,N_1439);
nand U2658 (N_2658,N_152,N_1172);
and U2659 (N_2659,N_1552,N_69);
or U2660 (N_2660,N_1993,N_1156);
or U2661 (N_2661,N_538,N_1672);
and U2662 (N_2662,N_1249,N_240);
nor U2663 (N_2663,N_1336,N_620);
nor U2664 (N_2664,N_1515,N_1645);
nand U2665 (N_2665,N_843,N_1876);
and U2666 (N_2666,N_1245,N_740);
nand U2667 (N_2667,N_232,N_1729);
nor U2668 (N_2668,N_975,N_815);
nor U2669 (N_2669,N_879,N_565);
nand U2670 (N_2670,N_27,N_1232);
nor U2671 (N_2671,N_1571,N_1640);
or U2672 (N_2672,N_866,N_1118);
nor U2673 (N_2673,N_1130,N_427);
nor U2674 (N_2674,N_1710,N_749);
or U2675 (N_2675,N_1122,N_1740);
and U2676 (N_2676,N_1615,N_1014);
nor U2677 (N_2677,N_1469,N_630);
nand U2678 (N_2678,N_319,N_1659);
nand U2679 (N_2679,N_235,N_1619);
nor U2680 (N_2680,N_340,N_945);
or U2681 (N_2681,N_760,N_1453);
nor U2682 (N_2682,N_589,N_386);
or U2683 (N_2683,N_1580,N_1230);
and U2684 (N_2684,N_239,N_1259);
nand U2685 (N_2685,N_30,N_1483);
and U2686 (N_2686,N_1433,N_1534);
and U2687 (N_2687,N_1963,N_1261);
nand U2688 (N_2688,N_737,N_184);
and U2689 (N_2689,N_1492,N_1989);
nand U2690 (N_2690,N_331,N_536);
or U2691 (N_2691,N_87,N_1985);
or U2692 (N_2692,N_1087,N_1247);
nor U2693 (N_2693,N_289,N_23);
or U2694 (N_2694,N_1417,N_702);
nor U2695 (N_2695,N_1496,N_118);
and U2696 (N_2696,N_696,N_1371);
nand U2697 (N_2697,N_705,N_1415);
and U2698 (N_2698,N_1755,N_1179);
nor U2699 (N_2699,N_1897,N_1391);
nor U2700 (N_2700,N_7,N_1348);
or U2701 (N_2701,N_667,N_510);
nor U2702 (N_2702,N_263,N_611);
or U2703 (N_2703,N_229,N_1974);
nand U2704 (N_2704,N_1587,N_1392);
nor U2705 (N_2705,N_1844,N_1826);
and U2706 (N_2706,N_990,N_48);
nand U2707 (N_2707,N_203,N_1349);
and U2708 (N_2708,N_180,N_1585);
nand U2709 (N_2709,N_639,N_502);
nor U2710 (N_2710,N_1980,N_941);
or U2711 (N_2711,N_486,N_347);
or U2712 (N_2712,N_1322,N_291);
nor U2713 (N_2713,N_1381,N_167);
or U2714 (N_2714,N_65,N_1696);
nand U2715 (N_2715,N_1227,N_551);
nor U2716 (N_2716,N_96,N_1604);
nor U2717 (N_2717,N_770,N_1237);
or U2718 (N_2718,N_388,N_962);
nor U2719 (N_2719,N_640,N_961);
nand U2720 (N_2720,N_677,N_1166);
nor U2721 (N_2721,N_1605,N_1714);
nor U2722 (N_2722,N_1003,N_1196);
and U2723 (N_2723,N_708,N_1578);
nor U2724 (N_2724,N_358,N_1028);
nor U2725 (N_2725,N_535,N_1549);
nand U2726 (N_2726,N_1829,N_1103);
nor U2727 (N_2727,N_1567,N_186);
nand U2728 (N_2728,N_559,N_1494);
and U2729 (N_2729,N_924,N_491);
nand U2730 (N_2730,N_882,N_1952);
nand U2731 (N_2731,N_1481,N_445);
nor U2732 (N_2732,N_718,N_694);
or U2733 (N_2733,N_1476,N_575);
nand U2734 (N_2734,N_1631,N_1350);
and U2735 (N_2735,N_225,N_1384);
and U2736 (N_2736,N_607,N_1149);
nand U2737 (N_2737,N_742,N_1142);
nand U2738 (N_2738,N_1938,N_1320);
and U2739 (N_2739,N_1814,N_1267);
and U2740 (N_2740,N_904,N_1545);
and U2741 (N_2741,N_785,N_969);
and U2742 (N_2742,N_726,N_524);
nor U2743 (N_2743,N_285,N_1275);
and U2744 (N_2744,N_233,N_920);
and U2745 (N_2745,N_1781,N_394);
nand U2746 (N_2746,N_350,N_309);
or U2747 (N_2747,N_1532,N_1553);
nand U2748 (N_2748,N_1568,N_463);
nand U2749 (N_2749,N_1354,N_1747);
nand U2750 (N_2750,N_1907,N_1593);
or U2751 (N_2751,N_1234,N_1891);
nor U2752 (N_2752,N_1036,N_1949);
nand U2753 (N_2753,N_574,N_780);
or U2754 (N_2754,N_972,N_419);
and U2755 (N_2755,N_1229,N_1285);
and U2756 (N_2756,N_850,N_1186);
nand U2757 (N_2757,N_568,N_1216);
nor U2758 (N_2758,N_1901,N_462);
and U2759 (N_2759,N_1096,N_1678);
and U2760 (N_2760,N_1119,N_921);
nor U2761 (N_2761,N_88,N_613);
and U2762 (N_2762,N_483,N_204);
and U2763 (N_2763,N_1423,N_944);
and U2764 (N_2764,N_1787,N_1987);
nand U2765 (N_2765,N_1375,N_1482);
or U2766 (N_2766,N_1394,N_1108);
nand U2767 (N_2767,N_1646,N_1104);
or U2768 (N_2768,N_1948,N_1051);
and U2769 (N_2769,N_1537,N_922);
nor U2770 (N_2770,N_601,N_408);
or U2771 (N_2771,N_894,N_1648);
and U2772 (N_2772,N_987,N_85);
and U2773 (N_2773,N_858,N_907);
xor U2774 (N_2774,N_83,N_1123);
or U2775 (N_2775,N_1526,N_1209);
nor U2776 (N_2776,N_963,N_458);
and U2777 (N_2777,N_508,N_1345);
nand U2778 (N_2778,N_985,N_1422);
xnor U2779 (N_2779,N_747,N_809);
or U2780 (N_2780,N_1959,N_1405);
nand U2781 (N_2781,N_624,N_1823);
and U2782 (N_2782,N_799,N_1973);
and U2783 (N_2783,N_682,N_218);
nor U2784 (N_2784,N_448,N_1536);
and U2785 (N_2785,N_369,N_1313);
or U2786 (N_2786,N_534,N_599);
nand U2787 (N_2787,N_1888,N_471);
nor U2788 (N_2788,N_1725,N_389);
nor U2789 (N_2789,N_1539,N_825);
nor U2790 (N_2790,N_247,N_557);
or U2791 (N_2791,N_1509,N_1506);
and U2792 (N_2792,N_497,N_986);
and U2793 (N_2793,N_1284,N_112);
or U2794 (N_2794,N_1002,N_1734);
xor U2795 (N_2795,N_1649,N_190);
nor U2796 (N_2796,N_1382,N_821);
nand U2797 (N_2797,N_66,N_877);
nand U2798 (N_2798,N_67,N_1436);
nand U2799 (N_2799,N_443,N_1054);
and U2800 (N_2800,N_16,N_912);
and U2801 (N_2801,N_1218,N_660);
nor U2802 (N_2802,N_806,N_1040);
and U2803 (N_2803,N_507,N_101);
nor U2804 (N_2804,N_1324,N_353);
nor U2805 (N_2805,N_1000,N_280);
nor U2806 (N_2806,N_1290,N_875);
nand U2807 (N_2807,N_2,N_857);
xnor U2808 (N_2808,N_1933,N_1479);
and U2809 (N_2809,N_1726,N_1169);
and U2810 (N_2810,N_1251,N_1945);
nand U2811 (N_2811,N_1491,N_238);
nor U2812 (N_2812,N_525,N_119);
nor U2813 (N_2813,N_1363,N_1830);
nand U2814 (N_2814,N_1835,N_73);
nor U2815 (N_2815,N_543,N_172);
or U2816 (N_2816,N_530,N_899);
and U2817 (N_2817,N_980,N_1673);
and U2818 (N_2818,N_913,N_1735);
nand U2819 (N_2819,N_1158,N_1641);
nand U2820 (N_2820,N_666,N_1109);
and U2821 (N_2821,N_1340,N_349);
nor U2822 (N_2822,N_95,N_929);
nand U2823 (N_2823,N_672,N_1018);
nand U2824 (N_2824,N_1931,N_177);
and U2825 (N_2825,N_1431,N_311);
and U2826 (N_2826,N_721,N_670);
nor U2827 (N_2827,N_504,N_207);
or U2828 (N_2828,N_1235,N_9);
nor U2829 (N_2829,N_370,N_654);
nand U2830 (N_2830,N_1798,N_1772);
or U2831 (N_2831,N_1463,N_1760);
nand U2832 (N_2832,N_596,N_874);
nor U2833 (N_2833,N_1519,N_1684);
and U2834 (N_2834,N_908,N_602);
and U2835 (N_2835,N_1465,N_1339);
or U2836 (N_2836,N_918,N_1037);
nor U2837 (N_2837,N_776,N_1455);
nand U2838 (N_2838,N_836,N_1444);
nand U2839 (N_2839,N_498,N_1012);
or U2840 (N_2840,N_363,N_823);
and U2841 (N_2841,N_136,N_398);
or U2842 (N_2842,N_1472,N_193);
nor U2843 (N_2843,N_75,N_1052);
nor U2844 (N_2844,N_219,N_1914);
nor U2845 (N_2845,N_569,N_374);
nand U2846 (N_2846,N_1331,N_1786);
and U2847 (N_2847,N_1095,N_1314);
or U2848 (N_2848,N_1124,N_1978);
and U2849 (N_2849,N_141,N_966);
or U2850 (N_2850,N_1435,N_1846);
or U2851 (N_2851,N_409,N_989);
and U2852 (N_2852,N_591,N_1202);
and U2853 (N_2853,N_1024,N_107);
nor U2854 (N_2854,N_926,N_1603);
nor U2855 (N_2855,N_80,N_1702);
xnor U2856 (N_2856,N_641,N_1395);
nand U2857 (N_2857,N_936,N_572);
nand U2858 (N_2858,N_902,N_1177);
or U2859 (N_2859,N_1326,N_1698);
and U2860 (N_2860,N_1362,N_597);
or U2861 (N_2861,N_1633,N_286);
nor U2862 (N_2862,N_813,N_317);
and U2863 (N_2863,N_1810,N_846);
nor U2864 (N_2864,N_637,N_673);
nand U2865 (N_2865,N_1926,N_1219);
or U2866 (N_2866,N_1185,N_1563);
or U2867 (N_2867,N_910,N_451);
and U2868 (N_2868,N_148,N_794);
nor U2869 (N_2869,N_1721,N_783);
and U2870 (N_2870,N_893,N_1572);
or U2871 (N_2871,N_1741,N_610);
and U2872 (N_2872,N_738,N_405);
nand U2873 (N_2873,N_1643,N_1841);
nand U2874 (N_2874,N_21,N_195);
or U2875 (N_2875,N_1946,N_438);
nand U2876 (N_2876,N_1253,N_76);
and U2877 (N_2877,N_1606,N_1937);
or U2878 (N_2878,N_645,N_1669);
or U2879 (N_2879,N_473,N_489);
nand U2880 (N_2880,N_1121,N_20);
xnor U2881 (N_2881,N_1677,N_1694);
or U2882 (N_2882,N_897,N_727);
and U2883 (N_2883,N_1407,N_871);
and U2884 (N_2884,N_1922,N_1703);
or U2885 (N_2885,N_1004,N_62);
and U2886 (N_2886,N_493,N_774);
nor U2887 (N_2887,N_1034,N_626);
or U2888 (N_2888,N_1916,N_643);
nor U2889 (N_2889,N_1424,N_1930);
or U2890 (N_2890,N_1214,N_1163);
and U2891 (N_2891,N_1610,N_296);
or U2892 (N_2892,N_1663,N_1263);
and U2893 (N_2893,N_1658,N_1790);
or U2894 (N_2894,N_1686,N_595);
and U2895 (N_2895,N_1462,N_1951);
nand U2896 (N_2896,N_847,N_173);
and U2897 (N_2897,N_169,N_970);
nand U2898 (N_2898,N_452,N_284);
nor U2899 (N_2899,N_1866,N_1293);
or U2900 (N_2900,N_418,N_1367);
nand U2901 (N_2901,N_1617,N_387);
nor U2902 (N_2902,N_827,N_1921);
or U2903 (N_2903,N_1120,N_222);
and U2904 (N_2904,N_579,N_736);
nor U2905 (N_2905,N_1047,N_724);
nand U2906 (N_2906,N_38,N_1632);
nor U2907 (N_2907,N_8,N_131);
and U2908 (N_2908,N_1007,N_971);
nor U2909 (N_2909,N_1988,N_1154);
or U2910 (N_2910,N_1715,N_1524);
nand U2911 (N_2911,N_786,N_1965);
nand U2912 (N_2912,N_399,N_1511);
nor U2913 (N_2913,N_878,N_1226);
nor U2914 (N_2914,N_337,N_422);
nand U2915 (N_2915,N_993,N_444);
nor U2916 (N_2916,N_714,N_1178);
or U2917 (N_2917,N_869,N_1583);
nor U2918 (N_2918,N_1685,N_657);
or U2919 (N_2919,N_1859,N_862);
and U2920 (N_2920,N_1164,N_1378);
nor U2921 (N_2921,N_1094,N_1068);
and U2922 (N_2922,N_355,N_63);
and U2923 (N_2923,N_1828,N_928);
nand U2924 (N_2924,N_779,N_265);
nand U2925 (N_2925,N_954,N_1960);
nand U2926 (N_2926,N_1856,N_39);
or U2927 (N_2927,N_442,N_722);
nor U2928 (N_2928,N_1626,N_1611);
nor U2929 (N_2929,N_1224,N_973);
nand U2930 (N_2930,N_1546,N_923);
or U2931 (N_2931,N_373,N_1300);
and U2932 (N_2932,N_573,N_1867);
or U2933 (N_2933,N_79,N_704);
nand U2934 (N_2934,N_1368,N_1732);
nor U2935 (N_2935,N_359,N_105);
and U2936 (N_2936,N_644,N_1738);
or U2937 (N_2937,N_984,N_1629);
nand U2938 (N_2938,N_1701,N_544);
or U2939 (N_2939,N_1903,N_344);
or U2940 (N_2940,N_1220,N_1420);
nand U2941 (N_2941,N_1357,N_1467);
nor U2942 (N_2942,N_1765,N_732);
or U2943 (N_2943,N_948,N_1709);
nor U2944 (N_2944,N_943,N_701);
nor U2945 (N_2945,N_1306,N_842);
nor U2946 (N_2946,N_348,N_1092);
and U2947 (N_2947,N_1401,N_965);
nand U2948 (N_2948,N_1145,N_860);
or U2949 (N_2949,N_828,N_547);
or U2950 (N_2950,N_915,N_1377);
nor U2951 (N_2951,N_1148,N_766);
nor U2952 (N_2952,N_739,N_1461);
nand U2953 (N_2953,N_1767,N_1181);
nor U2954 (N_2954,N_1591,N_566);
and U2955 (N_2955,N_976,N_949);
or U2956 (N_2956,N_1840,N_292);
nor U2957 (N_2957,N_646,N_1618);
or U2958 (N_2958,N_410,N_698);
and U2959 (N_2959,N_333,N_1412);
and U2960 (N_2960,N_1257,N_1356);
and U2961 (N_2961,N_807,N_844);
nand U2962 (N_2962,N_236,N_482);
nand U2963 (N_2963,N_1321,N_988);
nand U2964 (N_2964,N_503,N_931);
nand U2965 (N_2965,N_555,N_994);
nor U2966 (N_2966,N_1742,N_1927);
nor U2967 (N_2967,N_1540,N_876);
or U2968 (N_2968,N_142,N_765);
and U2969 (N_2969,N_1662,N_499);
or U2970 (N_2970,N_1998,N_516);
and U2971 (N_2971,N_1297,N_1062);
nor U2972 (N_2972,N_200,N_687);
or U2973 (N_2973,N_92,N_1739);
and U2974 (N_2974,N_466,N_1489);
or U2975 (N_2975,N_1091,N_1144);
nor U2976 (N_2976,N_1655,N_326);
nand U2977 (N_2977,N_1446,N_1200);
or U2978 (N_2978,N_1744,N_1852);
nor U2979 (N_2979,N_1291,N_1777);
or U2980 (N_2980,N_251,N_1886);
nand U2981 (N_2981,N_185,N_1936);
nand U2982 (N_2982,N_883,N_1380);
nand U2983 (N_2983,N_1566,N_757);
or U2984 (N_2984,N_1935,N_1881);
nand U2985 (N_2985,N_803,N_1064);
nand U2986 (N_2986,N_256,N_1402);
nor U2987 (N_2987,N_1029,N_1707);
or U2988 (N_2988,N_294,N_675);
nor U2989 (N_2989,N_1194,N_946);
or U2990 (N_2990,N_392,N_327);
or U2991 (N_2991,N_978,N_150);
and U2992 (N_2992,N_955,N_1495);
or U2993 (N_2993,N_481,N_1138);
and U2994 (N_2994,N_526,N_917);
nor U2995 (N_2995,N_1310,N_1210);
nor U2996 (N_2996,N_968,N_752);
or U2997 (N_2997,N_1575,N_903);
nor U2998 (N_2998,N_750,N_1723);
nand U2999 (N_2999,N_1080,N_1093);
nand U3000 (N_3000,N_651,N_458);
and U3001 (N_3001,N_1492,N_1594);
nand U3002 (N_3002,N_1040,N_289);
or U3003 (N_3003,N_401,N_75);
nand U3004 (N_3004,N_1919,N_595);
nor U3005 (N_3005,N_828,N_183);
and U3006 (N_3006,N_1710,N_1452);
nor U3007 (N_3007,N_1242,N_1032);
and U3008 (N_3008,N_1881,N_979);
nor U3009 (N_3009,N_1674,N_1673);
nor U3010 (N_3010,N_1675,N_680);
nor U3011 (N_3011,N_1710,N_1613);
and U3012 (N_3012,N_253,N_1029);
xor U3013 (N_3013,N_1305,N_1148);
and U3014 (N_3014,N_934,N_1378);
nand U3015 (N_3015,N_1709,N_306);
or U3016 (N_3016,N_1464,N_269);
and U3017 (N_3017,N_876,N_1146);
nand U3018 (N_3018,N_732,N_148);
and U3019 (N_3019,N_1166,N_41);
nor U3020 (N_3020,N_1936,N_1289);
nor U3021 (N_3021,N_313,N_1012);
or U3022 (N_3022,N_693,N_350);
nor U3023 (N_3023,N_1700,N_1764);
or U3024 (N_3024,N_788,N_884);
nand U3025 (N_3025,N_1628,N_1839);
nand U3026 (N_3026,N_1418,N_820);
and U3027 (N_3027,N_1122,N_1383);
nor U3028 (N_3028,N_640,N_1224);
nand U3029 (N_3029,N_1195,N_543);
or U3030 (N_3030,N_652,N_1752);
nand U3031 (N_3031,N_218,N_1482);
and U3032 (N_3032,N_276,N_1037);
nand U3033 (N_3033,N_1101,N_1739);
nand U3034 (N_3034,N_613,N_898);
or U3035 (N_3035,N_207,N_451);
or U3036 (N_3036,N_1008,N_1948);
nor U3037 (N_3037,N_1254,N_846);
or U3038 (N_3038,N_1811,N_1071);
or U3039 (N_3039,N_381,N_1544);
nand U3040 (N_3040,N_737,N_51);
or U3041 (N_3041,N_1748,N_1192);
nand U3042 (N_3042,N_692,N_1292);
nand U3043 (N_3043,N_1889,N_205);
nor U3044 (N_3044,N_922,N_1524);
and U3045 (N_3045,N_325,N_1938);
or U3046 (N_3046,N_697,N_1450);
nand U3047 (N_3047,N_1263,N_129);
nand U3048 (N_3048,N_669,N_885);
and U3049 (N_3049,N_1765,N_1316);
nor U3050 (N_3050,N_1376,N_442);
nor U3051 (N_3051,N_866,N_1856);
nand U3052 (N_3052,N_238,N_137);
and U3053 (N_3053,N_511,N_594);
or U3054 (N_3054,N_1459,N_277);
or U3055 (N_3055,N_354,N_267);
nand U3056 (N_3056,N_1429,N_1482);
nor U3057 (N_3057,N_145,N_38);
xnor U3058 (N_3058,N_200,N_925);
and U3059 (N_3059,N_161,N_1730);
nor U3060 (N_3060,N_643,N_1558);
and U3061 (N_3061,N_19,N_177);
or U3062 (N_3062,N_520,N_673);
and U3063 (N_3063,N_1364,N_758);
or U3064 (N_3064,N_1828,N_1362);
nor U3065 (N_3065,N_1707,N_1145);
and U3066 (N_3066,N_1135,N_1175);
and U3067 (N_3067,N_1717,N_856);
and U3068 (N_3068,N_727,N_528);
or U3069 (N_3069,N_1614,N_802);
nand U3070 (N_3070,N_1148,N_1545);
nor U3071 (N_3071,N_1802,N_576);
or U3072 (N_3072,N_1888,N_1303);
or U3073 (N_3073,N_819,N_1057);
or U3074 (N_3074,N_1462,N_584);
and U3075 (N_3075,N_1017,N_303);
or U3076 (N_3076,N_698,N_17);
nand U3077 (N_3077,N_1708,N_866);
or U3078 (N_3078,N_1033,N_1769);
and U3079 (N_3079,N_1534,N_386);
nand U3080 (N_3080,N_358,N_1004);
nand U3081 (N_3081,N_1744,N_1630);
nor U3082 (N_3082,N_550,N_1613);
nand U3083 (N_3083,N_1663,N_853);
and U3084 (N_3084,N_1577,N_508);
nor U3085 (N_3085,N_420,N_1212);
and U3086 (N_3086,N_916,N_1970);
nand U3087 (N_3087,N_841,N_571);
nand U3088 (N_3088,N_265,N_1915);
or U3089 (N_3089,N_1802,N_1029);
and U3090 (N_3090,N_1643,N_912);
or U3091 (N_3091,N_1104,N_1729);
nand U3092 (N_3092,N_523,N_1982);
or U3093 (N_3093,N_1422,N_1971);
nor U3094 (N_3094,N_409,N_892);
nand U3095 (N_3095,N_1451,N_1358);
nand U3096 (N_3096,N_141,N_1835);
nand U3097 (N_3097,N_1243,N_894);
nor U3098 (N_3098,N_1663,N_1835);
nor U3099 (N_3099,N_273,N_932);
nor U3100 (N_3100,N_74,N_773);
nand U3101 (N_3101,N_744,N_827);
nand U3102 (N_3102,N_1609,N_1655);
and U3103 (N_3103,N_738,N_1051);
nor U3104 (N_3104,N_1509,N_1487);
and U3105 (N_3105,N_1555,N_613);
or U3106 (N_3106,N_346,N_1705);
and U3107 (N_3107,N_1453,N_1839);
or U3108 (N_3108,N_339,N_592);
nor U3109 (N_3109,N_1536,N_65);
nor U3110 (N_3110,N_360,N_1751);
and U3111 (N_3111,N_933,N_1586);
or U3112 (N_3112,N_1831,N_1478);
nor U3113 (N_3113,N_638,N_1094);
and U3114 (N_3114,N_1590,N_220);
nor U3115 (N_3115,N_973,N_1632);
nand U3116 (N_3116,N_499,N_1407);
xor U3117 (N_3117,N_1088,N_1038);
xor U3118 (N_3118,N_1850,N_1409);
and U3119 (N_3119,N_1007,N_1351);
nand U3120 (N_3120,N_1911,N_1730);
and U3121 (N_3121,N_1329,N_972);
and U3122 (N_3122,N_1761,N_238);
nor U3123 (N_3123,N_1669,N_120);
nand U3124 (N_3124,N_1632,N_333);
nor U3125 (N_3125,N_475,N_1457);
nor U3126 (N_3126,N_327,N_290);
and U3127 (N_3127,N_904,N_349);
nor U3128 (N_3128,N_19,N_1146);
and U3129 (N_3129,N_1190,N_451);
nand U3130 (N_3130,N_1402,N_1287);
nor U3131 (N_3131,N_1001,N_1739);
nand U3132 (N_3132,N_441,N_271);
nand U3133 (N_3133,N_1633,N_1477);
and U3134 (N_3134,N_809,N_1195);
nor U3135 (N_3135,N_1486,N_1613);
and U3136 (N_3136,N_1622,N_682);
nor U3137 (N_3137,N_1412,N_325);
or U3138 (N_3138,N_1350,N_375);
and U3139 (N_3139,N_1158,N_180);
nand U3140 (N_3140,N_214,N_1825);
nand U3141 (N_3141,N_1241,N_97);
nand U3142 (N_3142,N_1013,N_1763);
xnor U3143 (N_3143,N_866,N_1490);
and U3144 (N_3144,N_1157,N_189);
or U3145 (N_3145,N_1526,N_1129);
nand U3146 (N_3146,N_1696,N_1024);
or U3147 (N_3147,N_24,N_172);
and U3148 (N_3148,N_623,N_846);
and U3149 (N_3149,N_957,N_1796);
nor U3150 (N_3150,N_1417,N_91);
nand U3151 (N_3151,N_1489,N_935);
nor U3152 (N_3152,N_1674,N_970);
or U3153 (N_3153,N_66,N_899);
xor U3154 (N_3154,N_1138,N_948);
nor U3155 (N_3155,N_568,N_624);
and U3156 (N_3156,N_1831,N_663);
and U3157 (N_3157,N_996,N_1198);
nor U3158 (N_3158,N_1579,N_52);
and U3159 (N_3159,N_570,N_974);
and U3160 (N_3160,N_870,N_1103);
nand U3161 (N_3161,N_1898,N_1978);
nand U3162 (N_3162,N_486,N_1933);
and U3163 (N_3163,N_811,N_1940);
nand U3164 (N_3164,N_1485,N_1001);
or U3165 (N_3165,N_394,N_1286);
nand U3166 (N_3166,N_1839,N_1143);
nand U3167 (N_3167,N_232,N_295);
nor U3168 (N_3168,N_1036,N_1156);
nand U3169 (N_3169,N_1857,N_607);
or U3170 (N_3170,N_100,N_764);
or U3171 (N_3171,N_447,N_62);
and U3172 (N_3172,N_1063,N_713);
nor U3173 (N_3173,N_128,N_1101);
and U3174 (N_3174,N_9,N_1977);
nor U3175 (N_3175,N_1010,N_1155);
and U3176 (N_3176,N_187,N_1306);
nor U3177 (N_3177,N_708,N_1066);
or U3178 (N_3178,N_1697,N_983);
and U3179 (N_3179,N_1922,N_507);
or U3180 (N_3180,N_1905,N_1113);
nand U3181 (N_3181,N_1298,N_1212);
nand U3182 (N_3182,N_1285,N_1959);
or U3183 (N_3183,N_1155,N_1462);
nand U3184 (N_3184,N_1888,N_257);
or U3185 (N_3185,N_448,N_1613);
nand U3186 (N_3186,N_1699,N_1404);
nor U3187 (N_3187,N_765,N_1104);
nor U3188 (N_3188,N_116,N_1132);
nor U3189 (N_3189,N_330,N_511);
nor U3190 (N_3190,N_1318,N_970);
nor U3191 (N_3191,N_77,N_1638);
nor U3192 (N_3192,N_727,N_1363);
and U3193 (N_3193,N_1194,N_1275);
and U3194 (N_3194,N_1276,N_1598);
and U3195 (N_3195,N_1989,N_1812);
nand U3196 (N_3196,N_1488,N_546);
nand U3197 (N_3197,N_1287,N_1708);
or U3198 (N_3198,N_1355,N_931);
and U3199 (N_3199,N_1157,N_1723);
nor U3200 (N_3200,N_496,N_88);
nor U3201 (N_3201,N_657,N_313);
and U3202 (N_3202,N_1593,N_1966);
nand U3203 (N_3203,N_159,N_387);
and U3204 (N_3204,N_1023,N_282);
or U3205 (N_3205,N_1849,N_1691);
nand U3206 (N_3206,N_681,N_44);
and U3207 (N_3207,N_1166,N_369);
and U3208 (N_3208,N_1588,N_1199);
nand U3209 (N_3209,N_1377,N_422);
nand U3210 (N_3210,N_840,N_712);
or U3211 (N_3211,N_302,N_306);
and U3212 (N_3212,N_1720,N_676);
and U3213 (N_3213,N_1699,N_1094);
and U3214 (N_3214,N_306,N_1625);
and U3215 (N_3215,N_908,N_1403);
and U3216 (N_3216,N_309,N_591);
nor U3217 (N_3217,N_206,N_1171);
nand U3218 (N_3218,N_367,N_235);
nor U3219 (N_3219,N_644,N_1576);
nor U3220 (N_3220,N_96,N_830);
and U3221 (N_3221,N_101,N_18);
nor U3222 (N_3222,N_1452,N_1307);
nand U3223 (N_3223,N_1118,N_1853);
nor U3224 (N_3224,N_515,N_513);
and U3225 (N_3225,N_531,N_1659);
nor U3226 (N_3226,N_1408,N_700);
and U3227 (N_3227,N_977,N_747);
and U3228 (N_3228,N_242,N_1218);
nor U3229 (N_3229,N_592,N_1391);
and U3230 (N_3230,N_744,N_761);
nor U3231 (N_3231,N_663,N_1315);
nor U3232 (N_3232,N_1858,N_1840);
nor U3233 (N_3233,N_168,N_1098);
and U3234 (N_3234,N_896,N_558);
and U3235 (N_3235,N_307,N_692);
nand U3236 (N_3236,N_1439,N_851);
nor U3237 (N_3237,N_1178,N_1331);
nor U3238 (N_3238,N_972,N_1753);
and U3239 (N_3239,N_1973,N_959);
nor U3240 (N_3240,N_1952,N_1128);
nor U3241 (N_3241,N_1465,N_1249);
nor U3242 (N_3242,N_1522,N_1552);
nor U3243 (N_3243,N_1280,N_658);
and U3244 (N_3244,N_384,N_1865);
nand U3245 (N_3245,N_1466,N_636);
or U3246 (N_3246,N_1396,N_1172);
nand U3247 (N_3247,N_1051,N_1377);
and U3248 (N_3248,N_1178,N_476);
nand U3249 (N_3249,N_320,N_875);
or U3250 (N_3250,N_1204,N_1378);
nand U3251 (N_3251,N_1679,N_1349);
nor U3252 (N_3252,N_1745,N_33);
nand U3253 (N_3253,N_1957,N_1447);
or U3254 (N_3254,N_1189,N_1370);
or U3255 (N_3255,N_1158,N_522);
or U3256 (N_3256,N_1104,N_1808);
and U3257 (N_3257,N_740,N_552);
nand U3258 (N_3258,N_1835,N_1487);
and U3259 (N_3259,N_1536,N_1855);
or U3260 (N_3260,N_124,N_1014);
nand U3261 (N_3261,N_103,N_1782);
nor U3262 (N_3262,N_1090,N_185);
nor U3263 (N_3263,N_151,N_1482);
or U3264 (N_3264,N_1326,N_1164);
nand U3265 (N_3265,N_335,N_815);
and U3266 (N_3266,N_1133,N_1522);
and U3267 (N_3267,N_1537,N_1495);
and U3268 (N_3268,N_1382,N_1271);
and U3269 (N_3269,N_893,N_1009);
and U3270 (N_3270,N_911,N_970);
nor U3271 (N_3271,N_1015,N_170);
nor U3272 (N_3272,N_1516,N_683);
or U3273 (N_3273,N_1656,N_1645);
nand U3274 (N_3274,N_1641,N_1822);
and U3275 (N_3275,N_414,N_1126);
and U3276 (N_3276,N_1225,N_34);
or U3277 (N_3277,N_281,N_82);
nand U3278 (N_3278,N_735,N_1836);
nand U3279 (N_3279,N_1639,N_949);
xnor U3280 (N_3280,N_789,N_86);
and U3281 (N_3281,N_379,N_781);
or U3282 (N_3282,N_1635,N_754);
or U3283 (N_3283,N_1813,N_1116);
nor U3284 (N_3284,N_202,N_1527);
nor U3285 (N_3285,N_1249,N_81);
xor U3286 (N_3286,N_409,N_883);
and U3287 (N_3287,N_889,N_606);
and U3288 (N_3288,N_1180,N_1983);
or U3289 (N_3289,N_1289,N_14);
and U3290 (N_3290,N_1761,N_100);
and U3291 (N_3291,N_289,N_1125);
and U3292 (N_3292,N_1117,N_551);
or U3293 (N_3293,N_302,N_645);
or U3294 (N_3294,N_1839,N_1793);
nor U3295 (N_3295,N_1340,N_779);
nand U3296 (N_3296,N_1762,N_813);
nand U3297 (N_3297,N_636,N_84);
or U3298 (N_3298,N_1437,N_113);
and U3299 (N_3299,N_546,N_395);
or U3300 (N_3300,N_1672,N_706);
or U3301 (N_3301,N_364,N_1769);
or U3302 (N_3302,N_314,N_36);
nor U3303 (N_3303,N_356,N_1234);
nor U3304 (N_3304,N_1233,N_188);
or U3305 (N_3305,N_262,N_756);
nand U3306 (N_3306,N_1951,N_346);
and U3307 (N_3307,N_452,N_1864);
and U3308 (N_3308,N_238,N_1083);
and U3309 (N_3309,N_191,N_487);
and U3310 (N_3310,N_570,N_1645);
and U3311 (N_3311,N_11,N_905);
nand U3312 (N_3312,N_317,N_658);
nand U3313 (N_3313,N_619,N_882);
and U3314 (N_3314,N_1603,N_121);
nand U3315 (N_3315,N_86,N_1609);
nand U3316 (N_3316,N_731,N_1647);
or U3317 (N_3317,N_15,N_1440);
nor U3318 (N_3318,N_96,N_786);
and U3319 (N_3319,N_1081,N_1380);
and U3320 (N_3320,N_1486,N_744);
nand U3321 (N_3321,N_1137,N_1432);
and U3322 (N_3322,N_404,N_307);
nor U3323 (N_3323,N_224,N_1418);
nor U3324 (N_3324,N_1440,N_1743);
and U3325 (N_3325,N_1064,N_504);
nor U3326 (N_3326,N_118,N_271);
or U3327 (N_3327,N_347,N_1730);
nand U3328 (N_3328,N_735,N_640);
nand U3329 (N_3329,N_1831,N_132);
nor U3330 (N_3330,N_622,N_1390);
and U3331 (N_3331,N_592,N_1233);
and U3332 (N_3332,N_389,N_1474);
nor U3333 (N_3333,N_950,N_316);
or U3334 (N_3334,N_1598,N_169);
xor U3335 (N_3335,N_1867,N_1766);
or U3336 (N_3336,N_462,N_1241);
nand U3337 (N_3337,N_697,N_660);
and U3338 (N_3338,N_1834,N_955);
nand U3339 (N_3339,N_208,N_1867);
or U3340 (N_3340,N_1308,N_119);
nand U3341 (N_3341,N_1037,N_1618);
nand U3342 (N_3342,N_61,N_1379);
and U3343 (N_3343,N_287,N_1651);
nand U3344 (N_3344,N_1658,N_1532);
nor U3345 (N_3345,N_1414,N_739);
and U3346 (N_3346,N_1145,N_713);
or U3347 (N_3347,N_310,N_233);
and U3348 (N_3348,N_512,N_109);
and U3349 (N_3349,N_1618,N_798);
and U3350 (N_3350,N_784,N_1811);
and U3351 (N_3351,N_270,N_119);
nand U3352 (N_3352,N_389,N_1463);
or U3353 (N_3353,N_1782,N_1563);
nor U3354 (N_3354,N_382,N_1497);
xor U3355 (N_3355,N_1239,N_921);
or U3356 (N_3356,N_1748,N_1193);
or U3357 (N_3357,N_227,N_1886);
nor U3358 (N_3358,N_913,N_384);
and U3359 (N_3359,N_1610,N_884);
nand U3360 (N_3360,N_991,N_796);
nand U3361 (N_3361,N_129,N_945);
nor U3362 (N_3362,N_572,N_1742);
and U3363 (N_3363,N_197,N_1678);
or U3364 (N_3364,N_549,N_1199);
and U3365 (N_3365,N_171,N_1729);
and U3366 (N_3366,N_1181,N_952);
nor U3367 (N_3367,N_1369,N_1150);
or U3368 (N_3368,N_1450,N_1253);
or U3369 (N_3369,N_541,N_218);
and U3370 (N_3370,N_516,N_1178);
nand U3371 (N_3371,N_1819,N_1659);
or U3372 (N_3372,N_356,N_270);
or U3373 (N_3373,N_877,N_204);
xnor U3374 (N_3374,N_1975,N_313);
nand U3375 (N_3375,N_1320,N_1746);
nand U3376 (N_3376,N_1081,N_1763);
nor U3377 (N_3377,N_1231,N_512);
or U3378 (N_3378,N_1459,N_561);
and U3379 (N_3379,N_847,N_1500);
nor U3380 (N_3380,N_1282,N_1013);
nand U3381 (N_3381,N_1500,N_1185);
or U3382 (N_3382,N_1420,N_1216);
nor U3383 (N_3383,N_707,N_1517);
and U3384 (N_3384,N_36,N_1463);
or U3385 (N_3385,N_346,N_873);
and U3386 (N_3386,N_1583,N_216);
and U3387 (N_3387,N_1495,N_191);
and U3388 (N_3388,N_663,N_1284);
nor U3389 (N_3389,N_1222,N_293);
nor U3390 (N_3390,N_605,N_1147);
or U3391 (N_3391,N_606,N_1845);
and U3392 (N_3392,N_441,N_689);
and U3393 (N_3393,N_1958,N_333);
nand U3394 (N_3394,N_1364,N_939);
and U3395 (N_3395,N_1408,N_18);
or U3396 (N_3396,N_1365,N_1119);
nor U3397 (N_3397,N_1999,N_505);
nand U3398 (N_3398,N_1352,N_235);
or U3399 (N_3399,N_368,N_60);
and U3400 (N_3400,N_800,N_1);
or U3401 (N_3401,N_1982,N_136);
and U3402 (N_3402,N_1292,N_776);
nand U3403 (N_3403,N_1412,N_867);
and U3404 (N_3404,N_1718,N_684);
or U3405 (N_3405,N_512,N_824);
and U3406 (N_3406,N_613,N_1161);
or U3407 (N_3407,N_413,N_1359);
and U3408 (N_3408,N_1460,N_350);
or U3409 (N_3409,N_1150,N_672);
nor U3410 (N_3410,N_543,N_597);
nor U3411 (N_3411,N_684,N_988);
nand U3412 (N_3412,N_226,N_1694);
and U3413 (N_3413,N_1476,N_1665);
or U3414 (N_3414,N_1972,N_1131);
nor U3415 (N_3415,N_1945,N_606);
and U3416 (N_3416,N_1731,N_711);
nor U3417 (N_3417,N_588,N_432);
nand U3418 (N_3418,N_1513,N_1270);
nor U3419 (N_3419,N_311,N_1);
and U3420 (N_3420,N_312,N_8);
nor U3421 (N_3421,N_810,N_1559);
nand U3422 (N_3422,N_519,N_1152);
nand U3423 (N_3423,N_1928,N_1591);
nor U3424 (N_3424,N_1581,N_1281);
nor U3425 (N_3425,N_720,N_1368);
or U3426 (N_3426,N_1552,N_1996);
and U3427 (N_3427,N_1629,N_785);
or U3428 (N_3428,N_979,N_81);
nand U3429 (N_3429,N_1528,N_1372);
nor U3430 (N_3430,N_425,N_1316);
and U3431 (N_3431,N_492,N_935);
nand U3432 (N_3432,N_1975,N_1652);
or U3433 (N_3433,N_57,N_1248);
nor U3434 (N_3434,N_1680,N_1647);
and U3435 (N_3435,N_704,N_1792);
and U3436 (N_3436,N_1592,N_884);
nor U3437 (N_3437,N_1415,N_909);
nor U3438 (N_3438,N_1488,N_225);
nor U3439 (N_3439,N_1885,N_1222);
and U3440 (N_3440,N_226,N_916);
nand U3441 (N_3441,N_1075,N_1307);
and U3442 (N_3442,N_1347,N_1551);
nor U3443 (N_3443,N_512,N_289);
or U3444 (N_3444,N_1291,N_1550);
nand U3445 (N_3445,N_1020,N_1718);
or U3446 (N_3446,N_1311,N_969);
and U3447 (N_3447,N_912,N_1631);
nand U3448 (N_3448,N_879,N_198);
nand U3449 (N_3449,N_615,N_1231);
and U3450 (N_3450,N_619,N_1692);
nand U3451 (N_3451,N_1432,N_1777);
or U3452 (N_3452,N_1778,N_722);
nor U3453 (N_3453,N_215,N_918);
nor U3454 (N_3454,N_334,N_583);
nand U3455 (N_3455,N_12,N_1474);
or U3456 (N_3456,N_1615,N_1673);
nand U3457 (N_3457,N_822,N_835);
or U3458 (N_3458,N_714,N_1819);
nand U3459 (N_3459,N_1475,N_875);
and U3460 (N_3460,N_1727,N_49);
nand U3461 (N_3461,N_1561,N_14);
or U3462 (N_3462,N_1237,N_1434);
nor U3463 (N_3463,N_48,N_739);
or U3464 (N_3464,N_915,N_1601);
or U3465 (N_3465,N_1104,N_874);
and U3466 (N_3466,N_98,N_545);
or U3467 (N_3467,N_1920,N_902);
or U3468 (N_3468,N_1303,N_1890);
nor U3469 (N_3469,N_1843,N_387);
nor U3470 (N_3470,N_1583,N_40);
and U3471 (N_3471,N_185,N_64);
nand U3472 (N_3472,N_1195,N_399);
nor U3473 (N_3473,N_176,N_696);
nor U3474 (N_3474,N_172,N_1983);
nand U3475 (N_3475,N_1839,N_65);
nand U3476 (N_3476,N_1558,N_1852);
nor U3477 (N_3477,N_1687,N_834);
nor U3478 (N_3478,N_1047,N_1998);
nand U3479 (N_3479,N_1584,N_812);
and U3480 (N_3480,N_735,N_1750);
nor U3481 (N_3481,N_340,N_1215);
and U3482 (N_3482,N_1643,N_614);
or U3483 (N_3483,N_714,N_1121);
and U3484 (N_3484,N_1217,N_1177);
nand U3485 (N_3485,N_892,N_266);
and U3486 (N_3486,N_757,N_1481);
nor U3487 (N_3487,N_938,N_515);
nand U3488 (N_3488,N_259,N_173);
nand U3489 (N_3489,N_792,N_1777);
or U3490 (N_3490,N_1420,N_836);
nand U3491 (N_3491,N_1403,N_1778);
nand U3492 (N_3492,N_1563,N_1456);
or U3493 (N_3493,N_506,N_1819);
nor U3494 (N_3494,N_43,N_501);
nor U3495 (N_3495,N_1390,N_710);
and U3496 (N_3496,N_716,N_1884);
and U3497 (N_3497,N_901,N_746);
or U3498 (N_3498,N_36,N_1294);
and U3499 (N_3499,N_1411,N_289);
and U3500 (N_3500,N_1866,N_66);
or U3501 (N_3501,N_1782,N_1227);
and U3502 (N_3502,N_983,N_1091);
nand U3503 (N_3503,N_1777,N_634);
nand U3504 (N_3504,N_1759,N_1835);
nor U3505 (N_3505,N_33,N_609);
and U3506 (N_3506,N_567,N_1635);
nor U3507 (N_3507,N_141,N_1690);
nand U3508 (N_3508,N_299,N_1718);
and U3509 (N_3509,N_1107,N_1624);
nor U3510 (N_3510,N_1222,N_1852);
nor U3511 (N_3511,N_1626,N_1444);
nor U3512 (N_3512,N_1519,N_12);
nand U3513 (N_3513,N_31,N_320);
nand U3514 (N_3514,N_1551,N_481);
nand U3515 (N_3515,N_511,N_921);
or U3516 (N_3516,N_246,N_1818);
xnor U3517 (N_3517,N_899,N_1805);
or U3518 (N_3518,N_498,N_1696);
or U3519 (N_3519,N_1051,N_1676);
or U3520 (N_3520,N_138,N_1322);
nor U3521 (N_3521,N_284,N_1418);
nor U3522 (N_3522,N_1051,N_1997);
nor U3523 (N_3523,N_1057,N_1079);
and U3524 (N_3524,N_19,N_82);
or U3525 (N_3525,N_740,N_742);
nor U3526 (N_3526,N_463,N_742);
and U3527 (N_3527,N_1461,N_130);
nor U3528 (N_3528,N_1016,N_315);
nand U3529 (N_3529,N_632,N_419);
nand U3530 (N_3530,N_366,N_1501);
or U3531 (N_3531,N_1039,N_1207);
or U3532 (N_3532,N_1171,N_748);
nor U3533 (N_3533,N_200,N_903);
nand U3534 (N_3534,N_1454,N_1212);
nor U3535 (N_3535,N_125,N_1680);
or U3536 (N_3536,N_1193,N_137);
or U3537 (N_3537,N_1244,N_1889);
nand U3538 (N_3538,N_1846,N_1288);
and U3539 (N_3539,N_1993,N_1610);
or U3540 (N_3540,N_1487,N_515);
nor U3541 (N_3541,N_166,N_1011);
or U3542 (N_3542,N_1460,N_54);
and U3543 (N_3543,N_627,N_667);
and U3544 (N_3544,N_929,N_595);
or U3545 (N_3545,N_1045,N_791);
nand U3546 (N_3546,N_1065,N_1527);
and U3547 (N_3547,N_1473,N_1578);
nand U3548 (N_3548,N_825,N_145);
and U3549 (N_3549,N_1734,N_53);
nor U3550 (N_3550,N_1689,N_323);
nand U3551 (N_3551,N_757,N_964);
or U3552 (N_3552,N_955,N_410);
and U3553 (N_3553,N_773,N_1186);
or U3554 (N_3554,N_1072,N_167);
and U3555 (N_3555,N_1132,N_1810);
nor U3556 (N_3556,N_1489,N_1746);
nor U3557 (N_3557,N_1237,N_1909);
nor U3558 (N_3558,N_158,N_1379);
or U3559 (N_3559,N_151,N_215);
nor U3560 (N_3560,N_1060,N_1929);
xor U3561 (N_3561,N_915,N_1347);
nor U3562 (N_3562,N_1472,N_1226);
and U3563 (N_3563,N_1708,N_1408);
or U3564 (N_3564,N_922,N_1461);
and U3565 (N_3565,N_353,N_689);
or U3566 (N_3566,N_107,N_1557);
or U3567 (N_3567,N_15,N_873);
nand U3568 (N_3568,N_508,N_1820);
nor U3569 (N_3569,N_1474,N_1417);
and U3570 (N_3570,N_702,N_1383);
nand U3571 (N_3571,N_961,N_1953);
nand U3572 (N_3572,N_1853,N_199);
nand U3573 (N_3573,N_550,N_155);
nand U3574 (N_3574,N_1502,N_1968);
and U3575 (N_3575,N_1038,N_488);
and U3576 (N_3576,N_651,N_802);
nand U3577 (N_3577,N_1688,N_1369);
and U3578 (N_3578,N_1172,N_686);
nor U3579 (N_3579,N_1235,N_916);
and U3580 (N_3580,N_341,N_1474);
nor U3581 (N_3581,N_710,N_1472);
and U3582 (N_3582,N_302,N_118);
nand U3583 (N_3583,N_1570,N_1544);
and U3584 (N_3584,N_273,N_1687);
and U3585 (N_3585,N_641,N_1863);
and U3586 (N_3586,N_769,N_66);
and U3587 (N_3587,N_1711,N_1301);
nor U3588 (N_3588,N_538,N_1247);
and U3589 (N_3589,N_505,N_1266);
and U3590 (N_3590,N_1671,N_791);
nor U3591 (N_3591,N_277,N_662);
nand U3592 (N_3592,N_407,N_400);
nand U3593 (N_3593,N_1098,N_758);
nor U3594 (N_3594,N_824,N_967);
or U3595 (N_3595,N_369,N_1580);
or U3596 (N_3596,N_1630,N_1887);
or U3597 (N_3597,N_1744,N_1629);
nor U3598 (N_3598,N_62,N_1479);
and U3599 (N_3599,N_1668,N_1272);
and U3600 (N_3600,N_577,N_1457);
or U3601 (N_3601,N_1672,N_1980);
or U3602 (N_3602,N_1819,N_1341);
or U3603 (N_3603,N_1390,N_331);
nor U3604 (N_3604,N_1796,N_592);
nor U3605 (N_3605,N_1577,N_1962);
nand U3606 (N_3606,N_1606,N_912);
and U3607 (N_3607,N_792,N_1074);
or U3608 (N_3608,N_904,N_275);
nor U3609 (N_3609,N_1340,N_1257);
or U3610 (N_3610,N_1006,N_437);
and U3611 (N_3611,N_1328,N_1219);
and U3612 (N_3612,N_1875,N_22);
or U3613 (N_3613,N_1065,N_1761);
nand U3614 (N_3614,N_294,N_946);
or U3615 (N_3615,N_1524,N_687);
nor U3616 (N_3616,N_847,N_741);
nor U3617 (N_3617,N_1479,N_1191);
or U3618 (N_3618,N_964,N_657);
nand U3619 (N_3619,N_1705,N_1450);
and U3620 (N_3620,N_624,N_1909);
nor U3621 (N_3621,N_544,N_632);
and U3622 (N_3622,N_1159,N_1941);
or U3623 (N_3623,N_1106,N_1759);
and U3624 (N_3624,N_1077,N_1946);
or U3625 (N_3625,N_1819,N_341);
xor U3626 (N_3626,N_187,N_1227);
or U3627 (N_3627,N_1141,N_1989);
nand U3628 (N_3628,N_1023,N_1288);
nor U3629 (N_3629,N_92,N_1865);
or U3630 (N_3630,N_1353,N_810);
nand U3631 (N_3631,N_1894,N_1291);
xor U3632 (N_3632,N_1735,N_620);
and U3633 (N_3633,N_1666,N_318);
and U3634 (N_3634,N_306,N_620);
xnor U3635 (N_3635,N_970,N_1475);
nor U3636 (N_3636,N_1817,N_190);
and U3637 (N_3637,N_1917,N_1079);
and U3638 (N_3638,N_1070,N_1773);
nand U3639 (N_3639,N_1306,N_1164);
or U3640 (N_3640,N_473,N_1951);
or U3641 (N_3641,N_1771,N_191);
and U3642 (N_3642,N_106,N_174);
or U3643 (N_3643,N_597,N_483);
nor U3644 (N_3644,N_267,N_678);
nor U3645 (N_3645,N_45,N_1527);
and U3646 (N_3646,N_1327,N_1188);
or U3647 (N_3647,N_181,N_435);
and U3648 (N_3648,N_819,N_299);
nor U3649 (N_3649,N_656,N_143);
nor U3650 (N_3650,N_230,N_1826);
nor U3651 (N_3651,N_1354,N_1539);
nor U3652 (N_3652,N_402,N_858);
nor U3653 (N_3653,N_742,N_117);
or U3654 (N_3654,N_143,N_6);
or U3655 (N_3655,N_1250,N_1868);
nor U3656 (N_3656,N_1788,N_1635);
nor U3657 (N_3657,N_1183,N_1976);
and U3658 (N_3658,N_1518,N_1181);
nor U3659 (N_3659,N_702,N_991);
or U3660 (N_3660,N_301,N_791);
and U3661 (N_3661,N_1508,N_485);
nand U3662 (N_3662,N_1720,N_150);
and U3663 (N_3663,N_1677,N_1916);
or U3664 (N_3664,N_1715,N_1546);
nor U3665 (N_3665,N_42,N_737);
nor U3666 (N_3666,N_205,N_1881);
and U3667 (N_3667,N_691,N_71);
nand U3668 (N_3668,N_17,N_1177);
nor U3669 (N_3669,N_1499,N_1208);
or U3670 (N_3670,N_1849,N_1791);
and U3671 (N_3671,N_936,N_664);
nor U3672 (N_3672,N_990,N_117);
and U3673 (N_3673,N_345,N_1380);
nor U3674 (N_3674,N_1776,N_1234);
nor U3675 (N_3675,N_858,N_1676);
or U3676 (N_3676,N_1777,N_114);
or U3677 (N_3677,N_910,N_872);
or U3678 (N_3678,N_843,N_1817);
and U3679 (N_3679,N_1357,N_1479);
nor U3680 (N_3680,N_636,N_55);
nor U3681 (N_3681,N_1977,N_1519);
nor U3682 (N_3682,N_1314,N_1564);
or U3683 (N_3683,N_800,N_1854);
or U3684 (N_3684,N_1522,N_974);
nand U3685 (N_3685,N_518,N_1737);
nand U3686 (N_3686,N_535,N_721);
nand U3687 (N_3687,N_1629,N_1557);
and U3688 (N_3688,N_226,N_855);
or U3689 (N_3689,N_1517,N_1373);
nand U3690 (N_3690,N_25,N_1208);
or U3691 (N_3691,N_1171,N_1825);
nor U3692 (N_3692,N_246,N_350);
or U3693 (N_3693,N_1707,N_792);
nand U3694 (N_3694,N_1319,N_1435);
and U3695 (N_3695,N_1654,N_1310);
nor U3696 (N_3696,N_1063,N_295);
xor U3697 (N_3697,N_1803,N_371);
nand U3698 (N_3698,N_1555,N_1352);
and U3699 (N_3699,N_1929,N_397);
or U3700 (N_3700,N_1958,N_1630);
nor U3701 (N_3701,N_1586,N_696);
or U3702 (N_3702,N_1783,N_1677);
nor U3703 (N_3703,N_110,N_558);
or U3704 (N_3704,N_632,N_1577);
and U3705 (N_3705,N_820,N_1866);
nor U3706 (N_3706,N_1335,N_1275);
nor U3707 (N_3707,N_881,N_573);
or U3708 (N_3708,N_859,N_1169);
and U3709 (N_3709,N_1895,N_983);
and U3710 (N_3710,N_78,N_130);
nand U3711 (N_3711,N_675,N_799);
nor U3712 (N_3712,N_1815,N_687);
nor U3713 (N_3713,N_422,N_1390);
nor U3714 (N_3714,N_1246,N_144);
nand U3715 (N_3715,N_1268,N_1756);
and U3716 (N_3716,N_1218,N_1254);
and U3717 (N_3717,N_112,N_1736);
nor U3718 (N_3718,N_912,N_506);
and U3719 (N_3719,N_457,N_554);
and U3720 (N_3720,N_167,N_1564);
or U3721 (N_3721,N_201,N_1108);
or U3722 (N_3722,N_1374,N_693);
or U3723 (N_3723,N_1354,N_1050);
and U3724 (N_3724,N_1739,N_1437);
and U3725 (N_3725,N_429,N_257);
nor U3726 (N_3726,N_1458,N_1501);
and U3727 (N_3727,N_1737,N_1572);
or U3728 (N_3728,N_1143,N_1834);
or U3729 (N_3729,N_1735,N_751);
nand U3730 (N_3730,N_801,N_1973);
and U3731 (N_3731,N_1837,N_927);
nand U3732 (N_3732,N_1083,N_608);
nand U3733 (N_3733,N_313,N_1074);
and U3734 (N_3734,N_706,N_1048);
nor U3735 (N_3735,N_552,N_243);
and U3736 (N_3736,N_1281,N_1519);
nor U3737 (N_3737,N_1634,N_99);
nand U3738 (N_3738,N_584,N_996);
and U3739 (N_3739,N_1157,N_259);
or U3740 (N_3740,N_1802,N_973);
nor U3741 (N_3741,N_1219,N_49);
nand U3742 (N_3742,N_421,N_337);
or U3743 (N_3743,N_624,N_996);
nand U3744 (N_3744,N_355,N_1137);
nor U3745 (N_3745,N_615,N_923);
nand U3746 (N_3746,N_998,N_984);
nand U3747 (N_3747,N_1364,N_1227);
or U3748 (N_3748,N_1804,N_1916);
nor U3749 (N_3749,N_1428,N_1347);
nand U3750 (N_3750,N_1477,N_612);
nor U3751 (N_3751,N_1836,N_1329);
nor U3752 (N_3752,N_112,N_1521);
nor U3753 (N_3753,N_967,N_1850);
and U3754 (N_3754,N_1648,N_665);
and U3755 (N_3755,N_372,N_1236);
and U3756 (N_3756,N_795,N_1226);
nor U3757 (N_3757,N_453,N_1168);
or U3758 (N_3758,N_89,N_1041);
nand U3759 (N_3759,N_147,N_762);
nand U3760 (N_3760,N_892,N_711);
and U3761 (N_3761,N_430,N_1917);
nor U3762 (N_3762,N_1513,N_1096);
nor U3763 (N_3763,N_203,N_89);
nor U3764 (N_3764,N_1128,N_1539);
nand U3765 (N_3765,N_634,N_308);
and U3766 (N_3766,N_723,N_1294);
nand U3767 (N_3767,N_1901,N_1112);
and U3768 (N_3768,N_1679,N_1667);
and U3769 (N_3769,N_329,N_767);
and U3770 (N_3770,N_677,N_58);
or U3771 (N_3771,N_197,N_1092);
and U3772 (N_3772,N_166,N_888);
xor U3773 (N_3773,N_1155,N_1679);
nand U3774 (N_3774,N_201,N_1963);
or U3775 (N_3775,N_1928,N_130);
nand U3776 (N_3776,N_1432,N_1572);
nor U3777 (N_3777,N_1904,N_596);
or U3778 (N_3778,N_273,N_1457);
or U3779 (N_3779,N_32,N_28);
and U3780 (N_3780,N_1976,N_693);
or U3781 (N_3781,N_430,N_1874);
nor U3782 (N_3782,N_738,N_1209);
nor U3783 (N_3783,N_45,N_1378);
or U3784 (N_3784,N_1618,N_981);
nor U3785 (N_3785,N_601,N_1717);
or U3786 (N_3786,N_1472,N_502);
or U3787 (N_3787,N_547,N_1083);
nand U3788 (N_3788,N_1184,N_1540);
or U3789 (N_3789,N_937,N_461);
or U3790 (N_3790,N_1256,N_41);
or U3791 (N_3791,N_1625,N_1709);
nor U3792 (N_3792,N_1701,N_787);
or U3793 (N_3793,N_234,N_298);
or U3794 (N_3794,N_1061,N_147);
nand U3795 (N_3795,N_1710,N_585);
nand U3796 (N_3796,N_421,N_1603);
nor U3797 (N_3797,N_84,N_901);
or U3798 (N_3798,N_1281,N_744);
nor U3799 (N_3799,N_1516,N_1394);
nor U3800 (N_3800,N_806,N_954);
and U3801 (N_3801,N_1582,N_1625);
nor U3802 (N_3802,N_109,N_1635);
and U3803 (N_3803,N_1953,N_1403);
or U3804 (N_3804,N_1550,N_1730);
and U3805 (N_3805,N_1361,N_1474);
and U3806 (N_3806,N_624,N_25);
and U3807 (N_3807,N_1664,N_1902);
nand U3808 (N_3808,N_991,N_779);
or U3809 (N_3809,N_174,N_555);
and U3810 (N_3810,N_1371,N_699);
and U3811 (N_3811,N_1845,N_1677);
or U3812 (N_3812,N_1802,N_1231);
nor U3813 (N_3813,N_1297,N_1278);
and U3814 (N_3814,N_885,N_1342);
xnor U3815 (N_3815,N_1912,N_218);
nand U3816 (N_3816,N_269,N_68);
or U3817 (N_3817,N_1067,N_139);
nor U3818 (N_3818,N_178,N_170);
nand U3819 (N_3819,N_1641,N_141);
and U3820 (N_3820,N_808,N_911);
nor U3821 (N_3821,N_1550,N_842);
and U3822 (N_3822,N_700,N_1791);
nor U3823 (N_3823,N_1522,N_233);
nand U3824 (N_3824,N_670,N_89);
and U3825 (N_3825,N_1393,N_223);
or U3826 (N_3826,N_1808,N_804);
nand U3827 (N_3827,N_471,N_930);
nand U3828 (N_3828,N_120,N_141);
or U3829 (N_3829,N_926,N_1951);
nand U3830 (N_3830,N_346,N_1467);
nand U3831 (N_3831,N_994,N_247);
nand U3832 (N_3832,N_612,N_619);
nand U3833 (N_3833,N_108,N_835);
and U3834 (N_3834,N_1366,N_1030);
and U3835 (N_3835,N_1207,N_344);
and U3836 (N_3836,N_939,N_567);
or U3837 (N_3837,N_891,N_1021);
nor U3838 (N_3838,N_385,N_623);
nor U3839 (N_3839,N_1425,N_1754);
nand U3840 (N_3840,N_1940,N_1070);
and U3841 (N_3841,N_1088,N_1119);
and U3842 (N_3842,N_252,N_291);
nor U3843 (N_3843,N_703,N_744);
or U3844 (N_3844,N_7,N_183);
nor U3845 (N_3845,N_588,N_1699);
nand U3846 (N_3846,N_1007,N_908);
and U3847 (N_3847,N_1408,N_1150);
nor U3848 (N_3848,N_1350,N_1029);
and U3849 (N_3849,N_1523,N_1567);
and U3850 (N_3850,N_419,N_828);
or U3851 (N_3851,N_1773,N_1646);
nand U3852 (N_3852,N_940,N_1376);
and U3853 (N_3853,N_1286,N_1952);
nor U3854 (N_3854,N_1307,N_1941);
nand U3855 (N_3855,N_677,N_274);
or U3856 (N_3856,N_944,N_324);
or U3857 (N_3857,N_1803,N_1864);
or U3858 (N_3858,N_1295,N_1880);
nand U3859 (N_3859,N_1239,N_931);
nor U3860 (N_3860,N_1342,N_1505);
or U3861 (N_3861,N_73,N_1908);
nand U3862 (N_3862,N_380,N_1838);
nand U3863 (N_3863,N_222,N_1005);
nor U3864 (N_3864,N_1613,N_948);
and U3865 (N_3865,N_1264,N_1750);
and U3866 (N_3866,N_811,N_516);
nor U3867 (N_3867,N_1854,N_1310);
or U3868 (N_3868,N_973,N_803);
nand U3869 (N_3869,N_1930,N_405);
or U3870 (N_3870,N_224,N_78);
nand U3871 (N_3871,N_165,N_1352);
nand U3872 (N_3872,N_1114,N_167);
and U3873 (N_3873,N_733,N_1763);
or U3874 (N_3874,N_736,N_484);
nand U3875 (N_3875,N_267,N_765);
nor U3876 (N_3876,N_503,N_1071);
and U3877 (N_3877,N_1639,N_69);
or U3878 (N_3878,N_1602,N_1056);
nand U3879 (N_3879,N_547,N_195);
nor U3880 (N_3880,N_1523,N_1209);
and U3881 (N_3881,N_208,N_482);
or U3882 (N_3882,N_379,N_1364);
or U3883 (N_3883,N_106,N_478);
nand U3884 (N_3884,N_801,N_538);
and U3885 (N_3885,N_1347,N_1649);
nand U3886 (N_3886,N_60,N_670);
nand U3887 (N_3887,N_688,N_1384);
nand U3888 (N_3888,N_305,N_667);
xor U3889 (N_3889,N_1966,N_570);
nor U3890 (N_3890,N_419,N_612);
nor U3891 (N_3891,N_722,N_221);
xor U3892 (N_3892,N_1479,N_1402);
or U3893 (N_3893,N_424,N_1915);
nor U3894 (N_3894,N_1859,N_1887);
nand U3895 (N_3895,N_320,N_1672);
nor U3896 (N_3896,N_1518,N_255);
nor U3897 (N_3897,N_202,N_1801);
nand U3898 (N_3898,N_861,N_469);
or U3899 (N_3899,N_1312,N_1868);
nor U3900 (N_3900,N_900,N_259);
and U3901 (N_3901,N_106,N_875);
or U3902 (N_3902,N_230,N_233);
nand U3903 (N_3903,N_828,N_1999);
and U3904 (N_3904,N_1099,N_41);
and U3905 (N_3905,N_259,N_533);
and U3906 (N_3906,N_24,N_1360);
nor U3907 (N_3907,N_883,N_89);
nor U3908 (N_3908,N_1873,N_257);
nand U3909 (N_3909,N_952,N_1600);
and U3910 (N_3910,N_657,N_880);
and U3911 (N_3911,N_1374,N_631);
and U3912 (N_3912,N_520,N_918);
nand U3913 (N_3913,N_585,N_917);
or U3914 (N_3914,N_1788,N_1477);
and U3915 (N_3915,N_233,N_557);
or U3916 (N_3916,N_540,N_801);
nand U3917 (N_3917,N_1938,N_773);
or U3918 (N_3918,N_265,N_1739);
nand U3919 (N_3919,N_1298,N_1476);
nor U3920 (N_3920,N_795,N_1086);
nor U3921 (N_3921,N_1794,N_1443);
nor U3922 (N_3922,N_352,N_304);
nand U3923 (N_3923,N_798,N_511);
or U3924 (N_3924,N_500,N_1911);
nor U3925 (N_3925,N_990,N_703);
or U3926 (N_3926,N_1770,N_1864);
nand U3927 (N_3927,N_712,N_332);
and U3928 (N_3928,N_1824,N_1856);
nor U3929 (N_3929,N_1003,N_1065);
xnor U3930 (N_3930,N_701,N_1135);
nand U3931 (N_3931,N_515,N_1976);
nand U3932 (N_3932,N_1746,N_1240);
nand U3933 (N_3933,N_158,N_595);
and U3934 (N_3934,N_21,N_1671);
nand U3935 (N_3935,N_1445,N_1978);
and U3936 (N_3936,N_67,N_1295);
and U3937 (N_3937,N_435,N_1085);
and U3938 (N_3938,N_1023,N_1763);
nor U3939 (N_3939,N_1836,N_1153);
or U3940 (N_3940,N_937,N_1890);
or U3941 (N_3941,N_1165,N_467);
or U3942 (N_3942,N_1259,N_296);
nor U3943 (N_3943,N_713,N_237);
nor U3944 (N_3944,N_554,N_281);
nor U3945 (N_3945,N_191,N_857);
nor U3946 (N_3946,N_982,N_384);
nor U3947 (N_3947,N_663,N_724);
and U3948 (N_3948,N_1659,N_1909);
nor U3949 (N_3949,N_1515,N_1022);
nand U3950 (N_3950,N_552,N_322);
nor U3951 (N_3951,N_405,N_1980);
or U3952 (N_3952,N_971,N_981);
nor U3953 (N_3953,N_1508,N_199);
nand U3954 (N_3954,N_49,N_1973);
or U3955 (N_3955,N_1701,N_1424);
nand U3956 (N_3956,N_1252,N_1038);
nor U3957 (N_3957,N_903,N_299);
nand U3958 (N_3958,N_533,N_302);
and U3959 (N_3959,N_1119,N_1641);
or U3960 (N_3960,N_1600,N_625);
or U3961 (N_3961,N_991,N_25);
nor U3962 (N_3962,N_1041,N_200);
and U3963 (N_3963,N_1912,N_1199);
and U3964 (N_3964,N_599,N_203);
nor U3965 (N_3965,N_222,N_310);
and U3966 (N_3966,N_360,N_1261);
nor U3967 (N_3967,N_463,N_1063);
and U3968 (N_3968,N_1908,N_1395);
nor U3969 (N_3969,N_1817,N_678);
and U3970 (N_3970,N_1116,N_168);
or U3971 (N_3971,N_546,N_1403);
nor U3972 (N_3972,N_1289,N_354);
nand U3973 (N_3973,N_1085,N_506);
and U3974 (N_3974,N_1642,N_280);
nand U3975 (N_3975,N_560,N_917);
and U3976 (N_3976,N_818,N_592);
nand U3977 (N_3977,N_1611,N_1673);
or U3978 (N_3978,N_1534,N_1267);
and U3979 (N_3979,N_1386,N_1987);
nand U3980 (N_3980,N_1585,N_1359);
and U3981 (N_3981,N_1692,N_1927);
and U3982 (N_3982,N_820,N_698);
or U3983 (N_3983,N_1107,N_1407);
nor U3984 (N_3984,N_1059,N_1994);
nand U3985 (N_3985,N_1626,N_1827);
nand U3986 (N_3986,N_1248,N_1874);
nand U3987 (N_3987,N_1203,N_1444);
nor U3988 (N_3988,N_1928,N_997);
or U3989 (N_3989,N_1367,N_1167);
nor U3990 (N_3990,N_1102,N_1067);
nand U3991 (N_3991,N_368,N_698);
nor U3992 (N_3992,N_160,N_1684);
or U3993 (N_3993,N_1925,N_999);
and U3994 (N_3994,N_1772,N_99);
and U3995 (N_3995,N_1848,N_332);
nand U3996 (N_3996,N_1732,N_1650);
nor U3997 (N_3997,N_882,N_853);
or U3998 (N_3998,N_1788,N_487);
and U3999 (N_3999,N_697,N_690);
and U4000 (N_4000,N_3527,N_2662);
or U4001 (N_4001,N_3362,N_3133);
nand U4002 (N_4002,N_2219,N_2546);
and U4003 (N_4003,N_2759,N_2770);
nand U4004 (N_4004,N_3454,N_2796);
or U4005 (N_4005,N_3152,N_2829);
and U4006 (N_4006,N_2808,N_2267);
or U4007 (N_4007,N_2297,N_2009);
nand U4008 (N_4008,N_3002,N_3483);
nor U4009 (N_4009,N_2221,N_3179);
or U4010 (N_4010,N_2892,N_2830);
xor U4011 (N_4011,N_2484,N_2855);
xor U4012 (N_4012,N_2817,N_2913);
or U4013 (N_4013,N_3931,N_2605);
nand U4014 (N_4014,N_2214,N_2055);
or U4015 (N_4015,N_2062,N_3218);
nor U4016 (N_4016,N_3741,N_2255);
and U4017 (N_4017,N_3350,N_2835);
and U4018 (N_4018,N_3269,N_2001);
nor U4019 (N_4019,N_2491,N_3544);
nand U4020 (N_4020,N_2399,N_3297);
or U4021 (N_4021,N_3719,N_3800);
and U4022 (N_4022,N_3558,N_2338);
and U4023 (N_4023,N_2740,N_2092);
nand U4024 (N_4024,N_3825,N_3986);
and U4025 (N_4025,N_2511,N_2564);
or U4026 (N_4026,N_3828,N_2436);
nand U4027 (N_4027,N_2642,N_3016);
and U4028 (N_4028,N_3457,N_2993);
nor U4029 (N_4029,N_2296,N_2198);
and U4030 (N_4030,N_2773,N_2037);
nand U4031 (N_4031,N_2164,N_2457);
nand U4032 (N_4032,N_3018,N_2506);
nor U4033 (N_4033,N_2695,N_2646);
and U4034 (N_4034,N_2456,N_3019);
and U4035 (N_4035,N_3170,N_2344);
and U4036 (N_4036,N_3492,N_3335);
nand U4037 (N_4037,N_2444,N_3441);
nand U4038 (N_4038,N_3522,N_2420);
or U4039 (N_4039,N_3562,N_2609);
or U4040 (N_4040,N_2868,N_2314);
and U4041 (N_4041,N_3949,N_2811);
nand U4042 (N_4042,N_3447,N_2096);
and U4043 (N_4043,N_3216,N_2772);
nand U4044 (N_4044,N_3981,N_3526);
and U4045 (N_4045,N_2714,N_2225);
nor U4046 (N_4046,N_2734,N_2348);
or U4047 (N_4047,N_2432,N_3320);
nor U4048 (N_4048,N_2885,N_3590);
or U4049 (N_4049,N_3213,N_3137);
nand U4050 (N_4050,N_3736,N_3337);
and U4051 (N_4051,N_3932,N_3649);
or U4052 (N_4052,N_3879,N_3980);
nand U4053 (N_4053,N_2015,N_3338);
or U4054 (N_4054,N_3095,N_3472);
or U4055 (N_4055,N_2223,N_2560);
or U4056 (N_4056,N_2746,N_2072);
or U4057 (N_4057,N_2732,N_2921);
nor U4058 (N_4058,N_3729,N_2794);
nor U4059 (N_4059,N_2032,N_3721);
or U4060 (N_4060,N_3596,N_3153);
nand U4061 (N_4061,N_3233,N_3129);
or U4062 (N_4062,N_3336,N_2115);
or U4063 (N_4063,N_3407,N_2607);
nor U4064 (N_4064,N_3554,N_3831);
nand U4065 (N_4065,N_3486,N_2720);
nor U4066 (N_4066,N_2659,N_3965);
nor U4067 (N_4067,N_2683,N_2899);
and U4068 (N_4068,N_2602,N_2128);
nor U4069 (N_4069,N_2136,N_2745);
nand U4070 (N_4070,N_3160,N_2922);
and U4071 (N_4071,N_2814,N_3571);
or U4072 (N_4072,N_3185,N_3126);
or U4073 (N_4073,N_3523,N_2983);
and U4074 (N_4074,N_2027,N_3164);
nand U4075 (N_4075,N_3491,N_2701);
nand U4076 (N_4076,N_3037,N_2345);
nand U4077 (N_4077,N_3263,N_2100);
nand U4078 (N_4078,N_2372,N_3911);
and U4079 (N_4079,N_2858,N_2328);
or U4080 (N_4080,N_2337,N_2448);
nand U4081 (N_4081,N_2961,N_2850);
nand U4082 (N_4082,N_2341,N_3592);
nor U4083 (N_4083,N_3833,N_3574);
nor U4084 (N_4084,N_2790,N_3538);
and U4085 (N_4085,N_2053,N_2269);
and U4086 (N_4086,N_2857,N_3070);
and U4087 (N_4087,N_2815,N_2586);
or U4088 (N_4088,N_3535,N_2180);
nor U4089 (N_4089,N_2631,N_2091);
nand U4090 (N_4090,N_2622,N_3021);
and U4091 (N_4091,N_2499,N_2893);
nand U4092 (N_4092,N_3174,N_2613);
nor U4093 (N_4093,N_2925,N_2901);
nor U4094 (N_4094,N_3244,N_3098);
and U4095 (N_4095,N_3498,N_2867);
nor U4096 (N_4096,N_2612,N_2936);
nand U4097 (N_4097,N_3915,N_2521);
nand U4098 (N_4098,N_2524,N_2633);
nor U4099 (N_4099,N_2283,N_2391);
nand U4100 (N_4100,N_3272,N_3248);
or U4101 (N_4101,N_2236,N_3751);
and U4102 (N_4102,N_3670,N_2816);
nor U4103 (N_4103,N_2856,N_2368);
nor U4104 (N_4104,N_2020,N_2119);
or U4105 (N_4105,N_3897,N_3893);
nor U4106 (N_4106,N_2923,N_3587);
and U4107 (N_4107,N_2805,N_2441);
nand U4108 (N_4108,N_3807,N_3062);
nand U4109 (N_4109,N_3926,N_2260);
nor U4110 (N_4110,N_3103,N_3092);
nand U4111 (N_4111,N_2292,N_2543);
and U4112 (N_4112,N_3977,N_3907);
nand U4113 (N_4113,N_2252,N_2628);
or U4114 (N_4114,N_2452,N_3579);
or U4115 (N_4115,N_2113,N_3165);
and U4116 (N_4116,N_2464,N_2016);
or U4117 (N_4117,N_3533,N_2208);
or U4118 (N_4118,N_3740,N_3324);
or U4119 (N_4119,N_2472,N_3642);
nand U4120 (N_4120,N_3270,N_2237);
nand U4121 (N_4121,N_2634,N_2266);
or U4122 (N_4122,N_3656,N_2625);
or U4123 (N_4123,N_2534,N_3359);
and U4124 (N_4124,N_2361,N_3341);
nand U4125 (N_4125,N_2851,N_3476);
or U4126 (N_4126,N_3291,N_3937);
and U4127 (N_4127,N_2183,N_2986);
and U4128 (N_4128,N_2501,N_3434);
or U4129 (N_4129,N_2308,N_2552);
nand U4130 (N_4130,N_3936,N_2496);
or U4131 (N_4131,N_3307,N_2247);
or U4132 (N_4132,N_2881,N_2764);
or U4133 (N_4133,N_3870,N_2199);
nand U4134 (N_4134,N_3022,N_2959);
or U4135 (N_4135,N_3795,N_2381);
nand U4136 (N_4136,N_3573,N_2486);
and U4137 (N_4137,N_3859,N_3525);
and U4138 (N_4138,N_2437,N_2778);
nor U4139 (N_4139,N_2042,N_2660);
nor U4140 (N_4140,N_3349,N_3867);
nand U4141 (N_4141,N_2044,N_3757);
nand U4142 (N_4142,N_2974,N_2641);
and U4143 (N_4143,N_3256,N_2752);
nor U4144 (N_4144,N_3032,N_3509);
and U4145 (N_4145,N_2782,N_3678);
and U4146 (N_4146,N_3763,N_3452);
nand U4147 (N_4147,N_3116,N_3396);
or U4148 (N_4148,N_3258,N_2415);
and U4149 (N_4149,N_2911,N_3553);
nand U4150 (N_4150,N_3329,N_2860);
nand U4151 (N_4151,N_3505,N_2476);
or U4152 (N_4152,N_3781,N_3626);
nand U4153 (N_4153,N_2271,N_3952);
or U4154 (N_4154,N_3245,N_2011);
nand U4155 (N_4155,N_2249,N_3632);
or U4156 (N_4156,N_3752,N_3882);
nor U4157 (N_4157,N_2987,N_3119);
nor U4158 (N_4158,N_3265,N_3809);
nor U4159 (N_4159,N_2008,N_3992);
and U4160 (N_4160,N_3207,N_3139);
xor U4161 (N_4161,N_3894,N_3344);
or U4162 (N_4162,N_2056,N_2114);
nand U4163 (N_4163,N_3797,N_3792);
nand U4164 (N_4164,N_3629,N_3841);
and U4165 (N_4165,N_2301,N_2919);
nor U4166 (N_4166,N_2175,N_2066);
or U4167 (N_4167,N_2801,N_3203);
nand U4168 (N_4168,N_2567,N_3123);
nand U4169 (N_4169,N_3730,N_3167);
nand U4170 (N_4170,N_3104,N_3765);
and U4171 (N_4171,N_3351,N_3438);
nand U4172 (N_4172,N_3379,N_2905);
and U4173 (N_4173,N_2243,N_2848);
nor U4174 (N_4174,N_2333,N_2562);
or U4175 (N_4175,N_3470,N_2654);
and U4176 (N_4176,N_3951,N_2258);
nand U4177 (N_4177,N_3237,N_2369);
nand U4178 (N_4178,N_2343,N_3542);
and U4179 (N_4179,N_2194,N_3517);
and U4180 (N_4180,N_2653,N_3617);
or U4181 (N_4181,N_2460,N_3520);
nand U4182 (N_4182,N_2742,N_2080);
or U4183 (N_4183,N_3051,N_3717);
nor U4184 (N_4184,N_3898,N_3425);
or U4185 (N_4185,N_3661,N_3724);
or U4186 (N_4186,N_2234,N_3727);
nor U4187 (N_4187,N_2733,N_3653);
and U4188 (N_4188,N_3837,N_3424);
nand U4189 (N_4189,N_3249,N_2182);
nand U4190 (N_4190,N_2173,N_3844);
nor U4191 (N_4191,N_3427,N_3159);
and U4192 (N_4192,N_3501,N_3246);
nor U4193 (N_4193,N_3300,N_3857);
or U4194 (N_4194,N_2294,N_3355);
or U4195 (N_4195,N_3384,N_3261);
nor U4196 (N_4196,N_2468,N_2412);
and U4197 (N_4197,N_3845,N_2085);
nand U4198 (N_4198,N_3530,N_3848);
and U4199 (N_4199,N_2865,N_3761);
nand U4200 (N_4200,N_3465,N_3776);
nor U4201 (N_4201,N_3439,N_3035);
or U4202 (N_4202,N_3577,N_2665);
and U4203 (N_4203,N_2050,N_3105);
nor U4204 (N_4204,N_2095,N_2540);
or U4205 (N_4205,N_3356,N_3658);
and U4206 (N_4206,N_3496,N_3923);
nor U4207 (N_4207,N_2087,N_3064);
or U4208 (N_4208,N_3340,N_2058);
nand U4209 (N_4209,N_3855,N_2135);
nand U4210 (N_4210,N_2282,N_2942);
or U4211 (N_4211,N_3777,N_3302);
nand U4212 (N_4212,N_2195,N_3918);
or U4213 (N_4213,N_3197,N_2580);
nor U4214 (N_4214,N_3330,N_3896);
or U4215 (N_4215,N_3838,N_2469);
or U4216 (N_4216,N_3947,N_3706);
or U4217 (N_4217,N_2226,N_3110);
or U4218 (N_4218,N_2075,N_3047);
nor U4219 (N_4219,N_3122,N_3753);
nor U4220 (N_4220,N_3933,N_2869);
nor U4221 (N_4221,N_2725,N_3108);
and U4222 (N_4222,N_3784,N_3823);
and U4223 (N_4223,N_2112,N_3860);
nor U4224 (N_4224,N_2021,N_2022);
and U4225 (N_4225,N_2853,N_2106);
or U4226 (N_4226,N_3488,N_2310);
nor U4227 (N_4227,N_2661,N_2006);
or U4228 (N_4228,N_2120,N_3059);
or U4229 (N_4229,N_3914,N_2263);
nor U4230 (N_4230,N_2786,N_2376);
or U4231 (N_4231,N_3429,N_2099);
or U4232 (N_4232,N_3886,N_3537);
xnor U4233 (N_4233,N_3487,N_3169);
nor U4234 (N_4234,N_3614,N_3917);
and U4235 (N_4235,N_2585,N_3696);
or U4236 (N_4236,N_2047,N_3690);
nor U4237 (N_4237,N_2411,N_3872);
and U4238 (N_4238,N_3830,N_3053);
nor U4239 (N_4239,N_3399,N_2902);
or U4240 (N_4240,N_3217,N_2553);
or U4241 (N_4241,N_3783,N_2823);
or U4242 (N_4242,N_3173,N_2466);
xor U4243 (N_4243,N_3404,N_3054);
nand U4244 (N_4244,N_3143,N_2317);
nor U4245 (N_4245,N_2272,N_3599);
nor U4246 (N_4246,N_2802,N_2677);
nand U4247 (N_4247,N_2880,N_3093);
nor U4248 (N_4248,N_2256,N_3728);
and U4249 (N_4249,N_3085,N_3497);
nor U4250 (N_4250,N_3227,N_3387);
nand U4251 (N_4251,N_3353,N_2211);
nand U4252 (N_4252,N_2969,N_2557);
or U4253 (N_4253,N_2280,N_2445);
and U4254 (N_4254,N_2556,N_2516);
nand U4255 (N_4255,N_2088,N_2862);
nor U4256 (N_4256,N_2700,N_3885);
nand U4257 (N_4257,N_3323,N_2680);
or U4258 (N_4258,N_3076,N_2825);
and U4259 (N_4259,N_3735,N_3725);
or U4260 (N_4260,N_2202,N_3023);
nor U4261 (N_4261,N_2629,N_2224);
and U4262 (N_4262,N_3257,N_2584);
nand U4263 (N_4263,N_3423,N_2155);
and U4264 (N_4264,N_3821,N_3887);
nor U4265 (N_4265,N_3166,N_3565);
and U4266 (N_4266,N_3625,N_3769);
nand U4267 (N_4267,N_2596,N_2005);
nor U4268 (N_4268,N_2941,N_2357);
or U4269 (N_4269,N_2065,N_2434);
and U4270 (N_4270,N_3140,N_3546);
or U4271 (N_4271,N_2757,N_3332);
and U4272 (N_4272,N_3645,N_3071);
and U4273 (N_4273,N_3552,N_3541);
or U4274 (N_4274,N_3682,N_2510);
nand U4275 (N_4275,N_3333,N_3118);
nor U4276 (N_4276,N_2209,N_3940);
and U4277 (N_4277,N_2064,N_2029);
and U4278 (N_4278,N_2687,N_3964);
nand U4279 (N_4279,N_3989,N_3087);
nand U4280 (N_4280,N_2396,N_3770);
nor U4281 (N_4281,N_3111,N_2821);
and U4282 (N_4282,N_3667,N_2531);
and U4283 (N_4283,N_2404,N_2723);
or U4284 (N_4284,N_2356,N_3467);
nand U4285 (N_4285,N_3292,N_2323);
and U4286 (N_4286,N_3874,N_3175);
and U4287 (N_4287,N_2528,N_3722);
nor U4288 (N_4288,N_3146,N_2471);
or U4289 (N_4289,N_2388,N_3268);
nand U4290 (N_4290,N_3827,N_3539);
nand U4291 (N_4291,N_3774,N_2241);
or U4292 (N_4292,N_3773,N_2306);
nor U4293 (N_4293,N_2244,N_2769);
nand U4294 (N_4294,N_2077,N_2409);
and U4295 (N_4295,N_3796,N_3178);
and U4296 (N_4296,N_3982,N_2929);
and U4297 (N_4297,N_2826,N_3061);
and U4298 (N_4298,N_2657,N_2229);
nor U4299 (N_4299,N_2274,N_2648);
nor U4300 (N_4300,N_2481,N_2141);
and U4301 (N_4301,N_2693,N_3365);
or U4302 (N_4302,N_2994,N_2390);
nor U4303 (N_4303,N_2889,N_3611);
or U4304 (N_4304,N_2908,N_2439);
nand U4305 (N_4305,N_3475,N_3073);
or U4306 (N_4306,N_3935,N_3694);
nand U4307 (N_4307,N_3556,N_3508);
and U4308 (N_4308,N_2614,N_3473);
nand U4309 (N_4309,N_3041,N_3666);
nand U4310 (N_4310,N_2799,N_2205);
or U4311 (N_4311,N_3102,N_3762);
and U4312 (N_4312,N_3230,N_3127);
or U4313 (N_4313,N_3704,N_3091);
nand U4314 (N_4314,N_3540,N_2218);
nor U4315 (N_4315,N_3929,N_2309);
or U4316 (N_4316,N_2101,N_2964);
and U4317 (N_4317,N_3842,N_3096);
nor U4318 (N_4318,N_2325,N_2321);
and U4319 (N_4319,N_3288,N_3331);
nor U4320 (N_4320,N_2918,N_3798);
nor U4321 (N_4321,N_2876,N_2474);
nand U4322 (N_4322,N_2378,N_2122);
and U4323 (N_4323,N_2952,N_3938);
nor U4324 (N_4324,N_3328,N_3843);
or U4325 (N_4325,N_2318,N_3089);
and U4326 (N_4326,N_2783,N_2289);
nand U4327 (N_4327,N_3601,N_2104);
nand U4328 (N_4328,N_2590,N_2842);
or U4329 (N_4329,N_3186,N_2386);
nand U4330 (N_4330,N_3416,N_2193);
and U4331 (N_4331,N_2281,N_3716);
nand U4332 (N_4332,N_3005,N_3036);
nor U4333 (N_4333,N_3279,N_2645);
nand U4334 (N_4334,N_2771,N_2618);
or U4335 (N_4335,N_3260,N_3731);
and U4336 (N_4336,N_2354,N_2026);
or U4337 (N_4337,N_2713,N_3188);
nor U4338 (N_4338,N_2569,N_3144);
and U4339 (N_4339,N_3619,N_2950);
and U4340 (N_4340,N_3668,N_2877);
or U4341 (N_4341,N_3689,N_2859);
nand U4342 (N_4342,N_2279,N_3247);
and U4343 (N_4343,N_2762,N_3634);
or U4344 (N_4344,N_2897,N_2558);
and U4345 (N_4345,N_2517,N_3495);
nor U4346 (N_4346,N_3060,N_3255);
nand U4347 (N_4347,N_2520,N_3132);
or U4348 (N_4348,N_3507,N_3313);
and U4349 (N_4349,N_3602,N_2571);
nand U4350 (N_4350,N_3504,N_3280);
or U4351 (N_4351,N_3976,N_3794);
and U4352 (N_4352,N_2477,N_2674);
nand U4353 (N_4353,N_2467,N_3945);
or U4354 (N_4354,N_2664,N_3606);
nand U4355 (N_4355,N_3615,N_2611);
or U4356 (N_4356,N_2672,N_2233);
nand U4357 (N_4357,N_3436,N_2383);
nor U4358 (N_4358,N_3589,N_3450);
nand U4359 (N_4359,N_2153,N_2615);
or U4360 (N_4360,N_3361,N_3881);
nand U4361 (N_4361,N_3223,N_2206);
or U4362 (N_4362,N_2573,N_2139);
nand U4363 (N_4363,N_2545,N_3618);
and U4364 (N_4364,N_3180,N_3622);
nand U4365 (N_4365,N_3339,N_3010);
nand U4366 (N_4366,N_3824,N_2691);
and U4367 (N_4367,N_3636,N_3851);
nand U4368 (N_4368,N_2428,N_2709);
nand U4369 (N_4369,N_2161,N_2960);
nand U4370 (N_4370,N_3250,N_2424);
and U4371 (N_4371,N_2400,N_3754);
nor U4372 (N_4372,N_2530,N_3393);
nand U4373 (N_4373,N_2313,N_2462);
nor U4374 (N_4374,N_2559,N_3275);
nand U4375 (N_4375,N_2675,N_3063);
nor U4376 (N_4376,N_2363,N_2103);
nor U4377 (N_4377,N_3580,N_2751);
nand U4378 (N_4378,N_3866,N_3397);
nor U4379 (N_4379,N_3746,N_3647);
xor U4380 (N_4380,N_2346,N_2600);
nor U4381 (N_4381,N_3009,N_2846);
and U4382 (N_4382,N_2666,N_3147);
or U4383 (N_4383,N_3162,N_3083);
nand U4384 (N_4384,N_2163,N_2597);
and U4385 (N_4385,N_3368,N_2152);
nand U4386 (N_4386,N_3832,N_2753);
or U4387 (N_4387,N_3518,N_2895);
nor U4388 (N_4388,N_3999,N_3806);
or U4389 (N_4389,N_2030,N_3942);
nor U4390 (N_4390,N_2362,N_2339);
nand U4391 (N_4391,N_2698,N_2638);
or U4392 (N_4392,N_2507,N_2920);
nand U4393 (N_4393,N_3304,N_3171);
nand U4394 (N_4394,N_3869,N_2930);
nand U4395 (N_4395,N_3478,N_2603);
or U4396 (N_4396,N_2380,N_2627);
nand U4397 (N_4397,N_2326,N_3354);
nor U4398 (N_4398,N_2991,N_2906);
and U4399 (N_4399,N_3299,N_2126);
nor U4400 (N_4400,N_2288,N_2957);
or U4401 (N_4401,N_3681,N_2111);
nand U4402 (N_4402,N_2210,N_3057);
or U4403 (N_4403,N_3386,N_2480);
nand U4404 (N_4404,N_3804,N_3639);
nor U4405 (N_4405,N_2954,N_2347);
nor U4406 (N_4406,N_3586,N_2433);
nand U4407 (N_4407,N_3748,N_2475);
or U4408 (N_4408,N_3998,N_2788);
nand U4409 (N_4409,N_2084,N_2440);
or U4410 (N_4410,N_2169,N_2744);
nand U4411 (N_4411,N_2777,N_2156);
and U4412 (N_4412,N_3364,N_3876);
nor U4413 (N_4413,N_3201,N_2818);
or U4414 (N_4414,N_2685,N_2054);
nand U4415 (N_4415,N_2013,N_3309);
nor U4416 (N_4416,N_2003,N_2048);
and U4417 (N_4417,N_2676,N_3853);
or U4418 (N_4418,N_2536,N_3377);
or U4419 (N_4419,N_3901,N_2747);
nand U4420 (N_4420,N_2765,N_3908);
or U4421 (N_4421,N_2217,N_3817);
nand U4422 (N_4422,N_3902,N_2105);
nand U4423 (N_4423,N_2542,N_3004);
nor U4424 (N_4424,N_2130,N_2541);
nor U4425 (N_4425,N_2191,N_3008);
or U4426 (N_4426,N_3904,N_2330);
and U4427 (N_4427,N_3996,N_3068);
nand U4428 (N_4428,N_3701,N_2010);
nor U4429 (N_4429,N_2538,N_2978);
or U4430 (N_4430,N_2512,N_3972);
or U4431 (N_4431,N_2593,N_2355);
nand U4432 (N_4432,N_3778,N_2839);
and U4433 (N_4433,N_2081,N_2264);
and U4434 (N_4434,N_2488,N_3380);
nand U4435 (N_4435,N_3563,N_3868);
nor U4436 (N_4436,N_2350,N_3308);
nor U4437 (N_4437,N_3529,N_2207);
and U4438 (N_4438,N_3381,N_3849);
or U4439 (N_4439,N_2490,N_3657);
nor U4440 (N_4440,N_3766,N_2358);
or U4441 (N_4441,N_2915,N_2425);
nand U4442 (N_4442,N_2150,N_2188);
or U4443 (N_4443,N_3613,N_3994);
nand U4444 (N_4444,N_2785,N_3506);
nor U4445 (N_4445,N_3097,N_2177);
and U4446 (N_4446,N_3455,N_3829);
nor U4447 (N_4447,N_2841,N_3814);
or U4448 (N_4448,N_3745,N_3081);
nor U4449 (N_4449,N_3531,N_3305);
and U4450 (N_4450,N_2470,N_2537);
nand U4451 (N_4451,N_3459,N_3759);
and U4452 (N_4452,N_2431,N_3576);
and U4453 (N_4453,N_3603,N_2623);
or U4454 (N_4454,N_3079,N_2485);
nor U4455 (N_4455,N_3077,N_2621);
or U4456 (N_4456,N_2566,N_2767);
or U4457 (N_4457,N_3643,N_3408);
and U4458 (N_4458,N_3259,N_2928);
nor U4459 (N_4459,N_3939,N_2423);
nor U4460 (N_4460,N_3718,N_2703);
or U4461 (N_4461,N_2756,N_3094);
nand U4462 (N_4462,N_2663,N_3030);
or U4463 (N_4463,N_3462,N_2133);
nand U4464 (N_4464,N_3409,N_3673);
nor U4465 (N_4465,N_2688,N_3148);
nor U4466 (N_4466,N_3225,N_3298);
and U4467 (N_4467,N_3732,N_3637);
and U4468 (N_4468,N_2966,N_3967);
or U4469 (N_4469,N_2232,N_2340);
nand U4470 (N_4470,N_2242,N_3708);
and U4471 (N_4471,N_3922,N_3948);
or U4472 (N_4472,N_3691,N_3873);
nand U4473 (N_4473,N_3241,N_3055);
nor U4474 (N_4474,N_2483,N_3569);
and U4475 (N_4475,N_3209,N_3243);
nor U4476 (N_4476,N_3418,N_2426);
and U4477 (N_4477,N_2360,N_3446);
nor U4478 (N_4478,N_2250,N_3510);
or U4479 (N_4479,N_2254,N_3480);
nor U4480 (N_4480,N_3818,N_2429);
and U4481 (N_4481,N_2148,N_3394);
and U4482 (N_4482,N_3193,N_3374);
nand U4483 (N_4483,N_2178,N_2827);
or U4484 (N_4484,N_3946,N_2043);
and U4485 (N_4485,N_3226,N_3371);
nand U4486 (N_4486,N_3229,N_2215);
and U4487 (N_4487,N_2729,N_2787);
and U4488 (N_4488,N_3663,N_3805);
or U4489 (N_4489,N_3543,N_3199);
and U4490 (N_4490,N_3865,N_3206);
nor U4491 (N_4491,N_2131,N_3802);
nand U4492 (N_4492,N_3316,N_2555);
or U4493 (N_4493,N_2063,N_3957);
or U4494 (N_4494,N_3034,N_2976);
or U4495 (N_4495,N_2179,N_3767);
nor U4496 (N_4496,N_2806,N_3052);
or U4497 (N_4497,N_2270,N_3084);
nor U4498 (N_4498,N_3950,N_2414);
nand U4499 (N_4499,N_2334,N_3327);
nor U4500 (N_4500,N_3107,N_2981);
and U4501 (N_4501,N_2840,N_3130);
or U4502 (N_4502,N_3712,N_3567);
nor U4503 (N_4503,N_2387,N_2327);
or U4504 (N_4504,N_2563,N_2682);
nand U4505 (N_4505,N_3685,N_2572);
nor U4506 (N_4506,N_3145,N_3700);
nor U4507 (N_4507,N_2982,N_3560);
and U4508 (N_4508,N_2743,N_3743);
nor U4509 (N_4509,N_2820,N_2227);
or U4510 (N_4510,N_2097,N_2040);
nor U4511 (N_4511,N_3934,N_2004);
nand U4512 (N_4512,N_2766,N_3990);
or U4513 (N_4513,N_2293,N_2626);
or U4514 (N_4514,N_3286,N_3966);
nand U4515 (N_4515,N_2172,N_3044);
nand U4516 (N_4516,N_3065,N_2392);
nor U4517 (N_4517,N_2946,N_2776);
and U4518 (N_4518,N_3750,N_2800);
nand U4519 (N_4519,N_2945,N_2953);
and U4520 (N_4520,N_3912,N_3378);
nor U4521 (N_4521,N_2014,N_2550);
and U4522 (N_4522,N_3775,N_2807);
or U4523 (N_4523,N_2539,N_2749);
nor U4524 (N_4524,N_2121,N_2886);
and U4525 (N_4525,N_3049,N_3909);
nor U4526 (N_4526,N_3676,N_3779);
and U4527 (N_4527,N_2532,N_2526);
and U4528 (N_4528,N_2079,N_2505);
and U4529 (N_4529,N_2722,N_2495);
or U4530 (N_4530,N_3638,N_2738);
nor U4531 (N_4531,N_3856,N_2527);
and U4532 (N_4532,N_2875,N_3836);
or U4533 (N_4533,N_2768,N_2699);
and U4534 (N_4534,N_3262,N_2649);
and U4535 (N_4535,N_2803,N_3686);
nor U4536 (N_4536,N_3568,N_2951);
nor U4537 (N_4537,N_3158,N_2838);
and U4538 (N_4538,N_2761,N_2076);
and U4539 (N_4539,N_3211,N_2696);
nand U4540 (N_4540,N_2498,N_3264);
nor U4541 (N_4541,N_3420,N_3630);
nand U4542 (N_4542,N_2154,N_3684);
nor U4543 (N_4543,N_3502,N_3277);
or U4544 (N_4544,N_3363,N_3195);
and U4545 (N_4545,N_3067,N_2937);
and U4546 (N_4546,N_3578,N_3295);
or U4547 (N_4547,N_3854,N_3451);
and U4548 (N_4548,N_3953,N_3598);
nand U4549 (N_4549,N_3955,N_2071);
and U4550 (N_4550,N_3888,N_2988);
nand U4551 (N_4551,N_2610,N_3974);
nor U4552 (N_4552,N_2741,N_3928);
nand U4553 (N_4553,N_2924,N_2870);
nor U4554 (N_4554,N_2366,N_3369);
nand U4555 (N_4555,N_2514,N_2192);
or U4556 (N_4556,N_3680,N_3528);
or U4557 (N_4557,N_2110,N_3954);
nor U4558 (N_4558,N_3402,N_3604);
nand U4559 (N_4559,N_2730,N_2727);
xor U4560 (N_4560,N_3597,N_3771);
or U4561 (N_4561,N_3204,N_3128);
nand U4562 (N_4562,N_2715,N_2132);
and U4563 (N_4563,N_3090,N_2939);
nand U4564 (N_4564,N_3555,N_2549);
and U4565 (N_4565,N_2834,N_3442);
nand U4566 (N_4566,N_3151,N_3956);
nand U4567 (N_4567,N_2909,N_3875);
or U4568 (N_4568,N_2019,N_3187);
nand U4569 (N_4569,N_3301,N_3720);
or U4570 (N_4570,N_2089,N_3747);
or U4571 (N_4571,N_2108,N_3366);
or U4572 (N_4572,N_3485,N_3285);
nor U4573 (N_4573,N_2094,N_2973);
or U4574 (N_4574,N_3086,N_3714);
nor U4575 (N_4575,N_3944,N_2465);
nor U4576 (N_4576,N_3612,N_3200);
and U4577 (N_4577,N_2508,N_2151);
nand U4578 (N_4578,N_2888,N_2137);
nor U4579 (N_4579,N_2938,N_2970);
or U4580 (N_4580,N_2917,N_3443);
xor U4581 (N_4581,N_2644,N_3400);
or U4582 (N_4582,N_3150,N_2797);
nor U4583 (N_4583,N_3605,N_2635);
nand U4584 (N_4584,N_3607,N_3627);
or U4585 (N_4585,N_3003,N_2997);
nand U4586 (N_4586,N_2833,N_3536);
and U4587 (N_4587,N_2394,N_3826);
or U4588 (N_4588,N_2033,N_3900);
nor U4589 (N_4589,N_3551,N_3534);
and U4590 (N_4590,N_2887,N_3993);
nor U4591 (N_4591,N_3760,N_2034);
nand U4592 (N_4592,N_3007,N_3600);
nor U4593 (N_4593,N_2074,N_3791);
and U4594 (N_4594,N_3687,N_2579);
nand U4595 (N_4595,N_2513,N_2138);
nand U4596 (N_4596,N_2295,N_2031);
or U4597 (N_4597,N_2102,N_3482);
xnor U4598 (N_4598,N_3042,N_3015);
and U4599 (N_4599,N_3168,N_3221);
nand U4600 (N_4600,N_3699,N_3240);
xor U4601 (N_4601,N_3303,N_3322);
nand U4602 (N_4602,N_3715,N_2287);
and U4603 (N_4603,N_2222,N_3190);
or U4604 (N_4604,N_3464,N_2619);
xor U4605 (N_4605,N_2450,N_3521);
nor U4606 (N_4606,N_3157,N_3742);
nand U4607 (N_4607,N_3516,N_3120);
nand U4608 (N_4608,N_3839,N_3705);
or U4609 (N_4609,N_3370,N_3822);
or U4610 (N_4610,N_3014,N_3281);
and U4611 (N_4611,N_3834,N_2791);
xor U4612 (N_4612,N_3479,N_2046);
nand U4613 (N_4613,N_2548,N_3609);
or U4614 (N_4614,N_2447,N_2760);
or U4615 (N_4615,N_2375,N_2461);
nand U4616 (N_4616,N_2186,N_3403);
nor U4617 (N_4617,N_3109,N_3212);
and U4618 (N_4618,N_2322,N_3758);
and U4619 (N_4619,N_2948,N_3652);
nor U4620 (N_4620,N_2052,N_3979);
nand U4621 (N_4621,N_3594,N_2828);
and U4622 (N_4622,N_2874,N_2518);
nor U4623 (N_4623,N_3326,N_3916);
or U4624 (N_4624,N_2230,N_2798);
nor U4625 (N_4625,N_2710,N_3711);
nor U4626 (N_4626,N_2554,N_3352);
nor U4627 (N_4627,N_2947,N_2410);
nor U4628 (N_4628,N_3983,N_3697);
or U4629 (N_4629,N_2878,N_3468);
nor U4630 (N_4630,N_3884,N_2458);
nand U4631 (N_4631,N_2482,N_3066);
nor U4632 (N_4632,N_2903,N_3906);
and U4633 (N_4633,N_2185,N_2863);
nor U4634 (N_4634,N_3082,N_3398);
nor U4635 (N_4635,N_3852,N_2246);
nor U4636 (N_4636,N_3910,N_2320);
nand U4637 (N_4637,N_3390,N_3358);
nor U4638 (N_4638,N_2721,N_2934);
nand U4639 (N_4639,N_2060,N_3660);
nand U4640 (N_4640,N_2265,N_3012);
nor U4641 (N_4641,N_3401,N_3392);
and U4642 (N_4642,N_2275,N_2669);
or U4643 (N_4643,N_2143,N_3435);
nor U4644 (N_4644,N_2812,N_3224);
or U4645 (N_4645,N_3723,N_3074);
nand U4646 (N_4646,N_3500,N_3820);
nand U4647 (N_4647,N_2231,N_3294);
nor U4648 (N_4648,N_2489,N_3222);
or U4649 (N_4649,N_3991,N_2979);
and U4650 (N_4650,N_2315,N_3445);
and U4651 (N_4651,N_2616,N_2303);
and U4652 (N_4652,N_3106,N_3131);
and U4653 (N_4653,N_2374,N_3460);
nor U4654 (N_4654,N_2712,N_3114);
and U4655 (N_4655,N_3978,N_2389);
or U4656 (N_4656,N_3310,N_3251);
or U4657 (N_4657,N_3026,N_3803);
nand U4658 (N_4658,N_3659,N_2395);
nor U4659 (N_4659,N_3707,N_2977);
or U4660 (N_4660,N_2726,N_3115);
or U4661 (N_4661,N_2884,N_2276);
nor U4662 (N_4662,N_2497,N_3357);
nor U4663 (N_4663,N_3348,N_2196);
nand U4664 (N_4664,N_3582,N_3880);
nand U4665 (N_4665,N_3321,N_3463);
nor U4666 (N_4666,N_2118,N_2671);
nand U4667 (N_4667,N_2502,N_3985);
and U4668 (N_4668,N_3235,N_2240);
and U4669 (N_4669,N_2529,N_2849);
nand U4670 (N_4670,N_3474,N_2995);
nand U4671 (N_4671,N_2204,N_3182);
nor U4672 (N_4672,N_2406,N_2678);
nor U4673 (N_4673,N_2750,N_2872);
nand U4674 (N_4674,N_2755,N_3628);
nor U4675 (N_4675,N_2160,N_3020);
or U4676 (N_4676,N_3710,N_2336);
nor U4677 (N_4677,N_3958,N_2781);
nor U4678 (N_4678,N_3426,N_3608);
and U4679 (N_4679,N_2083,N_2561);
nand U4680 (N_4680,N_2844,N_3739);
or U4681 (N_4681,N_3490,N_3489);
nor U4682 (N_4682,N_2958,N_2248);
and U4683 (N_4683,N_2630,N_2073);
or U4684 (N_4684,N_2117,N_3210);
nand U4685 (N_4685,N_2689,N_3466);
nor U4686 (N_4686,N_2583,N_3266);
nand U4687 (N_4687,N_3419,N_3183);
nor U4688 (N_4688,N_2568,N_2871);
nor U4689 (N_4689,N_3342,N_2176);
nand U4690 (N_4690,N_2962,N_2652);
nor U4691 (N_4691,N_2836,N_2774);
nand U4692 (N_4692,N_2402,N_3624);
or U4693 (N_4693,N_2473,N_2171);
nand U4694 (N_4694,N_3318,N_3347);
or U4695 (N_4695,N_2142,N_3456);
or U4696 (N_4696,N_2398,N_2397);
or U4697 (N_4697,N_3862,N_2819);
and U4698 (N_4698,N_2900,N_2589);
or U4699 (N_4699,N_3662,N_3017);
nor U4700 (N_4700,N_3616,N_2039);
or U4701 (N_4701,N_2382,N_3317);
nand U4702 (N_4702,N_2023,N_2384);
nor U4703 (N_4703,N_2165,N_3835);
and U4704 (N_4704,N_2927,N_2364);
nor U4705 (N_4705,N_2134,N_2494);
nor U4706 (N_4706,N_3252,N_3306);
nor U4707 (N_4707,N_3892,N_2896);
nand U4708 (N_4708,N_3417,N_3282);
or U4709 (N_4709,N_3088,N_3031);
nand U4710 (N_4710,N_3644,N_3811);
and U4711 (N_4711,N_3177,N_2446);
nand U4712 (N_4712,N_2127,N_3124);
nand U4713 (N_4713,N_2861,N_3149);
nor U4714 (N_4714,N_3877,N_3524);
nor U4715 (N_4715,N_2405,N_2018);
or U4716 (N_4716,N_3422,N_3709);
and U4717 (N_4717,N_3215,N_2890);
nor U4718 (N_4718,N_2147,N_2181);
nand U4719 (N_4719,N_2408,N_3768);
and U4720 (N_4720,N_2189,N_3278);
and U4721 (N_4721,N_2617,N_2684);
or U4722 (N_4722,N_2291,N_2679);
and U4723 (N_4723,N_3584,N_2810);
nand U4724 (N_4724,N_2697,N_2302);
and U4725 (N_4725,N_2162,N_3858);
nand U4726 (N_4726,N_2370,N_2793);
and U4727 (N_4727,N_3572,N_2706);
nand U4728 (N_4728,N_3575,N_3155);
and U4729 (N_4729,N_3654,N_2576);
nand U4730 (N_4730,N_3671,N_3101);
nand U4731 (N_4731,N_2601,N_3593);
or U4732 (N_4732,N_2582,N_2932);
nand U4733 (N_4733,N_3141,N_2916);
nor U4734 (N_4734,N_3788,N_2197);
nor U4735 (N_4735,N_3415,N_3620);
nand U4736 (N_4736,N_3383,N_2459);
nand U4737 (N_4737,N_2455,N_3372);
nor U4738 (N_4738,N_2305,N_3389);
or U4739 (N_4739,N_3315,N_3782);
or U4740 (N_4740,N_3273,N_3176);
or U4741 (N_4741,N_2000,N_3198);
nand U4742 (N_4742,N_2002,N_2707);
nand U4743 (N_4743,N_2184,N_2984);
nand U4744 (N_4744,N_2864,N_3142);
and U4745 (N_4745,N_3069,N_3674);
nor U4746 (N_4746,N_2804,N_3343);
or U4747 (N_4747,N_2748,N_2852);
and U4748 (N_4748,N_2201,N_3561);
and U4749 (N_4749,N_2972,N_2775);
nand U4750 (N_4750,N_3812,N_2157);
and U4751 (N_4751,N_2996,N_3078);
and U4752 (N_4752,N_2971,N_2591);
nor U4753 (N_4753,N_2949,N_3621);
nor U4754 (N_4754,N_3208,N_2332);
and U4755 (N_4755,N_3471,N_2643);
nand U4756 (N_4756,N_2891,N_2257);
xnor U4757 (N_4757,N_2620,N_2594);
xor U4758 (N_4758,N_2285,N_2335);
and U4759 (N_4759,N_2342,N_2311);
nor U4760 (N_4760,N_2598,N_2416);
nand U4761 (N_4761,N_2493,N_2278);
nand U4762 (N_4762,N_2167,N_2789);
or U4763 (N_4763,N_3314,N_3679);
nand U4764 (N_4764,N_2574,N_3391);
nor U4765 (N_4765,N_3360,N_2639);
nor U4766 (N_4766,N_3846,N_3234);
nand U4767 (N_4767,N_3648,N_2438);
nor U4768 (N_4768,N_3651,N_2082);
nor U4769 (N_4769,N_3112,N_2544);
and U4770 (N_4770,N_2690,N_3997);
nand U4771 (N_4771,N_3550,N_3987);
nand U4772 (N_4772,N_2166,N_2879);
and U4773 (N_4773,N_2624,N_3764);
or U4774 (N_4774,N_3433,N_2736);
or U4775 (N_4775,N_3231,N_2926);
nor U4776 (N_4776,N_3172,N_2286);
and U4777 (N_4777,N_3276,N_3484);
nor U4778 (N_4778,N_2717,N_3641);
and U4779 (N_4779,N_2588,N_3899);
or U4780 (N_4780,N_3513,N_3205);
or U4781 (N_4781,N_3011,N_2351);
nand U4782 (N_4782,N_3405,N_2200);
or U4783 (N_4783,N_3220,N_2090);
or U4784 (N_4784,N_3072,N_3790);
nand U4785 (N_4785,N_2724,N_2492);
nand U4786 (N_4786,N_3296,N_2655);
or U4787 (N_4787,N_2324,N_2419);
nor U4788 (N_4788,N_3345,N_2116);
or U4789 (N_4789,N_3181,N_3189);
nor U4790 (N_4790,N_3228,N_3799);
and U4791 (N_4791,N_3194,N_2203);
and U4792 (N_4792,N_2739,N_3737);
and U4793 (N_4793,N_3975,N_2413);
nand U4794 (N_4794,N_2443,N_3787);
or U4795 (N_4795,N_2418,N_2268);
or U4796 (N_4796,N_2454,N_3693);
and U4797 (N_4797,N_2329,N_2393);
and U4798 (N_4798,N_2866,N_3547);
and U4799 (N_4799,N_2421,N_3161);
or U4800 (N_4800,N_2124,N_2965);
or U4801 (N_4801,N_3570,N_3138);
nand U4802 (N_4802,N_2705,N_3665);
nand U4803 (N_4803,N_3850,N_3395);
nand U4804 (N_4804,N_2935,N_2028);
nor U4805 (N_4805,N_3410,N_2403);
nand U4806 (N_4806,N_3895,N_2578);
and U4807 (N_4807,N_3595,N_3925);
nor U4808 (N_4808,N_3028,N_2012);
nand U4809 (N_4809,N_3430,N_3962);
nor U4810 (N_4810,N_3267,N_2352);
or U4811 (N_4811,N_2824,N_2478);
nor U4812 (N_4812,N_2220,N_3847);
or U4813 (N_4813,N_2967,N_3738);
nand U4814 (N_4814,N_2290,N_2577);
and U4815 (N_4815,N_2795,N_2651);
nand U4816 (N_4816,N_3703,N_3274);
or U4817 (N_4817,N_3695,N_3232);
nand U4818 (N_4818,N_3412,N_3726);
or U4819 (N_4819,N_2235,N_3432);
nand U4820 (N_4820,N_2216,N_3135);
nor U4821 (N_4821,N_2067,N_3808);
or U4822 (N_4822,N_2109,N_2304);
and U4823 (N_4823,N_3029,N_2049);
or U4824 (N_4824,N_2453,N_2914);
nor U4825 (N_4825,N_2259,N_3924);
nand U4826 (N_4826,N_2479,N_3293);
or U4827 (N_4827,N_3024,N_3027);
xor U4828 (N_4828,N_3311,N_3514);
and U4829 (N_4829,N_3581,N_2035);
and U4830 (N_4830,N_2509,N_2041);
or U4831 (N_4831,N_3290,N_3861);
and U4832 (N_4832,N_3238,N_2284);
and U4833 (N_4833,N_2551,N_3920);
nor U4834 (N_4834,N_2442,N_2449);
nand U4835 (N_4835,N_2784,N_2061);
or U4836 (N_4836,N_2070,N_2832);
and U4837 (N_4837,N_2912,N_2525);
nor U4838 (N_4838,N_2968,N_2146);
nor U4839 (N_4839,N_2587,N_2158);
and U4840 (N_4840,N_2377,N_3271);
nor U4841 (N_4841,N_2038,N_3254);
nand U4842 (N_4842,N_3815,N_2581);
or U4843 (N_4843,N_2792,N_3780);
nor U4844 (N_4844,N_3913,N_2956);
and U4845 (N_4845,N_2898,N_3995);
nand U4846 (N_4846,N_2711,N_3744);
and U4847 (N_4847,N_2735,N_2637);
and U4848 (N_4848,N_3449,N_3236);
nor U4849 (N_4849,N_2763,N_3919);
or U4850 (N_4850,N_2847,N_2273);
and U4851 (N_4851,N_3367,N_3346);
and U4852 (N_4852,N_3154,N_2931);
and U4853 (N_4853,N_2504,N_2656);
and U4854 (N_4854,N_3388,N_3444);
nand U4855 (N_4855,N_3461,N_2123);
nand U4856 (N_4856,N_2599,N_2522);
nand U4857 (N_4857,N_2463,N_3564);
or U4858 (N_4858,N_3959,N_2822);
nand U4859 (N_4859,N_3646,N_2251);
nand U4860 (N_4860,N_3202,N_3819);
nand U4861 (N_4861,N_2963,N_3039);
nor U4862 (N_4862,N_2845,N_2904);
or U4863 (N_4863,N_2024,N_3121);
and U4864 (N_4864,N_2515,N_3664);
nand U4865 (N_4865,N_2882,N_2367);
nor U4866 (N_4866,N_2565,N_2989);
nand U4867 (N_4867,N_3756,N_2758);
or U4868 (N_4868,N_3963,N_3289);
or U4869 (N_4869,N_2245,N_3713);
nand U4870 (N_4870,N_3214,N_2955);
nand U4871 (N_4871,N_2093,N_3511);
nor U4872 (N_4872,N_3494,N_3219);
and U4873 (N_4873,N_3481,N_3650);
nand U4874 (N_4874,N_3789,N_3683);
nand U4875 (N_4875,N_2174,N_2068);
xor U4876 (N_4876,N_3334,N_2212);
or U4877 (N_4877,N_2673,N_3878);
or U4878 (N_4878,N_3312,N_2694);
nand U4879 (N_4879,N_2604,N_3050);
or U4880 (N_4880,N_3283,N_3113);
or U4881 (N_4881,N_2401,N_3414);
and U4882 (N_4882,N_3733,N_3640);
and U4883 (N_4883,N_3056,N_2681);
and U4884 (N_4884,N_2702,N_2813);
nand U4885 (N_4885,N_3075,N_2371);
nand U4886 (N_4886,N_3043,N_3755);
and U4887 (N_4887,N_2422,N_3428);
and U4888 (N_4888,N_3013,N_2843);
and U4889 (N_4889,N_2547,N_3099);
and U4890 (N_4890,N_2704,N_2261);
and U4891 (N_4891,N_3813,N_2992);
and U4892 (N_4892,N_2503,N_2299);
and U4893 (N_4893,N_3080,N_3191);
or U4894 (N_4894,N_2873,N_2300);
nor U4895 (N_4895,N_3448,N_3801);
nand U4896 (N_4896,N_3698,N_3905);
and U4897 (N_4897,N_2670,N_3376);
and U4898 (N_4898,N_3239,N_2883);
nor U4899 (N_4899,N_2238,N_3968);
nor U4900 (N_4900,N_3033,N_2535);
nor U4901 (N_4901,N_3440,N_2170);
and U4902 (N_4902,N_2570,N_2319);
nor U4903 (N_4903,N_2686,N_2907);
and U4904 (N_4904,N_2057,N_2894);
and U4905 (N_4905,N_2228,N_2854);
or U4906 (N_4906,N_2500,N_2606);
nor U4907 (N_4907,N_3437,N_3688);
nand U4908 (N_4908,N_3411,N_2407);
nor U4909 (N_4909,N_3038,N_2658);
nand U4910 (N_4910,N_2910,N_2999);
nand U4911 (N_4911,N_3382,N_2731);
nor U4912 (N_4912,N_2307,N_3477);
nor U4913 (N_4913,N_2435,N_2668);
nor U4914 (N_4914,N_2316,N_3785);
and U4915 (N_4915,N_2069,N_3493);
nor U4916 (N_4916,N_3941,N_2533);
and U4917 (N_4917,N_3058,N_2253);
nand U4918 (N_4918,N_3749,N_3512);
or U4919 (N_4919,N_3793,N_2331);
nor U4920 (N_4920,N_2487,N_2940);
and U4921 (N_4921,N_3840,N_2107);
xnor U4922 (N_4922,N_3583,N_2262);
and U4923 (N_4923,N_2025,N_3136);
nand U4924 (N_4924,N_3375,N_3515);
and U4925 (N_4925,N_2608,N_2373);
and U4926 (N_4926,N_2754,N_3325);
or U4927 (N_4927,N_3156,N_2632);
and U4928 (N_4928,N_3532,N_3040);
or U4929 (N_4929,N_3864,N_3469);
and U4930 (N_4930,N_3453,N_3196);
and U4931 (N_4931,N_3000,N_2098);
nand U4932 (N_4932,N_2190,N_3548);
nand U4933 (N_4933,N_3284,N_3045);
and U4934 (N_4934,N_3163,N_3863);
nand U4935 (N_4935,N_3889,N_3557);
nand U4936 (N_4936,N_2078,N_3585);
nand U4937 (N_4937,N_2708,N_3545);
nand U4938 (N_4938,N_3184,N_2213);
nand U4939 (N_4939,N_3921,N_3499);
and U4940 (N_4940,N_3566,N_3692);
and U4941 (N_4941,N_3253,N_3970);
nor U4942 (N_4942,N_3319,N_2837);
or U4943 (N_4943,N_2045,N_2728);
nor U4944 (N_4944,N_3242,N_2239);
nand U4945 (N_4945,N_3655,N_2007);
or U4946 (N_4946,N_2417,N_2379);
nor U4947 (N_4947,N_2831,N_2636);
and U4948 (N_4948,N_3669,N_2944);
nor U4949 (N_4949,N_3503,N_2159);
and U4950 (N_4950,N_2933,N_2086);
or U4951 (N_4951,N_2519,N_2779);
and U4952 (N_4952,N_2353,N_2059);
or U4953 (N_4953,N_2718,N_3702);
nand U4954 (N_4954,N_3734,N_3287);
and U4955 (N_4955,N_3930,N_3891);
nor U4956 (N_4956,N_2523,N_3125);
nand U4957 (N_4957,N_3610,N_2809);
nor U4958 (N_4958,N_3046,N_2125);
and U4959 (N_4959,N_3772,N_3786);
and U4960 (N_4960,N_3134,N_3406);
or U4961 (N_4961,N_3961,N_2719);
and U4962 (N_4962,N_3421,N_2647);
nand U4963 (N_4963,N_2277,N_3001);
or U4964 (N_4964,N_3192,N_2017);
and U4965 (N_4965,N_2980,N_3588);
or U4966 (N_4966,N_3943,N_3373);
nor U4967 (N_4967,N_3631,N_3903);
nand U4968 (N_4968,N_2975,N_3006);
nor U4969 (N_4969,N_2595,N_3969);
and U4970 (N_4970,N_2640,N_2943);
nand U4971 (N_4971,N_3385,N_3971);
nand U4972 (N_4972,N_3810,N_2187);
and U4973 (N_4973,N_3927,N_3431);
nand U4974 (N_4974,N_2430,N_3988);
and U4975 (N_4975,N_3635,N_3675);
and U4976 (N_4976,N_3677,N_2780);
and U4977 (N_4977,N_3960,N_3871);
nand U4978 (N_4978,N_2592,N_2349);
nor U4979 (N_4979,N_2385,N_2716);
nand U4980 (N_4980,N_3816,N_2451);
nor U4981 (N_4981,N_2737,N_3984);
or U4982 (N_4982,N_2168,N_2667);
and U4983 (N_4983,N_2140,N_3100);
nand U4984 (N_4984,N_2427,N_2359);
nor U4985 (N_4985,N_2129,N_2149);
nand U4986 (N_4986,N_2298,N_3591);
or U4987 (N_4987,N_3973,N_3672);
nand U4988 (N_4988,N_3413,N_2650);
xnor U4989 (N_4989,N_3883,N_2692);
nor U4990 (N_4990,N_3633,N_3117);
nor U4991 (N_4991,N_2990,N_3048);
nand U4992 (N_4992,N_2036,N_3890);
nand U4993 (N_4993,N_3549,N_2575);
nand U4994 (N_4994,N_2998,N_2365);
or U4995 (N_4995,N_3623,N_2144);
nor U4996 (N_4996,N_2051,N_3458);
nor U4997 (N_4997,N_2145,N_3559);
and U4998 (N_4998,N_3519,N_2985);
nand U4999 (N_4999,N_2312,N_3025);
or U5000 (N_5000,N_2907,N_3325);
nand U5001 (N_5001,N_2658,N_3984);
or U5002 (N_5002,N_3514,N_3735);
or U5003 (N_5003,N_3633,N_2270);
or U5004 (N_5004,N_3690,N_2768);
nand U5005 (N_5005,N_3544,N_2640);
nand U5006 (N_5006,N_3163,N_3723);
and U5007 (N_5007,N_2786,N_3637);
or U5008 (N_5008,N_2882,N_3721);
and U5009 (N_5009,N_3077,N_2709);
nor U5010 (N_5010,N_3908,N_2866);
or U5011 (N_5011,N_3202,N_2409);
nor U5012 (N_5012,N_3523,N_2076);
nor U5013 (N_5013,N_2854,N_2042);
and U5014 (N_5014,N_2623,N_2154);
or U5015 (N_5015,N_3191,N_3176);
or U5016 (N_5016,N_3582,N_2746);
nand U5017 (N_5017,N_2272,N_3828);
nand U5018 (N_5018,N_3822,N_2697);
nor U5019 (N_5019,N_2528,N_3328);
and U5020 (N_5020,N_3210,N_2969);
nor U5021 (N_5021,N_2684,N_2066);
nand U5022 (N_5022,N_3169,N_3758);
nor U5023 (N_5023,N_3973,N_2063);
or U5024 (N_5024,N_2210,N_3119);
nand U5025 (N_5025,N_3800,N_2625);
or U5026 (N_5026,N_3253,N_3477);
or U5027 (N_5027,N_2074,N_3904);
or U5028 (N_5028,N_3789,N_3500);
or U5029 (N_5029,N_3142,N_2152);
nor U5030 (N_5030,N_2782,N_2635);
or U5031 (N_5031,N_3229,N_3621);
and U5032 (N_5032,N_3668,N_3688);
and U5033 (N_5033,N_3326,N_2613);
and U5034 (N_5034,N_2111,N_3634);
nand U5035 (N_5035,N_3521,N_3919);
nor U5036 (N_5036,N_2951,N_2001);
nand U5037 (N_5037,N_2471,N_3503);
or U5038 (N_5038,N_2483,N_2199);
or U5039 (N_5039,N_2666,N_2402);
nand U5040 (N_5040,N_3754,N_2548);
nor U5041 (N_5041,N_3944,N_3403);
nand U5042 (N_5042,N_2172,N_3711);
and U5043 (N_5043,N_3995,N_2240);
nor U5044 (N_5044,N_3059,N_2592);
nand U5045 (N_5045,N_2579,N_3717);
or U5046 (N_5046,N_3434,N_3968);
nand U5047 (N_5047,N_3774,N_3918);
and U5048 (N_5048,N_3616,N_2398);
nor U5049 (N_5049,N_2862,N_3308);
nand U5050 (N_5050,N_3693,N_3232);
nand U5051 (N_5051,N_2649,N_2546);
and U5052 (N_5052,N_3894,N_3160);
nor U5053 (N_5053,N_2769,N_3794);
nor U5054 (N_5054,N_2099,N_3251);
and U5055 (N_5055,N_2784,N_3874);
or U5056 (N_5056,N_2425,N_3061);
or U5057 (N_5057,N_3525,N_2038);
and U5058 (N_5058,N_2782,N_3182);
or U5059 (N_5059,N_3793,N_2671);
nand U5060 (N_5060,N_2883,N_2006);
and U5061 (N_5061,N_2958,N_2715);
and U5062 (N_5062,N_3354,N_3043);
and U5063 (N_5063,N_3041,N_2971);
and U5064 (N_5064,N_3699,N_2656);
nor U5065 (N_5065,N_2054,N_3005);
nand U5066 (N_5066,N_3413,N_3537);
nand U5067 (N_5067,N_3799,N_3618);
nand U5068 (N_5068,N_2454,N_3971);
and U5069 (N_5069,N_3880,N_3175);
nand U5070 (N_5070,N_3443,N_3274);
nor U5071 (N_5071,N_3033,N_3281);
or U5072 (N_5072,N_3982,N_3838);
or U5073 (N_5073,N_2611,N_3802);
and U5074 (N_5074,N_2293,N_3658);
nor U5075 (N_5075,N_3463,N_2523);
nand U5076 (N_5076,N_2372,N_3544);
or U5077 (N_5077,N_3146,N_2358);
nand U5078 (N_5078,N_3235,N_2023);
or U5079 (N_5079,N_2030,N_2044);
nor U5080 (N_5080,N_3394,N_2648);
or U5081 (N_5081,N_3917,N_2255);
or U5082 (N_5082,N_3726,N_2072);
and U5083 (N_5083,N_2655,N_3502);
nor U5084 (N_5084,N_3064,N_2760);
nor U5085 (N_5085,N_3461,N_2870);
nor U5086 (N_5086,N_2297,N_2685);
or U5087 (N_5087,N_3219,N_2363);
xnor U5088 (N_5088,N_3566,N_3128);
or U5089 (N_5089,N_2134,N_2937);
or U5090 (N_5090,N_3158,N_3268);
or U5091 (N_5091,N_3396,N_2764);
or U5092 (N_5092,N_2762,N_3022);
nand U5093 (N_5093,N_2254,N_3919);
or U5094 (N_5094,N_3097,N_3416);
nand U5095 (N_5095,N_3965,N_2904);
nor U5096 (N_5096,N_3177,N_2049);
or U5097 (N_5097,N_2668,N_2734);
nor U5098 (N_5098,N_2685,N_2665);
and U5099 (N_5099,N_2722,N_3673);
nand U5100 (N_5100,N_3643,N_2500);
nor U5101 (N_5101,N_2898,N_2038);
nor U5102 (N_5102,N_3423,N_2862);
nand U5103 (N_5103,N_3445,N_2296);
nand U5104 (N_5104,N_3833,N_3792);
or U5105 (N_5105,N_3161,N_3697);
and U5106 (N_5106,N_2437,N_2340);
nand U5107 (N_5107,N_2209,N_3572);
or U5108 (N_5108,N_3265,N_3888);
or U5109 (N_5109,N_2108,N_3820);
nand U5110 (N_5110,N_3432,N_2931);
and U5111 (N_5111,N_2652,N_2386);
or U5112 (N_5112,N_2106,N_3961);
and U5113 (N_5113,N_3316,N_2154);
nand U5114 (N_5114,N_2649,N_2177);
or U5115 (N_5115,N_2836,N_2332);
or U5116 (N_5116,N_3455,N_3151);
or U5117 (N_5117,N_3564,N_3842);
and U5118 (N_5118,N_3427,N_2601);
or U5119 (N_5119,N_2404,N_3697);
or U5120 (N_5120,N_3502,N_3468);
nor U5121 (N_5121,N_3568,N_3165);
or U5122 (N_5122,N_3580,N_3335);
and U5123 (N_5123,N_2650,N_3965);
nand U5124 (N_5124,N_2368,N_3856);
nor U5125 (N_5125,N_3085,N_2673);
nand U5126 (N_5126,N_2216,N_2265);
nand U5127 (N_5127,N_2286,N_3367);
and U5128 (N_5128,N_3034,N_3383);
nor U5129 (N_5129,N_2684,N_3018);
nor U5130 (N_5130,N_2976,N_3824);
nand U5131 (N_5131,N_3322,N_2327);
nor U5132 (N_5132,N_2794,N_2542);
nor U5133 (N_5133,N_3844,N_3950);
nor U5134 (N_5134,N_3970,N_2627);
and U5135 (N_5135,N_2074,N_3347);
xor U5136 (N_5136,N_3583,N_3798);
or U5137 (N_5137,N_3186,N_2569);
nor U5138 (N_5138,N_3201,N_3182);
and U5139 (N_5139,N_3540,N_3851);
or U5140 (N_5140,N_3412,N_2712);
or U5141 (N_5141,N_3420,N_3993);
nor U5142 (N_5142,N_3990,N_3047);
or U5143 (N_5143,N_3273,N_3801);
and U5144 (N_5144,N_2392,N_2010);
xnor U5145 (N_5145,N_2172,N_3071);
or U5146 (N_5146,N_2924,N_2672);
nand U5147 (N_5147,N_2157,N_2247);
nand U5148 (N_5148,N_3616,N_2293);
nor U5149 (N_5149,N_2789,N_3863);
and U5150 (N_5150,N_3389,N_2339);
nor U5151 (N_5151,N_3809,N_2199);
or U5152 (N_5152,N_3872,N_2309);
nor U5153 (N_5153,N_3357,N_3535);
or U5154 (N_5154,N_3847,N_3477);
nand U5155 (N_5155,N_3474,N_3890);
nand U5156 (N_5156,N_2415,N_2849);
nor U5157 (N_5157,N_3061,N_2591);
nor U5158 (N_5158,N_2647,N_3268);
and U5159 (N_5159,N_3852,N_2376);
and U5160 (N_5160,N_2250,N_3314);
and U5161 (N_5161,N_2766,N_3099);
or U5162 (N_5162,N_3344,N_2677);
or U5163 (N_5163,N_2722,N_3203);
or U5164 (N_5164,N_3344,N_3836);
or U5165 (N_5165,N_2143,N_3675);
nand U5166 (N_5166,N_2260,N_3565);
or U5167 (N_5167,N_3619,N_3933);
nand U5168 (N_5168,N_3521,N_3396);
nand U5169 (N_5169,N_2975,N_2516);
nand U5170 (N_5170,N_3972,N_3017);
and U5171 (N_5171,N_3807,N_3071);
nand U5172 (N_5172,N_3398,N_3543);
nor U5173 (N_5173,N_3048,N_3474);
or U5174 (N_5174,N_3737,N_3976);
or U5175 (N_5175,N_2519,N_2932);
nand U5176 (N_5176,N_3730,N_2487);
and U5177 (N_5177,N_3189,N_2833);
or U5178 (N_5178,N_2823,N_2235);
or U5179 (N_5179,N_2476,N_2706);
or U5180 (N_5180,N_2439,N_3073);
or U5181 (N_5181,N_2840,N_3520);
nor U5182 (N_5182,N_3801,N_2880);
or U5183 (N_5183,N_2105,N_3354);
nand U5184 (N_5184,N_2507,N_3775);
nor U5185 (N_5185,N_2903,N_3858);
nand U5186 (N_5186,N_3606,N_2470);
or U5187 (N_5187,N_3385,N_2094);
and U5188 (N_5188,N_2305,N_3530);
nand U5189 (N_5189,N_2831,N_2323);
and U5190 (N_5190,N_2923,N_3763);
and U5191 (N_5191,N_2501,N_3774);
nand U5192 (N_5192,N_2249,N_3602);
and U5193 (N_5193,N_3991,N_3202);
or U5194 (N_5194,N_3429,N_2816);
nor U5195 (N_5195,N_3046,N_2637);
or U5196 (N_5196,N_2613,N_2162);
or U5197 (N_5197,N_2002,N_3188);
or U5198 (N_5198,N_3731,N_2490);
and U5199 (N_5199,N_3603,N_2055);
or U5200 (N_5200,N_3832,N_2389);
and U5201 (N_5201,N_2523,N_2203);
or U5202 (N_5202,N_3806,N_2713);
nand U5203 (N_5203,N_3684,N_2948);
or U5204 (N_5204,N_2672,N_2115);
nor U5205 (N_5205,N_3121,N_3748);
or U5206 (N_5206,N_3792,N_2696);
nand U5207 (N_5207,N_2675,N_2491);
and U5208 (N_5208,N_2795,N_2259);
nor U5209 (N_5209,N_3269,N_3804);
and U5210 (N_5210,N_3430,N_3794);
nor U5211 (N_5211,N_3160,N_3366);
nor U5212 (N_5212,N_2138,N_3302);
or U5213 (N_5213,N_2546,N_3229);
nor U5214 (N_5214,N_2040,N_3104);
and U5215 (N_5215,N_2458,N_2059);
nor U5216 (N_5216,N_2972,N_2280);
nand U5217 (N_5217,N_3227,N_2142);
or U5218 (N_5218,N_3529,N_3219);
nand U5219 (N_5219,N_3788,N_3766);
nor U5220 (N_5220,N_3232,N_2593);
nor U5221 (N_5221,N_3090,N_2551);
xnor U5222 (N_5222,N_2606,N_2944);
or U5223 (N_5223,N_2732,N_3527);
nand U5224 (N_5224,N_3804,N_3076);
or U5225 (N_5225,N_3102,N_2304);
or U5226 (N_5226,N_2379,N_2684);
or U5227 (N_5227,N_2726,N_3072);
or U5228 (N_5228,N_3558,N_2014);
or U5229 (N_5229,N_2904,N_3191);
and U5230 (N_5230,N_2710,N_2801);
nand U5231 (N_5231,N_2462,N_3837);
or U5232 (N_5232,N_2423,N_2316);
nor U5233 (N_5233,N_3398,N_3792);
and U5234 (N_5234,N_2953,N_2323);
or U5235 (N_5235,N_3026,N_2236);
or U5236 (N_5236,N_3704,N_3185);
and U5237 (N_5237,N_3679,N_2285);
and U5238 (N_5238,N_2891,N_3177);
nor U5239 (N_5239,N_3469,N_3870);
and U5240 (N_5240,N_3869,N_3433);
nor U5241 (N_5241,N_2418,N_2625);
and U5242 (N_5242,N_2562,N_3419);
and U5243 (N_5243,N_3805,N_3535);
or U5244 (N_5244,N_3266,N_3466);
or U5245 (N_5245,N_3914,N_2113);
nand U5246 (N_5246,N_2567,N_3417);
nor U5247 (N_5247,N_2733,N_2297);
nand U5248 (N_5248,N_2753,N_3021);
nor U5249 (N_5249,N_2139,N_3825);
or U5250 (N_5250,N_3269,N_3072);
or U5251 (N_5251,N_2586,N_2776);
nand U5252 (N_5252,N_2672,N_2010);
nor U5253 (N_5253,N_2473,N_3407);
nor U5254 (N_5254,N_2084,N_2288);
and U5255 (N_5255,N_3640,N_2020);
or U5256 (N_5256,N_2959,N_2157);
nand U5257 (N_5257,N_2701,N_3790);
and U5258 (N_5258,N_2188,N_3635);
nand U5259 (N_5259,N_3097,N_3086);
nor U5260 (N_5260,N_3052,N_2933);
nand U5261 (N_5261,N_3592,N_2100);
nor U5262 (N_5262,N_3516,N_3333);
or U5263 (N_5263,N_2389,N_2266);
nand U5264 (N_5264,N_3151,N_3066);
or U5265 (N_5265,N_3868,N_3051);
nand U5266 (N_5266,N_2128,N_3799);
and U5267 (N_5267,N_2788,N_3211);
or U5268 (N_5268,N_2269,N_2769);
or U5269 (N_5269,N_3149,N_3190);
nand U5270 (N_5270,N_2110,N_2052);
nand U5271 (N_5271,N_3079,N_3672);
or U5272 (N_5272,N_2891,N_2710);
or U5273 (N_5273,N_3629,N_2920);
and U5274 (N_5274,N_2560,N_3914);
nor U5275 (N_5275,N_3547,N_3470);
or U5276 (N_5276,N_2748,N_3926);
or U5277 (N_5277,N_3890,N_3430);
nor U5278 (N_5278,N_2843,N_3350);
or U5279 (N_5279,N_3128,N_3794);
nand U5280 (N_5280,N_2734,N_2338);
and U5281 (N_5281,N_2505,N_2851);
or U5282 (N_5282,N_3946,N_2541);
and U5283 (N_5283,N_2675,N_3128);
nor U5284 (N_5284,N_2430,N_2493);
and U5285 (N_5285,N_3340,N_2354);
and U5286 (N_5286,N_3317,N_2650);
or U5287 (N_5287,N_3125,N_2444);
nor U5288 (N_5288,N_2576,N_2867);
and U5289 (N_5289,N_2636,N_3254);
nor U5290 (N_5290,N_3098,N_2024);
and U5291 (N_5291,N_3042,N_3242);
nand U5292 (N_5292,N_2130,N_2748);
and U5293 (N_5293,N_3637,N_3360);
and U5294 (N_5294,N_3088,N_3119);
and U5295 (N_5295,N_2291,N_2027);
nor U5296 (N_5296,N_2098,N_3196);
nor U5297 (N_5297,N_2216,N_2285);
nor U5298 (N_5298,N_3343,N_3549);
or U5299 (N_5299,N_3271,N_3682);
or U5300 (N_5300,N_2460,N_3895);
nand U5301 (N_5301,N_2292,N_3035);
or U5302 (N_5302,N_3080,N_2260);
or U5303 (N_5303,N_2522,N_3982);
or U5304 (N_5304,N_2849,N_2561);
or U5305 (N_5305,N_3888,N_3875);
or U5306 (N_5306,N_3998,N_3232);
nor U5307 (N_5307,N_3495,N_3250);
or U5308 (N_5308,N_2165,N_3765);
or U5309 (N_5309,N_2827,N_2451);
nand U5310 (N_5310,N_2204,N_2977);
and U5311 (N_5311,N_3140,N_2890);
and U5312 (N_5312,N_3877,N_3375);
nor U5313 (N_5313,N_2149,N_3630);
nor U5314 (N_5314,N_2106,N_2606);
nand U5315 (N_5315,N_3318,N_2965);
and U5316 (N_5316,N_2401,N_3311);
or U5317 (N_5317,N_3477,N_2968);
and U5318 (N_5318,N_2705,N_3721);
nand U5319 (N_5319,N_2068,N_2810);
nor U5320 (N_5320,N_2947,N_3432);
and U5321 (N_5321,N_3643,N_2017);
nor U5322 (N_5322,N_2507,N_2307);
and U5323 (N_5323,N_3833,N_3739);
or U5324 (N_5324,N_2994,N_3270);
nor U5325 (N_5325,N_3935,N_2796);
nor U5326 (N_5326,N_3593,N_3423);
nand U5327 (N_5327,N_3563,N_3173);
and U5328 (N_5328,N_3977,N_2093);
nor U5329 (N_5329,N_2297,N_3113);
and U5330 (N_5330,N_2261,N_3842);
nor U5331 (N_5331,N_3162,N_2698);
nand U5332 (N_5332,N_3341,N_3726);
and U5333 (N_5333,N_3384,N_3487);
nand U5334 (N_5334,N_2337,N_2738);
or U5335 (N_5335,N_3803,N_3866);
or U5336 (N_5336,N_2814,N_2863);
or U5337 (N_5337,N_3527,N_2024);
nor U5338 (N_5338,N_2232,N_2217);
and U5339 (N_5339,N_2823,N_3098);
or U5340 (N_5340,N_3972,N_2712);
nor U5341 (N_5341,N_3024,N_2602);
xor U5342 (N_5342,N_2850,N_3756);
and U5343 (N_5343,N_3747,N_3227);
and U5344 (N_5344,N_2849,N_2329);
xnor U5345 (N_5345,N_2424,N_2738);
and U5346 (N_5346,N_2023,N_2825);
nor U5347 (N_5347,N_3884,N_2284);
or U5348 (N_5348,N_2152,N_3473);
and U5349 (N_5349,N_2195,N_3940);
or U5350 (N_5350,N_2112,N_2481);
nor U5351 (N_5351,N_3261,N_2361);
and U5352 (N_5352,N_2146,N_3461);
nand U5353 (N_5353,N_2271,N_3822);
nand U5354 (N_5354,N_2589,N_3359);
or U5355 (N_5355,N_2738,N_2383);
nor U5356 (N_5356,N_3851,N_3731);
nor U5357 (N_5357,N_2521,N_2803);
nor U5358 (N_5358,N_3476,N_2708);
and U5359 (N_5359,N_2466,N_2321);
or U5360 (N_5360,N_3965,N_2437);
or U5361 (N_5361,N_2748,N_2035);
nand U5362 (N_5362,N_3017,N_3589);
or U5363 (N_5363,N_3695,N_2209);
nor U5364 (N_5364,N_3968,N_3254);
nand U5365 (N_5365,N_3869,N_2600);
nor U5366 (N_5366,N_2708,N_2814);
and U5367 (N_5367,N_2012,N_3872);
nand U5368 (N_5368,N_3554,N_3492);
nand U5369 (N_5369,N_2169,N_2477);
and U5370 (N_5370,N_3032,N_3949);
nand U5371 (N_5371,N_3839,N_2301);
nand U5372 (N_5372,N_3947,N_2275);
and U5373 (N_5373,N_3770,N_3708);
nand U5374 (N_5374,N_3870,N_2151);
or U5375 (N_5375,N_3687,N_2064);
or U5376 (N_5376,N_3663,N_3630);
xor U5377 (N_5377,N_2746,N_2832);
or U5378 (N_5378,N_2522,N_3756);
nand U5379 (N_5379,N_2763,N_2707);
and U5380 (N_5380,N_2171,N_2330);
nand U5381 (N_5381,N_2909,N_3440);
nand U5382 (N_5382,N_2580,N_2249);
nand U5383 (N_5383,N_2305,N_2869);
and U5384 (N_5384,N_3256,N_3623);
and U5385 (N_5385,N_2098,N_3538);
nor U5386 (N_5386,N_2815,N_3930);
and U5387 (N_5387,N_3230,N_2779);
or U5388 (N_5388,N_3194,N_3405);
nand U5389 (N_5389,N_2060,N_2858);
nor U5390 (N_5390,N_3134,N_2621);
nor U5391 (N_5391,N_2102,N_2679);
nor U5392 (N_5392,N_2025,N_2614);
and U5393 (N_5393,N_2695,N_2165);
and U5394 (N_5394,N_3570,N_2013);
and U5395 (N_5395,N_3892,N_2928);
nor U5396 (N_5396,N_2578,N_2045);
nand U5397 (N_5397,N_3173,N_2530);
and U5398 (N_5398,N_3423,N_2268);
nor U5399 (N_5399,N_3657,N_3766);
nand U5400 (N_5400,N_3022,N_3907);
nor U5401 (N_5401,N_2059,N_2982);
nand U5402 (N_5402,N_3230,N_3267);
or U5403 (N_5403,N_3616,N_3990);
and U5404 (N_5404,N_3607,N_2318);
and U5405 (N_5405,N_2565,N_2920);
or U5406 (N_5406,N_2140,N_2312);
nor U5407 (N_5407,N_2620,N_2478);
or U5408 (N_5408,N_2335,N_2171);
nor U5409 (N_5409,N_3130,N_2067);
or U5410 (N_5410,N_2735,N_2937);
or U5411 (N_5411,N_2524,N_2642);
or U5412 (N_5412,N_2475,N_2592);
and U5413 (N_5413,N_2622,N_2483);
nand U5414 (N_5414,N_2277,N_2390);
nor U5415 (N_5415,N_3923,N_3916);
nand U5416 (N_5416,N_3718,N_3448);
or U5417 (N_5417,N_2496,N_3897);
or U5418 (N_5418,N_2581,N_2449);
or U5419 (N_5419,N_3784,N_3368);
nand U5420 (N_5420,N_3082,N_2208);
and U5421 (N_5421,N_3957,N_3020);
and U5422 (N_5422,N_2092,N_3176);
nor U5423 (N_5423,N_2827,N_2187);
nand U5424 (N_5424,N_2922,N_2565);
xor U5425 (N_5425,N_3785,N_3818);
and U5426 (N_5426,N_3792,N_2946);
nor U5427 (N_5427,N_3712,N_3743);
nor U5428 (N_5428,N_3393,N_3870);
nor U5429 (N_5429,N_2083,N_2500);
nand U5430 (N_5430,N_2232,N_3849);
or U5431 (N_5431,N_3250,N_3084);
and U5432 (N_5432,N_2999,N_2932);
and U5433 (N_5433,N_3367,N_3421);
nand U5434 (N_5434,N_2298,N_3909);
nand U5435 (N_5435,N_3975,N_2659);
and U5436 (N_5436,N_2079,N_2326);
nand U5437 (N_5437,N_2642,N_3007);
and U5438 (N_5438,N_3215,N_2394);
or U5439 (N_5439,N_3664,N_3750);
nand U5440 (N_5440,N_2274,N_3002);
or U5441 (N_5441,N_2075,N_3139);
or U5442 (N_5442,N_3478,N_3741);
nand U5443 (N_5443,N_2858,N_3615);
or U5444 (N_5444,N_2531,N_3433);
nand U5445 (N_5445,N_3977,N_3292);
or U5446 (N_5446,N_3721,N_2971);
and U5447 (N_5447,N_2122,N_2890);
nor U5448 (N_5448,N_2138,N_3081);
nand U5449 (N_5449,N_2113,N_2758);
nor U5450 (N_5450,N_3522,N_2687);
and U5451 (N_5451,N_3694,N_2960);
or U5452 (N_5452,N_2263,N_3036);
nor U5453 (N_5453,N_2205,N_2170);
and U5454 (N_5454,N_2766,N_3343);
and U5455 (N_5455,N_2154,N_2785);
or U5456 (N_5456,N_3714,N_2994);
nor U5457 (N_5457,N_2100,N_3741);
and U5458 (N_5458,N_3340,N_3402);
nand U5459 (N_5459,N_2412,N_2388);
or U5460 (N_5460,N_3490,N_2168);
nand U5461 (N_5461,N_3152,N_2034);
nor U5462 (N_5462,N_3796,N_3907);
nand U5463 (N_5463,N_3931,N_3779);
and U5464 (N_5464,N_2717,N_2451);
or U5465 (N_5465,N_2333,N_2347);
and U5466 (N_5466,N_2421,N_3376);
or U5467 (N_5467,N_3390,N_2839);
nor U5468 (N_5468,N_2357,N_2170);
and U5469 (N_5469,N_3200,N_3828);
and U5470 (N_5470,N_2782,N_3252);
nand U5471 (N_5471,N_2579,N_2696);
nand U5472 (N_5472,N_3503,N_2643);
nand U5473 (N_5473,N_2179,N_2173);
or U5474 (N_5474,N_3565,N_3965);
and U5475 (N_5475,N_2081,N_3221);
or U5476 (N_5476,N_2437,N_2364);
or U5477 (N_5477,N_2695,N_2823);
nor U5478 (N_5478,N_3673,N_3740);
nor U5479 (N_5479,N_2584,N_3107);
or U5480 (N_5480,N_3023,N_3100);
and U5481 (N_5481,N_3727,N_2851);
nand U5482 (N_5482,N_2156,N_3791);
nor U5483 (N_5483,N_2784,N_2377);
nor U5484 (N_5484,N_3923,N_2185);
nand U5485 (N_5485,N_3771,N_2711);
nor U5486 (N_5486,N_3256,N_3411);
and U5487 (N_5487,N_2805,N_2621);
nor U5488 (N_5488,N_3745,N_2014);
nand U5489 (N_5489,N_2534,N_3983);
nor U5490 (N_5490,N_3533,N_2850);
nand U5491 (N_5491,N_2210,N_2973);
nor U5492 (N_5492,N_3326,N_2884);
or U5493 (N_5493,N_3161,N_3072);
or U5494 (N_5494,N_2755,N_3763);
nor U5495 (N_5495,N_2856,N_2168);
nand U5496 (N_5496,N_3991,N_2500);
and U5497 (N_5497,N_2663,N_3121);
nor U5498 (N_5498,N_2920,N_2752);
and U5499 (N_5499,N_3493,N_3109);
and U5500 (N_5500,N_3352,N_2248);
nand U5501 (N_5501,N_3878,N_3992);
nand U5502 (N_5502,N_3783,N_3119);
or U5503 (N_5503,N_2251,N_3392);
and U5504 (N_5504,N_2551,N_2464);
nand U5505 (N_5505,N_2582,N_2375);
nor U5506 (N_5506,N_2712,N_2828);
nor U5507 (N_5507,N_3869,N_3461);
or U5508 (N_5508,N_3148,N_2222);
and U5509 (N_5509,N_3520,N_2586);
nor U5510 (N_5510,N_2443,N_3464);
or U5511 (N_5511,N_3931,N_2233);
nand U5512 (N_5512,N_3304,N_2894);
and U5513 (N_5513,N_3523,N_2658);
and U5514 (N_5514,N_2815,N_2289);
or U5515 (N_5515,N_2289,N_2198);
or U5516 (N_5516,N_3713,N_2759);
or U5517 (N_5517,N_2310,N_3396);
or U5518 (N_5518,N_3831,N_3976);
nor U5519 (N_5519,N_3793,N_2663);
nor U5520 (N_5520,N_3805,N_2068);
or U5521 (N_5521,N_3168,N_3219);
and U5522 (N_5522,N_2342,N_3976);
and U5523 (N_5523,N_3324,N_2647);
or U5524 (N_5524,N_3713,N_3496);
nor U5525 (N_5525,N_2232,N_2005);
nor U5526 (N_5526,N_3187,N_3653);
nand U5527 (N_5527,N_3353,N_3799);
or U5528 (N_5528,N_2462,N_2874);
nor U5529 (N_5529,N_3945,N_2817);
nand U5530 (N_5530,N_2738,N_2293);
and U5531 (N_5531,N_2825,N_2222);
and U5532 (N_5532,N_2750,N_2881);
nor U5533 (N_5533,N_2449,N_2438);
nor U5534 (N_5534,N_3005,N_2211);
nor U5535 (N_5535,N_3148,N_3815);
xnor U5536 (N_5536,N_3022,N_3559);
or U5537 (N_5537,N_2712,N_3370);
and U5538 (N_5538,N_2707,N_2512);
nand U5539 (N_5539,N_2725,N_3298);
nand U5540 (N_5540,N_2440,N_2612);
nor U5541 (N_5541,N_3283,N_2383);
or U5542 (N_5542,N_2395,N_2840);
nor U5543 (N_5543,N_3828,N_2482);
and U5544 (N_5544,N_2627,N_2044);
or U5545 (N_5545,N_2656,N_2696);
or U5546 (N_5546,N_3382,N_2792);
nor U5547 (N_5547,N_3546,N_3062);
nand U5548 (N_5548,N_3866,N_2967);
nor U5549 (N_5549,N_3864,N_2135);
and U5550 (N_5550,N_2600,N_2044);
and U5551 (N_5551,N_3173,N_3256);
nand U5552 (N_5552,N_3033,N_3547);
nor U5553 (N_5553,N_2059,N_2779);
nor U5554 (N_5554,N_3479,N_3368);
nor U5555 (N_5555,N_3704,N_3597);
or U5556 (N_5556,N_3621,N_3489);
nand U5557 (N_5557,N_2185,N_2126);
or U5558 (N_5558,N_3112,N_2562);
and U5559 (N_5559,N_3209,N_2497);
nor U5560 (N_5560,N_2737,N_2464);
or U5561 (N_5561,N_3801,N_3532);
nor U5562 (N_5562,N_3300,N_2897);
and U5563 (N_5563,N_2200,N_3422);
and U5564 (N_5564,N_3588,N_3657);
nand U5565 (N_5565,N_2303,N_3645);
or U5566 (N_5566,N_2091,N_2888);
nor U5567 (N_5567,N_2395,N_2217);
and U5568 (N_5568,N_2928,N_3679);
and U5569 (N_5569,N_3867,N_3869);
and U5570 (N_5570,N_2351,N_2276);
nand U5571 (N_5571,N_2531,N_2798);
or U5572 (N_5572,N_3102,N_2421);
xnor U5573 (N_5573,N_2963,N_2040);
nor U5574 (N_5574,N_2604,N_2322);
or U5575 (N_5575,N_2512,N_3886);
or U5576 (N_5576,N_3168,N_3845);
and U5577 (N_5577,N_2606,N_3436);
or U5578 (N_5578,N_3510,N_2976);
nand U5579 (N_5579,N_3873,N_2308);
nand U5580 (N_5580,N_2822,N_3425);
or U5581 (N_5581,N_3061,N_2298);
or U5582 (N_5582,N_2073,N_3238);
or U5583 (N_5583,N_3011,N_2499);
or U5584 (N_5584,N_2548,N_3141);
or U5585 (N_5585,N_2082,N_3519);
and U5586 (N_5586,N_2441,N_3091);
nand U5587 (N_5587,N_2824,N_3569);
nor U5588 (N_5588,N_3591,N_2847);
or U5589 (N_5589,N_2024,N_3729);
nor U5590 (N_5590,N_2273,N_2740);
or U5591 (N_5591,N_3601,N_2437);
nand U5592 (N_5592,N_2638,N_2477);
and U5593 (N_5593,N_2539,N_3763);
or U5594 (N_5594,N_3143,N_3688);
and U5595 (N_5595,N_3503,N_2563);
xor U5596 (N_5596,N_3699,N_2703);
nand U5597 (N_5597,N_3556,N_3587);
nand U5598 (N_5598,N_2607,N_3429);
and U5599 (N_5599,N_3525,N_2068);
nand U5600 (N_5600,N_2203,N_2417);
and U5601 (N_5601,N_3045,N_2400);
or U5602 (N_5602,N_3470,N_2313);
or U5603 (N_5603,N_2178,N_2983);
nand U5604 (N_5604,N_2210,N_3726);
nor U5605 (N_5605,N_3946,N_2874);
nor U5606 (N_5606,N_2733,N_3043);
or U5607 (N_5607,N_3016,N_2639);
nor U5608 (N_5608,N_3553,N_2056);
and U5609 (N_5609,N_3713,N_2642);
and U5610 (N_5610,N_3696,N_3196);
nor U5611 (N_5611,N_3770,N_2852);
nand U5612 (N_5612,N_3282,N_3529);
nor U5613 (N_5613,N_3473,N_2130);
and U5614 (N_5614,N_2430,N_3995);
or U5615 (N_5615,N_3399,N_2749);
and U5616 (N_5616,N_3698,N_3688);
and U5617 (N_5617,N_3067,N_3349);
nor U5618 (N_5618,N_2350,N_3357);
and U5619 (N_5619,N_3512,N_3333);
and U5620 (N_5620,N_2288,N_3539);
nor U5621 (N_5621,N_2969,N_3721);
or U5622 (N_5622,N_2140,N_3409);
nand U5623 (N_5623,N_2506,N_2706);
nor U5624 (N_5624,N_2948,N_2691);
and U5625 (N_5625,N_3574,N_3854);
or U5626 (N_5626,N_3770,N_3791);
and U5627 (N_5627,N_2348,N_3819);
and U5628 (N_5628,N_2639,N_3998);
nand U5629 (N_5629,N_3565,N_3393);
nor U5630 (N_5630,N_3616,N_2529);
nand U5631 (N_5631,N_3820,N_3558);
nor U5632 (N_5632,N_2838,N_3346);
or U5633 (N_5633,N_3041,N_3220);
or U5634 (N_5634,N_2777,N_3605);
nor U5635 (N_5635,N_2221,N_3219);
and U5636 (N_5636,N_2976,N_2087);
or U5637 (N_5637,N_3279,N_2074);
nand U5638 (N_5638,N_2574,N_3779);
nor U5639 (N_5639,N_2038,N_3601);
or U5640 (N_5640,N_3510,N_2666);
nor U5641 (N_5641,N_3227,N_2296);
and U5642 (N_5642,N_3135,N_2287);
and U5643 (N_5643,N_2008,N_2771);
nor U5644 (N_5644,N_2322,N_2176);
and U5645 (N_5645,N_3483,N_3057);
and U5646 (N_5646,N_3854,N_3893);
nor U5647 (N_5647,N_2976,N_3602);
nand U5648 (N_5648,N_2005,N_3911);
xor U5649 (N_5649,N_2222,N_3020);
or U5650 (N_5650,N_2109,N_2633);
and U5651 (N_5651,N_3931,N_3580);
or U5652 (N_5652,N_2978,N_2905);
and U5653 (N_5653,N_3044,N_2555);
and U5654 (N_5654,N_2515,N_2666);
nor U5655 (N_5655,N_2665,N_3450);
and U5656 (N_5656,N_2091,N_3339);
nand U5657 (N_5657,N_3330,N_3021);
nor U5658 (N_5658,N_2781,N_2574);
and U5659 (N_5659,N_2891,N_2905);
nand U5660 (N_5660,N_2440,N_2119);
nand U5661 (N_5661,N_2993,N_3234);
nand U5662 (N_5662,N_2409,N_2075);
and U5663 (N_5663,N_2520,N_2446);
nand U5664 (N_5664,N_2811,N_2353);
and U5665 (N_5665,N_2657,N_2771);
and U5666 (N_5666,N_2300,N_2550);
nand U5667 (N_5667,N_2597,N_3704);
nand U5668 (N_5668,N_3733,N_3101);
nor U5669 (N_5669,N_2886,N_3183);
and U5670 (N_5670,N_3417,N_2350);
or U5671 (N_5671,N_3638,N_2687);
nor U5672 (N_5672,N_2242,N_3046);
nor U5673 (N_5673,N_3989,N_3567);
nand U5674 (N_5674,N_2893,N_2735);
and U5675 (N_5675,N_3731,N_3452);
nor U5676 (N_5676,N_3779,N_2728);
or U5677 (N_5677,N_2536,N_3166);
or U5678 (N_5678,N_2163,N_3325);
and U5679 (N_5679,N_3911,N_2905);
and U5680 (N_5680,N_2227,N_2182);
or U5681 (N_5681,N_2333,N_3222);
nand U5682 (N_5682,N_2677,N_3301);
or U5683 (N_5683,N_3765,N_2341);
or U5684 (N_5684,N_2155,N_3198);
and U5685 (N_5685,N_3731,N_3422);
nor U5686 (N_5686,N_3296,N_3898);
xor U5687 (N_5687,N_3882,N_3272);
or U5688 (N_5688,N_3257,N_3992);
nor U5689 (N_5689,N_3321,N_3503);
nand U5690 (N_5690,N_3210,N_2895);
and U5691 (N_5691,N_3228,N_2343);
and U5692 (N_5692,N_2313,N_3286);
nand U5693 (N_5693,N_2510,N_3444);
nand U5694 (N_5694,N_3159,N_3211);
or U5695 (N_5695,N_2787,N_3946);
nand U5696 (N_5696,N_2669,N_3216);
nand U5697 (N_5697,N_3559,N_2882);
and U5698 (N_5698,N_2163,N_2820);
or U5699 (N_5699,N_2656,N_2693);
nor U5700 (N_5700,N_3527,N_3645);
nor U5701 (N_5701,N_2144,N_2348);
nand U5702 (N_5702,N_3996,N_3041);
nor U5703 (N_5703,N_2842,N_2835);
and U5704 (N_5704,N_3303,N_2657);
nand U5705 (N_5705,N_2155,N_2640);
or U5706 (N_5706,N_2853,N_3151);
nand U5707 (N_5707,N_3028,N_3126);
and U5708 (N_5708,N_2448,N_3807);
and U5709 (N_5709,N_3281,N_2083);
nor U5710 (N_5710,N_3846,N_3267);
or U5711 (N_5711,N_2055,N_2642);
nand U5712 (N_5712,N_2857,N_3369);
nand U5713 (N_5713,N_3760,N_2782);
nor U5714 (N_5714,N_3774,N_3442);
or U5715 (N_5715,N_3458,N_3770);
and U5716 (N_5716,N_3851,N_2877);
and U5717 (N_5717,N_3448,N_2715);
or U5718 (N_5718,N_3032,N_3827);
nand U5719 (N_5719,N_3593,N_3922);
nand U5720 (N_5720,N_3195,N_2767);
and U5721 (N_5721,N_2518,N_2754);
or U5722 (N_5722,N_2347,N_3550);
or U5723 (N_5723,N_2737,N_2666);
and U5724 (N_5724,N_3849,N_3050);
nand U5725 (N_5725,N_3865,N_3112);
nand U5726 (N_5726,N_2813,N_3283);
nand U5727 (N_5727,N_2657,N_3588);
nand U5728 (N_5728,N_2969,N_2596);
and U5729 (N_5729,N_3771,N_3892);
nor U5730 (N_5730,N_3457,N_2169);
or U5731 (N_5731,N_3552,N_2234);
or U5732 (N_5732,N_2512,N_2237);
and U5733 (N_5733,N_3928,N_3165);
nor U5734 (N_5734,N_3725,N_2601);
or U5735 (N_5735,N_3823,N_3124);
or U5736 (N_5736,N_2635,N_3532);
nor U5737 (N_5737,N_2580,N_2914);
and U5738 (N_5738,N_2587,N_3186);
nor U5739 (N_5739,N_3959,N_3103);
nand U5740 (N_5740,N_3342,N_2180);
and U5741 (N_5741,N_3436,N_2401);
and U5742 (N_5742,N_2157,N_3894);
and U5743 (N_5743,N_2572,N_3981);
nand U5744 (N_5744,N_3205,N_3872);
and U5745 (N_5745,N_2070,N_3460);
nor U5746 (N_5746,N_2863,N_2443);
nor U5747 (N_5747,N_2931,N_2269);
or U5748 (N_5748,N_2876,N_2551);
nand U5749 (N_5749,N_2763,N_3259);
or U5750 (N_5750,N_3462,N_3763);
or U5751 (N_5751,N_3593,N_2206);
nor U5752 (N_5752,N_3291,N_3048);
and U5753 (N_5753,N_3919,N_3782);
or U5754 (N_5754,N_2811,N_2699);
or U5755 (N_5755,N_3495,N_3558);
or U5756 (N_5756,N_3797,N_2822);
or U5757 (N_5757,N_3129,N_3341);
nor U5758 (N_5758,N_2399,N_2861);
nor U5759 (N_5759,N_3788,N_2212);
nand U5760 (N_5760,N_2850,N_2766);
nand U5761 (N_5761,N_3071,N_3050);
nand U5762 (N_5762,N_2319,N_2672);
or U5763 (N_5763,N_3676,N_3377);
and U5764 (N_5764,N_2021,N_3166);
nor U5765 (N_5765,N_3286,N_3458);
or U5766 (N_5766,N_2232,N_3252);
and U5767 (N_5767,N_3144,N_2286);
or U5768 (N_5768,N_2668,N_2652);
and U5769 (N_5769,N_2185,N_2777);
and U5770 (N_5770,N_2270,N_2365);
or U5771 (N_5771,N_2670,N_3160);
nor U5772 (N_5772,N_3565,N_3621);
nor U5773 (N_5773,N_3399,N_3124);
or U5774 (N_5774,N_2176,N_3494);
or U5775 (N_5775,N_3537,N_3247);
nor U5776 (N_5776,N_2779,N_3231);
or U5777 (N_5777,N_3592,N_2909);
nor U5778 (N_5778,N_3431,N_2502);
or U5779 (N_5779,N_3282,N_2306);
and U5780 (N_5780,N_2820,N_2234);
or U5781 (N_5781,N_3274,N_3623);
nor U5782 (N_5782,N_2272,N_3142);
or U5783 (N_5783,N_2915,N_2998);
nor U5784 (N_5784,N_3002,N_2484);
nor U5785 (N_5785,N_3172,N_2985);
nor U5786 (N_5786,N_2333,N_3628);
nand U5787 (N_5787,N_2005,N_2711);
nand U5788 (N_5788,N_2299,N_2513);
or U5789 (N_5789,N_2720,N_3118);
nand U5790 (N_5790,N_2290,N_3692);
nand U5791 (N_5791,N_3438,N_3375);
or U5792 (N_5792,N_2186,N_2314);
nand U5793 (N_5793,N_2744,N_2462);
or U5794 (N_5794,N_2290,N_3152);
or U5795 (N_5795,N_3780,N_2818);
nand U5796 (N_5796,N_2455,N_2054);
nor U5797 (N_5797,N_3423,N_2409);
or U5798 (N_5798,N_2314,N_3020);
and U5799 (N_5799,N_3100,N_2017);
and U5800 (N_5800,N_2458,N_3502);
nand U5801 (N_5801,N_3615,N_2031);
nor U5802 (N_5802,N_2104,N_2156);
and U5803 (N_5803,N_3800,N_3106);
nor U5804 (N_5804,N_3717,N_3721);
and U5805 (N_5805,N_3702,N_3509);
nand U5806 (N_5806,N_3018,N_2718);
nand U5807 (N_5807,N_3548,N_3336);
or U5808 (N_5808,N_3958,N_2139);
or U5809 (N_5809,N_3294,N_2162);
and U5810 (N_5810,N_2452,N_2564);
nor U5811 (N_5811,N_2221,N_2642);
and U5812 (N_5812,N_2892,N_3047);
nor U5813 (N_5813,N_3819,N_2005);
nor U5814 (N_5814,N_2890,N_3225);
and U5815 (N_5815,N_3913,N_3510);
nor U5816 (N_5816,N_2004,N_3419);
and U5817 (N_5817,N_2528,N_2791);
nand U5818 (N_5818,N_3509,N_3577);
or U5819 (N_5819,N_2332,N_3336);
nor U5820 (N_5820,N_2569,N_2044);
nand U5821 (N_5821,N_3733,N_3657);
nand U5822 (N_5822,N_2307,N_2885);
and U5823 (N_5823,N_2688,N_2893);
nor U5824 (N_5824,N_3665,N_3143);
nor U5825 (N_5825,N_2656,N_2596);
and U5826 (N_5826,N_3198,N_3938);
nand U5827 (N_5827,N_3971,N_2451);
nand U5828 (N_5828,N_3887,N_3823);
or U5829 (N_5829,N_2832,N_2531);
nand U5830 (N_5830,N_2064,N_3551);
and U5831 (N_5831,N_2877,N_3784);
nor U5832 (N_5832,N_2246,N_3334);
or U5833 (N_5833,N_2098,N_3774);
nand U5834 (N_5834,N_3241,N_2056);
and U5835 (N_5835,N_2533,N_3612);
or U5836 (N_5836,N_3382,N_3351);
and U5837 (N_5837,N_3833,N_2432);
and U5838 (N_5838,N_3873,N_3160);
and U5839 (N_5839,N_2677,N_2012);
nand U5840 (N_5840,N_2639,N_2629);
nand U5841 (N_5841,N_2855,N_2367);
nand U5842 (N_5842,N_3530,N_3280);
or U5843 (N_5843,N_3264,N_3568);
nand U5844 (N_5844,N_2425,N_3091);
or U5845 (N_5845,N_3373,N_2035);
or U5846 (N_5846,N_3410,N_3901);
nor U5847 (N_5847,N_2031,N_2548);
or U5848 (N_5848,N_2262,N_3537);
nand U5849 (N_5849,N_2796,N_3492);
nor U5850 (N_5850,N_3397,N_2081);
nand U5851 (N_5851,N_2136,N_2452);
nor U5852 (N_5852,N_3652,N_3177);
nor U5853 (N_5853,N_3581,N_2571);
nand U5854 (N_5854,N_3150,N_2321);
and U5855 (N_5855,N_3302,N_3561);
nand U5856 (N_5856,N_2148,N_3433);
and U5857 (N_5857,N_3614,N_2829);
and U5858 (N_5858,N_3757,N_3736);
nand U5859 (N_5859,N_3194,N_3399);
and U5860 (N_5860,N_2926,N_3869);
and U5861 (N_5861,N_3678,N_2555);
or U5862 (N_5862,N_2684,N_3891);
or U5863 (N_5863,N_2586,N_3977);
or U5864 (N_5864,N_3187,N_2326);
and U5865 (N_5865,N_3650,N_3057);
and U5866 (N_5866,N_3250,N_3810);
or U5867 (N_5867,N_2171,N_2526);
nand U5868 (N_5868,N_3207,N_3457);
nand U5869 (N_5869,N_3496,N_2231);
nor U5870 (N_5870,N_3961,N_2356);
and U5871 (N_5871,N_3486,N_2914);
and U5872 (N_5872,N_3141,N_2277);
nand U5873 (N_5873,N_2562,N_3288);
or U5874 (N_5874,N_3418,N_3203);
and U5875 (N_5875,N_2997,N_3455);
or U5876 (N_5876,N_2392,N_2984);
and U5877 (N_5877,N_2403,N_2021);
and U5878 (N_5878,N_2190,N_2599);
or U5879 (N_5879,N_3657,N_3412);
nor U5880 (N_5880,N_2564,N_2336);
or U5881 (N_5881,N_2709,N_3680);
or U5882 (N_5882,N_2082,N_2955);
and U5883 (N_5883,N_3396,N_3252);
nor U5884 (N_5884,N_2335,N_3472);
and U5885 (N_5885,N_2125,N_2657);
and U5886 (N_5886,N_2796,N_2893);
nand U5887 (N_5887,N_2865,N_2997);
or U5888 (N_5888,N_2439,N_3510);
nand U5889 (N_5889,N_2698,N_3179);
or U5890 (N_5890,N_2866,N_2702);
nor U5891 (N_5891,N_2952,N_2556);
or U5892 (N_5892,N_3026,N_2766);
nand U5893 (N_5893,N_3482,N_2696);
and U5894 (N_5894,N_3986,N_2053);
and U5895 (N_5895,N_2026,N_3013);
nand U5896 (N_5896,N_2011,N_2799);
nor U5897 (N_5897,N_2455,N_3000);
nor U5898 (N_5898,N_3548,N_3103);
nand U5899 (N_5899,N_2288,N_2113);
or U5900 (N_5900,N_3095,N_3763);
and U5901 (N_5901,N_3356,N_2196);
and U5902 (N_5902,N_3152,N_2382);
and U5903 (N_5903,N_2251,N_3585);
nor U5904 (N_5904,N_2027,N_3564);
or U5905 (N_5905,N_3665,N_3231);
nor U5906 (N_5906,N_2717,N_3716);
and U5907 (N_5907,N_3700,N_2550);
nand U5908 (N_5908,N_3385,N_3519);
or U5909 (N_5909,N_2157,N_2264);
or U5910 (N_5910,N_2695,N_2814);
nand U5911 (N_5911,N_2810,N_3110);
nand U5912 (N_5912,N_3611,N_3831);
nor U5913 (N_5913,N_3595,N_3023);
nor U5914 (N_5914,N_3859,N_2202);
nor U5915 (N_5915,N_2254,N_2052);
or U5916 (N_5916,N_2916,N_3185);
nor U5917 (N_5917,N_2466,N_3723);
and U5918 (N_5918,N_2646,N_3015);
nor U5919 (N_5919,N_2198,N_2692);
nor U5920 (N_5920,N_2271,N_2847);
and U5921 (N_5921,N_3145,N_3435);
nor U5922 (N_5922,N_3567,N_2827);
and U5923 (N_5923,N_2371,N_2453);
and U5924 (N_5924,N_3235,N_3231);
nand U5925 (N_5925,N_2328,N_2003);
nand U5926 (N_5926,N_3750,N_3518);
nor U5927 (N_5927,N_2927,N_3168);
nor U5928 (N_5928,N_2405,N_2065);
or U5929 (N_5929,N_3119,N_3036);
and U5930 (N_5930,N_3295,N_3761);
or U5931 (N_5931,N_3132,N_3992);
or U5932 (N_5932,N_3439,N_2622);
nand U5933 (N_5933,N_3051,N_3425);
and U5934 (N_5934,N_3624,N_2767);
and U5935 (N_5935,N_2985,N_3601);
and U5936 (N_5936,N_2289,N_3985);
and U5937 (N_5937,N_3765,N_2542);
and U5938 (N_5938,N_3012,N_3846);
and U5939 (N_5939,N_3514,N_2899);
and U5940 (N_5940,N_3379,N_3396);
nor U5941 (N_5941,N_2537,N_2525);
nand U5942 (N_5942,N_2253,N_2965);
nor U5943 (N_5943,N_2092,N_2320);
nand U5944 (N_5944,N_3167,N_3560);
and U5945 (N_5945,N_3792,N_3652);
and U5946 (N_5946,N_3072,N_3554);
nor U5947 (N_5947,N_2938,N_2231);
nand U5948 (N_5948,N_3089,N_3914);
nor U5949 (N_5949,N_2781,N_2248);
or U5950 (N_5950,N_2581,N_3036);
nand U5951 (N_5951,N_3728,N_3527);
and U5952 (N_5952,N_2031,N_2686);
nand U5953 (N_5953,N_3880,N_2420);
or U5954 (N_5954,N_3007,N_3495);
or U5955 (N_5955,N_3418,N_3130);
nand U5956 (N_5956,N_3276,N_2163);
xnor U5957 (N_5957,N_2493,N_2513);
nor U5958 (N_5958,N_2845,N_2415);
or U5959 (N_5959,N_3103,N_3180);
or U5960 (N_5960,N_2434,N_2991);
nor U5961 (N_5961,N_3502,N_2965);
and U5962 (N_5962,N_3732,N_3039);
and U5963 (N_5963,N_2146,N_3025);
and U5964 (N_5964,N_3227,N_3019);
nand U5965 (N_5965,N_3968,N_3071);
nand U5966 (N_5966,N_2872,N_3432);
and U5967 (N_5967,N_3237,N_3010);
nand U5968 (N_5968,N_2792,N_2976);
or U5969 (N_5969,N_2327,N_2364);
and U5970 (N_5970,N_3437,N_3116);
nor U5971 (N_5971,N_2169,N_2643);
or U5972 (N_5972,N_3450,N_2870);
nand U5973 (N_5973,N_2151,N_3617);
or U5974 (N_5974,N_3180,N_3821);
or U5975 (N_5975,N_3227,N_3859);
and U5976 (N_5976,N_2190,N_2356);
nor U5977 (N_5977,N_3513,N_2251);
nand U5978 (N_5978,N_3435,N_2248);
nand U5979 (N_5979,N_3839,N_2229);
nor U5980 (N_5980,N_3884,N_3610);
and U5981 (N_5981,N_3276,N_3800);
nand U5982 (N_5982,N_3577,N_2392);
and U5983 (N_5983,N_2124,N_3631);
xnor U5984 (N_5984,N_2765,N_3276);
nor U5985 (N_5985,N_2425,N_3614);
and U5986 (N_5986,N_2447,N_3693);
nand U5987 (N_5987,N_3011,N_3567);
or U5988 (N_5988,N_3096,N_3577);
or U5989 (N_5989,N_3543,N_3309);
nor U5990 (N_5990,N_2235,N_2392);
nor U5991 (N_5991,N_2181,N_2325);
nand U5992 (N_5992,N_2043,N_3834);
nand U5993 (N_5993,N_3365,N_3185);
nor U5994 (N_5994,N_2246,N_2197);
or U5995 (N_5995,N_2906,N_3436);
and U5996 (N_5996,N_2263,N_2422);
and U5997 (N_5997,N_2296,N_3770);
nand U5998 (N_5998,N_2791,N_3286);
nor U5999 (N_5999,N_2051,N_3009);
or U6000 (N_6000,N_4608,N_5838);
and U6001 (N_6001,N_5726,N_5764);
nor U6002 (N_6002,N_4393,N_4708);
or U6003 (N_6003,N_5735,N_4843);
or U6004 (N_6004,N_5930,N_5433);
or U6005 (N_6005,N_5058,N_4826);
xor U6006 (N_6006,N_5569,N_5293);
or U6007 (N_6007,N_5772,N_5851);
nand U6008 (N_6008,N_5744,N_4698);
or U6009 (N_6009,N_4602,N_5828);
nand U6010 (N_6010,N_4982,N_5814);
nand U6011 (N_6011,N_4274,N_4965);
nand U6012 (N_6012,N_5103,N_4131);
or U6013 (N_6013,N_4800,N_5129);
nor U6014 (N_6014,N_5820,N_5128);
nand U6015 (N_6015,N_4941,N_5414);
and U6016 (N_6016,N_4389,N_5046);
nor U6017 (N_6017,N_4864,N_5862);
xnor U6018 (N_6018,N_4366,N_4355);
or U6019 (N_6019,N_5776,N_5198);
nand U6020 (N_6020,N_4308,N_4600);
nand U6021 (N_6021,N_5054,N_4183);
nor U6022 (N_6022,N_5297,N_5605);
nand U6023 (N_6023,N_5403,N_5892);
nor U6024 (N_6024,N_4759,N_5543);
or U6025 (N_6025,N_4337,N_4762);
nand U6026 (N_6026,N_5727,N_5965);
nor U6027 (N_6027,N_5210,N_4169);
and U6028 (N_6028,N_5702,N_4012);
nand U6029 (N_6029,N_5205,N_5720);
nand U6030 (N_6030,N_5673,N_5999);
or U6031 (N_6031,N_5519,N_4089);
or U6032 (N_6032,N_5871,N_4410);
nand U6033 (N_6033,N_4589,N_4388);
nor U6034 (N_6034,N_4527,N_5746);
and U6035 (N_6035,N_4260,N_5259);
nor U6036 (N_6036,N_5879,N_4263);
nand U6037 (N_6037,N_4060,N_5283);
nand U6038 (N_6038,N_5540,N_5021);
or U6039 (N_6039,N_5284,N_5905);
and U6040 (N_6040,N_5171,N_5212);
or U6041 (N_6041,N_5802,N_4426);
nor U6042 (N_6042,N_4435,N_4372);
nor U6043 (N_6043,N_5958,N_4382);
and U6044 (N_6044,N_4996,N_5455);
nor U6045 (N_6045,N_5904,N_5339);
nand U6046 (N_6046,N_4760,N_4703);
nor U6047 (N_6047,N_4110,N_4367);
or U6048 (N_6048,N_4855,N_5131);
and U6049 (N_6049,N_5832,N_4559);
nand U6050 (N_6050,N_4117,N_4536);
nand U6051 (N_6051,N_4444,N_4515);
xnor U6052 (N_6052,N_5918,N_4324);
nor U6053 (N_6053,N_5754,N_5057);
nor U6054 (N_6054,N_5932,N_4926);
or U6055 (N_6055,N_5014,N_5773);
nand U6056 (N_6056,N_4599,N_4116);
nor U6057 (N_6057,N_4567,N_4670);
or U6058 (N_6058,N_4788,N_4310);
nand U6059 (N_6059,N_4883,N_5392);
nand U6060 (N_6060,N_5367,N_4139);
nand U6061 (N_6061,N_5602,N_4652);
and U6062 (N_6062,N_4043,N_5873);
nand U6063 (N_6063,N_5740,N_4962);
nand U6064 (N_6064,N_4576,N_4174);
or U6065 (N_6065,N_5739,N_5092);
and U6066 (N_6066,N_4838,N_4816);
nand U6067 (N_6067,N_4806,N_4176);
and U6068 (N_6068,N_4445,N_4297);
or U6069 (N_6069,N_5579,N_5537);
nand U6070 (N_6070,N_5565,N_4557);
or U6071 (N_6071,N_5886,N_4172);
and U6072 (N_6072,N_5416,N_4398);
nor U6073 (N_6073,N_4230,N_5557);
xor U6074 (N_6074,N_5115,N_5067);
and U6075 (N_6075,N_4924,N_4810);
nand U6076 (N_6076,N_5943,N_4828);
nand U6077 (N_6077,N_5812,N_4699);
or U6078 (N_6078,N_5803,N_5914);
or U6079 (N_6079,N_5531,N_4912);
xnor U6080 (N_6080,N_4119,N_4916);
and U6081 (N_6081,N_5227,N_5423);
nor U6082 (N_6082,N_4240,N_4848);
nand U6083 (N_6083,N_4009,N_5217);
nor U6084 (N_6084,N_5321,N_5829);
nor U6085 (N_6085,N_5162,N_5927);
and U6086 (N_6086,N_5571,N_5420);
and U6087 (N_6087,N_4207,N_5595);
or U6088 (N_6088,N_4636,N_4349);
nor U6089 (N_6089,N_5593,N_4632);
nor U6090 (N_6090,N_5143,N_4970);
or U6091 (N_6091,N_5608,N_5601);
nor U6092 (N_6092,N_5796,N_5575);
nor U6093 (N_6093,N_4231,N_5368);
or U6094 (N_6094,N_5265,N_5559);
or U6095 (N_6095,N_4879,N_4891);
or U6096 (N_6096,N_4854,N_5833);
and U6097 (N_6097,N_4930,N_4796);
nor U6098 (N_6098,N_4386,N_4819);
nand U6099 (N_6099,N_5859,N_5946);
and U6100 (N_6100,N_4002,N_4453);
or U6101 (N_6101,N_4877,N_4323);
and U6102 (N_6102,N_5426,N_5081);
xnor U6103 (N_6103,N_4190,N_5093);
xnor U6104 (N_6104,N_4540,N_4232);
and U6105 (N_6105,N_5948,N_5402);
nand U6106 (N_6106,N_4114,N_4691);
nor U6107 (N_6107,N_4302,N_5254);
nor U6108 (N_6108,N_4124,N_4049);
nand U6109 (N_6109,N_4211,N_4734);
nor U6110 (N_6110,N_5195,N_4038);
nor U6111 (N_6111,N_4693,N_5994);
or U6112 (N_6112,N_5363,N_5141);
nand U6113 (N_6113,N_4619,N_4106);
xnor U6114 (N_6114,N_5737,N_4665);
nor U6115 (N_6115,N_4330,N_5938);
and U6116 (N_6116,N_4784,N_5808);
nor U6117 (N_6117,N_5449,N_4503);
or U6118 (N_6118,N_5419,N_5199);
or U6119 (N_6119,N_5184,N_4897);
nand U6120 (N_6120,N_4121,N_4173);
and U6121 (N_6121,N_5604,N_4611);
and U6122 (N_6122,N_4082,N_4751);
nand U6123 (N_6123,N_4678,N_5424);
nor U6124 (N_6124,N_4776,N_4320);
or U6125 (N_6125,N_5916,N_5634);
and U6126 (N_6126,N_4747,N_4161);
nor U6127 (N_6127,N_5568,N_5885);
nor U6128 (N_6128,N_5157,N_5477);
nand U6129 (N_6129,N_4204,N_4625);
or U6130 (N_6130,N_4917,N_4166);
nand U6131 (N_6131,N_4409,N_5815);
nand U6132 (N_6132,N_5296,N_4309);
and U6133 (N_6133,N_4830,N_5194);
nand U6134 (N_6134,N_5759,N_5507);
nand U6135 (N_6135,N_5900,N_5896);
nand U6136 (N_6136,N_5797,N_5336);
nor U6137 (N_6137,N_4241,N_5708);
nor U6138 (N_6138,N_4006,N_4514);
nor U6139 (N_6139,N_5767,N_4675);
nand U6140 (N_6140,N_5113,N_5854);
nor U6141 (N_6141,N_5972,N_5233);
or U6142 (N_6142,N_4091,N_5091);
or U6143 (N_6143,N_5556,N_5677);
or U6144 (N_6144,N_4298,N_5226);
nand U6145 (N_6145,N_5350,N_4971);
and U6146 (N_6146,N_4150,N_5834);
nand U6147 (N_6147,N_4282,N_4072);
or U6148 (N_6148,N_5524,N_5077);
and U6149 (N_6149,N_4672,N_4414);
xor U6150 (N_6150,N_5635,N_4640);
nor U6151 (N_6151,N_5984,N_4687);
nor U6152 (N_6152,N_5782,N_4543);
and U6153 (N_6153,N_5170,N_4122);
nor U6154 (N_6154,N_5530,N_5730);
nand U6155 (N_6155,N_5039,N_5514);
nand U6156 (N_6156,N_4154,N_4815);
and U6157 (N_6157,N_5451,N_5752);
or U6158 (N_6158,N_4876,N_4521);
or U6159 (N_6159,N_4225,N_4785);
or U6160 (N_6160,N_4215,N_4909);
nand U6161 (N_6161,N_4904,N_5272);
or U6162 (N_6162,N_5732,N_5788);
nand U6163 (N_6163,N_4622,N_5799);
and U6164 (N_6164,N_4051,N_4763);
or U6165 (N_6165,N_4949,N_5022);
and U6166 (N_6166,N_4416,N_5709);
nor U6167 (N_6167,N_5515,N_5246);
or U6168 (N_6168,N_5358,N_5095);
nor U6169 (N_6169,N_4832,N_4755);
nor U6170 (N_6170,N_4710,N_5674);
and U6171 (N_6171,N_5983,N_4448);
nor U6172 (N_6172,N_5945,N_5496);
nor U6173 (N_6173,N_5098,N_5355);
and U6174 (N_6174,N_5700,N_4835);
nand U6175 (N_6175,N_5750,N_4406);
nor U6176 (N_6176,N_4723,N_5600);
nand U6177 (N_6177,N_4922,N_4782);
and U6178 (N_6178,N_5209,N_4075);
nand U6179 (N_6179,N_4220,N_5742);
nor U6180 (N_6180,N_5071,N_5382);
nor U6181 (N_6181,N_5895,N_4743);
nand U6182 (N_6182,N_5408,N_4590);
nand U6183 (N_6183,N_4849,N_5391);
nand U6184 (N_6184,N_5539,N_5388);
nand U6185 (N_6185,N_5572,N_4004);
nor U6186 (N_6186,N_5036,N_5631);
or U6187 (N_6187,N_4682,N_5073);
and U6188 (N_6188,N_5340,N_4945);
nor U6189 (N_6189,N_5399,N_5192);
nor U6190 (N_6190,N_4030,N_4679);
nor U6191 (N_6191,N_4192,N_4994);
or U6192 (N_6192,N_4680,N_4504);
or U6193 (N_6193,N_5224,N_4168);
nor U6194 (N_6194,N_4911,N_5670);
nand U6195 (N_6195,N_5292,N_5682);
and U6196 (N_6196,N_4947,N_4251);
or U6197 (N_6197,N_5791,N_4422);
and U6198 (N_6198,N_5055,N_4653);
nor U6199 (N_6199,N_5040,N_5500);
nand U6200 (N_6200,N_4713,N_5486);
and U6201 (N_6201,N_5641,N_5061);
nor U6202 (N_6202,N_4821,N_4532);
nand U6203 (N_6203,N_4431,N_4813);
nand U6204 (N_6204,N_4351,N_4558);
nor U6205 (N_6205,N_4766,N_4487);
and U6206 (N_6206,N_5454,N_5704);
and U6207 (N_6207,N_5405,N_4510);
nor U6208 (N_6208,N_4081,N_5146);
or U6209 (N_6209,N_5675,N_4040);
or U6210 (N_6210,N_5643,N_5109);
and U6211 (N_6211,N_4279,N_4860);
nand U6212 (N_6212,N_4048,N_5963);
or U6213 (N_6213,N_5723,N_5560);
nor U6214 (N_6214,N_5252,N_4221);
or U6215 (N_6215,N_4107,N_5268);
nand U6216 (N_6216,N_5487,N_4010);
or U6217 (N_6217,N_5733,N_4206);
nor U6218 (N_6218,N_4481,N_5415);
and U6219 (N_6219,N_4547,N_5661);
nor U6220 (N_6220,N_5889,N_5458);
nor U6221 (N_6221,N_4633,N_5019);
nor U6222 (N_6222,N_4775,N_5084);
or U6223 (N_6223,N_4118,N_4151);
or U6224 (N_6224,N_4530,N_5894);
nand U6225 (N_6225,N_4967,N_5887);
nand U6226 (N_6226,N_5235,N_5488);
nor U6227 (N_6227,N_5609,N_4780);
nor U6228 (N_6228,N_5182,N_4071);
nor U6229 (N_6229,N_4553,N_5187);
and U6230 (N_6230,N_4613,N_4457);
and U6231 (N_6231,N_5615,N_4379);
and U6232 (N_6232,N_4674,N_4973);
and U6233 (N_6233,N_4787,N_4099);
and U6234 (N_6234,N_5503,N_5956);
nand U6235 (N_6235,N_5206,N_4271);
or U6236 (N_6236,N_5654,N_5592);
nand U6237 (N_6237,N_4560,N_4023);
nor U6238 (N_6238,N_5305,N_5033);
nand U6239 (N_6239,N_4132,N_4129);
and U6240 (N_6240,N_4976,N_5981);
nor U6241 (N_6241,N_4722,N_4671);
nor U6242 (N_6242,N_4020,N_4783);
nor U6243 (N_6243,N_5010,N_5625);
nor U6244 (N_6244,N_4272,N_5218);
and U6245 (N_6245,N_5165,N_5714);
nand U6246 (N_6246,N_5979,N_5111);
nor U6247 (N_6247,N_4906,N_5903);
xor U6248 (N_6248,N_5304,N_5590);
and U6249 (N_6249,N_4688,N_5678);
nand U6250 (N_6250,N_5207,N_5324);
and U6251 (N_6251,N_5468,N_4342);
nor U6252 (N_6252,N_4027,N_5756);
nor U6253 (N_6253,N_4455,N_5237);
nor U6254 (N_6254,N_4656,N_5013);
or U6255 (N_6255,N_4396,N_5060);
nand U6256 (N_6256,N_4280,N_5729);
and U6257 (N_6257,N_5286,N_5869);
and U6258 (N_6258,N_5087,N_4307);
nand U6259 (N_6259,N_5401,N_5089);
or U6260 (N_6260,N_5505,N_5335);
nand U6261 (N_6261,N_4242,N_5883);
nand U6262 (N_6262,N_5476,N_5253);
nand U6263 (N_6263,N_4991,N_5683);
nand U6264 (N_6264,N_5491,N_4053);
and U6265 (N_6265,N_4208,N_5898);
nor U6266 (N_6266,N_5086,N_4436);
and U6267 (N_6267,N_5396,N_4474);
nand U6268 (N_6268,N_5941,N_4229);
and U6269 (N_6269,N_5623,N_4360);
nor U6270 (N_6270,N_4989,N_4163);
nor U6271 (N_6271,N_5464,N_4686);
or U6272 (N_6272,N_5660,N_5472);
or U6273 (N_6273,N_5317,N_5096);
and U6274 (N_6274,N_5422,N_5183);
nand U6275 (N_6275,N_4092,N_4634);
nand U6276 (N_6276,N_4079,N_5151);
nor U6277 (N_6277,N_5842,N_4073);
nand U6278 (N_6278,N_5045,N_4610);
or U6279 (N_6279,N_4077,N_5139);
nand U6280 (N_6280,N_4102,N_4178);
and U6281 (N_6281,N_5890,N_5450);
xnor U6282 (N_6282,N_4752,N_5511);
nor U6283 (N_6283,N_4715,N_4111);
nand U6284 (N_6284,N_4529,N_5784);
nand U6285 (N_6285,N_4791,N_4405);
nor U6286 (N_6286,N_4313,N_5164);
nand U6287 (N_6287,N_4998,N_5646);
or U6288 (N_6288,N_4463,N_4024);
or U6289 (N_6289,N_4494,N_5915);
and U6290 (N_6290,N_5931,N_4450);
nor U6291 (N_6291,N_4720,N_4765);
nand U6292 (N_6292,N_4411,N_4872);
and U6293 (N_6293,N_5000,N_5606);
and U6294 (N_6294,N_4718,N_4502);
and U6295 (N_6295,N_5993,N_4052);
nor U6296 (N_6296,N_5173,N_4862);
nand U6297 (N_6297,N_4321,N_5659);
and U6298 (N_6298,N_5875,N_5545);
nand U6299 (N_6299,N_5582,N_4370);
nor U6300 (N_6300,N_4205,N_5269);
nor U6301 (N_6301,N_4112,N_4095);
and U6302 (N_6302,N_4143,N_5690);
and U6303 (N_6303,N_5431,N_5452);
nor U6304 (N_6304,N_4239,N_5810);
or U6305 (N_6305,N_4562,N_5481);
nor U6306 (N_6306,N_5374,N_5755);
or U6307 (N_6307,N_4714,N_4852);
nand U6308 (N_6308,N_4654,N_4259);
or U6309 (N_6309,N_4655,N_4552);
nand U6310 (N_6310,N_5939,N_4988);
nor U6311 (N_6311,N_5749,N_4664);
or U6312 (N_6312,N_4820,N_5642);
or U6313 (N_6313,N_5371,N_4138);
nor U6314 (N_6314,N_5373,N_4197);
and U6315 (N_6315,N_5549,N_5824);
nand U6316 (N_6316,N_5413,N_5161);
nor U6317 (N_6317,N_4609,N_4014);
nand U6318 (N_6318,N_4517,N_4061);
nand U6319 (N_6319,N_4054,N_5957);
nor U6320 (N_6320,N_4381,N_4585);
nand U6321 (N_6321,N_4974,N_4226);
nor U6322 (N_6322,N_4730,N_4546);
nand U6323 (N_6323,N_4469,N_4789);
nor U6324 (N_6324,N_5006,N_5526);
and U6325 (N_6325,N_4918,N_5242);
nand U6326 (N_6326,N_4188,N_5504);
or U6327 (N_6327,N_5719,N_4088);
nand U6328 (N_6328,N_5163,N_5411);
or U6329 (N_6329,N_5322,N_4798);
xnor U6330 (N_6330,N_4062,N_4476);
or U6331 (N_6331,N_5996,N_4866);
or U6332 (N_6332,N_5562,N_5621);
nor U6333 (N_6333,N_4508,N_4771);
or U6334 (N_6334,N_4953,N_4203);
nand U6335 (N_6335,N_5418,N_5300);
nor U6336 (N_6336,N_4050,N_4607);
or U6337 (N_6337,N_4754,N_5248);
or U6338 (N_6338,N_5840,N_4200);
xnor U6339 (N_6339,N_5134,N_4036);
or U6340 (N_6340,N_5596,N_4193);
nand U6341 (N_6341,N_4291,N_4554);
or U6342 (N_6342,N_5301,N_5694);
and U6343 (N_6343,N_4373,N_4149);
and U6344 (N_6344,N_4339,N_4884);
and U6345 (N_6345,N_4856,N_4948);
nor U6346 (N_6346,N_4954,N_5955);
or U6347 (N_6347,N_4990,N_4356);
nand U6348 (N_6348,N_4268,N_4303);
nand U6349 (N_6349,N_5929,N_4046);
and U6350 (N_6350,N_4165,N_4773);
and U6351 (N_6351,N_4772,N_4960);
nand U6352 (N_6352,N_5064,N_4029);
nor U6353 (N_6353,N_4199,N_4972);
or U6354 (N_6354,N_5554,N_4160);
and U6355 (N_6355,N_5745,N_5778);
or U6356 (N_6356,N_4946,N_5591);
and U6357 (N_6357,N_5636,N_4807);
nor U6358 (N_6358,N_4981,N_5891);
or U6359 (N_6359,N_4721,N_4462);
nor U6360 (N_6360,N_5341,N_4017);
nor U6361 (N_6361,N_4368,N_5699);
nor U6362 (N_6362,N_5035,N_5587);
nor U6363 (N_6363,N_5123,N_5215);
and U6364 (N_6364,N_4564,N_5172);
nand U6365 (N_6365,N_5907,N_5011);
and U6366 (N_6366,N_5031,N_5586);
or U6367 (N_6367,N_5912,N_4364);
or U6368 (N_6368,N_4711,N_5474);
or U6369 (N_6369,N_4725,N_5313);
nor U6370 (N_6370,N_5968,N_4258);
or U6371 (N_6371,N_4353,N_4175);
nand U6372 (N_6372,N_4995,N_4374);
and U6373 (N_6373,N_5153,N_4246);
or U6374 (N_6374,N_4749,N_4064);
or U6375 (N_6375,N_5303,N_5817);
and U6376 (N_6376,N_4434,N_4887);
and U6377 (N_6377,N_5160,N_5628);
nor U6378 (N_6378,N_5835,N_4317);
or U6379 (N_6379,N_5188,N_5393);
or U6380 (N_6380,N_5349,N_4290);
nor U6381 (N_6381,N_4542,N_5508);
or U6382 (N_6382,N_5843,N_5223);
nor U6383 (N_6383,N_5620,N_4254);
nor U6384 (N_6384,N_5130,N_5960);
and U6385 (N_6385,N_4376,N_5516);
and U6386 (N_6386,N_4247,N_5934);
nand U6387 (N_6387,N_5489,N_4986);
and U6388 (N_6388,N_5546,N_4745);
nor U6389 (N_6389,N_4501,N_4329);
and U6390 (N_6390,N_5004,N_5364);
and U6391 (N_6391,N_5753,N_5229);
nor U6392 (N_6392,N_4395,N_4084);
nand U6393 (N_6393,N_5460,N_4498);
and U6394 (N_6394,N_4125,N_5584);
nand U6395 (N_6395,N_4415,N_5781);
nand U6396 (N_6396,N_5066,N_5271);
or U6397 (N_6397,N_5882,N_4753);
and U6398 (N_6398,N_5856,N_4375);
xor U6399 (N_6399,N_5015,N_4727);
nand U6400 (N_6400,N_4157,N_5342);
nor U6401 (N_6401,N_5348,N_4548);
or U6402 (N_6402,N_5083,N_5009);
nand U6403 (N_6403,N_4764,N_4758);
nand U6404 (N_6404,N_5610,N_5964);
or U6405 (N_6405,N_4584,N_4018);
and U6406 (N_6406,N_5012,N_5617);
and U6407 (N_6407,N_4978,N_4827);
and U6408 (N_6408,N_4195,N_4164);
nand U6409 (N_6409,N_5576,N_4300);
nor U6410 (N_6410,N_4871,N_5944);
nor U6411 (N_6411,N_4000,N_4189);
or U6412 (N_6412,N_4456,N_5465);
nor U6413 (N_6413,N_5521,N_5273);
nor U6414 (N_6414,N_4127,N_5649);
and U6415 (N_6415,N_5189,N_5809);
and U6416 (N_6416,N_4096,N_4705);
nand U6417 (N_6417,N_4979,N_4185);
or U6418 (N_6418,N_4620,N_4059);
and U6419 (N_6419,N_4063,N_4580);
nor U6420 (N_6420,N_4646,N_4539);
xnor U6421 (N_6421,N_5042,N_5913);
or U6422 (N_6422,N_5696,N_5716);
nor U6423 (N_6423,N_5332,N_4470);
nand U6424 (N_6424,N_4662,N_5658);
or U6425 (N_6425,N_4997,N_5566);
nand U6426 (N_6426,N_4359,N_5007);
nand U6427 (N_6427,N_5100,N_4278);
or U6428 (N_6428,N_5697,N_5236);
nor U6429 (N_6429,N_5107,N_4348);
nor U6430 (N_6430,N_5397,N_4446);
and U6431 (N_6431,N_4184,N_4041);
and U6432 (N_6432,N_5711,N_5053);
or U6433 (N_6433,N_5792,N_4180);
nor U6434 (N_6434,N_4253,N_4615);
nor U6435 (N_6435,N_4802,N_4683);
nand U6436 (N_6436,N_5552,N_4666);
nor U6437 (N_6437,N_5558,N_4093);
and U6438 (N_6438,N_4262,N_5406);
or U6439 (N_6439,N_5029,N_5655);
and U6440 (N_6440,N_5094,N_4859);
or U6441 (N_6441,N_4146,N_4812);
nand U6442 (N_6442,N_5074,N_4331);
or U6443 (N_6443,N_4465,N_5909);
nand U6444 (N_6444,N_4845,N_4344);
nor U6445 (N_6445,N_4987,N_5555);
or U6446 (N_6446,N_5417,N_4644);
and U6447 (N_6447,N_5149,N_5951);
or U6448 (N_6448,N_5108,N_5145);
nor U6449 (N_6449,N_5085,N_4322);
nand U6450 (N_6450,N_4248,N_4597);
xnor U6451 (N_6451,N_4840,N_5919);
nor U6452 (N_6452,N_5228,N_4735);
nand U6453 (N_6453,N_4327,N_5794);
and U6454 (N_6454,N_5806,N_4222);
nor U6455 (N_6455,N_4377,N_5208);
or U6456 (N_6456,N_5258,N_4555);
or U6457 (N_6457,N_4403,N_4397);
and U6458 (N_6458,N_4975,N_4459);
nor U6459 (N_6459,N_5247,N_4518);
nor U6460 (N_6460,N_5434,N_4867);
and U6461 (N_6461,N_5082,N_4433);
and U6462 (N_6462,N_4905,N_5002);
nand U6463 (N_6463,N_5523,N_5722);
and U6464 (N_6464,N_5822,N_4171);
and U6465 (N_6465,N_4829,N_4581);
nand U6466 (N_6466,N_5598,N_5461);
and U6467 (N_6467,N_4440,N_5068);
or U6468 (N_6468,N_4003,N_5785);
and U6469 (N_6469,N_5469,N_5447);
and U6470 (N_6470,N_4283,N_5354);
and U6471 (N_6471,N_4496,N_4427);
nor U6472 (N_6472,N_4732,N_5977);
nor U6473 (N_6473,N_4047,N_5619);
nor U6474 (N_6474,N_4202,N_4390);
or U6475 (N_6475,N_4078,N_5632);
nor U6476 (N_6476,N_5924,N_4575);
or U6477 (N_6477,N_4500,N_4085);
and U6478 (N_6478,N_5618,N_5701);
or U6479 (N_6479,N_5725,N_4583);
or U6480 (N_6480,N_5016,N_4522);
and U6481 (N_6481,N_4726,N_5386);
nand U6482 (N_6482,N_5219,N_5976);
nor U6483 (N_6483,N_5026,N_4598);
and U6484 (N_6484,N_4287,N_4591);
and U6485 (N_6485,N_4621,N_5037);
nor U6486 (N_6486,N_5717,N_5240);
nor U6487 (N_6487,N_5664,N_4296);
or U6488 (N_6488,N_5359,N_5573);
or U6489 (N_6489,N_5132,N_5110);
or U6490 (N_6490,N_4318,N_4865);
nand U6491 (N_6491,N_4538,N_4419);
or U6492 (N_6492,N_5088,N_5166);
nor U6493 (N_6493,N_5005,N_5482);
or U6494 (N_6494,N_4934,N_5928);
and U6495 (N_6495,N_5231,N_4624);
or U6496 (N_6496,N_5574,N_4643);
or U6497 (N_6497,N_5412,N_4108);
nor U6498 (N_6498,N_4736,N_4523);
or U6499 (N_6499,N_4980,N_4068);
or U6500 (N_6500,N_4777,N_4145);
and U6501 (N_6501,N_5935,N_4209);
nor U6502 (N_6502,N_5639,N_5456);
or U6503 (N_6503,N_4593,N_5312);
xor U6504 (N_6504,N_4289,N_4451);
or U6505 (N_6505,N_4236,N_5302);
and U6506 (N_6506,N_4927,N_5947);
or U6507 (N_6507,N_4639,N_5136);
and U6508 (N_6508,N_5230,N_5276);
or U6509 (N_6509,N_4822,N_5295);
nand U6510 (N_6510,N_4961,N_5116);
and U6511 (N_6511,N_4889,N_4495);
or U6512 (N_6512,N_5114,N_4034);
and U6513 (N_6513,N_5863,N_4198);
nand U6514 (N_6514,N_5762,N_5686);
or U6515 (N_6515,N_5721,N_5266);
and U6516 (N_6516,N_5329,N_5075);
and U6517 (N_6517,N_5627,N_4486);
nor U6518 (N_6518,N_5485,N_5398);
nand U6519 (N_6519,N_4424,N_5185);
and U6520 (N_6520,N_4213,N_5908);
nor U6521 (N_6521,N_4642,N_4690);
or U6522 (N_6522,N_4439,N_5379);
nor U6523 (N_6523,N_5320,N_4306);
nand U6524 (N_6524,N_5877,N_5866);
or U6525 (N_6525,N_4635,N_4479);
nor U6526 (N_6526,N_5541,N_4454);
and U6527 (N_6527,N_5680,N_4612);
and U6528 (N_6528,N_4658,N_4818);
nor U6529 (N_6529,N_5056,N_5048);
nor U6530 (N_6530,N_4648,N_5868);
and U6531 (N_6531,N_4281,N_5760);
and U6532 (N_6532,N_5527,N_5881);
nand U6533 (N_6533,N_5090,N_4605);
or U6534 (N_6534,N_4669,N_5220);
or U6535 (N_6535,N_5922,N_4288);
and U6536 (N_6536,N_4483,N_4724);
and U6537 (N_6537,N_4803,N_4958);
nor U6538 (N_6538,N_5375,N_5440);
nand U6539 (N_6539,N_4950,N_4779);
and U6540 (N_6540,N_5076,N_5360);
nor U6541 (N_6541,N_5119,N_4314);
nor U6542 (N_6542,N_5167,N_5685);
nor U6543 (N_6543,N_4269,N_4480);
nor U6544 (N_6544,N_4270,N_4423);
nand U6545 (N_6545,N_4556,N_5724);
and U6546 (N_6546,N_5695,N_5888);
nand U6547 (N_6547,N_5017,N_4768);
nor U6548 (N_6548,N_5616,N_5299);
nand U6549 (N_6549,N_4874,N_5243);
nor U6550 (N_6550,N_4842,N_5314);
nand U6551 (N_6551,N_5356,N_5651);
nand U6552 (N_6552,N_4275,N_5992);
nor U6553 (N_6553,N_4147,N_5512);
nand U6554 (N_6554,N_4781,N_5715);
or U6555 (N_6555,N_5971,N_4094);
nor U6556 (N_6556,N_5459,N_5933);
nand U6557 (N_6557,N_5949,N_4035);
nand U6558 (N_6558,N_4432,N_4315);
nor U6559 (N_6559,N_4295,N_5874);
nor U6560 (N_6560,N_5287,N_4767);
or U6561 (N_6561,N_4579,N_4345);
nor U6562 (N_6562,N_4616,N_4493);
and U6563 (N_6563,N_5671,N_5203);
and U6564 (N_6564,N_5471,N_4484);
or U6565 (N_6565,N_4086,N_4534);
nor U6566 (N_6566,N_4101,N_5501);
nand U6567 (N_6567,N_4628,N_4739);
nand U6568 (N_6568,N_5823,N_4659);
or U6569 (N_6569,N_5186,N_4223);
nor U6570 (N_6570,N_5837,N_5864);
and U6571 (N_6571,N_5848,N_5921);
or U6572 (N_6572,N_4429,N_5672);
or U6573 (N_6573,N_4863,N_5846);
and U6574 (N_6574,N_5008,N_4182);
nand U6575 (N_6575,N_4841,N_5544);
or U6576 (N_6576,N_4627,N_4234);
nor U6577 (N_6577,N_5973,N_4022);
nor U6578 (N_6578,N_4614,N_5347);
nor U6579 (N_6579,N_5280,N_5599);
nand U6580 (N_6580,N_5688,N_5743);
or U6581 (N_6581,N_5950,N_4592);
nor U6582 (N_6582,N_4074,N_5475);
and U6583 (N_6583,N_5389,N_5532);
nor U6584 (N_6584,N_4746,N_5990);
nor U6585 (N_6585,N_5277,N_5070);
nor U6586 (N_6586,N_4430,N_4244);
and U6587 (N_6587,N_4857,N_5032);
and U6588 (N_6588,N_5473,N_5926);
nor U6589 (N_6589,N_4008,N_5445);
or U6590 (N_6590,N_5370,N_4115);
nand U6591 (N_6591,N_4831,N_5917);
nor U6592 (N_6592,N_5346,N_4191);
nand U6593 (N_6593,N_5588,N_4380);
nor U6594 (N_6594,N_5849,N_4660);
and U6595 (N_6595,N_4201,N_5804);
nor U6596 (N_6596,N_4793,N_5536);
or U6597 (N_6597,N_5438,N_5122);
nor U6598 (N_6598,N_4033,N_4969);
nand U6599 (N_6599,N_5020,N_4770);
nor U6600 (N_6600,N_5380,N_4709);
and U6601 (N_6601,N_5997,N_5629);
nand U6602 (N_6602,N_4187,N_5624);
nand U6603 (N_6603,N_5897,N_4741);
nand U6604 (N_6604,N_5435,N_5633);
or U6605 (N_6605,N_4218,N_5535);
nor U6606 (N_6606,N_4181,N_4769);
and U6607 (N_6607,N_4511,N_5125);
or U6608 (N_6608,N_5638,N_5150);
or U6609 (N_6609,N_4606,N_5713);
and U6610 (N_6610,N_5241,N_4689);
nand U6611 (N_6611,N_4025,N_5816);
nor U6612 (N_6612,N_4384,N_4304);
nor U6613 (N_6613,N_4601,N_5078);
nand U6614 (N_6614,N_4362,N_5442);
nor U6615 (N_6615,N_5137,N_4537);
and U6616 (N_6616,N_4420,N_5255);
xnor U6617 (N_6617,N_5344,N_4134);
and U6618 (N_6618,N_5878,N_5826);
nand U6619 (N_6619,N_4507,N_4963);
nor U6620 (N_6620,N_4250,N_4249);
and U6621 (N_6621,N_5421,N_5147);
nor U6622 (N_6622,N_5567,N_4312);
or U6623 (N_6623,N_4482,N_5495);
nand U6624 (N_6624,N_5988,N_4013);
and U6625 (N_6625,N_4336,N_4923);
or U6626 (N_6626,N_5079,N_5428);
and U6627 (N_6627,N_5798,N_5333);
and U6628 (N_6628,N_4285,N_5191);
nor U6629 (N_6629,N_5594,N_5853);
nand U6630 (N_6630,N_5140,N_4738);
nand U6631 (N_6631,N_5528,N_5987);
or U6632 (N_6632,N_5630,N_4421);
or U6633 (N_6633,N_4369,N_5563);
nand U6634 (N_6634,N_4332,N_5159);
nand U6635 (N_6635,N_5260,N_4524);
or U6636 (N_6636,N_4673,N_5270);
or U6637 (N_6637,N_4833,N_5288);
or U6638 (N_6638,N_5385,N_5510);
nand U6639 (N_6639,N_5518,N_4478);
nor U6640 (N_6640,N_4886,N_4334);
nor U6641 (N_6641,N_5376,N_4335);
and U6642 (N_6642,N_5158,N_4028);
nand U6643 (N_6643,N_5334,N_4404);
and U6644 (N_6644,N_4596,N_5387);
or U6645 (N_6645,N_5479,N_4712);
nand U6646 (N_6646,N_5135,N_5692);
and U6647 (N_6647,N_5940,N_5404);
nand U6648 (N_6648,N_4097,N_5614);
nand U6649 (N_6649,N_4266,N_4786);
or U6650 (N_6650,N_4839,N_5542);
or U6651 (N_6651,N_4408,N_4574);
and U6652 (N_6652,N_5611,N_5911);
or U6653 (N_6653,N_4109,N_5793);
and U6654 (N_6654,N_5657,N_5378);
nand U6655 (N_6655,N_4528,N_4902);
and U6656 (N_6656,N_4105,N_4563);
nand U6657 (N_6657,N_5104,N_5640);
nand U6658 (N_6658,N_5962,N_5028);
and U6659 (N_6659,N_4243,N_5872);
nor U6660 (N_6660,N_5439,N_5275);
nand U6661 (N_6661,N_5954,N_5285);
nand U6662 (N_6662,N_4630,N_4519);
or U6663 (N_6663,N_5429,N_5942);
and U6664 (N_6664,N_5169,N_5771);
or U6665 (N_6665,N_5290,N_4778);
and U6666 (N_6666,N_5580,N_4506);
and U6667 (N_6667,N_4039,N_4080);
nand U6668 (N_6668,N_4333,N_4696);
or U6669 (N_6669,N_4066,N_4814);
nand U6670 (N_6670,N_5813,N_4264);
and U6671 (N_6671,N_5653,N_5024);
nand U6672 (N_6672,N_5261,N_5262);
or U6673 (N_6673,N_5534,N_5432);
and U6674 (N_6674,N_5043,N_5969);
nand U6675 (N_6675,N_5787,N_5705);
nand U6676 (N_6676,N_5050,N_5307);
and U6677 (N_6677,N_4649,N_5607);
or U6678 (N_6678,N_4497,N_5003);
nor U6679 (N_6679,N_4087,N_4512);
nor U6680 (N_6680,N_5779,N_5410);
and U6681 (N_6681,N_4123,N_5138);
and U6682 (N_6682,N_5986,N_5679);
nor U6683 (N_6683,N_5763,N_4549);
and U6684 (N_6684,N_5168,N_4944);
or U6685 (N_6685,N_4277,N_5238);
and U6686 (N_6686,N_4657,N_5650);
or U6687 (N_6687,N_5443,N_5827);
nand U6688 (N_6688,N_4900,N_5775);
nand U6689 (N_6689,N_4385,N_5731);
nor U6690 (N_6690,N_4358,N_4341);
xor U6691 (N_6691,N_4516,N_4210);
nand U6692 (N_6692,N_5001,N_5216);
nor U6693 (N_6693,N_5867,N_4392);
and U6694 (N_6694,N_4569,N_4032);
and U6695 (N_6695,N_5570,N_4015);
or U6696 (N_6696,N_4057,N_5506);
nor U6697 (N_6697,N_5457,N_4903);
xnor U6698 (N_6698,N_5847,N_5023);
and U6699 (N_6699,N_4186,N_5645);
and U6700 (N_6700,N_4354,N_5865);
nand U6701 (N_6701,N_4920,N_5970);
nor U6702 (N_6702,N_4113,N_5407);
and U6703 (N_6703,N_4007,N_4545);
or U6704 (N_6704,N_4586,N_4847);
and U6705 (N_6705,N_4892,N_5041);
and U6706 (N_6706,N_4350,N_5795);
or U6707 (N_6707,N_4179,N_5127);
nand U6708 (N_6708,N_4120,N_4956);
nand U6709 (N_6709,N_5667,N_4797);
or U6710 (N_6710,N_5648,N_5463);
nor U6711 (N_6711,N_4895,N_4697);
nor U6712 (N_6712,N_4731,N_4701);
or U6713 (N_6713,N_5492,N_5777);
or U6714 (N_6714,N_5770,N_5366);
and U6715 (N_6715,N_5681,N_4921);
or U6716 (N_6716,N_5202,N_4402);
nor U6717 (N_6717,N_5901,N_5427);
and U6718 (N_6718,N_4932,N_5597);
or U6719 (N_6719,N_5712,N_5264);
or U6720 (N_6720,N_4756,N_5807);
or U6721 (N_6721,N_5257,N_5178);
and U6722 (N_6722,N_4286,N_4162);
nand U6723 (N_6723,N_4794,N_5768);
nand U6724 (N_6724,N_5484,N_5538);
nor U6725 (N_6725,N_5839,N_4464);
or U6726 (N_6726,N_4449,N_5493);
or U6727 (N_6727,N_5430,N_5181);
nor U6728 (N_6728,N_5780,N_5499);
and U6729 (N_6729,N_5953,N_5361);
and U6730 (N_6730,N_5899,N_4401);
nor U6731 (N_6731,N_4144,N_5698);
and U6732 (N_6732,N_4551,N_5497);
or U6733 (N_6733,N_4299,N_4361);
or U6734 (N_6734,N_4925,N_5274);
nor U6735 (N_6735,N_5786,N_4407);
nor U6736 (N_6736,N_5316,N_4834);
nand U6737 (N_6737,N_5444,N_5728);
and U6738 (N_6738,N_4894,N_5613);
and U6739 (N_6739,N_4227,N_4316);
nor U6740 (N_6740,N_4214,N_4005);
nor U6741 (N_6741,N_4638,N_4985);
and U6742 (N_6742,N_5369,N_5502);
nor U6743 (N_6743,N_5263,N_4668);
nand U6744 (N_6744,N_4475,N_4676);
nor U6745 (N_6745,N_4090,N_4128);
nand U6746 (N_6746,N_5331,N_4016);
and U6747 (N_6747,N_4399,N_4792);
or U6748 (N_6748,N_5734,N_4265);
nor U6749 (N_6749,N_4878,N_5747);
nand U6750 (N_6750,N_4858,N_5466);
and U6751 (N_6751,N_4907,N_4733);
and U6752 (N_6752,N_5483,N_5372);
or U6753 (N_6753,N_4811,N_4383);
xnor U6754 (N_6754,N_5030,N_4603);
or U6755 (N_6755,N_5884,N_5470);
and U6756 (N_6756,N_4846,N_4742);
or U6757 (N_6757,N_4412,N_4056);
and U6758 (N_6758,N_4901,N_4156);
nor U6759 (N_6759,N_5703,N_4467);
nor U6760 (N_6760,N_5765,N_5989);
or U6761 (N_6761,N_4882,N_4159);
nor U6762 (N_6762,N_4196,N_4774);
nor U6763 (N_6763,N_5666,N_4126);
nand U6764 (N_6764,N_4400,N_4893);
nand U6765 (N_6765,N_4413,N_5603);
nand U6766 (N_6766,N_5256,N_5952);
xor U6767 (N_6767,N_5652,N_4799);
nor U6768 (N_6768,N_5741,N_4588);
nand U6769 (N_6769,N_4142,N_4566);
nand U6770 (N_6770,N_4936,N_5985);
and U6771 (N_6771,N_4728,N_5769);
or U6772 (N_6772,N_5923,N_5298);
or U6773 (N_6773,N_5676,N_5105);
or U6774 (N_6774,N_4964,N_5821);
or U6775 (N_6775,N_5520,N_4544);
nand U6776 (N_6776,N_5106,N_4256);
or U6777 (N_6777,N_5279,N_4042);
and U6778 (N_6778,N_5836,N_5800);
and U6779 (N_6779,N_4488,N_5494);
or U6780 (N_6780,N_5152,N_5684);
or U6781 (N_6781,N_5991,N_4472);
or U6782 (N_6782,N_5175,N_4570);
or U6783 (N_6783,N_4817,N_5906);
nand U6784 (N_6784,N_5323,N_4292);
nor U6785 (N_6785,N_5394,N_5059);
or U6786 (N_6786,N_4104,N_5319);
nor U6787 (N_6787,N_4070,N_5663);
nor U6788 (N_6788,N_4873,N_4853);
or U6789 (N_6789,N_4531,N_5338);
and U6790 (N_6790,N_4836,N_5974);
nand U6791 (N_6791,N_5748,N_5547);
or U6792 (N_6792,N_4795,N_5325);
nand U6793 (N_6793,N_4647,N_4363);
and U6794 (N_6794,N_4533,N_4293);
nor U6795 (N_6795,N_4929,N_4684);
nand U6796 (N_6796,N_5437,N_5467);
or U6797 (N_6797,N_5155,N_4717);
and U6798 (N_6798,N_4617,N_4338);
or U6799 (N_6799,N_4844,N_4442);
or U6800 (N_6800,N_4631,N_5844);
nand U6801 (N_6801,N_5736,N_5548);
nand U6802 (N_6802,N_4155,N_5148);
or U6803 (N_6803,N_4868,N_4252);
nand U6804 (N_6804,N_5062,N_5980);
nand U6805 (N_6805,N_4212,N_4908);
nor U6806 (N_6806,N_5478,N_5343);
or U6807 (N_6807,N_5453,N_5080);
nand U6808 (N_6808,N_4966,N_4626);
nand U6809 (N_6809,N_5327,N_5034);
nor U6810 (N_6810,N_5852,N_4573);
or U6811 (N_6811,N_5121,N_4550);
or U6812 (N_6812,N_4158,N_5910);
nand U6813 (N_6813,N_5311,N_5328);
and U6814 (N_6814,N_4951,N_5221);
or U6815 (N_6815,N_5498,N_5509);
or U6816 (N_6816,N_5517,N_4881);
nor U6817 (N_6817,N_5513,N_5811);
nand U6818 (N_6818,N_4418,N_4667);
nand U6819 (N_6819,N_5377,N_4267);
and U6820 (N_6820,N_4861,N_4037);
or U6821 (N_6821,N_4466,N_5049);
nor U6822 (N_6822,N_4425,N_4103);
nand U6823 (N_6823,N_5446,N_4216);
nand U6824 (N_6824,N_5310,N_5156);
nand U6825 (N_6825,N_4568,N_5662);
or U6826 (N_6826,N_4808,N_4357);
nor U6827 (N_6827,N_4940,N_4809);
nor U6828 (N_6828,N_5282,N_5200);
or U6829 (N_6829,N_4447,N_4983);
or U6830 (N_6830,N_4801,N_4098);
or U6831 (N_6831,N_5069,N_5400);
or U6832 (N_6832,N_5818,N_5693);
or U6833 (N_6833,N_4135,N_4019);
nand U6834 (N_6834,N_5176,N_4561);
or U6835 (N_6835,N_4460,N_4473);
nand U6836 (N_6836,N_4959,N_5177);
nand U6837 (N_6837,N_5831,N_4578);
nor U6838 (N_6838,N_5345,N_4067);
nor U6839 (N_6839,N_4461,N_5126);
nand U6840 (N_6840,N_5353,N_5790);
nand U6841 (N_6841,N_4870,N_5201);
or U6842 (N_6842,N_4869,N_5381);
or U6843 (N_6843,N_4441,N_4238);
nand U6844 (N_6844,N_4716,N_5937);
and U6845 (N_6845,N_4055,N_4898);
and U6846 (N_6846,N_4294,N_5281);
or U6847 (N_6847,N_5436,N_5522);
or U6848 (N_6848,N_4219,N_4623);
nand U6849 (N_6849,N_5982,N_4352);
nand U6850 (N_6850,N_5553,N_4257);
and U6851 (N_6851,N_4850,N_5845);
and U6852 (N_6852,N_4394,N_4011);
nor U6853 (N_6853,N_4952,N_4825);
and U6854 (N_6854,N_5101,N_5357);
and U6855 (N_6855,N_5018,N_5766);
or U6856 (N_6856,N_5044,N_5441);
nand U6857 (N_6857,N_5365,N_5637);
and U6858 (N_6858,N_4992,N_5665);
nor U6859 (N_6859,N_5102,N_5959);
xnor U6860 (N_6860,N_5352,N_5025);
nor U6861 (N_6861,N_4340,N_4391);
and U6862 (N_6862,N_5564,N_5936);
nor U6863 (N_6863,N_5462,N_5384);
and U6864 (N_6864,N_4452,N_5995);
and U6865 (N_6865,N_4058,N_5326);
or U6866 (N_6866,N_5330,N_5978);
and U6867 (N_6867,N_5052,N_5047);
nor U6868 (N_6868,N_4748,N_4880);
and U6869 (N_6869,N_4365,N_4729);
nand U6870 (N_6870,N_4663,N_5689);
nor U6871 (N_6871,N_5196,N_4477);
and U6872 (N_6872,N_4744,N_5051);
nand U6873 (N_6873,N_4021,N_4137);
or U6874 (N_6874,N_4999,N_4177);
nor U6875 (N_6875,N_4301,N_4737);
nor U6876 (N_6876,N_4977,N_4692);
nor U6877 (N_6877,N_4153,N_5861);
nor U6878 (N_6878,N_5860,N_4490);
and U6879 (N_6879,N_4650,N_4937);
nand U6880 (N_6880,N_4273,N_5306);
nor U6881 (N_6881,N_4681,N_5097);
and U6882 (N_6882,N_4489,N_5390);
and U6883 (N_6883,N_5757,N_5197);
or U6884 (N_6884,N_5214,N_4750);
or U6885 (N_6885,N_4245,N_5232);
nand U6886 (N_6886,N_5142,N_5578);
or U6887 (N_6887,N_4001,N_4919);
and U6888 (N_6888,N_5180,N_4888);
or U6889 (N_6889,N_5551,N_5710);
nand U6890 (N_6890,N_4311,N_5291);
nand U6891 (N_6891,N_5819,N_5876);
xnor U6892 (N_6892,N_4235,N_5925);
or U6893 (N_6893,N_4885,N_4896);
nor U6894 (N_6894,N_5612,N_4133);
nand U6895 (N_6895,N_4804,N_5647);
nor U6896 (N_6896,N_5718,N_5490);
or U6897 (N_6897,N_5789,N_5801);
and U6898 (N_6898,N_5669,N_4152);
and U6899 (N_6899,N_5855,N_4141);
and U6900 (N_6900,N_4938,N_4468);
nand U6901 (N_6901,N_4319,N_5550);
nor U6902 (N_6902,N_4491,N_4224);
nand U6903 (N_6903,N_5480,N_4572);
and U6904 (N_6904,N_4513,N_4824);
nand U6905 (N_6905,N_5144,N_5294);
nor U6906 (N_6906,N_4347,N_5902);
nor U6907 (N_6907,N_4148,N_4343);
and U6908 (N_6908,N_4677,N_4136);
nor U6909 (N_6909,N_4261,N_4378);
and U6910 (N_6910,N_4069,N_5783);
nand U6911 (N_6911,N_4587,N_5761);
and U6912 (N_6912,N_5213,N_4719);
nand U6913 (N_6913,N_4645,N_4492);
nor U6914 (N_6914,N_4694,N_4851);
and U6915 (N_6915,N_5583,N_4637);
and U6916 (N_6916,N_5707,N_4438);
nor U6917 (N_6917,N_4328,N_5309);
and U6918 (N_6918,N_5448,N_4984);
and U6919 (N_6919,N_4305,N_4641);
nand U6920 (N_6920,N_5533,N_4505);
nor U6921 (N_6921,N_5870,N_5211);
nand U6922 (N_6922,N_4276,N_4437);
nor U6923 (N_6923,N_4140,N_4935);
or U6924 (N_6924,N_5751,N_4823);
and U6925 (N_6925,N_4100,N_4955);
nand U6926 (N_6926,N_5825,N_4875);
nor U6927 (N_6927,N_5656,N_5193);
nor U6928 (N_6928,N_5626,N_5245);
or U6929 (N_6929,N_5966,N_5858);
nand U6930 (N_6930,N_4913,N_5204);
nor U6931 (N_6931,N_4194,N_5190);
or U6932 (N_6932,N_5561,N_4899);
nor U6933 (N_6933,N_4700,N_4428);
nor U6934 (N_6934,N_4702,N_4526);
and U6935 (N_6935,N_4130,N_5362);
nand U6936 (N_6936,N_5961,N_5318);
nand U6937 (N_6937,N_4704,N_5880);
nand U6938 (N_6938,N_4618,N_4837);
nor U6939 (N_6939,N_4170,N_5774);
nor U6940 (N_6940,N_4044,N_5289);
nor U6941 (N_6941,N_5998,N_4761);
and U6942 (N_6942,N_4387,N_5668);
or U6943 (N_6943,N_5133,N_4565);
and U6944 (N_6944,N_4968,N_5425);
xor U6945 (N_6945,N_4499,N_4915);
and U6946 (N_6946,N_5278,N_5244);
or U6947 (N_6947,N_4993,N_5585);
nand U6948 (N_6948,N_4509,N_4571);
nand U6949 (N_6949,N_5249,N_4707);
nor U6950 (N_6950,N_5893,N_5920);
and U6951 (N_6951,N_5409,N_5308);
nor U6952 (N_6952,N_5975,N_5687);
nor U6953 (N_6953,N_5065,N_4943);
nand U6954 (N_6954,N_5857,N_5850);
or U6955 (N_6955,N_4740,N_5525);
nor U6956 (N_6956,N_4910,N_4026);
nor U6957 (N_6957,N_4217,N_4325);
or U6958 (N_6958,N_5112,N_5239);
and U6959 (N_6959,N_4284,N_5622);
xnor U6960 (N_6960,N_5395,N_4326);
and U6961 (N_6961,N_5967,N_4594);
nand U6962 (N_6962,N_4443,N_5124);
or U6963 (N_6963,N_5581,N_5038);
or U6964 (N_6964,N_5337,N_5691);
nand U6965 (N_6965,N_4083,N_5644);
and U6966 (N_6966,N_4525,N_5027);
and U6967 (N_6967,N_4695,N_5234);
and U6968 (N_6968,N_4661,N_5120);
nand U6969 (N_6969,N_5351,N_4541);
and U6970 (N_6970,N_4805,N_4237);
nor U6971 (N_6971,N_4914,N_5841);
and U6972 (N_6972,N_4167,N_5179);
and U6973 (N_6973,N_5529,N_4933);
and U6974 (N_6974,N_5589,N_4928);
or U6975 (N_6975,N_4957,N_4485);
nor U6976 (N_6976,N_4045,N_4790);
nand U6977 (N_6977,N_4031,N_4065);
nand U6978 (N_6978,N_4076,N_5805);
or U6979 (N_6979,N_4890,N_5225);
or U6980 (N_6980,N_4417,N_4939);
or U6981 (N_6981,N_4255,N_5154);
nand U6982 (N_6982,N_5267,N_4685);
nor U6983 (N_6983,N_4228,N_5577);
or U6984 (N_6984,N_4346,N_5117);
nor U6985 (N_6985,N_5118,N_5099);
xnor U6986 (N_6986,N_5250,N_4604);
or U6987 (N_6987,N_4471,N_4942);
nand U6988 (N_6988,N_4371,N_4757);
nor U6989 (N_6989,N_5738,N_5706);
nand U6990 (N_6990,N_5758,N_4458);
nand U6991 (N_6991,N_4233,N_5063);
and U6992 (N_6992,N_4520,N_5072);
and U6993 (N_6993,N_5251,N_4931);
nand U6994 (N_6994,N_4651,N_4595);
or U6995 (N_6995,N_4535,N_5830);
nor U6996 (N_6996,N_5383,N_4582);
and U6997 (N_6997,N_4577,N_5315);
nor U6998 (N_6998,N_5222,N_5174);
or U6999 (N_6999,N_4629,N_4706);
nor U7000 (N_7000,N_4714,N_4587);
and U7001 (N_7001,N_5006,N_5463);
and U7002 (N_7002,N_5502,N_4625);
and U7003 (N_7003,N_5736,N_5401);
nor U7004 (N_7004,N_5911,N_4146);
or U7005 (N_7005,N_4625,N_5252);
nor U7006 (N_7006,N_5126,N_4290);
nand U7007 (N_7007,N_4929,N_4277);
nand U7008 (N_7008,N_5053,N_5823);
nand U7009 (N_7009,N_5222,N_5701);
or U7010 (N_7010,N_4016,N_4166);
nor U7011 (N_7011,N_4104,N_4965);
nand U7012 (N_7012,N_4611,N_4171);
nor U7013 (N_7013,N_5568,N_5255);
nor U7014 (N_7014,N_5203,N_5405);
nand U7015 (N_7015,N_4201,N_4280);
nor U7016 (N_7016,N_5882,N_4691);
or U7017 (N_7017,N_5653,N_4182);
nor U7018 (N_7018,N_4259,N_5147);
or U7019 (N_7019,N_5024,N_5747);
nand U7020 (N_7020,N_5053,N_5313);
nand U7021 (N_7021,N_4537,N_4084);
nand U7022 (N_7022,N_5652,N_5414);
nand U7023 (N_7023,N_4242,N_4188);
nand U7024 (N_7024,N_4966,N_4475);
nand U7025 (N_7025,N_4323,N_5144);
and U7026 (N_7026,N_5881,N_5251);
or U7027 (N_7027,N_5810,N_5299);
nand U7028 (N_7028,N_4937,N_5076);
nand U7029 (N_7029,N_5195,N_5761);
and U7030 (N_7030,N_5267,N_5690);
and U7031 (N_7031,N_4962,N_4396);
and U7032 (N_7032,N_5457,N_5644);
xnor U7033 (N_7033,N_4506,N_4475);
or U7034 (N_7034,N_5916,N_5371);
and U7035 (N_7035,N_5862,N_5844);
or U7036 (N_7036,N_5422,N_4189);
or U7037 (N_7037,N_4896,N_4542);
nor U7038 (N_7038,N_4319,N_4595);
and U7039 (N_7039,N_4847,N_5100);
nand U7040 (N_7040,N_4852,N_5309);
nor U7041 (N_7041,N_5318,N_5423);
or U7042 (N_7042,N_5807,N_4221);
or U7043 (N_7043,N_4494,N_5142);
xnor U7044 (N_7044,N_5791,N_5581);
and U7045 (N_7045,N_4260,N_5721);
nand U7046 (N_7046,N_5651,N_4045);
nand U7047 (N_7047,N_5006,N_4300);
nand U7048 (N_7048,N_5651,N_4682);
or U7049 (N_7049,N_4480,N_4080);
or U7050 (N_7050,N_4444,N_5364);
and U7051 (N_7051,N_4048,N_5158);
or U7052 (N_7052,N_4214,N_4433);
nand U7053 (N_7053,N_4160,N_5951);
and U7054 (N_7054,N_4945,N_5950);
and U7055 (N_7055,N_5857,N_5448);
and U7056 (N_7056,N_5789,N_5674);
nor U7057 (N_7057,N_4490,N_5230);
or U7058 (N_7058,N_4389,N_5129);
and U7059 (N_7059,N_5992,N_5726);
and U7060 (N_7060,N_5036,N_4781);
or U7061 (N_7061,N_5439,N_4571);
and U7062 (N_7062,N_5458,N_4113);
nor U7063 (N_7063,N_4249,N_4092);
and U7064 (N_7064,N_4281,N_4868);
and U7065 (N_7065,N_5848,N_4635);
nor U7066 (N_7066,N_5914,N_5411);
and U7067 (N_7067,N_4159,N_5707);
nor U7068 (N_7068,N_4810,N_5389);
nor U7069 (N_7069,N_4225,N_5585);
nand U7070 (N_7070,N_4959,N_5186);
or U7071 (N_7071,N_4244,N_5549);
and U7072 (N_7072,N_5040,N_5850);
or U7073 (N_7073,N_5760,N_5931);
or U7074 (N_7074,N_4648,N_4829);
nand U7075 (N_7075,N_5627,N_5824);
nor U7076 (N_7076,N_4123,N_5862);
nand U7077 (N_7077,N_5176,N_5538);
or U7078 (N_7078,N_4534,N_5894);
nor U7079 (N_7079,N_5829,N_4205);
and U7080 (N_7080,N_4884,N_4981);
nand U7081 (N_7081,N_4985,N_5844);
nand U7082 (N_7082,N_4691,N_5251);
nand U7083 (N_7083,N_4789,N_4909);
nor U7084 (N_7084,N_4263,N_4214);
and U7085 (N_7085,N_4178,N_5327);
nor U7086 (N_7086,N_4782,N_4771);
or U7087 (N_7087,N_5715,N_4866);
nand U7088 (N_7088,N_4188,N_4967);
and U7089 (N_7089,N_4653,N_4273);
nand U7090 (N_7090,N_5560,N_5729);
nand U7091 (N_7091,N_4230,N_4922);
nand U7092 (N_7092,N_4696,N_4288);
nor U7093 (N_7093,N_4227,N_5042);
nand U7094 (N_7094,N_5733,N_5802);
nand U7095 (N_7095,N_4292,N_4165);
nor U7096 (N_7096,N_5938,N_4744);
nor U7097 (N_7097,N_4282,N_4710);
nand U7098 (N_7098,N_4547,N_4045);
and U7099 (N_7099,N_5741,N_4002);
nand U7100 (N_7100,N_5801,N_5541);
or U7101 (N_7101,N_4968,N_5489);
nor U7102 (N_7102,N_4957,N_5889);
nor U7103 (N_7103,N_5161,N_4191);
and U7104 (N_7104,N_4052,N_4803);
or U7105 (N_7105,N_5269,N_5584);
nand U7106 (N_7106,N_5086,N_4349);
nor U7107 (N_7107,N_4992,N_5769);
nor U7108 (N_7108,N_5753,N_5134);
and U7109 (N_7109,N_5993,N_5690);
and U7110 (N_7110,N_4817,N_4166);
or U7111 (N_7111,N_5724,N_4052);
and U7112 (N_7112,N_5456,N_5154);
nand U7113 (N_7113,N_4865,N_5457);
or U7114 (N_7114,N_4491,N_5183);
or U7115 (N_7115,N_5073,N_4119);
xnor U7116 (N_7116,N_4833,N_5754);
and U7117 (N_7117,N_4654,N_4766);
nand U7118 (N_7118,N_5508,N_4676);
nand U7119 (N_7119,N_5915,N_5673);
and U7120 (N_7120,N_4949,N_5160);
nand U7121 (N_7121,N_5666,N_4294);
nor U7122 (N_7122,N_4236,N_4350);
nand U7123 (N_7123,N_5647,N_5250);
and U7124 (N_7124,N_4933,N_5943);
and U7125 (N_7125,N_5719,N_4852);
and U7126 (N_7126,N_5936,N_4265);
nor U7127 (N_7127,N_5960,N_5836);
and U7128 (N_7128,N_4963,N_4022);
nor U7129 (N_7129,N_4761,N_4110);
nor U7130 (N_7130,N_4634,N_4063);
or U7131 (N_7131,N_4568,N_4329);
and U7132 (N_7132,N_4491,N_4180);
or U7133 (N_7133,N_4758,N_5957);
or U7134 (N_7134,N_4230,N_4706);
nand U7135 (N_7135,N_4133,N_5652);
and U7136 (N_7136,N_5911,N_5805);
nand U7137 (N_7137,N_5499,N_4471);
nor U7138 (N_7138,N_5993,N_5122);
nor U7139 (N_7139,N_4438,N_5545);
nor U7140 (N_7140,N_5230,N_4947);
nor U7141 (N_7141,N_4082,N_4457);
and U7142 (N_7142,N_4337,N_4612);
or U7143 (N_7143,N_5256,N_4369);
nor U7144 (N_7144,N_5115,N_4050);
or U7145 (N_7145,N_5648,N_5555);
or U7146 (N_7146,N_4961,N_5826);
nand U7147 (N_7147,N_4539,N_5891);
nand U7148 (N_7148,N_5761,N_4867);
nor U7149 (N_7149,N_5114,N_4218);
nand U7150 (N_7150,N_4611,N_4427);
nand U7151 (N_7151,N_5182,N_5016);
nor U7152 (N_7152,N_5972,N_4185);
and U7153 (N_7153,N_4003,N_4743);
nand U7154 (N_7154,N_5200,N_4621);
or U7155 (N_7155,N_5771,N_4371);
or U7156 (N_7156,N_4703,N_4158);
nor U7157 (N_7157,N_4755,N_5436);
or U7158 (N_7158,N_5193,N_5407);
and U7159 (N_7159,N_5360,N_4917);
nor U7160 (N_7160,N_5391,N_4810);
nand U7161 (N_7161,N_4322,N_4589);
nor U7162 (N_7162,N_5690,N_5892);
nor U7163 (N_7163,N_5920,N_5337);
or U7164 (N_7164,N_5765,N_5034);
nand U7165 (N_7165,N_5677,N_5902);
nand U7166 (N_7166,N_4866,N_4349);
and U7167 (N_7167,N_5054,N_5989);
nor U7168 (N_7168,N_4602,N_5728);
nor U7169 (N_7169,N_5096,N_5945);
or U7170 (N_7170,N_5859,N_4696);
nand U7171 (N_7171,N_5145,N_5645);
or U7172 (N_7172,N_4794,N_4159);
nor U7173 (N_7173,N_5858,N_4074);
and U7174 (N_7174,N_5073,N_5594);
nor U7175 (N_7175,N_5210,N_4630);
nor U7176 (N_7176,N_4667,N_5700);
or U7177 (N_7177,N_5691,N_5124);
nand U7178 (N_7178,N_5871,N_4135);
nand U7179 (N_7179,N_5623,N_5541);
nand U7180 (N_7180,N_5717,N_5051);
nor U7181 (N_7181,N_5795,N_5199);
or U7182 (N_7182,N_4926,N_4161);
nand U7183 (N_7183,N_4113,N_5337);
and U7184 (N_7184,N_4966,N_5700);
nor U7185 (N_7185,N_5976,N_4564);
or U7186 (N_7186,N_4662,N_4350);
nor U7187 (N_7187,N_4869,N_5700);
nand U7188 (N_7188,N_5577,N_4566);
and U7189 (N_7189,N_4401,N_4753);
nand U7190 (N_7190,N_5303,N_4378);
nand U7191 (N_7191,N_5593,N_5553);
or U7192 (N_7192,N_4851,N_4480);
and U7193 (N_7193,N_5764,N_5897);
and U7194 (N_7194,N_5785,N_5210);
nand U7195 (N_7195,N_4088,N_5179);
and U7196 (N_7196,N_4179,N_5716);
or U7197 (N_7197,N_4003,N_4459);
nand U7198 (N_7198,N_5073,N_4294);
nand U7199 (N_7199,N_4179,N_5568);
and U7200 (N_7200,N_5005,N_5655);
or U7201 (N_7201,N_5136,N_5964);
or U7202 (N_7202,N_4947,N_5326);
nor U7203 (N_7203,N_4988,N_4157);
and U7204 (N_7204,N_5494,N_4245);
nor U7205 (N_7205,N_4468,N_5787);
nor U7206 (N_7206,N_5844,N_5460);
or U7207 (N_7207,N_5099,N_4373);
and U7208 (N_7208,N_5088,N_5049);
nor U7209 (N_7209,N_5375,N_4804);
or U7210 (N_7210,N_5719,N_4949);
nand U7211 (N_7211,N_4695,N_4861);
and U7212 (N_7212,N_5441,N_4183);
or U7213 (N_7213,N_4285,N_5316);
or U7214 (N_7214,N_4031,N_5453);
and U7215 (N_7215,N_4017,N_5741);
or U7216 (N_7216,N_4663,N_4113);
and U7217 (N_7217,N_5642,N_5767);
or U7218 (N_7218,N_5389,N_5081);
and U7219 (N_7219,N_4056,N_4425);
nand U7220 (N_7220,N_5139,N_4125);
and U7221 (N_7221,N_5965,N_5791);
xor U7222 (N_7222,N_5873,N_5874);
nand U7223 (N_7223,N_4998,N_4131);
nor U7224 (N_7224,N_4011,N_5269);
or U7225 (N_7225,N_5046,N_5329);
or U7226 (N_7226,N_4950,N_4802);
nand U7227 (N_7227,N_5101,N_5707);
and U7228 (N_7228,N_5078,N_4483);
and U7229 (N_7229,N_4025,N_4963);
nor U7230 (N_7230,N_4973,N_4847);
nand U7231 (N_7231,N_4118,N_5220);
nor U7232 (N_7232,N_4141,N_5414);
nand U7233 (N_7233,N_4950,N_4906);
or U7234 (N_7234,N_5026,N_4171);
nor U7235 (N_7235,N_5769,N_4415);
or U7236 (N_7236,N_5853,N_4570);
or U7237 (N_7237,N_4998,N_4246);
and U7238 (N_7238,N_4506,N_5296);
and U7239 (N_7239,N_5366,N_5239);
nor U7240 (N_7240,N_5585,N_5377);
nor U7241 (N_7241,N_4800,N_4121);
or U7242 (N_7242,N_4719,N_5907);
or U7243 (N_7243,N_5910,N_4317);
nor U7244 (N_7244,N_5749,N_4904);
and U7245 (N_7245,N_5752,N_5749);
or U7246 (N_7246,N_5447,N_4251);
or U7247 (N_7247,N_5403,N_4738);
nand U7248 (N_7248,N_5981,N_5920);
and U7249 (N_7249,N_5136,N_5395);
and U7250 (N_7250,N_5602,N_5449);
nand U7251 (N_7251,N_4457,N_4565);
nand U7252 (N_7252,N_4265,N_4865);
nor U7253 (N_7253,N_5358,N_5129);
nor U7254 (N_7254,N_4753,N_5686);
nand U7255 (N_7255,N_4380,N_5958);
or U7256 (N_7256,N_4593,N_4306);
and U7257 (N_7257,N_4056,N_5734);
or U7258 (N_7258,N_4344,N_5693);
nand U7259 (N_7259,N_4350,N_5650);
or U7260 (N_7260,N_5077,N_4761);
or U7261 (N_7261,N_4203,N_4423);
or U7262 (N_7262,N_5002,N_5223);
and U7263 (N_7263,N_4303,N_4144);
nor U7264 (N_7264,N_5719,N_4989);
nor U7265 (N_7265,N_5890,N_4417);
nand U7266 (N_7266,N_4324,N_4593);
and U7267 (N_7267,N_5061,N_5213);
nand U7268 (N_7268,N_4972,N_4726);
or U7269 (N_7269,N_5474,N_4575);
nor U7270 (N_7270,N_5006,N_4607);
nand U7271 (N_7271,N_4365,N_5515);
nor U7272 (N_7272,N_5204,N_5941);
and U7273 (N_7273,N_4016,N_4335);
nor U7274 (N_7274,N_4857,N_5265);
nand U7275 (N_7275,N_5942,N_5783);
nor U7276 (N_7276,N_5847,N_5884);
and U7277 (N_7277,N_4130,N_5148);
nor U7278 (N_7278,N_5845,N_4142);
xnor U7279 (N_7279,N_5281,N_4805);
nand U7280 (N_7280,N_4808,N_5346);
and U7281 (N_7281,N_4170,N_4639);
nand U7282 (N_7282,N_5646,N_4529);
nand U7283 (N_7283,N_5792,N_4651);
or U7284 (N_7284,N_5803,N_5023);
and U7285 (N_7285,N_5806,N_4579);
nor U7286 (N_7286,N_4570,N_5778);
nor U7287 (N_7287,N_5848,N_4179);
or U7288 (N_7288,N_4399,N_5748);
or U7289 (N_7289,N_5297,N_5740);
xnor U7290 (N_7290,N_5899,N_5368);
or U7291 (N_7291,N_5492,N_5728);
nand U7292 (N_7292,N_4933,N_4002);
and U7293 (N_7293,N_5153,N_4531);
or U7294 (N_7294,N_5792,N_4233);
nand U7295 (N_7295,N_4812,N_4411);
or U7296 (N_7296,N_5972,N_4751);
xnor U7297 (N_7297,N_5581,N_4264);
nor U7298 (N_7298,N_5779,N_4097);
or U7299 (N_7299,N_5909,N_5336);
nor U7300 (N_7300,N_5489,N_4251);
nor U7301 (N_7301,N_4260,N_4655);
nor U7302 (N_7302,N_5141,N_4444);
nor U7303 (N_7303,N_5392,N_5221);
or U7304 (N_7304,N_4061,N_4258);
nand U7305 (N_7305,N_4797,N_5539);
nand U7306 (N_7306,N_4838,N_4298);
and U7307 (N_7307,N_4039,N_4506);
and U7308 (N_7308,N_5896,N_5870);
and U7309 (N_7309,N_5859,N_5801);
nor U7310 (N_7310,N_4939,N_5810);
nand U7311 (N_7311,N_4000,N_4289);
or U7312 (N_7312,N_5738,N_5987);
and U7313 (N_7313,N_4906,N_4012);
nor U7314 (N_7314,N_5102,N_5464);
nor U7315 (N_7315,N_4842,N_4548);
and U7316 (N_7316,N_5091,N_5255);
nand U7317 (N_7317,N_4499,N_4707);
and U7318 (N_7318,N_5555,N_5891);
or U7319 (N_7319,N_4437,N_5226);
and U7320 (N_7320,N_4348,N_4886);
nand U7321 (N_7321,N_4992,N_5128);
and U7322 (N_7322,N_4231,N_5281);
nor U7323 (N_7323,N_5645,N_4338);
and U7324 (N_7324,N_4054,N_4432);
nand U7325 (N_7325,N_4253,N_5254);
nand U7326 (N_7326,N_5654,N_4502);
or U7327 (N_7327,N_5577,N_4872);
nor U7328 (N_7328,N_4430,N_5257);
or U7329 (N_7329,N_5010,N_4152);
or U7330 (N_7330,N_4184,N_5085);
and U7331 (N_7331,N_5365,N_5143);
or U7332 (N_7332,N_5467,N_4636);
nand U7333 (N_7333,N_4056,N_4715);
nor U7334 (N_7334,N_4849,N_5395);
and U7335 (N_7335,N_5779,N_4142);
nand U7336 (N_7336,N_4298,N_4347);
or U7337 (N_7337,N_5675,N_5138);
or U7338 (N_7338,N_4909,N_5151);
nor U7339 (N_7339,N_4539,N_4294);
nand U7340 (N_7340,N_5702,N_4921);
or U7341 (N_7341,N_5874,N_5150);
and U7342 (N_7342,N_5347,N_5948);
and U7343 (N_7343,N_4756,N_4317);
nand U7344 (N_7344,N_4528,N_5486);
and U7345 (N_7345,N_4757,N_5903);
or U7346 (N_7346,N_4628,N_4631);
and U7347 (N_7347,N_5841,N_5777);
and U7348 (N_7348,N_4186,N_4106);
or U7349 (N_7349,N_5544,N_5786);
nor U7350 (N_7350,N_5444,N_5835);
nor U7351 (N_7351,N_5440,N_5516);
nor U7352 (N_7352,N_5973,N_4333);
and U7353 (N_7353,N_4338,N_5911);
or U7354 (N_7354,N_5567,N_5526);
nor U7355 (N_7355,N_5208,N_5642);
nor U7356 (N_7356,N_4738,N_4789);
nand U7357 (N_7357,N_4138,N_5618);
nand U7358 (N_7358,N_5759,N_5407);
nor U7359 (N_7359,N_4078,N_5484);
or U7360 (N_7360,N_5153,N_5303);
and U7361 (N_7361,N_5789,N_5855);
nor U7362 (N_7362,N_5346,N_4816);
nand U7363 (N_7363,N_4366,N_4491);
and U7364 (N_7364,N_5810,N_5583);
and U7365 (N_7365,N_5851,N_5844);
and U7366 (N_7366,N_4538,N_5301);
nand U7367 (N_7367,N_4254,N_5739);
nand U7368 (N_7368,N_4433,N_5282);
or U7369 (N_7369,N_5640,N_4966);
and U7370 (N_7370,N_4483,N_4082);
or U7371 (N_7371,N_5153,N_5248);
nor U7372 (N_7372,N_5844,N_4116);
nor U7373 (N_7373,N_4813,N_4353);
nor U7374 (N_7374,N_5053,N_5832);
or U7375 (N_7375,N_5415,N_5100);
nand U7376 (N_7376,N_4288,N_5106);
nor U7377 (N_7377,N_4715,N_4256);
nand U7378 (N_7378,N_4015,N_5808);
and U7379 (N_7379,N_5572,N_5462);
nor U7380 (N_7380,N_5546,N_4893);
and U7381 (N_7381,N_5163,N_4060);
and U7382 (N_7382,N_4072,N_5630);
nand U7383 (N_7383,N_4439,N_4466);
and U7384 (N_7384,N_5521,N_5826);
nor U7385 (N_7385,N_5142,N_4939);
and U7386 (N_7386,N_4665,N_5842);
nor U7387 (N_7387,N_5031,N_5231);
or U7388 (N_7388,N_4327,N_5461);
and U7389 (N_7389,N_5863,N_5935);
nor U7390 (N_7390,N_4093,N_4709);
nor U7391 (N_7391,N_4462,N_5231);
and U7392 (N_7392,N_4411,N_4078);
or U7393 (N_7393,N_5235,N_4794);
nand U7394 (N_7394,N_5407,N_5669);
and U7395 (N_7395,N_4986,N_4737);
nand U7396 (N_7396,N_4879,N_4235);
nor U7397 (N_7397,N_4251,N_5471);
or U7398 (N_7398,N_5833,N_4019);
nor U7399 (N_7399,N_4883,N_4021);
nor U7400 (N_7400,N_5008,N_5703);
nor U7401 (N_7401,N_5888,N_5979);
and U7402 (N_7402,N_5274,N_4493);
and U7403 (N_7403,N_4779,N_4456);
nand U7404 (N_7404,N_5306,N_5156);
and U7405 (N_7405,N_4459,N_4588);
nor U7406 (N_7406,N_4865,N_4321);
nand U7407 (N_7407,N_4272,N_4488);
or U7408 (N_7408,N_4585,N_5148);
and U7409 (N_7409,N_5659,N_5484);
nor U7410 (N_7410,N_5645,N_5621);
and U7411 (N_7411,N_5313,N_5476);
nand U7412 (N_7412,N_5675,N_5668);
nor U7413 (N_7413,N_5747,N_4834);
nor U7414 (N_7414,N_5605,N_5090);
nand U7415 (N_7415,N_5862,N_5155);
nor U7416 (N_7416,N_4602,N_5835);
nand U7417 (N_7417,N_4032,N_5234);
or U7418 (N_7418,N_5827,N_5616);
nor U7419 (N_7419,N_5519,N_4592);
nand U7420 (N_7420,N_5952,N_4162);
nor U7421 (N_7421,N_5059,N_5589);
nor U7422 (N_7422,N_4961,N_5458);
nand U7423 (N_7423,N_5197,N_4251);
nand U7424 (N_7424,N_4317,N_4106);
nor U7425 (N_7425,N_5547,N_4605);
and U7426 (N_7426,N_5341,N_4432);
or U7427 (N_7427,N_5020,N_4239);
nor U7428 (N_7428,N_5222,N_4843);
nand U7429 (N_7429,N_5257,N_5234);
nor U7430 (N_7430,N_5086,N_5058);
nor U7431 (N_7431,N_4211,N_4506);
and U7432 (N_7432,N_4724,N_5686);
nand U7433 (N_7433,N_5569,N_5612);
nor U7434 (N_7434,N_4885,N_4626);
nand U7435 (N_7435,N_4140,N_4172);
and U7436 (N_7436,N_5146,N_4671);
nor U7437 (N_7437,N_5565,N_4678);
nand U7438 (N_7438,N_5597,N_5896);
nand U7439 (N_7439,N_4121,N_4862);
or U7440 (N_7440,N_4836,N_5786);
or U7441 (N_7441,N_5510,N_5137);
nor U7442 (N_7442,N_4366,N_4853);
nand U7443 (N_7443,N_4030,N_5067);
and U7444 (N_7444,N_4034,N_4536);
and U7445 (N_7445,N_4608,N_5624);
nand U7446 (N_7446,N_5576,N_4967);
nand U7447 (N_7447,N_5604,N_4865);
or U7448 (N_7448,N_4335,N_5232);
nand U7449 (N_7449,N_4825,N_5290);
nand U7450 (N_7450,N_4085,N_4066);
nor U7451 (N_7451,N_5025,N_5276);
and U7452 (N_7452,N_5416,N_4681);
nor U7453 (N_7453,N_4413,N_5717);
or U7454 (N_7454,N_5169,N_5036);
nand U7455 (N_7455,N_5936,N_4675);
and U7456 (N_7456,N_5633,N_4096);
nor U7457 (N_7457,N_4177,N_4608);
and U7458 (N_7458,N_5679,N_4568);
nor U7459 (N_7459,N_5465,N_5728);
or U7460 (N_7460,N_4322,N_4117);
or U7461 (N_7461,N_4473,N_5501);
nor U7462 (N_7462,N_4338,N_4015);
or U7463 (N_7463,N_5085,N_5289);
nand U7464 (N_7464,N_5503,N_4220);
nand U7465 (N_7465,N_4544,N_5606);
nand U7466 (N_7466,N_4525,N_4623);
or U7467 (N_7467,N_4419,N_5738);
nor U7468 (N_7468,N_5924,N_4404);
nor U7469 (N_7469,N_4545,N_4017);
or U7470 (N_7470,N_5463,N_5118);
or U7471 (N_7471,N_5731,N_5627);
or U7472 (N_7472,N_5438,N_5667);
nand U7473 (N_7473,N_5888,N_4856);
xor U7474 (N_7474,N_4464,N_4416);
and U7475 (N_7475,N_4224,N_4653);
or U7476 (N_7476,N_4493,N_5502);
and U7477 (N_7477,N_5608,N_4049);
nor U7478 (N_7478,N_5273,N_5820);
nand U7479 (N_7479,N_4736,N_4953);
and U7480 (N_7480,N_5048,N_4998);
nor U7481 (N_7481,N_5421,N_4200);
and U7482 (N_7482,N_5934,N_5807);
or U7483 (N_7483,N_4653,N_4772);
or U7484 (N_7484,N_4488,N_4342);
nor U7485 (N_7485,N_4231,N_4527);
nor U7486 (N_7486,N_4333,N_5299);
nor U7487 (N_7487,N_4259,N_4215);
or U7488 (N_7488,N_5249,N_5814);
nand U7489 (N_7489,N_5381,N_5299);
nand U7490 (N_7490,N_4640,N_4796);
nand U7491 (N_7491,N_5009,N_4344);
nor U7492 (N_7492,N_4846,N_4403);
and U7493 (N_7493,N_4990,N_4913);
nor U7494 (N_7494,N_5631,N_4814);
nand U7495 (N_7495,N_5406,N_4068);
and U7496 (N_7496,N_5392,N_5329);
and U7497 (N_7497,N_4382,N_5743);
or U7498 (N_7498,N_4082,N_5940);
or U7499 (N_7499,N_4013,N_5625);
nand U7500 (N_7500,N_4185,N_4362);
nor U7501 (N_7501,N_5740,N_5616);
and U7502 (N_7502,N_5646,N_4739);
or U7503 (N_7503,N_4865,N_5531);
nor U7504 (N_7504,N_4918,N_5317);
nor U7505 (N_7505,N_4427,N_5088);
nand U7506 (N_7506,N_4628,N_5211);
and U7507 (N_7507,N_5161,N_4586);
nor U7508 (N_7508,N_5285,N_4652);
nor U7509 (N_7509,N_4351,N_4666);
nor U7510 (N_7510,N_4769,N_4204);
nand U7511 (N_7511,N_4230,N_4855);
nand U7512 (N_7512,N_5368,N_5749);
nor U7513 (N_7513,N_5255,N_4241);
or U7514 (N_7514,N_5221,N_5458);
or U7515 (N_7515,N_4340,N_4023);
nand U7516 (N_7516,N_5134,N_5208);
nand U7517 (N_7517,N_4593,N_5829);
and U7518 (N_7518,N_5121,N_5742);
and U7519 (N_7519,N_4501,N_4933);
or U7520 (N_7520,N_5510,N_4494);
nor U7521 (N_7521,N_5980,N_5360);
nor U7522 (N_7522,N_4718,N_5939);
and U7523 (N_7523,N_5875,N_4196);
or U7524 (N_7524,N_5178,N_4356);
nor U7525 (N_7525,N_5495,N_5855);
and U7526 (N_7526,N_4141,N_5258);
nor U7527 (N_7527,N_5511,N_5287);
or U7528 (N_7528,N_4229,N_5277);
or U7529 (N_7529,N_5398,N_4764);
nor U7530 (N_7530,N_5458,N_4189);
and U7531 (N_7531,N_5943,N_5169);
nor U7532 (N_7532,N_5371,N_4346);
nor U7533 (N_7533,N_5761,N_5583);
nand U7534 (N_7534,N_5210,N_5478);
nor U7535 (N_7535,N_4265,N_4487);
and U7536 (N_7536,N_5497,N_4009);
or U7537 (N_7537,N_4829,N_5313);
nand U7538 (N_7538,N_4328,N_5885);
and U7539 (N_7539,N_5647,N_5475);
nand U7540 (N_7540,N_5943,N_4931);
and U7541 (N_7541,N_4699,N_5272);
nand U7542 (N_7542,N_5842,N_4338);
and U7543 (N_7543,N_5461,N_5818);
nor U7544 (N_7544,N_4010,N_4984);
nand U7545 (N_7545,N_5005,N_4475);
and U7546 (N_7546,N_4431,N_4364);
nor U7547 (N_7547,N_4281,N_4584);
nand U7548 (N_7548,N_4980,N_5227);
or U7549 (N_7549,N_5467,N_5615);
or U7550 (N_7550,N_4237,N_5669);
or U7551 (N_7551,N_5917,N_4057);
nand U7552 (N_7552,N_5392,N_5823);
and U7553 (N_7553,N_5604,N_4143);
and U7554 (N_7554,N_4345,N_5215);
nand U7555 (N_7555,N_4232,N_4153);
or U7556 (N_7556,N_4426,N_4548);
nand U7557 (N_7557,N_4387,N_5332);
or U7558 (N_7558,N_5922,N_4765);
and U7559 (N_7559,N_5490,N_5342);
and U7560 (N_7560,N_5191,N_5073);
nor U7561 (N_7561,N_4512,N_5026);
or U7562 (N_7562,N_5109,N_4793);
nor U7563 (N_7563,N_4422,N_5406);
nand U7564 (N_7564,N_4944,N_4671);
nor U7565 (N_7565,N_4517,N_5548);
nor U7566 (N_7566,N_4971,N_5570);
and U7567 (N_7567,N_4798,N_4456);
and U7568 (N_7568,N_5798,N_4050);
nor U7569 (N_7569,N_4224,N_5892);
nor U7570 (N_7570,N_5085,N_5309);
and U7571 (N_7571,N_4763,N_5841);
nor U7572 (N_7572,N_4128,N_5312);
and U7573 (N_7573,N_5967,N_4642);
nor U7574 (N_7574,N_4697,N_4492);
nand U7575 (N_7575,N_4729,N_5887);
nor U7576 (N_7576,N_5952,N_5090);
and U7577 (N_7577,N_5272,N_5599);
and U7578 (N_7578,N_5535,N_4449);
and U7579 (N_7579,N_4532,N_5293);
or U7580 (N_7580,N_4270,N_5247);
or U7581 (N_7581,N_5698,N_5481);
nor U7582 (N_7582,N_5938,N_4312);
nand U7583 (N_7583,N_4745,N_5639);
xor U7584 (N_7584,N_5440,N_5897);
or U7585 (N_7585,N_5594,N_5218);
nand U7586 (N_7586,N_5753,N_4124);
or U7587 (N_7587,N_5031,N_5466);
and U7588 (N_7588,N_5397,N_4019);
and U7589 (N_7589,N_5517,N_4621);
and U7590 (N_7590,N_4247,N_4486);
nor U7591 (N_7591,N_4357,N_5087);
nand U7592 (N_7592,N_5074,N_4636);
nor U7593 (N_7593,N_5000,N_4327);
or U7594 (N_7594,N_4492,N_4195);
nor U7595 (N_7595,N_4323,N_5603);
or U7596 (N_7596,N_4538,N_4349);
or U7597 (N_7597,N_4312,N_5736);
nor U7598 (N_7598,N_5081,N_5714);
nor U7599 (N_7599,N_5201,N_5146);
and U7600 (N_7600,N_4654,N_4116);
nand U7601 (N_7601,N_5991,N_5697);
nor U7602 (N_7602,N_5629,N_5478);
nor U7603 (N_7603,N_4856,N_4601);
or U7604 (N_7604,N_4954,N_4734);
or U7605 (N_7605,N_5189,N_4032);
nand U7606 (N_7606,N_5403,N_5002);
or U7607 (N_7607,N_5832,N_5730);
nand U7608 (N_7608,N_5227,N_4292);
nand U7609 (N_7609,N_5803,N_4555);
xnor U7610 (N_7610,N_5235,N_5620);
or U7611 (N_7611,N_4116,N_4133);
nor U7612 (N_7612,N_4624,N_5088);
nand U7613 (N_7613,N_5777,N_5509);
nor U7614 (N_7614,N_5938,N_4611);
or U7615 (N_7615,N_4765,N_4997);
nand U7616 (N_7616,N_4556,N_5412);
and U7617 (N_7617,N_4274,N_5358);
or U7618 (N_7618,N_4615,N_5789);
or U7619 (N_7619,N_5202,N_5873);
and U7620 (N_7620,N_4643,N_4725);
nand U7621 (N_7621,N_4406,N_4668);
or U7622 (N_7622,N_5827,N_5581);
nand U7623 (N_7623,N_4373,N_5407);
nand U7624 (N_7624,N_4471,N_4184);
nand U7625 (N_7625,N_4404,N_4065);
or U7626 (N_7626,N_4559,N_4755);
and U7627 (N_7627,N_5761,N_5819);
nor U7628 (N_7628,N_5181,N_5499);
xnor U7629 (N_7629,N_5289,N_4877);
nand U7630 (N_7630,N_5679,N_4147);
and U7631 (N_7631,N_5049,N_5061);
nand U7632 (N_7632,N_5023,N_5794);
or U7633 (N_7633,N_5399,N_5454);
and U7634 (N_7634,N_5938,N_5076);
nor U7635 (N_7635,N_5931,N_4332);
nor U7636 (N_7636,N_4339,N_4292);
xor U7637 (N_7637,N_4669,N_4769);
nor U7638 (N_7638,N_5196,N_4646);
and U7639 (N_7639,N_5489,N_5957);
nand U7640 (N_7640,N_4161,N_4071);
and U7641 (N_7641,N_5960,N_4373);
nor U7642 (N_7642,N_5877,N_5097);
or U7643 (N_7643,N_5116,N_4215);
nor U7644 (N_7644,N_4096,N_4000);
nand U7645 (N_7645,N_5627,N_5186);
nand U7646 (N_7646,N_5288,N_4248);
nand U7647 (N_7647,N_4834,N_4673);
nand U7648 (N_7648,N_5705,N_4826);
and U7649 (N_7649,N_4672,N_4381);
nor U7650 (N_7650,N_4065,N_4277);
nand U7651 (N_7651,N_5806,N_5900);
nand U7652 (N_7652,N_5224,N_5874);
or U7653 (N_7653,N_4638,N_4497);
and U7654 (N_7654,N_4840,N_4528);
nor U7655 (N_7655,N_5784,N_4970);
nor U7656 (N_7656,N_4658,N_4307);
or U7657 (N_7657,N_5873,N_5259);
or U7658 (N_7658,N_5379,N_5000);
or U7659 (N_7659,N_4506,N_4437);
nand U7660 (N_7660,N_4531,N_5026);
or U7661 (N_7661,N_4146,N_4465);
nor U7662 (N_7662,N_5202,N_5749);
nor U7663 (N_7663,N_5310,N_5697);
and U7664 (N_7664,N_5101,N_4320);
nand U7665 (N_7665,N_4180,N_5263);
nand U7666 (N_7666,N_4090,N_4923);
and U7667 (N_7667,N_5043,N_5883);
and U7668 (N_7668,N_5532,N_4453);
or U7669 (N_7669,N_5408,N_4083);
or U7670 (N_7670,N_5909,N_5254);
nor U7671 (N_7671,N_5522,N_4738);
and U7672 (N_7672,N_5838,N_4843);
nand U7673 (N_7673,N_4330,N_4553);
nor U7674 (N_7674,N_4714,N_4914);
nor U7675 (N_7675,N_5009,N_4898);
xor U7676 (N_7676,N_4367,N_5077);
nor U7677 (N_7677,N_5852,N_5176);
nand U7678 (N_7678,N_4553,N_4905);
nor U7679 (N_7679,N_4795,N_5362);
and U7680 (N_7680,N_5895,N_5966);
nand U7681 (N_7681,N_5279,N_4650);
and U7682 (N_7682,N_5713,N_4662);
nor U7683 (N_7683,N_5873,N_4720);
and U7684 (N_7684,N_4894,N_4520);
nand U7685 (N_7685,N_5233,N_5948);
nand U7686 (N_7686,N_5629,N_5624);
nand U7687 (N_7687,N_5758,N_4124);
nor U7688 (N_7688,N_5224,N_5369);
or U7689 (N_7689,N_5557,N_4921);
nor U7690 (N_7690,N_5589,N_4594);
nand U7691 (N_7691,N_5598,N_5387);
or U7692 (N_7692,N_5051,N_4670);
and U7693 (N_7693,N_4330,N_4246);
nor U7694 (N_7694,N_4817,N_5037);
and U7695 (N_7695,N_4061,N_4979);
nand U7696 (N_7696,N_5763,N_4724);
and U7697 (N_7697,N_5560,N_5569);
nor U7698 (N_7698,N_4908,N_5698);
and U7699 (N_7699,N_4127,N_4206);
and U7700 (N_7700,N_5896,N_4403);
or U7701 (N_7701,N_5721,N_4545);
and U7702 (N_7702,N_5910,N_5046);
nand U7703 (N_7703,N_4799,N_5611);
and U7704 (N_7704,N_4514,N_4293);
nor U7705 (N_7705,N_5853,N_5052);
and U7706 (N_7706,N_5591,N_4885);
and U7707 (N_7707,N_5616,N_4593);
or U7708 (N_7708,N_4429,N_4606);
nor U7709 (N_7709,N_4125,N_4097);
nor U7710 (N_7710,N_5833,N_5111);
nand U7711 (N_7711,N_5363,N_4982);
nor U7712 (N_7712,N_4133,N_4331);
or U7713 (N_7713,N_4859,N_4222);
or U7714 (N_7714,N_5873,N_5025);
nand U7715 (N_7715,N_5741,N_4553);
or U7716 (N_7716,N_5284,N_5810);
nand U7717 (N_7717,N_5391,N_5250);
and U7718 (N_7718,N_4444,N_5713);
or U7719 (N_7719,N_4503,N_4440);
nand U7720 (N_7720,N_5985,N_5727);
and U7721 (N_7721,N_5634,N_5666);
nand U7722 (N_7722,N_4228,N_5700);
or U7723 (N_7723,N_4969,N_5297);
nor U7724 (N_7724,N_4723,N_4824);
and U7725 (N_7725,N_4472,N_4408);
or U7726 (N_7726,N_4307,N_4278);
and U7727 (N_7727,N_4095,N_5129);
nand U7728 (N_7728,N_5075,N_4528);
nand U7729 (N_7729,N_5623,N_4522);
and U7730 (N_7730,N_4960,N_5992);
nand U7731 (N_7731,N_5979,N_4926);
nor U7732 (N_7732,N_4022,N_5055);
nor U7733 (N_7733,N_4272,N_5809);
nor U7734 (N_7734,N_4049,N_5921);
or U7735 (N_7735,N_4635,N_4219);
and U7736 (N_7736,N_5870,N_4185);
and U7737 (N_7737,N_4447,N_5772);
and U7738 (N_7738,N_4814,N_5920);
and U7739 (N_7739,N_5491,N_5223);
nor U7740 (N_7740,N_4632,N_5966);
nor U7741 (N_7741,N_4998,N_5137);
and U7742 (N_7742,N_4499,N_5631);
or U7743 (N_7743,N_5773,N_5643);
and U7744 (N_7744,N_4712,N_4077);
and U7745 (N_7745,N_5580,N_5748);
and U7746 (N_7746,N_5251,N_5428);
and U7747 (N_7747,N_4565,N_4791);
nor U7748 (N_7748,N_5407,N_4399);
or U7749 (N_7749,N_4254,N_5393);
nand U7750 (N_7750,N_4381,N_4133);
or U7751 (N_7751,N_4650,N_5702);
or U7752 (N_7752,N_4297,N_5782);
and U7753 (N_7753,N_5458,N_4540);
or U7754 (N_7754,N_4604,N_5383);
nand U7755 (N_7755,N_5625,N_5679);
or U7756 (N_7756,N_4828,N_4478);
and U7757 (N_7757,N_4039,N_5298);
nand U7758 (N_7758,N_4947,N_5737);
and U7759 (N_7759,N_5602,N_4006);
nand U7760 (N_7760,N_5615,N_4257);
or U7761 (N_7761,N_5049,N_4873);
nand U7762 (N_7762,N_4374,N_4761);
nand U7763 (N_7763,N_5024,N_5651);
and U7764 (N_7764,N_4357,N_5155);
nand U7765 (N_7765,N_5076,N_5550);
nand U7766 (N_7766,N_5920,N_5322);
and U7767 (N_7767,N_5337,N_5414);
nor U7768 (N_7768,N_5591,N_4084);
or U7769 (N_7769,N_5168,N_4783);
and U7770 (N_7770,N_5595,N_4872);
nand U7771 (N_7771,N_5736,N_5050);
nand U7772 (N_7772,N_5736,N_5126);
or U7773 (N_7773,N_5050,N_4264);
or U7774 (N_7774,N_4164,N_4252);
nor U7775 (N_7775,N_5884,N_5715);
or U7776 (N_7776,N_5191,N_4660);
nand U7777 (N_7777,N_5311,N_5504);
nand U7778 (N_7778,N_4822,N_5911);
and U7779 (N_7779,N_4277,N_4517);
and U7780 (N_7780,N_4248,N_5761);
or U7781 (N_7781,N_5845,N_5857);
and U7782 (N_7782,N_5848,N_4327);
nor U7783 (N_7783,N_5146,N_5883);
nor U7784 (N_7784,N_4358,N_4002);
nor U7785 (N_7785,N_5847,N_5408);
nand U7786 (N_7786,N_4972,N_4192);
nor U7787 (N_7787,N_5543,N_5015);
nand U7788 (N_7788,N_5593,N_5566);
and U7789 (N_7789,N_4432,N_5372);
nor U7790 (N_7790,N_5216,N_4415);
or U7791 (N_7791,N_5386,N_5339);
or U7792 (N_7792,N_5477,N_4913);
or U7793 (N_7793,N_5517,N_4398);
or U7794 (N_7794,N_4259,N_5198);
nand U7795 (N_7795,N_5874,N_4781);
and U7796 (N_7796,N_4847,N_4509);
nor U7797 (N_7797,N_5539,N_4428);
nand U7798 (N_7798,N_5232,N_4928);
or U7799 (N_7799,N_5541,N_5343);
nor U7800 (N_7800,N_5769,N_5891);
and U7801 (N_7801,N_5586,N_5549);
nor U7802 (N_7802,N_4597,N_4645);
or U7803 (N_7803,N_4772,N_5153);
nand U7804 (N_7804,N_5460,N_4104);
nand U7805 (N_7805,N_5927,N_5913);
nand U7806 (N_7806,N_5763,N_4154);
or U7807 (N_7807,N_5553,N_4539);
and U7808 (N_7808,N_4266,N_4549);
nand U7809 (N_7809,N_5804,N_4623);
or U7810 (N_7810,N_4213,N_4795);
nand U7811 (N_7811,N_4353,N_5721);
and U7812 (N_7812,N_5278,N_4252);
nor U7813 (N_7813,N_5977,N_4472);
and U7814 (N_7814,N_4750,N_4831);
or U7815 (N_7815,N_5641,N_4278);
nor U7816 (N_7816,N_4717,N_4111);
nand U7817 (N_7817,N_4060,N_4183);
xor U7818 (N_7818,N_4648,N_5567);
nor U7819 (N_7819,N_4283,N_4774);
or U7820 (N_7820,N_4165,N_4765);
and U7821 (N_7821,N_4803,N_5212);
or U7822 (N_7822,N_4546,N_4915);
nor U7823 (N_7823,N_5224,N_5935);
nor U7824 (N_7824,N_5348,N_4180);
and U7825 (N_7825,N_5868,N_5926);
or U7826 (N_7826,N_4964,N_5596);
nor U7827 (N_7827,N_5510,N_4180);
nand U7828 (N_7828,N_5882,N_5699);
nand U7829 (N_7829,N_4902,N_4883);
nand U7830 (N_7830,N_5815,N_4465);
and U7831 (N_7831,N_4751,N_5950);
nor U7832 (N_7832,N_4690,N_4410);
or U7833 (N_7833,N_5007,N_4598);
and U7834 (N_7834,N_4899,N_5771);
or U7835 (N_7835,N_5390,N_5124);
nand U7836 (N_7836,N_4632,N_4884);
and U7837 (N_7837,N_5853,N_5445);
nor U7838 (N_7838,N_4666,N_5814);
or U7839 (N_7839,N_5434,N_4833);
nor U7840 (N_7840,N_4599,N_5629);
or U7841 (N_7841,N_5654,N_5747);
and U7842 (N_7842,N_4363,N_4885);
and U7843 (N_7843,N_5605,N_4344);
nand U7844 (N_7844,N_5281,N_5165);
and U7845 (N_7845,N_4367,N_4507);
and U7846 (N_7846,N_4876,N_5691);
nor U7847 (N_7847,N_5044,N_5705);
and U7848 (N_7848,N_4470,N_4569);
or U7849 (N_7849,N_4070,N_5755);
nand U7850 (N_7850,N_5863,N_4699);
nor U7851 (N_7851,N_4457,N_4141);
and U7852 (N_7852,N_4515,N_5808);
nor U7853 (N_7853,N_4544,N_5880);
and U7854 (N_7854,N_4071,N_4255);
xnor U7855 (N_7855,N_5350,N_4177);
nand U7856 (N_7856,N_5426,N_4312);
nand U7857 (N_7857,N_5007,N_4272);
nor U7858 (N_7858,N_5841,N_5336);
nand U7859 (N_7859,N_4734,N_5100);
nor U7860 (N_7860,N_4292,N_5157);
or U7861 (N_7861,N_4983,N_4317);
and U7862 (N_7862,N_5907,N_5781);
or U7863 (N_7863,N_5339,N_4242);
nand U7864 (N_7864,N_5019,N_4187);
nor U7865 (N_7865,N_5141,N_5839);
nand U7866 (N_7866,N_5292,N_5041);
nor U7867 (N_7867,N_5881,N_5872);
and U7868 (N_7868,N_4129,N_4652);
and U7869 (N_7869,N_4975,N_4878);
and U7870 (N_7870,N_4006,N_4633);
nor U7871 (N_7871,N_5878,N_5709);
or U7872 (N_7872,N_4569,N_5423);
or U7873 (N_7873,N_5471,N_5437);
nand U7874 (N_7874,N_5430,N_5429);
nor U7875 (N_7875,N_4018,N_5984);
nand U7876 (N_7876,N_4662,N_5616);
or U7877 (N_7877,N_5332,N_5901);
nand U7878 (N_7878,N_4731,N_4276);
or U7879 (N_7879,N_5843,N_5903);
nor U7880 (N_7880,N_5175,N_4011);
nand U7881 (N_7881,N_4740,N_5682);
nand U7882 (N_7882,N_5662,N_5515);
nor U7883 (N_7883,N_5005,N_4799);
nand U7884 (N_7884,N_5413,N_4535);
or U7885 (N_7885,N_4747,N_5616);
or U7886 (N_7886,N_5843,N_4477);
nand U7887 (N_7887,N_5479,N_5351);
and U7888 (N_7888,N_5973,N_5447);
and U7889 (N_7889,N_4315,N_5083);
nand U7890 (N_7890,N_4345,N_4056);
or U7891 (N_7891,N_5363,N_5081);
or U7892 (N_7892,N_5723,N_4884);
nand U7893 (N_7893,N_5960,N_5217);
and U7894 (N_7894,N_5482,N_4184);
nor U7895 (N_7895,N_4170,N_5059);
or U7896 (N_7896,N_5955,N_5187);
nor U7897 (N_7897,N_4826,N_4346);
or U7898 (N_7898,N_5455,N_5308);
or U7899 (N_7899,N_4674,N_4935);
nor U7900 (N_7900,N_5006,N_5278);
and U7901 (N_7901,N_5403,N_4514);
nor U7902 (N_7902,N_4423,N_5517);
or U7903 (N_7903,N_4296,N_4506);
or U7904 (N_7904,N_5063,N_4387);
nor U7905 (N_7905,N_4106,N_5230);
and U7906 (N_7906,N_4050,N_5394);
or U7907 (N_7907,N_5932,N_5547);
nor U7908 (N_7908,N_5842,N_5073);
nor U7909 (N_7909,N_5948,N_5293);
or U7910 (N_7910,N_4430,N_5756);
nand U7911 (N_7911,N_5478,N_5746);
and U7912 (N_7912,N_5972,N_4061);
nand U7913 (N_7913,N_4778,N_5500);
and U7914 (N_7914,N_4337,N_4971);
or U7915 (N_7915,N_4821,N_4129);
nor U7916 (N_7916,N_4216,N_5706);
and U7917 (N_7917,N_5035,N_4393);
nand U7918 (N_7918,N_4471,N_5794);
nor U7919 (N_7919,N_4937,N_5592);
nand U7920 (N_7920,N_5627,N_4283);
nand U7921 (N_7921,N_4324,N_4584);
nor U7922 (N_7922,N_4736,N_5652);
nor U7923 (N_7923,N_5736,N_5714);
nor U7924 (N_7924,N_4444,N_4597);
and U7925 (N_7925,N_4570,N_4470);
and U7926 (N_7926,N_4093,N_4133);
or U7927 (N_7927,N_4484,N_5912);
or U7928 (N_7928,N_4954,N_4665);
nand U7929 (N_7929,N_4671,N_5604);
nor U7930 (N_7930,N_4228,N_4827);
nor U7931 (N_7931,N_4645,N_5218);
and U7932 (N_7932,N_4939,N_4588);
nand U7933 (N_7933,N_4193,N_5997);
or U7934 (N_7934,N_4902,N_4891);
nor U7935 (N_7935,N_4417,N_5667);
nor U7936 (N_7936,N_5885,N_5754);
and U7937 (N_7937,N_5102,N_4617);
nor U7938 (N_7938,N_4687,N_5723);
and U7939 (N_7939,N_5910,N_5590);
and U7940 (N_7940,N_5489,N_5288);
nand U7941 (N_7941,N_4669,N_5545);
nand U7942 (N_7942,N_5800,N_5275);
or U7943 (N_7943,N_5010,N_4038);
and U7944 (N_7944,N_4764,N_5518);
and U7945 (N_7945,N_4429,N_5948);
nor U7946 (N_7946,N_5791,N_4348);
nand U7947 (N_7947,N_5637,N_5159);
or U7948 (N_7948,N_4080,N_4657);
nand U7949 (N_7949,N_4193,N_4200);
or U7950 (N_7950,N_5456,N_4963);
or U7951 (N_7951,N_5281,N_5405);
nor U7952 (N_7952,N_5261,N_4000);
and U7953 (N_7953,N_4595,N_5361);
or U7954 (N_7954,N_5407,N_4305);
and U7955 (N_7955,N_5137,N_5568);
nor U7956 (N_7956,N_4594,N_5142);
nand U7957 (N_7957,N_4294,N_4673);
and U7958 (N_7958,N_5216,N_4528);
nor U7959 (N_7959,N_4282,N_4833);
or U7960 (N_7960,N_5973,N_4771);
xnor U7961 (N_7961,N_4610,N_5782);
or U7962 (N_7962,N_4011,N_4652);
nand U7963 (N_7963,N_5932,N_5412);
nor U7964 (N_7964,N_5321,N_4262);
nand U7965 (N_7965,N_4539,N_5945);
or U7966 (N_7966,N_4816,N_4138);
nand U7967 (N_7967,N_5065,N_4609);
and U7968 (N_7968,N_5847,N_5962);
nand U7969 (N_7969,N_5433,N_5628);
and U7970 (N_7970,N_5417,N_5937);
and U7971 (N_7971,N_4502,N_5512);
or U7972 (N_7972,N_4251,N_5826);
and U7973 (N_7973,N_4438,N_5891);
or U7974 (N_7974,N_5286,N_4457);
xor U7975 (N_7975,N_4128,N_5023);
nand U7976 (N_7976,N_4888,N_5403);
and U7977 (N_7977,N_4945,N_5682);
nand U7978 (N_7978,N_4147,N_4028);
and U7979 (N_7979,N_4053,N_5408);
xnor U7980 (N_7980,N_5279,N_4468);
or U7981 (N_7981,N_4498,N_4589);
and U7982 (N_7982,N_5285,N_5030);
nor U7983 (N_7983,N_5104,N_4426);
or U7984 (N_7984,N_4819,N_5555);
nand U7985 (N_7985,N_5622,N_4630);
nor U7986 (N_7986,N_4351,N_5851);
xnor U7987 (N_7987,N_5938,N_4068);
and U7988 (N_7988,N_4364,N_4946);
nor U7989 (N_7989,N_5679,N_4840);
and U7990 (N_7990,N_4086,N_4844);
nand U7991 (N_7991,N_5264,N_5901);
or U7992 (N_7992,N_5106,N_4799);
nor U7993 (N_7993,N_4852,N_5649);
or U7994 (N_7994,N_5879,N_5244);
and U7995 (N_7995,N_5708,N_4966);
nor U7996 (N_7996,N_4426,N_5060);
nand U7997 (N_7997,N_4316,N_5554);
nand U7998 (N_7998,N_4729,N_5302);
nand U7999 (N_7999,N_5491,N_4551);
nand U8000 (N_8000,N_6437,N_6157);
xor U8001 (N_8001,N_7890,N_7784);
nor U8002 (N_8002,N_6961,N_6251);
or U8003 (N_8003,N_6143,N_7945);
nand U8004 (N_8004,N_7187,N_6534);
and U8005 (N_8005,N_6795,N_7330);
and U8006 (N_8006,N_7824,N_7834);
nand U8007 (N_8007,N_7078,N_7052);
nand U8008 (N_8008,N_7669,N_6692);
and U8009 (N_8009,N_6225,N_6531);
nor U8010 (N_8010,N_7105,N_7268);
and U8011 (N_8011,N_7030,N_6834);
or U8012 (N_8012,N_7478,N_7167);
nor U8013 (N_8013,N_6425,N_7323);
nor U8014 (N_8014,N_7120,N_6129);
or U8015 (N_8015,N_6957,N_6621);
and U8016 (N_8016,N_7798,N_7009);
nor U8017 (N_8017,N_7370,N_6981);
or U8018 (N_8018,N_6641,N_7579);
nor U8019 (N_8019,N_7433,N_7211);
nand U8020 (N_8020,N_7244,N_6956);
and U8021 (N_8021,N_6459,N_6852);
and U8022 (N_8022,N_7879,N_7832);
and U8023 (N_8023,N_6636,N_6421);
nor U8024 (N_8024,N_6653,N_7852);
and U8025 (N_8025,N_7547,N_6120);
or U8026 (N_8026,N_6031,N_6438);
and U8027 (N_8027,N_7253,N_7762);
nand U8028 (N_8028,N_6618,N_6883);
nor U8029 (N_8029,N_7988,N_7247);
and U8030 (N_8030,N_7873,N_7492);
or U8031 (N_8031,N_7977,N_6044);
and U8032 (N_8032,N_7667,N_7168);
or U8033 (N_8033,N_6070,N_6314);
nand U8034 (N_8034,N_6212,N_6187);
and U8035 (N_8035,N_7942,N_6182);
and U8036 (N_8036,N_7399,N_7975);
nand U8037 (N_8037,N_6165,N_7348);
or U8038 (N_8038,N_7276,N_6483);
and U8039 (N_8039,N_7032,N_7599);
nand U8040 (N_8040,N_7170,N_7146);
and U8041 (N_8041,N_6985,N_7055);
and U8042 (N_8042,N_6853,N_7109);
and U8043 (N_8043,N_7713,N_6922);
or U8044 (N_8044,N_7930,N_6480);
nand U8045 (N_8045,N_7169,N_6519);
nor U8046 (N_8046,N_7031,N_6958);
nor U8047 (N_8047,N_7489,N_7225);
or U8048 (N_8048,N_6064,N_7519);
nor U8049 (N_8049,N_7668,N_7865);
nor U8050 (N_8050,N_7722,N_6654);
or U8051 (N_8051,N_6757,N_6499);
nor U8052 (N_8052,N_7926,N_7967);
nand U8053 (N_8053,N_6803,N_6105);
or U8054 (N_8054,N_7582,N_7110);
or U8055 (N_8055,N_6797,N_6918);
nand U8056 (N_8056,N_6805,N_6727);
or U8057 (N_8057,N_6171,N_6110);
and U8058 (N_8058,N_7261,N_7228);
nand U8059 (N_8059,N_7015,N_6948);
or U8060 (N_8060,N_6392,N_6050);
nor U8061 (N_8061,N_7158,N_6703);
nor U8062 (N_8062,N_6931,N_7781);
or U8063 (N_8063,N_6744,N_7178);
or U8064 (N_8064,N_6460,N_6203);
nor U8065 (N_8065,N_7946,N_6310);
and U8066 (N_8066,N_7269,N_6486);
nor U8067 (N_8067,N_7773,N_6631);
nand U8068 (N_8068,N_6742,N_6923);
and U8069 (N_8069,N_7687,N_6462);
nor U8070 (N_8070,N_6321,N_6357);
nor U8071 (N_8071,N_7822,N_6983);
and U8072 (N_8072,N_6214,N_6092);
or U8073 (N_8073,N_6262,N_6788);
or U8074 (N_8074,N_7462,N_6144);
nand U8075 (N_8075,N_7398,N_6525);
nand U8076 (N_8076,N_6152,N_7311);
and U8077 (N_8077,N_6794,N_6134);
or U8078 (N_8078,N_7750,N_6101);
nand U8079 (N_8079,N_7285,N_6432);
and U8080 (N_8080,N_6532,N_6719);
nor U8081 (N_8081,N_6585,N_6518);
nand U8082 (N_8082,N_6612,N_6146);
and U8083 (N_8083,N_7486,N_7809);
or U8084 (N_8084,N_7072,N_6232);
and U8085 (N_8085,N_6884,N_6975);
nor U8086 (N_8086,N_7223,N_6691);
or U8087 (N_8087,N_7801,N_7556);
nor U8088 (N_8088,N_7024,N_6091);
nor U8089 (N_8089,N_6205,N_6500);
nor U8090 (N_8090,N_7441,N_6294);
and U8091 (N_8091,N_7617,N_7405);
nand U8092 (N_8092,N_7037,N_6575);
or U8093 (N_8093,N_7724,N_7088);
and U8094 (N_8094,N_6115,N_7363);
or U8095 (N_8095,N_6769,N_7473);
nand U8096 (N_8096,N_6013,N_7565);
or U8097 (N_8097,N_6693,N_6060);
nor U8098 (N_8098,N_7603,N_7998);
and U8099 (N_8099,N_7983,N_6163);
nand U8100 (N_8100,N_7344,N_6337);
nand U8101 (N_8101,N_7665,N_6919);
nor U8102 (N_8102,N_6124,N_7346);
and U8103 (N_8103,N_6995,N_7915);
and U8104 (N_8104,N_6536,N_6130);
nand U8105 (N_8105,N_6153,N_7954);
nand U8106 (N_8106,N_7432,N_7270);
nand U8107 (N_8107,N_6002,N_7723);
and U8108 (N_8108,N_7540,N_7897);
and U8109 (N_8109,N_7561,N_7118);
nor U8110 (N_8110,N_6449,N_6676);
nor U8111 (N_8111,N_6396,N_6655);
nand U8112 (N_8112,N_7697,N_7746);
and U8113 (N_8113,N_6916,N_6327);
or U8114 (N_8114,N_7522,N_6541);
nor U8115 (N_8115,N_7586,N_7705);
nand U8116 (N_8116,N_6285,N_7510);
and U8117 (N_8117,N_7604,N_7876);
nand U8118 (N_8118,N_7925,N_6039);
nor U8119 (N_8119,N_7352,N_7690);
nand U8120 (N_8120,N_7191,N_6810);
and U8121 (N_8121,N_7036,N_6213);
nor U8122 (N_8122,N_7658,N_7921);
nand U8123 (N_8123,N_7494,N_7259);
nand U8124 (N_8124,N_7151,N_7091);
or U8125 (N_8125,N_6936,N_7403);
nand U8126 (N_8126,N_6180,N_6228);
and U8127 (N_8127,N_6823,N_6850);
xnor U8128 (N_8128,N_6287,N_6420);
or U8129 (N_8129,N_7631,N_6920);
and U8130 (N_8130,N_7855,N_7257);
or U8131 (N_8131,N_7601,N_6414);
or U8132 (N_8132,N_7161,N_6109);
nand U8133 (N_8133,N_7434,N_6424);
nand U8134 (N_8134,N_6763,N_6315);
nand U8135 (N_8135,N_7585,N_6629);
or U8136 (N_8136,N_6193,N_7020);
and U8137 (N_8137,N_7445,N_6955);
and U8138 (N_8138,N_7831,N_6147);
nor U8139 (N_8139,N_6684,N_7240);
or U8140 (N_8140,N_7867,N_6019);
nor U8141 (N_8141,N_6498,N_7797);
nand U8142 (N_8142,N_7113,N_6061);
nand U8143 (N_8143,N_7108,N_6054);
nor U8144 (N_8144,N_6409,N_6749);
and U8145 (N_8145,N_6448,N_6024);
and U8146 (N_8146,N_6501,N_7356);
nand U8147 (N_8147,N_6735,N_6240);
or U8148 (N_8148,N_6813,N_6700);
nor U8149 (N_8149,N_6762,N_6201);
nor U8150 (N_8150,N_7458,N_6894);
nor U8151 (N_8151,N_6177,N_6487);
or U8152 (N_8152,N_6907,N_7783);
nor U8153 (N_8153,N_6301,N_7207);
nand U8154 (N_8154,N_7581,N_7281);
or U8155 (N_8155,N_7325,N_7029);
and U8156 (N_8156,N_6765,N_7304);
or U8157 (N_8157,N_6974,N_6550);
and U8158 (N_8158,N_6325,N_6069);
or U8159 (N_8159,N_6309,N_7294);
nor U8160 (N_8160,N_7924,N_7107);
nand U8161 (N_8161,N_6045,N_7224);
nor U8162 (N_8162,N_7734,N_7076);
and U8163 (N_8163,N_7136,N_7466);
nand U8164 (N_8164,N_6634,N_6710);
and U8165 (N_8165,N_7950,N_7550);
and U8166 (N_8166,N_7386,N_6476);
nand U8167 (N_8167,N_6156,N_7771);
nand U8168 (N_8168,N_6914,N_7079);
nor U8169 (N_8169,N_6740,N_7551);
nor U8170 (N_8170,N_6485,N_7789);
or U8171 (N_8171,N_6046,N_6543);
and U8172 (N_8172,N_7452,N_6601);
or U8173 (N_8173,N_6697,N_6319);
nand U8174 (N_8174,N_6578,N_7912);
and U8175 (N_8175,N_7607,N_7575);
nand U8176 (N_8176,N_7058,N_6878);
nor U8177 (N_8177,N_7811,N_6018);
nand U8178 (N_8178,N_7471,N_7866);
and U8179 (N_8179,N_6354,N_7064);
and U8180 (N_8180,N_6638,N_6389);
nor U8181 (N_8181,N_7589,N_6554);
or U8182 (N_8182,N_6677,N_7212);
nand U8183 (N_8183,N_7678,N_6650);
nor U8184 (N_8184,N_7391,N_7358);
or U8185 (N_8185,N_7558,N_7780);
or U8186 (N_8186,N_7903,N_6741);
nor U8187 (N_8187,N_7862,N_6622);
nand U8188 (N_8188,N_7812,N_7731);
nor U8189 (N_8189,N_7173,N_6768);
nor U8190 (N_8190,N_6737,N_6510);
and U8191 (N_8191,N_7184,N_6912);
nor U8192 (N_8192,N_6140,N_6828);
or U8193 (N_8193,N_7028,N_6348);
nor U8194 (N_8194,N_6899,N_6860);
nand U8195 (N_8195,N_7958,N_7735);
and U8196 (N_8196,N_7769,N_7442);
nand U8197 (N_8197,N_6461,N_7626);
or U8198 (N_8198,N_7150,N_7680);
nand U8199 (N_8199,N_7538,N_7898);
nor U8200 (N_8200,N_6395,N_7414);
or U8201 (N_8201,N_6572,N_7996);
and U8202 (N_8202,N_6080,N_7083);
xor U8203 (N_8203,N_7310,N_7010);
and U8204 (N_8204,N_6305,N_7905);
nor U8205 (N_8205,N_7467,N_7190);
and U8206 (N_8206,N_7858,N_6141);
or U8207 (N_8207,N_6784,N_7124);
nor U8208 (N_8208,N_6355,N_6626);
nand U8209 (N_8209,N_6349,N_7104);
nor U8210 (N_8210,N_6248,N_6452);
nor U8211 (N_8211,N_7049,N_6383);
or U8212 (N_8212,N_7001,N_6973);
nor U8213 (N_8213,N_6652,N_6867);
nor U8214 (N_8214,N_6398,N_7699);
nand U8215 (N_8215,N_7666,N_6244);
and U8216 (N_8216,N_7464,N_7045);
nand U8217 (N_8217,N_7047,N_6154);
and U8218 (N_8218,N_6508,N_7140);
nor U8219 (N_8219,N_6989,N_6352);
xor U8220 (N_8220,N_7643,N_7900);
and U8221 (N_8221,N_7937,N_6714);
or U8222 (N_8222,N_7417,N_6647);
or U8223 (N_8223,N_7694,N_7251);
and U8224 (N_8224,N_7101,N_7162);
or U8225 (N_8225,N_6027,N_6218);
or U8226 (N_8226,N_6238,N_7154);
and U8227 (N_8227,N_6666,N_6090);
nand U8228 (N_8228,N_6084,N_6316);
or U8229 (N_8229,N_6509,N_7587);
or U8230 (N_8230,N_6411,N_7710);
nand U8231 (N_8231,N_7637,N_7062);
and U8232 (N_8232,N_6466,N_6880);
or U8233 (N_8233,N_6745,N_6303);
nand U8234 (N_8234,N_6739,N_7129);
nand U8235 (N_8235,N_6732,N_6811);
nor U8236 (N_8236,N_7814,N_6998);
or U8237 (N_8237,N_7636,N_6390);
and U8238 (N_8238,N_7883,N_7407);
nor U8239 (N_8239,N_7447,N_6104);
or U8240 (N_8240,N_6947,N_6410);
or U8241 (N_8241,N_6897,N_7704);
nor U8242 (N_8242,N_6293,N_7141);
or U8243 (N_8243,N_7588,N_7416);
and U8244 (N_8244,N_7701,N_6233);
nand U8245 (N_8245,N_6001,N_6529);
nand U8246 (N_8246,N_7102,N_6088);
or U8247 (N_8247,N_6237,N_7333);
nand U8248 (N_8248,N_6533,N_6846);
nand U8249 (N_8249,N_7267,N_6615);
and U8250 (N_8250,N_6387,N_7963);
and U8251 (N_8251,N_7265,N_6690);
nand U8252 (N_8252,N_6133,N_6126);
nor U8253 (N_8253,N_7514,N_7226);
or U8254 (N_8254,N_6016,N_6701);
xor U8255 (N_8255,N_7200,N_7402);
or U8256 (N_8256,N_7578,N_6669);
or U8257 (N_8257,N_7238,N_7870);
nor U8258 (N_8258,N_6453,N_7792);
nand U8259 (N_8259,N_6360,N_6605);
nor U8260 (N_8260,N_7851,N_7659);
nand U8261 (N_8261,N_7137,N_7194);
nand U8262 (N_8262,N_7515,N_7683);
and U8263 (N_8263,N_7470,N_6968);
nor U8264 (N_8264,N_6137,N_6535);
nor U8265 (N_8265,N_6925,N_7098);
and U8266 (N_8266,N_7737,N_6149);
or U8267 (N_8267,N_7299,N_7221);
or U8268 (N_8268,N_6750,N_6489);
xnor U8269 (N_8269,N_7035,N_6933);
and U8270 (N_8270,N_7766,N_6362);
nor U8271 (N_8271,N_6892,N_7175);
nor U8272 (N_8272,N_6011,N_7288);
and U8273 (N_8273,N_6785,N_7828);
and U8274 (N_8274,N_7069,N_6648);
nand U8275 (N_8275,N_7596,N_6668);
nand U8276 (N_8276,N_7689,N_7262);
nand U8277 (N_8277,N_6791,N_6953);
or U8278 (N_8278,N_6836,N_6940);
and U8279 (N_8279,N_7673,N_7071);
or U8280 (N_8280,N_7123,N_6216);
or U8281 (N_8281,N_6984,N_7159);
nand U8282 (N_8282,N_7785,N_7278);
and U8283 (N_8283,N_6217,N_7577);
nor U8284 (N_8284,N_6298,N_6567);
or U8285 (N_8285,N_6896,N_6552);
or U8286 (N_8286,N_6261,N_7183);
and U8287 (N_8287,N_6318,N_6145);
nand U8288 (N_8288,N_7249,N_7480);
nand U8289 (N_8289,N_6527,N_6043);
and U8290 (N_8290,N_7260,N_7034);
or U8291 (N_8291,N_6844,N_6635);
xor U8292 (N_8292,N_6747,N_6103);
nor U8293 (N_8293,N_7823,N_6503);
nor U8294 (N_8294,N_7755,N_6472);
nor U8295 (N_8295,N_6490,N_7531);
nor U8296 (N_8296,N_7564,N_7475);
nor U8297 (N_8297,N_7772,N_7641);
or U8298 (N_8298,N_6234,N_7317);
and U8299 (N_8299,N_7748,N_6708);
nand U8300 (N_8300,N_6291,N_6863);
nor U8301 (N_8301,N_7989,N_7424);
nor U8302 (N_8302,N_6748,N_7534);
or U8303 (N_8303,N_6308,N_6556);
nand U8304 (N_8304,N_6219,N_6731);
nand U8305 (N_8305,N_7006,N_6959);
or U8306 (N_8306,N_7728,N_7738);
or U8307 (N_8307,N_6664,N_6401);
or U8308 (N_8308,N_6997,N_6825);
and U8309 (N_8309,N_6704,N_6095);
or U8310 (N_8310,N_6003,N_6910);
nor U8311 (N_8311,N_6025,N_7796);
or U8312 (N_8312,N_6037,N_7490);
or U8313 (N_8313,N_6512,N_7340);
or U8314 (N_8314,N_6755,N_6833);
or U8315 (N_8315,N_6112,N_6426);
and U8316 (N_8316,N_7817,N_7324);
nor U8317 (N_8317,N_6271,N_7891);
nand U8318 (N_8318,N_7450,N_6670);
nand U8319 (N_8319,N_6331,N_6160);
or U8320 (N_8320,N_6840,N_7940);
or U8321 (N_8321,N_6761,N_7364);
or U8322 (N_8322,N_7974,N_7591);
or U8323 (N_8323,N_7176,N_6927);
and U8324 (N_8324,N_6530,N_6625);
or U8325 (N_8325,N_6876,N_6008);
and U8326 (N_8326,N_7732,N_7351);
nand U8327 (N_8327,N_6059,N_6372);
nand U8328 (N_8328,N_7920,N_7272);
or U8329 (N_8329,N_7916,N_7819);
or U8330 (N_8330,N_7574,N_7248);
or U8331 (N_8331,N_7273,N_6158);
nor U8332 (N_8332,N_7214,N_7662);
and U8333 (N_8333,N_7465,N_6712);
nand U8334 (N_8334,N_6941,N_6334);
or U8335 (N_8335,N_7090,N_7381);
nand U8336 (N_8336,N_7461,N_6772);
and U8337 (N_8337,N_6901,N_7695);
and U8338 (N_8338,N_6873,N_7182);
or U8339 (N_8339,N_6935,N_7496);
nand U8340 (N_8340,N_6168,N_7751);
nor U8341 (N_8341,N_7448,N_7508);
and U8342 (N_8342,N_6807,N_7051);
or U8343 (N_8343,N_7741,N_7672);
nand U8344 (N_8344,N_7544,N_7980);
nor U8345 (N_8345,N_6482,N_7087);
nand U8346 (N_8346,N_6970,N_7528);
or U8347 (N_8347,N_6790,N_7984);
or U8348 (N_8348,N_7861,N_6590);
and U8349 (N_8349,N_7499,N_7331);
and U8350 (N_8350,N_7663,N_6264);
nand U8351 (N_8351,N_7872,N_7854);
or U8352 (N_8352,N_6513,N_6364);
nor U8353 (N_8353,N_6333,N_6861);
and U8354 (N_8354,N_6824,N_6470);
and U8355 (N_8355,N_7733,N_6687);
nand U8356 (N_8356,N_7590,N_6882);
nand U8357 (N_8357,N_6614,N_6569);
nor U8358 (N_8358,N_6809,N_7463);
nand U8359 (N_8359,N_7932,N_6257);
or U8360 (N_8360,N_7453,N_7761);
or U8361 (N_8361,N_6779,N_6194);
and U8362 (N_8362,N_6107,N_6675);
nand U8363 (N_8363,N_6178,N_7982);
and U8364 (N_8364,N_7987,N_6464);
and U8365 (N_8365,N_6020,N_7990);
or U8366 (N_8366,N_7777,N_7838);
and U8367 (N_8367,N_6994,N_7795);
nand U8368 (N_8368,N_7130,N_6477);
and U8369 (N_8369,N_7745,N_7981);
nand U8370 (N_8370,N_7886,N_6726);
nand U8371 (N_8371,N_6633,N_7300);
nand U8372 (N_8372,N_6952,N_6938);
nor U8373 (N_8373,N_6123,N_6131);
and U8374 (N_8374,N_7995,N_7919);
nand U8375 (N_8375,N_7644,N_7793);
nor U8376 (N_8376,N_6292,N_7571);
nand U8377 (N_8377,N_7469,N_6017);
nor U8378 (N_8378,N_7147,N_7584);
xnor U8379 (N_8379,N_6546,N_7298);
nor U8380 (N_8380,N_6702,N_7100);
or U8381 (N_8381,N_7516,N_6138);
or U8382 (N_8382,N_6435,N_6777);
or U8383 (N_8383,N_6202,N_6843);
or U8384 (N_8384,N_6235,N_7612);
or U8385 (N_8385,N_7739,N_7054);
nand U8386 (N_8386,N_7057,N_7245);
or U8387 (N_8387,N_6760,N_7246);
and U8388 (N_8388,N_6055,N_7139);
nor U8389 (N_8389,N_6066,N_6800);
nor U8390 (N_8390,N_7715,N_6943);
and U8391 (N_8391,N_6999,N_6374);
nand U8392 (N_8392,N_7740,N_7548);
nor U8393 (N_8393,N_7497,N_6547);
nand U8394 (N_8394,N_6209,N_6734);
or U8395 (N_8395,N_7527,N_7700);
or U8396 (N_8396,N_6351,N_6538);
nand U8397 (N_8397,N_6619,N_7365);
nand U8398 (N_8398,N_6139,N_7965);
nor U8399 (N_8399,N_7218,N_7395);
or U8400 (N_8400,N_7804,N_6954);
nand U8401 (N_8401,N_6161,N_7112);
or U8402 (N_8402,N_7633,N_6042);
and U8403 (N_8403,N_6787,N_7457);
nand U8404 (N_8404,N_6608,N_6474);
or U8405 (N_8405,N_6239,N_7546);
nand U8406 (N_8406,N_7911,N_7569);
and U8407 (N_8407,N_6888,N_7959);
nand U8408 (N_8408,N_6818,N_6821);
nand U8409 (N_8409,N_7321,N_7291);
and U8410 (N_8410,N_7138,N_6125);
nor U8411 (N_8411,N_7947,N_7782);
nand U8412 (N_8412,N_7882,N_7166);
nor U8413 (N_8413,N_6408,N_7043);
or U8414 (N_8414,N_7653,N_7730);
or U8415 (N_8415,N_6300,N_6960);
nand U8416 (N_8416,N_7786,N_7708);
nor U8417 (N_8417,N_7345,N_7053);
or U8418 (N_8418,N_6344,N_6665);
or U8419 (N_8419,N_7266,N_6548);
and U8420 (N_8420,N_7908,N_6644);
or U8421 (N_8421,N_7359,N_7459);
and U8422 (N_8422,N_6048,N_6192);
nor U8423 (N_8423,N_6079,N_6847);
nand U8424 (N_8424,N_6320,N_7334);
nand U8425 (N_8425,N_6598,N_7605);
nor U8426 (N_8426,N_7338,N_7086);
nand U8427 (N_8427,N_6729,N_7316);
or U8428 (N_8428,N_6195,N_7134);
nand U8429 (N_8429,N_6877,N_7509);
or U8430 (N_8430,N_7976,N_6151);
nand U8431 (N_8431,N_6592,N_6199);
or U8432 (N_8432,N_6707,N_7611);
or U8433 (N_8433,N_7640,N_7639);
nor U8434 (N_8434,N_6493,N_6343);
nand U8435 (N_8435,N_6950,N_6210);
and U8436 (N_8436,N_6386,N_6346);
xor U8437 (N_8437,N_6932,N_6709);
and U8438 (N_8438,N_6979,N_6012);
nand U8439 (N_8439,N_6754,N_6400);
and U8440 (N_8440,N_7764,N_6589);
or U8441 (N_8441,N_7002,N_6705);
or U8442 (N_8442,N_6328,N_6211);
nor U8443 (N_8443,N_6051,N_6119);
or U8444 (N_8444,N_7092,N_6033);
and U8445 (N_8445,N_7839,N_6280);
or U8446 (N_8446,N_6093,N_7115);
and U8447 (N_8447,N_6976,N_7127);
nand U8448 (N_8448,N_6399,N_6100);
nand U8449 (N_8449,N_6671,N_6826);
or U8450 (N_8450,N_6097,N_6041);
or U8451 (N_8451,N_7089,N_6223);
nor U8452 (N_8452,N_7373,N_6200);
or U8453 (N_8453,N_7961,N_7389);
nor U8454 (N_8454,N_6864,N_7412);
nand U8455 (N_8455,N_7217,N_7018);
or U8456 (N_8456,N_6440,N_7027);
nand U8457 (N_8457,N_7802,N_6663);
or U8458 (N_8458,N_7252,N_7513);
or U8459 (N_8459,N_6699,N_6278);
and U8460 (N_8460,N_6875,N_7203);
nand U8461 (N_8461,N_6006,N_7435);
or U8462 (N_8462,N_6313,N_7095);
and U8463 (N_8463,N_7394,N_7973);
nand U8464 (N_8464,N_7293,N_6520);
or U8465 (N_8465,N_6269,N_7621);
nor U8466 (N_8466,N_6969,N_7408);
or U8467 (N_8467,N_6431,N_6593);
or U8468 (N_8468,N_6966,N_6559);
nand U8469 (N_8469,N_6595,N_7914);
and U8470 (N_8470,N_6297,N_7206);
nand U8471 (N_8471,N_6949,N_7231);
and U8472 (N_8472,N_6190,N_6555);
nor U8473 (N_8473,N_7320,N_7014);
nand U8474 (N_8474,N_7805,N_7679);
or U8475 (N_8475,N_6166,N_7744);
or U8476 (N_8476,N_6098,N_6746);
and U8477 (N_8477,N_7474,N_6394);
nor U8478 (N_8478,N_6266,N_6713);
and U8479 (N_8479,N_7688,N_7593);
and U8480 (N_8480,N_6723,N_7372);
and U8481 (N_8481,N_7749,N_7385);
nand U8482 (N_8482,N_7702,N_7401);
nand U8483 (N_8483,N_7536,N_7337);
nand U8484 (N_8484,N_6594,N_7966);
nand U8485 (N_8485,N_6730,N_7482);
nand U8486 (N_8486,N_6814,N_7479);
nand U8487 (N_8487,N_7254,N_6672);
nor U8488 (N_8488,N_7227,N_6176);
nor U8489 (N_8489,N_7116,N_7880);
and U8490 (N_8490,N_6111,N_7275);
nor U8491 (N_8491,N_7243,N_6607);
and U8492 (N_8492,N_6869,N_7613);
nor U8493 (N_8493,N_7437,N_7526);
nand U8494 (N_8494,N_7628,N_7301);
nand U8495 (N_8495,N_7844,N_7369);
or U8496 (N_8496,N_6560,N_6222);
nor U8497 (N_8497,N_7396,N_6247);
and U8498 (N_8498,N_7869,N_6767);
or U8499 (N_8499,N_7563,N_6915);
nand U8500 (N_8500,N_6573,N_7572);
xnor U8501 (N_8501,N_7444,N_6642);
or U8502 (N_8502,N_7815,N_7747);
or U8503 (N_8503,N_7488,N_6322);
and U8504 (N_8504,N_7199,N_6184);
or U8505 (N_8505,N_6304,N_6786);
nand U8506 (N_8506,N_7193,N_7555);
nand U8507 (N_8507,N_7033,N_7209);
nand U8508 (N_8508,N_7117,N_6254);
or U8509 (N_8509,N_6841,N_7380);
nand U8510 (N_8510,N_6574,N_7939);
and U8511 (N_8511,N_7718,N_7511);
or U8512 (N_8512,N_6577,N_7282);
nor U8513 (N_8513,N_7081,N_6359);
or U8514 (N_8514,N_7205,N_7234);
and U8515 (N_8515,N_6801,N_6491);
nand U8516 (N_8516,N_6430,N_6827);
nor U8517 (N_8517,N_7957,N_6167);
nor U8518 (N_8518,N_6770,N_7436);
and U8519 (N_8519,N_6402,N_6245);
or U8520 (N_8520,N_7884,N_6661);
or U8521 (N_8521,N_7557,N_7757);
nor U8522 (N_8522,N_7709,N_6356);
or U8523 (N_8523,N_6481,N_6288);
nor U8524 (N_8524,N_6689,N_7215);
or U8525 (N_8525,N_7362,N_7618);
nand U8526 (N_8526,N_6429,N_6268);
nor U8527 (N_8527,N_6312,N_6265);
or U8528 (N_8528,N_6926,N_7674);
nor U8529 (N_8529,N_7004,N_6204);
nor U8530 (N_8530,N_7650,N_7820);
nand U8531 (N_8531,N_6444,N_7430);
or U8532 (N_8532,N_6946,N_6259);
or U8533 (N_8533,N_6185,N_7893);
nor U8534 (N_8534,N_6385,N_7195);
nand U8535 (N_8535,N_7760,N_7242);
nor U8536 (N_8536,N_6964,N_6643);
or U8537 (N_8537,N_7366,N_6859);
nand U8538 (N_8538,N_6616,N_7856);
or U8539 (N_8539,N_6780,N_7378);
nand U8540 (N_8540,N_6673,N_7042);
nor U8541 (N_8541,N_6306,N_6053);
nand U8542 (N_8542,N_7910,N_6545);
nand U8543 (N_8543,N_7007,N_6422);
nand U8544 (N_8544,N_6255,N_6722);
nor U8545 (N_8545,N_7993,N_7477);
and U8546 (N_8546,N_7857,N_7622);
and U8547 (N_8547,N_7342,N_6542);
or U8548 (N_8548,N_7615,N_6522);
nor U8549 (N_8549,N_7198,N_7609);
and U8550 (N_8550,N_7440,N_6986);
or U8551 (N_8551,N_7425,N_7931);
xor U8552 (N_8552,N_6991,N_6067);
or U8553 (N_8553,N_6118,N_6524);
nand U8554 (N_8554,N_7239,N_7756);
nand U8555 (N_8555,N_6081,N_7070);
nor U8556 (N_8556,N_6911,N_7877);
nand U8557 (N_8557,N_7552,N_6068);
and U8558 (N_8558,N_7005,N_7778);
nor U8559 (N_8559,N_6407,N_6326);
and U8560 (N_8560,N_7332,N_7549);
and U8561 (N_8561,N_7502,N_6515);
nor U8562 (N_8562,N_7888,N_6808);
nand U8563 (N_8563,N_7286,N_6015);
nor U8564 (N_8564,N_7292,N_7901);
nor U8565 (N_8565,N_6189,N_7505);
nor U8566 (N_8566,N_7322,N_6488);
or U8567 (N_8567,N_7826,N_6014);
or U8568 (N_8568,N_7039,N_7602);
nand U8569 (N_8569,N_7818,N_7648);
and U8570 (N_8570,N_6816,N_6651);
or U8571 (N_8571,N_6822,N_6942);
or U8572 (N_8572,N_6889,N_6377);
or U8573 (N_8573,N_6307,N_7271);
nor U8574 (N_8574,N_6206,N_6227);
and U8575 (N_8575,N_6317,N_6368);
and U8576 (N_8576,N_6465,N_7314);
nand U8577 (N_8577,N_6913,N_7390);
and U8578 (N_8578,N_7375,N_7111);
nand U8579 (N_8579,N_7406,N_7885);
and U8580 (N_8580,N_7507,N_7026);
and U8581 (N_8581,N_6073,N_7692);
nand U8582 (N_8582,N_6871,N_7196);
and U8583 (N_8583,N_6094,N_6467);
or U8584 (N_8584,N_7923,N_6855);
or U8585 (N_8585,N_7994,N_7767);
and U8586 (N_8586,N_7660,N_6832);
or U8587 (N_8587,N_7313,N_7806);
nor U8588 (N_8588,N_7951,N_6010);
or U8589 (N_8589,N_6921,N_6568);
nand U8590 (N_8590,N_7779,N_6380);
nor U8591 (N_8591,N_6620,N_6497);
nand U8592 (N_8592,N_6135,N_6696);
nand U8593 (N_8593,N_7899,N_6365);
and U8594 (N_8594,N_6005,N_7279);
nor U8595 (N_8595,N_6230,N_6463);
or U8596 (N_8596,N_6738,N_7543);
nor U8597 (N_8597,N_6175,N_7156);
or U8598 (N_8598,N_7560,N_6062);
nor U8599 (N_8599,N_6142,N_6471);
and U8600 (N_8600,N_7106,N_7803);
nand U8601 (N_8601,N_7264,N_6891);
or U8602 (N_8602,N_6868,N_6371);
or U8603 (N_8603,N_7763,N_6829);
nor U8604 (N_8604,N_6056,N_7419);
nand U8605 (N_8605,N_6715,N_7922);
nor U8606 (N_8606,N_7800,N_6581);
nor U8607 (N_8607,N_6835,N_7759);
or U8608 (N_8608,N_6296,N_7307);
or U8609 (N_8609,N_6302,N_7295);
xnor U8610 (N_8610,N_7025,N_7754);
and U8611 (N_8611,N_6058,N_7237);
nand U8612 (N_8612,N_6934,N_6603);
nor U8613 (N_8613,N_7594,N_7638);
nand U8614 (N_8614,N_7788,N_6990);
nand U8615 (N_8615,N_7592,N_7343);
nand U8616 (N_8616,N_7060,N_7017);
and U8617 (N_8617,N_6817,N_7077);
or U8618 (N_8618,N_7657,N_6434);
nor U8619 (N_8619,N_6939,N_7179);
nand U8620 (N_8620,N_7097,N_6253);
and U8621 (N_8621,N_6526,N_7021);
nand U8622 (N_8622,N_7934,N_6982);
and U8623 (N_8623,N_7775,N_6842);
and U8624 (N_8624,N_7258,N_7318);
or U8625 (N_8625,N_7446,N_7483);
nor U8626 (N_8626,N_6627,N_7216);
and U8627 (N_8627,N_6759,N_6108);
or U8628 (N_8628,N_6281,N_6283);
and U8629 (N_8629,N_7329,N_7913);
nand U8630 (N_8630,N_7868,N_7685);
nor U8631 (N_8631,N_7274,N_6366);
nand U8632 (N_8632,N_7132,N_7864);
nor U8633 (N_8633,N_7308,N_7532);
nand U8634 (N_8634,N_7576,N_7208);
and U8635 (N_8635,N_7400,N_7493);
or U8636 (N_8636,N_7859,N_7830);
nand U8637 (N_8637,N_7562,N_6854);
or U8638 (N_8638,N_6267,N_6793);
and U8639 (N_8639,N_7355,N_7119);
nor U8640 (N_8640,N_6909,N_7336);
and U8641 (N_8641,N_7833,N_6725);
and U8642 (N_8642,N_7341,N_7451);
or U8643 (N_8643,N_6191,N_6282);
nand U8644 (N_8644,N_6628,N_7714);
nor U8645 (N_8645,N_7742,N_6207);
and U8646 (N_8646,N_7367,N_6951);
nor U8647 (N_8647,N_7427,N_7438);
nor U8648 (N_8648,N_6792,N_7933);
nor U8649 (N_8649,N_7691,N_6992);
or U8650 (N_8650,N_6681,N_7567);
nor U8651 (N_8651,N_6564,N_6886);
nand U8652 (N_8652,N_6295,N_7978);
or U8653 (N_8653,N_6539,N_6565);
or U8654 (N_8654,N_7056,N_6114);
nor U8655 (N_8655,N_7523,N_6468);
or U8656 (N_8656,N_7642,N_7681);
and U8657 (N_8657,N_7647,N_7808);
nor U8658 (N_8658,N_7941,N_6980);
nand U8659 (N_8659,N_6250,N_6658);
nand U8660 (N_8660,N_6405,N_7420);
nand U8661 (N_8661,N_6096,N_6369);
or U8662 (N_8662,N_7506,N_7085);
or U8663 (N_8663,N_7753,N_6469);
and U8664 (N_8664,N_7918,N_6035);
and U8665 (N_8665,N_6023,N_6865);
nor U8666 (N_8666,N_6905,N_6858);
or U8667 (N_8667,N_7835,N_6609);
nand U8668 (N_8668,N_7065,N_7131);
nand U8669 (N_8669,N_7960,N_7096);
nor U8670 (N_8670,N_7241,N_6071);
and U8671 (N_8671,N_7969,N_6971);
nand U8672 (N_8672,N_6517,N_7335);
nor U8673 (N_8673,N_6113,N_6174);
or U8674 (N_8674,N_7312,N_7174);
and U8675 (N_8675,N_6350,N_6667);
nand U8676 (N_8676,N_7656,N_6967);
nor U8677 (N_8677,N_6657,N_7630);
nor U8678 (N_8678,N_6582,N_6370);
and U8679 (N_8679,N_6341,N_6479);
nor U8680 (N_8680,N_6397,N_7729);
and U8681 (N_8681,N_6336,N_7986);
nand U8682 (N_8682,N_6454,N_6284);
nor U8683 (N_8683,N_6514,N_6127);
or U8684 (N_8684,N_7600,N_7887);
nand U8685 (N_8685,N_7379,N_7568);
and U8686 (N_8686,N_6799,N_7067);
nor U8687 (N_8687,N_6783,N_6427);
or U8688 (N_8688,N_7620,N_7810);
and U8689 (N_8689,N_6150,N_6403);
and U8690 (N_8690,N_6662,N_7794);
or U8691 (N_8691,N_6077,N_7696);
nand U8692 (N_8692,N_6428,N_6256);
nand U8693 (N_8693,N_6196,N_7693);
and U8694 (N_8694,N_7790,N_7384);
nand U8695 (N_8695,N_6169,N_6610);
or U8696 (N_8696,N_7664,N_7041);
and U8697 (N_8697,N_7881,N_6996);
nand U8698 (N_8698,N_6563,N_6446);
and U8699 (N_8699,N_7827,N_6367);
nand U8700 (N_8700,N_6812,N_6375);
xnor U8701 (N_8701,N_6423,N_6507);
nor U8702 (N_8702,N_6274,N_6776);
nand U8703 (N_8703,N_6221,N_7487);
and U8704 (N_8704,N_6277,N_6962);
nor U8705 (N_8705,N_7353,N_7387);
and U8706 (N_8706,N_6258,N_6226);
nor U8707 (N_8707,N_7491,N_7149);
nand U8708 (N_8708,N_6404,N_7171);
nor U8709 (N_8709,N_6751,N_7860);
nand U8710 (N_8710,N_6009,N_7180);
nand U8711 (N_8711,N_7936,N_7537);
or U8712 (N_8712,N_6345,N_7629);
nor U8713 (N_8713,N_6771,N_6323);
and U8714 (N_8714,N_6782,N_7727);
or U8715 (N_8715,N_7133,N_6887);
nor U8716 (N_8716,N_6361,N_6930);
nand U8717 (N_8717,N_6753,N_6562);
nor U8718 (N_8718,N_7906,N_6379);
nand U8719 (N_8719,N_6457,N_6243);
xor U8720 (N_8720,N_6695,N_7853);
and U8721 (N_8721,N_6972,N_7944);
or U8722 (N_8722,N_7371,N_6475);
and U8723 (N_8723,N_7404,N_7235);
nand U8724 (N_8724,N_6148,N_6773);
nand U8725 (N_8725,N_7846,N_6965);
or U8726 (N_8726,N_7374,N_6778);
and U8727 (N_8727,N_7063,N_7686);
nor U8728 (N_8728,N_7413,N_7177);
nand U8729 (N_8729,N_7411,N_6162);
nand U8730 (N_8730,N_7122,N_7084);
nand U8731 (N_8731,N_7962,N_6083);
nor U8732 (N_8732,N_7376,N_6611);
nor U8733 (N_8733,N_7992,N_7409);
nand U8734 (N_8734,N_6639,N_6384);
nand U8735 (N_8735,N_6736,N_6872);
xor U8736 (N_8736,N_7302,N_6335);
nand U8737 (N_8737,N_7917,N_7787);
and U8738 (N_8738,N_6898,N_6617);
nand U8739 (N_8739,N_7928,N_7066);
nor U8740 (N_8740,N_7813,N_7315);
or U8741 (N_8741,N_6516,N_6511);
nor U8742 (N_8742,N_7791,N_7046);
nand U8743 (N_8743,N_7675,N_6796);
nand U8744 (N_8744,N_6324,N_6260);
and U8745 (N_8745,N_7019,N_7943);
or U8746 (N_8746,N_7684,N_7529);
nand U8747 (N_8747,N_7073,N_6645);
nand U8748 (N_8748,N_7382,N_7712);
nand U8749 (N_8749,N_7719,N_6900);
nand U8750 (N_8750,N_6441,N_7422);
or U8751 (N_8751,N_7871,N_7220);
and U8752 (N_8752,N_7303,N_6393);
nor U8753 (N_8753,N_6558,N_6492);
and U8754 (N_8754,N_7968,N_6276);
or U8755 (N_8755,N_6040,N_6007);
or U8756 (N_8756,N_7553,N_6928);
nand U8757 (N_8757,N_6599,N_7711);
or U8758 (N_8758,N_6505,N_6236);
nor U8759 (N_8759,N_6540,N_7821);
or U8760 (N_8760,N_6624,N_6353);
and U8761 (N_8761,N_6155,N_6895);
nor U8762 (N_8762,N_6478,N_6252);
or U8763 (N_8763,N_7938,N_6373);
and U8764 (N_8764,N_6716,N_7624);
nor U8765 (N_8765,N_7012,N_6908);
and U8766 (N_8766,N_6557,N_7892);
and U8767 (N_8767,N_7155,N_6523);
or U8768 (N_8768,N_6458,N_6815);
and U8769 (N_8769,N_7186,N_6415);
nor U8770 (N_8770,N_6870,N_7126);
nor U8771 (N_8771,N_7256,N_7128);
nor U8772 (N_8772,N_6637,N_6085);
xor U8773 (N_8773,N_6831,N_7210);
and U8774 (N_8774,N_6977,N_7328);
nand U8775 (N_8775,N_7426,N_6032);
and U8776 (N_8776,N_6893,N_6286);
or U8777 (N_8777,N_7845,N_6198);
or U8778 (N_8778,N_7068,N_6683);
or U8779 (N_8779,N_7061,N_7580);
or U8780 (N_8780,N_7850,N_7201);
nor U8781 (N_8781,N_7476,N_7768);
and U8782 (N_8782,N_7717,N_6904);
or U8783 (N_8783,N_6376,N_6275);
nand U8784 (N_8784,N_6122,N_7774);
and U8785 (N_8785,N_6363,N_7520);
nor U8786 (N_8786,N_7284,N_6553);
nor U8787 (N_8787,N_7125,N_6456);
or U8788 (N_8788,N_7213,N_6078);
nand U8789 (N_8789,N_7598,N_7484);
nor U8790 (N_8790,N_7059,N_6682);
nor U8791 (N_8791,N_6381,N_7013);
or U8792 (N_8792,N_6613,N_6183);
or U8793 (N_8793,N_6775,N_6902);
and U8794 (N_8794,N_7619,N_7623);
or U8795 (N_8795,N_6774,N_7503);
nand U8796 (N_8796,N_6173,N_6249);
and U8797 (N_8797,N_7541,N_6418);
or U8798 (N_8798,N_7927,N_6065);
or U8799 (N_8799,N_7202,N_6413);
and U8800 (N_8800,N_7164,N_7902);
or U8801 (N_8801,N_7841,N_6406);
nand U8802 (N_8802,N_7319,N_6494);
and U8803 (N_8803,N_6566,N_7011);
nor U8804 (N_8804,N_7837,N_7114);
nand U8805 (N_8805,N_6229,N_7542);
or U8806 (N_8806,N_6988,N_6685);
nand U8807 (N_8807,N_7229,N_7481);
xor U8808 (N_8808,N_6186,N_6680);
nor U8809 (N_8809,N_7082,N_7677);
and U8810 (N_8810,N_6074,N_6679);
and U8811 (N_8811,N_6924,N_7608);
and U8812 (N_8812,N_6798,N_6874);
and U8813 (N_8813,N_7758,N_7495);
nand U8814 (N_8814,N_6241,N_7595);
nand U8815 (N_8815,N_7894,N_7410);
or U8816 (N_8816,N_7099,N_6433);
nor U8817 (N_8817,N_6038,N_7535);
nand U8818 (N_8818,N_7309,N_6678);
and U8819 (N_8819,N_6330,N_7661);
or U8820 (N_8820,N_6391,N_7521);
and U8821 (N_8821,N_6117,N_7443);
and U8822 (N_8822,N_6845,N_7703);
nand U8823 (N_8823,N_7625,N_6072);
nand U8824 (N_8824,N_7392,N_6502);
or U8825 (N_8825,N_7290,N_7044);
or U8826 (N_8826,N_7512,N_6358);
and U8827 (N_8827,N_7219,N_6586);
and U8828 (N_8828,N_6000,N_7165);
nand U8829 (N_8829,N_6451,N_7807);
and U8830 (N_8830,N_7878,N_6766);
or U8831 (N_8831,N_7439,N_6076);
nand U8832 (N_8832,N_7627,N_6717);
nor U8833 (N_8833,N_6879,N_7646);
or U8834 (N_8834,N_6806,N_7979);
and U8835 (N_8835,N_7289,N_7517);
or U8836 (N_8836,N_6602,N_6866);
nor U8837 (N_8837,N_6848,N_7970);
nor U8838 (N_8838,N_7360,N_7874);
xor U8839 (N_8839,N_6172,N_7848);
nor U8840 (N_8840,N_7000,N_6036);
nor U8841 (N_8841,N_6197,N_7350);
and U8842 (N_8842,N_6170,N_6820);
and U8843 (N_8843,N_7305,N_7904);
and U8844 (N_8844,N_6851,N_6052);
and U8845 (N_8845,N_7504,N_6116);
and U8846 (N_8846,N_7189,N_7255);
nand U8847 (N_8847,N_7614,N_6339);
or U8848 (N_8848,N_7896,N_6944);
and U8849 (N_8849,N_6447,N_6436);
or U8850 (N_8850,N_6837,N_6718);
nor U8851 (N_8851,N_7094,N_6106);
or U8852 (N_8852,N_7632,N_7847);
nand U8853 (N_8853,N_7971,N_6034);
or U8854 (N_8854,N_6270,N_6630);
and U8855 (N_8855,N_6987,N_6164);
or U8856 (N_8856,N_7354,N_7539);
and U8857 (N_8857,N_7533,N_6596);
or U8858 (N_8858,N_6089,N_7421);
and U8859 (N_8859,N_6496,N_6128);
nor U8860 (N_8860,N_6329,N_6591);
and U8861 (N_8861,N_7720,N_6993);
nor U8862 (N_8862,N_6724,N_6417);
nor U8863 (N_8863,N_7770,N_6028);
or U8864 (N_8864,N_6338,N_7706);
or U8865 (N_8865,N_6804,N_7233);
nor U8866 (N_8866,N_6382,N_7152);
nor U8867 (N_8867,N_7142,N_6830);
and U8868 (N_8868,N_7776,N_7236);
or U8869 (N_8869,N_7230,N_7197);
xor U8870 (N_8870,N_6789,N_7415);
nor U8871 (N_8871,N_6231,N_6694);
nor U8872 (N_8872,N_6764,N_7232);
nor U8873 (N_8873,N_6311,N_7559);
and U8874 (N_8874,N_7698,N_6576);
nor U8875 (N_8875,N_7525,N_6597);
nand U8876 (N_8876,N_6660,N_6881);
or U8877 (N_8877,N_6022,N_7181);
nor U8878 (N_8878,N_7368,N_7250);
nand U8879 (N_8879,N_7743,N_7524);
nand U8880 (N_8880,N_6906,N_6583);
and U8881 (N_8881,N_7875,N_7566);
or U8882 (N_8882,N_7075,N_6838);
and U8883 (N_8883,N_7829,N_7326);
and U8884 (N_8884,N_6728,N_7635);
nand U8885 (N_8885,N_6917,N_6455);
nand U8886 (N_8886,N_7048,N_7645);
or U8887 (N_8887,N_6047,N_7357);
and U8888 (N_8888,N_6450,N_6484);
or U8889 (N_8889,N_7895,N_7418);
or U8890 (N_8890,N_7889,N_6537);
nand U8891 (N_8891,N_6289,N_6606);
nand U8892 (N_8892,N_7455,N_6504);
nor U8893 (N_8893,N_7671,N_6272);
nor U8894 (N_8894,N_7397,N_7339);
or U8895 (N_8895,N_7349,N_6752);
nand U8896 (N_8896,N_7431,N_7148);
nand U8897 (N_8897,N_6600,N_6937);
or U8898 (N_8898,N_7956,N_6347);
nor U8899 (N_8899,N_7022,N_6242);
and U8900 (N_8900,N_6819,N_7283);
xnor U8901 (N_8901,N_6224,N_6416);
or U8902 (N_8902,N_7501,N_7172);
nor U8903 (N_8903,N_7583,N_6521);
and U8904 (N_8904,N_6340,N_7456);
nor U8905 (N_8905,N_7725,N_6929);
nand U8906 (N_8906,N_7016,N_7038);
nand U8907 (N_8907,N_6584,N_6528);
or U8908 (N_8908,N_6029,N_6963);
nor U8909 (N_8909,N_6758,N_6721);
nor U8910 (N_8910,N_7297,N_6332);
nor U8911 (N_8911,N_6075,N_7277);
nor U8912 (N_8912,N_6551,N_6049);
nand U8913 (N_8913,N_7530,N_7429);
and U8914 (N_8914,N_7654,N_7377);
xor U8915 (N_8915,N_7985,N_7597);
nor U8916 (N_8916,N_7842,N_7707);
xor U8917 (N_8917,N_6656,N_6443);
and U8918 (N_8918,N_6579,N_7093);
and U8919 (N_8919,N_7649,N_6378);
nor U8920 (N_8920,N_7616,N_7188);
and U8921 (N_8921,N_7554,N_7909);
nand U8922 (N_8922,N_6439,N_7682);
nor U8923 (N_8923,N_6473,N_7145);
nor U8924 (N_8924,N_7423,N_6588);
nor U8925 (N_8925,N_6419,N_7185);
nand U8926 (N_8926,N_7500,N_6026);
nand U8927 (N_8927,N_6802,N_7825);
or U8928 (N_8928,N_7610,N_6445);
and U8929 (N_8929,N_6646,N_7955);
nand U8930 (N_8930,N_7327,N_6781);
nand U8931 (N_8931,N_7736,N_7518);
or U8932 (N_8932,N_7676,N_6279);
nand U8933 (N_8933,N_7670,N_6839);
or U8934 (N_8934,N_7799,N_7428);
or U8935 (N_8935,N_6086,N_6549);
nor U8936 (N_8936,N_6674,N_7121);
and U8937 (N_8937,N_7726,N_6159);
and U8938 (N_8938,N_6649,N_7280);
or U8939 (N_8939,N_7953,N_6756);
nor U8940 (N_8940,N_7153,N_7383);
or U8941 (N_8941,N_7972,N_6849);
nand U8942 (N_8942,N_7222,N_7863);
nor U8943 (N_8943,N_6030,N_7192);
nand U8944 (N_8944,N_7752,N_7468);
nor U8945 (N_8945,N_6686,N_7287);
nor U8946 (N_8946,N_7843,N_6885);
or U8947 (N_8947,N_6273,N_7570);
and U8948 (N_8948,N_7144,N_7948);
nor U8949 (N_8949,N_6290,N_6632);
xnor U8950 (N_8950,N_7472,N_7573);
and U8951 (N_8951,N_7163,N_6706);
nor U8952 (N_8952,N_6890,N_6082);
and U8953 (N_8953,N_6102,N_7388);
or U8954 (N_8954,N_7949,N_7361);
nor U8955 (N_8955,N_6688,N_7454);
or U8956 (N_8956,N_7143,N_7652);
and U8957 (N_8957,N_6903,N_7816);
nand U8958 (N_8958,N_7498,N_6004);
or U8959 (N_8959,N_7655,N_7935);
nand U8960 (N_8960,N_6659,N_6544);
nor U8961 (N_8961,N_7634,N_7997);
and U8962 (N_8962,N_7135,N_6856);
or U8963 (N_8963,N_6220,N_7263);
nor U8964 (N_8964,N_6388,N_7485);
and U8965 (N_8965,N_6099,N_6495);
nand U8966 (N_8966,N_6506,N_6412);
nand U8967 (N_8967,N_6720,N_7003);
or U8968 (N_8968,N_7296,N_7836);
or U8969 (N_8969,N_7393,N_6136);
or U8970 (N_8970,N_6698,N_6021);
nor U8971 (N_8971,N_7991,N_6215);
nand U8972 (N_8972,N_7964,N_6263);
and U8973 (N_8973,N_6604,N_7204);
nor U8974 (N_8974,N_7074,N_6057);
or U8975 (N_8975,N_6623,N_7023);
nor U8976 (N_8976,N_7008,N_6587);
nand U8977 (N_8977,N_7306,N_6063);
nand U8978 (N_8978,N_7907,N_7606);
nor U8979 (N_8979,N_7721,N_6299);
nor U8980 (N_8980,N_6188,N_7716);
nand U8981 (N_8981,N_6945,N_7651);
or U8982 (N_8982,N_6733,N_6087);
or U8983 (N_8983,N_7040,N_6978);
nor U8984 (N_8984,N_6121,N_7545);
nor U8985 (N_8985,N_6442,N_6246);
nand U8986 (N_8986,N_7849,N_6181);
or U8987 (N_8987,N_7840,N_6571);
nor U8988 (N_8988,N_6179,N_6561);
and U8989 (N_8989,N_7460,N_6743);
nand U8990 (N_8990,N_6208,N_7952);
or U8991 (N_8991,N_7050,N_7103);
nor U8992 (N_8992,N_6640,N_7999);
or U8993 (N_8993,N_7347,N_7160);
and U8994 (N_8994,N_6862,N_6711);
nor U8995 (N_8995,N_6132,N_6570);
and U8996 (N_8996,N_7449,N_7080);
and U8997 (N_8997,N_6342,N_7929);
and U8998 (N_8998,N_6580,N_7765);
xnor U8999 (N_8999,N_6857,N_7157);
or U9000 (N_9000,N_6804,N_7381);
nor U9001 (N_9001,N_6815,N_6883);
and U9002 (N_9002,N_6801,N_7175);
or U9003 (N_9003,N_7035,N_6136);
or U9004 (N_9004,N_7961,N_7856);
or U9005 (N_9005,N_7689,N_7545);
nand U9006 (N_9006,N_7068,N_6864);
nand U9007 (N_9007,N_7823,N_6528);
or U9008 (N_9008,N_6684,N_6251);
and U9009 (N_9009,N_7617,N_6777);
and U9010 (N_9010,N_6898,N_7574);
nor U9011 (N_9011,N_6098,N_6937);
and U9012 (N_9012,N_6096,N_6364);
nand U9013 (N_9013,N_6689,N_7082);
nand U9014 (N_9014,N_7074,N_7187);
and U9015 (N_9015,N_7853,N_6522);
or U9016 (N_9016,N_7413,N_7637);
and U9017 (N_9017,N_6773,N_7209);
and U9018 (N_9018,N_7981,N_7995);
nand U9019 (N_9019,N_7609,N_7911);
or U9020 (N_9020,N_6356,N_6831);
and U9021 (N_9021,N_6072,N_6864);
or U9022 (N_9022,N_7297,N_7860);
nand U9023 (N_9023,N_6176,N_7106);
or U9024 (N_9024,N_7865,N_7085);
nand U9025 (N_9025,N_6873,N_7037);
nor U9026 (N_9026,N_6941,N_7675);
or U9027 (N_9027,N_7551,N_6436);
nor U9028 (N_9028,N_7376,N_6391);
and U9029 (N_9029,N_6420,N_7864);
nand U9030 (N_9030,N_7141,N_7968);
and U9031 (N_9031,N_7179,N_6273);
nand U9032 (N_9032,N_6584,N_6837);
and U9033 (N_9033,N_7403,N_6347);
nor U9034 (N_9034,N_7038,N_7504);
nor U9035 (N_9035,N_6689,N_7513);
nand U9036 (N_9036,N_6981,N_6137);
nor U9037 (N_9037,N_6817,N_7236);
and U9038 (N_9038,N_6165,N_7475);
nor U9039 (N_9039,N_6228,N_6005);
or U9040 (N_9040,N_7489,N_7708);
or U9041 (N_9041,N_6557,N_7084);
and U9042 (N_9042,N_6681,N_7331);
nand U9043 (N_9043,N_7978,N_6452);
nand U9044 (N_9044,N_7950,N_7268);
and U9045 (N_9045,N_7198,N_6390);
and U9046 (N_9046,N_6874,N_7340);
and U9047 (N_9047,N_6181,N_6546);
nor U9048 (N_9048,N_7596,N_6096);
nor U9049 (N_9049,N_7099,N_6614);
nand U9050 (N_9050,N_6873,N_6163);
nand U9051 (N_9051,N_7322,N_6036);
nand U9052 (N_9052,N_7124,N_7090);
and U9053 (N_9053,N_7471,N_6087);
and U9054 (N_9054,N_6808,N_6458);
nor U9055 (N_9055,N_7686,N_7019);
nand U9056 (N_9056,N_7522,N_7083);
nand U9057 (N_9057,N_6608,N_6642);
or U9058 (N_9058,N_7890,N_7430);
nor U9059 (N_9059,N_6583,N_6278);
nand U9060 (N_9060,N_7342,N_7658);
nand U9061 (N_9061,N_6573,N_6070);
or U9062 (N_9062,N_7158,N_6142);
and U9063 (N_9063,N_7048,N_6971);
or U9064 (N_9064,N_6070,N_7258);
and U9065 (N_9065,N_6981,N_6559);
or U9066 (N_9066,N_6133,N_6927);
or U9067 (N_9067,N_7153,N_7166);
and U9068 (N_9068,N_6431,N_6937);
and U9069 (N_9069,N_6934,N_7428);
and U9070 (N_9070,N_7959,N_7380);
and U9071 (N_9071,N_7219,N_7021);
and U9072 (N_9072,N_7503,N_7076);
nor U9073 (N_9073,N_6232,N_7212);
nor U9074 (N_9074,N_6807,N_6099);
and U9075 (N_9075,N_6019,N_7136);
and U9076 (N_9076,N_6409,N_7879);
or U9077 (N_9077,N_6521,N_7884);
or U9078 (N_9078,N_7929,N_7150);
nand U9079 (N_9079,N_6537,N_6200);
and U9080 (N_9080,N_7859,N_7572);
nor U9081 (N_9081,N_6316,N_6141);
nand U9082 (N_9082,N_7744,N_6062);
and U9083 (N_9083,N_7681,N_7624);
nor U9084 (N_9084,N_7787,N_6586);
and U9085 (N_9085,N_6967,N_7051);
and U9086 (N_9086,N_6855,N_7336);
nand U9087 (N_9087,N_6247,N_6184);
nor U9088 (N_9088,N_7006,N_7648);
nor U9089 (N_9089,N_7087,N_7332);
nor U9090 (N_9090,N_6402,N_7779);
nor U9091 (N_9091,N_7840,N_6053);
nand U9092 (N_9092,N_7342,N_7121);
nor U9093 (N_9093,N_6997,N_7050);
or U9094 (N_9094,N_6772,N_6703);
and U9095 (N_9095,N_7499,N_6365);
and U9096 (N_9096,N_7399,N_7613);
nand U9097 (N_9097,N_7889,N_7578);
and U9098 (N_9098,N_6415,N_6941);
nand U9099 (N_9099,N_7734,N_7417);
nand U9100 (N_9100,N_7506,N_6815);
nand U9101 (N_9101,N_6826,N_6732);
and U9102 (N_9102,N_6681,N_7246);
and U9103 (N_9103,N_7856,N_7373);
or U9104 (N_9104,N_6110,N_7984);
or U9105 (N_9105,N_6155,N_7667);
and U9106 (N_9106,N_6550,N_6936);
and U9107 (N_9107,N_6100,N_6171);
nor U9108 (N_9108,N_6311,N_6084);
nor U9109 (N_9109,N_7728,N_6032);
nand U9110 (N_9110,N_6274,N_7916);
or U9111 (N_9111,N_6264,N_6273);
or U9112 (N_9112,N_6042,N_7710);
nor U9113 (N_9113,N_7120,N_6833);
nor U9114 (N_9114,N_7626,N_7704);
nor U9115 (N_9115,N_7681,N_7193);
and U9116 (N_9116,N_6724,N_6953);
or U9117 (N_9117,N_7883,N_7419);
and U9118 (N_9118,N_6421,N_7881);
and U9119 (N_9119,N_6531,N_6865);
nand U9120 (N_9120,N_6538,N_7304);
nor U9121 (N_9121,N_6266,N_6260);
nor U9122 (N_9122,N_7432,N_6809);
and U9123 (N_9123,N_6632,N_6541);
nand U9124 (N_9124,N_7074,N_6857);
nand U9125 (N_9125,N_6041,N_6173);
nor U9126 (N_9126,N_6494,N_6630);
and U9127 (N_9127,N_7378,N_6552);
nor U9128 (N_9128,N_7222,N_6616);
nor U9129 (N_9129,N_6078,N_6516);
nor U9130 (N_9130,N_6595,N_6528);
and U9131 (N_9131,N_6036,N_7815);
and U9132 (N_9132,N_6038,N_6254);
and U9133 (N_9133,N_6270,N_6733);
and U9134 (N_9134,N_7025,N_6427);
and U9135 (N_9135,N_6002,N_6120);
nor U9136 (N_9136,N_7967,N_6114);
nand U9137 (N_9137,N_6238,N_7593);
nor U9138 (N_9138,N_7570,N_6231);
nand U9139 (N_9139,N_6578,N_7093);
or U9140 (N_9140,N_6219,N_6001);
nand U9141 (N_9141,N_7658,N_6697);
or U9142 (N_9142,N_6765,N_6209);
or U9143 (N_9143,N_6681,N_6579);
or U9144 (N_9144,N_7553,N_6927);
or U9145 (N_9145,N_7822,N_6276);
or U9146 (N_9146,N_6428,N_7915);
or U9147 (N_9147,N_6456,N_6814);
or U9148 (N_9148,N_6521,N_6647);
nor U9149 (N_9149,N_7383,N_7483);
nor U9150 (N_9150,N_7252,N_7068);
and U9151 (N_9151,N_6714,N_7339);
and U9152 (N_9152,N_7623,N_6374);
nor U9153 (N_9153,N_7862,N_7947);
nor U9154 (N_9154,N_6248,N_6650);
nand U9155 (N_9155,N_6933,N_6028);
nand U9156 (N_9156,N_6905,N_6426);
or U9157 (N_9157,N_6217,N_7230);
and U9158 (N_9158,N_7990,N_7602);
nand U9159 (N_9159,N_6870,N_7943);
nor U9160 (N_9160,N_6802,N_6973);
nand U9161 (N_9161,N_7906,N_6759);
nor U9162 (N_9162,N_6688,N_6149);
nor U9163 (N_9163,N_7455,N_6558);
and U9164 (N_9164,N_7910,N_6094);
nand U9165 (N_9165,N_7594,N_6405);
nor U9166 (N_9166,N_6288,N_6256);
and U9167 (N_9167,N_6244,N_7491);
or U9168 (N_9168,N_7735,N_6401);
nand U9169 (N_9169,N_7353,N_6199);
xor U9170 (N_9170,N_7554,N_6460);
nor U9171 (N_9171,N_6026,N_7096);
and U9172 (N_9172,N_7856,N_7383);
nand U9173 (N_9173,N_6507,N_7439);
and U9174 (N_9174,N_7412,N_7066);
nor U9175 (N_9175,N_6849,N_6434);
and U9176 (N_9176,N_6908,N_6938);
nand U9177 (N_9177,N_6669,N_6286);
nand U9178 (N_9178,N_7278,N_6331);
or U9179 (N_9179,N_7291,N_7840);
nand U9180 (N_9180,N_7878,N_7524);
or U9181 (N_9181,N_6346,N_7686);
nor U9182 (N_9182,N_6025,N_7815);
nor U9183 (N_9183,N_7593,N_7796);
and U9184 (N_9184,N_7601,N_6338);
nor U9185 (N_9185,N_6202,N_6740);
or U9186 (N_9186,N_7151,N_6899);
or U9187 (N_9187,N_6623,N_7437);
and U9188 (N_9188,N_6848,N_6436);
nor U9189 (N_9189,N_6464,N_6057);
or U9190 (N_9190,N_6029,N_6728);
nor U9191 (N_9191,N_7331,N_7051);
and U9192 (N_9192,N_7211,N_6819);
or U9193 (N_9193,N_6947,N_6615);
or U9194 (N_9194,N_6074,N_7792);
nor U9195 (N_9195,N_7785,N_6425);
nand U9196 (N_9196,N_6083,N_6026);
nand U9197 (N_9197,N_7979,N_6279);
or U9198 (N_9198,N_7974,N_6422);
nand U9199 (N_9199,N_7766,N_7474);
nand U9200 (N_9200,N_6875,N_6989);
and U9201 (N_9201,N_7655,N_6315);
nor U9202 (N_9202,N_7197,N_7809);
nor U9203 (N_9203,N_7906,N_7789);
and U9204 (N_9204,N_7736,N_7767);
and U9205 (N_9205,N_7699,N_7897);
and U9206 (N_9206,N_6782,N_6571);
and U9207 (N_9207,N_6642,N_7739);
nor U9208 (N_9208,N_7629,N_6323);
or U9209 (N_9209,N_7771,N_6688);
nor U9210 (N_9210,N_6464,N_6090);
nor U9211 (N_9211,N_6663,N_6711);
nor U9212 (N_9212,N_6844,N_6489);
nor U9213 (N_9213,N_6139,N_6558);
and U9214 (N_9214,N_6931,N_6481);
xor U9215 (N_9215,N_7786,N_6160);
and U9216 (N_9216,N_6551,N_6874);
nand U9217 (N_9217,N_7017,N_7675);
or U9218 (N_9218,N_7095,N_7958);
nor U9219 (N_9219,N_6254,N_7063);
nor U9220 (N_9220,N_6322,N_6913);
or U9221 (N_9221,N_7226,N_6005);
and U9222 (N_9222,N_7107,N_6187);
and U9223 (N_9223,N_7229,N_7396);
or U9224 (N_9224,N_6803,N_6239);
xnor U9225 (N_9225,N_6679,N_6845);
or U9226 (N_9226,N_7741,N_7410);
and U9227 (N_9227,N_7155,N_7299);
and U9228 (N_9228,N_6189,N_6056);
nor U9229 (N_9229,N_6553,N_7056);
nor U9230 (N_9230,N_6052,N_7286);
nand U9231 (N_9231,N_6183,N_6630);
nand U9232 (N_9232,N_6382,N_7994);
and U9233 (N_9233,N_7639,N_7456);
or U9234 (N_9234,N_6130,N_7606);
and U9235 (N_9235,N_6061,N_6404);
and U9236 (N_9236,N_7714,N_7945);
nand U9237 (N_9237,N_6980,N_6467);
nand U9238 (N_9238,N_7900,N_7775);
nand U9239 (N_9239,N_6054,N_7473);
or U9240 (N_9240,N_6797,N_7510);
nor U9241 (N_9241,N_6884,N_6766);
or U9242 (N_9242,N_6216,N_6300);
or U9243 (N_9243,N_7707,N_6679);
and U9244 (N_9244,N_7155,N_7929);
nor U9245 (N_9245,N_7316,N_6271);
or U9246 (N_9246,N_6749,N_7665);
nand U9247 (N_9247,N_6573,N_7931);
nor U9248 (N_9248,N_6116,N_6788);
or U9249 (N_9249,N_6618,N_7978);
nand U9250 (N_9250,N_6019,N_7201);
nor U9251 (N_9251,N_7553,N_6754);
nor U9252 (N_9252,N_6468,N_7290);
nand U9253 (N_9253,N_7572,N_6209);
or U9254 (N_9254,N_7344,N_7945);
or U9255 (N_9255,N_7394,N_7473);
nor U9256 (N_9256,N_7302,N_6734);
nand U9257 (N_9257,N_7724,N_7278);
nand U9258 (N_9258,N_6274,N_6904);
nor U9259 (N_9259,N_7040,N_7032);
or U9260 (N_9260,N_6820,N_6859);
nor U9261 (N_9261,N_6690,N_7215);
xor U9262 (N_9262,N_6912,N_7509);
and U9263 (N_9263,N_7020,N_6037);
nand U9264 (N_9264,N_7857,N_7869);
or U9265 (N_9265,N_7097,N_6598);
or U9266 (N_9266,N_6011,N_6461);
and U9267 (N_9267,N_7051,N_7321);
nand U9268 (N_9268,N_6532,N_6849);
nand U9269 (N_9269,N_6279,N_7190);
nand U9270 (N_9270,N_7984,N_6449);
nand U9271 (N_9271,N_6324,N_6890);
nor U9272 (N_9272,N_6418,N_7332);
nor U9273 (N_9273,N_7534,N_7454);
and U9274 (N_9274,N_6569,N_7708);
nor U9275 (N_9275,N_7952,N_6925);
nand U9276 (N_9276,N_6195,N_7863);
and U9277 (N_9277,N_7873,N_7797);
nor U9278 (N_9278,N_6919,N_6451);
or U9279 (N_9279,N_6662,N_7433);
and U9280 (N_9280,N_6117,N_6947);
and U9281 (N_9281,N_6828,N_7065);
nand U9282 (N_9282,N_7190,N_6763);
and U9283 (N_9283,N_6521,N_6311);
and U9284 (N_9284,N_7928,N_6318);
nand U9285 (N_9285,N_7569,N_7469);
nand U9286 (N_9286,N_6447,N_6346);
nand U9287 (N_9287,N_7412,N_7839);
and U9288 (N_9288,N_7647,N_7257);
nor U9289 (N_9289,N_7389,N_6856);
nor U9290 (N_9290,N_6530,N_7283);
and U9291 (N_9291,N_7458,N_6216);
or U9292 (N_9292,N_7537,N_7944);
xor U9293 (N_9293,N_7346,N_6307);
nor U9294 (N_9294,N_7218,N_6100);
nand U9295 (N_9295,N_7974,N_7416);
or U9296 (N_9296,N_7506,N_6420);
and U9297 (N_9297,N_7722,N_6991);
and U9298 (N_9298,N_7513,N_7654);
and U9299 (N_9299,N_6311,N_7796);
and U9300 (N_9300,N_6100,N_6831);
nand U9301 (N_9301,N_7889,N_7044);
and U9302 (N_9302,N_6161,N_7883);
nand U9303 (N_9303,N_7500,N_7551);
nand U9304 (N_9304,N_6905,N_7067);
and U9305 (N_9305,N_7986,N_6541);
and U9306 (N_9306,N_7990,N_7243);
nor U9307 (N_9307,N_7648,N_6681);
or U9308 (N_9308,N_7051,N_6088);
nand U9309 (N_9309,N_6561,N_7182);
nor U9310 (N_9310,N_6174,N_7594);
nand U9311 (N_9311,N_7596,N_7590);
and U9312 (N_9312,N_7309,N_6123);
or U9313 (N_9313,N_7711,N_7726);
nor U9314 (N_9314,N_7508,N_6684);
or U9315 (N_9315,N_7309,N_7544);
or U9316 (N_9316,N_7080,N_6758);
and U9317 (N_9317,N_7640,N_7595);
and U9318 (N_9318,N_7830,N_6726);
and U9319 (N_9319,N_6391,N_7665);
nor U9320 (N_9320,N_6779,N_6835);
and U9321 (N_9321,N_7994,N_6420);
nor U9322 (N_9322,N_7025,N_7408);
or U9323 (N_9323,N_7597,N_6901);
or U9324 (N_9324,N_7683,N_7752);
or U9325 (N_9325,N_6236,N_7133);
nand U9326 (N_9326,N_7372,N_7250);
and U9327 (N_9327,N_6366,N_7637);
nor U9328 (N_9328,N_6894,N_6760);
and U9329 (N_9329,N_6836,N_6006);
and U9330 (N_9330,N_7365,N_6267);
or U9331 (N_9331,N_7058,N_6001);
or U9332 (N_9332,N_6749,N_6816);
nand U9333 (N_9333,N_6845,N_7672);
or U9334 (N_9334,N_7906,N_7555);
or U9335 (N_9335,N_6840,N_7286);
nand U9336 (N_9336,N_6245,N_6478);
nand U9337 (N_9337,N_6307,N_6075);
nand U9338 (N_9338,N_7921,N_6935);
nor U9339 (N_9339,N_7150,N_6248);
or U9340 (N_9340,N_6544,N_7719);
or U9341 (N_9341,N_6065,N_7516);
nand U9342 (N_9342,N_7674,N_7166);
nand U9343 (N_9343,N_6559,N_7441);
nor U9344 (N_9344,N_6843,N_6400);
nand U9345 (N_9345,N_6473,N_6649);
nor U9346 (N_9346,N_6436,N_7492);
or U9347 (N_9347,N_6284,N_6801);
or U9348 (N_9348,N_7356,N_7779);
nand U9349 (N_9349,N_6974,N_7129);
nand U9350 (N_9350,N_6671,N_6874);
nor U9351 (N_9351,N_7426,N_6299);
or U9352 (N_9352,N_7727,N_6351);
nand U9353 (N_9353,N_6183,N_6078);
nor U9354 (N_9354,N_7837,N_7474);
nor U9355 (N_9355,N_6585,N_6027);
and U9356 (N_9356,N_6025,N_7245);
nand U9357 (N_9357,N_7041,N_7223);
nand U9358 (N_9358,N_7950,N_7209);
and U9359 (N_9359,N_6714,N_7338);
nand U9360 (N_9360,N_6569,N_7365);
and U9361 (N_9361,N_7859,N_6933);
nor U9362 (N_9362,N_6888,N_6889);
nand U9363 (N_9363,N_7420,N_6861);
nor U9364 (N_9364,N_7708,N_6120);
or U9365 (N_9365,N_7654,N_7972);
and U9366 (N_9366,N_7468,N_6324);
or U9367 (N_9367,N_6210,N_6951);
nor U9368 (N_9368,N_7932,N_7695);
or U9369 (N_9369,N_6238,N_6296);
or U9370 (N_9370,N_7698,N_7783);
nand U9371 (N_9371,N_6605,N_6388);
or U9372 (N_9372,N_6872,N_6572);
nor U9373 (N_9373,N_6487,N_6603);
or U9374 (N_9374,N_6537,N_6795);
and U9375 (N_9375,N_6132,N_7393);
or U9376 (N_9376,N_6358,N_7182);
and U9377 (N_9377,N_6742,N_6274);
or U9378 (N_9378,N_6539,N_7540);
nor U9379 (N_9379,N_6441,N_6859);
and U9380 (N_9380,N_7091,N_7113);
nor U9381 (N_9381,N_7870,N_6398);
nor U9382 (N_9382,N_6001,N_7512);
or U9383 (N_9383,N_7884,N_6313);
nor U9384 (N_9384,N_6256,N_6720);
or U9385 (N_9385,N_7296,N_7621);
nand U9386 (N_9386,N_7764,N_7007);
or U9387 (N_9387,N_6510,N_6528);
or U9388 (N_9388,N_6866,N_6082);
nor U9389 (N_9389,N_6717,N_6320);
nor U9390 (N_9390,N_6618,N_7690);
or U9391 (N_9391,N_7917,N_6316);
nand U9392 (N_9392,N_6269,N_6986);
and U9393 (N_9393,N_7235,N_6725);
nand U9394 (N_9394,N_6398,N_7812);
nand U9395 (N_9395,N_6351,N_6632);
and U9396 (N_9396,N_6706,N_7105);
xor U9397 (N_9397,N_6769,N_7479);
nor U9398 (N_9398,N_7007,N_6557);
xor U9399 (N_9399,N_6972,N_7101);
or U9400 (N_9400,N_7811,N_7365);
nand U9401 (N_9401,N_6503,N_6842);
and U9402 (N_9402,N_6950,N_7153);
or U9403 (N_9403,N_7586,N_6732);
nand U9404 (N_9404,N_6943,N_7348);
and U9405 (N_9405,N_6258,N_7582);
nand U9406 (N_9406,N_7667,N_6442);
and U9407 (N_9407,N_6576,N_6193);
nand U9408 (N_9408,N_7776,N_7667);
or U9409 (N_9409,N_6536,N_6702);
and U9410 (N_9410,N_7903,N_6949);
and U9411 (N_9411,N_6522,N_6872);
nand U9412 (N_9412,N_6109,N_6916);
nor U9413 (N_9413,N_6907,N_6104);
nor U9414 (N_9414,N_7283,N_6166);
or U9415 (N_9415,N_7872,N_7167);
or U9416 (N_9416,N_7805,N_6898);
and U9417 (N_9417,N_7584,N_7555);
nor U9418 (N_9418,N_7346,N_6479);
nand U9419 (N_9419,N_6981,N_7365);
nand U9420 (N_9420,N_7682,N_7164);
and U9421 (N_9421,N_6750,N_6087);
or U9422 (N_9422,N_7480,N_7868);
and U9423 (N_9423,N_6052,N_7970);
nand U9424 (N_9424,N_6123,N_7005);
or U9425 (N_9425,N_7378,N_7520);
nor U9426 (N_9426,N_6799,N_7696);
and U9427 (N_9427,N_7741,N_7823);
nand U9428 (N_9428,N_7719,N_7214);
nor U9429 (N_9429,N_6448,N_6780);
nand U9430 (N_9430,N_6741,N_6025);
nor U9431 (N_9431,N_7100,N_7070);
or U9432 (N_9432,N_7372,N_6467);
or U9433 (N_9433,N_6168,N_6576);
nand U9434 (N_9434,N_6634,N_6832);
nand U9435 (N_9435,N_6796,N_6387);
nor U9436 (N_9436,N_6738,N_7502);
nor U9437 (N_9437,N_7932,N_6199);
and U9438 (N_9438,N_6112,N_7659);
nor U9439 (N_9439,N_6553,N_6408);
nor U9440 (N_9440,N_7789,N_6447);
or U9441 (N_9441,N_6864,N_6992);
xor U9442 (N_9442,N_6925,N_6004);
and U9443 (N_9443,N_6952,N_7009);
nand U9444 (N_9444,N_6549,N_6269);
or U9445 (N_9445,N_6408,N_6593);
or U9446 (N_9446,N_7289,N_6523);
or U9447 (N_9447,N_6081,N_7720);
and U9448 (N_9448,N_7382,N_7443);
nand U9449 (N_9449,N_7278,N_7080);
or U9450 (N_9450,N_7892,N_6236);
or U9451 (N_9451,N_6300,N_6742);
or U9452 (N_9452,N_6900,N_7911);
nand U9453 (N_9453,N_7835,N_7414);
nor U9454 (N_9454,N_6438,N_6679);
or U9455 (N_9455,N_7170,N_7928);
nand U9456 (N_9456,N_6897,N_6245);
and U9457 (N_9457,N_7668,N_6881);
and U9458 (N_9458,N_7824,N_7247);
nand U9459 (N_9459,N_7917,N_7837);
and U9460 (N_9460,N_7857,N_6106);
and U9461 (N_9461,N_7960,N_7633);
nand U9462 (N_9462,N_7775,N_6623);
and U9463 (N_9463,N_6808,N_7711);
or U9464 (N_9464,N_7637,N_6654);
and U9465 (N_9465,N_7594,N_7491);
nor U9466 (N_9466,N_7151,N_7892);
or U9467 (N_9467,N_6312,N_6374);
or U9468 (N_9468,N_7717,N_7454);
nor U9469 (N_9469,N_6345,N_7785);
and U9470 (N_9470,N_6619,N_7582);
nand U9471 (N_9471,N_7176,N_6039);
or U9472 (N_9472,N_7118,N_6260);
and U9473 (N_9473,N_7415,N_7300);
and U9474 (N_9474,N_6743,N_7209);
or U9475 (N_9475,N_7716,N_6635);
and U9476 (N_9476,N_7527,N_6350);
nand U9477 (N_9477,N_7487,N_7411);
and U9478 (N_9478,N_6537,N_6530);
nand U9479 (N_9479,N_7389,N_7349);
nor U9480 (N_9480,N_6022,N_7853);
or U9481 (N_9481,N_6548,N_6049);
or U9482 (N_9482,N_6078,N_6004);
or U9483 (N_9483,N_7195,N_7025);
and U9484 (N_9484,N_6960,N_7242);
nand U9485 (N_9485,N_6156,N_6710);
nand U9486 (N_9486,N_6898,N_6536);
or U9487 (N_9487,N_6166,N_6736);
xnor U9488 (N_9488,N_7251,N_7461);
nor U9489 (N_9489,N_7949,N_6449);
and U9490 (N_9490,N_6452,N_6373);
nand U9491 (N_9491,N_7878,N_6032);
or U9492 (N_9492,N_6727,N_6954);
and U9493 (N_9493,N_6177,N_7092);
nor U9494 (N_9494,N_7143,N_6338);
nor U9495 (N_9495,N_7131,N_7368);
or U9496 (N_9496,N_6542,N_7408);
or U9497 (N_9497,N_7511,N_6031);
nand U9498 (N_9498,N_7307,N_6160);
or U9499 (N_9499,N_6677,N_6863);
nor U9500 (N_9500,N_7294,N_7034);
nor U9501 (N_9501,N_7951,N_7199);
and U9502 (N_9502,N_7190,N_7734);
nor U9503 (N_9503,N_6249,N_7277);
and U9504 (N_9504,N_6883,N_7463);
and U9505 (N_9505,N_7998,N_7208);
and U9506 (N_9506,N_7482,N_7172);
and U9507 (N_9507,N_6310,N_7151);
and U9508 (N_9508,N_7668,N_6479);
and U9509 (N_9509,N_7007,N_7971);
nor U9510 (N_9510,N_6637,N_7980);
or U9511 (N_9511,N_6493,N_7901);
nor U9512 (N_9512,N_6486,N_6530);
nor U9513 (N_9513,N_6962,N_6268);
or U9514 (N_9514,N_6604,N_6284);
nand U9515 (N_9515,N_6177,N_7337);
or U9516 (N_9516,N_6977,N_7696);
nand U9517 (N_9517,N_6886,N_6066);
nor U9518 (N_9518,N_6531,N_7580);
and U9519 (N_9519,N_6020,N_7001);
nand U9520 (N_9520,N_7029,N_6032);
or U9521 (N_9521,N_7656,N_7082);
nand U9522 (N_9522,N_7268,N_7500);
and U9523 (N_9523,N_7063,N_6243);
nor U9524 (N_9524,N_6732,N_6372);
nand U9525 (N_9525,N_7386,N_6355);
or U9526 (N_9526,N_7658,N_7606);
nand U9527 (N_9527,N_7434,N_7779);
nand U9528 (N_9528,N_7989,N_7065);
nor U9529 (N_9529,N_6967,N_7646);
or U9530 (N_9530,N_6323,N_7733);
and U9531 (N_9531,N_6265,N_6684);
and U9532 (N_9532,N_7711,N_7840);
nor U9533 (N_9533,N_6646,N_7014);
or U9534 (N_9534,N_6323,N_6462);
nand U9535 (N_9535,N_7694,N_7127);
and U9536 (N_9536,N_7456,N_6817);
nand U9537 (N_9537,N_7305,N_6013);
or U9538 (N_9538,N_6937,N_7073);
or U9539 (N_9539,N_7542,N_6613);
or U9540 (N_9540,N_7666,N_6535);
nor U9541 (N_9541,N_7299,N_6842);
and U9542 (N_9542,N_7418,N_6502);
nor U9543 (N_9543,N_6077,N_6787);
or U9544 (N_9544,N_6902,N_6075);
or U9545 (N_9545,N_6756,N_7607);
nand U9546 (N_9546,N_6084,N_7162);
or U9547 (N_9547,N_7824,N_7875);
or U9548 (N_9548,N_7778,N_6214);
and U9549 (N_9549,N_7651,N_6308);
and U9550 (N_9550,N_6109,N_7479);
nand U9551 (N_9551,N_7601,N_6477);
nand U9552 (N_9552,N_6741,N_7221);
and U9553 (N_9553,N_6357,N_6880);
nor U9554 (N_9554,N_7384,N_7036);
or U9555 (N_9555,N_7164,N_6884);
and U9556 (N_9556,N_6725,N_7373);
and U9557 (N_9557,N_6313,N_6361);
or U9558 (N_9558,N_7140,N_7754);
nand U9559 (N_9559,N_6185,N_6051);
nor U9560 (N_9560,N_7989,N_6550);
nor U9561 (N_9561,N_7849,N_6185);
nand U9562 (N_9562,N_6417,N_6582);
nand U9563 (N_9563,N_6768,N_7635);
and U9564 (N_9564,N_7639,N_7304);
or U9565 (N_9565,N_6910,N_7867);
or U9566 (N_9566,N_6022,N_6292);
and U9567 (N_9567,N_7667,N_7424);
nor U9568 (N_9568,N_7262,N_6408);
nand U9569 (N_9569,N_7727,N_7153);
or U9570 (N_9570,N_7930,N_7001);
nor U9571 (N_9571,N_7085,N_7228);
nand U9572 (N_9572,N_6740,N_7127);
and U9573 (N_9573,N_7644,N_6717);
nor U9574 (N_9574,N_7011,N_6698);
nand U9575 (N_9575,N_7752,N_7810);
nand U9576 (N_9576,N_7875,N_7696);
and U9577 (N_9577,N_7236,N_7099);
nor U9578 (N_9578,N_7461,N_6626);
nand U9579 (N_9579,N_6625,N_7161);
nor U9580 (N_9580,N_7611,N_6969);
nor U9581 (N_9581,N_7909,N_6281);
or U9582 (N_9582,N_7446,N_7154);
and U9583 (N_9583,N_6523,N_6435);
or U9584 (N_9584,N_6368,N_6473);
or U9585 (N_9585,N_6905,N_6403);
nor U9586 (N_9586,N_7238,N_6601);
and U9587 (N_9587,N_7792,N_7089);
nor U9588 (N_9588,N_7808,N_7925);
nand U9589 (N_9589,N_7188,N_7051);
or U9590 (N_9590,N_7971,N_6169);
nand U9591 (N_9591,N_6678,N_7288);
or U9592 (N_9592,N_6348,N_6382);
nor U9593 (N_9593,N_6551,N_7477);
and U9594 (N_9594,N_6380,N_7061);
and U9595 (N_9595,N_6642,N_6578);
nand U9596 (N_9596,N_6256,N_6998);
or U9597 (N_9597,N_6187,N_6557);
nand U9598 (N_9598,N_7700,N_7848);
or U9599 (N_9599,N_6482,N_6275);
and U9600 (N_9600,N_6312,N_7968);
xor U9601 (N_9601,N_6589,N_6559);
nand U9602 (N_9602,N_7278,N_6282);
and U9603 (N_9603,N_7582,N_7203);
and U9604 (N_9604,N_7846,N_7870);
or U9605 (N_9605,N_7229,N_7464);
xor U9606 (N_9606,N_7135,N_7786);
or U9607 (N_9607,N_6588,N_6566);
nand U9608 (N_9608,N_6288,N_6917);
nand U9609 (N_9609,N_6579,N_6797);
nor U9610 (N_9610,N_6614,N_6132);
nor U9611 (N_9611,N_7996,N_6146);
or U9612 (N_9612,N_7827,N_6381);
or U9613 (N_9613,N_6809,N_6985);
and U9614 (N_9614,N_7784,N_6241);
or U9615 (N_9615,N_6609,N_6497);
or U9616 (N_9616,N_6674,N_7530);
and U9617 (N_9617,N_7363,N_6299);
or U9618 (N_9618,N_7789,N_6620);
nand U9619 (N_9619,N_7394,N_6240);
or U9620 (N_9620,N_7512,N_7203);
nor U9621 (N_9621,N_6357,N_7447);
nor U9622 (N_9622,N_7736,N_7983);
and U9623 (N_9623,N_7236,N_6664);
nand U9624 (N_9624,N_6027,N_6508);
or U9625 (N_9625,N_7941,N_7108);
nor U9626 (N_9626,N_6775,N_7976);
nand U9627 (N_9627,N_7857,N_6737);
nand U9628 (N_9628,N_7259,N_7933);
or U9629 (N_9629,N_6892,N_6965);
nand U9630 (N_9630,N_7002,N_6486);
xor U9631 (N_9631,N_7913,N_7529);
nand U9632 (N_9632,N_7674,N_6631);
nor U9633 (N_9633,N_6856,N_7758);
nor U9634 (N_9634,N_6389,N_7400);
nor U9635 (N_9635,N_6072,N_6921);
nand U9636 (N_9636,N_6904,N_6471);
or U9637 (N_9637,N_7953,N_7727);
and U9638 (N_9638,N_7905,N_6988);
nor U9639 (N_9639,N_6284,N_6545);
nor U9640 (N_9640,N_7415,N_6130);
nor U9641 (N_9641,N_6511,N_7120);
or U9642 (N_9642,N_6986,N_6510);
and U9643 (N_9643,N_6856,N_7842);
nand U9644 (N_9644,N_6302,N_7583);
and U9645 (N_9645,N_7546,N_6365);
nand U9646 (N_9646,N_6858,N_7008);
and U9647 (N_9647,N_6499,N_6214);
and U9648 (N_9648,N_7730,N_7634);
and U9649 (N_9649,N_6585,N_6698);
nand U9650 (N_9650,N_7822,N_7221);
nor U9651 (N_9651,N_6839,N_6897);
or U9652 (N_9652,N_7171,N_7947);
or U9653 (N_9653,N_6523,N_7676);
or U9654 (N_9654,N_6803,N_6664);
nor U9655 (N_9655,N_7583,N_6145);
or U9656 (N_9656,N_6473,N_6133);
nand U9657 (N_9657,N_6646,N_7084);
and U9658 (N_9658,N_6179,N_6799);
nand U9659 (N_9659,N_7672,N_6661);
or U9660 (N_9660,N_7009,N_6437);
and U9661 (N_9661,N_7332,N_6265);
nor U9662 (N_9662,N_6468,N_6489);
and U9663 (N_9663,N_7474,N_7640);
or U9664 (N_9664,N_6063,N_6067);
nand U9665 (N_9665,N_7403,N_6324);
or U9666 (N_9666,N_6464,N_6270);
and U9667 (N_9667,N_6477,N_7077);
and U9668 (N_9668,N_7504,N_7828);
nand U9669 (N_9669,N_6629,N_7547);
and U9670 (N_9670,N_7256,N_7464);
nand U9671 (N_9671,N_7892,N_7152);
nand U9672 (N_9672,N_6211,N_7660);
and U9673 (N_9673,N_6192,N_7426);
and U9674 (N_9674,N_7713,N_7556);
or U9675 (N_9675,N_6504,N_6776);
and U9676 (N_9676,N_6644,N_7578);
nor U9677 (N_9677,N_6504,N_7066);
nor U9678 (N_9678,N_7784,N_7410);
nor U9679 (N_9679,N_6042,N_7746);
nand U9680 (N_9680,N_7655,N_7002);
or U9681 (N_9681,N_6700,N_6109);
nand U9682 (N_9682,N_6205,N_7203);
or U9683 (N_9683,N_7074,N_6191);
and U9684 (N_9684,N_7511,N_7715);
nor U9685 (N_9685,N_6952,N_6876);
or U9686 (N_9686,N_6892,N_7018);
nand U9687 (N_9687,N_7763,N_7679);
and U9688 (N_9688,N_7184,N_6413);
nand U9689 (N_9689,N_7858,N_6273);
nand U9690 (N_9690,N_6729,N_6855);
and U9691 (N_9691,N_7154,N_7522);
or U9692 (N_9692,N_7866,N_6500);
nor U9693 (N_9693,N_7986,N_7744);
nand U9694 (N_9694,N_6651,N_6846);
nand U9695 (N_9695,N_6557,N_6788);
or U9696 (N_9696,N_7033,N_7229);
nand U9697 (N_9697,N_6911,N_6199);
nand U9698 (N_9698,N_7903,N_7516);
and U9699 (N_9699,N_6163,N_6993);
or U9700 (N_9700,N_7242,N_7065);
and U9701 (N_9701,N_6457,N_6570);
and U9702 (N_9702,N_6835,N_7475);
nor U9703 (N_9703,N_7989,N_6756);
nor U9704 (N_9704,N_7062,N_6762);
or U9705 (N_9705,N_7066,N_6362);
and U9706 (N_9706,N_7638,N_7136);
or U9707 (N_9707,N_6708,N_7681);
or U9708 (N_9708,N_7566,N_6345);
nand U9709 (N_9709,N_6581,N_6544);
nand U9710 (N_9710,N_7458,N_7367);
nand U9711 (N_9711,N_7903,N_6749);
or U9712 (N_9712,N_6159,N_6968);
and U9713 (N_9713,N_6854,N_6075);
nand U9714 (N_9714,N_6887,N_6460);
or U9715 (N_9715,N_7114,N_7550);
or U9716 (N_9716,N_7091,N_6271);
nor U9717 (N_9717,N_6115,N_7299);
or U9718 (N_9718,N_6201,N_6192);
nand U9719 (N_9719,N_7931,N_6000);
or U9720 (N_9720,N_7598,N_6515);
nand U9721 (N_9721,N_7463,N_6619);
nand U9722 (N_9722,N_7793,N_7698);
or U9723 (N_9723,N_7602,N_7757);
and U9724 (N_9724,N_7057,N_7890);
nor U9725 (N_9725,N_6213,N_7443);
nor U9726 (N_9726,N_7363,N_6826);
and U9727 (N_9727,N_6383,N_7380);
and U9728 (N_9728,N_6043,N_7451);
nor U9729 (N_9729,N_7126,N_7253);
or U9730 (N_9730,N_7957,N_7593);
or U9731 (N_9731,N_7348,N_6363);
and U9732 (N_9732,N_7594,N_6952);
and U9733 (N_9733,N_6318,N_6161);
nand U9734 (N_9734,N_6128,N_7474);
nand U9735 (N_9735,N_7167,N_7289);
or U9736 (N_9736,N_6293,N_7691);
and U9737 (N_9737,N_7633,N_7654);
or U9738 (N_9738,N_7309,N_6627);
nor U9739 (N_9739,N_6921,N_7724);
and U9740 (N_9740,N_6496,N_6397);
xor U9741 (N_9741,N_6573,N_7464);
and U9742 (N_9742,N_7650,N_6909);
nand U9743 (N_9743,N_6966,N_6693);
or U9744 (N_9744,N_7654,N_7268);
nand U9745 (N_9745,N_6645,N_6194);
or U9746 (N_9746,N_7535,N_6630);
nand U9747 (N_9747,N_6406,N_7333);
nor U9748 (N_9748,N_6560,N_7551);
nand U9749 (N_9749,N_7254,N_6204);
nor U9750 (N_9750,N_7870,N_7686);
or U9751 (N_9751,N_6258,N_6421);
or U9752 (N_9752,N_7035,N_7528);
nand U9753 (N_9753,N_6571,N_6217);
nor U9754 (N_9754,N_6863,N_6346);
and U9755 (N_9755,N_7928,N_7826);
or U9756 (N_9756,N_7866,N_7075);
nor U9757 (N_9757,N_7036,N_7344);
xnor U9758 (N_9758,N_6976,N_7784);
nand U9759 (N_9759,N_6234,N_6355);
xor U9760 (N_9760,N_7774,N_7886);
nand U9761 (N_9761,N_7564,N_6629);
and U9762 (N_9762,N_7253,N_7171);
nor U9763 (N_9763,N_7688,N_6739);
nor U9764 (N_9764,N_7423,N_6737);
nand U9765 (N_9765,N_7098,N_7740);
and U9766 (N_9766,N_6934,N_7707);
nand U9767 (N_9767,N_7183,N_6473);
nand U9768 (N_9768,N_6482,N_6974);
nand U9769 (N_9769,N_7929,N_6908);
nand U9770 (N_9770,N_7206,N_6657);
nand U9771 (N_9771,N_7335,N_7689);
nand U9772 (N_9772,N_6563,N_7053);
and U9773 (N_9773,N_7555,N_7728);
nor U9774 (N_9774,N_7201,N_7640);
nor U9775 (N_9775,N_7950,N_6511);
nor U9776 (N_9776,N_7347,N_7022);
nand U9777 (N_9777,N_6848,N_7098);
nand U9778 (N_9778,N_6432,N_7973);
nand U9779 (N_9779,N_6386,N_6566);
nand U9780 (N_9780,N_7586,N_7445);
or U9781 (N_9781,N_6304,N_7718);
nor U9782 (N_9782,N_6685,N_7445);
or U9783 (N_9783,N_6996,N_6050);
or U9784 (N_9784,N_6076,N_6625);
nand U9785 (N_9785,N_7389,N_7461);
or U9786 (N_9786,N_6642,N_6577);
nand U9787 (N_9787,N_6935,N_7413);
and U9788 (N_9788,N_6019,N_6000);
nand U9789 (N_9789,N_6230,N_7490);
nor U9790 (N_9790,N_6082,N_7803);
and U9791 (N_9791,N_7802,N_7249);
nand U9792 (N_9792,N_7121,N_7168);
nor U9793 (N_9793,N_7806,N_7047);
xnor U9794 (N_9794,N_7635,N_6422);
or U9795 (N_9795,N_6302,N_7671);
nor U9796 (N_9796,N_6940,N_7558);
or U9797 (N_9797,N_6899,N_7047);
or U9798 (N_9798,N_6355,N_7025);
nor U9799 (N_9799,N_7459,N_7596);
nand U9800 (N_9800,N_7259,N_7986);
nand U9801 (N_9801,N_6750,N_7887);
nand U9802 (N_9802,N_7854,N_7532);
nor U9803 (N_9803,N_7776,N_6310);
nand U9804 (N_9804,N_7036,N_6693);
nand U9805 (N_9805,N_7876,N_6287);
nand U9806 (N_9806,N_6012,N_7891);
xor U9807 (N_9807,N_7954,N_7764);
nor U9808 (N_9808,N_7343,N_7895);
or U9809 (N_9809,N_6396,N_7609);
nor U9810 (N_9810,N_6656,N_6773);
and U9811 (N_9811,N_6081,N_7964);
and U9812 (N_9812,N_7603,N_7818);
or U9813 (N_9813,N_7339,N_7331);
nor U9814 (N_9814,N_6389,N_6986);
or U9815 (N_9815,N_6410,N_7269);
or U9816 (N_9816,N_7017,N_6750);
nand U9817 (N_9817,N_7787,N_6339);
nand U9818 (N_9818,N_7064,N_7347);
and U9819 (N_9819,N_6662,N_7966);
nor U9820 (N_9820,N_7846,N_6088);
nor U9821 (N_9821,N_6785,N_6136);
and U9822 (N_9822,N_6540,N_6422);
nand U9823 (N_9823,N_7697,N_7736);
nor U9824 (N_9824,N_6052,N_6862);
nand U9825 (N_9825,N_6493,N_6333);
and U9826 (N_9826,N_7292,N_6992);
nand U9827 (N_9827,N_7298,N_7561);
nand U9828 (N_9828,N_7399,N_7731);
and U9829 (N_9829,N_6865,N_7634);
nor U9830 (N_9830,N_6904,N_6285);
nand U9831 (N_9831,N_6088,N_7670);
or U9832 (N_9832,N_7036,N_6555);
nor U9833 (N_9833,N_7803,N_6188);
nor U9834 (N_9834,N_6777,N_6813);
and U9835 (N_9835,N_7385,N_6199);
nand U9836 (N_9836,N_7358,N_6389);
nand U9837 (N_9837,N_6788,N_6328);
or U9838 (N_9838,N_7490,N_6245);
or U9839 (N_9839,N_7765,N_6278);
and U9840 (N_9840,N_6312,N_6974);
and U9841 (N_9841,N_7794,N_6221);
nor U9842 (N_9842,N_6641,N_7482);
nor U9843 (N_9843,N_7625,N_7227);
or U9844 (N_9844,N_6847,N_7495);
and U9845 (N_9845,N_6975,N_6801);
and U9846 (N_9846,N_7376,N_7647);
or U9847 (N_9847,N_6838,N_6102);
or U9848 (N_9848,N_7720,N_7893);
nand U9849 (N_9849,N_7456,N_7532);
nor U9850 (N_9850,N_7725,N_6909);
nor U9851 (N_9851,N_7596,N_6518);
or U9852 (N_9852,N_6578,N_7899);
or U9853 (N_9853,N_6164,N_7583);
nand U9854 (N_9854,N_7562,N_7571);
nor U9855 (N_9855,N_6924,N_6024);
and U9856 (N_9856,N_6156,N_6875);
nand U9857 (N_9857,N_6253,N_7179);
or U9858 (N_9858,N_6233,N_7748);
nor U9859 (N_9859,N_6331,N_7846);
or U9860 (N_9860,N_6064,N_6975);
or U9861 (N_9861,N_7331,N_7020);
and U9862 (N_9862,N_7829,N_6249);
nor U9863 (N_9863,N_6434,N_6842);
nor U9864 (N_9864,N_6391,N_6732);
or U9865 (N_9865,N_7177,N_6876);
and U9866 (N_9866,N_6761,N_6465);
and U9867 (N_9867,N_7324,N_7027);
or U9868 (N_9868,N_7492,N_7024);
nor U9869 (N_9869,N_6026,N_6513);
or U9870 (N_9870,N_6834,N_7746);
nand U9871 (N_9871,N_7577,N_6711);
and U9872 (N_9872,N_7561,N_7751);
nand U9873 (N_9873,N_6031,N_7980);
or U9874 (N_9874,N_7417,N_6766);
nand U9875 (N_9875,N_7747,N_7529);
nor U9876 (N_9876,N_6191,N_7843);
nor U9877 (N_9877,N_7121,N_6369);
or U9878 (N_9878,N_6302,N_6911);
nor U9879 (N_9879,N_7549,N_6902);
and U9880 (N_9880,N_7633,N_6995);
or U9881 (N_9881,N_7002,N_7322);
nor U9882 (N_9882,N_6594,N_7432);
and U9883 (N_9883,N_7275,N_6282);
or U9884 (N_9884,N_7322,N_7226);
or U9885 (N_9885,N_7645,N_6923);
xnor U9886 (N_9886,N_7909,N_7634);
nor U9887 (N_9887,N_6342,N_6773);
or U9888 (N_9888,N_6311,N_7213);
or U9889 (N_9889,N_7506,N_6516);
nand U9890 (N_9890,N_7491,N_7575);
and U9891 (N_9891,N_6881,N_6449);
nor U9892 (N_9892,N_6322,N_6714);
nor U9893 (N_9893,N_7698,N_7878);
nor U9894 (N_9894,N_6549,N_6645);
nand U9895 (N_9895,N_6111,N_7518);
or U9896 (N_9896,N_7676,N_7553);
or U9897 (N_9897,N_6071,N_7813);
nor U9898 (N_9898,N_7690,N_6291);
nor U9899 (N_9899,N_7837,N_7304);
and U9900 (N_9900,N_7646,N_7593);
nand U9901 (N_9901,N_6252,N_6871);
and U9902 (N_9902,N_6398,N_7720);
and U9903 (N_9903,N_7653,N_6795);
or U9904 (N_9904,N_7153,N_6806);
or U9905 (N_9905,N_7296,N_6132);
nand U9906 (N_9906,N_7160,N_7810);
or U9907 (N_9907,N_7796,N_6163);
nand U9908 (N_9908,N_7137,N_7920);
nand U9909 (N_9909,N_7219,N_6475);
nand U9910 (N_9910,N_7267,N_7322);
and U9911 (N_9911,N_7007,N_6114);
nand U9912 (N_9912,N_7782,N_6011);
nor U9913 (N_9913,N_6617,N_7278);
nand U9914 (N_9914,N_6357,N_6250);
and U9915 (N_9915,N_7694,N_7071);
or U9916 (N_9916,N_6199,N_6219);
nor U9917 (N_9917,N_6518,N_6825);
and U9918 (N_9918,N_6877,N_7601);
or U9919 (N_9919,N_7199,N_7786);
nand U9920 (N_9920,N_7321,N_7491);
or U9921 (N_9921,N_7886,N_6806);
nand U9922 (N_9922,N_7436,N_6766);
and U9923 (N_9923,N_6377,N_6197);
and U9924 (N_9924,N_6916,N_7385);
nor U9925 (N_9925,N_6236,N_6429);
xor U9926 (N_9926,N_7251,N_6987);
or U9927 (N_9927,N_7579,N_7580);
nand U9928 (N_9928,N_7829,N_6410);
xor U9929 (N_9929,N_6798,N_6271);
nor U9930 (N_9930,N_7506,N_6838);
or U9931 (N_9931,N_7313,N_7138);
and U9932 (N_9932,N_7213,N_7103);
or U9933 (N_9933,N_6546,N_7815);
nor U9934 (N_9934,N_6693,N_6892);
nor U9935 (N_9935,N_6414,N_6615);
nor U9936 (N_9936,N_6264,N_7384);
and U9937 (N_9937,N_6644,N_6439);
nand U9938 (N_9938,N_7007,N_7863);
or U9939 (N_9939,N_6793,N_6968);
and U9940 (N_9940,N_6814,N_7710);
or U9941 (N_9941,N_7742,N_6034);
nor U9942 (N_9942,N_7141,N_7583);
nand U9943 (N_9943,N_7273,N_7926);
or U9944 (N_9944,N_6054,N_6228);
nor U9945 (N_9945,N_7116,N_7372);
nor U9946 (N_9946,N_6624,N_6754);
and U9947 (N_9947,N_6571,N_7484);
or U9948 (N_9948,N_6208,N_6376);
nor U9949 (N_9949,N_6083,N_7051);
or U9950 (N_9950,N_7017,N_7562);
nor U9951 (N_9951,N_7567,N_6078);
or U9952 (N_9952,N_6634,N_6813);
nor U9953 (N_9953,N_7797,N_7456);
nor U9954 (N_9954,N_6645,N_6530);
or U9955 (N_9955,N_6843,N_7670);
and U9956 (N_9956,N_6673,N_7608);
or U9957 (N_9957,N_6876,N_7196);
nand U9958 (N_9958,N_7267,N_6508);
nor U9959 (N_9959,N_7108,N_6495);
and U9960 (N_9960,N_6719,N_7254);
and U9961 (N_9961,N_7601,N_6939);
nor U9962 (N_9962,N_7250,N_6971);
and U9963 (N_9963,N_7274,N_7134);
or U9964 (N_9964,N_6814,N_7863);
nor U9965 (N_9965,N_7295,N_7187);
nor U9966 (N_9966,N_6565,N_7566);
or U9967 (N_9967,N_7383,N_6506);
nor U9968 (N_9968,N_7513,N_7665);
and U9969 (N_9969,N_6261,N_7951);
or U9970 (N_9970,N_6260,N_6342);
nor U9971 (N_9971,N_6107,N_6207);
and U9972 (N_9972,N_7219,N_6178);
or U9973 (N_9973,N_6534,N_7908);
and U9974 (N_9974,N_7027,N_7010);
and U9975 (N_9975,N_6668,N_6158);
and U9976 (N_9976,N_7168,N_7587);
nor U9977 (N_9977,N_6927,N_6996);
nor U9978 (N_9978,N_7281,N_6550);
or U9979 (N_9979,N_6522,N_6842);
and U9980 (N_9980,N_7924,N_6519);
nor U9981 (N_9981,N_7669,N_7547);
nand U9982 (N_9982,N_7536,N_7408);
and U9983 (N_9983,N_7575,N_6721);
nor U9984 (N_9984,N_6332,N_6358);
nand U9985 (N_9985,N_7909,N_6807);
nand U9986 (N_9986,N_6496,N_6373);
or U9987 (N_9987,N_7411,N_6254);
nor U9988 (N_9988,N_7295,N_7994);
xor U9989 (N_9989,N_7516,N_7201);
nor U9990 (N_9990,N_7323,N_6602);
or U9991 (N_9991,N_7150,N_6650);
or U9992 (N_9992,N_7229,N_6480);
xnor U9993 (N_9993,N_7124,N_7500);
or U9994 (N_9994,N_6274,N_7383);
or U9995 (N_9995,N_6264,N_6131);
nand U9996 (N_9996,N_6982,N_6682);
nor U9997 (N_9997,N_6052,N_7938);
nand U9998 (N_9998,N_7760,N_6951);
nor U9999 (N_9999,N_7438,N_7357);
xor U10000 (N_10000,N_9296,N_8291);
or U10001 (N_10001,N_8039,N_9607);
xnor U10002 (N_10002,N_9843,N_8565);
nor U10003 (N_10003,N_9897,N_9026);
nor U10004 (N_10004,N_9679,N_9173);
and U10005 (N_10005,N_8958,N_9440);
or U10006 (N_10006,N_8763,N_9832);
nand U10007 (N_10007,N_8793,N_9284);
nor U10008 (N_10008,N_9108,N_8718);
nor U10009 (N_10009,N_9677,N_9184);
nand U10010 (N_10010,N_9378,N_8824);
nor U10011 (N_10011,N_8308,N_9071);
and U10012 (N_10012,N_9760,N_9011);
or U10013 (N_10013,N_9165,N_8767);
or U10014 (N_10014,N_9403,N_8697);
nor U10015 (N_10015,N_8783,N_9512);
or U10016 (N_10016,N_9972,N_8096);
xor U10017 (N_10017,N_9935,N_8484);
or U10018 (N_10018,N_9393,N_8517);
nand U10019 (N_10019,N_8092,N_9475);
or U10020 (N_10020,N_9926,N_8263);
nor U10021 (N_10021,N_8908,N_9106);
nor U10022 (N_10022,N_9045,N_8315);
or U10023 (N_10023,N_8837,N_9836);
nor U10024 (N_10024,N_9453,N_9626);
nor U10025 (N_10025,N_8847,N_8164);
and U10026 (N_10026,N_9616,N_8500);
nor U10027 (N_10027,N_9846,N_8018);
nor U10028 (N_10028,N_9124,N_8639);
nor U10029 (N_10029,N_8266,N_9156);
nor U10030 (N_10030,N_8220,N_9375);
and U10031 (N_10031,N_9894,N_8141);
nor U10032 (N_10032,N_9931,N_8705);
nand U10033 (N_10033,N_9536,N_9898);
nor U10034 (N_10034,N_9125,N_8654);
or U10035 (N_10035,N_9492,N_9458);
nor U10036 (N_10036,N_9606,N_9987);
nor U10037 (N_10037,N_8350,N_9645);
nand U10038 (N_10038,N_8117,N_8632);
and U10039 (N_10039,N_8085,N_9338);
and U10040 (N_10040,N_8582,N_9650);
and U10041 (N_10041,N_8979,N_8984);
xnor U10042 (N_10042,N_8306,N_8228);
and U10043 (N_10043,N_9706,N_9831);
and U10044 (N_10044,N_8459,N_9759);
nor U10045 (N_10045,N_9945,N_8066);
and U10046 (N_10046,N_9300,N_8712);
or U10047 (N_10047,N_9291,N_8177);
nand U10048 (N_10048,N_9849,N_9752);
nand U10049 (N_10049,N_8448,N_8580);
and U10050 (N_10050,N_8441,N_9531);
nor U10051 (N_10051,N_8830,N_8260);
or U10052 (N_10052,N_8173,N_9658);
or U10053 (N_10053,N_8948,N_9326);
nor U10054 (N_10054,N_9663,N_9471);
or U10055 (N_10055,N_8785,N_9756);
nand U10056 (N_10056,N_9903,N_8419);
nor U10057 (N_10057,N_8098,N_9738);
nor U10058 (N_10058,N_9241,N_8934);
and U10059 (N_10059,N_8057,N_8577);
nor U10060 (N_10060,N_9714,N_9136);
nor U10061 (N_10061,N_8007,N_9358);
nand U10062 (N_10062,N_8485,N_9333);
or U10063 (N_10063,N_8715,N_8586);
or U10064 (N_10064,N_9632,N_8814);
nand U10065 (N_10065,N_8891,N_9457);
nand U10066 (N_10066,N_9075,N_8069);
nand U10067 (N_10067,N_8369,N_9301);
and U10068 (N_10068,N_9741,N_9621);
or U10069 (N_10069,N_8392,N_9070);
and U10070 (N_10070,N_8165,N_9044);
or U10071 (N_10071,N_8128,N_8197);
nand U10072 (N_10072,N_9352,N_8519);
nand U10073 (N_10073,N_9176,N_9057);
nor U10074 (N_10074,N_9964,N_9573);
and U10075 (N_10075,N_8820,N_8449);
nand U10076 (N_10076,N_9019,N_8467);
or U10077 (N_10077,N_9376,N_8095);
and U10078 (N_10078,N_8406,N_9162);
and U10079 (N_10079,N_9058,N_8156);
or U10080 (N_10080,N_9906,N_8765);
or U10081 (N_10081,N_9128,N_8277);
nand U10082 (N_10082,N_9370,N_9052);
and U10083 (N_10083,N_9302,N_8547);
and U10084 (N_10084,N_9719,N_8728);
and U10085 (N_10085,N_8460,N_8134);
or U10086 (N_10086,N_9984,N_8650);
and U10087 (N_10087,N_9013,N_9952);
and U10088 (N_10088,N_9895,N_9137);
or U10089 (N_10089,N_9971,N_8179);
nand U10090 (N_10090,N_9959,N_8180);
and U10091 (N_10091,N_9283,N_9918);
or U10092 (N_10092,N_8842,N_8115);
or U10093 (N_10093,N_9863,N_8829);
or U10094 (N_10094,N_8221,N_8218);
or U10095 (N_10095,N_8037,N_8653);
and U10096 (N_10096,N_8097,N_8290);
or U10097 (N_10097,N_8943,N_9881);
nor U10098 (N_10098,N_8275,N_8094);
and U10099 (N_10099,N_9637,N_8162);
nor U10100 (N_10100,N_9272,N_8594);
and U10101 (N_10101,N_9288,N_8844);
nand U10102 (N_10102,N_9819,N_8707);
or U10103 (N_10103,N_9802,N_8603);
nor U10104 (N_10104,N_9682,N_9309);
nand U10105 (N_10105,N_8910,N_8559);
nand U10106 (N_10106,N_8996,N_8677);
nor U10107 (N_10107,N_9979,N_9754);
or U10108 (N_10108,N_8967,N_8438);
and U10109 (N_10109,N_8530,N_9934);
nor U10110 (N_10110,N_9374,N_8243);
or U10111 (N_10111,N_9239,N_9280);
nand U10112 (N_10112,N_8019,N_8486);
and U10113 (N_10113,N_8285,N_8887);
nand U10114 (N_10114,N_8540,N_8643);
nor U10115 (N_10115,N_9068,N_8048);
or U10116 (N_10116,N_8481,N_8234);
nand U10117 (N_10117,N_9253,N_8231);
or U10118 (N_10118,N_9257,N_9155);
and U10119 (N_10119,N_8744,N_8772);
nand U10120 (N_10120,N_8739,N_8388);
nand U10121 (N_10121,N_8412,N_9647);
and U10122 (N_10122,N_8043,N_9537);
and U10123 (N_10123,N_8922,N_8751);
or U10124 (N_10124,N_8962,N_8619);
nand U10125 (N_10125,N_8950,N_9251);
and U10126 (N_10126,N_9657,N_9638);
and U10127 (N_10127,N_8430,N_8391);
and U10128 (N_10128,N_9785,N_8804);
nor U10129 (N_10129,N_9947,N_8384);
nand U10130 (N_10130,N_8940,N_8002);
nand U10131 (N_10131,N_9310,N_8900);
or U10132 (N_10132,N_9748,N_8379);
nor U10133 (N_10133,N_9414,N_8480);
and U10134 (N_10134,N_9604,N_8195);
nor U10135 (N_10135,N_9586,N_8349);
or U10136 (N_10136,N_9593,N_8640);
nand U10137 (N_10137,N_9481,N_9468);
and U10138 (N_10138,N_9639,N_8301);
nand U10139 (N_10139,N_9069,N_8074);
and U10140 (N_10140,N_8371,N_8012);
nand U10141 (N_10141,N_9902,N_9497);
nor U10142 (N_10142,N_8319,N_8009);
and U10143 (N_10143,N_9595,N_9042);
nor U10144 (N_10144,N_9523,N_9942);
nor U10145 (N_10145,N_8720,N_9498);
nor U10146 (N_10146,N_8644,N_9861);
nor U10147 (N_10147,N_9544,N_8364);
and U10148 (N_10148,N_8592,N_8143);
nand U10149 (N_10149,N_9149,N_8726);
or U10150 (N_10150,N_8759,N_9502);
or U10151 (N_10151,N_8854,N_8122);
nor U10152 (N_10152,N_8250,N_8811);
and U10153 (N_10153,N_8244,N_8883);
and U10154 (N_10154,N_8896,N_9147);
nor U10155 (N_10155,N_8733,N_8065);
and U10156 (N_10156,N_8158,N_8904);
nor U10157 (N_10157,N_8799,N_9331);
nor U10158 (N_10158,N_8911,N_9496);
and U10159 (N_10159,N_8025,N_9566);
nor U10160 (N_10160,N_9345,N_9189);
nor U10161 (N_10161,N_9179,N_8008);
nand U10162 (N_10162,N_9564,N_9190);
nand U10163 (N_10163,N_9691,N_8415);
nor U10164 (N_10164,N_8223,N_9804);
or U10165 (N_10165,N_9328,N_8865);
nand U10166 (N_10166,N_8169,N_9435);
and U10167 (N_10167,N_8602,N_8746);
nand U10168 (N_10168,N_9210,N_8023);
or U10169 (N_10169,N_9308,N_9033);
nand U10170 (N_10170,N_9693,N_8898);
nand U10171 (N_10171,N_8318,N_8638);
or U10172 (N_10172,N_9501,N_9919);
and U10173 (N_10173,N_9937,N_9776);
nor U10174 (N_10174,N_9551,N_8230);
or U10175 (N_10175,N_8954,N_8153);
and U10176 (N_10176,N_9643,N_8070);
or U10177 (N_10177,N_9713,N_8131);
nor U10178 (N_10178,N_9157,N_8708);
nand U10179 (N_10179,N_8067,N_9743);
xor U10180 (N_10180,N_8248,N_9871);
and U10181 (N_10181,N_8875,N_8300);
nand U10182 (N_10182,N_8426,N_8846);
nand U10183 (N_10183,N_9303,N_9107);
or U10184 (N_10184,N_9761,N_9427);
nor U10185 (N_10185,N_8732,N_9710);
nand U10186 (N_10186,N_8434,N_8044);
nor U10187 (N_10187,N_8274,N_8874);
or U10188 (N_10188,N_9887,N_8848);
nand U10189 (N_10189,N_8464,N_9782);
nand U10190 (N_10190,N_8510,N_8957);
nand U10191 (N_10191,N_8655,N_9431);
and U10192 (N_10192,N_9698,N_9290);
nor U10193 (N_10193,N_9342,N_9549);
or U10194 (N_10194,N_8951,N_9793);
and U10195 (N_10195,N_9390,N_9565);
or U10196 (N_10196,N_9437,N_8206);
and U10197 (N_10197,N_9164,N_8148);
and U10198 (N_10198,N_8505,N_8305);
or U10199 (N_10199,N_9229,N_8374);
or U10200 (N_10200,N_9172,N_8730);
nand U10201 (N_10201,N_8743,N_9269);
and U10202 (N_10202,N_9728,N_9605);
nand U10203 (N_10203,N_8154,N_9175);
nand U10204 (N_10204,N_8328,N_8462);
and U10205 (N_10205,N_8966,N_8150);
or U10206 (N_10206,N_9525,N_8667);
or U10207 (N_10207,N_8276,N_9079);
or U10208 (N_10208,N_9737,N_9362);
nor U10209 (N_10209,N_8139,N_8447);
nor U10210 (N_10210,N_8981,N_9998);
nand U10211 (N_10211,N_8104,N_9875);
nor U10212 (N_10212,N_8693,N_8803);
and U10213 (N_10213,N_9340,N_9783);
or U10214 (N_10214,N_9559,N_9656);
nor U10215 (N_10215,N_8443,N_8183);
nand U10216 (N_10216,N_8046,N_8719);
nand U10217 (N_10217,N_9419,N_8827);
nor U10218 (N_10218,N_8237,N_8365);
and U10219 (N_10219,N_9363,N_8279);
nand U10220 (N_10220,N_8112,N_8860);
nor U10221 (N_10221,N_9567,N_9965);
or U10222 (N_10222,N_9958,N_9751);
nor U10223 (N_10223,N_9215,N_9721);
nor U10224 (N_10224,N_8531,N_8816);
and U10225 (N_10225,N_8670,N_9348);
and U10226 (N_10226,N_8110,N_9794);
nand U10227 (N_10227,N_9874,N_9181);
nor U10228 (N_10228,N_9219,N_8532);
nor U10229 (N_10229,N_9319,N_8593);
and U10230 (N_10230,N_9775,N_8083);
nand U10231 (N_10231,N_9733,N_9542);
nor U10232 (N_10232,N_9410,N_9763);
nand U10233 (N_10233,N_9932,N_8993);
or U10234 (N_10234,N_8714,N_8612);
or U10235 (N_10235,N_8587,N_9975);
nand U10236 (N_10236,N_8855,N_8212);
and U10237 (N_10237,N_9493,N_8299);
and U10238 (N_10238,N_8506,N_8202);
or U10239 (N_10239,N_9202,N_8585);
or U10240 (N_10240,N_9177,N_9703);
or U10241 (N_10241,N_8287,N_8706);
nand U10242 (N_10242,N_8264,N_8633);
nand U10243 (N_10243,N_8872,N_9681);
nor U10244 (N_10244,N_9769,N_8787);
nor U10245 (N_10245,N_9977,N_9825);
xnor U10246 (N_10246,N_8529,N_9989);
or U10247 (N_10247,N_8217,N_8863);
or U10248 (N_10248,N_8440,N_8028);
nand U10249 (N_10249,N_8171,N_9985);
and U10250 (N_10250,N_9850,N_8229);
and U10251 (N_10251,N_9712,N_9767);
or U10252 (N_10252,N_8597,N_9032);
or U10253 (N_10253,N_9807,N_8895);
nor U10254 (N_10254,N_9571,N_8987);
nor U10255 (N_10255,N_9614,N_8659);
nand U10256 (N_10256,N_8596,N_8516);
nand U10257 (N_10257,N_8325,N_8133);
or U10258 (N_10258,N_9885,N_9034);
nand U10259 (N_10259,N_9174,N_8725);
nand U10260 (N_10260,N_9711,N_8105);
nor U10261 (N_10261,N_8889,N_9907);
nand U10262 (N_10262,N_9527,N_9815);
or U10263 (N_10263,N_8856,N_9109);
nor U10264 (N_10264,N_9364,N_9629);
and U10265 (N_10265,N_9355,N_8472);
nand U10266 (N_10266,N_9722,N_9306);
and U10267 (N_10267,N_9665,N_9298);
or U10268 (N_10268,N_9209,N_8601);
or U10269 (N_10269,N_9060,N_9091);
nor U10270 (N_10270,N_9329,N_9995);
nand U10271 (N_10271,N_8347,N_9216);
nor U10272 (N_10272,N_9939,N_9377);
or U10273 (N_10273,N_8488,N_9212);
nand U10274 (N_10274,N_9612,N_8172);
nand U10275 (N_10275,N_9867,N_9833);
nor U10276 (N_10276,N_9664,N_9267);
or U10277 (N_10277,N_8437,N_9951);
nor U10278 (N_10278,N_9050,N_8631);
nor U10279 (N_10279,N_9734,N_9242);
nor U10280 (N_10280,N_9557,N_8142);
nand U10281 (N_10281,N_8521,N_9888);
or U10282 (N_10282,N_9717,N_9009);
nand U10283 (N_10283,N_9387,N_8408);
nand U10284 (N_10284,N_8256,N_9287);
and U10285 (N_10285,N_8192,N_8523);
and U10286 (N_10286,N_9407,N_8986);
nor U10287 (N_10287,N_8791,N_8698);
and U10288 (N_10288,N_9892,N_8157);
nor U10289 (N_10289,N_8252,N_8571);
and U10290 (N_10290,N_9689,N_8961);
nand U10291 (N_10291,N_9725,N_9424);
nor U10292 (N_10292,N_9236,N_8797);
and U10293 (N_10293,N_9838,N_9430);
nor U10294 (N_10294,N_8808,N_8806);
nor U10295 (N_10295,N_8227,N_8817);
nor U10296 (N_10296,N_9126,N_9543);
nand U10297 (N_10297,N_8985,N_9896);
nand U10298 (N_10298,N_8402,N_9786);
or U10299 (N_10299,N_8953,N_8893);
or U10300 (N_10300,N_9074,N_8899);
nand U10301 (N_10301,N_8080,N_8129);
and U10302 (N_10302,N_8456,N_9411);
or U10303 (N_10303,N_9514,N_9749);
nand U10304 (N_10304,N_8064,N_8479);
or U10305 (N_10305,N_9705,N_8060);
nor U10306 (N_10306,N_8599,N_8702);
nor U10307 (N_10307,N_9562,N_9135);
nand U10308 (N_10308,N_8977,N_8209);
nand U10309 (N_10309,N_9094,N_9864);
or U10310 (N_10310,N_8906,N_9585);
and U10311 (N_10311,N_8344,N_9449);
nand U10312 (N_10312,N_8963,N_9762);
and U10313 (N_10313,N_9513,N_8998);
or U10314 (N_10314,N_9660,N_9193);
and U10315 (N_10315,N_9955,N_8870);
and U10316 (N_10316,N_9312,N_9988);
and U10317 (N_10317,N_9808,N_9443);
or U10318 (N_10318,N_8727,N_8515);
nand U10319 (N_10319,N_9796,N_9666);
or U10320 (N_10320,N_8045,N_8119);
and U10321 (N_10321,N_8182,N_8666);
nor U10322 (N_10322,N_8382,N_9357);
or U10323 (N_10323,N_8674,N_9930);
or U10324 (N_10324,N_8191,N_8376);
nand U10325 (N_10325,N_9653,N_8333);
nand U10326 (N_10326,N_9083,N_9774);
and U10327 (N_10327,N_8690,N_9716);
or U10328 (N_10328,N_9779,N_9161);
xor U10329 (N_10329,N_9813,N_9247);
nand U10330 (N_10330,N_8756,N_9360);
nor U10331 (N_10331,N_8433,N_9401);
nor U10332 (N_10332,N_8442,N_8648);
or U10333 (N_10333,N_9982,N_8781);
and U10334 (N_10334,N_9603,N_9787);
nand U10335 (N_10335,N_8036,N_8590);
nor U10336 (N_10336,N_8784,N_9275);
or U10337 (N_10337,N_9528,N_9915);
nor U10338 (N_10338,N_8343,N_8685);
nor U10339 (N_10339,N_9516,N_8723);
nor U10340 (N_10340,N_9000,N_8271);
and U10341 (N_10341,N_9686,N_9974);
and U10342 (N_10342,N_8113,N_9014);
and U10343 (N_10343,N_8903,N_8782);
and U10344 (N_10344,N_8750,N_9904);
nor U10345 (N_10345,N_9037,N_9311);
or U10346 (N_10346,N_8704,N_9791);
nand U10347 (N_10347,N_8973,N_9451);
nor U10348 (N_10348,N_9465,N_9067);
nor U10349 (N_10349,N_8838,N_9954);
nand U10350 (N_10350,N_8669,N_9858);
and U10351 (N_10351,N_8414,N_9581);
nand U10352 (N_10352,N_8929,N_9913);
and U10353 (N_10353,N_8949,N_9505);
xor U10354 (N_10354,N_9113,N_8575);
nor U10355 (N_10355,N_8058,N_9056);
nor U10356 (N_10356,N_9847,N_9004);
and U10357 (N_10357,N_8598,N_8327);
nor U10358 (N_10358,N_9857,N_9214);
xnor U10359 (N_10359,N_8923,N_9921);
and U10360 (N_10360,N_9388,N_9178);
nor U10361 (N_10361,N_8062,N_8205);
nor U10362 (N_10362,N_9917,N_8151);
nor U10363 (N_10363,N_9678,N_9144);
nor U10364 (N_10364,N_9598,N_9818);
nor U10365 (N_10365,N_8016,N_8608);
or U10366 (N_10366,N_9652,N_8637);
nor U10367 (N_10367,N_9556,N_9812);
and U10368 (N_10368,N_9321,N_9213);
nand U10369 (N_10369,N_9334,N_8056);
nand U10370 (N_10370,N_8160,N_9466);
nand U10371 (N_10371,N_8079,N_9346);
nand U10372 (N_10372,N_9690,N_8114);
nor U10373 (N_10373,N_9628,N_8316);
nand U10374 (N_10374,N_9294,N_8375);
nand U10375 (N_10375,N_9809,N_9574);
or U10376 (N_10376,N_9192,N_8332);
nor U10377 (N_10377,N_8695,N_8975);
nand U10378 (N_10378,N_8003,N_8032);
and U10379 (N_10379,N_8360,N_9285);
nand U10380 (N_10380,N_8946,N_9353);
nor U10381 (N_10381,N_8635,N_9318);
or U10382 (N_10382,N_8052,N_8563);
and U10383 (N_10383,N_9826,N_9234);
and U10384 (N_10384,N_8567,N_9563);
or U10385 (N_10385,N_9967,N_9495);
or U10386 (N_10386,N_9380,N_8242);
or U10387 (N_10387,N_9122,N_8673);
nand U10388 (N_10388,N_8584,N_9244);
nand U10389 (N_10389,N_8634,N_8859);
or U10390 (N_10390,N_8964,N_8175);
and U10391 (N_10391,N_8976,N_9010);
or U10392 (N_10392,N_9768,N_8542);
nand U10393 (N_10393,N_9266,N_8017);
or U10394 (N_10394,N_8630,N_9408);
or U10395 (N_10395,N_8915,N_8972);
nand U10396 (N_10396,N_8849,N_9535);
or U10397 (N_10397,N_9517,N_8184);
and U10398 (N_10398,N_9855,N_9018);
nor U10399 (N_10399,N_9609,N_8703);
nor U10400 (N_10400,N_8613,N_9596);
nor U10401 (N_10401,N_8609,N_9538);
or U10402 (N_10402,N_9359,N_8682);
nand U10403 (N_10403,N_9633,N_9391);
nor U10404 (N_10404,N_9694,N_8483);
or U10405 (N_10405,N_9781,N_8455);
nor U10406 (N_10406,N_8886,N_9158);
nand U10407 (N_10407,N_8983,N_9217);
nor U10408 (N_10408,N_9316,N_8478);
nand U10409 (N_10409,N_9064,N_9114);
nand U10410 (N_10410,N_8663,N_9669);
and U10411 (N_10411,N_8068,N_9405);
nor U10412 (N_10412,N_9720,N_8622);
or U10413 (N_10413,N_9697,N_8701);
nand U10414 (N_10414,N_8508,N_8736);
and U10415 (N_10415,N_8116,N_8210);
nand U10416 (N_10416,N_9262,N_9445);
or U10417 (N_10417,N_8541,N_9089);
nand U10418 (N_10418,N_8465,N_8268);
and U10419 (N_10419,N_9293,N_9095);
and U10420 (N_10420,N_8468,N_9432);
nand U10421 (N_10421,N_9188,N_8283);
nor U10422 (N_10422,N_8411,N_8550);
and U10423 (N_10423,N_8558,N_8748);
and U10424 (N_10424,N_9594,N_9065);
or U10425 (N_10425,N_8001,N_8245);
nand U10426 (N_10426,N_9166,N_8825);
nor U10427 (N_10427,N_9644,N_8099);
and U10428 (N_10428,N_9008,N_9088);
and U10429 (N_10429,N_9957,N_8762);
and U10430 (N_10430,N_9274,N_9642);
and U10431 (N_10431,N_8913,N_9911);
nor U10432 (N_10432,N_8564,N_9198);
and U10433 (N_10433,N_8780,N_9651);
and U10434 (N_10434,N_8554,N_8509);
and U10435 (N_10435,N_8713,N_9462);
nor U10436 (N_10436,N_8497,N_9385);
or U10437 (N_10437,N_9824,N_8029);
or U10438 (N_10438,N_8446,N_8463);
and U10439 (N_10439,N_8353,N_8304);
or U10440 (N_10440,N_8524,N_9619);
nor U10441 (N_10441,N_9099,N_8072);
and U10442 (N_10442,N_9470,N_8936);
or U10443 (N_10443,N_8649,N_9365);
or U10444 (N_10444,N_8651,N_8969);
and U10445 (N_10445,N_9503,N_9579);
nor U10446 (N_10446,N_9956,N_8932);
nand U10447 (N_10447,N_8569,N_8494);
or U10448 (N_10448,N_8314,N_9476);
nor U10449 (N_10449,N_8409,N_8270);
or U10450 (N_10450,N_8642,N_8387);
nand U10451 (N_10451,N_9646,N_8939);
nand U10452 (N_10452,N_9877,N_8520);
nand U10453 (N_10453,N_8288,N_9397);
nand U10454 (N_10454,N_8247,N_9232);
xnor U10455 (N_10455,N_8513,N_9670);
nor U10456 (N_10456,N_8454,N_9325);
or U10457 (N_10457,N_8310,N_9226);
and U10458 (N_10458,N_9715,N_8774);
or U10459 (N_10459,N_8111,N_8867);
nand U10460 (N_10460,N_9487,N_8439);
or U10461 (N_10461,N_9584,N_9803);
or U10462 (N_10462,N_8495,N_9671);
nor U10463 (N_10463,N_9820,N_8320);
and U10464 (N_10464,N_9920,N_8935);
nand U10465 (N_10465,N_8373,N_9938);
nand U10466 (N_10466,N_8760,N_8000);
nor U10467 (N_10467,N_8331,N_9928);
nor U10468 (N_10468,N_9016,N_8198);
or U10469 (N_10469,N_8185,N_9676);
nor U10470 (N_10470,N_8222,N_9383);
or U10471 (N_10471,N_8994,N_9700);
and U10472 (N_10472,N_8298,N_9675);
nand U10473 (N_10473,N_8978,N_8100);
and U10474 (N_10474,N_9530,N_9195);
nor U10475 (N_10475,N_9944,N_8710);
nor U10476 (N_10476,N_8011,N_9732);
nor U10477 (N_10477,N_8496,N_8386);
nor U10478 (N_10478,N_9927,N_8884);
or U10479 (N_10479,N_9059,N_9739);
and U10480 (N_10480,N_9171,N_9036);
or U10481 (N_10481,N_9848,N_9993);
nor U10482 (N_10482,N_9886,N_9943);
or U10483 (N_10483,N_8077,N_8920);
nand U10484 (N_10484,N_9382,N_8611);
nand U10485 (N_10485,N_8802,N_8108);
or U10486 (N_10486,N_8742,N_8082);
and U10487 (N_10487,N_9082,N_9541);
nor U10488 (N_10488,N_9191,N_8818);
nor U10489 (N_10489,N_9709,N_8167);
nor U10490 (N_10490,N_8137,N_8737);
nor U10491 (N_10491,N_8418,N_9096);
and U10492 (N_10492,N_9218,N_8552);
and U10493 (N_10493,N_9640,N_9687);
nor U10494 (N_10494,N_9139,N_8049);
nand U10495 (N_10495,N_8570,N_9608);
nor U10496 (N_10496,N_9684,N_9327);
and U10497 (N_10497,N_8711,N_9999);
nor U10498 (N_10498,N_8536,N_9572);
or U10499 (N_10499,N_9304,N_9829);
nand U10500 (N_10500,N_9230,N_9940);
or U10501 (N_10501,N_9617,N_8356);
and U10502 (N_10502,N_9587,N_9255);
nand U10503 (N_10503,N_9916,N_9238);
nand U10504 (N_10504,N_9463,N_9049);
nand U10505 (N_10505,N_8652,N_9908);
or U10506 (N_10506,N_8351,N_9592);
nor U10507 (N_10507,N_9780,N_9415);
nor U10508 (N_10508,N_9054,N_8716);
nor U10509 (N_10509,N_8297,N_8861);
nor U10510 (N_10510,N_9314,N_8955);
or U10511 (N_10511,N_9110,N_9250);
or U10512 (N_10512,N_9529,N_9893);
or U10513 (N_10513,N_9800,N_9766);
or U10514 (N_10514,N_8489,N_9024);
nor U10515 (N_10515,N_8005,N_8317);
nor U10516 (N_10516,N_9150,N_8193);
nor U10517 (N_10517,N_8502,N_9258);
nand U10518 (N_10518,N_9368,N_8687);
or U10519 (N_10519,N_8076,N_8401);
nand U10520 (N_10520,N_8071,N_9354);
and U10521 (N_10521,N_9474,N_9418);
nand U10522 (N_10522,N_9439,N_8562);
nor U10523 (N_10523,N_9256,N_8624);
and U10524 (N_10524,N_8421,N_8801);
or U10525 (N_10525,N_8417,N_8281);
or U10526 (N_10526,N_9151,N_8346);
and U10527 (N_10527,N_8342,N_8477);
or U10528 (N_10528,N_8924,N_8282);
nor U10529 (N_10529,N_9053,N_8031);
nor U10530 (N_10530,N_9610,N_8436);
nor U10531 (N_10531,N_9961,N_9655);
or U10532 (N_10532,N_8836,N_9649);
and U10533 (N_10533,N_9084,N_9797);
and U10534 (N_10534,N_8511,N_8851);
nand U10535 (N_10535,N_8776,N_8823);
nand U10536 (N_10536,N_8626,N_9035);
nor U10537 (N_10537,N_9990,N_9910);
nand U10538 (N_10538,N_9872,N_9121);
nor U10539 (N_10539,N_8168,N_8215);
nor U10540 (N_10540,N_9182,N_9757);
nor U10541 (N_10541,N_9118,N_9622);
and U10542 (N_10542,N_9844,N_8429);
nor U10543 (N_10543,N_9810,N_8845);
and U10544 (N_10544,N_9524,N_8499);
nor U10545 (N_10545,N_8938,N_9736);
nand U10546 (N_10546,N_9395,N_8013);
nand U10547 (N_10547,N_9901,N_8588);
or U10548 (N_10548,N_9112,N_8945);
nand U10549 (N_10549,N_9111,N_8309);
or U10550 (N_10550,N_8868,N_9526);
nor U10551 (N_10551,N_9292,N_9039);
or U10552 (N_10552,N_9221,N_9521);
and U10553 (N_10553,N_9701,N_9186);
and U10554 (N_10554,N_8930,N_9442);
xor U10555 (N_10555,N_9078,N_9337);
or U10556 (N_10556,N_9997,N_9727);
and U10557 (N_10557,N_9560,N_9520);
nand U10558 (N_10558,N_8757,N_8224);
and U10559 (N_10559,N_8933,N_9012);
and U10560 (N_10560,N_9086,N_8918);
nor U10561 (N_10561,N_9452,N_8813);
nand U10562 (N_10562,N_9891,N_8815);
nand U10563 (N_10563,N_9602,N_9207);
nor U10564 (N_10564,N_9146,N_9271);
and U10565 (N_10565,N_9960,N_8312);
xor U10566 (N_10566,N_9102,N_9454);
nor U10567 (N_10567,N_9792,N_8970);
and U10568 (N_10568,N_8188,N_8553);
nand U10569 (N_10569,N_8738,N_8914);
nor U10570 (N_10570,N_9180,N_8166);
or U10571 (N_10571,N_8284,N_8717);
and U10572 (N_10572,N_9167,N_9197);
nand U10573 (N_10573,N_8262,N_9772);
or U10574 (N_10574,N_9356,N_8432);
nand U10575 (N_10575,N_9140,N_9472);
nand U10576 (N_10576,N_8621,N_9143);
or U10577 (N_10577,N_9680,N_9396);
nor U10578 (N_10578,N_8676,N_9699);
nor U10579 (N_10579,N_9635,N_9381);
or U10580 (N_10580,N_9611,N_9723);
nand U10581 (N_10581,N_8537,N_8551);
and U10582 (N_10582,N_8395,N_8876);
nand U10583 (N_10583,N_8992,N_9260);
and U10584 (N_10584,N_8773,N_8345);
nand U10585 (N_10585,N_8947,N_9740);
or U10586 (N_10586,N_8393,N_8661);
nor U10587 (N_10587,N_8623,N_9636);
and U10588 (N_10588,N_8747,N_8361);
nor U10589 (N_10589,N_9413,N_8694);
and U10590 (N_10590,N_9624,N_9040);
and U10591 (N_10591,N_9554,N_9648);
and U10592 (N_10592,N_8683,N_9991);
and U10593 (N_10593,N_8684,N_8236);
nand U10594 (N_10594,N_9168,N_9880);
and U10595 (N_10595,N_8931,N_9771);
or U10596 (N_10596,N_8090,N_8348);
or U10597 (N_10597,N_9550,N_9994);
nor U10598 (N_10598,N_8595,N_9278);
or U10599 (N_10599,N_8261,N_8616);
nor U10600 (N_10600,N_9883,N_8323);
or U10601 (N_10601,N_8689,N_9518);
or U10602 (N_10602,N_9281,N_9969);
nor U10603 (N_10603,N_8798,N_9539);
nor U10604 (N_10604,N_9105,N_9350);
nor U10605 (N_10605,N_8161,N_9773);
and U10606 (N_10606,N_8675,N_8888);
nor U10607 (N_10607,N_9577,N_8579);
or U10608 (N_10608,N_8680,N_8549);
and U10609 (N_10609,N_9464,N_9591);
nor U10610 (N_10610,N_8239,N_9482);
nor U10611 (N_10611,N_9673,N_9038);
or U10612 (N_10612,N_9582,N_8038);
nor U10613 (N_10613,N_9924,N_8614);
or U10614 (N_10614,N_9547,N_9489);
and U10615 (N_10615,N_8127,N_9946);
nor U10616 (N_10616,N_8504,N_8201);
nor U10617 (N_10617,N_9225,N_9909);
nor U10618 (N_10618,N_9051,N_9702);
or U10619 (N_10619,N_8662,N_9268);
or U10620 (N_10620,N_9672,N_8890);
and U10621 (N_10621,N_8600,N_8761);
nor U10622 (N_10622,N_8163,N_9265);
nand U10623 (N_10623,N_8035,N_8424);
nor U10624 (N_10624,N_8989,N_9320);
and U10625 (N_10625,N_8469,N_8144);
or U10626 (N_10626,N_8370,N_9305);
or U10627 (N_10627,N_9522,N_9561);
or U10628 (N_10628,N_8404,N_8292);
or U10629 (N_10629,N_9460,N_8882);
nand U10630 (N_10630,N_9438,N_9141);
and U10631 (N_10631,N_9865,N_9343);
nand U10632 (N_10632,N_8233,N_9200);
and U10633 (N_10633,N_8871,N_9941);
nor U10634 (N_10634,N_8917,N_9222);
nand U10635 (N_10635,N_8396,N_9240);
nor U10636 (N_10636,N_8204,N_9087);
or U10637 (N_10637,N_8668,N_8809);
or U10638 (N_10638,N_8539,N_9409);
or U10639 (N_10639,N_9400,N_8858);
nor U10640 (N_10640,N_8503,N_9425);
or U10641 (N_10641,N_9862,N_9735);
nor U10642 (N_10642,N_9384,N_9264);
nor U10643 (N_10643,N_9821,N_9208);
or U10644 (N_10644,N_9978,N_8420);
nor U10645 (N_10645,N_9905,N_9570);
and U10646 (N_10646,N_9097,N_8959);
and U10647 (N_10647,N_9090,N_8091);
and U10648 (N_10648,N_9249,N_8453);
nand U10649 (N_10649,N_8878,N_9315);
and U10650 (N_10650,N_9163,N_8625);
and U10651 (N_10651,N_8610,N_8357);
and U10652 (N_10652,N_8377,N_9120);
nor U10653 (N_10653,N_9347,N_8894);
and U10654 (N_10654,N_9366,N_9478);
or U10655 (N_10655,N_8482,N_9668);
and U10656 (N_10656,N_8853,N_9873);
or U10657 (N_10657,N_9499,N_9822);
nor U10658 (N_10658,N_9131,N_9597);
nand U10659 (N_10659,N_9081,N_8794);
and U10660 (N_10660,N_8253,N_8557);
or U10661 (N_10661,N_8988,N_8336);
and U10662 (N_10662,N_8136,N_9817);
nand U10663 (N_10663,N_8902,N_9185);
or U10664 (N_10664,N_9983,N_9473);
nor U10665 (N_10665,N_8397,N_8941);
and U10666 (N_10666,N_8135,N_8213);
nand U10667 (N_10667,N_9750,N_8766);
nor U10668 (N_10668,N_8219,N_9504);
or U10669 (N_10669,N_8487,N_8641);
or U10670 (N_10670,N_9394,N_9765);
nor U10671 (N_10671,N_8416,N_8498);
or U10672 (N_10672,N_9142,N_8852);
nand U10673 (N_10673,N_8130,N_9361);
and U10674 (N_10674,N_9546,N_8004);
nor U10675 (N_10675,N_9286,N_8627);
and U10676 (N_10676,N_9970,N_8658);
or U10677 (N_10677,N_8833,N_8741);
nor U10678 (N_10678,N_8211,N_9259);
or U10679 (N_10679,N_8522,N_9404);
nor U10680 (N_10680,N_9170,N_8088);
nor U10681 (N_10681,N_8238,N_8721);
or U10682 (N_10682,N_9730,N_9589);
and U10683 (N_10683,N_9245,N_8543);
and U10684 (N_10684,N_8525,N_9001);
nand U10685 (N_10685,N_9441,N_9289);
nand U10686 (N_10686,N_8620,N_8995);
nor U10687 (N_10687,N_9076,N_8840);
or U10688 (N_10688,N_8771,N_9417);
and U10689 (N_10689,N_8514,N_8084);
nor U10690 (N_10690,N_9426,N_9133);
nand U10691 (N_10691,N_9726,N_8186);
and U10692 (N_10692,N_8330,N_9132);
and U10693 (N_10693,N_8389,N_9023);
or U10694 (N_10694,N_9925,N_9580);
nor U10695 (N_10695,N_8897,N_8645);
or U10696 (N_10696,N_8968,N_8629);
or U10697 (N_10697,N_9745,N_9981);
and U10698 (N_10698,N_8909,N_8444);
or U10699 (N_10699,N_8789,N_8006);
and U10700 (N_10700,N_8734,N_9480);
nand U10701 (N_10701,N_8390,N_8126);
or U10702 (N_10702,N_8646,N_9882);
and U10703 (N_10703,N_9235,N_8329);
xor U10704 (N_10704,N_9950,N_9422);
nor U10705 (N_10705,N_8805,N_9708);
and U10706 (N_10706,N_9349,N_9798);
nand U10707 (N_10707,N_8125,N_9299);
and U10708 (N_10708,N_8777,N_9790);
nor U10709 (N_10709,N_9588,N_9692);
nor U10710 (N_10710,N_8822,N_8403);
nand U10711 (N_10711,N_9890,N_9145);
nor U10712 (N_10712,N_8226,N_9854);
and U10713 (N_10713,N_8362,N_8267);
and U10714 (N_10714,N_9552,N_8832);
or U10715 (N_10715,N_8810,N_8583);
nand U10716 (N_10716,N_8826,N_8664);
nor U10717 (N_10717,N_9313,N_8779);
nand U10718 (N_10718,N_9339,N_8050);
and U10719 (N_10719,N_9704,N_8053);
and U10720 (N_10720,N_8873,N_9491);
and U10721 (N_10721,N_9695,N_8355);
nand U10722 (N_10722,N_8303,N_8014);
nand U10723 (N_10723,N_9183,N_8246);
or U10724 (N_10724,N_9856,N_8159);
nand U10725 (N_10725,N_9912,N_8507);
nor U10726 (N_10726,N_8030,N_8572);
or U10727 (N_10727,N_9211,N_9187);
and U10728 (N_10728,N_9130,N_9332);
and U10729 (N_10729,N_8059,N_9379);
nor U10730 (N_10730,N_9066,N_8578);
or U10731 (N_10731,N_8101,N_8181);
xnor U10732 (N_10732,N_8322,N_9201);
and U10733 (N_10733,N_9583,N_9899);
and U10734 (N_10734,N_9683,N_9770);
or U10735 (N_10735,N_9119,N_8337);
or U10736 (N_10736,N_8354,N_8843);
and U10737 (N_10737,N_8731,N_8121);
nor U10738 (N_10738,N_9889,N_8118);
or U10739 (N_10739,N_9373,N_8123);
nor U10740 (N_10740,N_8367,N_9273);
and U10741 (N_10741,N_9814,N_9806);
and U10742 (N_10742,N_8249,N_9223);
or U10743 (N_10743,N_9900,N_8971);
nand U10744 (N_10744,N_8535,N_8042);
or U10745 (N_10745,N_8754,N_9827);
nand U10746 (N_10746,N_8033,N_8660);
nand U10747 (N_10747,N_9237,N_9194);
nand U10748 (N_10748,N_8493,N_9519);
nor U10749 (N_10749,N_8269,N_9021);
and U10750 (N_10750,N_9022,N_8140);
or U10751 (N_10751,N_8041,N_9962);
or U10752 (N_10752,N_9152,N_9662);
nor U10753 (N_10753,N_8272,N_8081);
nand U10754 (N_10754,N_9688,N_9488);
and U10755 (N_10755,N_9322,N_8647);
nor U10756 (N_10756,N_8841,N_9227);
nor U10757 (N_10757,N_8302,N_8124);
nor U10758 (N_10758,N_9744,N_8474);
nand U10759 (N_10759,N_8753,N_8866);
nand U10760 (N_10760,N_8568,N_8352);
nor U10761 (N_10761,N_9620,N_9816);
or U10762 (N_10762,N_9048,N_9429);
and U10763 (N_10763,N_9992,N_8548);
nor U10764 (N_10764,N_9949,N_9876);
or U10765 (N_10765,N_9046,N_9515);
nor U10766 (N_10766,N_8334,N_9986);
or U10767 (N_10767,N_8490,N_8790);
nand U10768 (N_10768,N_9976,N_8307);
or U10769 (N_10769,N_9085,N_8189);
nand U10770 (N_10770,N_8199,N_9852);
and U10771 (N_10771,N_8363,N_8089);
nand U10772 (N_10772,N_9747,N_9402);
nand U10773 (N_10773,N_8225,N_9784);
or U10774 (N_10774,N_9731,N_8451);
or U10775 (N_10775,N_8061,N_9330);
nor U10776 (N_10776,N_9043,N_9459);
nand U10777 (N_10777,N_9228,N_8010);
and U10778 (N_10778,N_8740,N_9842);
nor U10779 (N_10779,N_9558,N_9553);
and U10780 (N_10780,N_8255,N_8452);
nor U10781 (N_10781,N_8607,N_8605);
nor U10782 (N_10782,N_9801,N_8208);
or U10783 (N_10783,N_9233,N_8170);
nor U10784 (N_10784,N_8696,N_9859);
and U10785 (N_10785,N_9263,N_8722);
or U10786 (N_10786,N_9840,N_8534);
nor U10787 (N_10787,N_9764,N_8665);
nor U10788 (N_10788,N_8991,N_8881);
nor U10789 (N_10789,N_8618,N_8916);
nand U10790 (N_10790,N_8240,N_8086);
or U10791 (N_10791,N_8445,N_8544);
nand U10792 (N_10792,N_8313,N_9667);
nand U10793 (N_10793,N_9031,N_8149);
nand U10794 (N_10794,N_9433,N_9661);
and U10795 (N_10795,N_9116,N_9015);
or U10796 (N_10796,N_9103,N_9483);
or U10797 (N_10797,N_9509,N_9618);
and U10798 (N_10798,N_8286,N_8422);
nand U10799 (N_10799,N_9196,N_9005);
nand U10800 (N_10800,N_9746,N_9160);
nor U10801 (N_10801,N_9555,N_8278);
and U10802 (N_10802,N_8850,N_9869);
and U10803 (N_10803,N_8410,N_8147);
nand U10804 (N_10804,N_9324,N_9297);
or U10805 (N_10805,N_8980,N_8775);
and U10806 (N_10806,N_8692,N_9839);
or U10807 (N_10807,N_8423,N_8216);
or U10808 (N_10808,N_9788,N_9386);
xnor U10809 (N_10809,N_8755,N_8073);
and U10810 (N_10810,N_9866,N_8792);
or U10811 (N_10811,N_8944,N_9002);
or U10812 (N_10812,N_9568,N_9444);
and U10813 (N_10813,N_8257,N_8235);
and U10814 (N_10814,N_9837,N_8200);
nand U10815 (N_10815,N_9870,N_9277);
or U10816 (N_10816,N_9025,N_8258);
nor U10817 (N_10817,N_9884,N_8768);
and U10818 (N_10818,N_9199,N_8699);
or U10819 (N_10819,N_8869,N_8321);
nor U10820 (N_10820,N_9868,N_9834);
nor U10821 (N_10821,N_8546,N_8729);
or U10822 (N_10822,N_8027,N_9630);
nand U10823 (N_10823,N_9317,N_9963);
and U10824 (N_10824,N_8518,N_9569);
nand U10825 (N_10825,N_8752,N_8138);
nor U10826 (N_10826,N_8691,N_8724);
or U10827 (N_10827,N_9789,N_8398);
nor U10828 (N_10828,N_8795,N_9576);
nor U10829 (N_10829,N_8606,N_9203);
nor U10830 (N_10830,N_8656,N_9966);
or U10831 (N_10831,N_9020,N_8187);
and U10832 (N_10832,N_8901,N_9613);
or U10833 (N_10833,N_9389,N_9003);
nand U10834 (N_10834,N_8591,N_8982);
and U10835 (N_10835,N_8907,N_9369);
nand U10836 (N_10836,N_8528,N_9455);
or U10837 (N_10837,N_8617,N_9795);
nand U10838 (N_10838,N_9922,N_8054);
or U10839 (N_10839,N_8063,N_8925);
nor U10840 (N_10840,N_8339,N_8102);
nor U10841 (N_10841,N_8928,N_8990);
and U10842 (N_10842,N_8232,N_9540);
nor U10843 (N_10843,N_8109,N_8735);
or U10844 (N_10844,N_9282,N_9416);
or U10845 (N_10845,N_9845,N_9707);
nand U10846 (N_10846,N_8047,N_8807);
xnor U10847 (N_10847,N_9344,N_8425);
and U10848 (N_10848,N_9371,N_9755);
or U10849 (N_10849,N_8997,N_9968);
nand U10850 (N_10850,N_9823,N_9412);
and U10851 (N_10851,N_9276,N_8407);
nor U10852 (N_10852,N_8176,N_8879);
nor U10853 (N_10853,N_9323,N_8581);
and U10854 (N_10854,N_8927,N_9270);
or U10855 (N_10855,N_8324,N_9134);
nand U10856 (N_10856,N_8657,N_8190);
and U10857 (N_10857,N_8251,N_8174);
nor U10858 (N_10858,N_9830,N_8254);
nor U10859 (N_10859,N_9246,N_9799);
and U10860 (N_10860,N_9027,N_8107);
nand U10861 (N_10861,N_8877,N_9098);
or U10862 (N_10862,N_9654,N_9484);
and U10863 (N_10863,N_9448,N_8194);
and U10864 (N_10864,N_9841,N_9507);
nor U10865 (N_10865,N_8492,N_8839);
nand U10866 (N_10866,N_9980,N_8615);
nand U10867 (N_10867,N_9685,N_8196);
nor U10868 (N_10868,N_9295,N_9948);
nor U10869 (N_10869,N_9148,N_9494);
or U10870 (N_10870,N_9590,N_9447);
nor U10871 (N_10871,N_9007,N_8241);
nand U10872 (N_10872,N_8778,N_8380);
nor U10873 (N_10873,N_8512,N_8672);
or U10874 (N_10874,N_8040,N_9154);
nand U10875 (N_10875,N_8952,N_8960);
or U10876 (N_10876,N_8155,N_9777);
nor U10877 (N_10877,N_8533,N_8120);
or U10878 (N_10878,N_8857,N_8628);
nand U10879 (N_10879,N_9072,N_8273);
nand U10880 (N_10880,N_8862,N_8786);
nand U10881 (N_10881,N_8999,N_9996);
nor U10882 (N_10882,N_8294,N_8458);
or U10883 (N_10883,N_9047,N_9123);
and U10884 (N_10884,N_8024,N_8473);
and U10885 (N_10885,N_9724,N_9063);
and U10886 (N_10886,N_8864,N_9061);
or U10887 (N_10887,N_8709,N_8471);
or U10888 (N_10888,N_8461,N_8470);
nand U10889 (N_10889,N_8427,N_8466);
or U10890 (N_10890,N_8526,N_8561);
nand U10891 (N_10891,N_9578,N_8055);
or U10892 (N_10892,N_8296,N_9500);
or U10893 (N_10893,N_9231,N_9077);
and U10894 (N_10894,N_8366,N_8700);
and U10895 (N_10895,N_9101,N_8132);
and U10896 (N_10896,N_9860,N_9115);
nand U10897 (N_10897,N_8259,N_9778);
and U10898 (N_10898,N_8589,N_8372);
nand U10899 (N_10899,N_8758,N_8745);
nor U10900 (N_10900,N_8974,N_8835);
or U10901 (N_10901,N_8476,N_8819);
or U10902 (N_10902,N_8926,N_9224);
or U10903 (N_10903,N_9615,N_8203);
and U10904 (N_10904,N_8293,N_8880);
nand U10905 (N_10905,N_9758,N_8501);
and U10906 (N_10906,N_9372,N_9129);
nor U10907 (N_10907,N_9805,N_8831);
nor U10908 (N_10908,N_8146,N_9914);
nor U10909 (N_10909,N_9092,N_8671);
nand U10910 (N_10910,N_9631,N_9421);
nand U10911 (N_10911,N_8087,N_9486);
nand U10912 (N_10912,N_8295,N_8770);
or U10913 (N_10913,N_8604,N_8265);
nand U10914 (N_10914,N_8026,N_8681);
nor U10915 (N_10915,N_8885,N_8152);
nor U10916 (N_10916,N_8905,N_8457);
nand U10917 (N_10917,N_9367,N_8942);
and U10918 (N_10918,N_9923,N_8545);
or U10919 (N_10919,N_8812,N_9545);
or U10920 (N_10920,N_8145,N_9252);
nand U10921 (N_10921,N_9169,N_9533);
xor U10922 (N_10922,N_9254,N_9279);
nor U10923 (N_10923,N_9485,N_9599);
xnor U10924 (N_10924,N_9835,N_9696);
nand U10925 (N_10925,N_9041,N_9674);
and U10926 (N_10926,N_8106,N_8921);
and U10927 (N_10927,N_8385,N_8491);
and U10928 (N_10928,N_8400,N_9456);
nor U10929 (N_10929,N_8764,N_9929);
nor U10930 (N_10930,N_9879,N_9220);
nand U10931 (N_10931,N_8178,N_8965);
and U10932 (N_10932,N_9508,N_8431);
xnor U10933 (N_10933,N_9548,N_9461);
and U10934 (N_10934,N_9428,N_9828);
or U10935 (N_10935,N_8769,N_9436);
nor U10936 (N_10936,N_9936,N_8311);
nand U10937 (N_10937,N_9398,N_9853);
or U10938 (N_10938,N_8207,N_8338);
nand U10939 (N_10939,N_8475,N_8359);
or U10940 (N_10940,N_8828,N_8749);
nor U10941 (N_10941,N_9017,N_8289);
nand U10942 (N_10942,N_9423,N_8937);
or U10943 (N_10943,N_8435,N_8020);
nand U10944 (N_10944,N_8078,N_8821);
nand U10945 (N_10945,N_8214,N_9625);
xnor U10946 (N_10946,N_8956,N_9073);
and U10947 (N_10947,N_8800,N_8919);
or U10948 (N_10948,N_9029,N_8555);
or U10949 (N_10949,N_8326,N_9153);
nand U10950 (N_10950,N_9100,N_9506);
and U10951 (N_10951,N_9420,N_8405);
or U10952 (N_10952,N_9634,N_8450);
and U10953 (N_10953,N_9534,N_8051);
or U10954 (N_10954,N_9093,N_9742);
or U10955 (N_10955,N_8788,N_9575);
nand U10956 (N_10956,N_8892,N_9718);
nand U10957 (N_10957,N_8678,N_9030);
or U10958 (N_10958,N_8413,N_9204);
or U10959 (N_10959,N_9127,N_8022);
nor U10960 (N_10960,N_9477,N_9104);
nand U10961 (N_10961,N_8399,N_9206);
nand U10962 (N_10962,N_9261,N_9851);
xor U10963 (N_10963,N_9080,N_8679);
nor U10964 (N_10964,N_9467,N_9973);
and U10965 (N_10965,N_8015,N_9510);
nand U10966 (N_10966,N_9307,N_9351);
nand U10967 (N_10967,N_9601,N_9659);
and U10968 (N_10968,N_9933,N_9446);
and U10969 (N_10969,N_8335,N_9205);
nor U10970 (N_10970,N_9341,N_9623);
nor U10971 (N_10971,N_8688,N_8556);
nand U10972 (N_10972,N_9434,N_8340);
or U10973 (N_10973,N_9450,N_8034);
or U10974 (N_10974,N_9641,N_8566);
and U10975 (N_10975,N_9336,N_8394);
nand U10976 (N_10976,N_8378,N_9138);
nand U10977 (N_10977,N_9878,N_8912);
nor U10978 (N_10978,N_9006,N_9532);
and U10979 (N_10979,N_8636,N_9479);
or U10980 (N_10980,N_8381,N_8103);
nor U10981 (N_10981,N_9600,N_9055);
or U10982 (N_10982,N_9511,N_8428);
or U10983 (N_10983,N_8358,N_8576);
or U10984 (N_10984,N_8538,N_9469);
or U10985 (N_10985,N_9490,N_8021);
nand U10986 (N_10986,N_8560,N_8368);
and U10987 (N_10987,N_8574,N_9406);
or U10988 (N_10988,N_9729,N_9627);
nand U10989 (N_10989,N_9028,N_9399);
and U10990 (N_10990,N_9243,N_9248);
nor U10991 (N_10991,N_9335,N_9062);
nor U10992 (N_10992,N_8093,N_8280);
or U10993 (N_10993,N_9159,N_8796);
and U10994 (N_10994,N_8573,N_8075);
and U10995 (N_10995,N_9953,N_8527);
and U10996 (N_10996,N_8341,N_8383);
nand U10997 (N_10997,N_8686,N_9117);
and U10998 (N_10998,N_9811,N_9392);
or U10999 (N_10999,N_8834,N_9753);
nand U11000 (N_11000,N_8440,N_8343);
nand U11001 (N_11001,N_8514,N_9973);
or U11002 (N_11002,N_8330,N_8382);
nand U11003 (N_11003,N_9221,N_9095);
nand U11004 (N_11004,N_8345,N_9052);
nand U11005 (N_11005,N_8178,N_8228);
or U11006 (N_11006,N_9003,N_8653);
and U11007 (N_11007,N_9088,N_8493);
nand U11008 (N_11008,N_8581,N_8605);
nand U11009 (N_11009,N_8110,N_8855);
and U11010 (N_11010,N_9452,N_8384);
and U11011 (N_11011,N_8711,N_9600);
nor U11012 (N_11012,N_8691,N_8546);
and U11013 (N_11013,N_8521,N_8104);
or U11014 (N_11014,N_9497,N_8453);
or U11015 (N_11015,N_8288,N_9365);
nor U11016 (N_11016,N_8323,N_8846);
nor U11017 (N_11017,N_9309,N_9345);
nor U11018 (N_11018,N_8681,N_8417);
nor U11019 (N_11019,N_8191,N_9452);
and U11020 (N_11020,N_9028,N_8299);
and U11021 (N_11021,N_8979,N_9519);
or U11022 (N_11022,N_9923,N_8098);
and U11023 (N_11023,N_8022,N_8024);
nand U11024 (N_11024,N_9152,N_9791);
nand U11025 (N_11025,N_8923,N_9118);
nor U11026 (N_11026,N_9865,N_8056);
nor U11027 (N_11027,N_9201,N_8389);
or U11028 (N_11028,N_9211,N_9019);
nand U11029 (N_11029,N_8092,N_8413);
nand U11030 (N_11030,N_8588,N_8919);
nor U11031 (N_11031,N_9834,N_9695);
and U11032 (N_11032,N_8158,N_9494);
and U11033 (N_11033,N_9491,N_8836);
nand U11034 (N_11034,N_9457,N_9782);
or U11035 (N_11035,N_9270,N_9177);
nand U11036 (N_11036,N_8300,N_9489);
nand U11037 (N_11037,N_8485,N_9210);
nand U11038 (N_11038,N_8602,N_8232);
nor U11039 (N_11039,N_9169,N_8621);
nand U11040 (N_11040,N_8353,N_9844);
nor U11041 (N_11041,N_8576,N_9272);
or U11042 (N_11042,N_9822,N_9701);
nand U11043 (N_11043,N_8755,N_9617);
or U11044 (N_11044,N_8372,N_9193);
nand U11045 (N_11045,N_8393,N_9557);
nor U11046 (N_11046,N_9213,N_8379);
nand U11047 (N_11047,N_8840,N_8531);
nor U11048 (N_11048,N_9157,N_8679);
and U11049 (N_11049,N_8700,N_9533);
or U11050 (N_11050,N_9894,N_9152);
nor U11051 (N_11051,N_9186,N_9821);
nor U11052 (N_11052,N_8721,N_9409);
nor U11053 (N_11053,N_8140,N_9671);
nor U11054 (N_11054,N_8981,N_8514);
nor U11055 (N_11055,N_9123,N_8548);
nand U11056 (N_11056,N_9401,N_8323);
or U11057 (N_11057,N_9933,N_8840);
and U11058 (N_11058,N_9855,N_9159);
or U11059 (N_11059,N_8048,N_8884);
and U11060 (N_11060,N_8943,N_9386);
nor U11061 (N_11061,N_8033,N_9261);
nor U11062 (N_11062,N_9873,N_9959);
nor U11063 (N_11063,N_8758,N_8911);
nand U11064 (N_11064,N_9105,N_9699);
nand U11065 (N_11065,N_8030,N_9718);
and U11066 (N_11066,N_8634,N_9062);
nand U11067 (N_11067,N_8033,N_8883);
or U11068 (N_11068,N_9912,N_8806);
nand U11069 (N_11069,N_8605,N_9685);
or U11070 (N_11070,N_9604,N_8777);
or U11071 (N_11071,N_9325,N_9134);
nor U11072 (N_11072,N_9029,N_9929);
nand U11073 (N_11073,N_9886,N_8211);
nand U11074 (N_11074,N_8206,N_9830);
nor U11075 (N_11075,N_8424,N_8494);
and U11076 (N_11076,N_8867,N_9164);
or U11077 (N_11077,N_8287,N_8872);
nand U11078 (N_11078,N_8295,N_8187);
nor U11079 (N_11079,N_8892,N_8090);
nor U11080 (N_11080,N_8745,N_8671);
and U11081 (N_11081,N_9900,N_8667);
nand U11082 (N_11082,N_9188,N_8751);
and U11083 (N_11083,N_8376,N_9440);
nand U11084 (N_11084,N_9607,N_8058);
and U11085 (N_11085,N_8086,N_8016);
nor U11086 (N_11086,N_8239,N_9914);
and U11087 (N_11087,N_9125,N_9330);
or U11088 (N_11088,N_8960,N_9134);
nor U11089 (N_11089,N_8470,N_8602);
nand U11090 (N_11090,N_8468,N_8648);
and U11091 (N_11091,N_8965,N_8424);
nor U11092 (N_11092,N_9382,N_9708);
nand U11093 (N_11093,N_9950,N_8907);
or U11094 (N_11094,N_8232,N_8130);
and U11095 (N_11095,N_8118,N_9666);
nand U11096 (N_11096,N_8326,N_8437);
nand U11097 (N_11097,N_9797,N_8408);
and U11098 (N_11098,N_9535,N_8832);
and U11099 (N_11099,N_8657,N_9805);
and U11100 (N_11100,N_8674,N_8594);
or U11101 (N_11101,N_8687,N_8732);
nand U11102 (N_11102,N_9730,N_9390);
nand U11103 (N_11103,N_8033,N_8950);
nand U11104 (N_11104,N_9476,N_9251);
nor U11105 (N_11105,N_8676,N_8990);
nor U11106 (N_11106,N_9183,N_9787);
nand U11107 (N_11107,N_8616,N_9622);
or U11108 (N_11108,N_8468,N_9448);
nor U11109 (N_11109,N_8087,N_8101);
or U11110 (N_11110,N_8958,N_9300);
nor U11111 (N_11111,N_8236,N_8847);
nand U11112 (N_11112,N_8961,N_8814);
nand U11113 (N_11113,N_8726,N_9879);
and U11114 (N_11114,N_8777,N_8240);
and U11115 (N_11115,N_8615,N_8614);
and U11116 (N_11116,N_9240,N_8315);
nor U11117 (N_11117,N_9159,N_8131);
or U11118 (N_11118,N_9133,N_9859);
or U11119 (N_11119,N_8286,N_9322);
nand U11120 (N_11120,N_9964,N_9172);
nand U11121 (N_11121,N_9364,N_8242);
or U11122 (N_11122,N_9789,N_9762);
nor U11123 (N_11123,N_9415,N_8118);
nor U11124 (N_11124,N_8461,N_8934);
nor U11125 (N_11125,N_8937,N_9067);
nand U11126 (N_11126,N_8483,N_8579);
or U11127 (N_11127,N_9214,N_8710);
nor U11128 (N_11128,N_8942,N_9745);
nor U11129 (N_11129,N_9263,N_9050);
nand U11130 (N_11130,N_8912,N_8678);
or U11131 (N_11131,N_8972,N_8385);
and U11132 (N_11132,N_9325,N_9606);
and U11133 (N_11133,N_9228,N_8462);
nor U11134 (N_11134,N_9223,N_9625);
or U11135 (N_11135,N_9771,N_8964);
nand U11136 (N_11136,N_9299,N_9330);
nand U11137 (N_11137,N_9561,N_8485);
or U11138 (N_11138,N_9290,N_9769);
or U11139 (N_11139,N_9984,N_8131);
or U11140 (N_11140,N_9281,N_8685);
and U11141 (N_11141,N_8111,N_8409);
or U11142 (N_11142,N_8464,N_8682);
or U11143 (N_11143,N_8344,N_9591);
and U11144 (N_11144,N_9624,N_9652);
nand U11145 (N_11145,N_8916,N_9284);
xor U11146 (N_11146,N_9078,N_9738);
nor U11147 (N_11147,N_8381,N_9684);
nor U11148 (N_11148,N_9448,N_8186);
nand U11149 (N_11149,N_8456,N_8010);
and U11150 (N_11150,N_9577,N_8076);
and U11151 (N_11151,N_8622,N_9795);
and U11152 (N_11152,N_8526,N_9149);
nand U11153 (N_11153,N_9620,N_9888);
and U11154 (N_11154,N_9449,N_8679);
nand U11155 (N_11155,N_8539,N_9446);
nand U11156 (N_11156,N_8772,N_8601);
nor U11157 (N_11157,N_8611,N_8271);
nand U11158 (N_11158,N_9488,N_9728);
or U11159 (N_11159,N_9430,N_8214);
and U11160 (N_11160,N_8005,N_9644);
nor U11161 (N_11161,N_9245,N_9994);
and U11162 (N_11162,N_8014,N_9939);
or U11163 (N_11163,N_9138,N_8014);
or U11164 (N_11164,N_9324,N_8574);
or U11165 (N_11165,N_9620,N_8565);
nor U11166 (N_11166,N_9281,N_8696);
nand U11167 (N_11167,N_9277,N_9400);
nand U11168 (N_11168,N_9767,N_9327);
or U11169 (N_11169,N_9557,N_8529);
and U11170 (N_11170,N_8178,N_8259);
nand U11171 (N_11171,N_9417,N_8417);
nand U11172 (N_11172,N_8483,N_9810);
and U11173 (N_11173,N_9953,N_8308);
or U11174 (N_11174,N_9666,N_8052);
nand U11175 (N_11175,N_8975,N_9439);
and U11176 (N_11176,N_8478,N_9711);
nor U11177 (N_11177,N_8831,N_9153);
nor U11178 (N_11178,N_9807,N_9182);
nand U11179 (N_11179,N_9248,N_8738);
nand U11180 (N_11180,N_9568,N_8630);
and U11181 (N_11181,N_8908,N_9393);
or U11182 (N_11182,N_8453,N_8094);
xnor U11183 (N_11183,N_9754,N_9319);
nand U11184 (N_11184,N_9584,N_8574);
or U11185 (N_11185,N_8008,N_9783);
and U11186 (N_11186,N_8374,N_9197);
nor U11187 (N_11187,N_8483,N_8474);
or U11188 (N_11188,N_9676,N_8675);
nand U11189 (N_11189,N_8621,N_8436);
or U11190 (N_11190,N_8022,N_9182);
nand U11191 (N_11191,N_9979,N_9007);
nand U11192 (N_11192,N_9733,N_8219);
and U11193 (N_11193,N_8848,N_9288);
and U11194 (N_11194,N_8921,N_9816);
nand U11195 (N_11195,N_9255,N_8892);
nor U11196 (N_11196,N_9136,N_8534);
nand U11197 (N_11197,N_8704,N_8976);
and U11198 (N_11198,N_9369,N_8260);
or U11199 (N_11199,N_8086,N_8353);
and U11200 (N_11200,N_9976,N_9314);
nor U11201 (N_11201,N_8029,N_8902);
nand U11202 (N_11202,N_9841,N_8960);
and U11203 (N_11203,N_9728,N_9480);
and U11204 (N_11204,N_8387,N_8627);
and U11205 (N_11205,N_8145,N_9564);
nand U11206 (N_11206,N_9624,N_8479);
nor U11207 (N_11207,N_8633,N_9142);
xor U11208 (N_11208,N_9518,N_9710);
or U11209 (N_11209,N_9854,N_9045);
or U11210 (N_11210,N_8525,N_9845);
nor U11211 (N_11211,N_9961,N_8895);
nor U11212 (N_11212,N_8907,N_8743);
nor U11213 (N_11213,N_8137,N_8082);
or U11214 (N_11214,N_9450,N_8039);
and U11215 (N_11215,N_8456,N_8484);
nor U11216 (N_11216,N_9103,N_9579);
nor U11217 (N_11217,N_8496,N_9869);
and U11218 (N_11218,N_9529,N_9021);
nor U11219 (N_11219,N_8204,N_8282);
nor U11220 (N_11220,N_9838,N_9131);
and U11221 (N_11221,N_8412,N_9128);
and U11222 (N_11222,N_8300,N_8457);
or U11223 (N_11223,N_8948,N_9305);
nand U11224 (N_11224,N_9778,N_8693);
nand U11225 (N_11225,N_9536,N_8223);
nand U11226 (N_11226,N_8141,N_8049);
nor U11227 (N_11227,N_8468,N_8647);
nand U11228 (N_11228,N_9551,N_9914);
or U11229 (N_11229,N_8148,N_9881);
nand U11230 (N_11230,N_9218,N_8998);
or U11231 (N_11231,N_8591,N_9840);
or U11232 (N_11232,N_8430,N_9651);
or U11233 (N_11233,N_9364,N_8580);
nor U11234 (N_11234,N_8613,N_8343);
nand U11235 (N_11235,N_8763,N_8039);
and U11236 (N_11236,N_8897,N_9917);
or U11237 (N_11237,N_8276,N_8703);
or U11238 (N_11238,N_8960,N_9403);
nor U11239 (N_11239,N_8865,N_9306);
xor U11240 (N_11240,N_8230,N_9981);
and U11241 (N_11241,N_9308,N_8544);
or U11242 (N_11242,N_8525,N_8222);
nand U11243 (N_11243,N_9427,N_9828);
and U11244 (N_11244,N_8517,N_9189);
and U11245 (N_11245,N_9881,N_8696);
and U11246 (N_11246,N_8796,N_8378);
nor U11247 (N_11247,N_8630,N_9537);
nor U11248 (N_11248,N_8950,N_9237);
or U11249 (N_11249,N_9931,N_8644);
nor U11250 (N_11250,N_8827,N_9172);
and U11251 (N_11251,N_9874,N_8696);
and U11252 (N_11252,N_9665,N_8849);
nand U11253 (N_11253,N_8104,N_9817);
or U11254 (N_11254,N_8018,N_8936);
nor U11255 (N_11255,N_8777,N_8873);
nand U11256 (N_11256,N_9832,N_9316);
nand U11257 (N_11257,N_9997,N_8436);
nor U11258 (N_11258,N_8107,N_9079);
nor U11259 (N_11259,N_8172,N_8810);
nand U11260 (N_11260,N_8475,N_8227);
and U11261 (N_11261,N_8648,N_8956);
and U11262 (N_11262,N_9648,N_8581);
or U11263 (N_11263,N_9115,N_9077);
and U11264 (N_11264,N_9190,N_9662);
nor U11265 (N_11265,N_8510,N_9854);
and U11266 (N_11266,N_9766,N_9053);
and U11267 (N_11267,N_9895,N_8627);
xnor U11268 (N_11268,N_9262,N_8033);
or U11269 (N_11269,N_9489,N_9810);
nor U11270 (N_11270,N_8427,N_8860);
nor U11271 (N_11271,N_9645,N_9999);
nor U11272 (N_11272,N_9940,N_8002);
nand U11273 (N_11273,N_8266,N_9725);
and U11274 (N_11274,N_8739,N_8665);
nand U11275 (N_11275,N_8041,N_8615);
nor U11276 (N_11276,N_9308,N_9195);
and U11277 (N_11277,N_9708,N_8774);
nor U11278 (N_11278,N_9280,N_9554);
or U11279 (N_11279,N_8496,N_9579);
nor U11280 (N_11280,N_9849,N_8546);
nor U11281 (N_11281,N_8701,N_9380);
and U11282 (N_11282,N_9391,N_9889);
nor U11283 (N_11283,N_8581,N_9094);
nand U11284 (N_11284,N_9085,N_8738);
nand U11285 (N_11285,N_9168,N_9430);
nor U11286 (N_11286,N_9464,N_8259);
nand U11287 (N_11287,N_9939,N_9117);
nand U11288 (N_11288,N_8764,N_8549);
xnor U11289 (N_11289,N_8863,N_8847);
or U11290 (N_11290,N_8487,N_9312);
or U11291 (N_11291,N_9953,N_8534);
and U11292 (N_11292,N_9098,N_9628);
nor U11293 (N_11293,N_9575,N_8206);
and U11294 (N_11294,N_8454,N_8244);
nor U11295 (N_11295,N_9276,N_8342);
or U11296 (N_11296,N_9615,N_8741);
nor U11297 (N_11297,N_8467,N_9571);
and U11298 (N_11298,N_8888,N_8941);
or U11299 (N_11299,N_8529,N_9132);
nand U11300 (N_11300,N_9041,N_9902);
nor U11301 (N_11301,N_8944,N_8964);
nand U11302 (N_11302,N_8779,N_8974);
and U11303 (N_11303,N_8836,N_8796);
and U11304 (N_11304,N_8116,N_9259);
nand U11305 (N_11305,N_9059,N_9089);
or U11306 (N_11306,N_9836,N_9143);
nand U11307 (N_11307,N_9681,N_9310);
or U11308 (N_11308,N_8890,N_8158);
or U11309 (N_11309,N_9019,N_8579);
nor U11310 (N_11310,N_9449,N_9392);
nand U11311 (N_11311,N_8740,N_9161);
nand U11312 (N_11312,N_9235,N_8877);
nor U11313 (N_11313,N_9088,N_9458);
nor U11314 (N_11314,N_8477,N_9095);
nor U11315 (N_11315,N_8346,N_9350);
nand U11316 (N_11316,N_8717,N_8869);
and U11317 (N_11317,N_8228,N_9487);
nand U11318 (N_11318,N_8388,N_9501);
or U11319 (N_11319,N_9253,N_9131);
nand U11320 (N_11320,N_8306,N_8003);
and U11321 (N_11321,N_9469,N_8307);
or U11322 (N_11322,N_9586,N_8085);
or U11323 (N_11323,N_8634,N_8620);
and U11324 (N_11324,N_9504,N_8051);
nor U11325 (N_11325,N_8702,N_9680);
and U11326 (N_11326,N_8821,N_8635);
and U11327 (N_11327,N_9991,N_8776);
nand U11328 (N_11328,N_9845,N_8163);
nor U11329 (N_11329,N_8651,N_8960);
and U11330 (N_11330,N_8290,N_9599);
and U11331 (N_11331,N_9722,N_8645);
nor U11332 (N_11332,N_9671,N_8752);
nor U11333 (N_11333,N_8365,N_8737);
or U11334 (N_11334,N_9588,N_9911);
nor U11335 (N_11335,N_9349,N_9952);
nand U11336 (N_11336,N_8387,N_9996);
and U11337 (N_11337,N_8828,N_9232);
nand U11338 (N_11338,N_8410,N_9129);
nor U11339 (N_11339,N_9817,N_9928);
nor U11340 (N_11340,N_8923,N_9449);
and U11341 (N_11341,N_8370,N_8423);
or U11342 (N_11342,N_8465,N_9240);
and U11343 (N_11343,N_8285,N_8132);
nand U11344 (N_11344,N_9338,N_8582);
and U11345 (N_11345,N_9282,N_9231);
nor U11346 (N_11346,N_8061,N_9743);
and U11347 (N_11347,N_8705,N_9842);
nor U11348 (N_11348,N_8520,N_9318);
or U11349 (N_11349,N_9197,N_9854);
nor U11350 (N_11350,N_8673,N_9014);
or U11351 (N_11351,N_9189,N_9097);
nand U11352 (N_11352,N_8599,N_8164);
nor U11353 (N_11353,N_9796,N_8891);
nor U11354 (N_11354,N_8787,N_8105);
or U11355 (N_11355,N_9011,N_9370);
nor U11356 (N_11356,N_9968,N_8071);
nor U11357 (N_11357,N_8002,N_9917);
nor U11358 (N_11358,N_9825,N_9422);
and U11359 (N_11359,N_9973,N_9158);
and U11360 (N_11360,N_9278,N_8292);
nand U11361 (N_11361,N_8831,N_8550);
nand U11362 (N_11362,N_9148,N_8889);
nor U11363 (N_11363,N_9851,N_9394);
and U11364 (N_11364,N_8787,N_9507);
or U11365 (N_11365,N_9407,N_9007);
and U11366 (N_11366,N_8925,N_9044);
nand U11367 (N_11367,N_9969,N_8548);
and U11368 (N_11368,N_9829,N_9524);
nor U11369 (N_11369,N_8484,N_8623);
nand U11370 (N_11370,N_9489,N_9525);
and U11371 (N_11371,N_8441,N_8473);
nand U11372 (N_11372,N_9862,N_8897);
nand U11373 (N_11373,N_9819,N_8944);
or U11374 (N_11374,N_9019,N_8711);
nand U11375 (N_11375,N_9756,N_8927);
nand U11376 (N_11376,N_8023,N_9766);
and U11377 (N_11377,N_9382,N_9471);
nand U11378 (N_11378,N_8454,N_8061);
or U11379 (N_11379,N_8910,N_8350);
or U11380 (N_11380,N_8218,N_9809);
or U11381 (N_11381,N_9228,N_9831);
and U11382 (N_11382,N_8375,N_8940);
nor U11383 (N_11383,N_9432,N_8237);
nor U11384 (N_11384,N_8957,N_8483);
xor U11385 (N_11385,N_8946,N_8017);
or U11386 (N_11386,N_9377,N_8998);
nand U11387 (N_11387,N_9894,N_9316);
and U11388 (N_11388,N_8475,N_8372);
nor U11389 (N_11389,N_8981,N_8292);
and U11390 (N_11390,N_9017,N_8524);
or U11391 (N_11391,N_8915,N_8857);
nand U11392 (N_11392,N_9424,N_8464);
nor U11393 (N_11393,N_8344,N_8319);
or U11394 (N_11394,N_9802,N_9258);
nand U11395 (N_11395,N_9028,N_9046);
nand U11396 (N_11396,N_8880,N_8580);
nor U11397 (N_11397,N_8490,N_8813);
or U11398 (N_11398,N_8844,N_8479);
or U11399 (N_11399,N_8643,N_8341);
or U11400 (N_11400,N_8685,N_8834);
nor U11401 (N_11401,N_8373,N_9521);
and U11402 (N_11402,N_9480,N_9865);
and U11403 (N_11403,N_8309,N_9849);
nand U11404 (N_11404,N_9398,N_9022);
nand U11405 (N_11405,N_9869,N_8939);
or U11406 (N_11406,N_8746,N_8012);
and U11407 (N_11407,N_9854,N_9264);
or U11408 (N_11408,N_8141,N_9597);
nor U11409 (N_11409,N_9222,N_9559);
and U11410 (N_11410,N_9537,N_9311);
or U11411 (N_11411,N_8184,N_8540);
nor U11412 (N_11412,N_8713,N_9326);
nor U11413 (N_11413,N_9497,N_9753);
and U11414 (N_11414,N_9739,N_8797);
or U11415 (N_11415,N_8201,N_8715);
nor U11416 (N_11416,N_9527,N_9590);
nand U11417 (N_11417,N_9249,N_8019);
nor U11418 (N_11418,N_8566,N_9033);
nand U11419 (N_11419,N_8245,N_8282);
nor U11420 (N_11420,N_9049,N_8381);
nor U11421 (N_11421,N_9281,N_9108);
nand U11422 (N_11422,N_9184,N_8918);
nand U11423 (N_11423,N_9358,N_8460);
nand U11424 (N_11424,N_9280,N_8609);
or U11425 (N_11425,N_9859,N_9388);
nand U11426 (N_11426,N_8631,N_8059);
or U11427 (N_11427,N_9576,N_8148);
and U11428 (N_11428,N_8153,N_9982);
nor U11429 (N_11429,N_8827,N_8245);
nor U11430 (N_11430,N_8134,N_8843);
nor U11431 (N_11431,N_8003,N_8289);
or U11432 (N_11432,N_9647,N_8397);
nand U11433 (N_11433,N_8279,N_8449);
and U11434 (N_11434,N_8169,N_8856);
or U11435 (N_11435,N_9801,N_9738);
nand U11436 (N_11436,N_9280,N_9972);
nor U11437 (N_11437,N_8688,N_8715);
and U11438 (N_11438,N_8088,N_8987);
nand U11439 (N_11439,N_9777,N_8118);
nor U11440 (N_11440,N_9418,N_8518);
nand U11441 (N_11441,N_8145,N_9201);
nand U11442 (N_11442,N_8061,N_9896);
nand U11443 (N_11443,N_9147,N_9249);
nand U11444 (N_11444,N_8773,N_9771);
or U11445 (N_11445,N_9380,N_9881);
and U11446 (N_11446,N_8566,N_9349);
or U11447 (N_11447,N_8787,N_8381);
or U11448 (N_11448,N_9465,N_9860);
and U11449 (N_11449,N_9930,N_8189);
and U11450 (N_11450,N_9558,N_9669);
and U11451 (N_11451,N_8696,N_9811);
or U11452 (N_11452,N_8004,N_9863);
and U11453 (N_11453,N_9003,N_9133);
or U11454 (N_11454,N_8350,N_8385);
nand U11455 (N_11455,N_9077,N_8275);
nand U11456 (N_11456,N_9551,N_8275);
nor U11457 (N_11457,N_9752,N_8444);
nand U11458 (N_11458,N_8277,N_8761);
nand U11459 (N_11459,N_8560,N_9114);
or U11460 (N_11460,N_8102,N_8564);
or U11461 (N_11461,N_9077,N_9782);
nor U11462 (N_11462,N_9912,N_8782);
and U11463 (N_11463,N_8081,N_8531);
or U11464 (N_11464,N_8119,N_8347);
or U11465 (N_11465,N_9459,N_8576);
or U11466 (N_11466,N_8912,N_9328);
and U11467 (N_11467,N_9224,N_9369);
and U11468 (N_11468,N_9177,N_9995);
and U11469 (N_11469,N_9550,N_8088);
nand U11470 (N_11470,N_8239,N_9255);
nor U11471 (N_11471,N_9258,N_8546);
nand U11472 (N_11472,N_9240,N_8263);
nor U11473 (N_11473,N_9415,N_8381);
or U11474 (N_11474,N_9878,N_9288);
and U11475 (N_11475,N_9318,N_9739);
nand U11476 (N_11476,N_9620,N_9937);
nand U11477 (N_11477,N_8142,N_9820);
nor U11478 (N_11478,N_8097,N_8740);
nor U11479 (N_11479,N_9191,N_9856);
nor U11480 (N_11480,N_9620,N_8479);
nand U11481 (N_11481,N_8536,N_9578);
nand U11482 (N_11482,N_9393,N_9290);
or U11483 (N_11483,N_9333,N_9427);
and U11484 (N_11484,N_9003,N_8016);
and U11485 (N_11485,N_9958,N_8478);
and U11486 (N_11486,N_9360,N_9603);
nor U11487 (N_11487,N_8747,N_9597);
or U11488 (N_11488,N_9568,N_8008);
or U11489 (N_11489,N_8553,N_9228);
or U11490 (N_11490,N_8626,N_9303);
nand U11491 (N_11491,N_8158,N_8059);
nand U11492 (N_11492,N_9556,N_8581);
nor U11493 (N_11493,N_9599,N_9296);
or U11494 (N_11494,N_8174,N_8449);
nand U11495 (N_11495,N_9502,N_8292);
nand U11496 (N_11496,N_9918,N_9142);
and U11497 (N_11497,N_9942,N_8794);
or U11498 (N_11498,N_9672,N_8507);
nand U11499 (N_11499,N_8414,N_8135);
and U11500 (N_11500,N_8197,N_9196);
nand U11501 (N_11501,N_9642,N_9397);
nand U11502 (N_11502,N_8696,N_8417);
nand U11503 (N_11503,N_9980,N_9534);
or U11504 (N_11504,N_8276,N_8091);
nand U11505 (N_11505,N_9829,N_8595);
nand U11506 (N_11506,N_9894,N_9752);
nor U11507 (N_11507,N_8981,N_8979);
nand U11508 (N_11508,N_8360,N_8415);
and U11509 (N_11509,N_8481,N_9233);
nor U11510 (N_11510,N_9984,N_9819);
or U11511 (N_11511,N_9439,N_9735);
nand U11512 (N_11512,N_9180,N_8838);
or U11513 (N_11513,N_8931,N_8085);
nand U11514 (N_11514,N_9968,N_8429);
nor U11515 (N_11515,N_8685,N_9636);
nand U11516 (N_11516,N_9039,N_9297);
nor U11517 (N_11517,N_9863,N_8503);
and U11518 (N_11518,N_9007,N_8617);
nor U11519 (N_11519,N_8487,N_8302);
nand U11520 (N_11520,N_9271,N_8638);
nand U11521 (N_11521,N_9752,N_9094);
nor U11522 (N_11522,N_9933,N_8936);
and U11523 (N_11523,N_9410,N_9492);
nor U11524 (N_11524,N_8081,N_9201);
nand U11525 (N_11525,N_8557,N_8673);
nor U11526 (N_11526,N_8173,N_9645);
and U11527 (N_11527,N_9725,N_8583);
or U11528 (N_11528,N_8420,N_8097);
or U11529 (N_11529,N_8613,N_9841);
and U11530 (N_11530,N_9995,N_8115);
nand U11531 (N_11531,N_8697,N_8550);
nor U11532 (N_11532,N_9714,N_9707);
and U11533 (N_11533,N_8196,N_9554);
nor U11534 (N_11534,N_9251,N_8297);
and U11535 (N_11535,N_9507,N_9198);
and U11536 (N_11536,N_8743,N_8555);
nand U11537 (N_11537,N_9238,N_8570);
and U11538 (N_11538,N_9806,N_8037);
and U11539 (N_11539,N_8565,N_8466);
nand U11540 (N_11540,N_9701,N_8989);
nand U11541 (N_11541,N_9809,N_8363);
nor U11542 (N_11542,N_8838,N_8427);
nand U11543 (N_11543,N_9551,N_8813);
nor U11544 (N_11544,N_8078,N_8682);
nor U11545 (N_11545,N_8615,N_8051);
and U11546 (N_11546,N_8112,N_9824);
nor U11547 (N_11547,N_8526,N_9061);
nand U11548 (N_11548,N_9453,N_8921);
or U11549 (N_11549,N_8633,N_9541);
nor U11550 (N_11550,N_8802,N_8939);
nand U11551 (N_11551,N_8661,N_8482);
or U11552 (N_11552,N_9027,N_8439);
and U11553 (N_11553,N_8911,N_9602);
nand U11554 (N_11554,N_8347,N_9163);
and U11555 (N_11555,N_9728,N_8439);
nor U11556 (N_11556,N_9582,N_9468);
or U11557 (N_11557,N_8788,N_9816);
and U11558 (N_11558,N_9322,N_8129);
xnor U11559 (N_11559,N_9859,N_9541);
and U11560 (N_11560,N_9299,N_8522);
nor U11561 (N_11561,N_8921,N_9057);
nor U11562 (N_11562,N_8154,N_9549);
or U11563 (N_11563,N_9331,N_9837);
and U11564 (N_11564,N_8724,N_8012);
or U11565 (N_11565,N_8334,N_8345);
or U11566 (N_11566,N_8376,N_9957);
and U11567 (N_11567,N_8272,N_8720);
nor U11568 (N_11568,N_8059,N_9487);
and U11569 (N_11569,N_9499,N_9666);
or U11570 (N_11570,N_8574,N_8207);
nand U11571 (N_11571,N_9534,N_9362);
or U11572 (N_11572,N_9150,N_8327);
or U11573 (N_11573,N_9149,N_9201);
nand U11574 (N_11574,N_9862,N_9604);
xor U11575 (N_11575,N_9412,N_8200);
and U11576 (N_11576,N_8889,N_9331);
and U11577 (N_11577,N_8954,N_9197);
nand U11578 (N_11578,N_9750,N_9552);
or U11579 (N_11579,N_9477,N_9691);
or U11580 (N_11580,N_8345,N_9743);
or U11581 (N_11581,N_9465,N_8762);
nand U11582 (N_11582,N_8277,N_8043);
or U11583 (N_11583,N_9236,N_9962);
and U11584 (N_11584,N_9406,N_9862);
nor U11585 (N_11585,N_8586,N_8415);
or U11586 (N_11586,N_9063,N_8306);
and U11587 (N_11587,N_8005,N_9394);
or U11588 (N_11588,N_8295,N_9796);
nand U11589 (N_11589,N_9063,N_8983);
xnor U11590 (N_11590,N_8242,N_9854);
or U11591 (N_11591,N_9781,N_8295);
nor U11592 (N_11592,N_8237,N_8302);
nand U11593 (N_11593,N_8302,N_8236);
nand U11594 (N_11594,N_9589,N_9489);
nand U11595 (N_11595,N_9955,N_8784);
nand U11596 (N_11596,N_9728,N_9755);
nor U11597 (N_11597,N_9342,N_8335);
nand U11598 (N_11598,N_9115,N_9446);
or U11599 (N_11599,N_8434,N_9340);
or U11600 (N_11600,N_8779,N_9102);
xnor U11601 (N_11601,N_8151,N_9078);
nor U11602 (N_11602,N_9957,N_8488);
nand U11603 (N_11603,N_8768,N_9030);
nand U11604 (N_11604,N_8393,N_9293);
xnor U11605 (N_11605,N_8658,N_9806);
nor U11606 (N_11606,N_8640,N_8737);
and U11607 (N_11607,N_9359,N_8138);
and U11608 (N_11608,N_8341,N_9583);
nor U11609 (N_11609,N_9314,N_9817);
nor U11610 (N_11610,N_9759,N_8418);
or U11611 (N_11611,N_8778,N_9146);
nand U11612 (N_11612,N_9668,N_8304);
nand U11613 (N_11613,N_8339,N_9113);
or U11614 (N_11614,N_9893,N_8487);
and U11615 (N_11615,N_8997,N_9952);
and U11616 (N_11616,N_9109,N_8757);
and U11617 (N_11617,N_9462,N_9384);
or U11618 (N_11618,N_8884,N_9460);
and U11619 (N_11619,N_8233,N_9885);
or U11620 (N_11620,N_9545,N_9379);
and U11621 (N_11621,N_8181,N_8321);
or U11622 (N_11622,N_9249,N_8232);
nor U11623 (N_11623,N_9104,N_9823);
nand U11624 (N_11624,N_8522,N_8598);
nand U11625 (N_11625,N_8326,N_8988);
nand U11626 (N_11626,N_9199,N_9304);
or U11627 (N_11627,N_8515,N_8272);
nand U11628 (N_11628,N_8069,N_9590);
or U11629 (N_11629,N_9953,N_9933);
nand U11630 (N_11630,N_8127,N_9098);
and U11631 (N_11631,N_9935,N_9053);
or U11632 (N_11632,N_8117,N_8328);
or U11633 (N_11633,N_9450,N_9578);
and U11634 (N_11634,N_9425,N_9671);
or U11635 (N_11635,N_9064,N_9875);
or U11636 (N_11636,N_8441,N_9765);
nor U11637 (N_11637,N_9688,N_9674);
nor U11638 (N_11638,N_9138,N_8320);
and U11639 (N_11639,N_9641,N_9351);
and U11640 (N_11640,N_8595,N_9003);
nand U11641 (N_11641,N_8724,N_8302);
and U11642 (N_11642,N_8090,N_8964);
or U11643 (N_11643,N_8391,N_9706);
or U11644 (N_11644,N_9203,N_9131);
or U11645 (N_11645,N_8869,N_9114);
and U11646 (N_11646,N_9210,N_8194);
nor U11647 (N_11647,N_9100,N_9595);
or U11648 (N_11648,N_9466,N_8266);
and U11649 (N_11649,N_9896,N_8696);
nor U11650 (N_11650,N_9682,N_8045);
nand U11651 (N_11651,N_8101,N_8121);
nand U11652 (N_11652,N_9234,N_9573);
nand U11653 (N_11653,N_8468,N_8779);
nor U11654 (N_11654,N_9292,N_9613);
or U11655 (N_11655,N_8354,N_8026);
and U11656 (N_11656,N_8591,N_8349);
nand U11657 (N_11657,N_9592,N_8690);
nand U11658 (N_11658,N_9174,N_8897);
nor U11659 (N_11659,N_9946,N_8099);
nor U11660 (N_11660,N_8078,N_8159);
nand U11661 (N_11661,N_8178,N_9983);
or U11662 (N_11662,N_9850,N_9396);
nor U11663 (N_11663,N_8438,N_8975);
or U11664 (N_11664,N_9678,N_9204);
nand U11665 (N_11665,N_9854,N_9984);
or U11666 (N_11666,N_8740,N_8657);
nor U11667 (N_11667,N_9558,N_8883);
or U11668 (N_11668,N_9683,N_8525);
nand U11669 (N_11669,N_9515,N_8001);
or U11670 (N_11670,N_9435,N_8777);
and U11671 (N_11671,N_8701,N_9202);
and U11672 (N_11672,N_8876,N_8369);
nand U11673 (N_11673,N_8641,N_8996);
nor U11674 (N_11674,N_8175,N_9654);
and U11675 (N_11675,N_8319,N_8911);
and U11676 (N_11676,N_8875,N_9511);
and U11677 (N_11677,N_8469,N_9928);
nand U11678 (N_11678,N_9005,N_9033);
and U11679 (N_11679,N_8259,N_9656);
nand U11680 (N_11680,N_8106,N_9859);
nand U11681 (N_11681,N_8965,N_9196);
and U11682 (N_11682,N_9235,N_9450);
nor U11683 (N_11683,N_9080,N_9100);
nor U11684 (N_11684,N_9340,N_8425);
or U11685 (N_11685,N_8878,N_9048);
nand U11686 (N_11686,N_9612,N_8264);
nor U11687 (N_11687,N_9984,N_9973);
and U11688 (N_11688,N_8545,N_8275);
nor U11689 (N_11689,N_9106,N_9285);
nand U11690 (N_11690,N_9659,N_9495);
and U11691 (N_11691,N_9867,N_9385);
and U11692 (N_11692,N_9624,N_9556);
or U11693 (N_11693,N_9269,N_8924);
xor U11694 (N_11694,N_8446,N_8859);
or U11695 (N_11695,N_9485,N_8930);
and U11696 (N_11696,N_9041,N_9823);
nor U11697 (N_11697,N_9896,N_8109);
nor U11698 (N_11698,N_9507,N_8604);
or U11699 (N_11699,N_9410,N_9738);
and U11700 (N_11700,N_8164,N_9351);
nand U11701 (N_11701,N_8615,N_8534);
and U11702 (N_11702,N_8750,N_8934);
nor U11703 (N_11703,N_9554,N_9521);
nor U11704 (N_11704,N_9031,N_9282);
nand U11705 (N_11705,N_9688,N_9390);
nand U11706 (N_11706,N_9125,N_9946);
or U11707 (N_11707,N_9253,N_8644);
or U11708 (N_11708,N_9997,N_8811);
or U11709 (N_11709,N_9906,N_8256);
or U11710 (N_11710,N_9766,N_8255);
nor U11711 (N_11711,N_8496,N_9734);
xnor U11712 (N_11712,N_8896,N_8384);
or U11713 (N_11713,N_8077,N_8307);
and U11714 (N_11714,N_9097,N_8384);
or U11715 (N_11715,N_9609,N_9198);
or U11716 (N_11716,N_9077,N_8450);
or U11717 (N_11717,N_9898,N_8706);
or U11718 (N_11718,N_9798,N_8681);
nand U11719 (N_11719,N_9612,N_9483);
or U11720 (N_11720,N_9150,N_9655);
and U11721 (N_11721,N_9426,N_9431);
or U11722 (N_11722,N_9720,N_9553);
nor U11723 (N_11723,N_9172,N_8160);
and U11724 (N_11724,N_8530,N_9313);
or U11725 (N_11725,N_9176,N_9084);
or U11726 (N_11726,N_9525,N_9281);
nand U11727 (N_11727,N_8443,N_8893);
nand U11728 (N_11728,N_9925,N_9069);
and U11729 (N_11729,N_9868,N_9280);
and U11730 (N_11730,N_8149,N_8966);
and U11731 (N_11731,N_8131,N_8833);
nand U11732 (N_11732,N_9752,N_9542);
nor U11733 (N_11733,N_8491,N_9482);
or U11734 (N_11734,N_9510,N_9307);
nand U11735 (N_11735,N_8836,N_8059);
nor U11736 (N_11736,N_8465,N_9566);
and U11737 (N_11737,N_8856,N_9004);
and U11738 (N_11738,N_8218,N_9482);
nor U11739 (N_11739,N_9098,N_8701);
or U11740 (N_11740,N_8958,N_8847);
or U11741 (N_11741,N_9436,N_8580);
nand U11742 (N_11742,N_9876,N_8521);
nand U11743 (N_11743,N_9141,N_9163);
nand U11744 (N_11744,N_8784,N_8556);
and U11745 (N_11745,N_9954,N_9346);
nand U11746 (N_11746,N_9354,N_8231);
or U11747 (N_11747,N_9151,N_9099);
nand U11748 (N_11748,N_9778,N_8723);
nand U11749 (N_11749,N_9757,N_9379);
and U11750 (N_11750,N_8510,N_9670);
nor U11751 (N_11751,N_9936,N_8037);
and U11752 (N_11752,N_8112,N_9828);
xnor U11753 (N_11753,N_8122,N_8643);
or U11754 (N_11754,N_8075,N_9740);
or U11755 (N_11755,N_9351,N_8029);
and U11756 (N_11756,N_9603,N_9160);
nand U11757 (N_11757,N_9211,N_9219);
and U11758 (N_11758,N_9804,N_9344);
nor U11759 (N_11759,N_9552,N_8538);
or U11760 (N_11760,N_8856,N_9080);
nand U11761 (N_11761,N_9018,N_9507);
and U11762 (N_11762,N_8731,N_8491);
nand U11763 (N_11763,N_8732,N_9833);
and U11764 (N_11764,N_9256,N_9584);
or U11765 (N_11765,N_8227,N_9364);
or U11766 (N_11766,N_8173,N_8960);
or U11767 (N_11767,N_8487,N_9940);
or U11768 (N_11768,N_8640,N_9652);
and U11769 (N_11769,N_9993,N_8166);
or U11770 (N_11770,N_8522,N_8294);
or U11771 (N_11771,N_8450,N_9379);
and U11772 (N_11772,N_9055,N_9487);
nand U11773 (N_11773,N_9023,N_8403);
nor U11774 (N_11774,N_9813,N_8781);
and U11775 (N_11775,N_9954,N_9575);
nor U11776 (N_11776,N_8970,N_8543);
or U11777 (N_11777,N_8329,N_8904);
or U11778 (N_11778,N_8178,N_8707);
or U11779 (N_11779,N_9123,N_8090);
or U11780 (N_11780,N_8930,N_8416);
nand U11781 (N_11781,N_8389,N_9511);
nor U11782 (N_11782,N_9458,N_9912);
and U11783 (N_11783,N_8890,N_9403);
and U11784 (N_11784,N_8575,N_9513);
nand U11785 (N_11785,N_9400,N_9312);
nor U11786 (N_11786,N_8882,N_9174);
or U11787 (N_11787,N_8912,N_9929);
or U11788 (N_11788,N_8933,N_8677);
or U11789 (N_11789,N_8701,N_9128);
nor U11790 (N_11790,N_9175,N_9746);
nor U11791 (N_11791,N_8415,N_8451);
nor U11792 (N_11792,N_8315,N_8673);
or U11793 (N_11793,N_8957,N_9235);
nand U11794 (N_11794,N_8873,N_8885);
and U11795 (N_11795,N_8620,N_8754);
or U11796 (N_11796,N_9242,N_8855);
or U11797 (N_11797,N_8708,N_9840);
or U11798 (N_11798,N_9450,N_9048);
nand U11799 (N_11799,N_9774,N_9647);
and U11800 (N_11800,N_9989,N_9473);
and U11801 (N_11801,N_8881,N_9161);
nand U11802 (N_11802,N_8458,N_9805);
nand U11803 (N_11803,N_9538,N_8417);
or U11804 (N_11804,N_9344,N_8214);
or U11805 (N_11805,N_9332,N_9604);
and U11806 (N_11806,N_9578,N_8162);
or U11807 (N_11807,N_9064,N_9739);
or U11808 (N_11808,N_9879,N_8678);
or U11809 (N_11809,N_8857,N_9525);
nand U11810 (N_11810,N_9892,N_8470);
or U11811 (N_11811,N_8309,N_9824);
and U11812 (N_11812,N_9328,N_9782);
nand U11813 (N_11813,N_8495,N_9983);
nand U11814 (N_11814,N_8859,N_9627);
and U11815 (N_11815,N_8561,N_9923);
nor U11816 (N_11816,N_9676,N_9885);
nand U11817 (N_11817,N_8500,N_8164);
xnor U11818 (N_11818,N_8013,N_8952);
nand U11819 (N_11819,N_8522,N_8130);
nor U11820 (N_11820,N_8863,N_9499);
or U11821 (N_11821,N_9102,N_9606);
nor U11822 (N_11822,N_8535,N_8012);
nand U11823 (N_11823,N_8687,N_9776);
nand U11824 (N_11824,N_8979,N_9909);
nand U11825 (N_11825,N_9030,N_9958);
and U11826 (N_11826,N_9464,N_8356);
nor U11827 (N_11827,N_8557,N_9857);
or U11828 (N_11828,N_9536,N_9061);
and U11829 (N_11829,N_8506,N_9417);
nand U11830 (N_11830,N_9570,N_9660);
nor U11831 (N_11831,N_8967,N_8103);
nand U11832 (N_11832,N_9933,N_9402);
and U11833 (N_11833,N_8593,N_9684);
or U11834 (N_11834,N_9624,N_9727);
and U11835 (N_11835,N_9947,N_9479);
nor U11836 (N_11836,N_9069,N_9506);
nor U11837 (N_11837,N_8340,N_8056);
nand U11838 (N_11838,N_9303,N_9494);
or U11839 (N_11839,N_8406,N_9618);
nor U11840 (N_11840,N_9851,N_9935);
nand U11841 (N_11841,N_8605,N_9316);
nor U11842 (N_11842,N_9702,N_9767);
nor U11843 (N_11843,N_9770,N_8929);
and U11844 (N_11844,N_8928,N_9272);
or U11845 (N_11845,N_9124,N_8518);
or U11846 (N_11846,N_9051,N_9843);
nand U11847 (N_11847,N_8350,N_8615);
or U11848 (N_11848,N_8463,N_9164);
or U11849 (N_11849,N_8800,N_8358);
nand U11850 (N_11850,N_9843,N_8083);
nor U11851 (N_11851,N_9490,N_9071);
or U11852 (N_11852,N_9711,N_8614);
or U11853 (N_11853,N_8606,N_9396);
nor U11854 (N_11854,N_8088,N_8845);
nand U11855 (N_11855,N_9412,N_9905);
nand U11856 (N_11856,N_8370,N_9240);
nor U11857 (N_11857,N_8599,N_8949);
nand U11858 (N_11858,N_8471,N_9583);
and U11859 (N_11859,N_9300,N_8485);
or U11860 (N_11860,N_9481,N_9292);
or U11861 (N_11861,N_8149,N_8941);
and U11862 (N_11862,N_8839,N_8607);
nand U11863 (N_11863,N_9309,N_9979);
nor U11864 (N_11864,N_9378,N_9317);
nor U11865 (N_11865,N_8809,N_8819);
nor U11866 (N_11866,N_8068,N_9955);
nand U11867 (N_11867,N_9150,N_8627);
nor U11868 (N_11868,N_8741,N_9145);
nor U11869 (N_11869,N_9331,N_8862);
and U11870 (N_11870,N_8642,N_9503);
nor U11871 (N_11871,N_8087,N_8717);
nand U11872 (N_11872,N_9952,N_9899);
or U11873 (N_11873,N_9993,N_8968);
nand U11874 (N_11874,N_8418,N_8618);
or U11875 (N_11875,N_9020,N_9950);
nor U11876 (N_11876,N_8637,N_9993);
nor U11877 (N_11877,N_8829,N_9679);
or U11878 (N_11878,N_9216,N_8028);
nand U11879 (N_11879,N_8955,N_8954);
nand U11880 (N_11880,N_9058,N_9051);
nand U11881 (N_11881,N_9240,N_8670);
nand U11882 (N_11882,N_8015,N_8884);
nor U11883 (N_11883,N_8314,N_8193);
or U11884 (N_11884,N_8027,N_9530);
nand U11885 (N_11885,N_8206,N_8137);
and U11886 (N_11886,N_8348,N_9109);
nand U11887 (N_11887,N_8538,N_8241);
and U11888 (N_11888,N_8571,N_9564);
or U11889 (N_11889,N_9308,N_9333);
nand U11890 (N_11890,N_8144,N_8284);
nor U11891 (N_11891,N_8404,N_8173);
or U11892 (N_11892,N_8339,N_8784);
and U11893 (N_11893,N_8557,N_9578);
and U11894 (N_11894,N_8853,N_8201);
nand U11895 (N_11895,N_9461,N_8874);
nor U11896 (N_11896,N_8570,N_9856);
nor U11897 (N_11897,N_9378,N_9921);
nand U11898 (N_11898,N_9054,N_8647);
or U11899 (N_11899,N_9001,N_8656);
nand U11900 (N_11900,N_9086,N_9755);
and U11901 (N_11901,N_9023,N_8992);
and U11902 (N_11902,N_9026,N_9797);
nor U11903 (N_11903,N_8636,N_9787);
or U11904 (N_11904,N_8359,N_8519);
or U11905 (N_11905,N_9242,N_8370);
or U11906 (N_11906,N_8496,N_9203);
or U11907 (N_11907,N_8173,N_9458);
nand U11908 (N_11908,N_8385,N_9526);
nor U11909 (N_11909,N_9017,N_8573);
nor U11910 (N_11910,N_9100,N_8891);
nand U11911 (N_11911,N_9129,N_9761);
and U11912 (N_11912,N_8892,N_9497);
nand U11913 (N_11913,N_9972,N_8660);
nand U11914 (N_11914,N_8248,N_9227);
nor U11915 (N_11915,N_8162,N_8914);
or U11916 (N_11916,N_8796,N_8650);
and U11917 (N_11917,N_8971,N_9006);
nand U11918 (N_11918,N_9254,N_8603);
and U11919 (N_11919,N_9027,N_9151);
nor U11920 (N_11920,N_8663,N_9298);
nor U11921 (N_11921,N_8695,N_8217);
nand U11922 (N_11922,N_9795,N_8741);
or U11923 (N_11923,N_9602,N_8755);
or U11924 (N_11924,N_8421,N_8254);
nand U11925 (N_11925,N_8870,N_9789);
nor U11926 (N_11926,N_9717,N_9870);
or U11927 (N_11927,N_9454,N_8109);
nor U11928 (N_11928,N_8148,N_8495);
or U11929 (N_11929,N_8963,N_8672);
or U11930 (N_11930,N_9853,N_9382);
and U11931 (N_11931,N_8095,N_8813);
nand U11932 (N_11932,N_9320,N_8917);
nand U11933 (N_11933,N_9174,N_9392);
and U11934 (N_11934,N_8857,N_9490);
and U11935 (N_11935,N_9758,N_9100);
nor U11936 (N_11936,N_8644,N_9632);
and U11937 (N_11937,N_8167,N_8501);
nand U11938 (N_11938,N_9247,N_9978);
nand U11939 (N_11939,N_9703,N_9672);
nor U11940 (N_11940,N_9736,N_8535);
nand U11941 (N_11941,N_8478,N_9329);
nand U11942 (N_11942,N_9905,N_8490);
and U11943 (N_11943,N_8752,N_8576);
or U11944 (N_11944,N_8902,N_8206);
xnor U11945 (N_11945,N_8963,N_8429);
nor U11946 (N_11946,N_8320,N_9508);
nand U11947 (N_11947,N_9455,N_9474);
and U11948 (N_11948,N_8915,N_8879);
nand U11949 (N_11949,N_8880,N_8328);
nand U11950 (N_11950,N_8040,N_9982);
and U11951 (N_11951,N_9006,N_8683);
and U11952 (N_11952,N_9073,N_8260);
nand U11953 (N_11953,N_9784,N_9966);
or U11954 (N_11954,N_8630,N_8587);
nor U11955 (N_11955,N_8656,N_8193);
and U11956 (N_11956,N_8624,N_8635);
and U11957 (N_11957,N_8045,N_9629);
nand U11958 (N_11958,N_9847,N_8843);
or U11959 (N_11959,N_8411,N_9729);
or U11960 (N_11960,N_9085,N_9832);
and U11961 (N_11961,N_8424,N_8858);
or U11962 (N_11962,N_8075,N_9776);
and U11963 (N_11963,N_9422,N_8060);
nor U11964 (N_11964,N_9079,N_9875);
nor U11965 (N_11965,N_9339,N_9661);
or U11966 (N_11966,N_8438,N_9218);
and U11967 (N_11967,N_8019,N_8853);
nor U11968 (N_11968,N_9409,N_9490);
nor U11969 (N_11969,N_9578,N_8170);
nor U11970 (N_11970,N_8703,N_9781);
nor U11971 (N_11971,N_8744,N_9693);
and U11972 (N_11972,N_8989,N_9922);
nor U11973 (N_11973,N_9313,N_8574);
nand U11974 (N_11974,N_9550,N_8972);
nor U11975 (N_11975,N_8416,N_9485);
and U11976 (N_11976,N_8147,N_9194);
nor U11977 (N_11977,N_8444,N_8718);
nand U11978 (N_11978,N_8469,N_9183);
and U11979 (N_11979,N_8602,N_9253);
or U11980 (N_11980,N_8946,N_9875);
and U11981 (N_11981,N_9881,N_8515);
or U11982 (N_11982,N_9518,N_8333);
nor U11983 (N_11983,N_8223,N_8994);
nand U11984 (N_11984,N_8704,N_8972);
and U11985 (N_11985,N_9082,N_9408);
and U11986 (N_11986,N_9284,N_8441);
or U11987 (N_11987,N_8625,N_8551);
and U11988 (N_11988,N_8192,N_8379);
or U11989 (N_11989,N_9759,N_8605);
nand U11990 (N_11990,N_9581,N_9301);
nor U11991 (N_11991,N_8415,N_8955);
nand U11992 (N_11992,N_8590,N_9193);
nor U11993 (N_11993,N_9125,N_8292);
nor U11994 (N_11994,N_9022,N_8688);
and U11995 (N_11995,N_9722,N_8479);
and U11996 (N_11996,N_9994,N_8518);
nor U11997 (N_11997,N_8248,N_8415);
and U11998 (N_11998,N_8702,N_8663);
or U11999 (N_11999,N_9656,N_9525);
nand U12000 (N_12000,N_10016,N_11980);
or U12001 (N_12001,N_10972,N_10284);
and U12002 (N_12002,N_10177,N_11212);
or U12003 (N_12003,N_10823,N_11329);
and U12004 (N_12004,N_11816,N_11840);
and U12005 (N_12005,N_10741,N_11657);
nand U12006 (N_12006,N_10857,N_11169);
nand U12007 (N_12007,N_10290,N_11286);
or U12008 (N_12008,N_11711,N_10360);
nand U12009 (N_12009,N_11650,N_10143);
nor U12010 (N_12010,N_10207,N_10710);
nand U12011 (N_12011,N_11892,N_11289);
and U12012 (N_12012,N_11791,N_10317);
or U12013 (N_12013,N_10017,N_11360);
nand U12014 (N_12014,N_10196,N_11949);
or U12015 (N_12015,N_11586,N_11667);
nand U12016 (N_12016,N_10154,N_10603);
xnor U12017 (N_12017,N_11740,N_11583);
nor U12018 (N_12018,N_10519,N_11691);
or U12019 (N_12019,N_10579,N_11889);
or U12020 (N_12020,N_10870,N_11839);
nand U12021 (N_12021,N_10530,N_11049);
or U12022 (N_12022,N_10155,N_11300);
nand U12023 (N_12023,N_11746,N_10783);
nor U12024 (N_12024,N_10630,N_10964);
and U12025 (N_12025,N_10420,N_10814);
or U12026 (N_12026,N_10755,N_10193);
and U12027 (N_12027,N_10550,N_11604);
nand U12028 (N_12028,N_10294,N_10858);
or U12029 (N_12029,N_11349,N_10141);
nor U12030 (N_12030,N_11793,N_10386);
or U12031 (N_12031,N_10331,N_11836);
nand U12032 (N_12032,N_11759,N_11718);
and U12033 (N_12033,N_10657,N_11419);
and U12034 (N_12034,N_11964,N_11525);
nand U12035 (N_12035,N_11488,N_10712);
and U12036 (N_12036,N_11426,N_10397);
and U12037 (N_12037,N_10558,N_10625);
nor U12038 (N_12038,N_10943,N_10693);
nor U12039 (N_12039,N_11995,N_11254);
nor U12040 (N_12040,N_11766,N_10371);
and U12041 (N_12041,N_10535,N_10374);
and U12042 (N_12042,N_10585,N_11203);
nor U12043 (N_12043,N_10847,N_11904);
nand U12044 (N_12044,N_11361,N_10075);
nor U12045 (N_12045,N_10663,N_11120);
and U12046 (N_12046,N_11809,N_11515);
nand U12047 (N_12047,N_10804,N_10165);
and U12048 (N_12048,N_11659,N_11493);
nand U12049 (N_12049,N_11784,N_10999);
or U12050 (N_12050,N_11270,N_11029);
and U12051 (N_12051,N_10615,N_10997);
or U12052 (N_12052,N_11383,N_10714);
and U12053 (N_12053,N_10572,N_10713);
or U12054 (N_12054,N_10895,N_11460);
xnor U12055 (N_12055,N_11292,N_11073);
or U12056 (N_12056,N_11854,N_11089);
or U12057 (N_12057,N_10327,N_11531);
nor U12058 (N_12058,N_11055,N_10656);
or U12059 (N_12059,N_10731,N_11577);
nor U12060 (N_12060,N_11370,N_10174);
and U12061 (N_12061,N_11883,N_11710);
and U12062 (N_12062,N_10012,N_10536);
nand U12063 (N_12063,N_10030,N_10853);
nand U12064 (N_12064,N_11037,N_10867);
nand U12065 (N_12065,N_11931,N_10215);
nand U12066 (N_12066,N_10932,N_11480);
nor U12067 (N_12067,N_10139,N_10977);
nor U12068 (N_12068,N_10310,N_10307);
and U12069 (N_12069,N_10130,N_11176);
or U12070 (N_12070,N_11000,N_11785);
or U12071 (N_12071,N_10481,N_11844);
nand U12072 (N_12072,N_10238,N_11496);
or U12073 (N_12073,N_10337,N_10808);
nor U12074 (N_12074,N_10072,N_10147);
and U12075 (N_12075,N_10569,N_11782);
or U12076 (N_12076,N_11162,N_10295);
and U12077 (N_12077,N_11396,N_10034);
nand U12078 (N_12078,N_10326,N_10864);
nand U12079 (N_12079,N_11321,N_11754);
and U12080 (N_12080,N_10476,N_10230);
and U12081 (N_12081,N_10396,N_11078);
or U12082 (N_12082,N_11533,N_11720);
and U12083 (N_12083,N_11502,N_11170);
or U12084 (N_12084,N_10559,N_10511);
and U12085 (N_12085,N_10753,N_11234);
and U12086 (N_12086,N_11530,N_11882);
nand U12087 (N_12087,N_11081,N_10865);
xnor U12088 (N_12088,N_10834,N_11783);
nor U12089 (N_12089,N_10276,N_10445);
or U12090 (N_12090,N_11192,N_10850);
and U12091 (N_12091,N_11975,N_11541);
nor U12092 (N_12092,N_11601,N_11977);
and U12093 (N_12093,N_10522,N_11544);
and U12094 (N_12094,N_11744,N_11699);
or U12095 (N_12095,N_10840,N_11005);
or U12096 (N_12096,N_11056,N_10925);
nor U12097 (N_12097,N_11510,N_10415);
and U12098 (N_12098,N_11859,N_11210);
and U12099 (N_12099,N_11163,N_10491);
or U12100 (N_12100,N_10115,N_11838);
xor U12101 (N_12101,N_10768,N_10869);
and U12102 (N_12102,N_10031,N_11171);
nand U12103 (N_12103,N_11907,N_10533);
nand U12104 (N_12104,N_10578,N_11774);
or U12105 (N_12105,N_11963,N_11211);
nand U12106 (N_12106,N_11725,N_11695);
and U12107 (N_12107,N_10939,N_10968);
nor U12108 (N_12108,N_10583,N_11933);
or U12109 (N_12109,N_11767,N_10844);
nand U12110 (N_12110,N_11866,N_11735);
nand U12111 (N_12111,N_11962,N_11296);
or U12112 (N_12112,N_11112,N_11214);
nor U12113 (N_12113,N_10984,N_10375);
nand U12114 (N_12114,N_10128,N_11334);
nor U12115 (N_12115,N_10313,N_10268);
nor U12116 (N_12116,N_10291,N_11602);
nor U12117 (N_12117,N_11475,N_10561);
and U12118 (N_12118,N_11989,N_10286);
nand U12119 (N_12119,N_10717,N_11034);
nor U12120 (N_12120,N_10863,N_11167);
and U12121 (N_12121,N_11679,N_10392);
or U12122 (N_12122,N_11158,N_10347);
nand U12123 (N_12123,N_11864,N_10759);
or U12124 (N_12124,N_10127,N_10500);
or U12125 (N_12125,N_10736,N_10330);
nor U12126 (N_12126,N_11527,N_10916);
and U12127 (N_12127,N_10354,N_11416);
nor U12128 (N_12128,N_11730,N_11431);
or U12129 (N_12129,N_10362,N_11960);
nand U12130 (N_12130,N_10711,N_11134);
or U12131 (N_12131,N_11812,N_10953);
nand U12132 (N_12132,N_10880,N_11654);
or U12133 (N_12133,N_10812,N_11757);
and U12134 (N_12134,N_10894,N_10624);
and U12135 (N_12135,N_11570,N_11803);
and U12136 (N_12136,N_11547,N_10325);
nand U12137 (N_12137,N_10049,N_11393);
nand U12138 (N_12138,N_10231,N_10746);
or U12139 (N_12139,N_11550,N_10541);
or U12140 (N_12140,N_10497,N_11568);
or U12141 (N_12141,N_11605,N_11154);
nor U12142 (N_12142,N_10233,N_11806);
nor U12143 (N_12143,N_10904,N_11756);
and U12144 (N_12144,N_11058,N_11312);
or U12145 (N_12145,N_11467,N_11161);
nand U12146 (N_12146,N_11362,N_11956);
nand U12147 (N_12147,N_10971,N_11436);
or U12148 (N_12148,N_11578,N_10660);
nand U12149 (N_12149,N_11445,N_11213);
and U12150 (N_12150,N_11748,N_10470);
nand U12151 (N_12151,N_11202,N_11378);
nor U12152 (N_12152,N_11469,N_11165);
nor U12153 (N_12153,N_11538,N_10239);
nand U12154 (N_12154,N_11672,N_10408);
nor U12155 (N_12155,N_10764,N_10503);
nor U12156 (N_12156,N_11596,N_10987);
nor U12157 (N_12157,N_10796,N_11109);
and U12158 (N_12158,N_10600,N_10906);
nor U12159 (N_12159,N_10223,N_10632);
nand U12160 (N_12160,N_11282,N_11841);
and U12161 (N_12161,N_10667,N_10209);
and U12162 (N_12162,N_11193,N_10947);
nor U12163 (N_12163,N_10794,N_10222);
and U12164 (N_12164,N_10555,N_11579);
nor U12165 (N_12165,N_11326,N_11022);
nor U12166 (N_12166,N_11208,N_11595);
nand U12167 (N_12167,N_11734,N_11339);
nand U12168 (N_12168,N_11603,N_11584);
nand U12169 (N_12169,N_10831,N_10664);
nand U12170 (N_12170,N_11015,N_11983);
or U12171 (N_12171,N_10696,N_10952);
and U12172 (N_12172,N_11622,N_10285);
nand U12173 (N_12173,N_11155,N_10817);
nand U12174 (N_12174,N_11855,N_11990);
or U12175 (N_12175,N_10961,N_10626);
nor U12176 (N_12176,N_11148,N_11144);
nor U12177 (N_12177,N_10591,N_10043);
or U12178 (N_12178,N_11072,N_10532);
nand U12179 (N_12179,N_10403,N_10169);
nor U12180 (N_12180,N_11412,N_11523);
and U12181 (N_12181,N_11441,N_10105);
or U12182 (N_12182,N_10227,N_10681);
nor U12183 (N_12183,N_10260,N_11149);
and U12184 (N_12184,N_11593,N_10734);
and U12185 (N_12185,N_10121,N_11986);
nand U12186 (N_12186,N_11130,N_10960);
or U12187 (N_12187,N_11779,N_10926);
and U12188 (N_12188,N_11094,N_10084);
or U12189 (N_12189,N_11035,N_11438);
and U12190 (N_12190,N_11115,N_11850);
nor U12191 (N_12191,N_11910,N_11944);
nand U12192 (N_12192,N_10885,N_11076);
nand U12193 (N_12193,N_10773,N_10526);
nand U12194 (N_12194,N_10502,N_11249);
nand U12195 (N_12195,N_10903,N_11722);
nor U12196 (N_12196,N_10039,N_11863);
nand U12197 (N_12197,N_10411,N_11733);
or U12198 (N_12198,N_11886,N_10190);
and U12199 (N_12199,N_10597,N_10252);
nor U12200 (N_12200,N_11898,N_10232);
or U12201 (N_12201,N_11253,N_10944);
nor U12202 (N_12202,N_11700,N_10750);
and U12203 (N_12203,N_10265,N_10152);
and U12204 (N_12204,N_10395,N_10671);
and U12205 (N_12205,N_11824,N_11002);
and U12206 (N_12206,N_11633,N_11057);
nand U12207 (N_12207,N_10669,N_11204);
and U12208 (N_12208,N_11209,N_11639);
and U12209 (N_12209,N_11505,N_11317);
or U12210 (N_12210,N_11755,N_10376);
nand U12211 (N_12211,N_11495,N_11887);
or U12212 (N_12212,N_10272,N_11999);
nor U12213 (N_12213,N_10157,N_10387);
nand U12214 (N_12214,N_10339,N_11994);
xor U12215 (N_12215,N_10905,N_11367);
nand U12216 (N_12216,N_11311,N_10274);
xnor U12217 (N_12217,N_10884,N_10319);
nand U12218 (N_12218,N_11379,N_11458);
or U12219 (N_12219,N_11860,N_11091);
or U12220 (N_12220,N_11871,N_11869);
or U12221 (N_12221,N_11542,N_11102);
nand U12222 (N_12222,N_10361,N_11125);
or U12223 (N_12223,N_11821,N_11008);
or U12224 (N_12224,N_10720,N_11357);
and U12225 (N_12225,N_10279,N_10547);
and U12226 (N_12226,N_11561,N_11265);
and U12227 (N_12227,N_11644,N_10336);
nand U12228 (N_12228,N_11512,N_10888);
nor U12229 (N_12229,N_10920,N_10056);
nor U12230 (N_12230,N_11786,N_11556);
xor U12231 (N_12231,N_10846,N_10173);
and U12232 (N_12232,N_11181,N_11314);
xor U12233 (N_12233,N_11566,N_10874);
and U12234 (N_12234,N_11724,N_11498);
or U12235 (N_12235,N_11677,N_11781);
nand U12236 (N_12236,N_10872,N_10088);
nand U12237 (N_12237,N_11385,N_10979);
and U12238 (N_12238,N_11492,N_10033);
or U12239 (N_12239,N_11937,N_10937);
and U12240 (N_12240,N_11683,N_11220);
nand U12241 (N_12241,N_10551,N_10060);
nand U12242 (N_12242,N_10311,N_10670);
and U12243 (N_12243,N_11662,N_10076);
nor U12244 (N_12244,N_11908,N_10191);
nand U12245 (N_12245,N_11301,N_11663);
nand U12246 (N_12246,N_10527,N_10614);
nand U12247 (N_12247,N_11688,N_10845);
nand U12248 (N_12248,N_10654,N_11477);
or U12249 (N_12249,N_11053,N_10728);
nor U12250 (N_12250,N_10422,N_11293);
and U12251 (N_12251,N_10214,N_10598);
or U12252 (N_12252,N_10269,N_11664);
nor U12253 (N_12253,N_10849,N_11111);
nor U12254 (N_12254,N_10504,N_11137);
or U12255 (N_12255,N_10228,N_10258);
nor U12256 (N_12256,N_11719,N_11074);
nor U12257 (N_12257,N_10062,N_10998);
nor U12258 (N_12258,N_10458,N_10004);
and U12259 (N_12259,N_10645,N_11923);
and U12260 (N_12260,N_10562,N_10065);
nand U12261 (N_12261,N_11952,N_10014);
nand U12262 (N_12262,N_10457,N_11777);
xnor U12263 (N_12263,N_10638,N_10086);
or U12264 (N_12264,N_10967,N_10661);
nor U12265 (N_12265,N_11592,N_10158);
nor U12266 (N_12266,N_10800,N_10119);
and U12267 (N_12267,N_10862,N_11518);
nor U12268 (N_12268,N_11743,N_10868);
nand U12269 (N_12269,N_11364,N_11397);
or U12270 (N_12270,N_10881,N_10048);
and U12271 (N_12271,N_11857,N_11447);
nor U12272 (N_12272,N_10015,N_10256);
nor U12273 (N_12273,N_11514,N_11197);
or U12274 (N_12274,N_10367,N_10003);
nor U12275 (N_12275,N_11375,N_10483);
nor U12276 (N_12276,N_11377,N_10795);
or U12277 (N_12277,N_10974,N_11105);
and U12278 (N_12278,N_11872,N_11064);
nor U12279 (N_12279,N_10827,N_10406);
and U12280 (N_12280,N_10404,N_10568);
nor U12281 (N_12281,N_10402,N_11909);
and U12282 (N_12282,N_10898,N_10582);
or U12283 (N_12283,N_11283,N_11307);
nor U12284 (N_12284,N_11299,N_10560);
nor U12285 (N_12285,N_10584,N_11951);
nand U12286 (N_12286,N_11351,N_10655);
nand U12287 (N_12287,N_10343,N_10006);
nor U12288 (N_12288,N_10702,N_10907);
and U12289 (N_12289,N_11415,N_11814);
nand U12290 (N_12290,N_10460,N_11372);
and U12291 (N_12291,N_11018,N_10142);
nand U12292 (N_12292,N_10125,N_10647);
or U12293 (N_12293,N_10349,N_10521);
or U12294 (N_12294,N_10097,N_11080);
and U12295 (N_12295,N_10213,N_10529);
nor U12296 (N_12296,N_10619,N_10698);
or U12297 (N_12297,N_11780,N_10303);
and U12298 (N_12298,N_10355,N_11084);
and U12299 (N_12299,N_11483,N_10855);
and U12300 (N_12300,N_11331,N_11770);
or U12301 (N_12301,N_11065,N_11571);
nor U12302 (N_12302,N_10724,N_10793);
nand U12303 (N_12303,N_11261,N_10927);
nor U12304 (N_12304,N_11304,N_10861);
nand U12305 (N_12305,N_10643,N_10449);
and U12306 (N_12306,N_11635,N_10455);
or U12307 (N_12307,N_10109,N_11276);
nor U12308 (N_12308,N_10520,N_11016);
nand U12309 (N_12309,N_11676,N_11520);
or U12310 (N_12310,N_11608,N_11340);
and U12311 (N_12311,N_10172,N_11052);
nor U12312 (N_12312,N_11096,N_10441);
nand U12313 (N_12313,N_11063,N_10292);
nor U12314 (N_12314,N_11926,N_10144);
or U12315 (N_12315,N_11215,N_11972);
and U12316 (N_12316,N_10554,N_11764);
nor U12317 (N_12317,N_10866,N_10766);
nand U12318 (N_12318,N_10994,N_11966);
or U12319 (N_12319,N_10924,N_10358);
nor U12320 (N_12320,N_10140,N_10480);
nand U12321 (N_12321,N_10672,N_11108);
and U12322 (N_12322,N_10391,N_10475);
and U12323 (N_12323,N_10225,N_10123);
and U12324 (N_12324,N_11686,N_10873);
nor U12325 (N_12325,N_11559,N_11189);
and U12326 (N_12326,N_10240,N_11801);
nor U12327 (N_12327,N_11858,N_11902);
and U12328 (N_12328,N_10694,N_10381);
nand U12329 (N_12329,N_10093,N_10778);
nand U12330 (N_12330,N_10691,N_11879);
xor U12331 (N_12331,N_11228,N_11600);
and U12332 (N_12332,N_11647,N_11621);
nand U12333 (N_12333,N_11328,N_11742);
and U12334 (N_12334,N_11519,N_10718);
nand U12335 (N_12335,N_10917,N_10416);
nand U12336 (N_12336,N_10452,N_10524);
and U12337 (N_12337,N_11625,N_11444);
nor U12338 (N_12338,N_11653,N_10236);
and U12339 (N_12339,N_10132,N_10627);
nand U12340 (N_12340,N_11930,N_10309);
and U12341 (N_12341,N_10482,N_11623);
nor U12342 (N_12342,N_11955,N_11051);
and U12343 (N_12343,N_10176,N_10891);
or U12344 (N_12344,N_10245,N_11443);
nand U12345 (N_12345,N_11403,N_10918);
and U12346 (N_12346,N_10803,N_10138);
or U12347 (N_12347,N_11924,N_10353);
nand U12348 (N_12348,N_10563,N_11086);
nor U12349 (N_12349,N_11732,N_10590);
or U12350 (N_12350,N_10675,N_11500);
and U12351 (N_12351,N_10604,N_11459);
nand U12352 (N_12352,N_11551,N_10574);
and U12353 (N_12353,N_10162,N_10267);
and U12354 (N_12354,N_10548,N_11287);
and U12355 (N_12355,N_11190,N_11819);
or U12356 (N_12356,N_11643,N_10243);
nor U12357 (N_12357,N_10911,N_10444);
or U12358 (N_12358,N_11017,N_11828);
nand U12359 (N_12359,N_11790,N_10565);
or U12360 (N_12360,N_10414,N_11979);
nand U12361 (N_12361,N_10807,N_10350);
and U12362 (N_12362,N_11545,N_11565);
or U12363 (N_12363,N_11888,N_10836);
nor U12364 (N_12364,N_10703,N_11151);
nand U12365 (N_12365,N_10463,N_10370);
and U12366 (N_12366,N_10606,N_11030);
nand U12367 (N_12367,N_11927,N_10447);
or U12368 (N_12368,N_11143,N_11395);
or U12369 (N_12369,N_11549,N_11354);
nor U12370 (N_12370,N_11697,N_11284);
and U12371 (N_12371,N_11591,N_10963);
or U12372 (N_12372,N_10499,N_10930);
or U12373 (N_12373,N_10875,N_10277);
or U12374 (N_12374,N_11713,N_11465);
and U12375 (N_12375,N_11087,N_10639);
nor U12376 (N_12376,N_11696,N_10423);
nand U12377 (N_12377,N_10421,N_10822);
nand U12378 (N_12378,N_10958,N_10087);
and U12379 (N_12379,N_11420,N_11487);
or U12380 (N_12380,N_10799,N_10296);
or U12381 (N_12381,N_11100,N_10393);
and U12382 (N_12382,N_10212,N_10512);
nor U12383 (N_12383,N_10612,N_11557);
and U12384 (N_12384,N_10593,N_11333);
and U12385 (N_12385,N_11342,N_10777);
nor U12386 (N_12386,N_11731,N_10767);
and U12387 (N_12387,N_11306,N_10107);
nand U12388 (N_12388,N_11618,N_11229);
or U12389 (N_12389,N_11433,N_11043);
nand U12390 (N_12390,N_11244,N_10271);
or U12391 (N_12391,N_11012,N_10095);
nand U12392 (N_12392,N_10024,N_10771);
and U12393 (N_12393,N_10431,N_11726);
and U12394 (N_12394,N_11666,N_10129);
and U12395 (N_12395,N_11238,N_10727);
or U12396 (N_12396,N_10709,N_11205);
nand U12397 (N_12397,N_11818,N_10915);
nor U12398 (N_12398,N_11421,N_11581);
nand U12399 (N_12399,N_11344,N_10506);
and U12400 (N_12400,N_10468,N_11552);
nor U12401 (N_12401,N_10513,N_11010);
xnor U12402 (N_12402,N_11124,N_10889);
nand U12403 (N_12403,N_11671,N_10020);
nor U12404 (N_12404,N_11524,N_11997);
nor U12405 (N_12405,N_11231,N_10025);
or U12406 (N_12406,N_11954,N_10453);
and U12407 (N_12407,N_10146,N_11142);
or U12408 (N_12408,N_10306,N_10580);
nand U12409 (N_12409,N_10534,N_10662);
nor U12410 (N_12410,N_11316,N_11745);
nand U12411 (N_12411,N_10485,N_11153);
and U12412 (N_12412,N_11437,N_10298);
nand U12413 (N_12413,N_11940,N_10465);
or U12414 (N_12414,N_10848,N_11322);
and U12415 (N_12415,N_11690,N_11895);
nor U12416 (N_12416,N_10743,N_11799);
nor U12417 (N_12417,N_11893,N_10544);
nor U12418 (N_12418,N_10249,N_10882);
nor U12419 (N_12419,N_10948,N_10488);
nor U12420 (N_12420,N_10659,N_11626);
nand U12421 (N_12421,N_10556,N_10929);
and U12422 (N_12422,N_10389,N_11281);
nor U12423 (N_12423,N_11548,N_10424);
or U12424 (N_12424,N_10137,N_10496);
and U12425 (N_12425,N_10970,N_10270);
nand U12426 (N_12426,N_11906,N_10305);
and U12427 (N_12427,N_10912,N_10321);
or U12428 (N_12428,N_10384,N_10705);
nor U12429 (N_12429,N_11262,N_11499);
or U12430 (N_12430,N_10022,N_11775);
and U12431 (N_12431,N_10312,N_10913);
and U12432 (N_12432,N_11598,N_10642);
nor U12433 (N_12433,N_11309,N_10540);
and U12434 (N_12434,N_11411,N_10380);
nor U12435 (N_12435,N_10697,N_11938);
nor U12436 (N_12436,N_11765,N_10262);
nand U12437 (N_12437,N_11380,N_11627);
nand U12438 (N_12438,N_10955,N_10721);
or U12439 (N_12439,N_10826,N_10641);
nand U12440 (N_12440,N_10378,N_10382);
and U12441 (N_12441,N_10013,N_11629);
nor U12442 (N_12442,N_10167,N_10346);
nor U12443 (N_12443,N_11652,N_10029);
nor U12444 (N_12444,N_10782,N_10108);
and U12445 (N_12445,N_10037,N_10185);
nand U12446 (N_12446,N_11714,N_10886);
and U12447 (N_12447,N_11760,N_10516);
nor U12448 (N_12448,N_10324,N_11389);
and U12449 (N_12449,N_11597,N_10852);
or U12450 (N_12450,N_11723,N_11269);
nand U12451 (N_12451,N_10435,N_10082);
nand U12452 (N_12452,N_11297,N_10484);
and U12453 (N_12453,N_10412,N_11381);
nand U12454 (N_12454,N_11223,N_11969);
or U12455 (N_12455,N_10204,N_11414);
or U12456 (N_12456,N_11862,N_11707);
nand U12457 (N_12457,N_11126,N_10234);
or U12458 (N_12458,N_10980,N_10220);
nand U12459 (N_12459,N_11615,N_11225);
and U12460 (N_12460,N_11885,N_10798);
or U12461 (N_12461,N_11646,N_11693);
and U12462 (N_12462,N_10035,N_10170);
or U12463 (N_12463,N_11028,N_10077);
or U12464 (N_12464,N_10893,N_11845);
or U12465 (N_12465,N_11182,N_10450);
nor U12466 (N_12466,N_10877,N_11092);
nor U12467 (N_12467,N_11939,N_10405);
or U12468 (N_12468,N_11484,N_11425);
and U12469 (N_12469,N_11356,N_10618);
nand U12470 (N_12470,N_11024,N_10890);
and U12471 (N_12471,N_10101,N_10007);
xnor U12472 (N_12472,N_11788,N_11698);
or U12473 (N_12473,N_11318,N_10079);
or U12474 (N_12474,N_11808,N_11494);
and U12475 (N_12475,N_10791,N_10195);
nand U12476 (N_12476,N_11992,N_10991);
or U12477 (N_12477,N_11922,N_10658);
nor U12478 (N_12478,N_11180,N_10250);
nor U12479 (N_12479,N_10477,N_10687);
or U12480 (N_12480,N_11852,N_11179);
nor U12481 (N_12481,N_10942,N_10951);
or U12482 (N_12482,N_11832,N_11874);
nand U12483 (N_12483,N_10308,N_11440);
and U12484 (N_12484,N_11807,N_11794);
nor U12485 (N_12485,N_10224,N_10011);
or U12486 (N_12486,N_11490,N_11829);
nand U12487 (N_12487,N_11474,N_11772);
and U12488 (N_12488,N_11656,N_10280);
and U12489 (N_12489,N_10100,N_11705);
nand U12490 (N_12490,N_10649,N_11408);
and U12491 (N_12491,N_10610,N_11422);
and U12492 (N_12492,N_10909,N_10809);
and U12493 (N_12493,N_10892,N_10828);
nand U12494 (N_12494,N_10957,N_10282);
nand U12495 (N_12495,N_11555,N_10134);
or U12496 (N_12496,N_11753,N_11513);
xnor U12497 (N_12497,N_10686,N_10027);
and U12498 (N_12498,N_11589,N_10175);
nand U12499 (N_12499,N_11061,N_10253);
nor U12500 (N_12500,N_11023,N_11201);
or U12501 (N_12501,N_11708,N_10990);
xor U12502 (N_12502,N_10928,N_11516);
and U12503 (N_12503,N_11925,N_11973);
or U12504 (N_12504,N_10426,N_10333);
nor U12505 (N_12505,N_11655,N_10797);
xor U12506 (N_12506,N_10473,N_10851);
and U12507 (N_12507,N_10495,N_10111);
nand U12508 (N_12508,N_10644,N_11264);
nor U12509 (N_12509,N_10388,N_11613);
and U12510 (N_12510,N_10525,N_10747);
or U12511 (N_12511,N_10543,N_10923);
and U12512 (N_12512,N_10456,N_11032);
nor U12513 (N_12513,N_11199,N_11594);
nor U12514 (N_12514,N_11567,N_11867);
nor U12515 (N_12515,N_11636,N_10676);
and U12516 (N_12516,N_11897,N_11302);
and U12517 (N_12517,N_10594,N_11588);
or U12518 (N_12518,N_11721,N_10390);
nor U12519 (N_12519,N_11160,N_11920);
nor U12520 (N_12520,N_10259,N_11394);
or U12521 (N_12521,N_11019,N_11576);
nor U12522 (N_12522,N_10611,N_11587);
nand U12523 (N_12523,N_11509,N_11097);
nand U12524 (N_12524,N_10090,N_10188);
and U12525 (N_12525,N_10439,N_11348);
and U12526 (N_12526,N_11325,N_11706);
nand U12527 (N_12527,N_11916,N_11186);
and U12528 (N_12528,N_11462,N_11082);
nor U12529 (N_12529,N_10651,N_11298);
nand U12530 (N_12530,N_10609,N_10364);
or U12531 (N_12531,N_10545,N_10623);
and U12532 (N_12532,N_11451,N_10498);
and U12533 (N_12533,N_10787,N_10567);
or U12534 (N_12534,N_11424,N_11407);
nor U12535 (N_12535,N_10443,N_11630);
or U12536 (N_12536,N_11401,N_11563);
xnor U12537 (N_12537,N_11868,N_11624);
or U12538 (N_12538,N_10640,N_11575);
or U12539 (N_12539,N_10581,N_11736);
or U12540 (N_12540,N_10092,N_10517);
nor U12541 (N_12541,N_11066,N_11062);
and U12542 (N_12542,N_10041,N_11040);
nor U12543 (N_12543,N_10936,N_10842);
xnor U12544 (N_12544,N_11684,N_10341);
nor U12545 (N_12545,N_10708,N_11106);
or U12546 (N_12546,N_11968,N_11027);
and U12547 (N_12547,N_11681,N_10599);
and U12548 (N_12548,N_10073,N_11773);
and U12549 (N_12549,N_11242,N_10433);
xnor U12550 (N_12550,N_10085,N_10613);
nor U12551 (N_12551,N_11914,N_11796);
nor U12552 (N_12552,N_11668,N_11665);
or U12553 (N_12553,N_11674,N_10254);
and U12554 (N_12554,N_10054,N_10689);
and U12555 (N_12555,N_10514,N_10418);
or U12556 (N_12556,N_11310,N_10634);
and U12557 (N_12557,N_10302,N_10762);
or U12558 (N_12558,N_11045,N_10275);
or U12559 (N_12559,N_11900,N_11763);
and U12560 (N_12560,N_11059,N_11258);
nor U12561 (N_12561,N_10348,N_11560);
or U12562 (N_12562,N_11390,N_10045);
or U12563 (N_12563,N_11917,N_10071);
or U12564 (N_12564,N_10780,N_10057);
and U12565 (N_12565,N_11752,N_11485);
nand U12566 (N_12566,N_11737,N_10156);
and U12567 (N_12567,N_10248,N_11337);
nor U12568 (N_12568,N_11178,N_11368);
nand U12569 (N_12569,N_11021,N_11478);
or U12570 (N_12570,N_10368,N_10163);
and U12571 (N_12571,N_11497,N_11044);
or U12572 (N_12572,N_11573,N_10908);
or U12573 (N_12573,N_10266,N_11582);
and U12574 (N_12574,N_11965,N_11685);
nor U12575 (N_12575,N_10345,N_11101);
nor U12576 (N_12576,N_11166,N_11184);
and U12577 (N_12577,N_10281,N_11574);
and U12578 (N_12578,N_10821,N_10815);
or U12579 (N_12579,N_11285,N_11822);
nand U12580 (N_12580,N_11508,N_10922);
nand U12581 (N_12581,N_11947,N_10946);
or U12582 (N_12582,N_10464,N_10607);
nand U12583 (N_12583,N_11305,N_11140);
or U12584 (N_12584,N_10036,N_11014);
nand U12585 (N_12585,N_10966,N_10106);
and U12586 (N_12586,N_11993,N_11827);
nand U12587 (N_12587,N_10287,N_10856);
nand U12588 (N_12588,N_10680,N_11905);
nand U12589 (N_12589,N_11453,N_11127);
nand U12590 (N_12590,N_11446,N_10841);
or U12591 (N_12591,N_11085,N_11946);
nor U12592 (N_12592,N_10226,N_10244);
or U12593 (N_12593,N_10096,N_11410);
nand U12594 (N_12594,N_11430,N_10854);
nand U12595 (N_12595,N_10050,N_10255);
and U12596 (N_12596,N_10148,N_10769);
and U12597 (N_12597,N_10344,N_11843);
and U12598 (N_12598,N_11507,N_10770);
and U12599 (N_12599,N_10471,N_10492);
nand U12600 (N_12600,N_11353,N_11792);
nor U12601 (N_12601,N_11536,N_10832);
nor U12602 (N_12602,N_11026,N_11849);
nor U12603 (N_12603,N_11945,N_11067);
and U12604 (N_12604,N_11392,N_11537);
nand U12605 (N_12605,N_11423,N_10472);
or U12606 (N_12606,N_11187,N_10487);
or U12607 (N_12607,N_11079,N_11366);
and U12608 (N_12608,N_11103,N_11255);
nor U12609 (N_12609,N_11164,N_10490);
nor U12610 (N_12610,N_10113,N_10192);
nor U12611 (N_12611,N_11246,N_10399);
nand U12612 (N_12612,N_11042,N_11984);
and U12613 (N_12613,N_11970,N_11694);
and U12614 (N_12614,N_11088,N_11384);
nand U12615 (N_12615,N_11833,N_11183);
nand U12616 (N_12616,N_10064,N_11768);
or U12617 (N_12617,N_11071,N_10810);
and U12618 (N_12618,N_11942,N_11248);
nor U12619 (N_12619,N_10181,N_11350);
nor U12620 (N_12620,N_10189,N_10825);
nor U12621 (N_12621,N_11041,N_10479);
or U12622 (N_12622,N_10273,N_11606);
and U12623 (N_12623,N_11069,N_10758);
and U12624 (N_12624,N_10945,N_11675);
and U12625 (N_12625,N_10571,N_11634);
and U12626 (N_12626,N_11168,N_11358);
and U12627 (N_12627,N_11457,N_10549);
nor U12628 (N_12628,N_11961,N_10959);
nand U12629 (N_12629,N_11987,N_11132);
nor U12630 (N_12630,N_10668,N_10186);
nor U12631 (N_12631,N_10754,N_10621);
or U12632 (N_12632,N_11013,N_10573);
nand U12633 (N_12633,N_10377,N_10328);
nand U12634 (N_12634,N_10701,N_11121);
and U12635 (N_12635,N_10900,N_11343);
or U12636 (N_12636,N_11107,N_10089);
nor U12637 (N_12637,N_11950,N_11658);
or U12638 (N_12638,N_11047,N_10819);
and U12639 (N_12639,N_10726,N_10159);
and U12640 (N_12640,N_11830,N_11476);
or U12641 (N_12641,N_11266,N_11175);
and U12642 (N_12642,N_10679,N_10740);
xnor U12643 (N_12643,N_10616,N_11728);
and U12644 (N_12644,N_11873,N_11463);
nand U12645 (N_12645,N_11243,N_10451);
or U12646 (N_12646,N_10428,N_11870);
and U12647 (N_12647,N_11159,N_10116);
and U12648 (N_12648,N_10216,N_11727);
nor U12649 (N_12649,N_10818,N_11196);
and U12650 (N_12650,N_10026,N_10501);
or U12651 (N_12651,N_11194,N_11750);
or U12652 (N_12652,N_11651,N_11891);
nor U12653 (N_12653,N_10779,N_11896);
or U12654 (N_12654,N_10021,N_11114);
nand U12655 (N_12655,N_11386,N_11405);
and U12656 (N_12656,N_11546,N_10595);
nand U12657 (N_12657,N_10334,N_10575);
and U12658 (N_12658,N_10198,N_10117);
nand U12659 (N_12659,N_11090,N_11252);
nand U12660 (N_12660,N_11580,N_11913);
and U12661 (N_12661,N_11116,N_11374);
nand U12662 (N_12662,N_10981,N_10899);
nor U12663 (N_12663,N_10992,N_10690);
or U12664 (N_12664,N_11957,N_11976);
or U12665 (N_12665,N_11486,N_10434);
or U12666 (N_12666,N_10985,N_11131);
nor U12667 (N_12667,N_10949,N_11251);
nand U12668 (N_12668,N_11461,N_10297);
and U12669 (N_12669,N_11915,N_10161);
or U12670 (N_12670,N_10914,N_11769);
nor U12671 (N_12671,N_10824,N_10973);
xor U12672 (N_12672,N_11207,N_11150);
and U12673 (N_12673,N_10058,N_11612);
xnor U12674 (N_12674,N_11875,N_11400);
and U12675 (N_12675,N_11232,N_11260);
and U12676 (N_12676,N_10941,N_11678);
nor U12677 (N_12677,N_11617,N_11230);
nand U12678 (N_12678,N_10805,N_10510);
or U12679 (N_12679,N_10131,N_11320);
and U12680 (N_12680,N_10542,N_11077);
or U12681 (N_12681,N_10744,N_11123);
nand U12682 (N_12682,N_10749,N_11152);
nand U12683 (N_12683,N_10739,N_11240);
or U12684 (N_12684,N_10789,N_11290);
nand U12685 (N_12685,N_11279,N_11614);
nand U12686 (N_12686,N_11826,N_10956);
nand U12687 (N_12687,N_10442,N_10774);
nand U12688 (N_12688,N_10217,N_11418);
nand U12689 (N_12689,N_10586,N_11271);
nor U12690 (N_12690,N_10467,N_10369);
nor U12691 (N_12691,N_11250,N_11771);
nor U12692 (N_12692,N_11585,N_11439);
nor U12693 (N_12693,N_10438,N_11749);
and U12694 (N_12694,N_11048,N_11632);
or U12695 (N_12695,N_10429,N_11813);
and U12696 (N_12696,N_10729,N_10776);
or U12697 (N_12697,N_10801,N_11856);
nand U12698 (N_12698,N_10461,N_10566);
or U12699 (N_12699,N_10136,N_11128);
nand U12700 (N_12700,N_10765,N_10419);
and U12701 (N_12701,N_10742,N_11454);
and U12702 (N_12702,N_11876,N_11741);
or U12703 (N_12703,N_10636,N_10066);
and U12704 (N_12704,N_11068,N_11095);
or U12705 (N_12705,N_10211,N_10518);
nor U12706 (N_12706,N_10761,N_10995);
and U12707 (N_12707,N_10737,N_10752);
or U12708 (N_12708,N_11842,N_10081);
or U12709 (N_12709,N_11098,N_10704);
nor U12710 (N_12710,N_11172,N_11974);
nand U12711 (N_12711,N_11288,N_10221);
or U12712 (N_12712,N_11303,N_10437);
nor U12713 (N_12713,N_11716,N_11256);
nor U12714 (N_12714,N_11173,N_11811);
xnor U12715 (N_12715,N_11391,N_10950);
nand U12716 (N_12716,N_10187,N_11899);
nor U12717 (N_12717,N_11135,N_11118);
or U12718 (N_12718,N_10047,N_10247);
or U12719 (N_12719,N_11185,N_11003);
or U12720 (N_12720,N_11113,N_10493);
nor U12721 (N_12721,N_11001,N_10897);
nor U12722 (N_12722,N_11359,N_11308);
nor U12723 (N_12723,N_11218,N_10962);
nand U12724 (N_12724,N_10829,N_10608);
and U12725 (N_12725,N_10053,N_10098);
and U12726 (N_12726,N_10383,N_10332);
or U12727 (N_12727,N_11104,N_11877);
and U12728 (N_12728,N_11259,N_10695);
nor U12729 (N_12729,N_10110,N_10577);
nor U12730 (N_12730,N_10379,N_11511);
and U12731 (N_12731,N_10748,N_10494);
nand U12732 (N_12732,N_10061,N_10871);
or U12733 (N_12733,N_11616,N_11738);
nand U12734 (N_12734,N_10055,N_10436);
nor U12735 (N_12735,N_10103,N_10678);
nand U12736 (N_12736,N_10425,N_10993);
or U12737 (N_12737,N_11145,N_11998);
or U12738 (N_12738,N_10261,N_11669);
nand U12739 (N_12739,N_10120,N_11689);
and U12740 (N_12740,N_10300,N_10241);
nor U12741 (N_12741,N_10359,N_11517);
or U12742 (N_12742,N_10646,N_11291);
or U12743 (N_12743,N_10180,N_11050);
nor U12744 (N_12744,N_10206,N_11245);
and U12745 (N_12745,N_10210,N_11528);
and U12746 (N_12746,N_10860,N_10813);
or U12747 (N_12747,N_11146,N_10725);
nor U12748 (N_12748,N_11399,N_10637);
and U12749 (N_12749,N_11427,N_10002);
nand U12750 (N_12750,N_11332,N_10199);
xnor U12751 (N_12751,N_10264,N_10446);
nand U12752 (N_12752,N_11715,N_11275);
and U12753 (N_12753,N_10673,N_10008);
nand U12754 (N_12754,N_10902,N_11805);
and U12755 (N_12755,N_11935,N_10507);
or U12756 (N_12756,N_10940,N_10104);
nand U12757 (N_12757,N_10935,N_11762);
and U12758 (N_12758,N_11607,N_11795);
or U12759 (N_12759,N_10682,N_10009);
and U12760 (N_12760,N_11376,N_11406);
or U12761 (N_12761,N_11543,N_11157);
and U12762 (N_12762,N_10219,N_10505);
nand U12763 (N_12763,N_11191,N_11890);
nor U12764 (N_12764,N_11797,N_10546);
nor U12765 (N_12765,N_11236,N_10757);
nor U12766 (N_12766,N_11619,N_11751);
or U12767 (N_12767,N_11369,N_11432);
and U12768 (N_12768,N_10620,N_10938);
xnor U12769 (N_12769,N_10965,N_11435);
nand U12770 (N_12770,N_11631,N_10700);
and U12771 (N_12771,N_11206,N_10257);
nand U12772 (N_12772,N_11198,N_10200);
nand U12773 (N_12773,N_11802,N_10149);
and U12774 (N_12774,N_11941,N_11472);
nor U12775 (N_12775,N_10069,N_10876);
or U12776 (N_12776,N_10531,N_10792);
or U12777 (N_12777,N_10168,N_10735);
nor U12778 (N_12778,N_10183,N_10208);
and U12779 (N_12779,N_10032,N_10094);
nand U12780 (N_12780,N_11263,N_10083);
nand U12781 (N_12781,N_10820,N_11978);
and U12782 (N_12782,N_10589,N_11119);
nor U12783 (N_12783,N_11429,N_11712);
nand U12784 (N_12784,N_11479,N_10723);
or U12785 (N_12785,N_10839,N_10242);
nor U12786 (N_12786,N_11122,N_11278);
and U12787 (N_12787,N_10046,N_10716);
and U12788 (N_12788,N_10398,N_11237);
nand U12789 (N_12789,N_11387,N_11628);
xnor U12790 (N_12790,N_10466,N_10205);
nor U12791 (N_12791,N_10665,N_10756);
and U12792 (N_12792,N_11848,N_11554);
and U12793 (N_12793,N_11503,N_11404);
and U12794 (N_12794,N_11470,N_11409);
nor U12795 (N_12795,N_11985,N_10440);
nor U12796 (N_12796,N_11363,N_10934);
and U12797 (N_12797,N_11934,N_11006);
or U12798 (N_12798,N_10806,N_10715);
nand U12799 (N_12799,N_11141,N_10954);
nand U12800 (N_12800,N_11295,N_10896);
nand U12801 (N_12801,N_11219,N_10772);
nor U12802 (N_12802,N_11880,N_11195);
nor U12803 (N_12803,N_11953,N_11011);
and U12804 (N_12804,N_10112,N_10363);
nand U12805 (N_12805,N_10454,N_11776);
xnor U12806 (N_12806,N_11046,N_11884);
xor U12807 (N_12807,N_10235,N_11943);
and U12808 (N_12808,N_10432,N_11506);
or U12809 (N_12809,N_11996,N_11060);
or U12810 (N_12810,N_11093,N_10552);
nand U12811 (N_12811,N_10080,N_10816);
nand U12812 (N_12812,N_10802,N_11640);
and U12813 (N_12813,N_11417,N_11919);
nor U12814 (N_12814,N_10879,N_11521);
nor U12815 (N_12815,N_10564,N_10001);
nor U12816 (N_12816,N_11981,N_10830);
or U12817 (N_12817,N_10837,N_10910);
or U12818 (N_12818,N_10751,N_10150);
and U12819 (N_12819,N_10719,N_10114);
or U12820 (N_12820,N_11031,N_11273);
nand U12821 (N_12821,N_10202,N_11673);
and U12822 (N_12822,N_10605,N_11526);
and U12823 (N_12823,N_10074,N_10601);
and U12824 (N_12824,N_10790,N_11489);
nand U12825 (N_12825,N_10763,N_11609);
nor U12826 (N_12826,N_10976,N_10588);
and U12827 (N_12827,N_11365,N_11804);
nand U12828 (N_12828,N_11761,N_11491);
nand U12829 (N_12829,N_10677,N_10000);
and U12830 (N_12830,N_11682,N_10289);
nand U12831 (N_12831,N_11442,N_11703);
nor U12832 (N_12832,N_10304,N_11865);
or U12833 (N_12833,N_11988,N_10509);
and U12834 (N_12834,N_11272,N_11083);
nor U12835 (N_12835,N_11936,N_11825);
or U12836 (N_12836,N_11569,N_10760);
and U12837 (N_12837,N_11227,N_10629);
nand U12838 (N_12838,N_10838,N_10528);
nand U12839 (N_12839,N_11336,N_11823);
or U12840 (N_12840,N_11638,N_10833);
nor U12841 (N_12841,N_10068,N_10570);
and U12842 (N_12842,N_10059,N_11739);
or U12843 (N_12843,N_11402,N_10151);
nor U12844 (N_12844,N_10474,N_10179);
and U12845 (N_12845,N_11553,N_11835);
nor U12846 (N_12846,N_10469,N_10338);
nor U12847 (N_12847,N_11649,N_10692);
nand U12848 (N_12848,N_11789,N_10251);
and U12849 (N_12849,N_11820,N_11319);
xnor U12850 (N_12850,N_10218,N_10099);
nor U12851 (N_12851,N_11341,N_10410);
nand U12852 (N_12852,N_10901,N_10356);
nand U12853 (N_12853,N_10323,N_10631);
or U12854 (N_12854,N_10996,N_11967);
nor U12855 (N_12855,N_10246,N_11466);
and U12856 (N_12856,N_10986,N_11901);
nor U12857 (N_12857,N_11787,N_10933);
nor U12858 (N_12858,N_10293,N_10229);
xnor U12859 (N_12859,N_11473,N_11729);
nand U12860 (N_12860,N_11324,N_10299);
nand U12861 (N_12861,N_10538,N_11222);
and U12862 (N_12862,N_11747,N_11471);
and U12863 (N_12863,N_11139,N_10357);
nor U12864 (N_12864,N_10164,N_11373);
and U12865 (N_12865,N_11177,N_10576);
or U12866 (N_12866,N_10508,N_10417);
or U12867 (N_12867,N_11233,N_10745);
nor U12868 (N_12868,N_10124,N_11239);
or U12869 (N_12869,N_10018,N_11529);
nor U12870 (N_12870,N_11448,N_10038);
and U12871 (N_12871,N_10010,N_10118);
nand U12872 (N_12872,N_10969,N_10329);
or U12873 (N_12873,N_10401,N_10318);
nor U12874 (N_12874,N_10462,N_10738);
and U12875 (N_12875,N_11717,N_11637);
and U12876 (N_12876,N_10314,N_11038);
nor U12877 (N_12877,N_10178,N_10182);
nor U12878 (N_12878,N_11020,N_10635);
nor U12879 (N_12879,N_11347,N_10166);
or U12880 (N_12880,N_11932,N_11709);
and U12881 (N_12881,N_11878,N_11540);
nor U12882 (N_12882,N_10982,N_10448);
nand U12883 (N_12883,N_11482,N_11642);
nor U12884 (N_12884,N_11280,N_10126);
or U12885 (N_12885,N_10557,N_11798);
nor U12886 (N_12886,N_11837,N_10919);
nand U12887 (N_12887,N_11928,N_10145);
and U12888 (N_12888,N_11257,N_10342);
or U12889 (N_12889,N_11452,N_11539);
or U12890 (N_12890,N_10063,N_11147);
nand U12891 (N_12891,N_11455,N_11504);
nor U12892 (N_12892,N_11501,N_11687);
nor U12893 (N_12893,N_10051,N_11831);
or U12894 (N_12894,N_11562,N_11355);
or U12895 (N_12895,N_11982,N_11235);
nand U12896 (N_12896,N_11188,N_10622);
nand U12897 (N_12897,N_11338,N_11778);
nor U12898 (N_12898,N_10859,N_10732);
nand U12899 (N_12899,N_11110,N_11226);
and U12900 (N_12900,N_10722,N_11661);
nor U12901 (N_12901,N_11054,N_10201);
or U12902 (N_12902,N_11817,N_10648);
nand U12903 (N_12903,N_11534,N_10102);
nor U12904 (N_12904,N_11241,N_10042);
nand U12905 (N_12905,N_10135,N_10352);
nand U12906 (N_12906,N_11912,N_10237);
or U12907 (N_12907,N_11641,N_10633);
and U12908 (N_12908,N_11468,N_10315);
and U12909 (N_12909,N_10385,N_11216);
and U12910 (N_12910,N_10983,N_10537);
and U12911 (N_12911,N_11881,N_10052);
and U12912 (N_12912,N_11327,N_10688);
nor U12913 (N_12913,N_11335,N_11611);
and U12914 (N_12914,N_10430,N_11133);
and U12915 (N_12915,N_11834,N_11991);
nor U12916 (N_12916,N_10316,N_10301);
and U12917 (N_12917,N_11645,N_10515);
or U12918 (N_12918,N_11434,N_10617);
nand U12919 (N_12919,N_11174,N_10288);
nor U12920 (N_12920,N_11572,N_10592);
nand U12921 (N_12921,N_10775,N_11039);
and U12922 (N_12922,N_10811,N_10707);
nor U12923 (N_12923,N_10489,N_11704);
and U12924 (N_12924,N_10023,N_11070);
or U12925 (N_12925,N_10133,N_11660);
or U12926 (N_12926,N_11117,N_11921);
nand U12927 (N_12927,N_10674,N_11346);
nand U12928 (N_12928,N_10685,N_10278);
nand U12929 (N_12929,N_10263,N_11004);
and U12930 (N_12930,N_10666,N_11610);
nand U12931 (N_12931,N_10365,N_11428);
and U12932 (N_12932,N_10067,N_10194);
nor U12933 (N_12933,N_10683,N_10373);
or U12934 (N_12934,N_11481,N_11099);
or U12935 (N_12935,N_10706,N_11247);
nand U12936 (N_12936,N_11800,N_11200);
nand U12937 (N_12937,N_10160,N_11221);
nor U12938 (N_12938,N_10887,N_11903);
or U12939 (N_12939,N_11620,N_10320);
or U12940 (N_12940,N_10340,N_10975);
nand U12941 (N_12941,N_10394,N_11911);
or U12942 (N_12942,N_11033,N_10366);
nand U12943 (N_12943,N_11564,N_11522);
and U12944 (N_12944,N_10788,N_11388);
or U12945 (N_12945,N_11277,N_10005);
nand U12946 (N_12946,N_11918,N_10733);
and U12947 (N_12947,N_11313,N_10028);
nor U12948 (N_12948,N_11382,N_10652);
nand U12949 (N_12949,N_11456,N_11323);
and U12950 (N_12950,N_10931,N_11274);
or U12951 (N_12951,N_10523,N_10153);
nor U12952 (N_12952,N_11853,N_11758);
and U12953 (N_12953,N_10335,N_10203);
nand U12954 (N_12954,N_11851,N_10602);
nand U12955 (N_12955,N_11670,N_11599);
nor U12956 (N_12956,N_11007,N_11450);
nand U12957 (N_12957,N_11959,N_10184);
nor U12958 (N_12958,N_11861,N_11449);
nand U12959 (N_12959,N_11701,N_11129);
and U12960 (N_12960,N_10539,N_10878);
or U12961 (N_12961,N_11413,N_11648);
nand U12962 (N_12962,N_11680,N_10883);
and U12963 (N_12963,N_10921,N_11929);
nor U12964 (N_12964,N_10628,N_11535);
nor U12965 (N_12965,N_11075,N_10122);
nor U12966 (N_12966,N_11846,N_10019);
or U12967 (N_12967,N_11294,N_11692);
and U12968 (N_12968,N_10459,N_10784);
or U12969 (N_12969,N_10478,N_11971);
and U12970 (N_12970,N_10372,N_10413);
nand U12971 (N_12971,N_11136,N_10078);
nor U12972 (N_12972,N_11025,N_10409);
or U12973 (N_12973,N_10835,N_11815);
nand U12974 (N_12974,N_10070,N_10988);
nor U12975 (N_12975,N_10427,N_10407);
and U12976 (N_12976,N_11558,N_11847);
or U12977 (N_12977,N_11948,N_10322);
and U12978 (N_12978,N_10171,N_11532);
or U12979 (N_12979,N_11590,N_10091);
nand U12980 (N_12980,N_11371,N_11138);
and U12981 (N_12981,N_10978,N_11036);
or U12982 (N_12982,N_11958,N_11398);
and U12983 (N_12983,N_11009,N_11217);
nand U12984 (N_12984,N_10197,N_11352);
and U12985 (N_12985,N_11315,N_10684);
nor U12986 (N_12986,N_10786,N_11810);
or U12987 (N_12987,N_10785,N_10989);
nor U12988 (N_12988,N_10351,N_10283);
nor U12989 (N_12989,N_11894,N_10843);
and U12990 (N_12990,N_10730,N_11224);
xnor U12991 (N_12991,N_10596,N_10653);
or U12992 (N_12992,N_10400,N_11267);
nand U12993 (N_12993,N_10699,N_11330);
nor U12994 (N_12994,N_11464,N_10044);
or U12995 (N_12995,N_11268,N_10486);
nand U12996 (N_12996,N_11156,N_11345);
and U12997 (N_12997,N_11702,N_10650);
nand U12998 (N_12998,N_10587,N_10553);
nand U12999 (N_12999,N_10040,N_10781);
or U13000 (N_13000,N_10661,N_11580);
or U13001 (N_13001,N_11982,N_11311);
nand U13002 (N_13002,N_10422,N_10675);
nand U13003 (N_13003,N_11514,N_10321);
or U13004 (N_13004,N_11715,N_10097);
nor U13005 (N_13005,N_10059,N_10323);
nor U13006 (N_13006,N_10373,N_10570);
nand U13007 (N_13007,N_11786,N_11825);
nand U13008 (N_13008,N_10434,N_10624);
nand U13009 (N_13009,N_10135,N_11389);
nand U13010 (N_13010,N_11711,N_10281);
or U13011 (N_13011,N_10429,N_10687);
or U13012 (N_13012,N_10569,N_10505);
nand U13013 (N_13013,N_11775,N_11029);
nand U13014 (N_13014,N_10156,N_10836);
and U13015 (N_13015,N_10737,N_11728);
nor U13016 (N_13016,N_10271,N_11691);
or U13017 (N_13017,N_11630,N_11491);
nand U13018 (N_13018,N_10890,N_11498);
nand U13019 (N_13019,N_10055,N_11046);
or U13020 (N_13020,N_10153,N_10808);
nand U13021 (N_13021,N_10951,N_11635);
and U13022 (N_13022,N_11429,N_10302);
nand U13023 (N_13023,N_10266,N_11297);
or U13024 (N_13024,N_10857,N_11979);
and U13025 (N_13025,N_10937,N_11246);
nand U13026 (N_13026,N_11460,N_10514);
or U13027 (N_13027,N_11250,N_10120);
and U13028 (N_13028,N_10760,N_11164);
nand U13029 (N_13029,N_10794,N_11682);
or U13030 (N_13030,N_10823,N_11595);
and U13031 (N_13031,N_10302,N_11172);
and U13032 (N_13032,N_11431,N_11803);
nor U13033 (N_13033,N_10123,N_11415);
nor U13034 (N_13034,N_10846,N_11143);
nand U13035 (N_13035,N_11741,N_11531);
nor U13036 (N_13036,N_10252,N_10322);
and U13037 (N_13037,N_11126,N_11204);
or U13038 (N_13038,N_10135,N_11634);
nand U13039 (N_13039,N_10934,N_10464);
nor U13040 (N_13040,N_11642,N_11647);
nand U13041 (N_13041,N_10030,N_11077);
and U13042 (N_13042,N_11180,N_11109);
nand U13043 (N_13043,N_11180,N_10189);
nor U13044 (N_13044,N_10825,N_11275);
nor U13045 (N_13045,N_10080,N_11804);
nor U13046 (N_13046,N_11897,N_11960);
nor U13047 (N_13047,N_11031,N_10800);
or U13048 (N_13048,N_10586,N_10493);
nand U13049 (N_13049,N_10320,N_10851);
and U13050 (N_13050,N_10569,N_11582);
or U13051 (N_13051,N_10386,N_10558);
and U13052 (N_13052,N_11213,N_11433);
nand U13053 (N_13053,N_10661,N_11310);
nor U13054 (N_13054,N_11232,N_11767);
or U13055 (N_13055,N_11922,N_10424);
nand U13056 (N_13056,N_11669,N_11163);
or U13057 (N_13057,N_10139,N_11514);
xor U13058 (N_13058,N_11704,N_11196);
or U13059 (N_13059,N_11941,N_10964);
nor U13060 (N_13060,N_11765,N_10752);
and U13061 (N_13061,N_10261,N_10410);
and U13062 (N_13062,N_10911,N_10135);
nand U13063 (N_13063,N_10400,N_10530);
nand U13064 (N_13064,N_11791,N_10616);
or U13065 (N_13065,N_10327,N_11947);
nor U13066 (N_13066,N_10869,N_10454);
or U13067 (N_13067,N_10429,N_10262);
nor U13068 (N_13068,N_10901,N_10382);
nor U13069 (N_13069,N_11620,N_11184);
nand U13070 (N_13070,N_11417,N_10085);
nand U13071 (N_13071,N_11471,N_10646);
nand U13072 (N_13072,N_11705,N_11508);
nand U13073 (N_13073,N_11106,N_10763);
nand U13074 (N_13074,N_11850,N_11899);
nand U13075 (N_13075,N_10830,N_10198);
nor U13076 (N_13076,N_11376,N_11194);
or U13077 (N_13077,N_11643,N_10019);
or U13078 (N_13078,N_10214,N_10494);
nor U13079 (N_13079,N_11007,N_10527);
and U13080 (N_13080,N_10553,N_11074);
nand U13081 (N_13081,N_10583,N_11763);
nand U13082 (N_13082,N_11627,N_10171);
and U13083 (N_13083,N_10682,N_10161);
nor U13084 (N_13084,N_11081,N_11838);
nand U13085 (N_13085,N_11753,N_10895);
nor U13086 (N_13086,N_11134,N_10640);
or U13087 (N_13087,N_10696,N_11309);
and U13088 (N_13088,N_11044,N_11024);
nand U13089 (N_13089,N_10732,N_11356);
nand U13090 (N_13090,N_11224,N_10197);
nand U13091 (N_13091,N_10908,N_11956);
or U13092 (N_13092,N_11985,N_10749);
or U13093 (N_13093,N_11950,N_10569);
and U13094 (N_13094,N_11062,N_11324);
nor U13095 (N_13095,N_10883,N_10427);
nand U13096 (N_13096,N_11690,N_11148);
nor U13097 (N_13097,N_11998,N_10752);
nor U13098 (N_13098,N_10379,N_11050);
or U13099 (N_13099,N_11429,N_10903);
nor U13100 (N_13100,N_10866,N_10634);
nand U13101 (N_13101,N_11571,N_11293);
or U13102 (N_13102,N_11716,N_10179);
or U13103 (N_13103,N_10028,N_11303);
nand U13104 (N_13104,N_10877,N_11603);
nand U13105 (N_13105,N_10898,N_10126);
or U13106 (N_13106,N_10821,N_10122);
and U13107 (N_13107,N_10077,N_10178);
or U13108 (N_13108,N_10658,N_11670);
nand U13109 (N_13109,N_10879,N_11239);
and U13110 (N_13110,N_10938,N_11365);
nand U13111 (N_13111,N_11724,N_10031);
nand U13112 (N_13112,N_10718,N_10442);
nand U13113 (N_13113,N_11155,N_11044);
nand U13114 (N_13114,N_10446,N_10230);
or U13115 (N_13115,N_10138,N_10750);
nand U13116 (N_13116,N_10732,N_11420);
and U13117 (N_13117,N_11211,N_11621);
nand U13118 (N_13118,N_10995,N_10164);
or U13119 (N_13119,N_11961,N_11968);
or U13120 (N_13120,N_11594,N_11762);
and U13121 (N_13121,N_11049,N_11883);
nand U13122 (N_13122,N_11086,N_10003);
or U13123 (N_13123,N_11403,N_10333);
or U13124 (N_13124,N_10439,N_10550);
nor U13125 (N_13125,N_11453,N_10193);
or U13126 (N_13126,N_11389,N_11508);
nor U13127 (N_13127,N_11242,N_11396);
or U13128 (N_13128,N_11783,N_10534);
nand U13129 (N_13129,N_11496,N_10142);
nor U13130 (N_13130,N_11579,N_10099);
nand U13131 (N_13131,N_11303,N_10679);
or U13132 (N_13132,N_10368,N_10889);
nor U13133 (N_13133,N_11247,N_10571);
nand U13134 (N_13134,N_10739,N_10156);
xor U13135 (N_13135,N_11802,N_11712);
nor U13136 (N_13136,N_11098,N_11778);
nor U13137 (N_13137,N_11145,N_10307);
and U13138 (N_13138,N_10362,N_10242);
and U13139 (N_13139,N_11835,N_11691);
nor U13140 (N_13140,N_10254,N_10760);
nand U13141 (N_13141,N_11666,N_10925);
nand U13142 (N_13142,N_10398,N_11108);
and U13143 (N_13143,N_11088,N_10130);
nor U13144 (N_13144,N_10173,N_11026);
or U13145 (N_13145,N_10367,N_11433);
nor U13146 (N_13146,N_11627,N_11632);
and U13147 (N_13147,N_11486,N_10890);
nand U13148 (N_13148,N_10962,N_11968);
nand U13149 (N_13149,N_10256,N_11695);
nand U13150 (N_13150,N_10932,N_10463);
or U13151 (N_13151,N_11702,N_11275);
or U13152 (N_13152,N_10562,N_11481);
or U13153 (N_13153,N_10743,N_11869);
and U13154 (N_13154,N_10877,N_11729);
nand U13155 (N_13155,N_11108,N_10029);
xor U13156 (N_13156,N_10469,N_11203);
nor U13157 (N_13157,N_11759,N_11571);
and U13158 (N_13158,N_10746,N_11042);
or U13159 (N_13159,N_11722,N_11855);
or U13160 (N_13160,N_11688,N_11394);
nor U13161 (N_13161,N_10598,N_10967);
or U13162 (N_13162,N_11490,N_10734);
nand U13163 (N_13163,N_10886,N_11291);
or U13164 (N_13164,N_11229,N_11562);
and U13165 (N_13165,N_10546,N_10052);
nor U13166 (N_13166,N_10470,N_11921);
or U13167 (N_13167,N_10177,N_10865);
or U13168 (N_13168,N_11741,N_11997);
nand U13169 (N_13169,N_11496,N_11531);
and U13170 (N_13170,N_10275,N_10095);
or U13171 (N_13171,N_10903,N_10803);
nand U13172 (N_13172,N_10970,N_11967);
nor U13173 (N_13173,N_10158,N_10885);
and U13174 (N_13174,N_11041,N_11782);
or U13175 (N_13175,N_11645,N_10683);
or U13176 (N_13176,N_11755,N_11943);
nand U13177 (N_13177,N_10607,N_11262);
or U13178 (N_13178,N_11925,N_10526);
and U13179 (N_13179,N_11637,N_11167);
nand U13180 (N_13180,N_11656,N_11519);
and U13181 (N_13181,N_11951,N_11490);
nor U13182 (N_13182,N_10935,N_11881);
or U13183 (N_13183,N_11698,N_11737);
or U13184 (N_13184,N_11624,N_10068);
nand U13185 (N_13185,N_10727,N_10676);
nor U13186 (N_13186,N_10704,N_10250);
nor U13187 (N_13187,N_11590,N_11715);
or U13188 (N_13188,N_10627,N_10473);
nand U13189 (N_13189,N_11176,N_10880);
and U13190 (N_13190,N_10103,N_10084);
or U13191 (N_13191,N_11194,N_10886);
xnor U13192 (N_13192,N_10870,N_11155);
xnor U13193 (N_13193,N_10133,N_11417);
and U13194 (N_13194,N_11619,N_10465);
nor U13195 (N_13195,N_11116,N_10290);
nor U13196 (N_13196,N_11178,N_11386);
or U13197 (N_13197,N_10925,N_10450);
or U13198 (N_13198,N_11925,N_10899);
or U13199 (N_13199,N_10350,N_11285);
and U13200 (N_13200,N_11810,N_10102);
and U13201 (N_13201,N_10924,N_10653);
nor U13202 (N_13202,N_11390,N_11844);
and U13203 (N_13203,N_10731,N_11881);
or U13204 (N_13204,N_10144,N_11898);
nand U13205 (N_13205,N_10359,N_10748);
and U13206 (N_13206,N_10402,N_10186);
and U13207 (N_13207,N_10315,N_10736);
nand U13208 (N_13208,N_10320,N_11924);
or U13209 (N_13209,N_10597,N_11547);
or U13210 (N_13210,N_11752,N_10277);
and U13211 (N_13211,N_11811,N_11577);
or U13212 (N_13212,N_10930,N_10836);
nand U13213 (N_13213,N_10608,N_10349);
or U13214 (N_13214,N_11902,N_10894);
nand U13215 (N_13215,N_11679,N_10293);
nor U13216 (N_13216,N_10212,N_11522);
and U13217 (N_13217,N_11130,N_10837);
nand U13218 (N_13218,N_11661,N_11396);
or U13219 (N_13219,N_11286,N_10531);
or U13220 (N_13220,N_11200,N_11516);
or U13221 (N_13221,N_11457,N_11791);
and U13222 (N_13222,N_11641,N_11675);
nand U13223 (N_13223,N_10392,N_10764);
or U13224 (N_13224,N_11774,N_11084);
nor U13225 (N_13225,N_11488,N_10580);
and U13226 (N_13226,N_11244,N_11364);
or U13227 (N_13227,N_11676,N_11222);
or U13228 (N_13228,N_10600,N_10737);
nand U13229 (N_13229,N_11109,N_10607);
or U13230 (N_13230,N_11097,N_10047);
nor U13231 (N_13231,N_10330,N_10173);
nand U13232 (N_13232,N_11983,N_10484);
nor U13233 (N_13233,N_11386,N_11966);
and U13234 (N_13234,N_10617,N_11891);
or U13235 (N_13235,N_11117,N_10220);
nand U13236 (N_13236,N_10399,N_11156);
or U13237 (N_13237,N_11559,N_10795);
nand U13238 (N_13238,N_11760,N_11198);
nand U13239 (N_13239,N_10472,N_10850);
nand U13240 (N_13240,N_10633,N_11842);
or U13241 (N_13241,N_11345,N_10025);
nor U13242 (N_13242,N_11083,N_11628);
and U13243 (N_13243,N_11002,N_11000);
nand U13244 (N_13244,N_10242,N_11778);
or U13245 (N_13245,N_11966,N_10162);
nor U13246 (N_13246,N_10023,N_10878);
or U13247 (N_13247,N_11907,N_11499);
or U13248 (N_13248,N_11327,N_10775);
nor U13249 (N_13249,N_11371,N_11230);
and U13250 (N_13250,N_11653,N_11732);
nand U13251 (N_13251,N_11649,N_10402);
and U13252 (N_13252,N_11961,N_10697);
nor U13253 (N_13253,N_11138,N_11298);
or U13254 (N_13254,N_11450,N_10789);
or U13255 (N_13255,N_11109,N_10052);
or U13256 (N_13256,N_10058,N_11013);
or U13257 (N_13257,N_10666,N_10081);
and U13258 (N_13258,N_10958,N_10987);
nand U13259 (N_13259,N_11442,N_10422);
nor U13260 (N_13260,N_10559,N_11142);
and U13261 (N_13261,N_11459,N_11854);
or U13262 (N_13262,N_10509,N_10223);
nor U13263 (N_13263,N_11088,N_11358);
nor U13264 (N_13264,N_11946,N_10121);
nand U13265 (N_13265,N_11138,N_11008);
nand U13266 (N_13266,N_10663,N_11487);
nor U13267 (N_13267,N_11505,N_10941);
nand U13268 (N_13268,N_11397,N_10053);
nand U13269 (N_13269,N_11744,N_10824);
or U13270 (N_13270,N_10778,N_10920);
or U13271 (N_13271,N_11070,N_10876);
nand U13272 (N_13272,N_11670,N_11618);
nand U13273 (N_13273,N_11361,N_10970);
nand U13274 (N_13274,N_10632,N_11454);
nand U13275 (N_13275,N_11980,N_10164);
and U13276 (N_13276,N_11142,N_10314);
nand U13277 (N_13277,N_10668,N_10940);
nor U13278 (N_13278,N_10005,N_11970);
nand U13279 (N_13279,N_11273,N_11458);
nand U13280 (N_13280,N_11150,N_11437);
and U13281 (N_13281,N_11440,N_11435);
nand U13282 (N_13282,N_10126,N_10478);
and U13283 (N_13283,N_10640,N_10964);
or U13284 (N_13284,N_10510,N_11464);
or U13285 (N_13285,N_11648,N_11279);
nand U13286 (N_13286,N_10382,N_11260);
or U13287 (N_13287,N_10891,N_10581);
nand U13288 (N_13288,N_11649,N_11780);
and U13289 (N_13289,N_10884,N_11375);
nor U13290 (N_13290,N_11506,N_10035);
and U13291 (N_13291,N_11429,N_11825);
and U13292 (N_13292,N_10357,N_10161);
or U13293 (N_13293,N_10308,N_10630);
or U13294 (N_13294,N_11149,N_11241);
nor U13295 (N_13295,N_11134,N_11882);
nor U13296 (N_13296,N_10821,N_11508);
nand U13297 (N_13297,N_10523,N_11245);
nand U13298 (N_13298,N_10336,N_11693);
nand U13299 (N_13299,N_10029,N_11838);
nand U13300 (N_13300,N_11301,N_11852);
nor U13301 (N_13301,N_10213,N_11398);
nor U13302 (N_13302,N_11314,N_10218);
or U13303 (N_13303,N_10717,N_11711);
and U13304 (N_13304,N_10977,N_11752);
nand U13305 (N_13305,N_10683,N_11191);
nand U13306 (N_13306,N_11776,N_10405);
nand U13307 (N_13307,N_11786,N_10474);
or U13308 (N_13308,N_11404,N_10048);
nand U13309 (N_13309,N_11809,N_10053);
nor U13310 (N_13310,N_11738,N_10206);
nand U13311 (N_13311,N_11171,N_10654);
nor U13312 (N_13312,N_11125,N_10693);
nand U13313 (N_13313,N_11862,N_11006);
or U13314 (N_13314,N_10996,N_10790);
nor U13315 (N_13315,N_11902,N_11690);
or U13316 (N_13316,N_11942,N_11739);
nor U13317 (N_13317,N_11965,N_11084);
nand U13318 (N_13318,N_11298,N_10792);
or U13319 (N_13319,N_10126,N_11032);
nor U13320 (N_13320,N_10565,N_10276);
nand U13321 (N_13321,N_11632,N_11986);
nor U13322 (N_13322,N_11601,N_11487);
nor U13323 (N_13323,N_11782,N_10923);
nand U13324 (N_13324,N_11060,N_11519);
nor U13325 (N_13325,N_10520,N_11836);
and U13326 (N_13326,N_11560,N_11864);
and U13327 (N_13327,N_10907,N_11985);
and U13328 (N_13328,N_11813,N_10824);
nand U13329 (N_13329,N_11530,N_10460);
nand U13330 (N_13330,N_11827,N_11373);
nor U13331 (N_13331,N_10493,N_11501);
or U13332 (N_13332,N_11672,N_11375);
or U13333 (N_13333,N_11070,N_11732);
nand U13334 (N_13334,N_11319,N_10201);
nand U13335 (N_13335,N_10678,N_10289);
and U13336 (N_13336,N_11226,N_10674);
or U13337 (N_13337,N_10626,N_10200);
and U13338 (N_13338,N_10009,N_11611);
nand U13339 (N_13339,N_11946,N_11119);
nor U13340 (N_13340,N_10034,N_10142);
or U13341 (N_13341,N_10373,N_11073);
and U13342 (N_13342,N_11439,N_11764);
nand U13343 (N_13343,N_10290,N_11089);
and U13344 (N_13344,N_11812,N_10769);
or U13345 (N_13345,N_10846,N_11569);
nor U13346 (N_13346,N_10362,N_10471);
and U13347 (N_13347,N_10183,N_10916);
or U13348 (N_13348,N_11324,N_11722);
nand U13349 (N_13349,N_10597,N_10331);
nor U13350 (N_13350,N_11778,N_10249);
or U13351 (N_13351,N_10643,N_10760);
and U13352 (N_13352,N_10362,N_11312);
and U13353 (N_13353,N_11776,N_10973);
nand U13354 (N_13354,N_10670,N_10209);
nor U13355 (N_13355,N_11828,N_10480);
nand U13356 (N_13356,N_10991,N_11658);
and U13357 (N_13357,N_10413,N_11801);
and U13358 (N_13358,N_11714,N_10907);
and U13359 (N_13359,N_10512,N_10330);
nor U13360 (N_13360,N_10432,N_10533);
nand U13361 (N_13361,N_11085,N_10692);
nand U13362 (N_13362,N_11164,N_11625);
nor U13363 (N_13363,N_10447,N_11519);
nor U13364 (N_13364,N_10958,N_10360);
nand U13365 (N_13365,N_10029,N_11634);
nand U13366 (N_13366,N_11384,N_11783);
nor U13367 (N_13367,N_10901,N_10831);
or U13368 (N_13368,N_10665,N_10361);
nor U13369 (N_13369,N_10456,N_10056);
or U13370 (N_13370,N_10672,N_11481);
nor U13371 (N_13371,N_10860,N_11912);
or U13372 (N_13372,N_11975,N_10089);
nor U13373 (N_13373,N_10895,N_10508);
nand U13374 (N_13374,N_10139,N_10224);
or U13375 (N_13375,N_11372,N_11210);
or U13376 (N_13376,N_11555,N_11455);
nand U13377 (N_13377,N_11568,N_11208);
or U13378 (N_13378,N_11719,N_10583);
nor U13379 (N_13379,N_10770,N_11825);
nand U13380 (N_13380,N_11152,N_11333);
nor U13381 (N_13381,N_10386,N_11552);
nand U13382 (N_13382,N_10828,N_11110);
or U13383 (N_13383,N_10881,N_11458);
nor U13384 (N_13384,N_10539,N_11024);
nor U13385 (N_13385,N_11077,N_11075);
and U13386 (N_13386,N_11983,N_11493);
nand U13387 (N_13387,N_10205,N_11724);
or U13388 (N_13388,N_11591,N_10499);
or U13389 (N_13389,N_11129,N_11298);
or U13390 (N_13390,N_10631,N_11627);
nor U13391 (N_13391,N_10054,N_10568);
or U13392 (N_13392,N_11469,N_10617);
nand U13393 (N_13393,N_10541,N_10695);
nor U13394 (N_13394,N_10741,N_10092);
and U13395 (N_13395,N_10993,N_10837);
nor U13396 (N_13396,N_11828,N_11385);
nand U13397 (N_13397,N_11659,N_10526);
nor U13398 (N_13398,N_10445,N_10221);
nand U13399 (N_13399,N_11039,N_11789);
nand U13400 (N_13400,N_11465,N_11811);
or U13401 (N_13401,N_11762,N_11844);
and U13402 (N_13402,N_10384,N_10306);
nand U13403 (N_13403,N_11377,N_10692);
or U13404 (N_13404,N_10202,N_11614);
or U13405 (N_13405,N_11064,N_11191);
nor U13406 (N_13406,N_10436,N_10999);
nand U13407 (N_13407,N_11488,N_10734);
and U13408 (N_13408,N_10741,N_10992);
nor U13409 (N_13409,N_10598,N_10386);
nand U13410 (N_13410,N_10704,N_10648);
and U13411 (N_13411,N_11238,N_11375);
or U13412 (N_13412,N_11017,N_11554);
and U13413 (N_13413,N_11153,N_11029);
nor U13414 (N_13414,N_11669,N_10218);
nand U13415 (N_13415,N_11586,N_10351);
nand U13416 (N_13416,N_11305,N_10874);
and U13417 (N_13417,N_11005,N_11615);
nor U13418 (N_13418,N_10119,N_10587);
and U13419 (N_13419,N_10824,N_10047);
or U13420 (N_13420,N_11899,N_11173);
or U13421 (N_13421,N_11033,N_10505);
nor U13422 (N_13422,N_10821,N_10937);
nand U13423 (N_13423,N_10505,N_10794);
nand U13424 (N_13424,N_11500,N_11349);
nor U13425 (N_13425,N_11813,N_11219);
xor U13426 (N_13426,N_11353,N_10878);
and U13427 (N_13427,N_11821,N_10537);
or U13428 (N_13428,N_11111,N_10329);
nor U13429 (N_13429,N_10796,N_11706);
or U13430 (N_13430,N_10039,N_10421);
nand U13431 (N_13431,N_11482,N_11735);
and U13432 (N_13432,N_11099,N_11377);
and U13433 (N_13433,N_10449,N_10788);
or U13434 (N_13434,N_11355,N_11922);
or U13435 (N_13435,N_10844,N_10151);
nand U13436 (N_13436,N_10882,N_11040);
and U13437 (N_13437,N_10707,N_11996);
nor U13438 (N_13438,N_10463,N_10484);
nand U13439 (N_13439,N_10584,N_11272);
nor U13440 (N_13440,N_11103,N_10581);
nor U13441 (N_13441,N_10691,N_11079);
nor U13442 (N_13442,N_10970,N_10661);
nand U13443 (N_13443,N_10203,N_11833);
nor U13444 (N_13444,N_11817,N_11975);
or U13445 (N_13445,N_11736,N_11720);
and U13446 (N_13446,N_10710,N_10356);
nor U13447 (N_13447,N_11712,N_10222);
and U13448 (N_13448,N_10607,N_10435);
nand U13449 (N_13449,N_10393,N_10149);
and U13450 (N_13450,N_11038,N_10928);
nand U13451 (N_13451,N_11959,N_10465);
or U13452 (N_13452,N_11804,N_10360);
nor U13453 (N_13453,N_10252,N_10734);
or U13454 (N_13454,N_11211,N_11842);
nor U13455 (N_13455,N_11646,N_10268);
and U13456 (N_13456,N_11240,N_11186);
or U13457 (N_13457,N_10984,N_11628);
nor U13458 (N_13458,N_10205,N_10669);
or U13459 (N_13459,N_10104,N_11183);
nand U13460 (N_13460,N_10410,N_11362);
nand U13461 (N_13461,N_10827,N_10394);
xor U13462 (N_13462,N_11491,N_10895);
and U13463 (N_13463,N_11986,N_10334);
nand U13464 (N_13464,N_10703,N_11178);
or U13465 (N_13465,N_11334,N_11670);
or U13466 (N_13466,N_11260,N_11247);
nor U13467 (N_13467,N_11087,N_10312);
xnor U13468 (N_13468,N_11563,N_11579);
or U13469 (N_13469,N_11450,N_10887);
nor U13470 (N_13470,N_10835,N_10734);
and U13471 (N_13471,N_10506,N_10588);
nor U13472 (N_13472,N_11615,N_11201);
or U13473 (N_13473,N_11547,N_11100);
nand U13474 (N_13474,N_10522,N_10168);
xnor U13475 (N_13475,N_11166,N_11558);
nand U13476 (N_13476,N_10030,N_10232);
nor U13477 (N_13477,N_11362,N_11291);
nand U13478 (N_13478,N_10675,N_10581);
nor U13479 (N_13479,N_11095,N_10086);
nand U13480 (N_13480,N_10288,N_11694);
or U13481 (N_13481,N_11076,N_11501);
nand U13482 (N_13482,N_11468,N_11169);
nand U13483 (N_13483,N_11662,N_11589);
or U13484 (N_13484,N_10236,N_11240);
and U13485 (N_13485,N_11970,N_11531);
nor U13486 (N_13486,N_10669,N_11756);
or U13487 (N_13487,N_10271,N_10033);
nand U13488 (N_13488,N_11380,N_11890);
nand U13489 (N_13489,N_10512,N_11565);
or U13490 (N_13490,N_11857,N_10005);
and U13491 (N_13491,N_10705,N_11026);
or U13492 (N_13492,N_10389,N_10039);
or U13493 (N_13493,N_11619,N_11346);
or U13494 (N_13494,N_11368,N_11626);
nand U13495 (N_13495,N_11548,N_11449);
nand U13496 (N_13496,N_10543,N_11847);
or U13497 (N_13497,N_10318,N_11250);
and U13498 (N_13498,N_10716,N_11455);
nor U13499 (N_13499,N_11839,N_10767);
or U13500 (N_13500,N_11990,N_11415);
nor U13501 (N_13501,N_10368,N_10278);
or U13502 (N_13502,N_11638,N_10601);
nand U13503 (N_13503,N_10761,N_11264);
and U13504 (N_13504,N_11692,N_10828);
and U13505 (N_13505,N_10671,N_11481);
and U13506 (N_13506,N_10185,N_11654);
or U13507 (N_13507,N_10411,N_11110);
or U13508 (N_13508,N_10733,N_10829);
and U13509 (N_13509,N_11833,N_11610);
or U13510 (N_13510,N_10869,N_11971);
or U13511 (N_13511,N_11124,N_11564);
or U13512 (N_13512,N_11359,N_10202);
nor U13513 (N_13513,N_11685,N_10440);
nor U13514 (N_13514,N_10140,N_10805);
nor U13515 (N_13515,N_10988,N_11283);
or U13516 (N_13516,N_10593,N_11297);
and U13517 (N_13517,N_10917,N_11577);
or U13518 (N_13518,N_11977,N_11674);
nand U13519 (N_13519,N_10189,N_11725);
nor U13520 (N_13520,N_11325,N_11375);
or U13521 (N_13521,N_10589,N_10242);
nand U13522 (N_13522,N_10475,N_11261);
xor U13523 (N_13523,N_11134,N_10394);
and U13524 (N_13524,N_10572,N_11593);
and U13525 (N_13525,N_11859,N_10805);
nand U13526 (N_13526,N_10864,N_10661);
or U13527 (N_13527,N_11247,N_11771);
xnor U13528 (N_13528,N_11349,N_11887);
xor U13529 (N_13529,N_10990,N_11339);
nor U13530 (N_13530,N_10070,N_10842);
and U13531 (N_13531,N_10784,N_11055);
nor U13532 (N_13532,N_11841,N_11009);
xor U13533 (N_13533,N_11742,N_10970);
nor U13534 (N_13534,N_10482,N_11921);
or U13535 (N_13535,N_10364,N_11625);
nand U13536 (N_13536,N_10547,N_11987);
or U13537 (N_13537,N_10810,N_10423);
and U13538 (N_13538,N_11702,N_11164);
or U13539 (N_13539,N_11918,N_11007);
xor U13540 (N_13540,N_10267,N_11562);
or U13541 (N_13541,N_11154,N_11446);
nand U13542 (N_13542,N_11156,N_10286);
and U13543 (N_13543,N_10975,N_11165);
or U13544 (N_13544,N_11206,N_10879);
xor U13545 (N_13545,N_11307,N_11377);
nand U13546 (N_13546,N_11043,N_10998);
or U13547 (N_13547,N_10817,N_11339);
nor U13548 (N_13548,N_11643,N_10817);
or U13549 (N_13549,N_10536,N_10494);
nand U13550 (N_13550,N_10297,N_10239);
or U13551 (N_13551,N_11303,N_11523);
nand U13552 (N_13552,N_10611,N_10539);
or U13553 (N_13553,N_11717,N_10588);
nand U13554 (N_13554,N_10046,N_11362);
nor U13555 (N_13555,N_10239,N_11924);
and U13556 (N_13556,N_10050,N_10982);
nor U13557 (N_13557,N_10541,N_10288);
nor U13558 (N_13558,N_11797,N_11868);
and U13559 (N_13559,N_10291,N_11424);
nand U13560 (N_13560,N_11328,N_10249);
and U13561 (N_13561,N_10239,N_10775);
nand U13562 (N_13562,N_10881,N_10642);
and U13563 (N_13563,N_11751,N_11504);
nand U13564 (N_13564,N_11543,N_11217);
nand U13565 (N_13565,N_10805,N_10606);
nand U13566 (N_13566,N_10143,N_10974);
nor U13567 (N_13567,N_11713,N_11426);
or U13568 (N_13568,N_11785,N_11991);
and U13569 (N_13569,N_10660,N_10558);
and U13570 (N_13570,N_10269,N_11765);
nor U13571 (N_13571,N_10695,N_10360);
nor U13572 (N_13572,N_11375,N_11017);
and U13573 (N_13573,N_10725,N_11016);
nor U13574 (N_13574,N_10215,N_10180);
and U13575 (N_13575,N_11587,N_11861);
nor U13576 (N_13576,N_10851,N_11158);
nor U13577 (N_13577,N_11976,N_11696);
or U13578 (N_13578,N_10466,N_10976);
and U13579 (N_13579,N_11572,N_10399);
and U13580 (N_13580,N_10555,N_11684);
nor U13581 (N_13581,N_11163,N_10859);
or U13582 (N_13582,N_10946,N_10165);
and U13583 (N_13583,N_11501,N_11084);
or U13584 (N_13584,N_10990,N_11431);
nor U13585 (N_13585,N_11037,N_10610);
and U13586 (N_13586,N_11983,N_10349);
nand U13587 (N_13587,N_11695,N_11796);
or U13588 (N_13588,N_10908,N_11304);
and U13589 (N_13589,N_11116,N_10771);
nand U13590 (N_13590,N_10992,N_11974);
nor U13591 (N_13591,N_10822,N_10671);
or U13592 (N_13592,N_10783,N_11860);
nand U13593 (N_13593,N_11580,N_10810);
and U13594 (N_13594,N_11729,N_10557);
and U13595 (N_13595,N_11323,N_11080);
nand U13596 (N_13596,N_11661,N_11543);
nor U13597 (N_13597,N_11047,N_11690);
nor U13598 (N_13598,N_10964,N_10878);
or U13599 (N_13599,N_11400,N_10629);
nor U13600 (N_13600,N_10938,N_10283);
nor U13601 (N_13601,N_10373,N_10751);
nand U13602 (N_13602,N_11994,N_11559);
nand U13603 (N_13603,N_11076,N_10169);
nand U13604 (N_13604,N_11143,N_10800);
nand U13605 (N_13605,N_10639,N_11225);
or U13606 (N_13606,N_10949,N_11950);
and U13607 (N_13607,N_11880,N_11231);
or U13608 (N_13608,N_10395,N_10023);
and U13609 (N_13609,N_10774,N_10909);
nand U13610 (N_13610,N_11400,N_11734);
nor U13611 (N_13611,N_10477,N_10928);
nor U13612 (N_13612,N_11366,N_11282);
nand U13613 (N_13613,N_10846,N_10378);
nor U13614 (N_13614,N_10056,N_10104);
nor U13615 (N_13615,N_10318,N_10495);
and U13616 (N_13616,N_10404,N_10124);
nor U13617 (N_13617,N_11493,N_11070);
or U13618 (N_13618,N_10779,N_10863);
nand U13619 (N_13619,N_11859,N_11680);
and U13620 (N_13620,N_11518,N_10606);
or U13621 (N_13621,N_10517,N_10934);
and U13622 (N_13622,N_11316,N_10507);
nor U13623 (N_13623,N_10490,N_10241);
or U13624 (N_13624,N_11768,N_11909);
nand U13625 (N_13625,N_10119,N_10665);
nor U13626 (N_13626,N_11743,N_11057);
or U13627 (N_13627,N_11002,N_11603);
nor U13628 (N_13628,N_11855,N_11073);
and U13629 (N_13629,N_11381,N_10128);
or U13630 (N_13630,N_10612,N_10876);
nand U13631 (N_13631,N_11879,N_11073);
and U13632 (N_13632,N_10911,N_10174);
nor U13633 (N_13633,N_10421,N_10593);
nand U13634 (N_13634,N_11756,N_11440);
and U13635 (N_13635,N_11251,N_11249);
nand U13636 (N_13636,N_11542,N_11349);
nor U13637 (N_13637,N_11162,N_11640);
nand U13638 (N_13638,N_11780,N_10268);
nor U13639 (N_13639,N_11516,N_10519);
nand U13640 (N_13640,N_10645,N_11278);
xnor U13641 (N_13641,N_10075,N_10001);
or U13642 (N_13642,N_11835,N_11970);
nor U13643 (N_13643,N_11054,N_10221);
nor U13644 (N_13644,N_10695,N_11612);
or U13645 (N_13645,N_11669,N_11688);
nor U13646 (N_13646,N_11528,N_10337);
or U13647 (N_13647,N_11560,N_10857);
or U13648 (N_13648,N_11117,N_10267);
or U13649 (N_13649,N_11107,N_11783);
nand U13650 (N_13650,N_10728,N_11110);
and U13651 (N_13651,N_10381,N_11523);
or U13652 (N_13652,N_10206,N_11244);
nor U13653 (N_13653,N_10602,N_11411);
and U13654 (N_13654,N_10235,N_11599);
nand U13655 (N_13655,N_11892,N_10518);
nand U13656 (N_13656,N_11630,N_10921);
nor U13657 (N_13657,N_11980,N_11583);
xor U13658 (N_13658,N_11242,N_10114);
or U13659 (N_13659,N_11142,N_10750);
nand U13660 (N_13660,N_10884,N_11742);
and U13661 (N_13661,N_10138,N_11847);
nand U13662 (N_13662,N_11095,N_11770);
or U13663 (N_13663,N_10373,N_10138);
nor U13664 (N_13664,N_11432,N_11406);
nor U13665 (N_13665,N_11218,N_11995);
or U13666 (N_13666,N_11231,N_10863);
nor U13667 (N_13667,N_11916,N_11943);
nor U13668 (N_13668,N_11766,N_10019);
nor U13669 (N_13669,N_10738,N_10940);
nor U13670 (N_13670,N_11620,N_10722);
and U13671 (N_13671,N_10986,N_11151);
or U13672 (N_13672,N_11239,N_10692);
nand U13673 (N_13673,N_11820,N_10814);
nor U13674 (N_13674,N_11509,N_10094);
nor U13675 (N_13675,N_10343,N_11919);
and U13676 (N_13676,N_11671,N_10352);
or U13677 (N_13677,N_11816,N_11608);
nor U13678 (N_13678,N_10643,N_11076);
or U13679 (N_13679,N_10545,N_11093);
and U13680 (N_13680,N_11173,N_10240);
and U13681 (N_13681,N_11132,N_10647);
nand U13682 (N_13682,N_11511,N_11278);
or U13683 (N_13683,N_10260,N_10909);
or U13684 (N_13684,N_10216,N_11267);
nor U13685 (N_13685,N_11337,N_11631);
nand U13686 (N_13686,N_11786,N_11761);
nand U13687 (N_13687,N_11188,N_11322);
nand U13688 (N_13688,N_10548,N_10417);
or U13689 (N_13689,N_11981,N_10710);
nand U13690 (N_13690,N_11769,N_11045);
nand U13691 (N_13691,N_11978,N_10478);
and U13692 (N_13692,N_11879,N_10224);
or U13693 (N_13693,N_11256,N_11723);
nor U13694 (N_13694,N_11991,N_10913);
nand U13695 (N_13695,N_10431,N_11785);
or U13696 (N_13696,N_11062,N_11273);
nor U13697 (N_13697,N_11628,N_11954);
nand U13698 (N_13698,N_10492,N_11628);
or U13699 (N_13699,N_10905,N_10480);
nor U13700 (N_13700,N_11083,N_11689);
and U13701 (N_13701,N_11991,N_10559);
nand U13702 (N_13702,N_10530,N_10472);
nand U13703 (N_13703,N_11635,N_10325);
nor U13704 (N_13704,N_11139,N_11913);
nand U13705 (N_13705,N_10523,N_10166);
nand U13706 (N_13706,N_10056,N_10050);
nor U13707 (N_13707,N_10868,N_11082);
or U13708 (N_13708,N_10685,N_10607);
and U13709 (N_13709,N_11234,N_11587);
or U13710 (N_13710,N_10626,N_11404);
or U13711 (N_13711,N_10788,N_11497);
nor U13712 (N_13712,N_11011,N_11401);
and U13713 (N_13713,N_11528,N_10325);
xnor U13714 (N_13714,N_10743,N_11593);
and U13715 (N_13715,N_10932,N_10432);
or U13716 (N_13716,N_11527,N_10658);
nand U13717 (N_13717,N_11626,N_11423);
and U13718 (N_13718,N_11348,N_10979);
and U13719 (N_13719,N_11975,N_11178);
nor U13720 (N_13720,N_10818,N_10557);
nor U13721 (N_13721,N_10750,N_11186);
or U13722 (N_13722,N_10856,N_10791);
or U13723 (N_13723,N_10795,N_11627);
or U13724 (N_13724,N_10192,N_10777);
nor U13725 (N_13725,N_11926,N_11774);
nor U13726 (N_13726,N_10108,N_11849);
nor U13727 (N_13727,N_11965,N_10265);
and U13728 (N_13728,N_10677,N_10205);
and U13729 (N_13729,N_10158,N_10027);
and U13730 (N_13730,N_10302,N_10261);
or U13731 (N_13731,N_11645,N_10666);
and U13732 (N_13732,N_11167,N_11141);
nand U13733 (N_13733,N_10498,N_11971);
and U13734 (N_13734,N_10495,N_10971);
nor U13735 (N_13735,N_10517,N_11535);
or U13736 (N_13736,N_11154,N_10858);
nand U13737 (N_13737,N_11957,N_10643);
nand U13738 (N_13738,N_11900,N_10377);
or U13739 (N_13739,N_11657,N_11065);
and U13740 (N_13740,N_10218,N_11298);
and U13741 (N_13741,N_10991,N_11931);
nor U13742 (N_13742,N_10364,N_11090);
nor U13743 (N_13743,N_11408,N_10296);
and U13744 (N_13744,N_11216,N_10991);
or U13745 (N_13745,N_11720,N_11257);
nand U13746 (N_13746,N_10582,N_10928);
and U13747 (N_13747,N_10973,N_10572);
nand U13748 (N_13748,N_11630,N_10710);
or U13749 (N_13749,N_10414,N_11372);
or U13750 (N_13750,N_10037,N_10008);
nand U13751 (N_13751,N_10599,N_11667);
or U13752 (N_13752,N_11623,N_11734);
nand U13753 (N_13753,N_10574,N_10921);
and U13754 (N_13754,N_11020,N_10917);
nor U13755 (N_13755,N_11860,N_11162);
or U13756 (N_13756,N_11167,N_11531);
nor U13757 (N_13757,N_10960,N_11002);
nand U13758 (N_13758,N_10164,N_10496);
and U13759 (N_13759,N_11387,N_11414);
or U13760 (N_13760,N_10108,N_10438);
nor U13761 (N_13761,N_11383,N_10220);
or U13762 (N_13762,N_11205,N_11843);
or U13763 (N_13763,N_10677,N_10334);
nor U13764 (N_13764,N_11947,N_11333);
and U13765 (N_13765,N_10311,N_11614);
and U13766 (N_13766,N_11045,N_10075);
nor U13767 (N_13767,N_11539,N_11943);
or U13768 (N_13768,N_11542,N_11301);
nand U13769 (N_13769,N_10415,N_10045);
and U13770 (N_13770,N_10435,N_10325);
and U13771 (N_13771,N_11091,N_10648);
or U13772 (N_13772,N_11235,N_11911);
nor U13773 (N_13773,N_11522,N_11621);
nand U13774 (N_13774,N_11627,N_11643);
or U13775 (N_13775,N_10432,N_10956);
or U13776 (N_13776,N_11540,N_10642);
or U13777 (N_13777,N_11765,N_10762);
nand U13778 (N_13778,N_11435,N_10793);
or U13779 (N_13779,N_10207,N_10136);
or U13780 (N_13780,N_10449,N_11159);
nand U13781 (N_13781,N_11642,N_11873);
nand U13782 (N_13782,N_11128,N_10585);
and U13783 (N_13783,N_11204,N_11078);
and U13784 (N_13784,N_10748,N_10133);
nor U13785 (N_13785,N_11383,N_10771);
nor U13786 (N_13786,N_10986,N_11301);
and U13787 (N_13787,N_10253,N_10900);
nand U13788 (N_13788,N_10058,N_11801);
or U13789 (N_13789,N_11918,N_11796);
nand U13790 (N_13790,N_11589,N_11703);
or U13791 (N_13791,N_10574,N_10694);
nand U13792 (N_13792,N_11655,N_10549);
nor U13793 (N_13793,N_11299,N_10137);
or U13794 (N_13794,N_11280,N_10011);
nand U13795 (N_13795,N_11579,N_11903);
nand U13796 (N_13796,N_10858,N_11455);
or U13797 (N_13797,N_10757,N_11051);
or U13798 (N_13798,N_10381,N_11267);
and U13799 (N_13799,N_10664,N_11363);
nand U13800 (N_13800,N_11836,N_11393);
nand U13801 (N_13801,N_11552,N_10536);
or U13802 (N_13802,N_11752,N_11623);
or U13803 (N_13803,N_11969,N_10143);
or U13804 (N_13804,N_10787,N_10302);
nor U13805 (N_13805,N_10785,N_10908);
or U13806 (N_13806,N_11256,N_10451);
nand U13807 (N_13807,N_10677,N_11601);
nor U13808 (N_13808,N_11298,N_11384);
nand U13809 (N_13809,N_11625,N_10133);
and U13810 (N_13810,N_10646,N_10752);
and U13811 (N_13811,N_10750,N_11808);
or U13812 (N_13812,N_11496,N_10312);
and U13813 (N_13813,N_10038,N_10729);
nand U13814 (N_13814,N_10055,N_11215);
nor U13815 (N_13815,N_10434,N_11080);
nor U13816 (N_13816,N_10647,N_10884);
or U13817 (N_13817,N_11231,N_10579);
and U13818 (N_13818,N_11707,N_10483);
or U13819 (N_13819,N_10190,N_11440);
and U13820 (N_13820,N_10586,N_11739);
and U13821 (N_13821,N_11249,N_10311);
or U13822 (N_13822,N_11577,N_10926);
or U13823 (N_13823,N_11775,N_11741);
nor U13824 (N_13824,N_10890,N_11876);
and U13825 (N_13825,N_10191,N_11587);
and U13826 (N_13826,N_10513,N_10312);
nand U13827 (N_13827,N_11643,N_10671);
or U13828 (N_13828,N_11322,N_10970);
and U13829 (N_13829,N_11226,N_11351);
nand U13830 (N_13830,N_10906,N_11722);
or U13831 (N_13831,N_11631,N_11305);
nand U13832 (N_13832,N_10526,N_10083);
nand U13833 (N_13833,N_11471,N_11728);
or U13834 (N_13834,N_10027,N_11551);
or U13835 (N_13835,N_11210,N_10393);
or U13836 (N_13836,N_10717,N_11008);
nand U13837 (N_13837,N_11780,N_11987);
or U13838 (N_13838,N_11528,N_10069);
or U13839 (N_13839,N_10117,N_11468);
nand U13840 (N_13840,N_10962,N_11764);
or U13841 (N_13841,N_10545,N_10606);
and U13842 (N_13842,N_10972,N_10943);
nand U13843 (N_13843,N_11274,N_10879);
nor U13844 (N_13844,N_10718,N_11431);
nor U13845 (N_13845,N_11172,N_10916);
and U13846 (N_13846,N_10211,N_10225);
and U13847 (N_13847,N_11210,N_10633);
nand U13848 (N_13848,N_11499,N_10018);
and U13849 (N_13849,N_11916,N_10205);
nand U13850 (N_13850,N_11482,N_11689);
or U13851 (N_13851,N_10213,N_10602);
and U13852 (N_13852,N_10852,N_11912);
nor U13853 (N_13853,N_10134,N_10498);
nand U13854 (N_13854,N_11855,N_10414);
and U13855 (N_13855,N_10041,N_10845);
or U13856 (N_13856,N_11842,N_11269);
nand U13857 (N_13857,N_11297,N_11579);
and U13858 (N_13858,N_11724,N_10507);
nand U13859 (N_13859,N_11854,N_10970);
nor U13860 (N_13860,N_10272,N_10535);
nor U13861 (N_13861,N_11402,N_10803);
and U13862 (N_13862,N_11672,N_10022);
nand U13863 (N_13863,N_11562,N_10789);
and U13864 (N_13864,N_11381,N_11157);
and U13865 (N_13865,N_11955,N_11348);
and U13866 (N_13866,N_10830,N_10454);
nor U13867 (N_13867,N_11838,N_10692);
or U13868 (N_13868,N_10372,N_10256);
nand U13869 (N_13869,N_10303,N_11148);
or U13870 (N_13870,N_10239,N_10323);
nand U13871 (N_13871,N_10593,N_11248);
and U13872 (N_13872,N_10396,N_11657);
or U13873 (N_13873,N_10716,N_11442);
or U13874 (N_13874,N_11271,N_11263);
or U13875 (N_13875,N_11765,N_10883);
and U13876 (N_13876,N_10765,N_10925);
nand U13877 (N_13877,N_10767,N_10828);
nor U13878 (N_13878,N_10765,N_11385);
nand U13879 (N_13879,N_10613,N_10061);
nor U13880 (N_13880,N_10480,N_10039);
and U13881 (N_13881,N_10074,N_11688);
nor U13882 (N_13882,N_10838,N_11196);
nand U13883 (N_13883,N_10758,N_11722);
or U13884 (N_13884,N_11248,N_10102);
and U13885 (N_13885,N_10416,N_11901);
and U13886 (N_13886,N_11773,N_11833);
nand U13887 (N_13887,N_11830,N_11949);
nor U13888 (N_13888,N_10992,N_11547);
nand U13889 (N_13889,N_10784,N_11890);
and U13890 (N_13890,N_10107,N_10855);
nand U13891 (N_13891,N_11209,N_11206);
nand U13892 (N_13892,N_10177,N_11655);
and U13893 (N_13893,N_11665,N_10646);
nand U13894 (N_13894,N_11289,N_11972);
and U13895 (N_13895,N_10498,N_11448);
or U13896 (N_13896,N_10402,N_10701);
nand U13897 (N_13897,N_10697,N_10746);
nor U13898 (N_13898,N_11284,N_11828);
nor U13899 (N_13899,N_11610,N_10762);
or U13900 (N_13900,N_11117,N_11358);
nor U13901 (N_13901,N_11304,N_10355);
nand U13902 (N_13902,N_11924,N_10225);
nand U13903 (N_13903,N_11706,N_11114);
nor U13904 (N_13904,N_11764,N_10157);
or U13905 (N_13905,N_10191,N_11858);
or U13906 (N_13906,N_11231,N_11969);
nand U13907 (N_13907,N_10667,N_11102);
xor U13908 (N_13908,N_10903,N_11857);
and U13909 (N_13909,N_11276,N_11134);
nand U13910 (N_13910,N_11461,N_11675);
nor U13911 (N_13911,N_10654,N_11427);
nand U13912 (N_13912,N_10222,N_11847);
nand U13913 (N_13913,N_11103,N_10266);
and U13914 (N_13914,N_10751,N_10108);
or U13915 (N_13915,N_11376,N_10702);
nor U13916 (N_13916,N_10979,N_10121);
and U13917 (N_13917,N_10295,N_11183);
or U13918 (N_13918,N_10759,N_10546);
or U13919 (N_13919,N_11338,N_10910);
and U13920 (N_13920,N_10635,N_10582);
nand U13921 (N_13921,N_10881,N_10356);
nand U13922 (N_13922,N_11835,N_10629);
nor U13923 (N_13923,N_11443,N_11251);
nor U13924 (N_13924,N_11195,N_10830);
nand U13925 (N_13925,N_11768,N_11042);
and U13926 (N_13926,N_10499,N_11569);
and U13927 (N_13927,N_11559,N_11041);
nand U13928 (N_13928,N_10247,N_11039);
nand U13929 (N_13929,N_11994,N_10302);
nand U13930 (N_13930,N_10151,N_10476);
and U13931 (N_13931,N_10195,N_11321);
nor U13932 (N_13932,N_11002,N_11773);
nand U13933 (N_13933,N_11367,N_10012);
or U13934 (N_13934,N_10569,N_10244);
or U13935 (N_13935,N_11151,N_11200);
and U13936 (N_13936,N_10438,N_10370);
or U13937 (N_13937,N_11970,N_11828);
nor U13938 (N_13938,N_10348,N_10750);
or U13939 (N_13939,N_10776,N_10811);
nor U13940 (N_13940,N_10058,N_10491);
or U13941 (N_13941,N_11981,N_10174);
or U13942 (N_13942,N_10377,N_11155);
nand U13943 (N_13943,N_10862,N_10760);
or U13944 (N_13944,N_10669,N_11095);
nand U13945 (N_13945,N_10112,N_10924);
nand U13946 (N_13946,N_11793,N_10903);
nor U13947 (N_13947,N_10025,N_10572);
and U13948 (N_13948,N_11336,N_10660);
nor U13949 (N_13949,N_11693,N_10941);
nand U13950 (N_13950,N_11737,N_10834);
and U13951 (N_13951,N_10135,N_10400);
or U13952 (N_13952,N_10004,N_11842);
nor U13953 (N_13953,N_11755,N_10531);
nor U13954 (N_13954,N_10845,N_11619);
and U13955 (N_13955,N_11657,N_10027);
or U13956 (N_13956,N_11223,N_10193);
and U13957 (N_13957,N_10980,N_11598);
nor U13958 (N_13958,N_10781,N_10578);
nand U13959 (N_13959,N_11184,N_11147);
nor U13960 (N_13960,N_10018,N_11447);
and U13961 (N_13961,N_11826,N_11557);
and U13962 (N_13962,N_11217,N_11772);
and U13963 (N_13963,N_11842,N_10575);
and U13964 (N_13964,N_10757,N_10658);
nor U13965 (N_13965,N_10121,N_11110);
or U13966 (N_13966,N_10320,N_10739);
or U13967 (N_13967,N_10943,N_10594);
or U13968 (N_13968,N_10006,N_11171);
and U13969 (N_13969,N_11864,N_11680);
and U13970 (N_13970,N_10639,N_10930);
and U13971 (N_13971,N_11968,N_11546);
and U13972 (N_13972,N_10283,N_10895);
nor U13973 (N_13973,N_11675,N_10941);
nor U13974 (N_13974,N_11916,N_11932);
or U13975 (N_13975,N_11294,N_11522);
or U13976 (N_13976,N_11074,N_10286);
nand U13977 (N_13977,N_11124,N_10746);
and U13978 (N_13978,N_11697,N_10702);
or U13979 (N_13979,N_10816,N_11420);
or U13980 (N_13980,N_11048,N_10023);
nor U13981 (N_13981,N_11786,N_10214);
nand U13982 (N_13982,N_11947,N_11398);
and U13983 (N_13983,N_11829,N_10996);
nor U13984 (N_13984,N_10527,N_10157);
or U13985 (N_13985,N_10127,N_11628);
nor U13986 (N_13986,N_11137,N_10664);
or U13987 (N_13987,N_11460,N_10840);
or U13988 (N_13988,N_11548,N_10528);
nand U13989 (N_13989,N_10517,N_11931);
and U13990 (N_13990,N_10168,N_11485);
nor U13991 (N_13991,N_10057,N_10509);
and U13992 (N_13992,N_10245,N_10076);
nor U13993 (N_13993,N_11777,N_10750);
or U13994 (N_13994,N_10921,N_11826);
nor U13995 (N_13995,N_10959,N_11685);
nor U13996 (N_13996,N_11310,N_11286);
or U13997 (N_13997,N_10258,N_10551);
or U13998 (N_13998,N_11859,N_11650);
and U13999 (N_13999,N_11254,N_10722);
nor U14000 (N_14000,N_12294,N_13196);
nand U14001 (N_14001,N_13054,N_13862);
or U14002 (N_14002,N_13357,N_12896);
nor U14003 (N_14003,N_12146,N_13016);
nor U14004 (N_14004,N_12767,N_12353);
and U14005 (N_14005,N_12555,N_13596);
nand U14006 (N_14006,N_12153,N_12817);
nand U14007 (N_14007,N_13132,N_13377);
or U14008 (N_14008,N_12542,N_12168);
and U14009 (N_14009,N_12221,N_12184);
nand U14010 (N_14010,N_12999,N_13190);
nand U14011 (N_14011,N_13847,N_13457);
or U14012 (N_14012,N_13694,N_12070);
nor U14013 (N_14013,N_13979,N_12578);
and U14014 (N_14014,N_13333,N_13871);
and U14015 (N_14015,N_13358,N_13763);
nand U14016 (N_14016,N_13512,N_13602);
and U14017 (N_14017,N_12741,N_12994);
nor U14018 (N_14018,N_13989,N_13469);
nand U14019 (N_14019,N_13254,N_12851);
nor U14020 (N_14020,N_13153,N_12998);
and U14021 (N_14021,N_13137,N_12382);
nor U14022 (N_14022,N_13405,N_13232);
or U14023 (N_14023,N_12076,N_12937);
nor U14024 (N_14024,N_13946,N_13026);
and U14025 (N_14025,N_12085,N_12003);
nand U14026 (N_14026,N_13453,N_12406);
nor U14027 (N_14027,N_13777,N_13362);
and U14028 (N_14028,N_13423,N_12758);
nand U14029 (N_14029,N_13073,N_13613);
or U14030 (N_14030,N_12032,N_13143);
nand U14031 (N_14031,N_13677,N_12704);
nand U14032 (N_14032,N_13755,N_12694);
and U14033 (N_14033,N_13265,N_12540);
nand U14034 (N_14034,N_12558,N_12254);
and U14035 (N_14035,N_13240,N_13919);
nor U14036 (N_14036,N_12652,N_12264);
nand U14037 (N_14037,N_13985,N_12666);
and U14038 (N_14038,N_12709,N_13787);
nand U14039 (N_14039,N_12503,N_12728);
nand U14040 (N_14040,N_13242,N_13491);
nand U14041 (N_14041,N_12585,N_12706);
nand U14042 (N_14042,N_12436,N_13536);
and U14043 (N_14043,N_12904,N_13388);
nand U14044 (N_14044,N_12380,N_13443);
nand U14045 (N_14045,N_12017,N_13526);
or U14046 (N_14046,N_12965,N_13781);
and U14047 (N_14047,N_13560,N_13421);
nor U14048 (N_14048,N_13138,N_12049);
and U14049 (N_14049,N_12266,N_13625);
or U14050 (N_14050,N_12393,N_12403);
and U14051 (N_14051,N_13223,N_12968);
and U14052 (N_14052,N_12040,N_12243);
nand U14053 (N_14053,N_13945,N_12592);
nand U14054 (N_14054,N_12966,N_12396);
or U14055 (N_14055,N_13622,N_13730);
or U14056 (N_14056,N_12148,N_13898);
nor U14057 (N_14057,N_13752,N_12330);
and U14058 (N_14058,N_12807,N_13692);
nor U14059 (N_14059,N_13316,N_13340);
or U14060 (N_14060,N_12082,N_13507);
or U14061 (N_14061,N_13222,N_12499);
or U14062 (N_14062,N_13515,N_12844);
and U14063 (N_14063,N_12385,N_13581);
nand U14064 (N_14064,N_13637,N_12210);
nand U14065 (N_14065,N_13228,N_12496);
and U14066 (N_14066,N_12888,N_13765);
nand U14067 (N_14067,N_12402,N_13575);
or U14068 (N_14068,N_13773,N_13426);
or U14069 (N_14069,N_13470,N_12283);
or U14070 (N_14070,N_12489,N_13970);
nand U14071 (N_14071,N_13539,N_12957);
nor U14072 (N_14072,N_13798,N_13125);
and U14073 (N_14073,N_12880,N_13088);
nand U14074 (N_14074,N_13354,N_13929);
and U14075 (N_14075,N_12260,N_13936);
nand U14076 (N_14076,N_13455,N_13084);
nand U14077 (N_14077,N_13049,N_12103);
or U14078 (N_14078,N_12952,N_12799);
or U14079 (N_14079,N_12322,N_12716);
nor U14080 (N_14080,N_13447,N_13029);
nand U14081 (N_14081,N_13211,N_13135);
nand U14082 (N_14082,N_12375,N_12151);
nand U14083 (N_14083,N_13425,N_13010);
and U14084 (N_14084,N_13188,N_13605);
nand U14085 (N_14085,N_13661,N_12123);
xor U14086 (N_14086,N_12849,N_13077);
or U14087 (N_14087,N_12836,N_13550);
nand U14088 (N_14088,N_13434,N_12480);
nor U14089 (N_14089,N_12869,N_13626);
and U14090 (N_14090,N_13294,N_12864);
and U14091 (N_14091,N_12078,N_12627);
and U14092 (N_14092,N_12596,N_13187);
and U14093 (N_14093,N_13905,N_13683);
nor U14094 (N_14094,N_12793,N_12001);
or U14095 (N_14095,N_12095,N_13900);
nand U14096 (N_14096,N_12356,N_13156);
or U14097 (N_14097,N_12399,N_13206);
nor U14098 (N_14098,N_12868,N_13090);
nor U14099 (N_14099,N_13805,N_12919);
or U14100 (N_14100,N_12613,N_12363);
and U14101 (N_14101,N_13967,N_12346);
and U14102 (N_14102,N_13731,N_13636);
nand U14103 (N_14103,N_12006,N_13503);
or U14104 (N_14104,N_12282,N_13315);
or U14105 (N_14105,N_12622,N_12617);
and U14106 (N_14106,N_12140,N_12909);
or U14107 (N_14107,N_12191,N_13344);
nor U14108 (N_14108,N_13573,N_13348);
nand U14109 (N_14109,N_12347,N_12944);
nor U14110 (N_14110,N_12659,N_13809);
nand U14111 (N_14111,N_13591,N_12201);
nand U14112 (N_14112,N_12673,N_13243);
nor U14113 (N_14113,N_12843,N_12926);
and U14114 (N_14114,N_13392,N_12335);
nor U14115 (N_14115,N_12536,N_12788);
nand U14116 (N_14116,N_13619,N_12316);
nor U14117 (N_14117,N_12386,N_12566);
or U14118 (N_14118,N_12111,N_12114);
nand U14119 (N_14119,N_13947,N_12400);
nor U14120 (N_14120,N_12634,N_12731);
xnor U14121 (N_14121,N_12593,N_12862);
nor U14122 (N_14122,N_13982,N_13704);
nand U14123 (N_14123,N_13725,N_12832);
nor U14124 (N_14124,N_13885,N_13972);
or U14125 (N_14125,N_12630,N_12005);
or U14126 (N_14126,N_13075,N_13247);
nand U14127 (N_14127,N_12182,N_13177);
nand U14128 (N_14128,N_13008,N_13118);
xor U14129 (N_14129,N_13909,N_13456);
nor U14130 (N_14130,N_13363,N_13230);
and U14131 (N_14131,N_13908,N_12068);
or U14132 (N_14132,N_13480,N_12284);
or U14133 (N_14133,N_12211,N_13767);
xnor U14134 (N_14134,N_13514,N_13145);
or U14135 (N_14135,N_13493,N_13364);
or U14136 (N_14136,N_12199,N_12742);
nor U14137 (N_14137,N_13925,N_13290);
xnor U14138 (N_14138,N_13399,N_12572);
and U14139 (N_14139,N_13673,N_13404);
nand U14140 (N_14140,N_12513,N_12218);
nand U14141 (N_14141,N_13018,N_12415);
nor U14142 (N_14142,N_13600,N_12478);
nand U14143 (N_14143,N_12829,N_12521);
and U14144 (N_14144,N_12544,N_13033);
nand U14145 (N_14145,N_13269,N_12167);
nand U14146 (N_14146,N_13727,N_12112);
nor U14147 (N_14147,N_12147,N_13041);
or U14148 (N_14148,N_12786,N_13039);
nand U14149 (N_14149,N_12384,N_13003);
and U14150 (N_14150,N_13617,N_12495);
and U14151 (N_14151,N_13858,N_12635);
or U14152 (N_14152,N_12669,N_12351);
nor U14153 (N_14153,N_12823,N_13886);
and U14154 (N_14154,N_13586,N_12682);
and U14155 (N_14155,N_13565,N_12019);
nor U14156 (N_14156,N_13562,N_13672);
nand U14157 (N_14157,N_12369,N_12686);
nor U14158 (N_14158,N_12993,N_13748);
or U14159 (N_14159,N_13971,N_13343);
nand U14160 (N_14160,N_12603,N_12859);
nand U14161 (N_14161,N_12238,N_13563);
or U14162 (N_14162,N_12214,N_13571);
and U14163 (N_14163,N_13771,N_13115);
and U14164 (N_14164,N_13367,N_12502);
and U14165 (N_14165,N_12787,N_13258);
nor U14166 (N_14166,N_12413,N_12454);
nand U14167 (N_14167,N_13747,N_12708);
nor U14168 (N_14168,N_13653,N_13834);
nor U14169 (N_14169,N_12421,N_13183);
nand U14170 (N_14170,N_13058,N_12860);
and U14171 (N_14171,N_13328,N_12087);
or U14172 (N_14172,N_13802,N_12277);
nor U14173 (N_14173,N_12714,N_12511);
nand U14174 (N_14174,N_12975,N_12154);
nor U14175 (N_14175,N_13484,N_13783);
and U14176 (N_14176,N_12650,N_13352);
and U14177 (N_14177,N_13784,N_12121);
or U14178 (N_14178,N_12929,N_12169);
and U14179 (N_14179,N_13915,N_12552);
xor U14180 (N_14180,N_12162,N_13131);
nand U14181 (N_14181,N_12805,N_12763);
and U14182 (N_14182,N_13511,N_13454);
nand U14183 (N_14183,N_12133,N_12341);
nor U14184 (N_14184,N_12246,N_13022);
nand U14185 (N_14185,N_13304,N_12483);
and U14186 (N_14186,N_12281,N_12762);
nand U14187 (N_14187,N_12698,N_12989);
nor U14188 (N_14188,N_13686,N_12317);
nand U14189 (N_14189,N_13610,N_13656);
and U14190 (N_14190,N_13698,N_12826);
or U14191 (N_14191,N_13418,N_13116);
nand U14192 (N_14192,N_13816,N_12370);
and U14193 (N_14193,N_12876,N_12395);
nor U14194 (N_14194,N_13827,N_13890);
or U14195 (N_14195,N_12209,N_12835);
or U14196 (N_14196,N_12345,N_13204);
nand U14197 (N_14197,N_12453,N_13452);
nand U14198 (N_14198,N_12446,N_13225);
nor U14199 (N_14199,N_13843,N_13920);
or U14200 (N_14200,N_13293,N_13554);
nand U14201 (N_14201,N_13824,N_13059);
nand U14202 (N_14202,N_12770,N_12924);
nand U14203 (N_14203,N_12379,N_13272);
nand U14204 (N_14204,N_13180,N_12273);
and U14205 (N_14205,N_13370,N_13440);
nor U14206 (N_14206,N_12389,N_12561);
nand U14207 (N_14207,N_12173,N_13549);
nor U14208 (N_14208,N_12515,N_13096);
nand U14209 (N_14209,N_12105,N_12307);
and U14210 (N_14210,N_13048,N_12098);
and U14211 (N_14211,N_12978,N_12658);
nand U14212 (N_14212,N_13815,N_12715);
nand U14213 (N_14213,N_12806,N_13313);
and U14214 (N_14214,N_13275,N_13848);
and U14215 (N_14215,N_12776,N_12271);
or U14216 (N_14216,N_13774,N_12769);
or U14217 (N_14217,N_13064,N_12094);
nor U14218 (N_14218,N_12204,N_12853);
and U14219 (N_14219,N_13921,N_13838);
or U14220 (N_14220,N_12619,N_12481);
nand U14221 (N_14221,N_12426,N_13935);
nor U14222 (N_14222,N_13066,N_12107);
nor U14223 (N_14223,N_13445,N_12202);
nand U14224 (N_14224,N_12913,N_12189);
and U14225 (N_14225,N_12150,N_12229);
nand U14226 (N_14226,N_12309,N_13845);
or U14227 (N_14227,N_12756,N_13589);
nor U14228 (N_14228,N_12482,N_13050);
or U14229 (N_14229,N_13220,N_12620);
nor U14230 (N_14230,N_12933,N_12663);
nand U14231 (N_14231,N_12618,N_13708);
nand U14232 (N_14232,N_12839,N_13969);
or U14233 (N_14233,N_13530,N_12774);
xor U14234 (N_14234,N_12736,N_12041);
and U14235 (N_14235,N_12348,N_13331);
nand U14236 (N_14236,N_13629,N_13253);
or U14237 (N_14237,N_13829,N_12404);
nand U14238 (N_14238,N_12137,N_12522);
or U14239 (N_14239,N_12996,N_12611);
xor U14240 (N_14240,N_13942,N_13281);
or U14241 (N_14241,N_12644,N_13014);
nor U14242 (N_14242,N_13006,N_12304);
and U14243 (N_14243,N_12104,N_12872);
nand U14244 (N_14244,N_12308,N_12754);
nand U14245 (N_14245,N_12329,N_12764);
and U14246 (N_14246,N_13410,N_13311);
nor U14247 (N_14247,N_12713,N_13988);
or U14248 (N_14248,N_13182,N_12240);
and U14249 (N_14249,N_12035,N_13594);
nand U14250 (N_14250,N_12349,N_12936);
nor U14251 (N_14251,N_12466,N_12675);
nand U14252 (N_14252,N_12056,N_12960);
and U14253 (N_14253,N_12165,N_13561);
or U14254 (N_14254,N_12546,N_13711);
nand U14255 (N_14255,N_13390,N_13795);
nand U14256 (N_14256,N_12615,N_13743);
nand U14257 (N_14257,N_12156,N_13938);
nor U14258 (N_14258,N_12647,N_13701);
and U14259 (N_14259,N_13011,N_13648);
nor U14260 (N_14260,N_13044,N_12641);
nor U14261 (N_14261,N_13104,N_12877);
and U14262 (N_14262,N_12719,N_13406);
and U14263 (N_14263,N_12073,N_13466);
nand U14264 (N_14264,N_12100,N_13351);
or U14265 (N_14265,N_12895,N_13065);
nand U14266 (N_14266,N_12905,N_12463);
or U14267 (N_14267,N_12693,N_13785);
nand U14268 (N_14268,N_13583,N_12985);
nor U14269 (N_14269,N_13608,N_13811);
nand U14270 (N_14270,N_12607,N_12205);
and U14271 (N_14271,N_12430,N_12038);
nand U14272 (N_14272,N_12576,N_13793);
and U14273 (N_14273,N_13288,N_13537);
nor U14274 (N_14274,N_13844,N_12725);
nor U14275 (N_14275,N_12458,N_12161);
and U14276 (N_14276,N_12573,N_12560);
and U14277 (N_14277,N_12488,N_13611);
nor U14278 (N_14278,N_12871,N_12126);
nand U14279 (N_14279,N_13121,N_12373);
xnor U14280 (N_14280,N_12724,N_12122);
nand U14281 (N_14281,N_13195,N_13218);
and U14282 (N_14282,N_13531,N_12310);
nand U14283 (N_14283,N_13667,N_13036);
nand U14284 (N_14284,N_13689,N_13252);
or U14285 (N_14285,N_13569,N_13857);
or U14286 (N_14286,N_13172,N_13807);
and U14287 (N_14287,N_13740,N_13607);
nor U14288 (N_14288,N_13310,N_13117);
and U14289 (N_14289,N_13152,N_13389);
or U14290 (N_14290,N_12881,N_13212);
nand U14291 (N_14291,N_13564,N_13579);
nor U14292 (N_14292,N_13662,N_12323);
nor U14293 (N_14293,N_12866,N_12350);
nor U14294 (N_14294,N_12911,N_12293);
nand U14295 (N_14295,N_12730,N_12722);
and U14296 (N_14296,N_12569,N_12670);
nand U14297 (N_14297,N_12688,N_13797);
or U14298 (N_14298,N_13161,N_13061);
nand U14299 (N_14299,N_12071,N_13770);
nand U14300 (N_14300,N_13820,N_12231);
nand U14301 (N_14301,N_12811,N_12442);
nand U14302 (N_14302,N_13160,N_12397);
nor U14303 (N_14303,N_13882,N_12366);
and U14304 (N_14304,N_13801,N_13374);
or U14305 (N_14305,N_12311,N_13422);
nand U14306 (N_14306,N_12196,N_13162);
and U14307 (N_14307,N_13158,N_12270);
nor U14308 (N_14308,N_13499,N_13407);
or U14309 (N_14309,N_13490,N_12128);
or U14310 (N_14310,N_12075,N_12759);
and U14311 (N_14311,N_13063,N_13235);
nor U14312 (N_14312,N_13168,N_12172);
nor U14313 (N_14313,N_13734,N_12320);
or U14314 (N_14314,N_12452,N_12012);
or U14315 (N_14315,N_13199,N_13669);
or U14316 (N_14316,N_13017,N_13699);
and U14317 (N_14317,N_13387,N_12459);
nand U14318 (N_14318,N_13910,N_13893);
and U14319 (N_14319,N_12465,N_13430);
nor U14320 (N_14320,N_13438,N_13080);
and U14321 (N_14321,N_13663,N_13419);
and U14322 (N_14322,N_12574,N_12990);
nor U14323 (N_14323,N_12955,N_13754);
or U14324 (N_14324,N_12987,N_12791);
nor U14325 (N_14325,N_13892,N_13492);
and U14326 (N_14326,N_13442,N_12239);
and U14327 (N_14327,N_13208,N_13529);
nor U14328 (N_14328,N_12761,N_12633);
nand U14329 (N_14329,N_13504,N_12707);
nor U14330 (N_14330,N_13751,N_13170);
and U14331 (N_14331,N_13100,N_13489);
or U14332 (N_14332,N_13585,N_12781);
nand U14333 (N_14333,N_13994,N_13749);
nand U14334 (N_14334,N_12941,N_13639);
nor U14335 (N_14335,N_12557,N_12800);
nand U14336 (N_14336,N_12250,N_13301);
or U14337 (N_14337,N_13334,N_13186);
and U14338 (N_14338,N_12149,N_13286);
nor U14339 (N_14339,N_13513,N_13993);
or U14340 (N_14340,N_12738,N_13013);
and U14341 (N_14341,N_12614,N_12241);
nor U14342 (N_14342,N_12882,N_12512);
and U14343 (N_14343,N_12015,N_13157);
or U14344 (N_14344,N_12841,N_13913);
nor U14345 (N_14345,N_13391,N_13723);
nor U14346 (N_14346,N_13558,N_12610);
nand U14347 (N_14347,N_12291,N_12778);
nor U14348 (N_14348,N_13174,N_13974);
or U14349 (N_14349,N_12449,N_12890);
or U14350 (N_14350,N_13148,N_12117);
or U14351 (N_14351,N_13069,N_12796);
and U14352 (N_14352,N_13034,N_13070);
or U14353 (N_14353,N_12185,N_12176);
and U14354 (N_14354,N_13082,N_12568);
nor U14355 (N_14355,N_13592,N_12498);
nand U14356 (N_14356,N_12684,N_12437);
and U14357 (N_14357,N_13498,N_13192);
nand U14358 (N_14358,N_13666,N_12803);
nand U14359 (N_14359,N_12470,N_13085);
or U14360 (N_14360,N_12609,N_12821);
nor U14361 (N_14361,N_13401,N_13139);
and U14362 (N_14362,N_13287,N_12702);
or U14363 (N_14363,N_12755,N_12562);
nand U14364 (N_14364,N_12979,N_12197);
or U14365 (N_14365,N_13707,N_12834);
nand U14366 (N_14366,N_13710,N_12157);
and U14367 (N_14367,N_13191,N_13649);
and U14368 (N_14368,N_13541,N_12276);
nand U14369 (N_14369,N_13769,N_12414);
and U14370 (N_14370,N_12314,N_12054);
and U14371 (N_14371,N_13122,N_13780);
and U14372 (N_14372,N_13046,N_13806);
nor U14373 (N_14373,N_12678,N_13215);
and U14374 (N_14374,N_13911,N_13580);
nand U14375 (N_14375,N_12712,N_12080);
and U14376 (N_14376,N_12431,N_13828);
nor U14377 (N_14377,N_12267,N_13072);
and U14378 (N_14378,N_13519,N_13523);
nor U14379 (N_14379,N_12847,N_13912);
nand U14380 (N_14380,N_13567,N_13154);
nand U14381 (N_14381,N_13574,N_13759);
and U14382 (N_14382,N_12377,N_13133);
and U14383 (N_14383,N_12765,N_13163);
nor U14384 (N_14384,N_13194,N_12043);
or U14385 (N_14385,N_13381,N_13103);
nand U14386 (N_14386,N_13300,N_12226);
nor U14387 (N_14387,N_12563,N_13201);
nand U14388 (N_14388,N_13329,N_12280);
nand U14389 (N_14389,N_13899,N_12018);
nor U14390 (N_14390,N_12188,N_12654);
or U14391 (N_14391,N_13478,N_12170);
and U14392 (N_14392,N_13856,N_12579);
nand U14393 (N_14393,N_12766,N_13548);
nor U14394 (N_14394,N_13079,N_13339);
nand U14395 (N_14395,N_12494,N_13271);
and U14396 (N_14396,N_13895,N_13146);
or U14397 (N_14397,N_12656,N_13872);
and U14398 (N_14398,N_12288,N_13958);
nor U14399 (N_14399,N_13198,N_13217);
nand U14400 (N_14400,N_12000,N_13149);
nand U14401 (N_14401,N_13397,N_13479);
and U14402 (N_14402,N_13880,N_12268);
nand U14403 (N_14403,N_12381,N_12261);
or U14404 (N_14404,N_12639,N_12789);
nor U14405 (N_14405,N_13144,N_12474);
nor U14406 (N_14406,N_12186,N_12444);
nor U14407 (N_14407,N_12934,N_12740);
nand U14408 (N_14408,N_13630,N_13818);
nand U14409 (N_14409,N_13214,N_13250);
or U14410 (N_14410,N_13705,N_13327);
nor U14411 (N_14411,N_13505,N_13476);
nor U14412 (N_14412,N_12305,N_12674);
and U14413 (N_14413,N_13000,N_13962);
nor U14414 (N_14414,N_12838,N_12491);
and U14415 (N_14415,N_13112,N_13261);
or U14416 (N_14416,N_13094,N_12248);
or U14417 (N_14417,N_13823,N_12321);
nor U14418 (N_14418,N_12178,N_13471);
nand U14419 (N_14419,N_13928,N_12166);
nand U14420 (N_14420,N_12837,N_13709);
nor U14421 (N_14421,N_13995,N_13833);
nand U14422 (N_14422,N_12069,N_12507);
nand U14423 (N_14423,N_13169,N_12528);
or U14424 (N_14424,N_12412,N_13609);
nor U14425 (N_14425,N_12677,N_12245);
nand U14426 (N_14426,N_12024,N_12409);
or U14427 (N_14427,N_13166,N_13732);
nor U14428 (N_14428,N_13446,N_13907);
nor U14429 (N_14429,N_13557,N_12125);
and U14430 (N_14430,N_12700,N_12490);
and U14431 (N_14431,N_12200,N_13245);
or U14432 (N_14432,N_12810,N_12870);
and U14433 (N_14433,N_12134,N_12206);
nor U14434 (N_14434,N_12464,N_12244);
nor U14435 (N_14435,N_12626,N_12976);
nor U14436 (N_14436,N_13477,N_12279);
nor U14437 (N_14437,N_13123,N_13814);
nand U14438 (N_14438,N_13739,N_12954);
and U14439 (N_14439,N_13668,N_12064);
nor U14440 (N_14440,N_13433,N_12886);
nor U14441 (N_14441,N_12629,N_13796);
or U14442 (N_14442,N_12815,N_12879);
or U14443 (N_14443,N_12263,N_12171);
nor U14444 (N_14444,N_12822,N_12598);
nor U14445 (N_14445,N_13257,N_13922);
nor U14446 (N_14446,N_12720,N_12334);
nor U14447 (N_14447,N_13873,N_13291);
or U14448 (N_14448,N_13472,N_13099);
and U14449 (N_14449,N_13142,N_13326);
nand U14450 (N_14450,N_13961,N_12804);
nor U14451 (N_14451,N_13954,N_13980);
or U14452 (N_14452,N_12368,N_12339);
nand U14453 (N_14453,N_12152,N_13950);
and U14454 (N_14454,N_13804,N_12031);
nor U14455 (N_14455,N_13312,N_12110);
nand U14456 (N_14456,N_12432,N_12195);
or U14457 (N_14457,N_12216,N_13598);
nor U14458 (N_14458,N_12548,N_12779);
nand U14459 (N_14459,N_13234,N_13508);
nor U14460 (N_14460,N_12359,N_12131);
and U14461 (N_14461,N_12009,N_12492);
and U14462 (N_14462,N_12388,N_13179);
and U14463 (N_14463,N_12067,N_12451);
or U14464 (N_14464,N_13884,N_12717);
and U14465 (N_14465,N_13572,N_12749);
nand U14466 (N_14466,N_12514,N_13839);
or U14467 (N_14467,N_13266,N_12113);
and U14468 (N_14468,N_13712,N_13128);
and U14469 (N_14469,N_12771,N_13361);
nand U14470 (N_14470,N_13495,N_12477);
or U14471 (N_14471,N_12831,N_13051);
and U14472 (N_14472,N_12225,N_13007);
nand U14473 (N_14473,N_13852,N_12052);
and U14474 (N_14474,N_12021,N_13887);
nor U14475 (N_14475,N_13289,N_13114);
and U14476 (N_14476,N_12753,N_12435);
nor U14477 (N_14477,N_13098,N_13632);
and U14478 (N_14478,N_13321,N_13808);
or U14479 (N_14479,N_12144,N_13292);
and U14480 (N_14480,N_12797,N_13259);
or U14481 (N_14481,N_13497,N_13917);
and U14482 (N_14482,N_12252,N_12943);
nor U14483 (N_14483,N_12930,N_13408);
nand U14484 (N_14484,N_13951,N_12473);
nor U14485 (N_14485,N_13067,N_13924);
nand U14486 (N_14486,N_12772,N_12475);
and U14487 (N_14487,N_13060,N_13934);
xnor U14488 (N_14488,N_12668,N_12892);
nand U14489 (N_14489,N_12407,N_12063);
nor U14490 (N_14490,N_12595,N_13015);
nand U14491 (N_14491,N_12692,N_12660);
nand U14492 (N_14492,N_12504,N_12416);
nand U14493 (N_14493,N_12274,N_13959);
nand U14494 (N_14494,N_12798,N_12604);
nand U14495 (N_14495,N_12139,N_13424);
and U14496 (N_14496,N_12262,N_12194);
and U14497 (N_14497,N_12441,N_12600);
or U14498 (N_14498,N_12648,N_13800);
or U14499 (N_14499,N_13108,N_12234);
and U14500 (N_14500,N_12516,N_13398);
or U14501 (N_14501,N_12986,N_13027);
nand U14502 (N_14502,N_12801,N_13510);
nand U14503 (N_14503,N_12939,N_12013);
and U14504 (N_14504,N_12995,N_13700);
xor U14505 (N_14505,N_13119,N_13772);
nor U14506 (N_14506,N_13535,N_12591);
nand U14507 (N_14507,N_12961,N_13317);
nand U14508 (N_14508,N_13056,N_12319);
nor U14509 (N_14509,N_13178,N_12088);
nand U14510 (N_14510,N_13322,N_12181);
nand U14511 (N_14511,N_13628,N_12649);
and U14512 (N_14512,N_12072,N_12750);
or U14513 (N_14513,N_13427,N_12391);
nor U14514 (N_14514,N_13750,N_13249);
and U14515 (N_14515,N_12907,N_12703);
and U14516 (N_14516,N_12751,N_12057);
or U14517 (N_14517,N_13926,N_13342);
or U14518 (N_14518,N_13200,N_13227);
and U14519 (N_14519,N_13366,N_12981);
nor U14520 (N_14520,N_12116,N_13324);
nor U14521 (N_14521,N_12155,N_12460);
or U14522 (N_14522,N_12527,N_12735);
and U14523 (N_14523,N_13944,N_13246);
nand U14524 (N_14524,N_13889,N_13385);
or U14525 (N_14525,N_12963,N_12325);
and U14526 (N_14526,N_13428,N_13369);
or U14527 (N_14527,N_12295,N_12093);
or U14528 (N_14528,N_12324,N_12020);
nor U14529 (N_14529,N_12136,N_13140);
nor U14530 (N_14530,N_12340,N_12780);
or U14531 (N_14531,N_13937,N_12858);
nand U14532 (N_14532,N_12129,N_13603);
or U14533 (N_14533,N_13518,N_13356);
or U14534 (N_14534,N_12352,N_13376);
nand U14535 (N_14535,N_13778,N_12632);
nand U14536 (N_14536,N_12903,N_13465);
nand U14537 (N_14537,N_13411,N_13810);
or U14538 (N_14538,N_13233,N_13053);
nor U14539 (N_14539,N_12079,N_13753);
or U14540 (N_14540,N_13577,N_13713);
or U14541 (N_14541,N_12265,N_13282);
nand U14542 (N_14542,N_12917,N_12865);
nor U14543 (N_14543,N_12973,N_13687);
or U14544 (N_14544,N_13830,N_12120);
nand U14545 (N_14545,N_12982,N_12300);
nand U14546 (N_14546,N_12951,N_12729);
and U14547 (N_14547,N_13981,N_12795);
nor U14548 (N_14548,N_13955,N_12493);
nand U14549 (N_14549,N_12914,N_12338);
nor U14550 (N_14550,N_13097,N_13719);
nor U14551 (N_14551,N_13997,N_13551);
and U14552 (N_14552,N_13975,N_13803);
nand U14553 (N_14553,N_13320,N_13207);
nand U14554 (N_14554,N_13714,N_12457);
nor U14555 (N_14555,N_12208,N_12467);
nor U14556 (N_14556,N_13881,N_13538);
and U14557 (N_14557,N_12687,N_13684);
nor U14558 (N_14558,N_12824,N_12143);
nor U14559 (N_14559,N_13646,N_13299);
and U14560 (N_14560,N_12737,N_12177);
or U14561 (N_14561,N_13102,N_13615);
and U14562 (N_14562,N_13396,N_12028);
nand U14563 (N_14563,N_13570,N_13870);
or U14564 (N_14564,N_13832,N_12680);
nand U14565 (N_14565,N_13500,N_13078);
nand U14566 (N_14566,N_13120,N_13081);
nor U14567 (N_14567,N_12543,N_13991);
and U14568 (N_14568,N_12550,N_12861);
nand U14569 (N_14569,N_13597,N_12551);
or U14570 (N_14570,N_12401,N_12394);
nand U14571 (N_14571,N_12327,N_12476);
and U14572 (N_14572,N_13879,N_12681);
nor U14573 (N_14573,N_12783,N_12053);
nor U14574 (N_14574,N_13028,N_13262);
and U14575 (N_14575,N_12662,N_13841);
and U14576 (N_14576,N_13378,N_13213);
or U14577 (N_14577,N_12378,N_12940);
nand U14578 (N_14578,N_13875,N_13164);
nand U14579 (N_14579,N_13415,N_12683);
and U14580 (N_14580,N_13024,N_12058);
nand U14581 (N_14581,N_12605,N_13840);
or U14582 (N_14582,N_12902,N_13520);
and U14583 (N_14583,N_12883,N_12946);
nand U14584 (N_14584,N_13429,N_13963);
or U14585 (N_14585,N_12599,N_12570);
xor U14586 (N_14586,N_13635,N_13052);
nand U14587 (N_14587,N_13651,N_13556);
nor U14588 (N_14588,N_12857,N_13604);
xnor U14589 (N_14589,N_13717,N_13525);
and U14590 (N_14590,N_12697,N_12445);
nor U14591 (N_14591,N_12636,N_13973);
nor U14592 (N_14592,N_13221,N_12631);
or U14593 (N_14593,N_13021,N_12927);
nand U14594 (N_14594,N_13949,N_13502);
nor U14595 (N_14595,N_13486,N_13546);
and U14596 (N_14596,N_12343,N_13393);
and U14597 (N_14597,N_13948,N_12333);
and U14598 (N_14598,N_13644,N_13319);
or U14599 (N_14599,N_13267,N_12667);
nor U14600 (N_14600,N_12768,N_12743);
nor U14601 (N_14601,N_13547,N_13268);
or U14602 (N_14602,N_12042,N_12623);
xnor U14603 (N_14603,N_13459,N_13101);
nand U14604 (N_14604,N_12419,N_13332);
or U14605 (N_14605,N_13932,N_13409);
nor U14606 (N_14606,N_13193,N_12091);
and U14607 (N_14607,N_12533,N_13189);
or U14608 (N_14608,N_12898,N_13371);
nor U14609 (N_14609,N_13185,N_12690);
nor U14610 (N_14610,N_12242,N_13030);
or U14611 (N_14611,N_13745,N_12645);
and U14612 (N_14612,N_13057,N_12518);
or U14613 (N_14613,N_13664,N_12701);
and U14614 (N_14614,N_13853,N_13702);
and U14615 (N_14615,N_13501,N_12108);
or U14616 (N_14616,N_12289,N_13431);
or U14617 (N_14617,N_12387,N_13576);
nor U14618 (N_14618,N_12501,N_13256);
nand U14619 (N_14619,N_13458,N_12469);
or U14620 (N_14620,N_13545,N_12956);
nor U14621 (N_14621,N_12935,N_12727);
nor U14622 (N_14622,N_13134,N_12571);
and U14623 (N_14623,N_13314,N_13239);
and U14624 (N_14624,N_13107,N_13931);
xnor U14625 (N_14625,N_12942,N_13297);
or U14626 (N_14626,N_12034,N_12535);
nand U14627 (N_14627,N_12422,N_12567);
nor U14628 (N_14628,N_12893,N_12418);
or U14629 (N_14629,N_12306,N_13766);
and U14630 (N_14630,N_13903,N_13355);
nand U14631 (N_14631,N_13658,N_12734);
or U14632 (N_14632,N_13318,N_13867);
or U14633 (N_14633,N_12062,N_12487);
or U14634 (N_14634,N_13276,N_13055);
or U14635 (N_14635,N_13682,N_13306);
or U14636 (N_14636,N_12411,N_12757);
or U14637 (N_14637,N_12084,N_13209);
nand U14638 (N_14638,N_12183,N_13341);
nand U14639 (N_14639,N_12228,N_12580);
nand U14640 (N_14640,N_13461,N_12900);
nand U14641 (N_14641,N_12594,N_13812);
nand U14642 (N_14642,N_12710,N_12037);
nand U14643 (N_14643,N_13616,N_13606);
nor U14644 (N_14644,N_13280,N_13768);
nand U14645 (N_14645,N_12213,N_12665);
or U14646 (N_14646,N_13516,N_12597);
and U14647 (N_14647,N_13403,N_13086);
nand U14648 (N_14648,N_12785,N_12711);
and U14649 (N_14649,N_12564,N_13894);
or U14650 (N_14650,N_12141,N_12219);
or U14651 (N_14651,N_13638,N_13023);
nor U14652 (N_14652,N_13849,N_12640);
and U14653 (N_14653,N_13861,N_12545);
and U14654 (N_14654,N_12587,N_12971);
nor U14655 (N_14655,N_13851,N_12179);
nand U14656 (N_14656,N_13302,N_12655);
or U14657 (N_14657,N_12287,N_13733);
nor U14658 (N_14658,N_12447,N_13675);
nand U14659 (N_14659,N_13109,N_13353);
and U14660 (N_14660,N_12180,N_13402);
or U14661 (N_14661,N_13744,N_12485);
nand U14662 (N_14662,N_12253,N_12554);
nor U14663 (N_14663,N_13141,N_13706);
nand U14664 (N_14664,N_12486,N_13716);
nor U14665 (N_14665,N_13718,N_13106);
nand U14666 (N_14666,N_12964,N_13680);
or U14667 (N_14667,N_12047,N_13448);
and U14668 (N_14668,N_12390,N_12423);
nor U14669 (N_14669,N_12337,N_13216);
nor U14670 (N_14670,N_12657,N_13968);
nand U14671 (N_14671,N_12651,N_13590);
and U14672 (N_14672,N_12891,N_12559);
or U14673 (N_14673,N_13004,N_12429);
nor U14674 (N_14674,N_12376,N_12606);
and U14675 (N_14675,N_12988,N_12297);
and U14676 (N_14676,N_13864,N_12203);
or U14677 (N_14677,N_13042,N_13775);
nand U14678 (N_14678,N_13741,N_12468);
nor U14679 (N_14679,N_13365,N_12685);
nand U14680 (N_14680,N_13437,N_12664);
nor U14681 (N_14681,N_12777,N_13978);
nor U14682 (N_14682,N_13742,N_13043);
and U14683 (N_14683,N_13544,N_12582);
nor U14684 (N_14684,N_13624,N_13336);
nand U14685 (N_14685,N_12792,N_13093);
nand U14686 (N_14686,N_12362,N_12109);
nor U14687 (N_14687,N_13124,N_13496);
or U14688 (N_14688,N_12696,N_13826);
nand U14689 (N_14689,N_13309,N_13960);
or U14690 (N_14690,N_12251,N_13308);
nor U14691 (N_14691,N_12257,N_12207);
or U14692 (N_14692,N_13860,N_12539);
nand U14693 (N_14693,N_12531,N_13736);
and U14694 (N_14694,N_13799,N_13940);
nand U14695 (N_14695,N_12292,N_12198);
nor U14696 (N_14696,N_12959,N_13618);
xor U14697 (N_14697,N_13219,N_13241);
nor U14698 (N_14698,N_13005,N_13203);
and U14699 (N_14699,N_13031,N_12889);
nor U14700 (N_14700,N_12510,N_12671);
or U14701 (N_14701,N_13918,N_12901);
and U14702 (N_14702,N_13721,N_12643);
and U14703 (N_14703,N_12255,N_12237);
or U14704 (N_14704,N_12193,N_13383);
and U14705 (N_14705,N_12022,N_13210);
nor U14706 (N_14706,N_13386,N_12608);
nand U14707 (N_14707,N_13165,N_12331);
and U14708 (N_14708,N_13593,N_13620);
nand U14709 (N_14709,N_12312,N_12760);
and U14710 (N_14710,N_13776,N_12299);
nand U14711 (N_14711,N_12802,N_13916);
xnor U14712 (N_14712,N_12530,N_13762);
or U14713 (N_14713,N_13835,N_13678);
nand U14714 (N_14714,N_12127,N_12672);
nor U14715 (N_14715,N_12479,N_13002);
nand U14716 (N_14716,N_13642,N_13229);
and U14717 (N_14717,N_12290,N_13037);
and U14718 (N_14718,N_12991,N_12164);
nor U14719 (N_14719,N_13126,N_12081);
nor U14720 (N_14720,N_12653,N_13679);
or U14721 (N_14721,N_12928,N_13020);
nor U14722 (N_14722,N_13822,N_12086);
or U14723 (N_14723,N_12679,N_13035);
and U14724 (N_14724,N_13914,N_12819);
or U14725 (N_14725,N_13380,N_13786);
or U14726 (N_14726,N_13284,N_12354);
or U14727 (N_14727,N_12296,N_12520);
nor U14728 (N_14728,N_13986,N_12855);
nor U14729 (N_14729,N_13083,N_12301);
nor U14730 (N_14730,N_13983,N_12044);
or U14731 (N_14731,N_13521,N_13640);
nor U14732 (N_14732,N_12509,N_12361);
nor U14733 (N_14733,N_12119,N_13791);
nand U14734 (N_14734,N_12718,N_12010);
nand U14735 (N_14735,N_13657,N_12752);
nand U14736 (N_14736,N_13467,N_13517);
nor U14737 (N_14737,N_13868,N_13127);
nand U14738 (N_14738,N_12055,N_12025);
and U14739 (N_14739,N_12918,N_12854);
and U14740 (N_14740,N_13226,N_12433);
and U14741 (N_14741,N_12538,N_13697);
nor U14742 (N_14742,N_12586,N_13836);
nor U14743 (N_14743,N_12059,N_12472);
nand U14744 (N_14744,N_13451,N_13506);
and U14745 (N_14745,N_12285,N_12405);
nand U14746 (N_14746,N_13695,N_13176);
nand U14747 (N_14747,N_13939,N_12118);
nor U14748 (N_14748,N_12318,N_13599);
or U14749 (N_14749,N_12408,N_13990);
nor U14750 (N_14750,N_12833,N_13688);
xor U14751 (N_14751,N_12899,N_13621);
xor U14752 (N_14752,N_12074,N_12820);
nand U14753 (N_14753,N_12046,N_13588);
or U14754 (N_14754,N_12142,N_12256);
and U14755 (N_14755,N_13643,N_12060);
nor U14756 (N_14756,N_12227,N_12581);
and U14757 (N_14757,N_12355,N_12002);
nand U14758 (N_14758,N_12365,N_12050);
nor U14759 (N_14759,N_12008,N_13821);
nor U14760 (N_14760,N_13543,N_12588);
or U14761 (N_14761,N_12602,N_13113);
nand U14762 (N_14762,N_12825,N_13439);
nand U14763 (N_14763,N_13110,N_12417);
and U14764 (N_14764,N_12816,N_13485);
nor U14765 (N_14765,N_12970,N_13416);
nor U14766 (N_14766,N_13349,N_12138);
nor U14767 (N_14767,N_12033,N_13345);
or U14768 (N_14768,N_13129,N_13674);
nor U14769 (N_14769,N_13474,N_13159);
or U14770 (N_14770,N_12947,N_12974);
and U14771 (N_14771,N_12455,N_13236);
nor U14772 (N_14772,N_13463,N_13896);
nor U14773 (N_14773,N_12016,N_13450);
or U14774 (N_14774,N_12878,N_12048);
or U14775 (N_14775,N_12233,N_13488);
nor U14776 (N_14776,N_13237,N_12036);
nand U14777 (N_14777,N_12235,N_13902);
and U14778 (N_14778,N_13338,N_12497);
and U14779 (N_14779,N_12326,N_12222);
nor U14780 (N_14780,N_12175,N_13631);
nand U14781 (N_14781,N_13601,N_13482);
nand U14782 (N_14782,N_13987,N_13325);
nor U14783 (N_14783,N_12584,N_13670);
nor U14784 (N_14784,N_12958,N_13789);
nand U14785 (N_14785,N_13966,N_13414);
and U14786 (N_14786,N_12556,N_12969);
and U14787 (N_14787,N_12163,N_13263);
and U14788 (N_14788,N_13943,N_13952);
nand U14789 (N_14789,N_13693,N_13650);
nand U14790 (N_14790,N_13038,N_13136);
or U14791 (N_14791,N_13155,N_13175);
nand U14792 (N_14792,N_12967,N_13859);
nor U14793 (N_14793,N_12925,N_12328);
and U14794 (N_14794,N_12906,N_12910);
nor U14795 (N_14795,N_12007,N_12534);
and U14796 (N_14796,N_12286,N_12332);
and U14797 (N_14797,N_12932,N_13930);
and U14798 (N_14798,N_13435,N_12874);
nand U14799 (N_14799,N_12827,N_13897);
nor U14800 (N_14800,N_12525,N_12357);
nand U14801 (N_14801,N_13953,N_12410);
and U14802 (N_14802,N_13998,N_12027);
or U14803 (N_14803,N_12950,N_12814);
nor U14804 (N_14804,N_13647,N_12863);
or U14805 (N_14805,N_12590,N_12077);
nor U14806 (N_14806,N_12980,N_13509);
and U14807 (N_14807,N_13025,N_12541);
nand U14808 (N_14808,N_13202,N_13273);
and U14809 (N_14809,N_12726,N_13587);
nand U14810 (N_14810,N_12224,N_12462);
or U14811 (N_14811,N_12775,N_13764);
nand U14812 (N_14812,N_12784,N_13087);
and U14813 (N_14813,N_12962,N_12984);
or U14814 (N_14814,N_13372,N_13473);
or U14815 (N_14815,N_13846,N_13032);
and U14816 (N_14816,N_12850,N_13906);
nand U14817 (N_14817,N_13019,N_12739);
nor U14818 (N_14818,N_13654,N_13307);
nand U14819 (N_14819,N_12014,N_13147);
and U14820 (N_14820,N_12661,N_12532);
and U14821 (N_14821,N_13375,N_13788);
and U14822 (N_14822,N_13197,N_13726);
nand U14823 (N_14823,N_12438,N_13384);
or U14824 (N_14824,N_13522,N_13012);
and U14825 (N_14825,N_12004,N_12099);
or U14826 (N_14826,N_12374,N_13641);
and U14827 (N_14827,N_12732,N_13001);
nand U14828 (N_14828,N_12842,N_12508);
nand U14829 (N_14829,N_13475,N_12721);
and U14830 (N_14830,N_13652,N_13584);
and U14831 (N_14831,N_13111,N_12637);
or U14832 (N_14832,N_13837,N_12097);
nand U14833 (N_14833,N_13559,N_12733);
nand U14834 (N_14834,N_13076,N_12398);
nand U14835 (N_14835,N_13298,N_13779);
nand U14836 (N_14836,N_12689,N_13441);
nand U14837 (N_14837,N_13095,N_12269);
nor U14838 (N_14838,N_13181,N_12921);
or U14839 (N_14839,N_12448,N_12336);
and U14840 (N_14840,N_12537,N_13360);
and U14841 (N_14841,N_13255,N_13432);
or U14842 (N_14842,N_13295,N_12030);
nand U14843 (N_14843,N_12549,N_12873);
xor U14844 (N_14844,N_13542,N_13184);
and U14845 (N_14845,N_13062,N_12628);
and U14846 (N_14846,N_12065,N_13244);
nor U14847 (N_14847,N_13413,N_12130);
or U14848 (N_14848,N_13092,N_12931);
nand U14849 (N_14849,N_12790,N_12439);
nand U14850 (N_14850,N_12115,N_12158);
nor U14851 (N_14851,N_13468,N_12887);
nand U14852 (N_14852,N_12589,N_13045);
nand U14853 (N_14853,N_12096,N_12160);
nand U14854 (N_14854,N_13901,N_13279);
or U14855 (N_14855,N_12315,N_13270);
nor U14856 (N_14856,N_13724,N_13368);
nor U14857 (N_14857,N_13655,N_12948);
nor U14858 (N_14858,N_12691,N_13231);
or U14859 (N_14859,N_13068,N_12367);
or U14860 (N_14860,N_12443,N_13382);
xnor U14861 (N_14861,N_12190,N_12232);
or U14862 (N_14862,N_12212,N_13850);
nor U14863 (N_14863,N_13792,N_13956);
and U14864 (N_14864,N_13464,N_12089);
and U14865 (N_14865,N_12553,N_12621);
nor U14866 (N_14866,N_12360,N_13595);
nand U14867 (N_14867,N_13996,N_13040);
and U14868 (N_14868,N_12577,N_12461);
nand U14869 (N_14869,N_13831,N_13260);
and U14870 (N_14870,N_13337,N_13379);
nand U14871 (N_14871,N_12875,N_12174);
and U14872 (N_14872,N_13869,N_13746);
or U14873 (N_14873,N_12747,N_12051);
or U14874 (N_14874,N_13394,N_13728);
or U14875 (N_14875,N_13854,N_13305);
nand U14876 (N_14876,N_13323,N_13933);
nor U14877 (N_14877,N_12145,N_13436);
or U14878 (N_14878,N_12744,N_13941);
and U14879 (N_14879,N_12526,N_12920);
and U14880 (N_14880,N_13524,N_13790);
nor U14881 (N_14881,N_13634,N_12220);
and U14882 (N_14882,N_12428,N_12583);
nor U14883 (N_14883,N_13487,N_13794);
nor U14884 (N_14884,N_13761,N_13335);
nand U14885 (N_14885,N_12923,N_12192);
and U14886 (N_14886,N_13760,N_12102);
and U14887 (N_14887,N_13238,N_12612);
nor U14888 (N_14888,N_13825,N_12215);
nor U14889 (N_14889,N_12601,N_13460);
nor U14890 (N_14890,N_13412,N_12342);
nand U14891 (N_14891,N_13696,N_12364);
and U14892 (N_14892,N_12748,N_12302);
nor U14893 (N_14893,N_13715,N_12471);
and U14894 (N_14894,N_12997,N_13957);
or U14895 (N_14895,N_12427,N_13553);
nor U14896 (N_14896,N_12484,N_13285);
or U14897 (N_14897,N_13346,N_12813);
nand U14898 (N_14898,N_12023,N_12259);
nor U14899 (N_14899,N_12132,N_13923);
or U14900 (N_14900,N_12809,N_13866);
nor U14901 (N_14901,N_13566,N_12344);
or U14902 (N_14902,N_13483,N_13047);
or U14903 (N_14903,N_12922,N_13855);
nor U14904 (N_14904,N_12026,N_12011);
and U14905 (N_14905,N_12061,N_12506);
nand U14906 (N_14906,N_13665,N_13676);
and U14907 (N_14907,N_13167,N_13527);
and U14908 (N_14908,N_12523,N_12845);
nor U14909 (N_14909,N_13251,N_13874);
nor U14910 (N_14910,N_13296,N_13876);
xor U14911 (N_14911,N_13729,N_12090);
nand U14912 (N_14912,N_12705,N_12852);
nor U14913 (N_14913,N_13278,N_13999);
or U14914 (N_14914,N_12945,N_12949);
nand U14915 (N_14915,N_12456,N_12642);
nand U14916 (N_14916,N_13984,N_13722);
nor U14917 (N_14917,N_13883,N_12045);
or U14918 (N_14918,N_13224,N_12187);
xnor U14919 (N_14919,N_12773,N_12897);
or U14920 (N_14920,N_13813,N_12092);
nor U14921 (N_14921,N_12624,N_12247);
and U14922 (N_14922,N_13737,N_13685);
nor U14923 (N_14923,N_12383,N_12124);
or U14924 (N_14924,N_13359,N_12529);
nand U14925 (N_14925,N_13400,N_13540);
and U14926 (N_14926,N_12782,N_12983);
and U14927 (N_14927,N_12818,N_13150);
nand U14928 (N_14928,N_13274,N_12840);
or U14929 (N_14929,N_13614,N_13533);
nand U14930 (N_14930,N_12848,N_12695);
or U14931 (N_14931,N_12830,N_13555);
and U14932 (N_14932,N_13494,N_13782);
nand U14933 (N_14933,N_12908,N_12230);
nand U14934 (N_14934,N_13659,N_12812);
nor U14935 (N_14935,N_13627,N_13888);
nor U14936 (N_14936,N_12159,N_12392);
or U14937 (N_14937,N_12565,N_13105);
or U14938 (N_14938,N_13568,N_12884);
and U14939 (N_14939,N_12699,N_13089);
nor U14940 (N_14940,N_12616,N_13205);
nor U14941 (N_14941,N_13444,N_13660);
nor U14942 (N_14942,N_12575,N_13532);
or U14943 (N_14943,N_13735,N_12646);
nor U14944 (N_14944,N_13965,N_13417);
nor U14945 (N_14945,N_13481,N_13074);
nand U14946 (N_14946,N_12794,N_12272);
nor U14947 (N_14947,N_12372,N_12424);
or U14948 (N_14948,N_13633,N_12885);
or U14949 (N_14949,N_13691,N_12275);
nand U14950 (N_14950,N_13645,N_13863);
nand U14951 (N_14951,N_12517,N_13703);
and U14952 (N_14952,N_13552,N_13758);
or U14953 (N_14953,N_12298,N_12039);
nand U14954 (N_14954,N_13690,N_12440);
nand U14955 (N_14955,N_12972,N_13303);
nor U14956 (N_14956,N_12894,N_13151);
nand U14957 (N_14957,N_12278,N_13350);
and U14958 (N_14958,N_13130,N_12083);
nor U14959 (N_14959,N_13462,N_13842);
nand U14960 (N_14960,N_12420,N_12358);
or U14961 (N_14961,N_12217,N_13992);
nor U14962 (N_14962,N_12953,N_13091);
and U14963 (N_14963,N_12303,N_12371);
or U14964 (N_14964,N_13449,N_12856);
nor U14965 (N_14965,N_12992,N_12313);
or U14966 (N_14966,N_12258,N_13420);
nor U14967 (N_14967,N_13877,N_13277);
nand U14968 (N_14968,N_13865,N_12450);
xnor U14969 (N_14969,N_12846,N_12519);
and U14970 (N_14970,N_12867,N_13977);
nor U14971 (N_14971,N_12249,N_13612);
nand U14972 (N_14972,N_13671,N_13623);
or U14973 (N_14973,N_13347,N_12029);
and U14974 (N_14974,N_13578,N_12915);
and U14975 (N_14975,N_12746,N_13927);
nor U14976 (N_14976,N_13819,N_13757);
nor U14977 (N_14977,N_13071,N_12828);
nor U14978 (N_14978,N_12977,N_13248);
and U14979 (N_14979,N_13330,N_13173);
and U14980 (N_14980,N_13891,N_12676);
or U14981 (N_14981,N_13534,N_13817);
and U14982 (N_14982,N_12808,N_12638);
and U14983 (N_14983,N_12425,N_12101);
nand U14984 (N_14984,N_12745,N_12500);
or U14985 (N_14985,N_12236,N_13373);
nand U14986 (N_14986,N_12723,N_12434);
or U14987 (N_14987,N_12912,N_13009);
nor U14988 (N_14988,N_13171,N_13528);
nand U14989 (N_14989,N_13681,N_13582);
nand U14990 (N_14990,N_13878,N_13964);
or U14991 (N_14991,N_13264,N_12938);
or U14992 (N_14992,N_12625,N_13904);
nand U14993 (N_14993,N_12066,N_12524);
and U14994 (N_14994,N_12135,N_12106);
or U14995 (N_14995,N_13283,N_12505);
or U14996 (N_14996,N_13720,N_12547);
nor U14997 (N_14997,N_13738,N_12916);
and U14998 (N_14998,N_13756,N_13976);
nor U14999 (N_14999,N_12223,N_13395);
nor U15000 (N_15000,N_12326,N_12718);
or U15001 (N_15001,N_13334,N_13973);
and U15002 (N_15002,N_12992,N_12947);
nand U15003 (N_15003,N_13662,N_12083);
or U15004 (N_15004,N_13946,N_13967);
nand U15005 (N_15005,N_13329,N_12941);
or U15006 (N_15006,N_12110,N_13929);
nor U15007 (N_15007,N_12881,N_12087);
and U15008 (N_15008,N_12521,N_12567);
or U15009 (N_15009,N_13475,N_12172);
nor U15010 (N_15010,N_13125,N_12491);
nor U15011 (N_15011,N_13561,N_13074);
nor U15012 (N_15012,N_13166,N_13683);
nand U15013 (N_15013,N_13105,N_12834);
or U15014 (N_15014,N_13170,N_13763);
or U15015 (N_15015,N_13573,N_12342);
nand U15016 (N_15016,N_13969,N_13819);
nor U15017 (N_15017,N_13890,N_12052);
or U15018 (N_15018,N_12000,N_13590);
or U15019 (N_15019,N_13575,N_13849);
nor U15020 (N_15020,N_12083,N_12827);
or U15021 (N_15021,N_13760,N_12177);
and U15022 (N_15022,N_13868,N_12493);
nand U15023 (N_15023,N_13694,N_12490);
and U15024 (N_15024,N_12540,N_12542);
nand U15025 (N_15025,N_12395,N_12233);
and U15026 (N_15026,N_13717,N_12723);
nor U15027 (N_15027,N_12354,N_13535);
nand U15028 (N_15028,N_13546,N_12074);
nor U15029 (N_15029,N_13193,N_13568);
or U15030 (N_15030,N_13718,N_13199);
nand U15031 (N_15031,N_13117,N_13351);
nor U15032 (N_15032,N_13496,N_13284);
and U15033 (N_15033,N_13004,N_12147);
xnor U15034 (N_15034,N_12326,N_12242);
nand U15035 (N_15035,N_13076,N_13866);
or U15036 (N_15036,N_13393,N_13622);
and U15037 (N_15037,N_12099,N_12783);
or U15038 (N_15038,N_12421,N_12273);
or U15039 (N_15039,N_12165,N_13540);
and U15040 (N_15040,N_13320,N_12686);
nor U15041 (N_15041,N_13930,N_13055);
or U15042 (N_15042,N_13362,N_13722);
nand U15043 (N_15043,N_13445,N_13580);
or U15044 (N_15044,N_13420,N_13999);
or U15045 (N_15045,N_12799,N_12812);
or U15046 (N_15046,N_13732,N_12379);
nand U15047 (N_15047,N_12203,N_13004);
nand U15048 (N_15048,N_13762,N_13846);
or U15049 (N_15049,N_12809,N_12175);
nor U15050 (N_15050,N_12641,N_13894);
nor U15051 (N_15051,N_12931,N_13656);
nor U15052 (N_15052,N_13627,N_13876);
or U15053 (N_15053,N_13530,N_12596);
nor U15054 (N_15054,N_13801,N_12247);
nand U15055 (N_15055,N_12859,N_13267);
and U15056 (N_15056,N_13094,N_12724);
nand U15057 (N_15057,N_12804,N_13241);
nor U15058 (N_15058,N_13052,N_13506);
or U15059 (N_15059,N_12220,N_12287);
nor U15060 (N_15060,N_12407,N_12454);
or U15061 (N_15061,N_13021,N_13734);
or U15062 (N_15062,N_12999,N_13413);
nand U15063 (N_15063,N_13683,N_13570);
and U15064 (N_15064,N_13441,N_13497);
nand U15065 (N_15065,N_13560,N_12772);
nor U15066 (N_15066,N_12634,N_13054);
nand U15067 (N_15067,N_13040,N_12475);
nor U15068 (N_15068,N_12104,N_12757);
or U15069 (N_15069,N_13008,N_13070);
nand U15070 (N_15070,N_13310,N_12468);
nand U15071 (N_15071,N_13508,N_12972);
and U15072 (N_15072,N_12848,N_13155);
or U15073 (N_15073,N_13765,N_12070);
or U15074 (N_15074,N_13119,N_13043);
or U15075 (N_15075,N_12373,N_12948);
or U15076 (N_15076,N_12110,N_12752);
and U15077 (N_15077,N_12375,N_13717);
nand U15078 (N_15078,N_12149,N_12462);
nor U15079 (N_15079,N_12075,N_12054);
nor U15080 (N_15080,N_12083,N_12456);
or U15081 (N_15081,N_12346,N_12270);
nand U15082 (N_15082,N_13362,N_12320);
and U15083 (N_15083,N_13011,N_12169);
and U15084 (N_15084,N_13189,N_12035);
or U15085 (N_15085,N_13958,N_12405);
or U15086 (N_15086,N_13496,N_12045);
and U15087 (N_15087,N_12356,N_12605);
or U15088 (N_15088,N_13310,N_12465);
or U15089 (N_15089,N_13473,N_13811);
or U15090 (N_15090,N_13794,N_12889);
or U15091 (N_15091,N_12980,N_12134);
nand U15092 (N_15092,N_13358,N_12440);
nand U15093 (N_15093,N_13981,N_13082);
nand U15094 (N_15094,N_12940,N_13019);
nand U15095 (N_15095,N_12246,N_12009);
or U15096 (N_15096,N_13508,N_13764);
and U15097 (N_15097,N_12410,N_12635);
nand U15098 (N_15098,N_12498,N_12712);
or U15099 (N_15099,N_13756,N_12534);
and U15100 (N_15100,N_13173,N_13794);
or U15101 (N_15101,N_13778,N_12150);
and U15102 (N_15102,N_12449,N_13023);
and U15103 (N_15103,N_12474,N_13096);
and U15104 (N_15104,N_13362,N_12966);
and U15105 (N_15105,N_12761,N_13561);
and U15106 (N_15106,N_13732,N_12479);
or U15107 (N_15107,N_13412,N_12486);
and U15108 (N_15108,N_13866,N_13125);
nand U15109 (N_15109,N_13371,N_12374);
nor U15110 (N_15110,N_12855,N_13249);
nand U15111 (N_15111,N_12637,N_12501);
or U15112 (N_15112,N_12418,N_12638);
or U15113 (N_15113,N_12725,N_12141);
and U15114 (N_15114,N_13560,N_12631);
and U15115 (N_15115,N_12953,N_12148);
nor U15116 (N_15116,N_12665,N_13767);
and U15117 (N_15117,N_13480,N_12107);
nor U15118 (N_15118,N_13500,N_13856);
and U15119 (N_15119,N_13219,N_12986);
nand U15120 (N_15120,N_13798,N_13560);
or U15121 (N_15121,N_13356,N_13663);
or U15122 (N_15122,N_13364,N_12913);
and U15123 (N_15123,N_12089,N_13466);
nor U15124 (N_15124,N_13698,N_12237);
nand U15125 (N_15125,N_12888,N_12659);
and U15126 (N_15126,N_12994,N_12125);
or U15127 (N_15127,N_12734,N_12113);
nor U15128 (N_15128,N_12492,N_13096);
or U15129 (N_15129,N_12689,N_12354);
nand U15130 (N_15130,N_13440,N_12100);
nand U15131 (N_15131,N_12312,N_13645);
nand U15132 (N_15132,N_13960,N_12475);
nor U15133 (N_15133,N_12538,N_12325);
or U15134 (N_15134,N_12662,N_12801);
nand U15135 (N_15135,N_12817,N_12136);
nor U15136 (N_15136,N_13753,N_13648);
xor U15137 (N_15137,N_13385,N_12215);
nor U15138 (N_15138,N_12896,N_13570);
nor U15139 (N_15139,N_13808,N_12486);
or U15140 (N_15140,N_13896,N_13596);
or U15141 (N_15141,N_12936,N_12230);
nor U15142 (N_15142,N_12113,N_12857);
nor U15143 (N_15143,N_13724,N_12731);
and U15144 (N_15144,N_13915,N_13408);
or U15145 (N_15145,N_13029,N_12664);
and U15146 (N_15146,N_13635,N_12139);
nor U15147 (N_15147,N_13120,N_13859);
nand U15148 (N_15148,N_12258,N_13923);
or U15149 (N_15149,N_12797,N_12206);
and U15150 (N_15150,N_13920,N_12884);
and U15151 (N_15151,N_12297,N_13701);
and U15152 (N_15152,N_13921,N_13407);
and U15153 (N_15153,N_12236,N_12397);
nor U15154 (N_15154,N_13773,N_12427);
and U15155 (N_15155,N_13378,N_13617);
nand U15156 (N_15156,N_12473,N_12881);
nand U15157 (N_15157,N_13926,N_12762);
xnor U15158 (N_15158,N_13498,N_13327);
nand U15159 (N_15159,N_13403,N_13621);
nor U15160 (N_15160,N_12302,N_13416);
or U15161 (N_15161,N_13220,N_12280);
or U15162 (N_15162,N_13248,N_13727);
or U15163 (N_15163,N_13852,N_12010);
nand U15164 (N_15164,N_13017,N_12855);
and U15165 (N_15165,N_13169,N_12851);
nor U15166 (N_15166,N_12238,N_13867);
and U15167 (N_15167,N_12655,N_13525);
nand U15168 (N_15168,N_13211,N_13262);
nand U15169 (N_15169,N_13126,N_12910);
and U15170 (N_15170,N_12850,N_12796);
and U15171 (N_15171,N_13326,N_13152);
and U15172 (N_15172,N_12571,N_13277);
nor U15173 (N_15173,N_12541,N_12334);
nor U15174 (N_15174,N_12565,N_12043);
nand U15175 (N_15175,N_12539,N_12286);
or U15176 (N_15176,N_12295,N_12101);
nand U15177 (N_15177,N_12636,N_12496);
or U15178 (N_15178,N_12983,N_13494);
and U15179 (N_15179,N_13722,N_12177);
and U15180 (N_15180,N_13754,N_13238);
nor U15181 (N_15181,N_12653,N_12954);
nor U15182 (N_15182,N_12226,N_13551);
nor U15183 (N_15183,N_13821,N_12438);
nand U15184 (N_15184,N_13717,N_12226);
nand U15185 (N_15185,N_13842,N_12621);
or U15186 (N_15186,N_13280,N_12171);
or U15187 (N_15187,N_13005,N_12653);
nand U15188 (N_15188,N_12599,N_12309);
and U15189 (N_15189,N_12489,N_13942);
nand U15190 (N_15190,N_12256,N_13822);
and U15191 (N_15191,N_13439,N_12900);
nand U15192 (N_15192,N_12895,N_13870);
and U15193 (N_15193,N_12762,N_13637);
nand U15194 (N_15194,N_12081,N_13055);
or U15195 (N_15195,N_13351,N_12937);
or U15196 (N_15196,N_12014,N_13361);
nor U15197 (N_15197,N_12143,N_13462);
nand U15198 (N_15198,N_13458,N_12668);
and U15199 (N_15199,N_12974,N_13216);
or U15200 (N_15200,N_12064,N_13340);
nor U15201 (N_15201,N_13502,N_12189);
nor U15202 (N_15202,N_13079,N_13524);
nor U15203 (N_15203,N_12049,N_13494);
and U15204 (N_15204,N_13186,N_12301);
or U15205 (N_15205,N_13622,N_13466);
nor U15206 (N_15206,N_13496,N_12007);
and U15207 (N_15207,N_12725,N_13563);
or U15208 (N_15208,N_12455,N_13414);
nand U15209 (N_15209,N_12352,N_12871);
or U15210 (N_15210,N_12971,N_12481);
and U15211 (N_15211,N_12860,N_12088);
and U15212 (N_15212,N_12521,N_13055);
xnor U15213 (N_15213,N_13767,N_12160);
nand U15214 (N_15214,N_13442,N_13897);
nand U15215 (N_15215,N_12031,N_13451);
and U15216 (N_15216,N_13243,N_13516);
nor U15217 (N_15217,N_12972,N_13874);
or U15218 (N_15218,N_13754,N_13939);
nand U15219 (N_15219,N_13020,N_12923);
nor U15220 (N_15220,N_13479,N_12144);
nand U15221 (N_15221,N_12630,N_13553);
nor U15222 (N_15222,N_12310,N_12848);
or U15223 (N_15223,N_12466,N_12207);
and U15224 (N_15224,N_12312,N_13580);
and U15225 (N_15225,N_12484,N_12399);
nand U15226 (N_15226,N_13261,N_13641);
nor U15227 (N_15227,N_12434,N_12487);
nand U15228 (N_15228,N_12600,N_12689);
and U15229 (N_15229,N_12022,N_13497);
and U15230 (N_15230,N_12475,N_12416);
and U15231 (N_15231,N_13791,N_12572);
or U15232 (N_15232,N_13606,N_13936);
and U15233 (N_15233,N_13705,N_13095);
xnor U15234 (N_15234,N_13802,N_12385);
and U15235 (N_15235,N_13574,N_12585);
nand U15236 (N_15236,N_12009,N_13098);
nor U15237 (N_15237,N_12188,N_13252);
or U15238 (N_15238,N_12509,N_12962);
nor U15239 (N_15239,N_13951,N_12146);
or U15240 (N_15240,N_13846,N_13646);
nor U15241 (N_15241,N_12611,N_13236);
or U15242 (N_15242,N_12105,N_13616);
or U15243 (N_15243,N_13149,N_13979);
or U15244 (N_15244,N_12144,N_13857);
nand U15245 (N_15245,N_13359,N_12503);
nor U15246 (N_15246,N_13221,N_13671);
or U15247 (N_15247,N_12183,N_13381);
or U15248 (N_15248,N_12736,N_13756);
nor U15249 (N_15249,N_12137,N_12960);
and U15250 (N_15250,N_12540,N_12140);
and U15251 (N_15251,N_12382,N_13158);
or U15252 (N_15252,N_13667,N_12802);
or U15253 (N_15253,N_12282,N_12122);
and U15254 (N_15254,N_12267,N_12284);
and U15255 (N_15255,N_12811,N_13805);
nor U15256 (N_15256,N_12715,N_12419);
nor U15257 (N_15257,N_12866,N_12266);
nand U15258 (N_15258,N_13300,N_12865);
nand U15259 (N_15259,N_13906,N_13865);
and U15260 (N_15260,N_13228,N_13577);
or U15261 (N_15261,N_12875,N_12500);
and U15262 (N_15262,N_13603,N_13542);
and U15263 (N_15263,N_12690,N_13497);
and U15264 (N_15264,N_12049,N_12193);
and U15265 (N_15265,N_12887,N_12726);
nand U15266 (N_15266,N_13642,N_12326);
and U15267 (N_15267,N_12368,N_13481);
nor U15268 (N_15268,N_12442,N_13163);
nor U15269 (N_15269,N_12915,N_12736);
or U15270 (N_15270,N_12858,N_13518);
or U15271 (N_15271,N_12984,N_12569);
and U15272 (N_15272,N_12607,N_13129);
or U15273 (N_15273,N_13859,N_13552);
nand U15274 (N_15274,N_13636,N_12442);
and U15275 (N_15275,N_13935,N_13815);
or U15276 (N_15276,N_13942,N_12949);
and U15277 (N_15277,N_12968,N_12305);
nor U15278 (N_15278,N_13901,N_13443);
or U15279 (N_15279,N_12274,N_13549);
nor U15280 (N_15280,N_13626,N_12906);
or U15281 (N_15281,N_13321,N_13311);
nand U15282 (N_15282,N_12131,N_13298);
nand U15283 (N_15283,N_12441,N_13826);
or U15284 (N_15284,N_13435,N_12272);
and U15285 (N_15285,N_12761,N_12238);
and U15286 (N_15286,N_13733,N_13224);
and U15287 (N_15287,N_13479,N_13056);
or U15288 (N_15288,N_12592,N_12070);
or U15289 (N_15289,N_13349,N_13142);
or U15290 (N_15290,N_13358,N_12807);
nor U15291 (N_15291,N_13541,N_12359);
or U15292 (N_15292,N_12909,N_13451);
and U15293 (N_15293,N_13726,N_13525);
nand U15294 (N_15294,N_12510,N_13795);
xnor U15295 (N_15295,N_12033,N_13126);
nor U15296 (N_15296,N_13562,N_12147);
or U15297 (N_15297,N_12304,N_13501);
and U15298 (N_15298,N_12904,N_12767);
nand U15299 (N_15299,N_12667,N_13980);
nor U15300 (N_15300,N_13942,N_13065);
nor U15301 (N_15301,N_13118,N_13104);
or U15302 (N_15302,N_13281,N_12255);
and U15303 (N_15303,N_13306,N_13592);
nand U15304 (N_15304,N_12678,N_13194);
and U15305 (N_15305,N_13266,N_12541);
or U15306 (N_15306,N_13797,N_13246);
nand U15307 (N_15307,N_13411,N_12131);
or U15308 (N_15308,N_12905,N_13210);
nand U15309 (N_15309,N_12250,N_12735);
nor U15310 (N_15310,N_12680,N_13900);
or U15311 (N_15311,N_12123,N_13870);
nand U15312 (N_15312,N_13040,N_12252);
and U15313 (N_15313,N_13073,N_13479);
or U15314 (N_15314,N_13865,N_13751);
nand U15315 (N_15315,N_13948,N_12398);
and U15316 (N_15316,N_13096,N_12431);
or U15317 (N_15317,N_12101,N_12895);
nor U15318 (N_15318,N_13551,N_12654);
or U15319 (N_15319,N_13463,N_13722);
nand U15320 (N_15320,N_13748,N_12667);
or U15321 (N_15321,N_13171,N_12636);
nand U15322 (N_15322,N_12813,N_12248);
nand U15323 (N_15323,N_12759,N_12224);
nand U15324 (N_15324,N_13777,N_13881);
xor U15325 (N_15325,N_13639,N_12269);
nor U15326 (N_15326,N_13287,N_12247);
nand U15327 (N_15327,N_12782,N_13078);
and U15328 (N_15328,N_13452,N_13508);
nor U15329 (N_15329,N_12589,N_12651);
nand U15330 (N_15330,N_13134,N_12530);
nor U15331 (N_15331,N_12190,N_12946);
nor U15332 (N_15332,N_13743,N_13422);
nand U15333 (N_15333,N_13827,N_12758);
nor U15334 (N_15334,N_12065,N_12173);
nor U15335 (N_15335,N_12625,N_12066);
nand U15336 (N_15336,N_13145,N_12946);
and U15337 (N_15337,N_13768,N_13627);
and U15338 (N_15338,N_13002,N_12293);
or U15339 (N_15339,N_13384,N_13468);
nor U15340 (N_15340,N_13974,N_12944);
nand U15341 (N_15341,N_13729,N_12499);
or U15342 (N_15342,N_13651,N_13107);
nor U15343 (N_15343,N_12365,N_13974);
or U15344 (N_15344,N_13277,N_12136);
and U15345 (N_15345,N_13901,N_12705);
or U15346 (N_15346,N_13476,N_12577);
or U15347 (N_15347,N_13126,N_13169);
and U15348 (N_15348,N_12604,N_12481);
and U15349 (N_15349,N_13173,N_13916);
nand U15350 (N_15350,N_12489,N_12595);
nand U15351 (N_15351,N_13152,N_13386);
nand U15352 (N_15352,N_13222,N_12662);
nor U15353 (N_15353,N_13435,N_12111);
or U15354 (N_15354,N_13946,N_13615);
nor U15355 (N_15355,N_12924,N_13014);
nor U15356 (N_15356,N_13001,N_12657);
nand U15357 (N_15357,N_13313,N_12836);
or U15358 (N_15358,N_13738,N_13272);
nand U15359 (N_15359,N_13129,N_12117);
nand U15360 (N_15360,N_12718,N_12927);
nor U15361 (N_15361,N_13785,N_13237);
and U15362 (N_15362,N_13472,N_13950);
and U15363 (N_15363,N_12390,N_13079);
nor U15364 (N_15364,N_12701,N_12735);
nand U15365 (N_15365,N_12583,N_13671);
nor U15366 (N_15366,N_12892,N_13863);
and U15367 (N_15367,N_13516,N_13897);
or U15368 (N_15368,N_12926,N_12131);
nand U15369 (N_15369,N_12144,N_13467);
and U15370 (N_15370,N_12934,N_13434);
and U15371 (N_15371,N_12530,N_13168);
or U15372 (N_15372,N_13233,N_12784);
and U15373 (N_15373,N_12257,N_12762);
and U15374 (N_15374,N_12542,N_12959);
nor U15375 (N_15375,N_12639,N_12697);
nand U15376 (N_15376,N_12366,N_13818);
and U15377 (N_15377,N_13773,N_13396);
nor U15378 (N_15378,N_12800,N_12541);
nand U15379 (N_15379,N_13758,N_13284);
nand U15380 (N_15380,N_12877,N_13959);
nor U15381 (N_15381,N_13229,N_12624);
or U15382 (N_15382,N_13902,N_13279);
nor U15383 (N_15383,N_13266,N_12554);
nor U15384 (N_15384,N_13218,N_13479);
nand U15385 (N_15385,N_13623,N_12862);
or U15386 (N_15386,N_13797,N_12870);
nor U15387 (N_15387,N_12657,N_12832);
nor U15388 (N_15388,N_12367,N_13007);
nand U15389 (N_15389,N_12562,N_13087);
nand U15390 (N_15390,N_13181,N_12768);
and U15391 (N_15391,N_12931,N_13914);
and U15392 (N_15392,N_13185,N_12158);
and U15393 (N_15393,N_12741,N_13074);
or U15394 (N_15394,N_12118,N_13297);
nand U15395 (N_15395,N_12282,N_13132);
xnor U15396 (N_15396,N_12119,N_12333);
nand U15397 (N_15397,N_12500,N_12040);
nor U15398 (N_15398,N_12888,N_12690);
nor U15399 (N_15399,N_12582,N_13994);
and U15400 (N_15400,N_12714,N_13735);
or U15401 (N_15401,N_12704,N_13096);
or U15402 (N_15402,N_12316,N_12947);
nand U15403 (N_15403,N_13636,N_12413);
nor U15404 (N_15404,N_13016,N_12924);
nand U15405 (N_15405,N_12705,N_13482);
or U15406 (N_15406,N_13986,N_13594);
nand U15407 (N_15407,N_13920,N_13777);
and U15408 (N_15408,N_12027,N_12177);
nor U15409 (N_15409,N_12053,N_13871);
or U15410 (N_15410,N_12232,N_12510);
or U15411 (N_15411,N_12772,N_13847);
nand U15412 (N_15412,N_12502,N_13036);
nand U15413 (N_15413,N_13238,N_12100);
nor U15414 (N_15414,N_13316,N_12343);
or U15415 (N_15415,N_12194,N_12741);
or U15416 (N_15416,N_13830,N_13618);
nand U15417 (N_15417,N_12939,N_12569);
or U15418 (N_15418,N_13280,N_13926);
or U15419 (N_15419,N_13506,N_13573);
nand U15420 (N_15420,N_12558,N_13011);
nand U15421 (N_15421,N_13341,N_12893);
or U15422 (N_15422,N_13523,N_12856);
xor U15423 (N_15423,N_12872,N_12865);
nor U15424 (N_15424,N_13236,N_12916);
or U15425 (N_15425,N_12560,N_12230);
nor U15426 (N_15426,N_12479,N_12053);
nor U15427 (N_15427,N_12323,N_12611);
xor U15428 (N_15428,N_12152,N_13199);
and U15429 (N_15429,N_12081,N_12979);
and U15430 (N_15430,N_12564,N_12495);
and U15431 (N_15431,N_12755,N_13543);
or U15432 (N_15432,N_12049,N_13962);
nand U15433 (N_15433,N_12759,N_12506);
or U15434 (N_15434,N_13786,N_13195);
or U15435 (N_15435,N_12206,N_12040);
or U15436 (N_15436,N_13467,N_12142);
or U15437 (N_15437,N_13844,N_12351);
nor U15438 (N_15438,N_12963,N_12716);
nor U15439 (N_15439,N_12543,N_12160);
and U15440 (N_15440,N_13635,N_13240);
nand U15441 (N_15441,N_13766,N_13187);
nor U15442 (N_15442,N_13977,N_12702);
nand U15443 (N_15443,N_12549,N_12611);
or U15444 (N_15444,N_13121,N_12330);
and U15445 (N_15445,N_13153,N_13672);
or U15446 (N_15446,N_12989,N_13267);
and U15447 (N_15447,N_13729,N_13644);
nand U15448 (N_15448,N_13968,N_13355);
and U15449 (N_15449,N_12237,N_13890);
or U15450 (N_15450,N_12123,N_12512);
and U15451 (N_15451,N_13717,N_12227);
and U15452 (N_15452,N_13377,N_12347);
nand U15453 (N_15453,N_12625,N_13346);
or U15454 (N_15454,N_13599,N_12755);
nand U15455 (N_15455,N_13628,N_13463);
nor U15456 (N_15456,N_12914,N_13619);
nor U15457 (N_15457,N_12158,N_12723);
nor U15458 (N_15458,N_12264,N_12890);
nor U15459 (N_15459,N_13240,N_12954);
nor U15460 (N_15460,N_13893,N_12575);
and U15461 (N_15461,N_13510,N_12467);
nor U15462 (N_15462,N_12094,N_13254);
nor U15463 (N_15463,N_12417,N_12720);
or U15464 (N_15464,N_13724,N_12558);
and U15465 (N_15465,N_13666,N_13002);
or U15466 (N_15466,N_13513,N_13599);
or U15467 (N_15467,N_12434,N_13358);
nor U15468 (N_15468,N_12640,N_13747);
nand U15469 (N_15469,N_12568,N_13758);
nand U15470 (N_15470,N_12626,N_12217);
and U15471 (N_15471,N_12291,N_13456);
or U15472 (N_15472,N_13660,N_13707);
nor U15473 (N_15473,N_12005,N_13532);
nor U15474 (N_15474,N_12072,N_12295);
or U15475 (N_15475,N_12670,N_12466);
and U15476 (N_15476,N_13015,N_13786);
or U15477 (N_15477,N_12981,N_12128);
nor U15478 (N_15478,N_13434,N_13282);
and U15479 (N_15479,N_13703,N_12270);
or U15480 (N_15480,N_12853,N_13319);
or U15481 (N_15481,N_13126,N_13743);
and U15482 (N_15482,N_13453,N_13910);
or U15483 (N_15483,N_13781,N_12716);
nor U15484 (N_15484,N_13554,N_13098);
and U15485 (N_15485,N_13430,N_13884);
or U15486 (N_15486,N_13754,N_13425);
or U15487 (N_15487,N_12209,N_13966);
nor U15488 (N_15488,N_12503,N_12326);
and U15489 (N_15489,N_12843,N_12320);
nor U15490 (N_15490,N_12826,N_12073);
or U15491 (N_15491,N_12900,N_13654);
nor U15492 (N_15492,N_12244,N_12018);
nand U15493 (N_15493,N_13709,N_12929);
and U15494 (N_15494,N_12810,N_13348);
nor U15495 (N_15495,N_12229,N_12564);
and U15496 (N_15496,N_12334,N_13974);
nor U15497 (N_15497,N_12219,N_13750);
and U15498 (N_15498,N_12776,N_13386);
nor U15499 (N_15499,N_12571,N_13789);
or U15500 (N_15500,N_12210,N_12254);
or U15501 (N_15501,N_12569,N_13542);
nor U15502 (N_15502,N_12302,N_13034);
and U15503 (N_15503,N_13808,N_13504);
or U15504 (N_15504,N_13804,N_13618);
and U15505 (N_15505,N_13134,N_12346);
nor U15506 (N_15506,N_12267,N_12834);
or U15507 (N_15507,N_12693,N_12068);
nand U15508 (N_15508,N_13628,N_12861);
or U15509 (N_15509,N_13098,N_13681);
or U15510 (N_15510,N_12869,N_13967);
or U15511 (N_15511,N_12088,N_12775);
and U15512 (N_15512,N_12235,N_12192);
nor U15513 (N_15513,N_13791,N_13201);
nand U15514 (N_15514,N_12534,N_13470);
and U15515 (N_15515,N_13589,N_13227);
nor U15516 (N_15516,N_12608,N_12258);
or U15517 (N_15517,N_12291,N_13472);
and U15518 (N_15518,N_12219,N_13546);
or U15519 (N_15519,N_13213,N_12261);
nand U15520 (N_15520,N_12502,N_12148);
nor U15521 (N_15521,N_12051,N_12437);
and U15522 (N_15522,N_13073,N_12018);
or U15523 (N_15523,N_13108,N_13912);
and U15524 (N_15524,N_12911,N_12693);
nand U15525 (N_15525,N_12265,N_12773);
nand U15526 (N_15526,N_13680,N_12247);
and U15527 (N_15527,N_12190,N_13201);
or U15528 (N_15528,N_13252,N_13187);
and U15529 (N_15529,N_12413,N_12690);
nand U15530 (N_15530,N_13964,N_12791);
nand U15531 (N_15531,N_12984,N_13278);
and U15532 (N_15532,N_13961,N_12077);
and U15533 (N_15533,N_12371,N_12342);
and U15534 (N_15534,N_12806,N_13913);
nor U15535 (N_15535,N_13830,N_13021);
or U15536 (N_15536,N_12173,N_12465);
and U15537 (N_15537,N_13772,N_12454);
or U15538 (N_15538,N_12876,N_12953);
nand U15539 (N_15539,N_13190,N_13768);
and U15540 (N_15540,N_13208,N_13366);
nor U15541 (N_15541,N_12982,N_12909);
or U15542 (N_15542,N_13347,N_13230);
and U15543 (N_15543,N_13460,N_13798);
and U15544 (N_15544,N_13069,N_12145);
nor U15545 (N_15545,N_13864,N_12179);
and U15546 (N_15546,N_13210,N_13707);
nor U15547 (N_15547,N_13075,N_12631);
nor U15548 (N_15548,N_13358,N_12191);
nand U15549 (N_15549,N_13802,N_13332);
nand U15550 (N_15550,N_13820,N_13266);
nand U15551 (N_15551,N_12961,N_13418);
or U15552 (N_15552,N_12516,N_12267);
nand U15553 (N_15553,N_12988,N_13619);
and U15554 (N_15554,N_12761,N_13598);
and U15555 (N_15555,N_12154,N_12850);
nand U15556 (N_15556,N_12257,N_13031);
nand U15557 (N_15557,N_12024,N_13652);
or U15558 (N_15558,N_12124,N_12549);
and U15559 (N_15559,N_13148,N_13596);
nand U15560 (N_15560,N_12679,N_13979);
nor U15561 (N_15561,N_12153,N_13672);
or U15562 (N_15562,N_13241,N_12911);
or U15563 (N_15563,N_12548,N_13199);
nor U15564 (N_15564,N_13662,N_12246);
and U15565 (N_15565,N_13199,N_12388);
nor U15566 (N_15566,N_13116,N_13023);
or U15567 (N_15567,N_12899,N_13088);
and U15568 (N_15568,N_13103,N_12676);
nor U15569 (N_15569,N_12696,N_13020);
and U15570 (N_15570,N_12825,N_12640);
nand U15571 (N_15571,N_12465,N_12593);
and U15572 (N_15572,N_12401,N_13436);
nand U15573 (N_15573,N_13719,N_12810);
nor U15574 (N_15574,N_12882,N_13934);
and U15575 (N_15575,N_12982,N_13283);
and U15576 (N_15576,N_12009,N_12363);
nand U15577 (N_15577,N_12612,N_12470);
or U15578 (N_15578,N_13495,N_13905);
nor U15579 (N_15579,N_13096,N_13232);
nand U15580 (N_15580,N_12370,N_13293);
or U15581 (N_15581,N_12922,N_13259);
nor U15582 (N_15582,N_12161,N_13775);
nor U15583 (N_15583,N_12563,N_13894);
or U15584 (N_15584,N_13836,N_13065);
nand U15585 (N_15585,N_12649,N_12288);
and U15586 (N_15586,N_13232,N_13744);
and U15587 (N_15587,N_12740,N_13974);
nor U15588 (N_15588,N_13099,N_12576);
and U15589 (N_15589,N_13699,N_13919);
nor U15590 (N_15590,N_13419,N_12771);
nor U15591 (N_15591,N_12587,N_12155);
and U15592 (N_15592,N_12166,N_12967);
or U15593 (N_15593,N_13835,N_13968);
and U15594 (N_15594,N_12437,N_13585);
or U15595 (N_15595,N_13349,N_13414);
nand U15596 (N_15596,N_13823,N_12341);
nand U15597 (N_15597,N_13434,N_13286);
or U15598 (N_15598,N_13196,N_13735);
or U15599 (N_15599,N_13941,N_13855);
and U15600 (N_15600,N_13343,N_13455);
or U15601 (N_15601,N_13712,N_13446);
and U15602 (N_15602,N_13416,N_13832);
and U15603 (N_15603,N_13865,N_12561);
or U15604 (N_15604,N_12995,N_13765);
and U15605 (N_15605,N_13091,N_13250);
nand U15606 (N_15606,N_13009,N_12224);
nor U15607 (N_15607,N_12662,N_13777);
nand U15608 (N_15608,N_12507,N_13739);
or U15609 (N_15609,N_12664,N_13159);
nand U15610 (N_15610,N_13118,N_13905);
nand U15611 (N_15611,N_12968,N_13478);
and U15612 (N_15612,N_12476,N_13703);
nor U15613 (N_15613,N_13668,N_12801);
and U15614 (N_15614,N_13271,N_13005);
and U15615 (N_15615,N_13442,N_12321);
nor U15616 (N_15616,N_12981,N_13817);
nor U15617 (N_15617,N_12924,N_12423);
or U15618 (N_15618,N_13472,N_12498);
or U15619 (N_15619,N_13494,N_13688);
nand U15620 (N_15620,N_13144,N_13716);
and U15621 (N_15621,N_13443,N_13218);
or U15622 (N_15622,N_13373,N_13585);
nand U15623 (N_15623,N_13589,N_13228);
and U15624 (N_15624,N_12622,N_12078);
nor U15625 (N_15625,N_12790,N_13243);
nor U15626 (N_15626,N_13807,N_13642);
nand U15627 (N_15627,N_12113,N_12478);
or U15628 (N_15628,N_13893,N_13025);
nor U15629 (N_15629,N_13894,N_12138);
nand U15630 (N_15630,N_12912,N_13154);
or U15631 (N_15631,N_12051,N_12895);
nor U15632 (N_15632,N_12077,N_12899);
or U15633 (N_15633,N_13092,N_13093);
nor U15634 (N_15634,N_12854,N_12906);
and U15635 (N_15635,N_12093,N_13399);
and U15636 (N_15636,N_12269,N_13330);
nor U15637 (N_15637,N_12455,N_12990);
or U15638 (N_15638,N_13979,N_13015);
and U15639 (N_15639,N_13059,N_12755);
nor U15640 (N_15640,N_13270,N_13480);
or U15641 (N_15641,N_12070,N_12406);
nor U15642 (N_15642,N_13351,N_12151);
and U15643 (N_15643,N_12041,N_12184);
nor U15644 (N_15644,N_12040,N_12865);
nand U15645 (N_15645,N_13906,N_12274);
nand U15646 (N_15646,N_13373,N_12728);
nor U15647 (N_15647,N_12283,N_12005);
or U15648 (N_15648,N_13833,N_12615);
and U15649 (N_15649,N_12936,N_13999);
and U15650 (N_15650,N_12860,N_12913);
nor U15651 (N_15651,N_12739,N_13814);
and U15652 (N_15652,N_12449,N_13254);
and U15653 (N_15653,N_13856,N_12029);
nand U15654 (N_15654,N_13828,N_12466);
nor U15655 (N_15655,N_13119,N_12617);
nor U15656 (N_15656,N_12013,N_13831);
and U15657 (N_15657,N_12325,N_13871);
nor U15658 (N_15658,N_13247,N_13683);
and U15659 (N_15659,N_12601,N_12387);
and U15660 (N_15660,N_12875,N_13640);
nor U15661 (N_15661,N_12687,N_12000);
or U15662 (N_15662,N_13717,N_13104);
or U15663 (N_15663,N_13639,N_13977);
nand U15664 (N_15664,N_12536,N_12540);
and U15665 (N_15665,N_13482,N_13873);
and U15666 (N_15666,N_12084,N_12973);
or U15667 (N_15667,N_13703,N_12025);
nor U15668 (N_15668,N_12105,N_13794);
nor U15669 (N_15669,N_13082,N_12514);
nand U15670 (N_15670,N_12712,N_13545);
and U15671 (N_15671,N_12740,N_12029);
nor U15672 (N_15672,N_13070,N_13240);
nor U15673 (N_15673,N_13518,N_13928);
or U15674 (N_15674,N_12457,N_12739);
and U15675 (N_15675,N_13994,N_13952);
or U15676 (N_15676,N_12654,N_12494);
or U15677 (N_15677,N_12002,N_12964);
nand U15678 (N_15678,N_13160,N_12230);
nand U15679 (N_15679,N_13718,N_12463);
or U15680 (N_15680,N_12423,N_13166);
nor U15681 (N_15681,N_13319,N_13896);
nand U15682 (N_15682,N_12721,N_13010);
nor U15683 (N_15683,N_13068,N_13923);
nand U15684 (N_15684,N_13481,N_12725);
nand U15685 (N_15685,N_13076,N_13670);
nand U15686 (N_15686,N_13173,N_13406);
or U15687 (N_15687,N_13136,N_13702);
xor U15688 (N_15688,N_12228,N_13411);
nor U15689 (N_15689,N_13169,N_12253);
and U15690 (N_15690,N_13282,N_13767);
xnor U15691 (N_15691,N_13022,N_13973);
xor U15692 (N_15692,N_12067,N_13203);
or U15693 (N_15693,N_13496,N_13266);
nand U15694 (N_15694,N_12133,N_12855);
or U15695 (N_15695,N_12246,N_12155);
nand U15696 (N_15696,N_13867,N_12419);
and U15697 (N_15697,N_12471,N_12817);
and U15698 (N_15698,N_12193,N_13590);
nor U15699 (N_15699,N_12503,N_12285);
and U15700 (N_15700,N_13513,N_12350);
nor U15701 (N_15701,N_13635,N_13447);
and U15702 (N_15702,N_12924,N_12975);
nor U15703 (N_15703,N_13860,N_13434);
or U15704 (N_15704,N_12656,N_13459);
and U15705 (N_15705,N_12986,N_12668);
or U15706 (N_15706,N_13007,N_12874);
nand U15707 (N_15707,N_13206,N_12405);
nand U15708 (N_15708,N_13617,N_12209);
and U15709 (N_15709,N_13378,N_12556);
nand U15710 (N_15710,N_13788,N_12452);
or U15711 (N_15711,N_13299,N_13580);
nand U15712 (N_15712,N_13939,N_13251);
nor U15713 (N_15713,N_12592,N_13758);
nand U15714 (N_15714,N_12183,N_12879);
and U15715 (N_15715,N_12677,N_12925);
and U15716 (N_15716,N_12601,N_12708);
or U15717 (N_15717,N_12685,N_12598);
or U15718 (N_15718,N_13861,N_12517);
nor U15719 (N_15719,N_13959,N_12521);
or U15720 (N_15720,N_13740,N_13931);
nand U15721 (N_15721,N_12738,N_13127);
or U15722 (N_15722,N_12145,N_12148);
or U15723 (N_15723,N_13901,N_12603);
nand U15724 (N_15724,N_12252,N_13244);
nand U15725 (N_15725,N_13362,N_12919);
or U15726 (N_15726,N_13994,N_12464);
nor U15727 (N_15727,N_13317,N_12462);
nand U15728 (N_15728,N_12755,N_12862);
nand U15729 (N_15729,N_12684,N_13583);
nand U15730 (N_15730,N_13210,N_13448);
and U15731 (N_15731,N_13567,N_13330);
nor U15732 (N_15732,N_13849,N_13511);
and U15733 (N_15733,N_12079,N_12878);
and U15734 (N_15734,N_12205,N_12912);
nor U15735 (N_15735,N_13910,N_13865);
nor U15736 (N_15736,N_12361,N_12076);
nand U15737 (N_15737,N_12021,N_13902);
and U15738 (N_15738,N_12752,N_12440);
or U15739 (N_15739,N_12532,N_12064);
and U15740 (N_15740,N_12478,N_13031);
nand U15741 (N_15741,N_12389,N_13846);
and U15742 (N_15742,N_13504,N_12711);
nor U15743 (N_15743,N_13632,N_12333);
nor U15744 (N_15744,N_13128,N_13708);
and U15745 (N_15745,N_13157,N_13160);
nor U15746 (N_15746,N_12340,N_13839);
or U15747 (N_15747,N_12332,N_12328);
nor U15748 (N_15748,N_13538,N_12035);
nand U15749 (N_15749,N_12630,N_12671);
nor U15750 (N_15750,N_12681,N_12162);
or U15751 (N_15751,N_13087,N_12334);
nand U15752 (N_15752,N_12495,N_12412);
or U15753 (N_15753,N_13897,N_12837);
nor U15754 (N_15754,N_13270,N_12072);
or U15755 (N_15755,N_12134,N_12023);
and U15756 (N_15756,N_12487,N_12931);
and U15757 (N_15757,N_13987,N_13756);
or U15758 (N_15758,N_12875,N_12968);
nand U15759 (N_15759,N_13820,N_12123);
nor U15760 (N_15760,N_12120,N_12376);
or U15761 (N_15761,N_13999,N_12430);
and U15762 (N_15762,N_13673,N_13924);
nor U15763 (N_15763,N_13370,N_13580);
and U15764 (N_15764,N_13984,N_12384);
and U15765 (N_15765,N_12366,N_12128);
nand U15766 (N_15766,N_12534,N_13492);
nand U15767 (N_15767,N_12661,N_12285);
nand U15768 (N_15768,N_12371,N_12945);
nand U15769 (N_15769,N_12949,N_13203);
nand U15770 (N_15770,N_12904,N_12044);
nand U15771 (N_15771,N_12762,N_12537);
and U15772 (N_15772,N_13594,N_12139);
and U15773 (N_15773,N_12615,N_12157);
and U15774 (N_15774,N_13842,N_13527);
nor U15775 (N_15775,N_12457,N_13161);
nor U15776 (N_15776,N_13620,N_13245);
nor U15777 (N_15777,N_12910,N_13328);
and U15778 (N_15778,N_12634,N_13949);
and U15779 (N_15779,N_13000,N_13760);
and U15780 (N_15780,N_13066,N_12057);
nor U15781 (N_15781,N_13758,N_12541);
or U15782 (N_15782,N_13309,N_13273);
and U15783 (N_15783,N_13332,N_13346);
nand U15784 (N_15784,N_12575,N_13087);
and U15785 (N_15785,N_12141,N_12308);
nor U15786 (N_15786,N_12302,N_12000);
nor U15787 (N_15787,N_13598,N_13983);
and U15788 (N_15788,N_13953,N_13132);
or U15789 (N_15789,N_12747,N_13198);
nand U15790 (N_15790,N_12805,N_13721);
nand U15791 (N_15791,N_12598,N_13365);
nand U15792 (N_15792,N_13507,N_13657);
nor U15793 (N_15793,N_12532,N_12278);
xnor U15794 (N_15794,N_12569,N_13959);
and U15795 (N_15795,N_12177,N_12945);
or U15796 (N_15796,N_12767,N_13012);
nor U15797 (N_15797,N_12987,N_13315);
nor U15798 (N_15798,N_13525,N_12401);
nand U15799 (N_15799,N_12542,N_12232);
nand U15800 (N_15800,N_12597,N_13135);
nor U15801 (N_15801,N_12360,N_13687);
and U15802 (N_15802,N_12484,N_12782);
nor U15803 (N_15803,N_13128,N_13588);
or U15804 (N_15804,N_12555,N_13076);
and U15805 (N_15805,N_13962,N_13201);
nand U15806 (N_15806,N_12215,N_12401);
nor U15807 (N_15807,N_13145,N_12400);
nand U15808 (N_15808,N_13522,N_13040);
nand U15809 (N_15809,N_13392,N_13620);
nand U15810 (N_15810,N_12974,N_13029);
and U15811 (N_15811,N_12567,N_12378);
and U15812 (N_15812,N_13460,N_13308);
nand U15813 (N_15813,N_13019,N_13629);
and U15814 (N_15814,N_13269,N_13102);
or U15815 (N_15815,N_12436,N_12778);
or U15816 (N_15816,N_12467,N_12724);
nor U15817 (N_15817,N_12213,N_13351);
or U15818 (N_15818,N_12514,N_13883);
or U15819 (N_15819,N_13809,N_13285);
and U15820 (N_15820,N_13299,N_13805);
and U15821 (N_15821,N_13901,N_13445);
or U15822 (N_15822,N_13387,N_12424);
or U15823 (N_15823,N_13264,N_13698);
and U15824 (N_15824,N_13763,N_12213);
nor U15825 (N_15825,N_13544,N_13881);
nor U15826 (N_15826,N_12321,N_13136);
nor U15827 (N_15827,N_13109,N_12590);
or U15828 (N_15828,N_12468,N_12025);
and U15829 (N_15829,N_12185,N_12026);
and U15830 (N_15830,N_13383,N_13430);
nor U15831 (N_15831,N_13448,N_12379);
and U15832 (N_15832,N_12027,N_12553);
nand U15833 (N_15833,N_13328,N_13075);
and U15834 (N_15834,N_12861,N_13392);
nor U15835 (N_15835,N_12585,N_12582);
nor U15836 (N_15836,N_12362,N_13637);
or U15837 (N_15837,N_13840,N_12083);
nor U15838 (N_15838,N_12311,N_13922);
nor U15839 (N_15839,N_12160,N_13070);
and U15840 (N_15840,N_12830,N_13680);
nand U15841 (N_15841,N_12803,N_12084);
nor U15842 (N_15842,N_12124,N_13123);
and U15843 (N_15843,N_13534,N_12104);
nand U15844 (N_15844,N_13632,N_12385);
or U15845 (N_15845,N_12536,N_12020);
or U15846 (N_15846,N_13341,N_13280);
nor U15847 (N_15847,N_13494,N_13056);
or U15848 (N_15848,N_12889,N_13770);
xor U15849 (N_15849,N_12240,N_12500);
or U15850 (N_15850,N_12160,N_12794);
nand U15851 (N_15851,N_13388,N_12556);
or U15852 (N_15852,N_12484,N_13064);
and U15853 (N_15853,N_12336,N_13247);
nand U15854 (N_15854,N_12954,N_12592);
and U15855 (N_15855,N_13482,N_12054);
and U15856 (N_15856,N_13004,N_12588);
nor U15857 (N_15857,N_13902,N_12217);
and U15858 (N_15858,N_12005,N_13030);
and U15859 (N_15859,N_13496,N_13465);
or U15860 (N_15860,N_12245,N_13469);
nor U15861 (N_15861,N_12194,N_12622);
or U15862 (N_15862,N_12959,N_12408);
and U15863 (N_15863,N_13910,N_13647);
and U15864 (N_15864,N_13838,N_12119);
nand U15865 (N_15865,N_13006,N_13690);
and U15866 (N_15866,N_13443,N_12802);
or U15867 (N_15867,N_13193,N_12076);
nor U15868 (N_15868,N_12432,N_13702);
and U15869 (N_15869,N_12782,N_13749);
or U15870 (N_15870,N_12137,N_13301);
and U15871 (N_15871,N_13978,N_12544);
nand U15872 (N_15872,N_12509,N_12281);
and U15873 (N_15873,N_12057,N_12656);
or U15874 (N_15874,N_12336,N_12896);
or U15875 (N_15875,N_12815,N_13397);
nand U15876 (N_15876,N_13431,N_12823);
nor U15877 (N_15877,N_13139,N_13593);
nand U15878 (N_15878,N_12176,N_13565);
or U15879 (N_15879,N_13433,N_13587);
and U15880 (N_15880,N_12172,N_12369);
or U15881 (N_15881,N_13726,N_12347);
and U15882 (N_15882,N_12718,N_13742);
nor U15883 (N_15883,N_13746,N_13208);
nor U15884 (N_15884,N_13134,N_12508);
nor U15885 (N_15885,N_12971,N_13705);
and U15886 (N_15886,N_12064,N_12016);
nor U15887 (N_15887,N_13886,N_12745);
or U15888 (N_15888,N_13279,N_12137);
and U15889 (N_15889,N_13653,N_13629);
nand U15890 (N_15890,N_13350,N_12125);
and U15891 (N_15891,N_13821,N_12693);
or U15892 (N_15892,N_13262,N_13567);
nor U15893 (N_15893,N_13991,N_13717);
nand U15894 (N_15894,N_13423,N_12172);
nor U15895 (N_15895,N_12362,N_13823);
nand U15896 (N_15896,N_13003,N_12832);
xnor U15897 (N_15897,N_13738,N_12453);
nand U15898 (N_15898,N_13953,N_13742);
nand U15899 (N_15899,N_12312,N_13520);
or U15900 (N_15900,N_12271,N_12187);
nor U15901 (N_15901,N_13063,N_12811);
xor U15902 (N_15902,N_13019,N_13556);
nand U15903 (N_15903,N_13494,N_12879);
and U15904 (N_15904,N_13615,N_13690);
nor U15905 (N_15905,N_13828,N_12987);
or U15906 (N_15906,N_13530,N_12435);
nand U15907 (N_15907,N_13354,N_12528);
nand U15908 (N_15908,N_13272,N_13187);
or U15909 (N_15909,N_13455,N_13063);
or U15910 (N_15910,N_13540,N_12726);
nand U15911 (N_15911,N_12182,N_13624);
nor U15912 (N_15912,N_13999,N_13366);
and U15913 (N_15913,N_12863,N_12903);
or U15914 (N_15914,N_12971,N_12773);
nor U15915 (N_15915,N_13760,N_13925);
or U15916 (N_15916,N_13563,N_12318);
nor U15917 (N_15917,N_12312,N_13171);
nand U15918 (N_15918,N_13913,N_12939);
or U15919 (N_15919,N_13889,N_13613);
or U15920 (N_15920,N_13792,N_12831);
or U15921 (N_15921,N_12442,N_13870);
and U15922 (N_15922,N_12439,N_13498);
or U15923 (N_15923,N_13030,N_12119);
or U15924 (N_15924,N_13317,N_12734);
or U15925 (N_15925,N_12235,N_12329);
nand U15926 (N_15926,N_12081,N_13462);
nand U15927 (N_15927,N_12732,N_12989);
or U15928 (N_15928,N_12384,N_12553);
nand U15929 (N_15929,N_13160,N_12262);
or U15930 (N_15930,N_13163,N_12643);
nand U15931 (N_15931,N_13068,N_12922);
nor U15932 (N_15932,N_12395,N_13528);
nor U15933 (N_15933,N_13138,N_13929);
nor U15934 (N_15934,N_13248,N_12546);
xor U15935 (N_15935,N_12506,N_12781);
and U15936 (N_15936,N_12482,N_12411);
nor U15937 (N_15937,N_12821,N_13920);
nand U15938 (N_15938,N_12616,N_12806);
and U15939 (N_15939,N_12314,N_12304);
and U15940 (N_15940,N_13946,N_12420);
nand U15941 (N_15941,N_13101,N_12726);
or U15942 (N_15942,N_12680,N_12484);
nand U15943 (N_15943,N_13325,N_12216);
and U15944 (N_15944,N_12969,N_12563);
nand U15945 (N_15945,N_13624,N_12870);
and U15946 (N_15946,N_12093,N_13636);
nor U15947 (N_15947,N_12129,N_13840);
or U15948 (N_15948,N_13556,N_12340);
and U15949 (N_15949,N_13084,N_12674);
nand U15950 (N_15950,N_13339,N_13935);
nor U15951 (N_15951,N_13710,N_12629);
nand U15952 (N_15952,N_12502,N_13769);
and U15953 (N_15953,N_12507,N_12171);
and U15954 (N_15954,N_13142,N_12540);
nor U15955 (N_15955,N_12759,N_13074);
nor U15956 (N_15956,N_12281,N_12839);
and U15957 (N_15957,N_12344,N_12339);
nand U15958 (N_15958,N_13161,N_12521);
or U15959 (N_15959,N_13040,N_12041);
and U15960 (N_15960,N_13900,N_12301);
and U15961 (N_15961,N_12173,N_12393);
or U15962 (N_15962,N_12559,N_12629);
nand U15963 (N_15963,N_13670,N_13524);
and U15964 (N_15964,N_13432,N_12684);
nor U15965 (N_15965,N_12967,N_13350);
nor U15966 (N_15966,N_12907,N_13638);
nand U15967 (N_15967,N_12917,N_13090);
or U15968 (N_15968,N_13632,N_13309);
nand U15969 (N_15969,N_12389,N_13384);
and U15970 (N_15970,N_12240,N_12234);
or U15971 (N_15971,N_13625,N_12028);
and U15972 (N_15972,N_13342,N_13824);
and U15973 (N_15973,N_12410,N_13315);
or U15974 (N_15974,N_13731,N_13903);
nand U15975 (N_15975,N_12225,N_12200);
nor U15976 (N_15976,N_12308,N_12911);
nor U15977 (N_15977,N_13268,N_13375);
nor U15978 (N_15978,N_13918,N_12304);
and U15979 (N_15979,N_13689,N_12849);
and U15980 (N_15980,N_13445,N_12956);
nor U15981 (N_15981,N_12051,N_12037);
nor U15982 (N_15982,N_12766,N_12437);
and U15983 (N_15983,N_13835,N_12264);
or U15984 (N_15984,N_13860,N_12158);
and U15985 (N_15985,N_13340,N_12780);
nand U15986 (N_15986,N_12068,N_12559);
nand U15987 (N_15987,N_12746,N_12481);
nor U15988 (N_15988,N_13489,N_13401);
or U15989 (N_15989,N_13024,N_13585);
nand U15990 (N_15990,N_12646,N_13601);
or U15991 (N_15991,N_13943,N_12702);
nand U15992 (N_15992,N_13032,N_12675);
nor U15993 (N_15993,N_12622,N_13065);
nand U15994 (N_15994,N_13407,N_13866);
or U15995 (N_15995,N_12753,N_12276);
nand U15996 (N_15996,N_13919,N_13578);
nor U15997 (N_15997,N_13633,N_13550);
nand U15998 (N_15998,N_12452,N_13535);
nor U15999 (N_15999,N_12671,N_12657);
nor U16000 (N_16000,N_15042,N_14959);
nor U16001 (N_16001,N_14188,N_14659);
nor U16002 (N_16002,N_14708,N_14610);
or U16003 (N_16003,N_14908,N_15041);
nand U16004 (N_16004,N_14231,N_14912);
nor U16005 (N_16005,N_14219,N_14596);
nand U16006 (N_16006,N_15023,N_14128);
nor U16007 (N_16007,N_15822,N_15239);
or U16008 (N_16008,N_14005,N_14733);
and U16009 (N_16009,N_15353,N_15018);
or U16010 (N_16010,N_14837,N_14754);
nand U16011 (N_16011,N_15801,N_15603);
nor U16012 (N_16012,N_14558,N_14867);
or U16013 (N_16013,N_15676,N_15745);
nor U16014 (N_16014,N_15525,N_15807);
or U16015 (N_16015,N_15918,N_15098);
nor U16016 (N_16016,N_15794,N_15096);
and U16017 (N_16017,N_14215,N_14491);
or U16018 (N_16018,N_15003,N_15388);
nand U16019 (N_16019,N_14429,N_15590);
nor U16020 (N_16020,N_14747,N_14858);
or U16021 (N_16021,N_15437,N_15470);
nor U16022 (N_16022,N_14566,N_15981);
or U16023 (N_16023,N_15117,N_15644);
or U16024 (N_16024,N_15521,N_14939);
nand U16025 (N_16025,N_15138,N_15402);
nand U16026 (N_16026,N_14518,N_15725);
or U16027 (N_16027,N_15899,N_14926);
or U16028 (N_16028,N_15963,N_15548);
nor U16029 (N_16029,N_15333,N_15339);
nand U16030 (N_16030,N_14704,N_14412);
nand U16031 (N_16031,N_14721,N_14540);
nor U16032 (N_16032,N_15379,N_15244);
nand U16033 (N_16033,N_15088,N_15990);
nand U16034 (N_16034,N_14948,N_15334);
nand U16035 (N_16035,N_14725,N_15208);
nand U16036 (N_16036,N_15457,N_15775);
nor U16037 (N_16037,N_14986,N_15874);
and U16038 (N_16038,N_14451,N_14592);
nand U16039 (N_16039,N_14149,N_15136);
nor U16040 (N_16040,N_15202,N_14668);
nor U16041 (N_16041,N_14812,N_15558);
and U16042 (N_16042,N_14861,N_15902);
xnor U16043 (N_16043,N_14306,N_15130);
nand U16044 (N_16044,N_14878,N_14587);
nor U16045 (N_16045,N_14119,N_14259);
nor U16046 (N_16046,N_15272,N_14515);
or U16047 (N_16047,N_15040,N_14390);
nand U16048 (N_16048,N_14968,N_14262);
and U16049 (N_16049,N_14041,N_14370);
nand U16050 (N_16050,N_15375,N_14321);
nand U16051 (N_16051,N_15795,N_14696);
nand U16052 (N_16052,N_14473,N_15120);
or U16053 (N_16053,N_14862,N_15915);
or U16054 (N_16054,N_14474,N_15620);
or U16055 (N_16055,N_14191,N_14143);
nor U16056 (N_16056,N_15116,N_14138);
nand U16057 (N_16057,N_15065,N_14172);
nor U16058 (N_16058,N_14101,N_15154);
nand U16059 (N_16059,N_14165,N_15103);
nor U16060 (N_16060,N_15496,N_15193);
nand U16061 (N_16061,N_14365,N_15783);
nand U16062 (N_16062,N_15473,N_14269);
and U16063 (N_16063,N_14726,N_15081);
and U16064 (N_16064,N_14007,N_14360);
nand U16065 (N_16065,N_14617,N_15476);
nand U16066 (N_16066,N_14109,N_14573);
and U16067 (N_16067,N_14205,N_14913);
nor U16068 (N_16068,N_14675,N_14834);
nand U16069 (N_16069,N_14546,N_15812);
and U16070 (N_16070,N_15692,N_15764);
nand U16071 (N_16071,N_15786,N_15967);
nand U16072 (N_16072,N_15084,N_15734);
nand U16073 (N_16073,N_14703,N_15100);
or U16074 (N_16074,N_15598,N_14588);
or U16075 (N_16075,N_15608,N_15937);
and U16076 (N_16076,N_14386,N_14485);
nor U16077 (N_16077,N_15210,N_14871);
and U16078 (N_16078,N_14795,N_14481);
and U16079 (N_16079,N_14380,N_15415);
nand U16080 (N_16080,N_14411,N_14802);
or U16081 (N_16081,N_14415,N_14970);
and U16082 (N_16082,N_14560,N_14161);
nand U16083 (N_16083,N_14100,N_14953);
or U16084 (N_16084,N_14103,N_15724);
and U16085 (N_16085,N_15428,N_14378);
and U16086 (N_16086,N_14294,N_14649);
nand U16087 (N_16087,N_14579,N_15896);
or U16088 (N_16088,N_15176,N_14001);
and U16089 (N_16089,N_14826,N_14775);
nand U16090 (N_16090,N_15566,N_15797);
or U16091 (N_16091,N_14767,N_14062);
nor U16092 (N_16092,N_14801,N_15925);
nor U16093 (N_16093,N_14264,N_14927);
xnor U16094 (N_16094,N_15730,N_14771);
or U16095 (N_16095,N_15221,N_14655);
and U16096 (N_16096,N_15622,N_14279);
xor U16097 (N_16097,N_14718,N_14176);
and U16098 (N_16098,N_14192,N_14366);
and U16099 (N_16099,N_15431,N_14050);
nor U16100 (N_16100,N_15557,N_14142);
nor U16101 (N_16101,N_14432,N_15816);
and U16102 (N_16102,N_14002,N_15288);
and U16103 (N_16103,N_14293,N_14427);
and U16104 (N_16104,N_15107,N_15573);
nor U16105 (N_16105,N_15790,N_14152);
or U16106 (N_16106,N_14909,N_14436);
nand U16107 (N_16107,N_15593,N_14541);
nor U16108 (N_16108,N_15440,N_14538);
and U16109 (N_16109,N_15450,N_14509);
or U16110 (N_16110,N_14793,N_15867);
nor U16111 (N_16111,N_14200,N_14778);
nand U16112 (N_16112,N_14028,N_14097);
nor U16113 (N_16113,N_15094,N_15536);
nor U16114 (N_16114,N_14032,N_15849);
and U16115 (N_16115,N_14875,N_15382);
or U16116 (N_16116,N_14717,N_14864);
and U16117 (N_16117,N_15840,N_14088);
nor U16118 (N_16118,N_14449,N_14608);
or U16119 (N_16119,N_14236,N_14283);
or U16120 (N_16120,N_15549,N_14693);
nor U16121 (N_16121,N_14616,N_15389);
or U16122 (N_16122,N_15323,N_15973);
nor U16123 (N_16123,N_14857,N_14877);
nand U16124 (N_16124,N_14990,N_14995);
nand U16125 (N_16125,N_14214,N_15351);
or U16126 (N_16126,N_14140,N_15747);
nor U16127 (N_16127,N_14460,N_14487);
or U16128 (N_16128,N_14414,N_15252);
nand U16129 (N_16129,N_14590,N_15662);
or U16130 (N_16130,N_15586,N_14393);
or U16131 (N_16131,N_15327,N_14835);
nor U16132 (N_16132,N_14237,N_14510);
nand U16133 (N_16133,N_15577,N_15019);
nor U16134 (N_16134,N_15992,N_14500);
nor U16135 (N_16135,N_15913,N_15308);
and U16136 (N_16136,N_14893,N_15196);
and U16137 (N_16137,N_15599,N_15302);
or U16138 (N_16138,N_15419,N_15984);
or U16139 (N_16139,N_14830,N_14578);
nand U16140 (N_16140,N_15988,N_14863);
or U16141 (N_16141,N_14357,N_15082);
nand U16142 (N_16142,N_14288,N_15928);
and U16143 (N_16143,N_15032,N_15987);
or U16144 (N_16144,N_15448,N_14484);
nor U16145 (N_16145,N_14364,N_14713);
or U16146 (N_16146,N_14853,N_14091);
nor U16147 (N_16147,N_15506,N_15818);
nand U16148 (N_16148,N_14526,N_14544);
or U16149 (N_16149,N_14054,N_15943);
nor U16150 (N_16150,N_15850,N_14804);
and U16151 (N_16151,N_15109,N_14599);
and U16152 (N_16152,N_14277,N_14439);
or U16153 (N_16153,N_14208,N_14823);
nor U16154 (N_16154,N_14533,N_15634);
or U16155 (N_16155,N_15214,N_15534);
nor U16156 (N_16156,N_14320,N_15270);
nand U16157 (N_16157,N_14446,N_14388);
or U16158 (N_16158,N_15736,N_14348);
nor U16159 (N_16159,N_14160,N_15097);
nand U16160 (N_16160,N_14465,N_15106);
and U16161 (N_16161,N_14682,N_15505);
or U16162 (N_16162,N_15914,N_15746);
or U16163 (N_16163,N_15962,N_15219);
and U16164 (N_16164,N_15134,N_14477);
and U16165 (N_16165,N_14574,N_15254);
or U16166 (N_16166,N_15364,N_15013);
nand U16167 (N_16167,N_14313,N_15520);
or U16168 (N_16168,N_15187,N_15365);
or U16169 (N_16169,N_14445,N_14911);
or U16170 (N_16170,N_14016,N_15059);
and U16171 (N_16171,N_15459,N_15901);
nand U16172 (N_16172,N_14554,N_15828);
nand U16173 (N_16173,N_15631,N_14282);
or U16174 (N_16174,N_15737,N_15971);
nor U16175 (N_16175,N_14023,N_15927);
or U16176 (N_16176,N_15649,N_14611);
nand U16177 (N_16177,N_14121,N_15556);
and U16178 (N_16178,N_14698,N_14132);
nand U16179 (N_16179,N_15063,N_14168);
or U16180 (N_16180,N_14255,N_14890);
and U16181 (N_16181,N_14821,N_14941);
and U16182 (N_16182,N_15378,N_14490);
nor U16183 (N_16183,N_14329,N_15658);
nor U16184 (N_16184,N_15681,N_15894);
nor U16185 (N_16185,N_15882,N_14692);
nor U16186 (N_16186,N_14431,N_14768);
nand U16187 (N_16187,N_14331,N_15145);
nand U16188 (N_16188,N_15263,N_14466);
and U16189 (N_16189,N_14618,N_14117);
nor U16190 (N_16190,N_14094,N_15251);
nor U16191 (N_16191,N_15183,N_15515);
nor U16192 (N_16192,N_14918,N_15555);
nand U16193 (N_16193,N_15144,N_15685);
nand U16194 (N_16194,N_15160,N_15275);
nor U16195 (N_16195,N_14225,N_15741);
and U16196 (N_16196,N_14268,N_15424);
or U16197 (N_16197,N_14632,N_14372);
nor U16198 (N_16198,N_14650,N_15953);
and U16199 (N_16199,N_14104,N_15640);
nor U16200 (N_16200,N_14882,N_14010);
and U16201 (N_16201,N_14253,N_14563);
nand U16202 (N_16202,N_15695,N_15427);
or U16203 (N_16203,N_14936,N_15934);
or U16204 (N_16204,N_14345,N_15854);
nor U16205 (N_16205,N_15209,N_15195);
or U16206 (N_16206,N_14102,N_14951);
or U16207 (N_16207,N_14346,N_14794);
or U16208 (N_16208,N_14433,N_15580);
and U16209 (N_16209,N_15680,N_15921);
or U16210 (N_16210,N_14800,N_15380);
and U16211 (N_16211,N_14731,N_14772);
or U16212 (N_16212,N_15115,N_15618);
or U16213 (N_16213,N_14084,N_15889);
or U16214 (N_16214,N_14956,N_14782);
or U16215 (N_16215,N_14565,N_15529);
and U16216 (N_16216,N_14620,N_15340);
and U16217 (N_16217,N_15814,N_15859);
or U16218 (N_16218,N_15728,N_14919);
or U16219 (N_16219,N_14859,N_15666);
nor U16220 (N_16220,N_15488,N_14110);
nand U16221 (N_16221,N_14250,N_15776);
nand U16222 (N_16222,N_14443,N_14315);
nand U16223 (N_16223,N_15164,N_14979);
and U16224 (N_16224,N_14124,N_14764);
nor U16225 (N_16225,N_15985,N_14706);
or U16226 (N_16226,N_14932,N_14502);
nand U16227 (N_16227,N_15352,N_14737);
or U16228 (N_16228,N_15014,N_15876);
nand U16229 (N_16229,N_15661,N_14811);
nand U16230 (N_16230,N_14732,N_14855);
or U16231 (N_16231,N_15390,N_14261);
nor U16232 (N_16232,N_14568,N_14266);
nor U16233 (N_16233,N_14749,N_14173);
or U16234 (N_16234,N_15011,N_15757);
or U16235 (N_16235,N_14923,N_14082);
and U16236 (N_16236,N_14644,N_14730);
nor U16237 (N_16237,N_14711,N_14111);
or U16238 (N_16238,N_15223,N_14786);
nor U16239 (N_16239,N_14743,N_14906);
nor U16240 (N_16240,N_15030,N_14729);
and U16241 (N_16241,N_15768,N_15702);
nor U16242 (N_16242,N_15931,N_15245);
or U16243 (N_16243,N_15989,N_15460);
nand U16244 (N_16244,N_14507,N_15941);
or U16245 (N_16245,N_15262,N_14963);
and U16246 (N_16246,N_15242,N_14946);
nor U16247 (N_16247,N_14435,N_15501);
nand U16248 (N_16248,N_14419,N_14854);
nand U16249 (N_16249,N_14162,N_14265);
or U16250 (N_16250,N_15182,N_15968);
nand U16251 (N_16251,N_14263,N_15298);
nor U16252 (N_16252,N_15975,N_14238);
or U16253 (N_16253,N_14816,N_14006);
nor U16254 (N_16254,N_14407,N_15759);
nand U16255 (N_16255,N_15192,N_15163);
or U16256 (N_16256,N_14137,N_14326);
nor U16257 (N_16257,N_15713,N_14420);
or U16258 (N_16258,N_15624,N_14080);
or U16259 (N_16259,N_15143,N_14305);
nor U16260 (N_16260,N_15360,N_15838);
and U16261 (N_16261,N_14133,N_14907);
or U16262 (N_16262,N_15717,N_14874);
and U16263 (N_16263,N_14086,N_14457);
or U16264 (N_16264,N_15295,N_15420);
or U16265 (N_16265,N_14651,N_15587);
or U16266 (N_16266,N_14513,N_14150);
and U16267 (N_16267,N_14202,N_14680);
and U16268 (N_16268,N_14889,N_15315);
nor U16269 (N_16269,N_14008,N_15655);
nor U16270 (N_16270,N_15504,N_15386);
nor U16271 (N_16271,N_14003,N_15359);
nor U16272 (N_16272,N_14580,N_14840);
and U16273 (N_16273,N_14634,N_14130);
nand U16274 (N_16274,N_15951,N_15070);
and U16275 (N_16275,N_15132,N_14781);
or U16276 (N_16276,N_15118,N_15810);
or U16277 (N_16277,N_15220,N_15743);
nor U16278 (N_16278,N_15227,N_15682);
and U16279 (N_16279,N_14021,N_15799);
nor U16280 (N_16280,N_15231,N_14595);
nand U16281 (N_16281,N_14604,N_15922);
or U16282 (N_16282,N_14181,N_15996);
and U16283 (N_16283,N_15819,N_15016);
or U16284 (N_16284,N_14447,N_14280);
or U16285 (N_16285,N_15399,N_15878);
nor U16286 (N_16286,N_15756,N_15170);
nand U16287 (N_16287,N_14702,N_15835);
nand U16288 (N_16288,N_14289,N_14019);
or U16289 (N_16289,N_15654,N_15924);
nor U16290 (N_16290,N_14850,N_15146);
or U16291 (N_16291,N_14085,N_14543);
nor U16292 (N_16292,N_14391,N_15129);
nor U16293 (N_16293,N_14641,N_14645);
nand U16294 (N_16294,N_15369,N_14482);
or U16295 (N_16295,N_14803,N_14516);
nand U16296 (N_16296,N_15621,N_15900);
and U16297 (N_16297,N_14083,N_14093);
or U16298 (N_16298,N_14339,N_14492);
nor U16299 (N_16299,N_15821,N_15303);
and U16300 (N_16300,N_15524,N_15248);
nor U16301 (N_16301,N_14969,N_14809);
nor U16302 (N_16302,N_14359,N_15543);
nand U16303 (N_16303,N_15372,N_14309);
and U16304 (N_16304,N_15993,N_14066);
nand U16305 (N_16305,N_14052,N_15320);
nor U16306 (N_16306,N_15995,N_15074);
and U16307 (N_16307,N_15553,N_15665);
nand U16308 (N_16308,N_15149,N_14697);
or U16309 (N_16309,N_15343,N_14709);
nand U16310 (N_16310,N_14351,N_15688);
or U16311 (N_16311,N_15647,N_14937);
or U16312 (N_16312,N_15212,N_15385);
nand U16313 (N_16313,N_14405,N_14349);
nor U16314 (N_16314,N_15413,N_15811);
or U16315 (N_16315,N_15766,N_15178);
or U16316 (N_16316,N_14413,N_15443);
nand U16317 (N_16317,N_14243,N_15526);
nand U16318 (N_16318,N_14136,N_15704);
nor U16319 (N_16319,N_15346,N_14756);
nor U16320 (N_16320,N_15997,N_14727);
or U16321 (N_16321,N_14135,N_15090);
nand U16322 (N_16322,N_15628,N_15294);
nor U16323 (N_16323,N_14389,N_14623);
or U16324 (N_16324,N_14735,N_15978);
nand U16325 (N_16325,N_14656,N_14057);
nand U16326 (N_16326,N_14227,N_15228);
nor U16327 (N_16327,N_15514,N_15157);
nand U16328 (N_16328,N_14015,N_15664);
and U16329 (N_16329,N_14751,N_14824);
nand U16330 (N_16330,N_15260,N_14493);
or U16331 (N_16331,N_14661,N_15397);
nand U16332 (N_16332,N_14978,N_14636);
and U16333 (N_16333,N_15261,N_14209);
nand U16334 (N_16334,N_15847,N_14159);
or U16335 (N_16335,N_14387,N_14640);
and U16336 (N_16336,N_14187,N_15305);
nor U16337 (N_16337,N_14417,N_14361);
and U16338 (N_16338,N_14684,N_15562);
nand U16339 (N_16339,N_15559,N_14637);
nand U16340 (N_16340,N_14017,N_15255);
nand U16341 (N_16341,N_15336,N_15276);
and U16342 (N_16342,N_14553,N_14865);
or U16343 (N_16343,N_14814,N_14228);
or U16344 (N_16344,N_15020,N_14042);
nand U16345 (N_16345,N_15366,N_15158);
and U16346 (N_16346,N_14998,N_15449);
or U16347 (N_16347,N_15863,N_15919);
nor U16348 (N_16348,N_15108,N_14459);
and U16349 (N_16349,N_15721,N_14131);
and U16350 (N_16350,N_14683,N_14317);
nand U16351 (N_16351,N_15815,N_14434);
nor U16352 (N_16352,N_14822,N_14025);
nor U16353 (N_16353,N_14197,N_15588);
and U16354 (N_16354,N_15738,N_15024);
and U16355 (N_16355,N_15763,N_15509);
nand U16356 (N_16356,N_14099,N_15483);
nand U16357 (N_16357,N_14755,N_14256);
and U16358 (N_16358,N_15328,N_14489);
xnor U16359 (N_16359,N_15304,N_14815);
or U16360 (N_16360,N_14367,N_15279);
and U16361 (N_16361,N_14601,N_15619);
and U16362 (N_16362,N_14354,N_15545);
and U16363 (N_16363,N_14217,N_15857);
nor U16364 (N_16364,N_15769,N_14338);
or U16365 (N_16365,N_15762,N_14190);
and U16366 (N_16366,N_14053,N_14886);
or U16367 (N_16367,N_15958,N_14750);
nor U16368 (N_16368,N_15405,N_14638);
and U16369 (N_16369,N_15007,N_15241);
xor U16370 (N_16370,N_14462,N_14375);
nand U16371 (N_16371,N_14072,N_14895);
or U16372 (N_16372,N_15885,N_15139);
nor U16373 (N_16373,N_15249,N_15773);
nand U16374 (N_16374,N_15886,N_15701);
nor U16375 (N_16375,N_14004,N_15581);
nor U16376 (N_16376,N_15433,N_14146);
or U16377 (N_16377,N_14189,N_14258);
and U16378 (N_16378,N_14274,N_15152);
nor U16379 (N_16379,N_15319,N_15870);
nor U16380 (N_16380,N_15168,N_14198);
nand U16381 (N_16381,N_14746,N_15151);
or U16382 (N_16382,N_15920,N_14308);
nand U16383 (N_16383,N_15265,N_14527);
nor U16384 (N_16384,N_15156,N_15641);
nor U16385 (N_16385,N_15435,N_15726);
or U16386 (N_16386,N_14307,N_15530);
and U16387 (N_16387,N_15770,N_15974);
nand U16388 (N_16388,N_14058,N_15938);
or U16389 (N_16389,N_15837,N_14043);
nand U16390 (N_16390,N_14270,N_15078);
or U16391 (N_16391,N_14896,N_15284);
nor U16392 (N_16392,N_15771,N_15462);
or U16393 (N_16393,N_15479,N_14056);
and U16394 (N_16394,N_14866,N_15945);
or U16395 (N_16395,N_15412,N_15293);
or U16396 (N_16396,N_14783,N_15213);
and U16397 (N_16397,N_14037,N_14224);
nor U16398 (N_16398,N_15401,N_14728);
or U16399 (N_16399,N_14127,N_14770);
nor U16400 (N_16400,N_14744,N_14839);
and U16401 (N_16401,N_14833,N_15637);
nor U16402 (N_16402,N_14720,N_15817);
and U16403 (N_16403,N_14440,N_15888);
and U16404 (N_16404,N_15689,N_15053);
nor U16405 (N_16405,N_15377,N_15777);
or U16406 (N_16406,N_14593,N_15595);
nand U16407 (N_16407,N_14660,N_15426);
or U16408 (N_16408,N_14324,N_14070);
and U16409 (N_16409,N_15691,N_14705);
nor U16410 (N_16410,N_14810,N_15949);
or U16411 (N_16411,N_15273,N_14201);
nand U16412 (N_16412,N_14472,N_14983);
and U16413 (N_16413,N_15578,N_15696);
nor U16414 (N_16414,N_15511,N_15936);
or U16415 (N_16415,N_15012,N_14156);
nor U16416 (N_16416,N_15001,N_14022);
or U16417 (N_16417,N_15602,N_14860);
nand U16418 (N_16418,N_15610,N_15036);
nand U16419 (N_16419,N_15086,N_15186);
and U16420 (N_16420,N_14395,N_14891);
or U16421 (N_16421,N_14922,N_14561);
and U16422 (N_16422,N_15856,N_14597);
or U16423 (N_16423,N_15607,N_15475);
nor U16424 (N_16424,N_15191,N_14557);
or U16425 (N_16425,N_15029,N_15583);
nand U16426 (N_16426,N_15535,N_15541);
nand U16427 (N_16427,N_15684,N_14991);
nand U16428 (N_16428,N_15446,N_14758);
or U16429 (N_16429,N_14676,N_14233);
and U16430 (N_16430,N_15652,N_14379);
or U16431 (N_16431,N_15947,N_15224);
or U16432 (N_16432,N_14461,N_15616);
nand U16433 (N_16433,N_14679,N_14843);
nand U16434 (N_16434,N_14740,N_14079);
or U16435 (N_16435,N_14455,N_14504);
nor U16436 (N_16436,N_14757,N_15111);
or U16437 (N_16437,N_15820,N_14397);
or U16438 (N_16438,N_14899,N_14126);
or U16439 (N_16439,N_14399,N_14673);
and U16440 (N_16440,N_14444,N_15406);
and U16441 (N_16441,N_14322,N_14615);
nand U16442 (N_16442,N_15394,N_15671);
and U16443 (N_16443,N_14602,N_14511);
nand U16444 (N_16444,N_15230,N_15335);
nor U16445 (N_16445,N_15274,N_15675);
or U16446 (N_16446,N_15056,N_15050);
nor U16447 (N_16447,N_14993,N_14063);
and U16448 (N_16448,N_15961,N_14020);
and U16449 (N_16449,N_14404,N_14068);
or U16450 (N_16450,N_14869,N_15080);
or U16451 (N_16451,N_15396,N_15141);
or U16452 (N_16452,N_15229,N_15269);
or U16453 (N_16453,N_15656,N_14373);
or U16454 (N_16454,N_15128,N_14218);
and U16455 (N_16455,N_15999,N_15357);
or U16456 (N_16456,N_15546,N_14416);
or U16457 (N_16457,N_15233,N_15179);
nor U16458 (N_16458,N_15418,N_14738);
and U16459 (N_16459,N_15374,N_15875);
or U16460 (N_16460,N_14591,N_15166);
xor U16461 (N_16461,N_15916,N_15347);
or U16462 (N_16462,N_14067,N_14807);
nand U16463 (N_16463,N_15678,N_15648);
nor U16464 (N_16464,N_14323,N_14271);
nor U16465 (N_16465,N_14776,N_15071);
nand U16466 (N_16466,N_15632,N_14163);
nor U16467 (N_16467,N_14508,N_14522);
nor U16468 (N_16468,N_15006,N_14710);
or U16469 (N_16469,N_15547,N_15271);
nand U16470 (N_16470,N_15832,N_15309);
and U16471 (N_16471,N_15868,N_14987);
and U16472 (N_16472,N_14402,N_14545);
nand U16473 (N_16473,N_14957,N_15986);
nand U16474 (N_16474,N_14988,N_14343);
and U16475 (N_16475,N_14030,N_14520);
nor U16476 (N_16476,N_15940,N_14276);
nand U16477 (N_16477,N_15722,N_14355);
nand U16478 (N_16478,N_15533,N_14362);
and U16479 (N_16479,N_15126,N_15732);
or U16480 (N_16480,N_14619,N_15864);
or U16481 (N_16481,N_15564,N_14235);
or U16482 (N_16482,N_14938,N_15492);
and U16483 (N_16483,N_15860,N_15234);
or U16484 (N_16484,N_14630,N_15839);
or U16485 (N_16485,N_14870,N_15027);
nor U16486 (N_16486,N_14844,N_14442);
and U16487 (N_16487,N_15257,N_14382);
and U16488 (N_16488,N_15091,N_15760);
and U16489 (N_16489,N_14894,N_15341);
and U16490 (N_16490,N_14048,N_15058);
nor U16491 (N_16491,N_14049,N_14248);
nand U16492 (N_16492,N_14542,N_14628);
nor U16493 (N_16493,N_15465,N_15758);
and U16494 (N_16494,N_14752,N_14700);
nor U16495 (N_16495,N_15697,N_14852);
xor U16496 (N_16496,N_14064,N_14944);
or U16497 (N_16497,N_14183,N_15625);
and U16498 (N_16498,N_14027,N_15171);
and U16499 (N_16499,N_15976,N_15826);
or U16500 (N_16500,N_14966,N_15398);
or U16501 (N_16501,N_15453,N_15709);
nor U16502 (N_16502,N_15055,N_15663);
nand U16503 (N_16503,N_14977,N_14920);
nand U16504 (N_16504,N_15466,N_15392);
nand U16505 (N_16505,N_15674,N_15623);
and U16506 (N_16506,N_15148,N_15079);
or U16507 (N_16507,N_15190,N_14040);
nand U16508 (N_16508,N_15329,N_14376);
or U16509 (N_16509,N_14494,N_14363);
nor U16510 (N_16510,N_15381,N_15004);
nor U16511 (N_16511,N_15487,N_15932);
nand U16512 (N_16512,N_15296,N_15517);
nor U16513 (N_16513,N_14425,N_14295);
nor U16514 (N_16514,N_15076,N_15606);
nor U16515 (N_16515,N_15322,N_15708);
xnor U16516 (N_16516,N_15824,N_14199);
and U16517 (N_16517,N_15869,N_15354);
and U16518 (N_16518,N_14196,N_14910);
or U16519 (N_16519,N_14879,N_15836);
nand U16520 (N_16520,N_15280,N_15613);
or U16521 (N_16521,N_15668,N_14984);
or U16522 (N_16522,N_15643,N_14069);
or U16523 (N_16523,N_14626,N_15044);
or U16524 (N_16524,N_14796,N_15751);
or U16525 (N_16525,N_15189,N_14724);
or U16526 (N_16526,N_15314,N_14643);
or U16527 (N_16527,N_15253,N_15403);
and U16528 (N_16528,N_14169,N_15387);
xnor U16529 (N_16529,N_14642,N_15877);
nand U16530 (N_16530,N_14622,N_14765);
nor U16531 (N_16531,N_15125,N_14471);
nor U16532 (N_16532,N_15710,N_15017);
and U16533 (N_16533,N_15539,N_14836);
nor U16534 (N_16534,N_14352,N_14564);
or U16535 (N_16535,N_14213,N_15008);
and U16536 (N_16536,N_15247,N_14092);
or U16537 (N_16537,N_14337,N_14779);
or U16538 (N_16538,N_14774,N_15672);
and U16539 (N_16539,N_15235,N_15414);
nand U16540 (N_16540,N_15358,N_14577);
or U16541 (N_16541,N_15800,N_15218);
and U16542 (N_16542,N_15310,N_15421);
or U16543 (N_16543,N_15646,N_15142);
and U16544 (N_16544,N_14635,N_15423);
nand U16545 (N_16545,N_15754,N_14029);
and U16546 (N_16546,N_14333,N_14689);
or U16547 (N_16547,N_15774,N_15266);
nor U16548 (N_16548,N_14572,N_15324);
or U16549 (N_16549,N_14831,N_14905);
nor U16550 (N_16550,N_15455,N_15707);
nor U16551 (N_16551,N_14467,N_15679);
or U16552 (N_16552,N_14613,N_15808);
or U16553 (N_16553,N_15368,N_15180);
nor U16554 (N_16554,N_14761,N_14498);
nor U16555 (N_16555,N_15225,N_15761);
nor U16556 (N_16556,N_15803,N_15735);
nand U16557 (N_16557,N_15604,N_15851);
nor U16558 (N_16558,N_15285,N_15612);
and U16559 (N_16559,N_15910,N_14917);
nand U16560 (N_16560,N_14887,N_15742);
and U16561 (N_16561,N_14658,N_14701);
and U16562 (N_16562,N_14452,N_15873);
nand U16563 (N_16563,N_15095,N_14845);
or U16564 (N_16564,N_15373,N_15411);
or U16565 (N_16565,N_15893,N_15845);
or U16566 (N_16566,N_14303,N_14076);
or U16567 (N_16567,N_14521,N_15660);
nand U16568 (N_16568,N_14589,N_15300);
and U16569 (N_16569,N_14286,N_14448);
and U16570 (N_16570,N_15485,N_15124);
or U16571 (N_16571,N_15299,N_15174);
nand U16572 (N_16572,N_14164,N_15456);
or U16573 (N_16573,N_14106,N_14739);
and U16574 (N_16574,N_14356,N_14114);
and U16575 (N_16575,N_15325,N_15172);
or U16576 (N_16576,N_15731,N_15898);
nor U16577 (N_16577,N_14598,N_14885);
or U16578 (N_16578,N_15057,N_14244);
or U16579 (N_16579,N_15215,N_14478);
nand U16580 (N_16580,N_15633,N_15830);
and U16581 (N_16581,N_14284,N_15425);
nand U16582 (N_16582,N_14797,N_15463);
nand U16583 (N_16583,N_14657,N_14206);
nor U16584 (N_16584,N_14335,N_14901);
xnor U16585 (N_16585,N_14631,N_14952);
nor U16586 (N_16586,N_14633,N_14234);
and U16587 (N_16587,N_15544,N_14422);
nand U16588 (N_16588,N_14147,N_15054);
or U16589 (N_16589,N_15908,N_15240);
nor U16590 (N_16590,N_15510,N_14898);
nand U16591 (N_16591,N_14145,N_15561);
nand U16592 (N_16592,N_15211,N_14961);
xnor U16593 (N_16593,N_15638,N_15497);
and U16594 (N_16594,N_15286,N_15706);
and U16595 (N_16595,N_14033,N_15935);
or U16596 (N_16596,N_15503,N_15112);
or U16597 (N_16597,N_14394,N_15015);
nor U16598 (N_16598,N_15579,N_15653);
and U16599 (N_16599,N_15923,N_15862);
or U16600 (N_16600,N_15495,N_14787);
nand U16601 (N_16601,N_14344,N_14166);
nand U16602 (N_16602,N_15842,N_14583);
and U16603 (N_16603,N_15667,N_14872);
nor U16604 (N_16604,N_15567,N_14646);
nor U16605 (N_16605,N_15002,N_14074);
nand U16606 (N_16606,N_14061,N_14400);
and U16607 (N_16607,N_14203,N_14975);
nor U16608 (N_16608,N_15025,N_14805);
and U16609 (N_16609,N_15568,N_14496);
or U16610 (N_16610,N_14667,N_15716);
nand U16611 (N_16611,N_15110,N_15611);
or U16612 (N_16612,N_15563,N_14240);
and U16613 (N_16613,N_14994,N_14691);
nand U16614 (N_16614,N_15461,N_14639);
nand U16615 (N_16615,N_15371,N_14418);
nor U16616 (N_16616,N_15683,N_14669);
nor U16617 (N_16617,N_14784,N_14267);
or U16618 (N_16618,N_15045,N_15574);
nor U16619 (N_16619,N_14529,N_14971);
or U16620 (N_16620,N_14275,N_15034);
nand U16621 (N_16621,N_15217,N_15290);
or U16622 (N_16622,N_15767,N_14505);
or U16623 (N_16623,N_15802,N_15184);
xnor U16624 (N_16624,N_15972,N_14819);
nand U16625 (N_16625,N_15400,N_14475);
nand U16626 (N_16626,N_14556,N_15494);
or U16627 (N_16627,N_14059,N_14934);
and U16628 (N_16628,N_15205,N_15306);
and U16629 (N_16629,N_15113,N_14624);
or U16630 (N_16630,N_15391,N_15518);
or U16631 (N_16631,N_15355,N_14330);
and U16632 (N_16632,N_15085,N_15206);
or U16633 (N_16633,N_15010,N_15484);
and U16634 (N_16634,N_14325,N_14464);
and U16635 (N_16635,N_14018,N_15477);
or U16636 (N_16636,N_14385,N_14071);
and U16637 (N_16637,N_14954,N_14534);
nor U16638 (N_16638,N_14759,N_15153);
and U16639 (N_16639,N_14523,N_14828);
nor U16640 (N_16640,N_14229,N_15264);
nor U16641 (N_16641,N_14087,N_14112);
nor U16642 (N_16642,N_15123,N_14654);
or U16643 (N_16643,N_14671,N_15778);
or U16644 (N_16644,N_14653,N_15052);
and U16645 (N_16645,N_14532,N_14065);
nand U16646 (N_16646,N_14401,N_15946);
and U16647 (N_16647,N_14681,N_14585);
and U16648 (N_16648,N_14790,N_14013);
or U16649 (N_16649,N_14962,N_14690);
nor U16650 (N_16650,N_14535,N_14715);
or U16651 (N_16651,N_14848,N_14582);
and U16652 (N_16652,N_15788,N_14047);
and U16653 (N_16653,N_15825,N_15796);
nor U16654 (N_16654,N_15852,N_14549);
and U16655 (N_16655,N_14426,N_14290);
nor U16656 (N_16656,N_15204,N_15150);
and U16657 (N_16657,N_14955,N_15474);
and U16658 (N_16658,N_15283,N_15292);
nand U16659 (N_16659,N_15592,N_14495);
or U16660 (N_16660,N_14141,N_15554);
nand U16661 (N_16661,N_15552,N_14785);
nor U16662 (N_16662,N_14423,N_14753);
xnor U16663 (N_16663,N_14118,N_15693);
nor U16664 (N_16664,N_14999,N_14011);
or U16665 (N_16665,N_14904,N_15383);
or U16666 (N_16666,N_14576,N_14888);
and U16667 (N_16667,N_15912,N_15502);
nand U16668 (N_16668,N_14483,N_14665);
and U16669 (N_16669,N_15119,N_14806);
nand U16670 (N_16670,N_15942,N_14239);
nor U16671 (N_16671,N_15114,N_15642);
and U16672 (N_16672,N_15538,N_14695);
and U16673 (N_16673,N_14627,N_15712);
and U16674 (N_16674,N_14550,N_14925);
nand U16675 (N_16675,N_14531,N_14108);
nand U16676 (N_16676,N_14486,N_15659);
and U16677 (N_16677,N_15855,N_15237);
or U16678 (N_16678,N_15865,N_14369);
or U16679 (N_16679,N_15551,N_14396);
and U16680 (N_16680,N_15445,N_14548);
nand U16681 (N_16681,N_14060,N_15792);
and U16682 (N_16682,N_14122,N_15793);
nand U16683 (N_16683,N_14186,N_14763);
nor U16684 (N_16684,N_15956,N_14943);
nor U16685 (N_16685,N_14972,N_14838);
xnor U16686 (N_16686,N_15441,N_15222);
nor U16687 (N_16687,N_15791,N_15362);
or U16688 (N_16688,N_14629,N_15043);
nor U16689 (N_16689,N_14298,N_15159);
nand U16690 (N_16690,N_14437,N_15570);
or U16691 (N_16691,N_14151,N_15356);
or U16692 (N_16692,N_15363,N_15104);
or U16693 (N_16693,N_15858,N_15532);
or U16694 (N_16694,N_14299,N_15384);
nand U16695 (N_16695,N_14341,N_15733);
nand U16696 (N_16696,N_14868,N_14915);
and U16697 (N_16697,N_14575,N_14144);
nand U16698 (N_16698,N_14945,N_14916);
nand U16699 (N_16699,N_14347,N_15831);
nand U16700 (N_16700,N_15236,N_15991);
xnor U16701 (N_16701,N_15565,N_14982);
nand U16702 (N_16702,N_15926,N_14736);
nor U16703 (N_16703,N_15952,N_14195);
nor U16704 (N_16704,N_15782,N_15313);
nand U16705 (N_16705,N_14662,N_15047);
and U16706 (N_16706,N_15594,N_15954);
or U16707 (N_16707,N_15979,N_14377);
or U16708 (N_16708,N_14381,N_15188);
nor U16709 (N_16709,N_15829,N_15165);
or U16710 (N_16710,N_15201,N_15370);
nor U16711 (N_16711,N_15367,N_14272);
nand U16712 (N_16712,N_14254,N_15349);
nor U16713 (N_16713,N_15167,N_14328);
nor U16714 (N_16714,N_14180,N_15651);
nor U16715 (N_16715,N_15805,N_15307);
nand U16716 (N_16716,N_15844,N_15500);
nand U16717 (N_16717,N_15780,N_14762);
nor U16718 (N_16718,N_15256,N_15585);
or U16719 (N_16719,N_14780,N_14612);
and U16720 (N_16720,N_14552,N_14410);
nand U16721 (N_16721,N_14158,N_14989);
nor U16722 (N_16722,N_15282,N_15438);
and U16723 (N_16723,N_15744,N_14278);
and U16724 (N_16724,N_15584,N_14976);
and U16725 (N_16725,N_14096,N_14035);
nand U16726 (N_16726,N_14678,N_15809);
or U16727 (N_16727,N_15226,N_15035);
nand U16728 (N_16728,N_15291,N_14115);
nand U16729 (N_16729,N_14712,N_14480);
nand U16730 (N_16730,N_14009,N_15571);
and U16731 (N_16731,N_14318,N_15911);
nand U16732 (N_16732,N_15073,N_14211);
and U16733 (N_16733,N_14216,N_14327);
nor U16734 (N_16734,N_14832,N_14567);
nor U16735 (N_16735,N_14469,N_15361);
nand U16736 (N_16736,N_14514,N_14933);
or U16737 (N_16737,N_15326,N_15895);
nand U16738 (N_16738,N_14766,N_14113);
nand U16739 (N_16739,N_14519,N_15853);
nand U16740 (N_16740,N_14134,N_14967);
nand U16741 (N_16741,N_15348,N_14849);
nand U16742 (N_16742,N_14903,N_15458);
and U16743 (N_16743,N_15944,N_15994);
nand U16744 (N_16744,N_14123,N_14045);
nand U16745 (N_16745,N_14409,N_14000);
or U16746 (N_16746,N_15866,N_15444);
and U16747 (N_16747,N_15321,N_15471);
nor U16748 (N_16748,N_15560,N_14012);
and U16749 (N_16749,N_14741,N_15454);
or U16750 (N_16750,N_14929,N_15122);
or U16751 (N_16751,N_14584,N_15137);
and U16752 (N_16752,N_14392,N_14245);
nor U16753 (N_16753,N_14226,N_15629);
or U16754 (N_16754,N_14463,N_14311);
nand U16755 (N_16755,N_14551,N_14078);
or U16756 (N_16756,N_15432,N_15331);
or U16757 (N_16757,N_14421,N_14876);
nor U16758 (N_16758,N_14846,N_15140);
nand U16759 (N_16759,N_15338,N_14300);
xnor U16760 (N_16760,N_14297,N_15410);
and U16761 (N_16761,N_15522,N_15711);
and U16762 (N_16762,N_14536,N_15719);
and U16763 (N_16763,N_14586,N_15903);
or U16764 (N_16764,N_14319,N_14316);
and U16765 (N_16765,N_15977,N_14734);
and U16766 (N_16766,N_14605,N_15033);
xnor U16767 (N_16767,N_14194,N_15022);
nand U16768 (N_16768,N_14827,N_14742);
and U16769 (N_16769,N_14260,N_14207);
nand U16770 (N_16770,N_14251,N_15798);
and U16771 (N_16771,N_14204,N_15089);
nand U16772 (N_16772,N_15481,N_15752);
or U16773 (N_16773,N_14296,N_15469);
or U16774 (N_16774,N_15422,N_15092);
and U16775 (N_16775,N_14095,N_15447);
nor U16776 (N_16776,N_15959,N_15135);
or U16777 (N_16777,N_15246,N_14177);
nor U16778 (N_16778,N_15970,N_15350);
or U16779 (N_16779,N_14688,N_15232);
and U16780 (N_16780,N_14497,N_15700);
nand U16781 (N_16781,N_14090,N_14924);
or U16782 (N_16782,N_15478,N_14788);
and U16783 (N_16783,N_15026,N_14791);
nor U16784 (N_16784,N_14539,N_14981);
and U16785 (N_16785,N_15267,N_14044);
and U16786 (N_16786,N_15442,N_15301);
and U16787 (N_16787,N_15051,N_14829);
nand U16788 (N_16788,N_14880,N_14046);
xor U16789 (N_16789,N_14175,N_14430);
and U16790 (N_16790,N_15203,N_15705);
and U16791 (N_16791,N_14851,N_14892);
and U16792 (N_16792,N_14488,N_15318);
nor U16793 (N_16793,N_15480,N_15527);
and U16794 (N_16794,N_14997,N_15881);
nor U16795 (N_16795,N_14285,N_14073);
nand U16796 (N_16796,N_15173,N_15207);
or U16797 (N_16797,N_15600,N_15905);
nand U16798 (N_16798,N_15243,N_14530);
or U16799 (N_16799,N_15781,N_14773);
and U16800 (N_16800,N_14506,N_14257);
xor U16801 (N_16801,N_15630,N_14342);
nor U16802 (N_16802,N_14273,N_14222);
nand U16803 (N_16803,N_15093,N_14707);
and U16804 (N_16804,N_15194,N_15259);
nand U16805 (N_16805,N_15729,N_15393);
nand U16806 (N_16806,N_15133,N_14232);
or U16807 (N_16807,N_15105,N_15601);
nor U16808 (N_16808,N_14428,N_14687);
nand U16809 (N_16809,N_14479,N_15983);
nand U16810 (N_16810,N_15131,N_14350);
and U16811 (N_16811,N_14178,N_15582);
nand U16812 (N_16812,N_15884,N_14570);
and U16813 (N_16813,N_14406,N_14914);
or U16814 (N_16814,N_15964,N_15748);
nand U16815 (N_16815,N_15429,N_15846);
nor U16816 (N_16816,N_15519,N_14036);
nor U16817 (N_16817,N_15486,N_15686);
and U16818 (N_16818,N_15102,N_14291);
xnor U16819 (N_16819,N_14314,N_15550);
nor U16820 (N_16820,N_15861,N_14098);
nand U16821 (N_16821,N_15121,N_15009);
xor U16822 (N_16822,N_14384,N_15749);
nand U16823 (N_16823,N_14398,N_15572);
nor U16824 (N_16824,N_14185,N_15407);
nand U16825 (N_16825,N_15451,N_14930);
and U16826 (N_16826,N_15489,N_15982);
nand U16827 (N_16827,N_15332,N_15161);
nor U16828 (N_16828,N_14603,N_15467);
nand U16829 (N_16829,N_14249,N_15779);
or U16830 (N_16830,N_15765,N_15417);
or U16831 (N_16831,N_15617,N_14621);
nor U16832 (N_16832,N_15715,N_15342);
nor U16833 (N_16833,N_15703,N_14748);
nor U16834 (N_16834,N_15087,N_15162);
nor U16835 (N_16835,N_15589,N_15669);
or U16836 (N_16836,N_14625,N_15039);
nand U16837 (N_16837,N_14973,N_15677);
and U16838 (N_16838,N_15739,N_15575);
nand U16839 (N_16839,N_14212,N_15287);
or U16840 (N_16840,N_15005,N_14992);
and U16841 (N_16841,N_14745,N_15038);
and U16842 (N_16842,N_14039,N_15099);
nor U16843 (N_16843,N_15482,N_14722);
nand U16844 (N_16844,N_15046,N_15966);
and U16845 (N_16845,N_14714,N_14301);
and U16846 (N_16846,N_15626,N_14154);
and U16847 (N_16847,N_14374,N_14818);
nand U16848 (N_16848,N_14441,N_14358);
or U16849 (N_16849,N_14841,N_14081);
or U16850 (N_16850,N_15277,N_14935);
or U16851 (N_16851,N_14468,N_15216);
and U16852 (N_16852,N_15909,N_15969);
nand U16853 (N_16853,N_14677,N_14694);
and U16854 (N_16854,N_14902,N_15028);
nor U16855 (N_16855,N_14581,N_14996);
or U16856 (N_16856,N_14302,N_14798);
or U16857 (N_16857,N_14310,N_14537);
nand U16858 (N_16858,N_14026,N_14129);
or U16859 (N_16859,N_14246,N_15804);
or U16860 (N_16860,N_15833,N_14897);
nor U16861 (N_16861,N_14312,N_14453);
and U16862 (N_16862,N_15917,N_14940);
or U16863 (N_16863,N_14120,N_15075);
and U16864 (N_16864,N_15289,N_15531);
nor U16865 (N_16865,N_15843,N_14242);
and U16866 (N_16866,N_15784,N_15887);
and U16867 (N_16867,N_15906,N_15069);
nand U16868 (N_16868,N_15337,N_14555);
and U16869 (N_16869,N_14820,N_14528);
nor U16870 (N_16870,N_14663,N_15597);
or U16871 (N_16871,N_15181,N_14371);
and U16872 (N_16872,N_15077,N_15891);
nand U16873 (N_16873,N_14847,N_14014);
and U16874 (N_16874,N_15436,N_15434);
or U16875 (N_16875,N_14501,N_15960);
nor U16876 (N_16876,N_15609,N_14949);
nand U16877 (N_16877,N_14942,N_15871);
nor U16878 (N_16878,N_15699,N_15491);
or U16879 (N_16879,N_15537,N_14517);
and U16880 (N_16880,N_15528,N_15718);
nor U16881 (N_16881,N_14368,N_14340);
nand U16882 (N_16882,N_15929,N_15376);
or U16883 (N_16883,N_15890,N_14928);
nor U16884 (N_16884,N_15950,N_14438);
or U16885 (N_16885,N_15490,N_14031);
nand U16886 (N_16886,N_15690,N_14179);
nor U16887 (N_16887,N_15720,N_15468);
nor U16888 (N_16888,N_15650,N_14672);
or U16889 (N_16889,N_14974,N_15848);
nand U16890 (N_16890,N_15408,N_14155);
nand U16891 (N_16891,N_15897,N_15827);
nor U16892 (N_16892,N_14808,N_14075);
and U16893 (N_16893,N_15980,N_15879);
and U16894 (N_16894,N_14960,N_14921);
nor U16895 (N_16895,N_15591,N_14958);
and U16896 (N_16896,N_14525,N_14499);
nor U16897 (N_16897,N_15740,N_15066);
nor U16898 (N_16898,N_14900,N_14792);
and U16899 (N_16899,N_15061,N_14148);
and U16900 (N_16900,N_15452,N_14980);
nand U16901 (N_16901,N_15907,N_15636);
nor U16902 (N_16902,N_14055,N_15687);
and U16903 (N_16903,N_15297,N_15955);
and U16904 (N_16904,N_15198,N_14777);
nand U16905 (N_16905,N_14281,N_15067);
nor U16906 (N_16906,N_14353,N_15516);
and U16907 (N_16907,N_14403,N_15199);
nor U16908 (N_16908,N_14334,N_14985);
xor U16909 (N_16909,N_15596,N_14456);
or U16910 (N_16910,N_15614,N_14157);
nand U16911 (N_16911,N_15670,N_15499);
and U16912 (N_16912,N_15472,N_14184);
and U16913 (N_16913,N_14931,N_15892);
and U16914 (N_16914,N_14813,N_14470);
or U16915 (N_16915,N_14292,N_14664);
nand U16916 (N_16916,N_14789,N_14089);
and U16917 (N_16917,N_15316,N_14193);
nor U16918 (N_16918,N_15645,N_14699);
or U16919 (N_16919,N_15523,N_15049);
or U16920 (N_16920,N_15930,N_15344);
nor U16921 (N_16921,N_15068,N_14686);
and U16922 (N_16922,N_15540,N_14223);
nand U16923 (N_16923,N_14116,N_15694);
nor U16924 (N_16924,N_15439,N_14950);
or U16925 (N_16925,N_14167,N_15200);
or U16926 (N_16926,N_15493,N_14024);
nor U16927 (N_16927,N_14182,N_15127);
or U16928 (N_16928,N_14719,N_15698);
and U16929 (N_16929,N_14170,N_15806);
nand U16930 (N_16930,N_14600,N_14408);
or U16931 (N_16931,N_15635,N_15395);
nor U16932 (N_16932,N_15787,N_15311);
or U16933 (N_16933,N_14171,N_15498);
nor U16934 (N_16934,N_14674,N_14964);
nand U16935 (N_16935,N_14769,N_15841);
nor U16936 (N_16936,N_15657,N_15155);
nand U16937 (N_16937,N_15512,N_15772);
and U16938 (N_16938,N_14571,N_15605);
or U16939 (N_16939,N_15723,N_14856);
or U16940 (N_16940,N_15998,N_15072);
nor U16941 (N_16941,N_14458,N_14559);
and U16942 (N_16942,N_15753,N_14230);
nor U16943 (N_16943,N_14760,N_14666);
nand U16944 (N_16944,N_14647,N_14304);
nor U16945 (N_16945,N_14241,N_14609);
and U16946 (N_16946,N_14648,N_15404);
or U16947 (N_16947,N_15904,N_15048);
nor U16948 (N_16948,N_15031,N_15147);
or U16949 (N_16949,N_14332,N_14125);
nor U16950 (N_16950,N_15278,N_15576);
nor U16951 (N_16951,N_14716,N_14873);
nand U16952 (N_16952,N_15789,N_14336);
nand U16953 (N_16953,N_15281,N_15615);
nand U16954 (N_16954,N_14825,N_15169);
and U16955 (N_16955,N_15268,N_15785);
nor U16956 (N_16956,N_15872,N_14884);
nand U16957 (N_16957,N_15639,N_14723);
nor U16958 (N_16958,N_15727,N_15037);
and U16959 (N_16959,N_15175,N_15197);
and U16960 (N_16960,N_14153,N_14685);
or U16961 (N_16961,N_14614,N_15000);
and U16962 (N_16962,N_15513,N_14562);
nand U16963 (N_16963,N_15965,N_14652);
nor U16964 (N_16964,N_15250,N_15238);
and U16965 (N_16965,N_15507,N_15750);
and U16966 (N_16966,N_14221,N_15813);
and U16967 (N_16967,N_15755,N_15508);
nand U16968 (N_16968,N_15569,N_15101);
and U16969 (N_16969,N_15823,N_14883);
and U16970 (N_16970,N_14210,N_14252);
and U16971 (N_16971,N_15430,N_15957);
or U16972 (N_16972,N_14965,N_14547);
or U16973 (N_16973,N_15258,N_15345);
nand U16974 (N_16974,N_14105,N_14947);
nand U16975 (N_16975,N_14881,N_14569);
and U16976 (N_16976,N_15177,N_15185);
nand U16977 (N_16977,N_15714,N_15021);
and U16978 (N_16978,N_14034,N_14051);
or U16979 (N_16979,N_14842,N_14817);
nand U16980 (N_16980,N_15627,N_14799);
or U16981 (N_16981,N_15330,N_14077);
or U16982 (N_16982,N_14594,N_15834);
nor U16983 (N_16983,N_14606,N_15673);
nand U16984 (N_16984,N_15312,N_15062);
nor U16985 (N_16985,N_14607,N_14174);
nand U16986 (N_16986,N_15883,N_15542);
or U16987 (N_16987,N_14139,N_14287);
or U16988 (N_16988,N_14503,N_15416);
nand U16989 (N_16989,N_14424,N_14383);
nand U16990 (N_16990,N_15083,N_14512);
and U16991 (N_16991,N_14450,N_14454);
nor U16992 (N_16992,N_15933,N_14247);
nand U16993 (N_16993,N_15880,N_15317);
nor U16994 (N_16994,N_14038,N_14107);
nand U16995 (N_16995,N_15064,N_14670);
and U16996 (N_16996,N_14524,N_15060);
or U16997 (N_16997,N_14220,N_15948);
and U16998 (N_16998,N_14476,N_15464);
or U16999 (N_16999,N_15409,N_15939);
nor U17000 (N_17000,N_14007,N_14945);
or U17001 (N_17001,N_14763,N_14320);
and U17002 (N_17002,N_14652,N_15450);
nand U17003 (N_17003,N_14132,N_14433);
nand U17004 (N_17004,N_15926,N_14756);
and U17005 (N_17005,N_14610,N_14775);
nor U17006 (N_17006,N_15305,N_14064);
or U17007 (N_17007,N_14189,N_14935);
nor U17008 (N_17008,N_14401,N_14934);
nand U17009 (N_17009,N_14777,N_15200);
nand U17010 (N_17010,N_15310,N_15918);
and U17011 (N_17011,N_15367,N_15462);
or U17012 (N_17012,N_14687,N_14336);
nand U17013 (N_17013,N_14361,N_15563);
and U17014 (N_17014,N_15771,N_14080);
and U17015 (N_17015,N_15806,N_15975);
or U17016 (N_17016,N_15097,N_14762);
nor U17017 (N_17017,N_14043,N_15742);
and U17018 (N_17018,N_15034,N_14513);
or U17019 (N_17019,N_14061,N_15151);
nand U17020 (N_17020,N_15556,N_14389);
nor U17021 (N_17021,N_15708,N_15683);
nand U17022 (N_17022,N_14190,N_14599);
nor U17023 (N_17023,N_15270,N_14455);
or U17024 (N_17024,N_14745,N_15610);
nor U17025 (N_17025,N_15975,N_14022);
nor U17026 (N_17026,N_14782,N_14776);
nand U17027 (N_17027,N_15727,N_15838);
nor U17028 (N_17028,N_14970,N_14283);
nand U17029 (N_17029,N_14000,N_14585);
and U17030 (N_17030,N_14009,N_14113);
or U17031 (N_17031,N_14173,N_15425);
nor U17032 (N_17032,N_14285,N_15478);
and U17033 (N_17033,N_15038,N_14929);
nor U17034 (N_17034,N_15083,N_15195);
and U17035 (N_17035,N_15253,N_15420);
or U17036 (N_17036,N_14670,N_15611);
or U17037 (N_17037,N_14955,N_15203);
nor U17038 (N_17038,N_15304,N_15954);
and U17039 (N_17039,N_15192,N_15147);
or U17040 (N_17040,N_14199,N_14881);
and U17041 (N_17041,N_14479,N_15191);
nand U17042 (N_17042,N_14259,N_14669);
and U17043 (N_17043,N_14565,N_14533);
or U17044 (N_17044,N_15589,N_15948);
nand U17045 (N_17045,N_14089,N_15916);
nor U17046 (N_17046,N_15408,N_14325);
and U17047 (N_17047,N_14813,N_14861);
or U17048 (N_17048,N_14658,N_15135);
or U17049 (N_17049,N_15271,N_14142);
nand U17050 (N_17050,N_15501,N_15525);
nand U17051 (N_17051,N_14951,N_14810);
nor U17052 (N_17052,N_14506,N_15009);
and U17053 (N_17053,N_15521,N_15633);
or U17054 (N_17054,N_14310,N_15149);
and U17055 (N_17055,N_14486,N_15969);
nor U17056 (N_17056,N_14279,N_15899);
or U17057 (N_17057,N_14308,N_14015);
or U17058 (N_17058,N_15805,N_15453);
and U17059 (N_17059,N_14343,N_14030);
or U17060 (N_17060,N_14118,N_14217);
or U17061 (N_17061,N_15262,N_14944);
nand U17062 (N_17062,N_14881,N_15932);
or U17063 (N_17063,N_15834,N_15524);
or U17064 (N_17064,N_14145,N_14078);
and U17065 (N_17065,N_14146,N_14420);
or U17066 (N_17066,N_14843,N_15752);
and U17067 (N_17067,N_14577,N_14721);
and U17068 (N_17068,N_15398,N_14470);
nand U17069 (N_17069,N_14627,N_15695);
or U17070 (N_17070,N_14772,N_15141);
nand U17071 (N_17071,N_15121,N_15487);
and U17072 (N_17072,N_14520,N_14077);
nand U17073 (N_17073,N_14576,N_14798);
nand U17074 (N_17074,N_14424,N_14134);
nor U17075 (N_17075,N_14724,N_14574);
and U17076 (N_17076,N_14924,N_14873);
or U17077 (N_17077,N_14150,N_14161);
and U17078 (N_17078,N_15008,N_14778);
nor U17079 (N_17079,N_14739,N_14599);
nand U17080 (N_17080,N_14573,N_14599);
nor U17081 (N_17081,N_15777,N_14667);
nor U17082 (N_17082,N_15070,N_15196);
nand U17083 (N_17083,N_14845,N_14836);
and U17084 (N_17084,N_14459,N_14010);
nor U17085 (N_17085,N_15653,N_14030);
and U17086 (N_17086,N_14238,N_14713);
or U17087 (N_17087,N_15854,N_14903);
or U17088 (N_17088,N_14423,N_14948);
or U17089 (N_17089,N_15153,N_14081);
or U17090 (N_17090,N_15406,N_14018);
or U17091 (N_17091,N_14182,N_15812);
nand U17092 (N_17092,N_15821,N_15882);
or U17093 (N_17093,N_15859,N_15753);
nor U17094 (N_17094,N_14353,N_14566);
and U17095 (N_17095,N_15230,N_15708);
nor U17096 (N_17096,N_15424,N_14466);
nand U17097 (N_17097,N_15740,N_14804);
nor U17098 (N_17098,N_15171,N_15392);
nor U17099 (N_17099,N_14543,N_15132);
nor U17100 (N_17100,N_14601,N_14094);
nand U17101 (N_17101,N_15444,N_14872);
and U17102 (N_17102,N_14153,N_15139);
nand U17103 (N_17103,N_15603,N_15659);
xnor U17104 (N_17104,N_15975,N_15953);
or U17105 (N_17105,N_15160,N_15433);
nand U17106 (N_17106,N_14087,N_14137);
nand U17107 (N_17107,N_15858,N_15662);
nor U17108 (N_17108,N_15967,N_14851);
and U17109 (N_17109,N_15133,N_15119);
nand U17110 (N_17110,N_14117,N_14151);
or U17111 (N_17111,N_15375,N_14021);
and U17112 (N_17112,N_15126,N_14177);
and U17113 (N_17113,N_14628,N_14071);
or U17114 (N_17114,N_14204,N_15307);
and U17115 (N_17115,N_15770,N_14152);
and U17116 (N_17116,N_15851,N_14989);
and U17117 (N_17117,N_15138,N_15847);
nand U17118 (N_17118,N_14203,N_15476);
and U17119 (N_17119,N_14042,N_15824);
nor U17120 (N_17120,N_14763,N_14788);
nand U17121 (N_17121,N_15751,N_15797);
nand U17122 (N_17122,N_14367,N_15590);
and U17123 (N_17123,N_15354,N_14072);
nand U17124 (N_17124,N_15576,N_14456);
and U17125 (N_17125,N_15546,N_14590);
and U17126 (N_17126,N_15752,N_15126);
nor U17127 (N_17127,N_15354,N_14791);
and U17128 (N_17128,N_14708,N_14705);
nand U17129 (N_17129,N_15483,N_14123);
nand U17130 (N_17130,N_15821,N_14564);
nor U17131 (N_17131,N_15338,N_14617);
nand U17132 (N_17132,N_15712,N_15346);
nor U17133 (N_17133,N_14280,N_14939);
nor U17134 (N_17134,N_14029,N_15950);
nand U17135 (N_17135,N_15910,N_15846);
nor U17136 (N_17136,N_14889,N_15710);
nand U17137 (N_17137,N_15931,N_14203);
nor U17138 (N_17138,N_14548,N_15860);
nand U17139 (N_17139,N_15179,N_14459);
nor U17140 (N_17140,N_14738,N_15809);
and U17141 (N_17141,N_15153,N_14938);
nor U17142 (N_17142,N_15969,N_14510);
nor U17143 (N_17143,N_14917,N_14825);
and U17144 (N_17144,N_14522,N_15502);
nand U17145 (N_17145,N_14565,N_15860);
nand U17146 (N_17146,N_15092,N_15810);
and U17147 (N_17147,N_15321,N_15194);
and U17148 (N_17148,N_14010,N_14474);
nand U17149 (N_17149,N_14744,N_15292);
nand U17150 (N_17150,N_14943,N_14015);
or U17151 (N_17151,N_15870,N_14907);
or U17152 (N_17152,N_14706,N_14514);
nor U17153 (N_17153,N_15409,N_15816);
or U17154 (N_17154,N_15805,N_15371);
and U17155 (N_17155,N_15875,N_15339);
or U17156 (N_17156,N_14032,N_14190);
and U17157 (N_17157,N_14512,N_14778);
nor U17158 (N_17158,N_14495,N_15241);
or U17159 (N_17159,N_14564,N_15586);
nor U17160 (N_17160,N_15023,N_14660);
or U17161 (N_17161,N_14919,N_14676);
or U17162 (N_17162,N_14591,N_15803);
and U17163 (N_17163,N_14117,N_15495);
xor U17164 (N_17164,N_15903,N_14121);
nor U17165 (N_17165,N_15757,N_15330);
or U17166 (N_17166,N_15035,N_14826);
nand U17167 (N_17167,N_15495,N_14613);
nand U17168 (N_17168,N_15058,N_14556);
nand U17169 (N_17169,N_15562,N_15323);
nand U17170 (N_17170,N_15660,N_14699);
and U17171 (N_17171,N_15719,N_15927);
nand U17172 (N_17172,N_14405,N_15339);
nand U17173 (N_17173,N_15916,N_15255);
and U17174 (N_17174,N_14687,N_15348);
nor U17175 (N_17175,N_15512,N_14999);
and U17176 (N_17176,N_14869,N_15995);
or U17177 (N_17177,N_15199,N_14087);
nand U17178 (N_17178,N_15025,N_14928);
nand U17179 (N_17179,N_15275,N_15196);
nand U17180 (N_17180,N_15464,N_15020);
xnor U17181 (N_17181,N_14514,N_15925);
nand U17182 (N_17182,N_15200,N_14589);
or U17183 (N_17183,N_15186,N_15399);
nor U17184 (N_17184,N_14880,N_14991);
nand U17185 (N_17185,N_15058,N_15879);
nor U17186 (N_17186,N_14003,N_15264);
nand U17187 (N_17187,N_14716,N_14988);
nand U17188 (N_17188,N_14567,N_14834);
and U17189 (N_17189,N_14117,N_15927);
or U17190 (N_17190,N_15942,N_14935);
and U17191 (N_17191,N_14881,N_15791);
nor U17192 (N_17192,N_14280,N_14630);
nor U17193 (N_17193,N_14104,N_14040);
nand U17194 (N_17194,N_15922,N_14963);
or U17195 (N_17195,N_15282,N_15583);
nand U17196 (N_17196,N_15275,N_15922);
nand U17197 (N_17197,N_14085,N_14250);
nand U17198 (N_17198,N_15278,N_14449);
or U17199 (N_17199,N_15287,N_15520);
or U17200 (N_17200,N_14450,N_14845);
or U17201 (N_17201,N_15516,N_15519);
nand U17202 (N_17202,N_14889,N_15622);
or U17203 (N_17203,N_15337,N_14222);
or U17204 (N_17204,N_15587,N_14149);
nor U17205 (N_17205,N_15416,N_14352);
nor U17206 (N_17206,N_15533,N_14822);
nor U17207 (N_17207,N_15286,N_14958);
nor U17208 (N_17208,N_15958,N_14332);
nor U17209 (N_17209,N_15238,N_14699);
and U17210 (N_17210,N_14505,N_15079);
or U17211 (N_17211,N_14766,N_14337);
nand U17212 (N_17212,N_14628,N_14515);
nand U17213 (N_17213,N_14882,N_15846);
nand U17214 (N_17214,N_15294,N_14948);
nor U17215 (N_17215,N_15433,N_15822);
and U17216 (N_17216,N_14960,N_15755);
and U17217 (N_17217,N_14561,N_14668);
or U17218 (N_17218,N_15068,N_15930);
nor U17219 (N_17219,N_14885,N_14678);
nand U17220 (N_17220,N_14778,N_15230);
or U17221 (N_17221,N_14963,N_15192);
nor U17222 (N_17222,N_15513,N_15464);
or U17223 (N_17223,N_14818,N_14558);
and U17224 (N_17224,N_14581,N_14337);
or U17225 (N_17225,N_15869,N_15290);
nand U17226 (N_17226,N_14532,N_14697);
and U17227 (N_17227,N_14672,N_15844);
nand U17228 (N_17228,N_15124,N_15694);
nand U17229 (N_17229,N_14664,N_15752);
nor U17230 (N_17230,N_14542,N_15996);
nand U17231 (N_17231,N_15659,N_14436);
nand U17232 (N_17232,N_15344,N_14236);
and U17233 (N_17233,N_14146,N_14598);
or U17234 (N_17234,N_14377,N_15354);
and U17235 (N_17235,N_15489,N_14294);
nor U17236 (N_17236,N_14205,N_15837);
and U17237 (N_17237,N_14306,N_15184);
or U17238 (N_17238,N_15346,N_14491);
or U17239 (N_17239,N_14118,N_15102);
or U17240 (N_17240,N_14774,N_14662);
or U17241 (N_17241,N_15132,N_14240);
nand U17242 (N_17242,N_14947,N_14682);
or U17243 (N_17243,N_15613,N_15957);
nor U17244 (N_17244,N_15814,N_15443);
nor U17245 (N_17245,N_15242,N_15717);
nand U17246 (N_17246,N_15776,N_15993);
and U17247 (N_17247,N_14129,N_14504);
nor U17248 (N_17248,N_15376,N_14734);
nand U17249 (N_17249,N_14614,N_15260);
or U17250 (N_17250,N_15320,N_15286);
nand U17251 (N_17251,N_15080,N_15604);
nand U17252 (N_17252,N_14854,N_15603);
and U17253 (N_17253,N_15186,N_14707);
nand U17254 (N_17254,N_15716,N_15143);
and U17255 (N_17255,N_15156,N_15352);
and U17256 (N_17256,N_14874,N_14877);
nand U17257 (N_17257,N_14364,N_14785);
nor U17258 (N_17258,N_14994,N_15423);
and U17259 (N_17259,N_14235,N_14953);
and U17260 (N_17260,N_15920,N_14297);
or U17261 (N_17261,N_14869,N_15425);
and U17262 (N_17262,N_15037,N_15497);
nand U17263 (N_17263,N_15205,N_14121);
or U17264 (N_17264,N_14772,N_14478);
nand U17265 (N_17265,N_15367,N_14033);
nor U17266 (N_17266,N_15456,N_14204);
nor U17267 (N_17267,N_14870,N_14686);
nor U17268 (N_17268,N_14968,N_15831);
and U17269 (N_17269,N_14659,N_15508);
nand U17270 (N_17270,N_14074,N_14833);
nor U17271 (N_17271,N_15399,N_14618);
or U17272 (N_17272,N_15788,N_15752);
or U17273 (N_17273,N_14459,N_15985);
nor U17274 (N_17274,N_14179,N_14772);
nand U17275 (N_17275,N_14295,N_14071);
or U17276 (N_17276,N_15261,N_14108);
or U17277 (N_17277,N_15058,N_14069);
nand U17278 (N_17278,N_15126,N_14375);
or U17279 (N_17279,N_14392,N_15875);
or U17280 (N_17280,N_15230,N_15254);
nand U17281 (N_17281,N_15532,N_14325);
xor U17282 (N_17282,N_14964,N_14769);
nand U17283 (N_17283,N_14821,N_14612);
nor U17284 (N_17284,N_15543,N_15685);
nor U17285 (N_17285,N_14226,N_15573);
and U17286 (N_17286,N_14771,N_15212);
or U17287 (N_17287,N_14125,N_15714);
nand U17288 (N_17288,N_14886,N_15447);
or U17289 (N_17289,N_15098,N_15265);
nand U17290 (N_17290,N_15095,N_14348);
nor U17291 (N_17291,N_14521,N_15812);
or U17292 (N_17292,N_15051,N_15518);
nand U17293 (N_17293,N_14425,N_15281);
nor U17294 (N_17294,N_15440,N_14447);
nand U17295 (N_17295,N_14420,N_14951);
nor U17296 (N_17296,N_14093,N_14603);
xnor U17297 (N_17297,N_15442,N_15009);
nand U17298 (N_17298,N_15271,N_14798);
or U17299 (N_17299,N_15446,N_15731);
nand U17300 (N_17300,N_15912,N_15607);
or U17301 (N_17301,N_14249,N_15918);
or U17302 (N_17302,N_15390,N_15197);
or U17303 (N_17303,N_15452,N_14193);
xnor U17304 (N_17304,N_15541,N_14142);
or U17305 (N_17305,N_14795,N_14187);
or U17306 (N_17306,N_15744,N_15999);
nand U17307 (N_17307,N_14533,N_15643);
nand U17308 (N_17308,N_15955,N_14284);
nor U17309 (N_17309,N_14430,N_14802);
and U17310 (N_17310,N_15817,N_15757);
nand U17311 (N_17311,N_14092,N_14647);
nand U17312 (N_17312,N_14807,N_14686);
and U17313 (N_17313,N_15018,N_15675);
nand U17314 (N_17314,N_15529,N_14294);
and U17315 (N_17315,N_14749,N_15263);
or U17316 (N_17316,N_15510,N_15595);
or U17317 (N_17317,N_15970,N_15921);
nand U17318 (N_17318,N_15508,N_14809);
or U17319 (N_17319,N_15269,N_15971);
nor U17320 (N_17320,N_15544,N_15445);
nor U17321 (N_17321,N_15600,N_14412);
and U17322 (N_17322,N_15003,N_14067);
nand U17323 (N_17323,N_14496,N_14642);
and U17324 (N_17324,N_15270,N_14382);
nand U17325 (N_17325,N_14643,N_14085);
or U17326 (N_17326,N_15821,N_15735);
nand U17327 (N_17327,N_14498,N_14543);
and U17328 (N_17328,N_15781,N_15196);
or U17329 (N_17329,N_15467,N_14094);
nor U17330 (N_17330,N_14125,N_14249);
and U17331 (N_17331,N_15549,N_15300);
nor U17332 (N_17332,N_15618,N_14342);
and U17333 (N_17333,N_15532,N_15568);
or U17334 (N_17334,N_14017,N_15203);
nand U17335 (N_17335,N_15347,N_14491);
nor U17336 (N_17336,N_14597,N_15814);
or U17337 (N_17337,N_14077,N_15897);
or U17338 (N_17338,N_15715,N_14784);
nand U17339 (N_17339,N_14857,N_14049);
nor U17340 (N_17340,N_14703,N_15123);
and U17341 (N_17341,N_14290,N_14631);
and U17342 (N_17342,N_14895,N_15920);
or U17343 (N_17343,N_15955,N_14520);
and U17344 (N_17344,N_15712,N_14127);
or U17345 (N_17345,N_14902,N_15390);
nand U17346 (N_17346,N_14778,N_15491);
nand U17347 (N_17347,N_15273,N_15149);
nand U17348 (N_17348,N_14291,N_14695);
nor U17349 (N_17349,N_14129,N_14477);
and U17350 (N_17350,N_15811,N_15750);
or U17351 (N_17351,N_14019,N_14377);
nor U17352 (N_17352,N_15212,N_15732);
nand U17353 (N_17353,N_14584,N_15311);
nor U17354 (N_17354,N_15429,N_15369);
and U17355 (N_17355,N_15940,N_14000);
nor U17356 (N_17356,N_15945,N_15573);
or U17357 (N_17357,N_14324,N_14216);
and U17358 (N_17358,N_14500,N_15203);
or U17359 (N_17359,N_15786,N_15660);
or U17360 (N_17360,N_15076,N_14453);
nor U17361 (N_17361,N_14617,N_15620);
nand U17362 (N_17362,N_14235,N_14296);
and U17363 (N_17363,N_14940,N_15790);
or U17364 (N_17364,N_14424,N_15461);
nand U17365 (N_17365,N_14568,N_14309);
or U17366 (N_17366,N_14114,N_15987);
nor U17367 (N_17367,N_14437,N_14400);
nand U17368 (N_17368,N_14608,N_14112);
and U17369 (N_17369,N_15896,N_14056);
nor U17370 (N_17370,N_15840,N_14180);
or U17371 (N_17371,N_14409,N_15301);
and U17372 (N_17372,N_14476,N_15166);
and U17373 (N_17373,N_15118,N_14704);
nand U17374 (N_17374,N_15146,N_15287);
nand U17375 (N_17375,N_14786,N_15077);
or U17376 (N_17376,N_15474,N_14164);
and U17377 (N_17377,N_15784,N_14298);
nand U17378 (N_17378,N_14082,N_14461);
or U17379 (N_17379,N_15611,N_14341);
nor U17380 (N_17380,N_14085,N_14906);
nand U17381 (N_17381,N_15258,N_15188);
and U17382 (N_17382,N_15132,N_15270);
nor U17383 (N_17383,N_15273,N_14034);
and U17384 (N_17384,N_15516,N_15959);
nor U17385 (N_17385,N_14738,N_14031);
nor U17386 (N_17386,N_15885,N_15441);
or U17387 (N_17387,N_15929,N_14514);
and U17388 (N_17388,N_15747,N_14082);
and U17389 (N_17389,N_15303,N_15198);
nor U17390 (N_17390,N_14556,N_15404);
or U17391 (N_17391,N_15235,N_15266);
or U17392 (N_17392,N_14176,N_14018);
nor U17393 (N_17393,N_14124,N_15145);
or U17394 (N_17394,N_15048,N_14221);
nor U17395 (N_17395,N_14821,N_14594);
nor U17396 (N_17396,N_14244,N_15433);
and U17397 (N_17397,N_15504,N_15795);
and U17398 (N_17398,N_15731,N_15333);
nor U17399 (N_17399,N_14252,N_15370);
nand U17400 (N_17400,N_14991,N_15370);
nand U17401 (N_17401,N_14609,N_14924);
or U17402 (N_17402,N_14713,N_14706);
or U17403 (N_17403,N_15266,N_14000);
or U17404 (N_17404,N_15326,N_15694);
and U17405 (N_17405,N_14339,N_14965);
and U17406 (N_17406,N_14631,N_15321);
nor U17407 (N_17407,N_15558,N_14528);
nand U17408 (N_17408,N_14095,N_15399);
or U17409 (N_17409,N_14244,N_14532);
nand U17410 (N_17410,N_14331,N_14879);
nor U17411 (N_17411,N_15630,N_14169);
or U17412 (N_17412,N_15750,N_15852);
xor U17413 (N_17413,N_15139,N_15822);
nand U17414 (N_17414,N_15780,N_15343);
nor U17415 (N_17415,N_14240,N_14859);
nor U17416 (N_17416,N_15110,N_14079);
nor U17417 (N_17417,N_15252,N_15788);
and U17418 (N_17418,N_14372,N_14466);
or U17419 (N_17419,N_14337,N_14482);
or U17420 (N_17420,N_14912,N_14717);
xnor U17421 (N_17421,N_14215,N_15920);
and U17422 (N_17422,N_14382,N_14021);
or U17423 (N_17423,N_15321,N_14953);
nor U17424 (N_17424,N_15714,N_15166);
nor U17425 (N_17425,N_15871,N_15829);
or U17426 (N_17426,N_14502,N_14282);
or U17427 (N_17427,N_14489,N_14303);
or U17428 (N_17428,N_14225,N_15580);
nor U17429 (N_17429,N_15021,N_14236);
nor U17430 (N_17430,N_14889,N_14337);
nor U17431 (N_17431,N_15230,N_15380);
nor U17432 (N_17432,N_15932,N_14239);
and U17433 (N_17433,N_15487,N_15100);
nand U17434 (N_17434,N_15652,N_14426);
nor U17435 (N_17435,N_14735,N_14369);
nor U17436 (N_17436,N_15297,N_14397);
nand U17437 (N_17437,N_15176,N_14573);
nand U17438 (N_17438,N_15685,N_14164);
nor U17439 (N_17439,N_15857,N_15352);
or U17440 (N_17440,N_15344,N_15434);
nand U17441 (N_17441,N_14042,N_15403);
or U17442 (N_17442,N_15377,N_14342);
and U17443 (N_17443,N_15627,N_15886);
nor U17444 (N_17444,N_14516,N_14274);
nor U17445 (N_17445,N_15032,N_14371);
nor U17446 (N_17446,N_14495,N_15914);
and U17447 (N_17447,N_14697,N_14363);
and U17448 (N_17448,N_15390,N_14472);
or U17449 (N_17449,N_14874,N_15886);
and U17450 (N_17450,N_14708,N_14481);
nor U17451 (N_17451,N_14178,N_15853);
or U17452 (N_17452,N_14164,N_14339);
and U17453 (N_17453,N_14474,N_15469);
or U17454 (N_17454,N_14589,N_15077);
nor U17455 (N_17455,N_15513,N_14355);
nand U17456 (N_17456,N_15936,N_14552);
nor U17457 (N_17457,N_15022,N_14996);
nor U17458 (N_17458,N_15633,N_14920);
and U17459 (N_17459,N_14884,N_15923);
nand U17460 (N_17460,N_14720,N_15170);
xor U17461 (N_17461,N_14034,N_14020);
and U17462 (N_17462,N_14537,N_14976);
nor U17463 (N_17463,N_15772,N_15353);
and U17464 (N_17464,N_15852,N_14573);
nand U17465 (N_17465,N_14662,N_15273);
nor U17466 (N_17466,N_14979,N_15452);
nor U17467 (N_17467,N_14582,N_15383);
nand U17468 (N_17468,N_14569,N_15106);
xnor U17469 (N_17469,N_15291,N_15719);
nor U17470 (N_17470,N_14087,N_14623);
or U17471 (N_17471,N_14768,N_14740);
or U17472 (N_17472,N_14214,N_15846);
nand U17473 (N_17473,N_15532,N_15004);
nand U17474 (N_17474,N_14444,N_15627);
or U17475 (N_17475,N_14265,N_15406);
nor U17476 (N_17476,N_15972,N_14201);
or U17477 (N_17477,N_15334,N_14478);
and U17478 (N_17478,N_15391,N_14631);
nor U17479 (N_17479,N_15304,N_15953);
nand U17480 (N_17480,N_14119,N_15355);
nand U17481 (N_17481,N_15255,N_15229);
or U17482 (N_17482,N_14657,N_14202);
and U17483 (N_17483,N_15262,N_14598);
nand U17484 (N_17484,N_14422,N_14355);
nand U17485 (N_17485,N_15965,N_15057);
nand U17486 (N_17486,N_14013,N_15945);
and U17487 (N_17487,N_14699,N_15658);
and U17488 (N_17488,N_14369,N_14783);
or U17489 (N_17489,N_14780,N_15678);
or U17490 (N_17490,N_14323,N_14034);
nand U17491 (N_17491,N_15311,N_15185);
and U17492 (N_17492,N_14190,N_15901);
nand U17493 (N_17493,N_15872,N_15059);
nand U17494 (N_17494,N_15136,N_14633);
or U17495 (N_17495,N_14177,N_15945);
or U17496 (N_17496,N_15355,N_15095);
or U17497 (N_17497,N_14709,N_15490);
nand U17498 (N_17498,N_15758,N_15505);
or U17499 (N_17499,N_14781,N_15662);
or U17500 (N_17500,N_15130,N_14559);
nor U17501 (N_17501,N_15315,N_14329);
nor U17502 (N_17502,N_15636,N_15876);
or U17503 (N_17503,N_14061,N_14538);
nand U17504 (N_17504,N_15301,N_15754);
nand U17505 (N_17505,N_14474,N_14319);
nor U17506 (N_17506,N_15416,N_15868);
nand U17507 (N_17507,N_15920,N_14379);
nand U17508 (N_17508,N_15455,N_14117);
and U17509 (N_17509,N_15871,N_14197);
nand U17510 (N_17510,N_14443,N_15209);
nor U17511 (N_17511,N_15819,N_14038);
nand U17512 (N_17512,N_15339,N_14934);
or U17513 (N_17513,N_15348,N_14945);
and U17514 (N_17514,N_14422,N_14223);
or U17515 (N_17515,N_14390,N_14789);
and U17516 (N_17516,N_15703,N_15055);
nor U17517 (N_17517,N_15064,N_15094);
nor U17518 (N_17518,N_15085,N_14306);
or U17519 (N_17519,N_15584,N_15618);
or U17520 (N_17520,N_15122,N_14452);
nor U17521 (N_17521,N_14912,N_14480);
nand U17522 (N_17522,N_15078,N_14754);
or U17523 (N_17523,N_15812,N_15278);
or U17524 (N_17524,N_14105,N_14520);
and U17525 (N_17525,N_15042,N_15783);
nand U17526 (N_17526,N_15264,N_14371);
and U17527 (N_17527,N_14512,N_15637);
nand U17528 (N_17528,N_14015,N_15786);
nand U17529 (N_17529,N_14278,N_15163);
or U17530 (N_17530,N_15692,N_15446);
or U17531 (N_17531,N_14933,N_14280);
or U17532 (N_17532,N_15708,N_15651);
nor U17533 (N_17533,N_14360,N_15850);
or U17534 (N_17534,N_14014,N_15793);
nand U17535 (N_17535,N_15754,N_15007);
and U17536 (N_17536,N_14007,N_14220);
and U17537 (N_17537,N_15270,N_14786);
or U17538 (N_17538,N_15254,N_14633);
nand U17539 (N_17539,N_15981,N_15815);
or U17540 (N_17540,N_15929,N_14763);
nor U17541 (N_17541,N_15168,N_14720);
nor U17542 (N_17542,N_14759,N_15627);
and U17543 (N_17543,N_15587,N_14050);
and U17544 (N_17544,N_14108,N_14786);
and U17545 (N_17545,N_14874,N_14835);
or U17546 (N_17546,N_14956,N_15404);
or U17547 (N_17547,N_15144,N_14542);
and U17548 (N_17548,N_15661,N_15718);
and U17549 (N_17549,N_14188,N_14705);
and U17550 (N_17550,N_14203,N_14966);
nor U17551 (N_17551,N_14557,N_14452);
or U17552 (N_17552,N_14709,N_15477);
or U17553 (N_17553,N_14729,N_14295);
or U17554 (N_17554,N_15150,N_15469);
nand U17555 (N_17555,N_15550,N_14599);
and U17556 (N_17556,N_14842,N_15657);
nor U17557 (N_17557,N_14348,N_14982);
nand U17558 (N_17558,N_15458,N_15632);
nor U17559 (N_17559,N_15957,N_15130);
and U17560 (N_17560,N_14025,N_14653);
nor U17561 (N_17561,N_15278,N_14626);
nor U17562 (N_17562,N_15489,N_14611);
or U17563 (N_17563,N_14356,N_15679);
nand U17564 (N_17564,N_14821,N_14582);
or U17565 (N_17565,N_14198,N_15142);
or U17566 (N_17566,N_15140,N_15354);
nand U17567 (N_17567,N_14522,N_14865);
and U17568 (N_17568,N_15949,N_14405);
and U17569 (N_17569,N_15119,N_14310);
and U17570 (N_17570,N_15571,N_15382);
nand U17571 (N_17571,N_15947,N_15971);
and U17572 (N_17572,N_15114,N_14545);
or U17573 (N_17573,N_15080,N_15989);
or U17574 (N_17574,N_14681,N_15600);
nand U17575 (N_17575,N_14864,N_14450);
or U17576 (N_17576,N_14193,N_14119);
or U17577 (N_17577,N_15445,N_14953);
or U17578 (N_17578,N_15795,N_15810);
or U17579 (N_17579,N_14828,N_15368);
and U17580 (N_17580,N_15277,N_15979);
nand U17581 (N_17581,N_14274,N_15639);
or U17582 (N_17582,N_14772,N_15424);
nand U17583 (N_17583,N_14744,N_14554);
and U17584 (N_17584,N_14127,N_15134);
and U17585 (N_17585,N_15983,N_15614);
and U17586 (N_17586,N_14517,N_15630);
nor U17587 (N_17587,N_14771,N_15467);
and U17588 (N_17588,N_15205,N_15633);
nor U17589 (N_17589,N_14999,N_14877);
and U17590 (N_17590,N_15531,N_14450);
nand U17591 (N_17591,N_14699,N_15427);
xnor U17592 (N_17592,N_14849,N_14915);
nand U17593 (N_17593,N_14944,N_15452);
or U17594 (N_17594,N_14399,N_14649);
or U17595 (N_17595,N_15881,N_14356);
nand U17596 (N_17596,N_14979,N_15022);
and U17597 (N_17597,N_14458,N_15077);
or U17598 (N_17598,N_14233,N_15219);
or U17599 (N_17599,N_14855,N_14566);
nor U17600 (N_17600,N_15357,N_15488);
nor U17601 (N_17601,N_14901,N_15564);
and U17602 (N_17602,N_15382,N_15835);
nand U17603 (N_17603,N_15559,N_15264);
nor U17604 (N_17604,N_14099,N_14952);
and U17605 (N_17605,N_15354,N_15422);
and U17606 (N_17606,N_14862,N_14793);
nor U17607 (N_17607,N_14307,N_15393);
nor U17608 (N_17608,N_15752,N_15515);
and U17609 (N_17609,N_14830,N_14087);
and U17610 (N_17610,N_14785,N_14555);
or U17611 (N_17611,N_15832,N_15386);
or U17612 (N_17612,N_15986,N_14885);
nor U17613 (N_17613,N_15377,N_14049);
or U17614 (N_17614,N_15384,N_15393);
nand U17615 (N_17615,N_15013,N_15960);
nand U17616 (N_17616,N_14993,N_15823);
or U17617 (N_17617,N_14536,N_15463);
nor U17618 (N_17618,N_14105,N_15383);
or U17619 (N_17619,N_14683,N_15060);
and U17620 (N_17620,N_15509,N_14507);
nand U17621 (N_17621,N_14048,N_15225);
and U17622 (N_17622,N_15049,N_15409);
and U17623 (N_17623,N_14976,N_15272);
xor U17624 (N_17624,N_15097,N_15469);
and U17625 (N_17625,N_14845,N_14585);
or U17626 (N_17626,N_15956,N_15780);
nor U17627 (N_17627,N_14897,N_15380);
nand U17628 (N_17628,N_14213,N_14376);
nor U17629 (N_17629,N_14876,N_15738);
and U17630 (N_17630,N_15240,N_14267);
nand U17631 (N_17631,N_15899,N_14413);
and U17632 (N_17632,N_15424,N_14603);
and U17633 (N_17633,N_14206,N_15672);
nor U17634 (N_17634,N_14896,N_14532);
nand U17635 (N_17635,N_15366,N_15536);
nand U17636 (N_17636,N_15530,N_14728);
and U17637 (N_17637,N_15988,N_15906);
nor U17638 (N_17638,N_14339,N_15075);
xor U17639 (N_17639,N_14133,N_15852);
nor U17640 (N_17640,N_15930,N_14471);
or U17641 (N_17641,N_14797,N_15504);
nor U17642 (N_17642,N_15480,N_15750);
and U17643 (N_17643,N_15630,N_15016);
and U17644 (N_17644,N_14176,N_14489);
or U17645 (N_17645,N_14613,N_15419);
and U17646 (N_17646,N_15181,N_14259);
nor U17647 (N_17647,N_14311,N_15972);
and U17648 (N_17648,N_15713,N_14003);
and U17649 (N_17649,N_15899,N_15843);
or U17650 (N_17650,N_15322,N_14905);
and U17651 (N_17651,N_15995,N_15778);
nor U17652 (N_17652,N_14110,N_14663);
or U17653 (N_17653,N_14938,N_15590);
nor U17654 (N_17654,N_14855,N_14724);
or U17655 (N_17655,N_14951,N_14945);
or U17656 (N_17656,N_15230,N_14377);
or U17657 (N_17657,N_14355,N_15210);
nor U17658 (N_17658,N_14660,N_15271);
nand U17659 (N_17659,N_14898,N_14170);
nor U17660 (N_17660,N_15981,N_14964);
nand U17661 (N_17661,N_15957,N_15050);
and U17662 (N_17662,N_15410,N_15332);
and U17663 (N_17663,N_14754,N_15478);
or U17664 (N_17664,N_15355,N_15755);
nor U17665 (N_17665,N_14367,N_15301);
or U17666 (N_17666,N_15709,N_14211);
or U17667 (N_17667,N_15233,N_14656);
xor U17668 (N_17668,N_14235,N_14067);
or U17669 (N_17669,N_14826,N_14130);
and U17670 (N_17670,N_14692,N_15234);
and U17671 (N_17671,N_15255,N_15656);
and U17672 (N_17672,N_15847,N_15975);
and U17673 (N_17673,N_14231,N_14128);
nand U17674 (N_17674,N_14638,N_14371);
nand U17675 (N_17675,N_14699,N_14835);
or U17676 (N_17676,N_14533,N_14858);
and U17677 (N_17677,N_14916,N_14472);
nor U17678 (N_17678,N_15065,N_15643);
nand U17679 (N_17679,N_14960,N_14530);
nor U17680 (N_17680,N_15617,N_15131);
or U17681 (N_17681,N_15051,N_14187);
and U17682 (N_17682,N_14036,N_14619);
and U17683 (N_17683,N_14735,N_15542);
nor U17684 (N_17684,N_14324,N_15353);
or U17685 (N_17685,N_15543,N_14407);
and U17686 (N_17686,N_14153,N_15672);
or U17687 (N_17687,N_14031,N_14646);
nand U17688 (N_17688,N_14672,N_14792);
nand U17689 (N_17689,N_14570,N_14922);
or U17690 (N_17690,N_14814,N_15175);
nor U17691 (N_17691,N_14229,N_14858);
and U17692 (N_17692,N_15960,N_15813);
and U17693 (N_17693,N_15963,N_14542);
and U17694 (N_17694,N_15684,N_15097);
nand U17695 (N_17695,N_14138,N_14761);
nand U17696 (N_17696,N_15991,N_14556);
nor U17697 (N_17697,N_14666,N_14549);
and U17698 (N_17698,N_14546,N_15183);
and U17699 (N_17699,N_15964,N_14301);
nor U17700 (N_17700,N_14734,N_14050);
or U17701 (N_17701,N_15086,N_15030);
nand U17702 (N_17702,N_15551,N_14265);
and U17703 (N_17703,N_15614,N_14771);
nor U17704 (N_17704,N_14017,N_15094);
and U17705 (N_17705,N_14021,N_15854);
and U17706 (N_17706,N_15415,N_14879);
and U17707 (N_17707,N_15332,N_15507);
and U17708 (N_17708,N_14128,N_15843);
and U17709 (N_17709,N_15842,N_15064);
and U17710 (N_17710,N_14545,N_14306);
nor U17711 (N_17711,N_15965,N_15138);
nand U17712 (N_17712,N_14748,N_14335);
nand U17713 (N_17713,N_14520,N_15853);
or U17714 (N_17714,N_14797,N_14259);
nand U17715 (N_17715,N_15281,N_14128);
or U17716 (N_17716,N_14818,N_15519);
or U17717 (N_17717,N_15428,N_14630);
nand U17718 (N_17718,N_15321,N_14869);
and U17719 (N_17719,N_15595,N_14865);
or U17720 (N_17720,N_15327,N_15179);
and U17721 (N_17721,N_15217,N_15177);
or U17722 (N_17722,N_14783,N_15342);
and U17723 (N_17723,N_15321,N_15709);
and U17724 (N_17724,N_14435,N_14355);
or U17725 (N_17725,N_15980,N_15869);
or U17726 (N_17726,N_14665,N_14949);
and U17727 (N_17727,N_15188,N_15358);
nand U17728 (N_17728,N_15784,N_15745);
or U17729 (N_17729,N_15028,N_14676);
and U17730 (N_17730,N_15716,N_14579);
nand U17731 (N_17731,N_14342,N_14804);
nor U17732 (N_17732,N_14382,N_14006);
nor U17733 (N_17733,N_14023,N_14379);
and U17734 (N_17734,N_14371,N_15564);
and U17735 (N_17735,N_15957,N_15330);
and U17736 (N_17736,N_15731,N_14758);
nor U17737 (N_17737,N_14230,N_14403);
nand U17738 (N_17738,N_15096,N_15396);
and U17739 (N_17739,N_15297,N_14097);
or U17740 (N_17740,N_14796,N_14807);
nor U17741 (N_17741,N_14872,N_14970);
and U17742 (N_17742,N_15179,N_14366);
or U17743 (N_17743,N_15895,N_15144);
and U17744 (N_17744,N_15205,N_15350);
or U17745 (N_17745,N_14724,N_15441);
nor U17746 (N_17746,N_15629,N_15715);
nand U17747 (N_17747,N_15286,N_15625);
nor U17748 (N_17748,N_15728,N_14728);
and U17749 (N_17749,N_15362,N_15508);
nand U17750 (N_17750,N_15065,N_15409);
nand U17751 (N_17751,N_15689,N_14178);
and U17752 (N_17752,N_15180,N_14275);
nand U17753 (N_17753,N_14399,N_14311);
or U17754 (N_17754,N_14932,N_14960);
nand U17755 (N_17755,N_14688,N_14158);
and U17756 (N_17756,N_14471,N_14975);
nor U17757 (N_17757,N_14912,N_15328);
or U17758 (N_17758,N_15284,N_14751);
nand U17759 (N_17759,N_14462,N_15959);
nor U17760 (N_17760,N_14494,N_14214);
or U17761 (N_17761,N_14470,N_14092);
nand U17762 (N_17762,N_14814,N_14266);
nor U17763 (N_17763,N_15274,N_14139);
and U17764 (N_17764,N_14497,N_15980);
nand U17765 (N_17765,N_15777,N_14613);
nand U17766 (N_17766,N_15931,N_15960);
and U17767 (N_17767,N_15722,N_15363);
nand U17768 (N_17768,N_14245,N_14446);
and U17769 (N_17769,N_15453,N_14520);
or U17770 (N_17770,N_15239,N_15919);
and U17771 (N_17771,N_14913,N_15830);
nand U17772 (N_17772,N_15727,N_14496);
or U17773 (N_17773,N_14129,N_15546);
nand U17774 (N_17774,N_15083,N_14184);
nand U17775 (N_17775,N_15823,N_15032);
nand U17776 (N_17776,N_14902,N_14935);
and U17777 (N_17777,N_15329,N_14322);
nand U17778 (N_17778,N_14662,N_14783);
and U17779 (N_17779,N_15852,N_14515);
or U17780 (N_17780,N_14725,N_15855);
nand U17781 (N_17781,N_15151,N_14163);
or U17782 (N_17782,N_15283,N_14399);
and U17783 (N_17783,N_15543,N_14920);
nor U17784 (N_17784,N_14181,N_15673);
nand U17785 (N_17785,N_14489,N_14869);
and U17786 (N_17786,N_14447,N_14819);
nand U17787 (N_17787,N_15305,N_15403);
nor U17788 (N_17788,N_15881,N_15688);
and U17789 (N_17789,N_14565,N_15406);
and U17790 (N_17790,N_14362,N_14804);
nand U17791 (N_17791,N_15281,N_15502);
nor U17792 (N_17792,N_15613,N_15107);
nand U17793 (N_17793,N_15745,N_14866);
nand U17794 (N_17794,N_14155,N_14944);
or U17795 (N_17795,N_15109,N_15016);
and U17796 (N_17796,N_15545,N_14961);
and U17797 (N_17797,N_14972,N_14745);
or U17798 (N_17798,N_15471,N_14499);
or U17799 (N_17799,N_14520,N_14675);
or U17800 (N_17800,N_14133,N_15456);
and U17801 (N_17801,N_15430,N_15461);
nor U17802 (N_17802,N_14259,N_15244);
and U17803 (N_17803,N_15743,N_15980);
or U17804 (N_17804,N_15961,N_14377);
and U17805 (N_17805,N_14855,N_15050);
or U17806 (N_17806,N_15308,N_15783);
nor U17807 (N_17807,N_15221,N_15540);
nor U17808 (N_17808,N_14126,N_15068);
nor U17809 (N_17809,N_15498,N_14562);
or U17810 (N_17810,N_15662,N_14405);
nor U17811 (N_17811,N_15377,N_15114);
or U17812 (N_17812,N_14028,N_14889);
nor U17813 (N_17813,N_14618,N_15596);
nand U17814 (N_17814,N_15858,N_14631);
and U17815 (N_17815,N_14059,N_15475);
and U17816 (N_17816,N_15298,N_15572);
nor U17817 (N_17817,N_14591,N_14421);
nand U17818 (N_17818,N_14655,N_14105);
nor U17819 (N_17819,N_14627,N_15917);
nand U17820 (N_17820,N_15715,N_15339);
or U17821 (N_17821,N_14040,N_14218);
nand U17822 (N_17822,N_15109,N_14432);
nor U17823 (N_17823,N_14929,N_15911);
nand U17824 (N_17824,N_14244,N_15477);
and U17825 (N_17825,N_15261,N_14648);
nor U17826 (N_17826,N_15894,N_14580);
or U17827 (N_17827,N_15112,N_14092);
and U17828 (N_17828,N_14389,N_15530);
nand U17829 (N_17829,N_15353,N_15069);
nor U17830 (N_17830,N_15768,N_14572);
nand U17831 (N_17831,N_15524,N_15418);
or U17832 (N_17832,N_14521,N_15221);
and U17833 (N_17833,N_15964,N_15402);
nor U17834 (N_17834,N_14615,N_15760);
or U17835 (N_17835,N_14749,N_15184);
nor U17836 (N_17836,N_14258,N_15294);
and U17837 (N_17837,N_15078,N_14795);
and U17838 (N_17838,N_14117,N_15152);
nor U17839 (N_17839,N_15394,N_14629);
nor U17840 (N_17840,N_14520,N_14946);
nor U17841 (N_17841,N_15151,N_14663);
and U17842 (N_17842,N_15883,N_14751);
nand U17843 (N_17843,N_15799,N_14209);
and U17844 (N_17844,N_14600,N_15439);
or U17845 (N_17845,N_14585,N_14948);
nand U17846 (N_17846,N_15164,N_15110);
nand U17847 (N_17847,N_15340,N_14123);
or U17848 (N_17848,N_15696,N_14012);
nor U17849 (N_17849,N_14194,N_15249);
nand U17850 (N_17850,N_15504,N_14165);
nor U17851 (N_17851,N_14044,N_15120);
and U17852 (N_17852,N_15893,N_14545);
and U17853 (N_17853,N_15092,N_14219);
nand U17854 (N_17854,N_14408,N_15128);
nand U17855 (N_17855,N_14131,N_15794);
nor U17856 (N_17856,N_15158,N_14429);
nor U17857 (N_17857,N_15903,N_14405);
or U17858 (N_17858,N_14132,N_15756);
or U17859 (N_17859,N_15819,N_14820);
or U17860 (N_17860,N_14522,N_15088);
nand U17861 (N_17861,N_14677,N_15056);
nand U17862 (N_17862,N_15068,N_15573);
nand U17863 (N_17863,N_15798,N_15894);
nor U17864 (N_17864,N_15975,N_15233);
or U17865 (N_17865,N_14752,N_15029);
or U17866 (N_17866,N_15294,N_14006);
or U17867 (N_17867,N_14491,N_15900);
or U17868 (N_17868,N_14371,N_15999);
nand U17869 (N_17869,N_15018,N_14953);
or U17870 (N_17870,N_15627,N_15774);
or U17871 (N_17871,N_14117,N_14672);
and U17872 (N_17872,N_14955,N_15756);
and U17873 (N_17873,N_15942,N_14670);
nand U17874 (N_17874,N_14172,N_14922);
nor U17875 (N_17875,N_14638,N_14506);
and U17876 (N_17876,N_15911,N_15144);
nand U17877 (N_17877,N_15134,N_14734);
or U17878 (N_17878,N_15208,N_15525);
or U17879 (N_17879,N_14633,N_14982);
nand U17880 (N_17880,N_15834,N_15174);
and U17881 (N_17881,N_14526,N_14830);
nand U17882 (N_17882,N_14305,N_15420);
or U17883 (N_17883,N_15693,N_14238);
and U17884 (N_17884,N_15173,N_15704);
nand U17885 (N_17885,N_14583,N_15941);
nor U17886 (N_17886,N_14004,N_14767);
nand U17887 (N_17887,N_14272,N_15466);
nand U17888 (N_17888,N_15669,N_15337);
and U17889 (N_17889,N_14484,N_15357);
or U17890 (N_17890,N_14249,N_14768);
nor U17891 (N_17891,N_14341,N_14369);
or U17892 (N_17892,N_15455,N_14122);
nand U17893 (N_17893,N_15114,N_14456);
and U17894 (N_17894,N_15897,N_15573);
nor U17895 (N_17895,N_15711,N_14687);
nand U17896 (N_17896,N_15279,N_14396);
nor U17897 (N_17897,N_15690,N_15580);
nor U17898 (N_17898,N_15176,N_15191);
nor U17899 (N_17899,N_14280,N_14718);
nand U17900 (N_17900,N_15046,N_14826);
nand U17901 (N_17901,N_14460,N_15665);
and U17902 (N_17902,N_15187,N_15835);
and U17903 (N_17903,N_14244,N_15083);
nor U17904 (N_17904,N_15609,N_14052);
or U17905 (N_17905,N_15434,N_14373);
nor U17906 (N_17906,N_14623,N_15323);
nor U17907 (N_17907,N_15880,N_14118);
nand U17908 (N_17908,N_15413,N_14010);
nand U17909 (N_17909,N_15292,N_14021);
or U17910 (N_17910,N_14962,N_14251);
nor U17911 (N_17911,N_14307,N_14034);
nand U17912 (N_17912,N_15756,N_14390);
or U17913 (N_17913,N_14858,N_15873);
nor U17914 (N_17914,N_14995,N_14623);
nor U17915 (N_17915,N_15336,N_15296);
nand U17916 (N_17916,N_15317,N_15312);
and U17917 (N_17917,N_15917,N_15946);
or U17918 (N_17918,N_15440,N_14655);
nor U17919 (N_17919,N_15088,N_15714);
nand U17920 (N_17920,N_15568,N_14904);
nor U17921 (N_17921,N_15928,N_14009);
or U17922 (N_17922,N_15009,N_14802);
nand U17923 (N_17923,N_15870,N_15824);
and U17924 (N_17924,N_14199,N_15718);
nand U17925 (N_17925,N_14824,N_14427);
nor U17926 (N_17926,N_14385,N_15030);
and U17927 (N_17927,N_14000,N_14968);
nor U17928 (N_17928,N_15423,N_14348);
nand U17929 (N_17929,N_14569,N_15948);
nand U17930 (N_17930,N_14660,N_15496);
or U17931 (N_17931,N_14607,N_15264);
nor U17932 (N_17932,N_15443,N_15579);
nand U17933 (N_17933,N_14955,N_14210);
or U17934 (N_17934,N_14487,N_14231);
or U17935 (N_17935,N_15634,N_14273);
and U17936 (N_17936,N_14842,N_15062);
and U17937 (N_17937,N_15432,N_14284);
and U17938 (N_17938,N_14804,N_14807);
nor U17939 (N_17939,N_15204,N_14719);
or U17940 (N_17940,N_14479,N_15993);
nand U17941 (N_17941,N_14662,N_14463);
nor U17942 (N_17942,N_15690,N_14664);
nor U17943 (N_17943,N_14418,N_15835);
nor U17944 (N_17944,N_15194,N_14453);
nor U17945 (N_17945,N_15065,N_14774);
or U17946 (N_17946,N_14416,N_14938);
nor U17947 (N_17947,N_14451,N_15864);
or U17948 (N_17948,N_14427,N_14178);
or U17949 (N_17949,N_14053,N_14616);
or U17950 (N_17950,N_15272,N_15705);
and U17951 (N_17951,N_14678,N_14077);
and U17952 (N_17952,N_14099,N_14431);
nand U17953 (N_17953,N_14547,N_14596);
nor U17954 (N_17954,N_14883,N_15440);
nor U17955 (N_17955,N_15670,N_14745);
xor U17956 (N_17956,N_15549,N_15592);
nor U17957 (N_17957,N_14741,N_15710);
and U17958 (N_17958,N_14860,N_14479);
or U17959 (N_17959,N_15419,N_14541);
nand U17960 (N_17960,N_14079,N_14298);
or U17961 (N_17961,N_15430,N_14270);
nor U17962 (N_17962,N_14619,N_15861);
and U17963 (N_17963,N_14875,N_15884);
and U17964 (N_17964,N_15932,N_14252);
or U17965 (N_17965,N_14872,N_15121);
and U17966 (N_17966,N_14384,N_15430);
nor U17967 (N_17967,N_14466,N_14478);
and U17968 (N_17968,N_15553,N_15165);
nor U17969 (N_17969,N_14851,N_14724);
nor U17970 (N_17970,N_15539,N_14786);
nor U17971 (N_17971,N_15934,N_15506);
or U17972 (N_17972,N_15462,N_14632);
and U17973 (N_17973,N_15344,N_14821);
nand U17974 (N_17974,N_14575,N_14896);
or U17975 (N_17975,N_15061,N_15290);
nand U17976 (N_17976,N_15262,N_14303);
or U17977 (N_17977,N_14065,N_15984);
or U17978 (N_17978,N_15106,N_15797);
or U17979 (N_17979,N_15324,N_15992);
and U17980 (N_17980,N_15585,N_14062);
xor U17981 (N_17981,N_15326,N_14935);
nor U17982 (N_17982,N_15897,N_14530);
nor U17983 (N_17983,N_15673,N_14552);
or U17984 (N_17984,N_15832,N_15032);
nor U17985 (N_17985,N_14487,N_14155);
nand U17986 (N_17986,N_14058,N_15969);
or U17987 (N_17987,N_15101,N_15323);
or U17988 (N_17988,N_14751,N_14983);
or U17989 (N_17989,N_15166,N_15135);
nor U17990 (N_17990,N_15123,N_14164);
or U17991 (N_17991,N_14343,N_14612);
and U17992 (N_17992,N_15543,N_15034);
nor U17993 (N_17993,N_14769,N_15216);
and U17994 (N_17994,N_15918,N_15870);
nor U17995 (N_17995,N_14955,N_14906);
nor U17996 (N_17996,N_14315,N_15061);
nor U17997 (N_17997,N_15152,N_15797);
nor U17998 (N_17998,N_15993,N_15844);
or U17999 (N_17999,N_14317,N_14075);
nor U18000 (N_18000,N_17931,N_16428);
or U18001 (N_18001,N_17212,N_16031);
nor U18002 (N_18002,N_16487,N_17864);
and U18003 (N_18003,N_17224,N_16764);
nand U18004 (N_18004,N_17687,N_17877);
or U18005 (N_18005,N_17738,N_16909);
nand U18006 (N_18006,N_16264,N_16113);
or U18007 (N_18007,N_17091,N_17068);
nand U18008 (N_18008,N_16825,N_17645);
nor U18009 (N_18009,N_16730,N_17934);
nand U18010 (N_18010,N_17265,N_16279);
or U18011 (N_18011,N_17794,N_17708);
or U18012 (N_18012,N_17462,N_17707);
and U18013 (N_18013,N_17333,N_16745);
and U18014 (N_18014,N_16337,N_17317);
nand U18015 (N_18015,N_16843,N_16767);
and U18016 (N_18016,N_16396,N_17267);
nand U18017 (N_18017,N_16787,N_16658);
or U18018 (N_18018,N_16102,N_17587);
and U18019 (N_18019,N_17613,N_16725);
or U18020 (N_18020,N_17621,N_17731);
nand U18021 (N_18021,N_17325,N_17921);
nor U18022 (N_18022,N_17434,N_17320);
nor U18023 (N_18023,N_17505,N_17421);
nor U18024 (N_18024,N_17319,N_17906);
nand U18025 (N_18025,N_17277,N_16702);
nand U18026 (N_18026,N_16245,N_16535);
and U18027 (N_18027,N_16806,N_16752);
or U18028 (N_18028,N_17947,N_16613);
nor U18029 (N_18029,N_16800,N_16871);
xor U18030 (N_18030,N_16099,N_17274);
and U18031 (N_18031,N_17053,N_17468);
nand U18032 (N_18032,N_17933,N_17562);
nor U18033 (N_18033,N_16551,N_16014);
nand U18034 (N_18034,N_17964,N_17181);
and U18035 (N_18035,N_17611,N_16324);
and U18036 (N_18036,N_17177,N_16603);
or U18037 (N_18037,N_16118,N_16706);
and U18038 (N_18038,N_17340,N_16075);
and U18039 (N_18039,N_16254,N_16778);
nand U18040 (N_18040,N_16464,N_17482);
and U18041 (N_18041,N_16561,N_17595);
nand U18042 (N_18042,N_17733,N_16729);
nand U18043 (N_18043,N_17169,N_16583);
nor U18044 (N_18044,N_17927,N_17291);
or U18045 (N_18045,N_17492,N_17284);
nor U18046 (N_18046,N_16612,N_16876);
nor U18047 (N_18047,N_16802,N_17263);
and U18048 (N_18048,N_17522,N_16173);
or U18049 (N_18049,N_17994,N_17406);
and U18050 (N_18050,N_16799,N_16445);
or U18051 (N_18051,N_17454,N_17629);
or U18052 (N_18052,N_17984,N_16369);
nor U18053 (N_18053,N_16441,N_16013);
nor U18054 (N_18054,N_17074,N_17575);
nor U18055 (N_18055,N_17923,N_17771);
nor U18056 (N_18056,N_16247,N_17376);
nand U18057 (N_18057,N_16550,N_17513);
nand U18058 (N_18058,N_17281,N_16309);
or U18059 (N_18059,N_17205,N_16544);
nor U18060 (N_18060,N_16125,N_16440);
or U18061 (N_18061,N_17891,N_16683);
nor U18062 (N_18062,N_16720,N_17915);
and U18063 (N_18063,N_16162,N_16616);
nand U18064 (N_18064,N_17533,N_17515);
or U18065 (N_18065,N_16803,N_16911);
or U18066 (N_18066,N_16766,N_17573);
and U18067 (N_18067,N_16169,N_17742);
or U18068 (N_18068,N_16686,N_17061);
nand U18069 (N_18069,N_17678,N_17179);
or U18070 (N_18070,N_17432,N_16626);
nor U18071 (N_18071,N_16176,N_17913);
nor U18072 (N_18072,N_16357,N_16466);
nor U18073 (N_18073,N_17694,N_17809);
nand U18074 (N_18074,N_17067,N_17995);
nor U18075 (N_18075,N_17386,N_17171);
or U18076 (N_18076,N_16444,N_17056);
nor U18077 (N_18077,N_16775,N_16220);
and U18078 (N_18078,N_17506,N_17118);
nand U18079 (N_18079,N_16159,N_17588);
and U18080 (N_18080,N_17829,N_16793);
or U18081 (N_18081,N_16966,N_17960);
and U18082 (N_18082,N_17688,N_17236);
nand U18083 (N_18083,N_17559,N_17627);
nor U18084 (N_18084,N_16788,N_17603);
nor U18085 (N_18085,N_17303,N_17502);
or U18086 (N_18086,N_17845,N_16841);
and U18087 (N_18087,N_16414,N_16387);
and U18088 (N_18088,N_17422,N_16978);
and U18089 (N_18089,N_17431,N_17347);
nand U18090 (N_18090,N_16804,N_16281);
or U18091 (N_18091,N_16164,N_16867);
nand U18092 (N_18092,N_17836,N_16827);
or U18093 (N_18093,N_16680,N_17956);
nand U18094 (N_18094,N_17088,N_16557);
or U18095 (N_18095,N_16826,N_16252);
and U18096 (N_18096,N_17175,N_17199);
nor U18097 (N_18097,N_16060,N_16861);
or U18098 (N_18098,N_17736,N_16079);
nand U18099 (N_18099,N_16246,N_16709);
or U18100 (N_18100,N_16988,N_17709);
nor U18101 (N_18101,N_16455,N_16366);
nor U18102 (N_18102,N_17391,N_17498);
nand U18103 (N_18103,N_16289,N_17814);
nor U18104 (N_18104,N_17804,N_16740);
or U18105 (N_18105,N_16157,N_16419);
nand U18106 (N_18106,N_16644,N_17894);
nor U18107 (N_18107,N_16738,N_17965);
nand U18108 (N_18108,N_16580,N_17892);
and U18109 (N_18109,N_16648,N_16393);
nor U18110 (N_18110,N_16772,N_17474);
nor U18111 (N_18111,N_16870,N_17677);
nand U18112 (N_18112,N_17527,N_17381);
nand U18113 (N_18113,N_16552,N_16615);
nor U18114 (N_18114,N_16748,N_16307);
nand U18115 (N_18115,N_17970,N_16946);
nand U18116 (N_18116,N_17801,N_16574);
nand U18117 (N_18117,N_16833,N_17624);
nand U18118 (N_18118,N_16822,N_16558);
and U18119 (N_18119,N_17125,N_17747);
or U18120 (N_18120,N_16878,N_16992);
or U18121 (N_18121,N_17959,N_17282);
and U18122 (N_18122,N_16923,N_16111);
nand U18123 (N_18123,N_16659,N_16210);
nor U18124 (N_18124,N_17697,N_17403);
and U18125 (N_18125,N_17919,N_17417);
nor U18126 (N_18126,N_17461,N_16668);
and U18127 (N_18127,N_16547,N_17252);
or U18128 (N_18128,N_17117,N_17479);
nor U18129 (N_18129,N_16081,N_16652);
nor U18130 (N_18130,N_17626,N_17761);
nand U18131 (N_18131,N_17321,N_17350);
nand U18132 (N_18132,N_17718,N_16721);
and U18133 (N_18133,N_16965,N_16782);
nor U18134 (N_18134,N_17285,N_17076);
and U18135 (N_18135,N_16527,N_16314);
nor U18136 (N_18136,N_16065,N_16687);
nor U18137 (N_18137,N_16071,N_17485);
nand U18138 (N_18138,N_17180,N_16947);
or U18139 (N_18139,N_16585,N_17210);
nor U18140 (N_18140,N_16678,N_17589);
or U18141 (N_18141,N_16776,N_17401);
and U18142 (N_18142,N_16724,N_17765);
nor U18143 (N_18143,N_16167,N_16614);
nand U18144 (N_18144,N_17246,N_16633);
nand U18145 (N_18145,N_16136,N_17021);
nor U18146 (N_18146,N_17800,N_17726);
nand U18147 (N_18147,N_16926,N_17193);
nand U18148 (N_18148,N_16589,N_16402);
nand U18149 (N_18149,N_17173,N_17574);
nand U18150 (N_18150,N_16274,N_17930);
xnor U18151 (N_18151,N_17135,N_16215);
nand U18152 (N_18152,N_16945,N_16912);
nor U18153 (N_18153,N_17238,N_17602);
or U18154 (N_18154,N_16622,N_17618);
nand U18155 (N_18155,N_16261,N_16781);
nor U18156 (N_18156,N_17969,N_16045);
xnor U18157 (N_18157,N_16001,N_17767);
and U18158 (N_18158,N_17751,N_17090);
or U18159 (N_18159,N_16650,N_17055);
nor U18160 (N_18160,N_17197,N_16457);
and U18161 (N_18161,N_17693,N_17571);
nand U18162 (N_18162,N_16395,N_16762);
and U18163 (N_18163,N_17614,N_17288);
and U18164 (N_18164,N_17393,N_16932);
or U18165 (N_18165,N_16524,N_17245);
nor U18166 (N_18166,N_16592,N_16479);
nor U18167 (N_18167,N_16488,N_17107);
nand U18168 (N_18168,N_16999,N_16222);
nor U18169 (N_18169,N_17858,N_17052);
and U18170 (N_18170,N_16098,N_16231);
nor U18171 (N_18171,N_16342,N_16877);
nand U18172 (N_18172,N_16134,N_16760);
nor U18173 (N_18173,N_16105,N_17990);
and U18174 (N_18174,N_17341,N_16278);
nand U18175 (N_18175,N_17841,N_17186);
or U18176 (N_18176,N_16543,N_17172);
or U18177 (N_18177,N_17248,N_17781);
and U18178 (N_18178,N_16373,N_16830);
and U18179 (N_18179,N_17371,N_16838);
or U18180 (N_18180,N_17062,N_17988);
nand U18181 (N_18181,N_17951,N_16052);
nor U18182 (N_18182,N_17483,N_17811);
or U18183 (N_18183,N_16186,N_16602);
nor U18184 (N_18184,N_16203,N_17441);
nand U18185 (N_18185,N_16413,N_16801);
nand U18186 (N_18186,N_16979,N_16914);
nand U18187 (N_18187,N_16447,N_17493);
or U18188 (N_18188,N_16213,N_17328);
and U18189 (N_18189,N_16795,N_17685);
or U18190 (N_18190,N_16915,N_17047);
nand U18191 (N_18191,N_17475,N_17878);
or U18192 (N_18192,N_16200,N_16392);
or U18193 (N_18193,N_16175,N_17208);
and U18194 (N_18194,N_16107,N_16423);
or U18195 (N_18195,N_17779,N_17191);
and U18196 (N_18196,N_16416,N_16991);
or U18197 (N_18197,N_16636,N_16785);
or U18198 (N_18198,N_16844,N_16901);
nand U18199 (N_18199,N_17057,N_17636);
nor U18200 (N_18200,N_16707,N_16860);
xor U18201 (N_18201,N_17598,N_16061);
nor U18202 (N_18202,N_17564,N_16197);
nor U18203 (N_18203,N_16382,N_17108);
nand U18204 (N_18204,N_16759,N_16670);
nand U18205 (N_18205,N_17448,N_17665);
and U18206 (N_18206,N_17433,N_17999);
and U18207 (N_18207,N_16989,N_16091);
nor U18208 (N_18208,N_17937,N_17360);
nor U18209 (N_18209,N_16971,N_17223);
or U18210 (N_18210,N_16051,N_17194);
and U18211 (N_18211,N_17259,N_17842);
and U18212 (N_18212,N_17338,N_16501);
nor U18213 (N_18213,N_17049,N_16831);
xor U18214 (N_18214,N_16009,N_17080);
nand U18215 (N_18215,N_17949,N_16886);
nand U18216 (N_18216,N_16913,N_17922);
nor U18217 (N_18217,N_17854,N_16238);
nand U18218 (N_18218,N_16887,N_17983);
nor U18219 (N_18219,N_17550,N_17002);
nand U18220 (N_18220,N_16437,N_17942);
nor U18221 (N_18221,N_17046,N_17941);
and U18222 (N_18222,N_17012,N_16828);
and U18223 (N_18223,N_17287,N_17565);
and U18224 (N_18224,N_17901,N_17762);
nand U18225 (N_18225,N_17240,N_16951);
nand U18226 (N_18226,N_16773,N_16267);
nor U18227 (N_18227,N_16746,N_17227);
nor U18228 (N_18228,N_17642,N_17528);
nand U18229 (N_18229,N_16899,N_16076);
and U18230 (N_18230,N_17330,N_16536);
nor U18231 (N_18231,N_17170,N_16798);
nor U18232 (N_18232,N_16345,N_17536);
nor U18233 (N_18233,N_16150,N_17404);
xnor U18234 (N_18234,N_16146,N_16884);
or U18235 (N_18235,N_16360,N_17644);
nand U18236 (N_18236,N_16634,N_17250);
nor U18237 (N_18237,N_17048,N_16185);
or U18238 (N_18238,N_17608,N_17022);
or U18239 (N_18239,N_16655,N_16050);
and U18240 (N_18240,N_16205,N_17799);
and U18241 (N_18241,N_17982,N_16832);
or U18242 (N_18242,N_17398,N_17719);
and U18243 (N_18243,N_16008,N_17791);
nor U18244 (N_18244,N_17980,N_17449);
and U18245 (N_18245,N_16599,N_17129);
and U18246 (N_18246,N_16684,N_16755);
nand U18247 (N_18247,N_17145,N_17016);
or U18248 (N_18248,N_17152,N_17416);
and U18249 (N_18249,N_16212,N_16119);
nor U18250 (N_18250,N_16969,N_16509);
nand U18251 (N_18251,N_17499,N_16930);
or U18252 (N_18252,N_17324,N_16500);
and U18253 (N_18253,N_17774,N_17123);
nand U18254 (N_18254,N_17552,N_16862);
nand U18255 (N_18255,N_16041,N_17534);
and U18256 (N_18256,N_16957,N_17063);
and U18257 (N_18257,N_17429,N_17342);
or U18258 (N_18258,N_16904,N_16704);
and U18259 (N_18259,N_17201,N_17030);
and U18260 (N_18260,N_16528,N_16410);
nor U18261 (N_18261,N_17759,N_17702);
nor U18262 (N_18262,N_17509,N_16713);
nor U18263 (N_18263,N_16718,N_16619);
nand U18264 (N_18264,N_17083,N_17716);
nand U18265 (N_18265,N_17355,N_16866);
or U18266 (N_18266,N_17242,N_16556);
or U18267 (N_18267,N_17008,N_16179);
nor U18268 (N_18268,N_17436,N_16232);
or U18269 (N_18269,N_16386,N_16390);
and U18270 (N_18270,N_17489,N_16977);
and U18271 (N_18271,N_17549,N_17737);
or U18272 (N_18272,N_17418,N_17467);
and U18273 (N_18273,N_16350,N_16259);
nor U18274 (N_18274,N_17495,N_16019);
nor U18275 (N_18275,N_17308,N_16303);
and U18276 (N_18276,N_17997,N_17953);
nand U18277 (N_18277,N_16888,N_17655);
and U18278 (N_18278,N_16943,N_16056);
nand U18279 (N_18279,N_16430,N_16266);
nand U18280 (N_18280,N_17300,N_16600);
nand U18281 (N_18281,N_17302,N_16216);
or U18282 (N_18282,N_17810,N_17542);
nor U18283 (N_18283,N_17860,N_16406);
and U18284 (N_18284,N_16623,N_17200);
and U18285 (N_18285,N_17748,N_17184);
and U18286 (N_18286,N_16021,N_17093);
and U18287 (N_18287,N_16834,N_16515);
xnor U18288 (N_18288,N_17615,N_17396);
or U18289 (N_18289,N_16507,N_16288);
or U18290 (N_18290,N_16950,N_17410);
nand U18291 (N_18291,N_16554,N_16319);
and U18292 (N_18292,N_17299,N_16399);
nand U18293 (N_18293,N_17554,N_16074);
nor U18294 (N_18294,N_16123,N_16070);
or U18295 (N_18295,N_16273,N_17222);
and U18296 (N_18296,N_17204,N_17440);
and U18297 (N_18297,N_16473,N_17745);
nand U18298 (N_18298,N_17374,N_16058);
and U18299 (N_18299,N_17657,N_17546);
or U18300 (N_18300,N_17698,N_17981);
or U18301 (N_18301,N_17018,N_17815);
or U18302 (N_18302,N_16953,N_17419);
nor U18303 (N_18303,N_16864,N_17523);
nor U18304 (N_18304,N_16491,N_16715);
or U18305 (N_18305,N_16218,N_17189);
or U18306 (N_18306,N_17666,N_17312);
nand U18307 (N_18307,N_16891,N_17793);
and U18308 (N_18308,N_17798,N_17974);
and U18309 (N_18309,N_16100,N_17544);
or U18310 (N_18310,N_17221,N_16331);
or U18311 (N_18311,N_17889,N_17682);
and U18312 (N_18312,N_17789,N_17161);
and U18313 (N_18313,N_17622,N_17477);
nand U18314 (N_18314,N_17442,N_16918);
nand U18315 (N_18315,N_17060,N_16133);
nand U18316 (N_18316,N_16598,N_17273);
nand U18317 (N_18317,N_16874,N_16629);
or U18318 (N_18318,N_17881,N_16510);
nor U18319 (N_18319,N_17993,N_16171);
nand U18320 (N_18320,N_16757,N_16090);
nand U18321 (N_18321,N_17961,N_17917);
or U18322 (N_18322,N_17986,N_17343);
nor U18323 (N_18323,N_17547,N_16809);
nand U18324 (N_18324,N_16627,N_17451);
and U18325 (N_18325,N_17672,N_17024);
or U18326 (N_18326,N_16810,N_17887);
and U18327 (N_18327,N_16868,N_17111);
nor U18328 (N_18328,N_16865,N_16442);
nand U18329 (N_18329,N_17309,N_16676);
and U18330 (N_18330,N_16010,N_17757);
or U18331 (N_18331,N_16401,N_17078);
or U18332 (N_18332,N_17846,N_17648);
and U18333 (N_18333,N_17213,N_17883);
nor U18334 (N_18334,N_16240,N_17151);
and U18335 (N_18335,N_17220,N_17459);
or U18336 (N_18336,N_16845,N_17137);
and U18337 (N_18337,N_17103,N_17604);
and U18338 (N_18338,N_16304,N_16114);
or U18339 (N_18339,N_16370,N_16165);
nor U18340 (N_18340,N_17476,N_17367);
or U18341 (N_18341,N_17007,N_17607);
nor U18342 (N_18342,N_17813,N_16849);
and U18343 (N_18343,N_16086,N_16421);
and U18344 (N_18344,N_17992,N_17163);
and U18345 (N_18345,N_17714,N_17428);
nor U18346 (N_18346,N_16316,N_16642);
nand U18347 (N_18347,N_17147,N_17700);
nor U18348 (N_18348,N_16062,N_16937);
nor U18349 (N_18349,N_16483,N_16910);
and U18350 (N_18350,N_16753,N_17821);
and U18351 (N_18351,N_17397,N_17668);
nand U18352 (N_18352,N_17834,N_16530);
or U18353 (N_18353,N_16756,N_16028);
nor U18354 (N_18354,N_17795,N_16939);
or U18355 (N_18355,N_17950,N_16270);
or U18356 (N_18356,N_17031,N_17262);
or U18357 (N_18357,N_17085,N_16587);
nor U18358 (N_18358,N_17732,N_16198);
nor U18359 (N_18359,N_16540,N_17148);
nor U18360 (N_18360,N_16452,N_16078);
nand U18361 (N_18361,N_17803,N_17863);
nor U18362 (N_18362,N_16996,N_17026);
and U18363 (N_18363,N_16941,N_16701);
or U18364 (N_18364,N_17596,N_16879);
nor U18365 (N_18365,N_16195,N_17674);
nor U18366 (N_18366,N_17207,N_16496);
and U18367 (N_18367,N_17069,N_16570);
nand U18368 (N_18368,N_17383,N_17802);
and U18369 (N_18369,N_17211,N_17132);
and U18370 (N_18370,N_16381,N_17070);
or U18371 (N_18371,N_17870,N_16434);
or U18372 (N_18372,N_17165,N_16258);
or U18373 (N_18373,N_17399,N_16117);
and U18374 (N_18374,N_17192,N_17258);
nor U18375 (N_18375,N_17480,N_17849);
and U18376 (N_18376,N_16694,N_16958);
nand U18377 (N_18377,N_17743,N_17890);
nand U18378 (N_18378,N_17297,N_17124);
or U18379 (N_18379,N_16840,N_16448);
nor U18380 (N_18380,N_16533,N_16476);
or U18381 (N_18381,N_17412,N_17038);
or U18382 (N_18382,N_17840,N_17364);
nand U18383 (N_18383,N_16549,N_16362);
and U18384 (N_18384,N_16542,N_16204);
and U18385 (N_18385,N_16330,N_16214);
and U18386 (N_18386,N_16974,N_16007);
and U18387 (N_18387,N_16039,N_17149);
nand U18388 (N_18388,N_17345,N_17365);
nor U18389 (N_18389,N_16815,N_16068);
or U18390 (N_18390,N_16379,N_17833);
nor U18391 (N_18391,N_16905,N_17957);
and U18392 (N_18392,N_16161,N_16225);
and U18393 (N_18393,N_16053,N_16997);
or U18394 (N_18394,N_17033,N_17897);
nand U18395 (N_18395,N_16143,N_16618);
or U18396 (N_18396,N_16588,N_16226);
nand U18397 (N_18397,N_16127,N_17384);
nor U18398 (N_18398,N_17918,N_17253);
or U18399 (N_18399,N_16523,N_16120);
and U18400 (N_18400,N_17156,N_16727);
nor U18401 (N_18401,N_16579,N_17827);
nor U18402 (N_18402,N_16178,N_17879);
or U18403 (N_18403,N_17042,N_16451);
and U18404 (N_18404,N_16145,N_17592);
and U18405 (N_18405,N_16504,N_16191);
nor U18406 (N_18406,N_17243,N_17543);
nor U18407 (N_18407,N_17017,N_16454);
nand U18408 (N_18408,N_17576,N_16881);
nand U18409 (N_18409,N_17867,N_17099);
nand U18410 (N_18410,N_17120,N_17154);
nand U18411 (N_18411,N_17659,N_16708);
nor U18412 (N_18412,N_17235,N_17643);
and U18413 (N_18413,N_17444,N_17348);
nor U18414 (N_18414,N_17209,N_16903);
nor U18415 (N_18415,N_16073,N_16995);
nand U18416 (N_18416,N_16697,N_16621);
nor U18417 (N_18417,N_16131,N_17473);
nand U18418 (N_18418,N_16181,N_17712);
nor U18419 (N_18419,N_17039,N_17978);
or U18420 (N_18420,N_17553,N_16080);
nand U18421 (N_18421,N_16148,N_17368);
or U18422 (N_18422,N_16325,N_16377);
and U18423 (N_18423,N_16223,N_16765);
nor U18424 (N_18424,N_16519,N_16332);
and U18425 (N_18425,N_16716,N_17301);
and U18426 (N_18426,N_17128,N_17112);
nor U18427 (N_18427,N_16987,N_17435);
or U18428 (N_18428,N_16272,N_16320);
and U18429 (N_18429,N_17455,N_16894);
nand U18430 (N_18430,N_17102,N_17405);
or U18431 (N_18431,N_17239,N_17739);
nor U18432 (N_18432,N_16057,N_17071);
or U18433 (N_18433,N_16734,N_16217);
or U18434 (N_18434,N_16567,N_16235);
nand U18435 (N_18435,N_16166,N_17295);
nor U18436 (N_18436,N_17187,N_16449);
nor U18437 (N_18437,N_17050,N_16532);
and U18438 (N_18438,N_16959,N_17443);
or U18439 (N_18439,N_16685,N_16088);
or U18440 (N_18440,N_16172,N_17486);
or U18441 (N_18441,N_17020,N_16135);
nand U18442 (N_18442,N_16571,N_17585);
nand U18443 (N_18443,N_16002,N_16671);
nand U18444 (N_18444,N_16949,N_17601);
nor U18445 (N_18445,N_16572,N_17681);
xnor U18446 (N_18446,N_16842,N_17667);
nand U18447 (N_18447,N_16372,N_17457);
or U18448 (N_18448,N_16016,N_17975);
and U18449 (N_18449,N_17530,N_17121);
or U18450 (N_18450,N_16494,N_16326);
nand U18451 (N_18451,N_17059,N_16174);
or U18452 (N_18452,N_17723,N_16461);
nand U18453 (N_18453,N_17520,N_16339);
or U18454 (N_18454,N_17658,N_17126);
or U18455 (N_18455,N_16749,N_17283);
and U18456 (N_18456,N_17280,N_16679);
nor U18457 (N_18457,N_17407,N_16450);
or U18458 (N_18458,N_17230,N_16696);
nor U18459 (N_18459,N_16968,N_16639);
nor U18460 (N_18460,N_17635,N_17825);
or U18461 (N_18461,N_16285,N_17684);
nor U18462 (N_18462,N_17649,N_17855);
or U18463 (N_18463,N_16541,N_16993);
and U18464 (N_18464,N_16420,N_16722);
nand U18465 (N_18465,N_17661,N_17402);
nor U18466 (N_18466,N_16812,N_17939);
nand U18467 (N_18467,N_16431,N_16147);
or U18468 (N_18468,N_17127,N_16893);
nand U18469 (N_18469,N_17948,N_17054);
and U18470 (N_18470,N_17247,N_16385);
and U18471 (N_18471,N_16699,N_16485);
or U18472 (N_18472,N_16689,N_17721);
and U18473 (N_18473,N_16230,N_17786);
or U18474 (N_18474,N_16083,N_17569);
nand U18475 (N_18475,N_16106,N_16069);
and U18476 (N_18476,N_17269,N_16375);
or U18477 (N_18477,N_17298,N_17812);
or U18478 (N_18478,N_16383,N_16816);
or U18479 (N_18479,N_16768,N_17178);
and U18480 (N_18480,N_16952,N_17346);
nand U18481 (N_18481,N_17518,N_16705);
or U18482 (N_18482,N_17326,N_17414);
or U18483 (N_18483,N_16460,N_17164);
and U18484 (N_18484,N_17058,N_17647);
and U18485 (N_18485,N_16737,N_17219);
nor U18486 (N_18486,N_16415,N_17514);
nand U18487 (N_18487,N_17260,N_17377);
nor U18488 (N_18488,N_17734,N_16286);
or U18489 (N_18489,N_16525,N_16066);
nand U18490 (N_18490,N_17578,N_16620);
or U18491 (N_18491,N_16265,N_17689);
and U18492 (N_18492,N_17293,N_16249);
nor U18493 (N_18493,N_16020,N_16934);
and U18494 (N_18494,N_17653,N_17214);
nor U18495 (N_18495,N_16469,N_16139);
xor U18496 (N_18496,N_17563,N_16731);
nand U18497 (N_18497,N_16835,N_17362);
nor U18498 (N_18498,N_16856,N_16624);
and U18499 (N_18499,N_16703,N_17160);
nor U18500 (N_18500,N_17032,N_16486);
or U18501 (N_18501,N_17000,N_17472);
and U18502 (N_18502,N_17579,N_16022);
nand U18503 (N_18503,N_17512,N_16417);
nand U18504 (N_18504,N_16365,N_16408);
nand U18505 (N_18505,N_17869,N_17634);
and U18506 (N_18506,N_17828,N_16610);
or U18507 (N_18507,N_16004,N_17532);
nor U18508 (N_18508,N_17884,N_16733);
and U18509 (N_18509,N_16294,N_16649);
nand U18510 (N_18510,N_16817,N_16608);
nand U18511 (N_18511,N_17760,N_17851);
and U18512 (N_18512,N_17508,N_16889);
nor U18513 (N_18513,N_17469,N_17307);
or U18514 (N_18514,N_17914,N_17797);
and U18515 (N_18515,N_17511,N_16682);
nand U18516 (N_18516,N_17491,N_16346);
or U18517 (N_18517,N_16654,N_17226);
nor U18518 (N_18518,N_16981,N_17591);
and U18519 (N_18519,N_17380,N_17976);
nand U18520 (N_18520,N_17713,N_16575);
or U18521 (N_18521,N_16468,N_16282);
and U18522 (N_18522,N_17847,N_17203);
or U18523 (N_18523,N_17305,N_16935);
nand U18524 (N_18524,N_17599,N_16628);
or U18525 (N_18525,N_17967,N_17837);
and U18526 (N_18526,N_17727,N_16499);
nand U18527 (N_18527,N_16582,N_16333);
and U18528 (N_18528,N_16154,N_16902);
nand U18529 (N_18529,N_16153,N_16662);
nor U18530 (N_18530,N_17616,N_16681);
and U18531 (N_18531,N_17873,N_17640);
or U18532 (N_18532,N_16436,N_17823);
and U18533 (N_18533,N_17857,N_16044);
and U18534 (N_18534,N_16569,N_17133);
nor U18535 (N_18535,N_17671,N_16677);
nor U18536 (N_18536,N_16596,N_16783);
or U18537 (N_18537,N_16617,N_16474);
nand U18538 (N_18538,N_16409,N_16818);
and U18539 (N_18539,N_17865,N_16811);
and U18540 (N_18540,N_17216,N_16368);
and U18541 (N_18541,N_17232,N_16189);
or U18542 (N_18542,N_16710,N_16666);
and U18543 (N_18543,N_17159,N_16023);
and U18544 (N_18544,N_17670,N_16269);
or U18545 (N_18545,N_17540,N_17989);
nor U18546 (N_18546,N_17507,N_17037);
or U18547 (N_18547,N_16163,N_16660);
and U18548 (N_18548,N_17484,N_17095);
nand U18549 (N_18549,N_17334,N_16526);
or U18550 (N_18550,N_17379,N_16643);
nand U18551 (N_18551,N_17787,N_16298);
or U18552 (N_18552,N_16789,N_17217);
nor U18553 (N_18553,N_16590,N_17251);
or U18554 (N_18554,N_16607,N_17490);
nand U18555 (N_18555,N_17357,N_16182);
and U18556 (N_18556,N_16609,N_16371);
nand U18557 (N_18557,N_17415,N_16211);
nand U18558 (N_18558,N_16378,N_16097);
or U18559 (N_18559,N_16072,N_17072);
or U18560 (N_18560,N_17354,N_17051);
nor U18561 (N_18561,N_17991,N_17369);
nand U18562 (N_18562,N_17503,N_16647);
and U18563 (N_18563,N_16597,N_16638);
nor U18564 (N_18564,N_17775,N_16446);
nand U18565 (N_18565,N_17504,N_16391);
nand U18566 (N_18566,N_16805,N_17423);
and U18567 (N_18567,N_16857,N_17086);
and U18568 (N_18568,N_17977,N_16924);
and U18569 (N_18569,N_17409,N_17703);
and U18570 (N_18570,N_17706,N_17438);
nand U18571 (N_18571,N_16354,N_17231);
nor U18572 (N_18572,N_17390,N_16892);
nand U18573 (N_18573,N_16741,N_17692);
and U18574 (N_18574,N_17521,N_17646);
and U18575 (N_18575,N_17639,N_16443);
or U18576 (N_18576,N_16975,N_17594);
or U18577 (N_18577,N_16439,N_17567);
nor U18578 (N_18578,N_17876,N_16819);
nor U18579 (N_18579,N_17710,N_16201);
and U18580 (N_18580,N_17044,N_17625);
nand U18581 (N_18581,N_17660,N_16328);
or U18582 (N_18582,N_16955,N_17335);
nand U18583 (N_18583,N_16898,N_17763);
nand U18584 (N_18584,N_16553,N_16035);
or U18585 (N_18585,N_16714,N_17104);
and U18586 (N_18586,N_16290,N_16922);
and U18587 (N_18587,N_17788,N_17065);
and U18588 (N_18588,N_17385,N_16064);
and U18589 (N_18589,N_16531,N_16712);
and U18590 (N_18590,N_16435,N_17339);
and U18591 (N_18591,N_16239,N_16492);
or U18592 (N_18592,N_16471,N_17704);
nand U18593 (N_18593,N_16661,N_17623);
or U18594 (N_18594,N_17106,N_16093);
nand U18595 (N_18595,N_17420,N_16140);
and U18596 (N_18596,N_17525,N_16555);
or U18597 (N_18597,N_16637,N_16854);
and U18598 (N_18598,N_17754,N_16095);
and U18599 (N_18599,N_17306,N_17555);
or U18600 (N_18600,N_17075,N_16846);
and U18601 (N_18601,N_16944,N_16851);
nor U18602 (N_18602,N_17905,N_16276);
nor U18603 (N_18603,N_17264,N_16970);
or U18604 (N_18604,N_16347,N_17304);
nand U18605 (N_18605,N_17749,N_16132);
or U18606 (N_18606,N_17773,N_17673);
nor U18607 (N_18607,N_17885,N_17735);
or U18608 (N_18608,N_17370,N_17874);
nor U18609 (N_18609,N_17935,N_17497);
nand U18610 (N_18610,N_16017,N_16026);
nand U18611 (N_18611,N_16277,N_17566);
nand U18612 (N_18612,N_17966,N_17105);
or U18613 (N_18613,N_17336,N_16190);
and U18614 (N_18614,N_17463,N_17144);
or U18615 (N_18615,N_16361,N_17958);
nor U18616 (N_18616,N_17850,N_16293);
or U18617 (N_18617,N_16635,N_17551);
and U18618 (N_18618,N_17537,N_16335);
and U18619 (N_18619,N_16769,N_16824);
nor U18620 (N_18620,N_17375,N_17830);
or U18621 (N_18621,N_16962,N_16470);
or U18622 (N_18622,N_17630,N_16334);
nor U18623 (N_18623,N_17822,N_17899);
nor U18624 (N_18624,N_16480,N_16537);
or U18625 (N_18625,N_17651,N_16438);
and U18626 (N_18626,N_17316,N_17859);
or U18627 (N_18627,N_16593,N_16750);
nand U18628 (N_18628,N_17278,N_16233);
or U18629 (N_18629,N_17926,N_17359);
nand U18630 (N_18630,N_17073,N_17331);
nor U18631 (N_18631,N_17349,N_16604);
and U18632 (N_18632,N_17122,N_16576);
or U18633 (N_18633,N_17029,N_16717);
or U18634 (N_18634,N_17817,N_16241);
nand U18635 (N_18635,N_16518,N_16158);
nor U18636 (N_18636,N_17089,N_16327);
nand U18637 (N_18637,N_17447,N_17971);
or U18638 (N_18638,N_16046,N_16092);
or U18639 (N_18639,N_17777,N_16084);
and U18640 (N_18640,N_16219,N_16318);
nand U18641 (N_18641,N_16770,N_16156);
nand U18642 (N_18642,N_17494,N_16126);
or U18643 (N_18643,N_16508,N_17488);
nor U18644 (N_18644,N_17952,N_16790);
nor U18645 (N_18645,N_16493,N_16433);
or U18646 (N_18646,N_16183,N_16358);
nor U18647 (N_18647,N_17344,N_17453);
nor U18648 (N_18648,N_17456,N_16594);
nand U18649 (N_18649,N_17272,N_16641);
nor U18650 (N_18650,N_16367,N_16196);
or U18651 (N_18651,N_17526,N_16115);
nor U18652 (N_18652,N_17844,N_16927);
or U18653 (N_18653,N_16306,N_17916);
nor U18654 (N_18654,N_17987,N_17577);
or U18655 (N_18655,N_16723,N_16963);
and U18656 (N_18656,N_17198,N_17938);
nor U18657 (N_18657,N_16498,N_17437);
nor U18658 (N_18658,N_16049,N_16412);
and U18659 (N_18659,N_16025,N_17556);
nor U18660 (N_18660,N_17755,N_16771);
xor U18661 (N_18661,N_17425,N_16227);
nor U18662 (N_18662,N_16895,N_17696);
or U18663 (N_18663,N_16037,N_17943);
or U18664 (N_18664,N_16400,N_17650);
nand U18665 (N_18665,N_17818,N_16122);
and U18666 (N_18666,N_17541,N_16085);
and U18667 (N_18667,N_16458,N_16630);
nand U18668 (N_18668,N_17750,N_17619);
nor U18669 (N_18669,N_17464,N_16137);
nor U18670 (N_18670,N_16465,N_17167);
nand U18671 (N_18671,N_16961,N_17924);
nor U18672 (N_18672,N_17932,N_17327);
and U18673 (N_18673,N_16983,N_17256);
nand U18674 (N_18674,N_17676,N_17158);
nand U18675 (N_18675,N_16268,N_16209);
nand U18676 (N_18676,N_16384,N_17780);
nand U18677 (N_18677,N_16796,N_16967);
or U18678 (N_18678,N_16728,N_16692);
or U18679 (N_18679,N_17168,N_17558);
nand U18680 (N_18680,N_17866,N_17389);
or U18681 (N_18681,N_17356,N_17322);
nand U18682 (N_18682,N_16631,N_17332);
xnor U18683 (N_18683,N_17925,N_17531);
nor U18684 (N_18684,N_16024,N_16513);
nand U18685 (N_18685,N_16726,N_17820);
and U18686 (N_18686,N_16459,N_17446);
nor U18687 (N_18687,N_16792,N_16168);
and U18688 (N_18688,N_16149,N_16380);
or U18689 (N_18689,N_17560,N_16006);
nor U18690 (N_18690,N_16883,N_16732);
and U18691 (N_18691,N_17430,N_16917);
and U18692 (N_18692,N_16152,N_16497);
and U18693 (N_18693,N_17234,N_17580);
nor U18694 (N_18694,N_16869,N_16012);
nand U18695 (N_18695,N_16315,N_17257);
nor U18696 (N_18696,N_16038,N_16916);
nand U18697 (N_18697,N_16047,N_17758);
nand U18698 (N_18698,N_16960,N_17139);
and U18699 (N_18699,N_16940,N_16780);
nand U18700 (N_18700,N_16151,N_17311);
nand U18701 (N_18701,N_16651,N_16398);
nand U18702 (N_18702,N_16807,N_16018);
and U18703 (N_18703,N_16177,N_16467);
nand U18704 (N_18704,N_16674,N_16043);
or U18705 (N_18705,N_17146,N_17772);
nand U18706 (N_18706,N_17119,N_17077);
nand U18707 (N_18707,N_17826,N_17911);
nand U18708 (N_18708,N_16973,N_16925);
nand U18709 (N_18709,N_17411,N_16427);
nand U18710 (N_18710,N_17768,N_17084);
nand U18711 (N_18711,N_17286,N_16984);
nor U18712 (N_18712,N_17912,N_16193);
nand U18713 (N_18713,N_17557,N_16170);
nand U18714 (N_18714,N_17011,N_16251);
nor U18715 (N_18715,N_17395,N_17519);
nor U18716 (N_18716,N_16994,N_17568);
or U18717 (N_18717,N_16067,N_16343);
nand U18718 (N_18718,N_16284,N_17378);
or U18719 (N_18719,N_16321,N_16094);
nor U18720 (N_18720,N_17944,N_17294);
and U18721 (N_18721,N_17015,N_16128);
or U18722 (N_18722,N_17664,N_17097);
nor U18723 (N_18723,N_17861,N_17096);
nand U18724 (N_18724,N_16850,N_16322);
nand U18725 (N_18725,N_16972,N_16356);
nand U18726 (N_18726,N_17394,N_17806);
and U18727 (N_18727,N_16029,N_16929);
nor U18728 (N_18728,N_17631,N_16820);
and U18729 (N_18729,N_17848,N_16489);
nand U18730 (N_18730,N_16605,N_16144);
nor U18731 (N_18731,N_17450,N_17756);
and U18732 (N_18732,N_17190,N_16242);
and U18733 (N_18733,N_16688,N_16908);
or U18734 (N_18734,N_16188,N_17581);
nor U18735 (N_18735,N_17517,N_17606);
nand U18736 (N_18736,N_16938,N_17109);
nand U18737 (N_18737,N_17400,N_16089);
and U18738 (N_18738,N_16669,N_17720);
and U18739 (N_18739,N_17632,N_16980);
or U18740 (N_18740,N_17496,N_17142);
and U18741 (N_18741,N_16657,N_16863);
nand U18742 (N_18742,N_17153,N_17439);
and U18743 (N_18743,N_17202,N_17680);
nor U18744 (N_18744,N_16890,N_16852);
nor U18745 (N_18745,N_17796,N_16287);
nand U18746 (N_18746,N_16300,N_17136);
nor U18747 (N_18747,N_17510,N_16275);
or U18748 (N_18748,N_17832,N_17289);
or U18749 (N_18749,N_16928,N_17155);
and U18750 (N_18750,N_17353,N_16034);
nor U18751 (N_18751,N_16711,N_16853);
nand U18752 (N_18752,N_16990,N_17638);
nand U18753 (N_18753,N_17195,N_16184);
nand U18754 (N_18754,N_16040,N_16224);
or U18755 (N_18755,N_17516,N_17729);
or U18756 (N_18756,N_16581,N_17466);
and U18757 (N_18757,N_16698,N_17426);
and U18758 (N_18758,N_16921,N_16244);
nor U18759 (N_18759,N_16665,N_17373);
nor U18760 (N_18760,N_17705,N_16942);
nand U18761 (N_18761,N_17004,N_16794);
and U18762 (N_18762,N_17752,N_16397);
or U18763 (N_18763,N_17764,N_16426);
or U18764 (N_18764,N_16048,N_17679);
nor U18765 (N_18765,N_16155,N_16221);
nand U18766 (N_18766,N_16747,N_16207);
and U18767 (N_18767,N_16104,N_17633);
xnor U18768 (N_18768,N_17722,N_16763);
nand U18769 (N_18769,N_16885,N_17290);
nor U18770 (N_18770,N_16077,N_16063);
nor U18771 (N_18771,N_16411,N_17620);
nand U18772 (N_18772,N_16129,N_16003);
nor U18773 (N_18773,N_17101,N_17296);
or U18774 (N_18774,N_16664,N_17535);
nand U18775 (N_18775,N_17157,N_17313);
or U18776 (N_18776,N_16055,N_16472);
and U18777 (N_18777,N_17996,N_16341);
and U18778 (N_18778,N_16394,N_16663);
nand U18779 (N_18779,N_17092,N_16425);
nor U18780 (N_18780,N_17529,N_17465);
nor U18781 (N_18781,N_17249,N_16336);
and U18782 (N_18782,N_16562,N_16310);
or U18783 (N_18783,N_16595,N_16234);
and U18784 (N_18784,N_17920,N_17701);
or U18785 (N_18785,N_16042,N_16859);
or U18786 (N_18786,N_16253,N_17746);
nor U18787 (N_18787,N_17783,N_17605);
and U18788 (N_18788,N_17902,N_17233);
or U18789 (N_18789,N_17424,N_16407);
xnor U18790 (N_18790,N_16456,N_17675);
nor U18791 (N_18791,N_16897,N_17228);
nand U18792 (N_18792,N_16514,N_16693);
or U18793 (N_18793,N_17586,N_16566);
xor U18794 (N_18794,N_16813,N_16463);
or U18795 (N_18795,N_17637,N_16735);
nor U18796 (N_18796,N_16291,N_17363);
or U18797 (N_18797,N_17215,N_16087);
nand U18798 (N_18798,N_17946,N_17458);
and U18799 (N_18799,N_16280,N_16511);
nor U18800 (N_18800,N_16920,N_17140);
and U18801 (N_18801,N_17741,N_16138);
and U18802 (N_18802,N_16349,N_17907);
nor U18803 (N_18803,N_16404,N_16299);
and U18804 (N_18804,N_17100,N_17271);
nor U18805 (N_18805,N_17110,N_16237);
nand U18806 (N_18806,N_16005,N_16858);
or U18807 (N_18807,N_16559,N_16255);
or U18808 (N_18808,N_16640,N_17725);
and U18809 (N_18809,N_17003,N_17176);
nor U18810 (N_18810,N_16096,N_17856);
nand U18811 (N_18811,N_16363,N_16534);
and U18812 (N_18812,N_16954,N_17617);
or U18813 (N_18813,N_17805,N_16453);
or U18814 (N_18814,N_17593,N_16142);
nand U18815 (N_18815,N_16141,N_17904);
or U18816 (N_18816,N_16338,N_16656);
nor U18817 (N_18817,N_17583,N_17244);
nand U18818 (N_18818,N_16847,N_16082);
nand U18819 (N_18819,N_17275,N_17597);
nand U18820 (N_18820,N_17041,N_16855);
and U18821 (N_18821,N_16317,N_17500);
nand U18822 (N_18822,N_17728,N_17785);
or U18823 (N_18823,N_16632,N_17009);
and U18824 (N_18824,N_17115,N_16586);
nand U18825 (N_18825,N_17955,N_16872);
nand U18826 (N_18826,N_17027,N_16986);
and U18827 (N_18827,N_17408,N_17388);
nand U18828 (N_18828,N_17656,N_16301);
nand U18829 (N_18829,N_16283,N_16584);
nor U18830 (N_18830,N_17188,N_17162);
xor U18831 (N_18831,N_17366,N_16672);
nor U18832 (N_18832,N_17382,N_17998);
or U18833 (N_18833,N_17064,N_17372);
and U18834 (N_18834,N_17695,N_17337);
nor U18835 (N_18835,N_16564,N_16563);
or U18836 (N_18836,N_17318,N_17196);
or U18837 (N_18837,N_16353,N_17843);
and U18838 (N_18838,N_16229,N_17979);
nor U18839 (N_18839,N_16364,N_16208);
and U18840 (N_18840,N_16429,N_16116);
or U18841 (N_18841,N_16295,N_16568);
nor U18842 (N_18842,N_16565,N_17237);
and U18843 (N_18843,N_16548,N_16403);
and U18844 (N_18844,N_16744,N_17896);
nand U18845 (N_18845,N_17831,N_17717);
nand U18846 (N_18846,N_16573,N_17910);
nor U18847 (N_18847,N_17361,N_17351);
nand U18848 (N_18848,N_17036,N_16839);
or U18849 (N_18849,N_16538,N_16808);
and U18850 (N_18850,N_17909,N_17663);
and U18851 (N_18851,N_16121,N_16482);
nand U18852 (N_18852,N_16187,N_16560);
nand U18853 (N_18853,N_17824,N_17183);
or U18854 (N_18854,N_17206,N_17835);
nor U18855 (N_18855,N_17392,N_17839);
and U18856 (N_18856,N_17808,N_17005);
nor U18857 (N_18857,N_17928,N_16505);
nand U18858 (N_18858,N_16522,N_16124);
and U18859 (N_18859,N_17582,N_16985);
nand U18860 (N_18860,N_17862,N_16919);
nand U18861 (N_18861,N_16206,N_16192);
nor U18862 (N_18862,N_16296,N_16312);
nand U18863 (N_18863,N_17968,N_17413);
or U18864 (N_18864,N_17903,N_16262);
or U18865 (N_18865,N_16103,N_16719);
nor U18866 (N_18866,N_17600,N_16936);
nand U18867 (N_18867,N_16271,N_16374);
xor U18868 (N_18868,N_17292,N_17255);
and U18869 (N_18869,N_17770,N_16030);
nor U18870 (N_18870,N_17730,N_17740);
nor U18871 (N_18871,N_16673,N_17628);
or U18872 (N_18872,N_16194,N_17006);
or U18873 (N_18873,N_16355,N_16340);
nand U18874 (N_18874,N_17985,N_17141);
and U18875 (N_18875,N_17784,N_16424);
and U18876 (N_18876,N_16263,N_17143);
and U18877 (N_18877,N_17315,N_17066);
and U18878 (N_18878,N_17261,N_16875);
nor U18879 (N_18879,N_16248,N_17875);
and U18880 (N_18880,N_17501,N_16512);
and U18881 (N_18881,N_16761,N_16742);
nor U18882 (N_18882,N_16130,N_16821);
nor U18883 (N_18883,N_16352,N_17470);
xor U18884 (N_18884,N_17166,N_17218);
nand U18885 (N_18885,N_17538,N_16545);
and U18886 (N_18886,N_16521,N_16956);
nand U18887 (N_18887,N_16256,N_16577);
nor U18888 (N_18888,N_17113,N_16475);
and U18889 (N_18889,N_16976,N_17683);
or U18890 (N_18890,N_16257,N_16250);
nor U18891 (N_18891,N_16477,N_16606);
nand U18892 (N_18892,N_16503,N_17310);
nor U18893 (N_18893,N_16376,N_17539);
nor U18894 (N_18894,N_17898,N_17776);
nor U18895 (N_18895,N_16645,N_17225);
or U18896 (N_18896,N_16027,N_16653);
and U18897 (N_18897,N_17174,N_17753);
and U18898 (N_18898,N_17766,N_17572);
nand U18899 (N_18899,N_17744,N_16112);
nand U18900 (N_18900,N_16743,N_16506);
nor U18901 (N_18901,N_17570,N_17098);
and U18902 (N_18902,N_16109,N_16059);
nand U18903 (N_18903,N_17025,N_17279);
nor U18904 (N_18904,N_16348,N_17028);
or U18905 (N_18905,N_17524,N_16529);
nand U18906 (N_18906,N_17852,N_17868);
and U18907 (N_18907,N_16297,N_16751);
and U18908 (N_18908,N_16490,N_17853);
nor U18909 (N_18909,N_17807,N_16033);
or U18910 (N_18910,N_16389,N_17945);
or U18911 (N_18911,N_17254,N_17724);
or U18912 (N_18912,N_16495,N_17045);
nor U18913 (N_18913,N_17314,N_16313);
and U18914 (N_18914,N_16736,N_17035);
nor U18915 (N_18915,N_17138,N_16982);
nand U18916 (N_18916,N_16202,N_16779);
or U18917 (N_18917,N_17116,N_17134);
nor U18918 (N_18918,N_17094,N_17182);
and U18919 (N_18919,N_16948,N_17893);
or U18920 (N_18920,N_17612,N_17131);
nor U18921 (N_18921,N_16814,N_16896);
nor U18922 (N_18922,N_16032,N_17561);
and U18923 (N_18923,N_17900,N_16236);
or U18924 (N_18924,N_17819,N_16691);
and U18925 (N_18925,N_16110,N_17778);
nor U18926 (N_18926,N_17929,N_16758);
and U18927 (N_18927,N_16180,N_16388);
nand U18928 (N_18928,N_16754,N_16054);
nand U18929 (N_18929,N_17641,N_16308);
nor U18930 (N_18930,N_17081,N_17452);
or U18931 (N_18931,N_17609,N_17792);
nand U18932 (N_18932,N_16880,N_17888);
or U18933 (N_18933,N_17940,N_17872);
and U18934 (N_18934,N_16520,N_17936);
and U18935 (N_18935,N_16964,N_16422);
and U18936 (N_18936,N_17548,N_17087);
nor U18937 (N_18937,N_17023,N_17352);
nand U18938 (N_18938,N_16199,N_16591);
or U18939 (N_18939,N_16667,N_17229);
nand U18940 (N_18940,N_16774,N_16323);
or U18941 (N_18941,N_17445,N_16797);
or U18942 (N_18942,N_17387,N_16539);
nand U18943 (N_18943,N_17711,N_16829);
or U18944 (N_18944,N_17323,N_16243);
or U18945 (N_18945,N_17662,N_16478);
nor U18946 (N_18946,N_17545,N_17973);
or U18947 (N_18947,N_16836,N_17329);
nor U18948 (N_18948,N_16873,N_16516);
or U18949 (N_18949,N_17471,N_17769);
nor U18950 (N_18950,N_17019,N_16228);
nor U18951 (N_18951,N_16837,N_16462);
nand U18952 (N_18952,N_17908,N_17358);
and U18953 (N_18953,N_16432,N_17691);
nor U18954 (N_18954,N_17082,N_16578);
or U18955 (N_18955,N_16739,N_16302);
nand U18956 (N_18956,N_16359,N_16405);
or U18957 (N_18957,N_17686,N_16418);
nor U18958 (N_18958,N_17010,N_16517);
or U18959 (N_18959,N_16784,N_16015);
or U18960 (N_18960,N_16690,N_16036);
nor U18961 (N_18961,N_16998,N_16848);
nand U18962 (N_18962,N_16675,N_16777);
nand U18963 (N_18963,N_16695,N_16160);
nor U18964 (N_18964,N_17954,N_16646);
or U18965 (N_18965,N_16101,N_16786);
nand U18966 (N_18966,N_16305,N_16601);
nor U18967 (N_18967,N_16700,N_16823);
nand U18968 (N_18968,N_16011,N_16611);
and U18969 (N_18969,N_17481,N_17816);
nor U18970 (N_18970,N_16311,N_17043);
nand U18971 (N_18971,N_17895,N_17001);
or U18972 (N_18972,N_17654,N_16546);
and U18973 (N_18973,N_16344,N_17268);
nor U18974 (N_18974,N_17962,N_16882);
or U18975 (N_18975,N_17963,N_16292);
or U18976 (N_18976,N_17130,N_17040);
and U18977 (N_18977,N_17669,N_17427);
xnor U18978 (N_18978,N_17886,N_17871);
nand U18979 (N_18979,N_16502,N_17782);
or U18980 (N_18980,N_17652,N_16484);
nand U18981 (N_18981,N_16906,N_16933);
or U18982 (N_18982,N_17014,N_17880);
nand U18983 (N_18983,N_16791,N_17276);
or U18984 (N_18984,N_17185,N_16351);
or U18985 (N_18985,N_17690,N_17266);
and U18986 (N_18986,N_17079,N_17270);
nand U18987 (N_18987,N_17838,N_16481);
and U18988 (N_18988,N_16625,N_17699);
or U18989 (N_18989,N_16907,N_17790);
nor U18990 (N_18990,N_17478,N_17487);
and U18991 (N_18991,N_17150,N_17034);
nor U18992 (N_18992,N_17114,N_17013);
nand U18993 (N_18993,N_16329,N_17610);
and U18994 (N_18994,N_17460,N_17590);
or U18995 (N_18995,N_17972,N_17715);
nand U18996 (N_18996,N_16108,N_16000);
nand U18997 (N_18997,N_16931,N_16900);
or U18998 (N_18998,N_17882,N_17584);
or U18999 (N_18999,N_17241,N_16260);
or U19000 (N_19000,N_17019,N_16740);
nand U19001 (N_19001,N_16834,N_17132);
and U19002 (N_19002,N_17014,N_16250);
and U19003 (N_19003,N_16283,N_17950);
nand U19004 (N_19004,N_17053,N_16236);
or U19005 (N_19005,N_17289,N_16556);
or U19006 (N_19006,N_17778,N_17492);
and U19007 (N_19007,N_16856,N_17347);
nor U19008 (N_19008,N_17534,N_16536);
or U19009 (N_19009,N_17851,N_16399);
nor U19010 (N_19010,N_17756,N_17791);
or U19011 (N_19011,N_16911,N_16617);
and U19012 (N_19012,N_17614,N_17172);
nor U19013 (N_19013,N_16029,N_17028);
nand U19014 (N_19014,N_16786,N_16496);
and U19015 (N_19015,N_16541,N_16184);
nor U19016 (N_19016,N_16127,N_17668);
nor U19017 (N_19017,N_17935,N_16114);
nand U19018 (N_19018,N_17852,N_16799);
nand U19019 (N_19019,N_17160,N_17048);
or U19020 (N_19020,N_17124,N_16832);
nand U19021 (N_19021,N_17996,N_17191);
or U19022 (N_19022,N_16446,N_16138);
or U19023 (N_19023,N_17982,N_17135);
nor U19024 (N_19024,N_16968,N_16219);
and U19025 (N_19025,N_16409,N_16101);
nor U19026 (N_19026,N_17549,N_16434);
nand U19027 (N_19027,N_17723,N_16523);
or U19028 (N_19028,N_16696,N_16800);
nand U19029 (N_19029,N_16482,N_16458);
or U19030 (N_19030,N_16081,N_16764);
or U19031 (N_19031,N_16262,N_17003);
nor U19032 (N_19032,N_16859,N_16566);
and U19033 (N_19033,N_17535,N_17336);
nand U19034 (N_19034,N_17647,N_17576);
or U19035 (N_19035,N_17529,N_17414);
and U19036 (N_19036,N_17664,N_17449);
or U19037 (N_19037,N_16872,N_17412);
nor U19038 (N_19038,N_17467,N_16640);
nor U19039 (N_19039,N_17745,N_17218);
or U19040 (N_19040,N_16812,N_16265);
nor U19041 (N_19041,N_16941,N_16211);
or U19042 (N_19042,N_17136,N_17503);
nand U19043 (N_19043,N_16538,N_17471);
nand U19044 (N_19044,N_17149,N_17215);
and U19045 (N_19045,N_16494,N_16207);
and U19046 (N_19046,N_16521,N_16434);
and U19047 (N_19047,N_16912,N_17923);
and U19048 (N_19048,N_17678,N_16727);
nand U19049 (N_19049,N_17067,N_17267);
or U19050 (N_19050,N_16302,N_16779);
or U19051 (N_19051,N_17415,N_16387);
and U19052 (N_19052,N_16879,N_17527);
nand U19053 (N_19053,N_17912,N_17793);
nand U19054 (N_19054,N_16146,N_16847);
nand U19055 (N_19055,N_17647,N_17723);
nor U19056 (N_19056,N_16723,N_17921);
or U19057 (N_19057,N_16783,N_17793);
or U19058 (N_19058,N_16866,N_17123);
nor U19059 (N_19059,N_17235,N_17029);
nor U19060 (N_19060,N_17912,N_16701);
or U19061 (N_19061,N_16787,N_16236);
nor U19062 (N_19062,N_16443,N_16161);
and U19063 (N_19063,N_16844,N_17022);
or U19064 (N_19064,N_16876,N_16689);
or U19065 (N_19065,N_17642,N_17224);
and U19066 (N_19066,N_17925,N_16902);
nand U19067 (N_19067,N_16408,N_16204);
nor U19068 (N_19068,N_16852,N_17415);
nor U19069 (N_19069,N_16691,N_16457);
nor U19070 (N_19070,N_16743,N_17496);
or U19071 (N_19071,N_16353,N_17949);
and U19072 (N_19072,N_17947,N_16324);
and U19073 (N_19073,N_16466,N_16149);
nand U19074 (N_19074,N_17814,N_17545);
or U19075 (N_19075,N_16575,N_17601);
xnor U19076 (N_19076,N_16280,N_16049);
nor U19077 (N_19077,N_17736,N_16189);
or U19078 (N_19078,N_17358,N_17877);
nand U19079 (N_19079,N_16709,N_16162);
or U19080 (N_19080,N_16482,N_16409);
and U19081 (N_19081,N_16606,N_16697);
nor U19082 (N_19082,N_17695,N_17022);
nand U19083 (N_19083,N_16681,N_17064);
nand U19084 (N_19084,N_17054,N_16008);
or U19085 (N_19085,N_16115,N_16138);
nand U19086 (N_19086,N_16139,N_17578);
or U19087 (N_19087,N_17132,N_16972);
and U19088 (N_19088,N_16214,N_16788);
nand U19089 (N_19089,N_17136,N_17684);
xor U19090 (N_19090,N_17064,N_17700);
nor U19091 (N_19091,N_16240,N_16791);
or U19092 (N_19092,N_17767,N_16944);
nor U19093 (N_19093,N_16340,N_17995);
and U19094 (N_19094,N_16619,N_16984);
nand U19095 (N_19095,N_17676,N_17010);
or U19096 (N_19096,N_17877,N_17166);
nor U19097 (N_19097,N_17185,N_17387);
nor U19098 (N_19098,N_17333,N_16156);
nor U19099 (N_19099,N_17620,N_17205);
nand U19100 (N_19100,N_17430,N_17754);
nor U19101 (N_19101,N_16045,N_16386);
or U19102 (N_19102,N_16054,N_17044);
nor U19103 (N_19103,N_16877,N_17499);
or U19104 (N_19104,N_16282,N_16916);
or U19105 (N_19105,N_17150,N_17709);
and U19106 (N_19106,N_16448,N_17352);
and U19107 (N_19107,N_16102,N_16972);
and U19108 (N_19108,N_17756,N_16574);
nand U19109 (N_19109,N_16129,N_17750);
and U19110 (N_19110,N_16683,N_17958);
or U19111 (N_19111,N_16600,N_16948);
nor U19112 (N_19112,N_17630,N_16923);
and U19113 (N_19113,N_16566,N_17158);
or U19114 (N_19114,N_17524,N_16933);
or U19115 (N_19115,N_17872,N_17432);
nor U19116 (N_19116,N_16769,N_16186);
xnor U19117 (N_19117,N_17183,N_17226);
and U19118 (N_19118,N_16345,N_17052);
and U19119 (N_19119,N_16349,N_17929);
nor U19120 (N_19120,N_16382,N_16658);
nor U19121 (N_19121,N_17259,N_17438);
nand U19122 (N_19122,N_17236,N_17985);
or U19123 (N_19123,N_16833,N_16682);
nor U19124 (N_19124,N_17306,N_16287);
and U19125 (N_19125,N_16342,N_16341);
and U19126 (N_19126,N_17904,N_17618);
or U19127 (N_19127,N_16820,N_17689);
and U19128 (N_19128,N_17430,N_17319);
nor U19129 (N_19129,N_17673,N_16797);
and U19130 (N_19130,N_16054,N_17500);
or U19131 (N_19131,N_16767,N_17162);
nor U19132 (N_19132,N_17785,N_16698);
or U19133 (N_19133,N_17309,N_17688);
and U19134 (N_19134,N_16552,N_17328);
nand U19135 (N_19135,N_16215,N_17898);
and U19136 (N_19136,N_17810,N_17229);
nor U19137 (N_19137,N_16536,N_16234);
nor U19138 (N_19138,N_16913,N_16980);
nand U19139 (N_19139,N_16895,N_17999);
nor U19140 (N_19140,N_16115,N_17656);
and U19141 (N_19141,N_17873,N_16121);
and U19142 (N_19142,N_16429,N_17266);
or U19143 (N_19143,N_16021,N_17719);
nor U19144 (N_19144,N_17924,N_17147);
nand U19145 (N_19145,N_16034,N_16820);
or U19146 (N_19146,N_16350,N_17079);
nand U19147 (N_19147,N_17253,N_17118);
nor U19148 (N_19148,N_16286,N_16436);
and U19149 (N_19149,N_16549,N_16758);
and U19150 (N_19150,N_17417,N_17760);
and U19151 (N_19151,N_16343,N_17422);
nand U19152 (N_19152,N_17260,N_17284);
and U19153 (N_19153,N_16008,N_16285);
nor U19154 (N_19154,N_17562,N_17604);
nor U19155 (N_19155,N_16769,N_16388);
and U19156 (N_19156,N_16542,N_17214);
and U19157 (N_19157,N_17166,N_17176);
xor U19158 (N_19158,N_16933,N_16664);
nor U19159 (N_19159,N_16265,N_16775);
or U19160 (N_19160,N_17431,N_16762);
and U19161 (N_19161,N_16453,N_16071);
nand U19162 (N_19162,N_17178,N_16409);
nor U19163 (N_19163,N_17163,N_16311);
nor U19164 (N_19164,N_17531,N_16086);
nor U19165 (N_19165,N_16105,N_17967);
nor U19166 (N_19166,N_17863,N_16065);
nor U19167 (N_19167,N_17000,N_17786);
nand U19168 (N_19168,N_17020,N_17545);
nor U19169 (N_19169,N_16727,N_16793);
nand U19170 (N_19170,N_16310,N_17723);
or U19171 (N_19171,N_17621,N_16903);
nand U19172 (N_19172,N_16918,N_16244);
nor U19173 (N_19173,N_17257,N_16135);
nor U19174 (N_19174,N_16501,N_17064);
nor U19175 (N_19175,N_16538,N_16081);
nand U19176 (N_19176,N_17308,N_16685);
or U19177 (N_19177,N_16979,N_17371);
and U19178 (N_19178,N_16009,N_17918);
and U19179 (N_19179,N_17163,N_16106);
or U19180 (N_19180,N_16048,N_16822);
nor U19181 (N_19181,N_17804,N_17889);
or U19182 (N_19182,N_16498,N_16244);
or U19183 (N_19183,N_17885,N_16774);
and U19184 (N_19184,N_16094,N_17688);
or U19185 (N_19185,N_17444,N_17411);
nor U19186 (N_19186,N_17587,N_16180);
nor U19187 (N_19187,N_16114,N_16375);
nor U19188 (N_19188,N_16953,N_16122);
nand U19189 (N_19189,N_17225,N_17627);
nand U19190 (N_19190,N_16003,N_16330);
nand U19191 (N_19191,N_16973,N_16172);
nand U19192 (N_19192,N_17749,N_16806);
and U19193 (N_19193,N_16945,N_17323);
and U19194 (N_19194,N_16729,N_16568);
and U19195 (N_19195,N_16137,N_17373);
nor U19196 (N_19196,N_16094,N_16995);
and U19197 (N_19197,N_16685,N_16944);
or U19198 (N_19198,N_17985,N_16530);
nor U19199 (N_19199,N_17640,N_17540);
or U19200 (N_19200,N_16957,N_17087);
nor U19201 (N_19201,N_17173,N_16534);
nand U19202 (N_19202,N_17336,N_16209);
nor U19203 (N_19203,N_17644,N_17335);
nand U19204 (N_19204,N_16758,N_16030);
and U19205 (N_19205,N_16159,N_16971);
or U19206 (N_19206,N_16086,N_17821);
nor U19207 (N_19207,N_17522,N_16027);
nor U19208 (N_19208,N_16693,N_16958);
nor U19209 (N_19209,N_16955,N_16377);
or U19210 (N_19210,N_16521,N_16605);
and U19211 (N_19211,N_16690,N_17922);
and U19212 (N_19212,N_16150,N_16556);
nor U19213 (N_19213,N_16179,N_16665);
or U19214 (N_19214,N_17166,N_17361);
nor U19215 (N_19215,N_17429,N_16905);
and U19216 (N_19216,N_17857,N_16259);
and U19217 (N_19217,N_16828,N_16856);
nand U19218 (N_19218,N_16806,N_17921);
and U19219 (N_19219,N_17069,N_17541);
or U19220 (N_19220,N_17343,N_17885);
nand U19221 (N_19221,N_16215,N_17376);
and U19222 (N_19222,N_17625,N_17052);
nor U19223 (N_19223,N_17672,N_16151);
nor U19224 (N_19224,N_16711,N_17806);
nor U19225 (N_19225,N_16901,N_17323);
nand U19226 (N_19226,N_17470,N_16254);
or U19227 (N_19227,N_16643,N_17381);
and U19228 (N_19228,N_17776,N_16616);
or U19229 (N_19229,N_16949,N_17746);
or U19230 (N_19230,N_16016,N_17967);
or U19231 (N_19231,N_16299,N_16463);
or U19232 (N_19232,N_17314,N_16646);
nor U19233 (N_19233,N_17886,N_17218);
or U19234 (N_19234,N_16948,N_16334);
nor U19235 (N_19235,N_16578,N_17222);
or U19236 (N_19236,N_16550,N_17589);
or U19237 (N_19237,N_17635,N_17095);
or U19238 (N_19238,N_16128,N_16704);
nor U19239 (N_19239,N_16559,N_16335);
or U19240 (N_19240,N_16661,N_17558);
nor U19241 (N_19241,N_17270,N_16188);
or U19242 (N_19242,N_16651,N_16601);
nand U19243 (N_19243,N_17642,N_16565);
nand U19244 (N_19244,N_17759,N_16538);
nand U19245 (N_19245,N_17165,N_16094);
nor U19246 (N_19246,N_17406,N_17164);
and U19247 (N_19247,N_17218,N_17834);
and U19248 (N_19248,N_17050,N_17271);
nor U19249 (N_19249,N_16721,N_17789);
and U19250 (N_19250,N_16764,N_17517);
nor U19251 (N_19251,N_16230,N_16102);
nand U19252 (N_19252,N_16545,N_16654);
nand U19253 (N_19253,N_17883,N_17823);
nand U19254 (N_19254,N_17411,N_17217);
and U19255 (N_19255,N_17950,N_17612);
nand U19256 (N_19256,N_17153,N_16987);
nor U19257 (N_19257,N_17475,N_16429);
nand U19258 (N_19258,N_17715,N_17554);
nor U19259 (N_19259,N_17377,N_17132);
or U19260 (N_19260,N_17955,N_17230);
nand U19261 (N_19261,N_16889,N_17636);
nand U19262 (N_19262,N_17858,N_16704);
nor U19263 (N_19263,N_16550,N_17044);
and U19264 (N_19264,N_17001,N_16917);
or U19265 (N_19265,N_16132,N_16296);
xor U19266 (N_19266,N_16498,N_17728);
and U19267 (N_19267,N_17198,N_17415);
or U19268 (N_19268,N_16893,N_16608);
nor U19269 (N_19269,N_16464,N_16729);
and U19270 (N_19270,N_16612,N_16290);
nand U19271 (N_19271,N_16265,N_16800);
or U19272 (N_19272,N_16766,N_16564);
or U19273 (N_19273,N_16726,N_16951);
and U19274 (N_19274,N_17411,N_17185);
nor U19275 (N_19275,N_16679,N_16887);
nor U19276 (N_19276,N_16815,N_16375);
nand U19277 (N_19277,N_16912,N_17105);
and U19278 (N_19278,N_16999,N_16580);
nor U19279 (N_19279,N_16319,N_17453);
or U19280 (N_19280,N_16657,N_17426);
nand U19281 (N_19281,N_16435,N_17301);
nor U19282 (N_19282,N_17065,N_16874);
and U19283 (N_19283,N_16372,N_17879);
xor U19284 (N_19284,N_16769,N_17534);
nand U19285 (N_19285,N_17274,N_16347);
or U19286 (N_19286,N_16020,N_16964);
nor U19287 (N_19287,N_16637,N_17436);
nand U19288 (N_19288,N_17905,N_17711);
or U19289 (N_19289,N_17309,N_16190);
or U19290 (N_19290,N_16530,N_16028);
and U19291 (N_19291,N_16618,N_17624);
nor U19292 (N_19292,N_16012,N_17738);
nor U19293 (N_19293,N_16367,N_16777);
nand U19294 (N_19294,N_16971,N_16870);
and U19295 (N_19295,N_17984,N_17673);
or U19296 (N_19296,N_17985,N_16725);
and U19297 (N_19297,N_17521,N_17159);
and U19298 (N_19298,N_17204,N_16724);
nand U19299 (N_19299,N_17095,N_16745);
and U19300 (N_19300,N_16069,N_17216);
nand U19301 (N_19301,N_17299,N_17632);
nor U19302 (N_19302,N_16357,N_16785);
and U19303 (N_19303,N_17565,N_16092);
or U19304 (N_19304,N_16215,N_16391);
and U19305 (N_19305,N_17265,N_16014);
and U19306 (N_19306,N_16331,N_17147);
nand U19307 (N_19307,N_17180,N_17800);
or U19308 (N_19308,N_16497,N_16722);
nor U19309 (N_19309,N_17473,N_16754);
and U19310 (N_19310,N_16424,N_16808);
or U19311 (N_19311,N_17278,N_17205);
nand U19312 (N_19312,N_16558,N_16419);
or U19313 (N_19313,N_16979,N_17283);
nand U19314 (N_19314,N_17976,N_17677);
nor U19315 (N_19315,N_16482,N_17281);
and U19316 (N_19316,N_17016,N_16498);
nand U19317 (N_19317,N_17768,N_16025);
nor U19318 (N_19318,N_17758,N_16663);
or U19319 (N_19319,N_16779,N_16298);
nor U19320 (N_19320,N_16717,N_16567);
nor U19321 (N_19321,N_16764,N_17091);
nor U19322 (N_19322,N_16962,N_16128);
or U19323 (N_19323,N_17156,N_17748);
nor U19324 (N_19324,N_17640,N_16110);
and U19325 (N_19325,N_16528,N_16212);
or U19326 (N_19326,N_16750,N_16924);
and U19327 (N_19327,N_16660,N_16970);
nand U19328 (N_19328,N_16224,N_16929);
nand U19329 (N_19329,N_17395,N_17103);
or U19330 (N_19330,N_16447,N_17437);
and U19331 (N_19331,N_16230,N_16158);
nand U19332 (N_19332,N_16240,N_16382);
or U19333 (N_19333,N_16764,N_17134);
nor U19334 (N_19334,N_16336,N_17269);
nor U19335 (N_19335,N_17670,N_17981);
or U19336 (N_19336,N_16354,N_17302);
nand U19337 (N_19337,N_16434,N_16815);
and U19338 (N_19338,N_16311,N_16611);
nand U19339 (N_19339,N_17166,N_17605);
nor U19340 (N_19340,N_17382,N_17072);
or U19341 (N_19341,N_16277,N_16403);
and U19342 (N_19342,N_16475,N_17412);
nand U19343 (N_19343,N_16714,N_16425);
and U19344 (N_19344,N_17650,N_16130);
nor U19345 (N_19345,N_17086,N_17534);
nor U19346 (N_19346,N_17256,N_16445);
nor U19347 (N_19347,N_16306,N_16714);
and U19348 (N_19348,N_17470,N_16553);
nor U19349 (N_19349,N_17363,N_17247);
nand U19350 (N_19350,N_16625,N_17280);
or U19351 (N_19351,N_16757,N_17782);
nand U19352 (N_19352,N_17981,N_17484);
or U19353 (N_19353,N_16454,N_17160);
nand U19354 (N_19354,N_17673,N_17878);
nand U19355 (N_19355,N_16013,N_16145);
and U19356 (N_19356,N_17180,N_16049);
nor U19357 (N_19357,N_16422,N_16556);
and U19358 (N_19358,N_17063,N_16232);
nor U19359 (N_19359,N_17062,N_17208);
nor U19360 (N_19360,N_16633,N_16022);
or U19361 (N_19361,N_17478,N_17632);
nand U19362 (N_19362,N_17379,N_17602);
nand U19363 (N_19363,N_16763,N_17669);
nand U19364 (N_19364,N_16833,N_16896);
nand U19365 (N_19365,N_17373,N_16555);
and U19366 (N_19366,N_16383,N_16607);
or U19367 (N_19367,N_16952,N_16632);
nor U19368 (N_19368,N_16440,N_17686);
nor U19369 (N_19369,N_17923,N_17878);
and U19370 (N_19370,N_16511,N_17371);
or U19371 (N_19371,N_17984,N_16612);
and U19372 (N_19372,N_17213,N_16854);
nor U19373 (N_19373,N_17993,N_17975);
nand U19374 (N_19374,N_17412,N_17538);
or U19375 (N_19375,N_16815,N_16737);
and U19376 (N_19376,N_16716,N_17516);
nor U19377 (N_19377,N_16118,N_17825);
nor U19378 (N_19378,N_16485,N_17811);
nor U19379 (N_19379,N_17724,N_16844);
and U19380 (N_19380,N_16318,N_16291);
and U19381 (N_19381,N_16630,N_17449);
or U19382 (N_19382,N_16753,N_16260);
and U19383 (N_19383,N_16791,N_16958);
and U19384 (N_19384,N_16963,N_16329);
nor U19385 (N_19385,N_16205,N_17756);
nand U19386 (N_19386,N_16441,N_17590);
nand U19387 (N_19387,N_16656,N_17543);
nor U19388 (N_19388,N_17926,N_16534);
nand U19389 (N_19389,N_17373,N_16227);
nand U19390 (N_19390,N_17895,N_17436);
nor U19391 (N_19391,N_16498,N_17369);
nor U19392 (N_19392,N_16475,N_17574);
or U19393 (N_19393,N_16193,N_16213);
nor U19394 (N_19394,N_16833,N_16184);
nor U19395 (N_19395,N_16840,N_16834);
and U19396 (N_19396,N_17116,N_17030);
nor U19397 (N_19397,N_17762,N_16357);
or U19398 (N_19398,N_17520,N_17480);
and U19399 (N_19399,N_17527,N_17163);
nand U19400 (N_19400,N_17047,N_17323);
or U19401 (N_19401,N_17303,N_16826);
and U19402 (N_19402,N_17600,N_17033);
or U19403 (N_19403,N_17799,N_16445);
nand U19404 (N_19404,N_17668,N_17892);
nor U19405 (N_19405,N_17132,N_16319);
nor U19406 (N_19406,N_16633,N_16867);
or U19407 (N_19407,N_16109,N_17157);
nor U19408 (N_19408,N_16178,N_16060);
nand U19409 (N_19409,N_17102,N_16403);
nand U19410 (N_19410,N_17757,N_17537);
nand U19411 (N_19411,N_17005,N_17972);
nor U19412 (N_19412,N_17084,N_17828);
nor U19413 (N_19413,N_17905,N_17104);
and U19414 (N_19414,N_17464,N_17462);
nor U19415 (N_19415,N_16138,N_17242);
nor U19416 (N_19416,N_16839,N_17388);
or U19417 (N_19417,N_17589,N_16268);
nor U19418 (N_19418,N_16460,N_16780);
and U19419 (N_19419,N_16157,N_16877);
or U19420 (N_19420,N_16524,N_16732);
nand U19421 (N_19421,N_16011,N_17906);
and U19422 (N_19422,N_17453,N_16042);
and U19423 (N_19423,N_16413,N_17978);
nor U19424 (N_19424,N_16572,N_17474);
nand U19425 (N_19425,N_17338,N_16539);
and U19426 (N_19426,N_16223,N_16738);
nand U19427 (N_19427,N_16938,N_17226);
and U19428 (N_19428,N_17246,N_16973);
nor U19429 (N_19429,N_17727,N_16807);
and U19430 (N_19430,N_17725,N_16438);
or U19431 (N_19431,N_17889,N_16564);
nor U19432 (N_19432,N_17208,N_17035);
nor U19433 (N_19433,N_16448,N_16014);
and U19434 (N_19434,N_17607,N_16993);
nor U19435 (N_19435,N_17880,N_17381);
nor U19436 (N_19436,N_16388,N_16751);
or U19437 (N_19437,N_17887,N_17851);
nand U19438 (N_19438,N_16163,N_17008);
nor U19439 (N_19439,N_16389,N_17438);
and U19440 (N_19440,N_17312,N_16086);
and U19441 (N_19441,N_17412,N_17462);
nor U19442 (N_19442,N_17924,N_17312);
nand U19443 (N_19443,N_16371,N_17567);
or U19444 (N_19444,N_17006,N_17026);
nor U19445 (N_19445,N_17083,N_17916);
nor U19446 (N_19446,N_17509,N_16372);
or U19447 (N_19447,N_16537,N_16371);
nor U19448 (N_19448,N_16476,N_16524);
nor U19449 (N_19449,N_16639,N_17802);
and U19450 (N_19450,N_16601,N_17397);
or U19451 (N_19451,N_16629,N_17659);
or U19452 (N_19452,N_16179,N_16899);
nand U19453 (N_19453,N_17535,N_16397);
and U19454 (N_19454,N_17363,N_16839);
nor U19455 (N_19455,N_16890,N_16411);
nor U19456 (N_19456,N_16825,N_17132);
and U19457 (N_19457,N_16988,N_17156);
xor U19458 (N_19458,N_16520,N_16969);
and U19459 (N_19459,N_17606,N_16250);
or U19460 (N_19460,N_17155,N_17380);
or U19461 (N_19461,N_17492,N_16935);
xor U19462 (N_19462,N_16948,N_17774);
or U19463 (N_19463,N_16640,N_16886);
nand U19464 (N_19464,N_17642,N_16751);
nand U19465 (N_19465,N_17152,N_17150);
nand U19466 (N_19466,N_16414,N_16578);
or U19467 (N_19467,N_16501,N_16410);
nor U19468 (N_19468,N_17649,N_16432);
or U19469 (N_19469,N_17829,N_16639);
nor U19470 (N_19470,N_16114,N_17509);
nand U19471 (N_19471,N_16823,N_17349);
and U19472 (N_19472,N_17097,N_16943);
nand U19473 (N_19473,N_16389,N_17769);
and U19474 (N_19474,N_16399,N_17731);
nand U19475 (N_19475,N_16384,N_17652);
or U19476 (N_19476,N_17871,N_16312);
and U19477 (N_19477,N_17441,N_17530);
nor U19478 (N_19478,N_17805,N_17676);
or U19479 (N_19479,N_16329,N_16812);
or U19480 (N_19480,N_16190,N_16639);
nand U19481 (N_19481,N_17011,N_17437);
or U19482 (N_19482,N_17216,N_17690);
nor U19483 (N_19483,N_16063,N_17253);
nor U19484 (N_19484,N_17474,N_16834);
nor U19485 (N_19485,N_17772,N_16797);
nor U19486 (N_19486,N_16670,N_16184);
or U19487 (N_19487,N_17582,N_16285);
and U19488 (N_19488,N_16690,N_16687);
nor U19489 (N_19489,N_17448,N_17498);
nor U19490 (N_19490,N_17157,N_16226);
nor U19491 (N_19491,N_16006,N_17598);
or U19492 (N_19492,N_16860,N_16178);
nand U19493 (N_19493,N_16775,N_16283);
and U19494 (N_19494,N_17330,N_16447);
or U19495 (N_19495,N_16438,N_16348);
nand U19496 (N_19496,N_16320,N_17446);
nor U19497 (N_19497,N_17412,N_17291);
nand U19498 (N_19498,N_16915,N_17587);
and U19499 (N_19499,N_16258,N_17854);
nand U19500 (N_19500,N_17638,N_17558);
nor U19501 (N_19501,N_17537,N_16992);
and U19502 (N_19502,N_16801,N_17486);
or U19503 (N_19503,N_17267,N_16433);
and U19504 (N_19504,N_17404,N_16782);
nor U19505 (N_19505,N_16409,N_16419);
or U19506 (N_19506,N_16987,N_17594);
nor U19507 (N_19507,N_16677,N_17356);
nor U19508 (N_19508,N_17579,N_16861);
or U19509 (N_19509,N_17595,N_16295);
and U19510 (N_19510,N_17892,N_16542);
or U19511 (N_19511,N_17553,N_17251);
or U19512 (N_19512,N_17512,N_16004);
and U19513 (N_19513,N_17178,N_17383);
and U19514 (N_19514,N_17214,N_17809);
and U19515 (N_19515,N_17528,N_16878);
and U19516 (N_19516,N_17660,N_17595);
or U19517 (N_19517,N_16037,N_16587);
nor U19518 (N_19518,N_17046,N_16680);
or U19519 (N_19519,N_17914,N_17896);
nor U19520 (N_19520,N_16890,N_17089);
or U19521 (N_19521,N_16915,N_17279);
and U19522 (N_19522,N_17698,N_17214);
nand U19523 (N_19523,N_16741,N_17932);
nor U19524 (N_19524,N_16554,N_16214);
nand U19525 (N_19525,N_17976,N_17924);
nor U19526 (N_19526,N_17061,N_17492);
or U19527 (N_19527,N_17966,N_17126);
nor U19528 (N_19528,N_17250,N_16520);
nor U19529 (N_19529,N_16345,N_17639);
nand U19530 (N_19530,N_16367,N_17319);
or U19531 (N_19531,N_16585,N_17016);
or U19532 (N_19532,N_16269,N_16457);
or U19533 (N_19533,N_16912,N_16656);
or U19534 (N_19534,N_16643,N_17281);
nor U19535 (N_19535,N_17483,N_17954);
nor U19536 (N_19536,N_17398,N_17658);
nand U19537 (N_19537,N_17705,N_17116);
nand U19538 (N_19538,N_16511,N_16283);
nor U19539 (N_19539,N_17602,N_16674);
nand U19540 (N_19540,N_17053,N_16660);
or U19541 (N_19541,N_16463,N_17859);
or U19542 (N_19542,N_17392,N_16155);
nand U19543 (N_19543,N_16279,N_17499);
nand U19544 (N_19544,N_17927,N_16088);
and U19545 (N_19545,N_17942,N_17830);
nand U19546 (N_19546,N_16780,N_17497);
or U19547 (N_19547,N_17693,N_16579);
and U19548 (N_19548,N_17929,N_17429);
or U19549 (N_19549,N_17623,N_17361);
nand U19550 (N_19550,N_16281,N_17593);
nor U19551 (N_19551,N_17594,N_17562);
or U19552 (N_19552,N_17937,N_17058);
nand U19553 (N_19553,N_17694,N_17055);
or U19554 (N_19554,N_16115,N_17803);
and U19555 (N_19555,N_16647,N_16557);
nand U19556 (N_19556,N_17347,N_16858);
and U19557 (N_19557,N_16686,N_17219);
nand U19558 (N_19558,N_17131,N_16146);
nor U19559 (N_19559,N_16234,N_16192);
nor U19560 (N_19560,N_16477,N_17750);
nand U19561 (N_19561,N_16909,N_16873);
nor U19562 (N_19562,N_17463,N_17609);
nor U19563 (N_19563,N_17881,N_16539);
nand U19564 (N_19564,N_17456,N_17373);
nor U19565 (N_19565,N_17030,N_16198);
and U19566 (N_19566,N_16896,N_17658);
nor U19567 (N_19567,N_17446,N_16693);
nor U19568 (N_19568,N_16682,N_16766);
nor U19569 (N_19569,N_17300,N_17830);
nor U19570 (N_19570,N_16106,N_17683);
nor U19571 (N_19571,N_16666,N_17536);
nand U19572 (N_19572,N_16292,N_17105);
and U19573 (N_19573,N_16656,N_17840);
nand U19574 (N_19574,N_17014,N_16754);
nand U19575 (N_19575,N_17679,N_17571);
nor U19576 (N_19576,N_17673,N_16686);
or U19577 (N_19577,N_16570,N_16985);
nand U19578 (N_19578,N_16978,N_17152);
nor U19579 (N_19579,N_16807,N_16749);
and U19580 (N_19580,N_16220,N_17962);
nor U19581 (N_19581,N_17112,N_16461);
nand U19582 (N_19582,N_16254,N_16761);
nor U19583 (N_19583,N_17257,N_17822);
or U19584 (N_19584,N_16088,N_16217);
or U19585 (N_19585,N_16254,N_16932);
nand U19586 (N_19586,N_16305,N_16186);
nor U19587 (N_19587,N_17117,N_16913);
and U19588 (N_19588,N_17821,N_16231);
or U19589 (N_19589,N_16661,N_16492);
nor U19590 (N_19590,N_17658,N_16120);
and U19591 (N_19591,N_16541,N_17534);
nor U19592 (N_19592,N_17378,N_17308);
and U19593 (N_19593,N_16438,N_17372);
nor U19594 (N_19594,N_16937,N_17782);
or U19595 (N_19595,N_17601,N_17425);
nor U19596 (N_19596,N_16304,N_17491);
and U19597 (N_19597,N_16650,N_17738);
or U19598 (N_19598,N_16089,N_16217);
and U19599 (N_19599,N_16076,N_16703);
and U19600 (N_19600,N_17572,N_16510);
nor U19601 (N_19601,N_16547,N_17772);
nand U19602 (N_19602,N_17485,N_16661);
nor U19603 (N_19603,N_17488,N_17300);
nand U19604 (N_19604,N_17153,N_16507);
nand U19605 (N_19605,N_17398,N_17005);
and U19606 (N_19606,N_16266,N_16009);
or U19607 (N_19607,N_16416,N_16116);
nor U19608 (N_19608,N_17871,N_17894);
nor U19609 (N_19609,N_17971,N_17947);
or U19610 (N_19610,N_17969,N_17367);
nor U19611 (N_19611,N_17612,N_16196);
and U19612 (N_19612,N_16990,N_17102);
nand U19613 (N_19613,N_16498,N_17224);
and U19614 (N_19614,N_17748,N_17136);
nand U19615 (N_19615,N_16414,N_16349);
nand U19616 (N_19616,N_17127,N_16057);
and U19617 (N_19617,N_16111,N_17870);
nand U19618 (N_19618,N_16377,N_16171);
nor U19619 (N_19619,N_16055,N_17811);
nand U19620 (N_19620,N_17912,N_17611);
nor U19621 (N_19621,N_17172,N_16945);
nand U19622 (N_19622,N_16958,N_16186);
or U19623 (N_19623,N_17191,N_16870);
and U19624 (N_19624,N_17622,N_16362);
and U19625 (N_19625,N_17594,N_16999);
nor U19626 (N_19626,N_16410,N_16522);
nor U19627 (N_19627,N_17515,N_16906);
and U19628 (N_19628,N_16216,N_16907);
nand U19629 (N_19629,N_17955,N_16111);
and U19630 (N_19630,N_17352,N_16500);
nor U19631 (N_19631,N_16228,N_17816);
nand U19632 (N_19632,N_16513,N_16972);
xnor U19633 (N_19633,N_16103,N_16311);
or U19634 (N_19634,N_17077,N_17836);
or U19635 (N_19635,N_17038,N_16705);
nor U19636 (N_19636,N_16946,N_16927);
nand U19637 (N_19637,N_16885,N_17993);
nor U19638 (N_19638,N_17821,N_16334);
nand U19639 (N_19639,N_17464,N_16650);
nand U19640 (N_19640,N_17088,N_17097);
nand U19641 (N_19641,N_16269,N_17103);
nand U19642 (N_19642,N_17166,N_17429);
and U19643 (N_19643,N_17419,N_16215);
nand U19644 (N_19644,N_16208,N_17844);
nand U19645 (N_19645,N_16086,N_17333);
nor U19646 (N_19646,N_16043,N_17803);
or U19647 (N_19647,N_16553,N_16622);
nand U19648 (N_19648,N_16930,N_17869);
nor U19649 (N_19649,N_17724,N_16070);
nor U19650 (N_19650,N_17263,N_16878);
nor U19651 (N_19651,N_17929,N_16767);
or U19652 (N_19652,N_17724,N_16422);
or U19653 (N_19653,N_16443,N_17959);
and U19654 (N_19654,N_16996,N_16903);
and U19655 (N_19655,N_16137,N_17786);
nor U19656 (N_19656,N_16527,N_16812);
and U19657 (N_19657,N_16581,N_17171);
or U19658 (N_19658,N_17663,N_17837);
and U19659 (N_19659,N_17582,N_16414);
and U19660 (N_19660,N_17684,N_16368);
and U19661 (N_19661,N_16138,N_17669);
and U19662 (N_19662,N_16481,N_16769);
nor U19663 (N_19663,N_17531,N_17919);
nand U19664 (N_19664,N_16352,N_17094);
nand U19665 (N_19665,N_16029,N_16617);
nor U19666 (N_19666,N_16358,N_16804);
nand U19667 (N_19667,N_17921,N_17966);
nor U19668 (N_19668,N_17002,N_17976);
and U19669 (N_19669,N_16459,N_16687);
and U19670 (N_19670,N_16998,N_16001);
and U19671 (N_19671,N_17757,N_16344);
and U19672 (N_19672,N_16556,N_16919);
xnor U19673 (N_19673,N_16320,N_17058);
nor U19674 (N_19674,N_17422,N_17837);
nand U19675 (N_19675,N_16603,N_17875);
or U19676 (N_19676,N_17790,N_17727);
nor U19677 (N_19677,N_16268,N_16730);
and U19678 (N_19678,N_16356,N_16037);
nor U19679 (N_19679,N_17162,N_17841);
nor U19680 (N_19680,N_16244,N_17440);
nor U19681 (N_19681,N_16194,N_17071);
and U19682 (N_19682,N_16321,N_16295);
or U19683 (N_19683,N_17467,N_17436);
nand U19684 (N_19684,N_17535,N_16209);
or U19685 (N_19685,N_17831,N_16473);
nor U19686 (N_19686,N_16125,N_16139);
and U19687 (N_19687,N_17075,N_17345);
or U19688 (N_19688,N_17972,N_17673);
or U19689 (N_19689,N_17875,N_17858);
nor U19690 (N_19690,N_16423,N_16269);
nand U19691 (N_19691,N_16901,N_17370);
nor U19692 (N_19692,N_16221,N_16965);
nor U19693 (N_19693,N_17980,N_17303);
nor U19694 (N_19694,N_16322,N_17236);
nand U19695 (N_19695,N_16911,N_16258);
nand U19696 (N_19696,N_17766,N_17914);
nor U19697 (N_19697,N_17348,N_16792);
nor U19698 (N_19698,N_17408,N_17474);
nand U19699 (N_19699,N_17934,N_16814);
nor U19700 (N_19700,N_17413,N_17240);
nor U19701 (N_19701,N_16990,N_17418);
and U19702 (N_19702,N_17800,N_16171);
nand U19703 (N_19703,N_17507,N_16657);
nor U19704 (N_19704,N_16173,N_16752);
and U19705 (N_19705,N_17455,N_16832);
nor U19706 (N_19706,N_16518,N_16654);
nand U19707 (N_19707,N_16901,N_16375);
and U19708 (N_19708,N_16214,N_17818);
and U19709 (N_19709,N_17258,N_16493);
nor U19710 (N_19710,N_17972,N_16676);
nor U19711 (N_19711,N_16058,N_16721);
or U19712 (N_19712,N_17477,N_17759);
nor U19713 (N_19713,N_16897,N_16155);
nor U19714 (N_19714,N_17354,N_17249);
or U19715 (N_19715,N_17876,N_16772);
nor U19716 (N_19716,N_16990,N_16926);
nor U19717 (N_19717,N_16074,N_16578);
and U19718 (N_19718,N_17461,N_16852);
nand U19719 (N_19719,N_16203,N_17829);
or U19720 (N_19720,N_17344,N_16227);
or U19721 (N_19721,N_17361,N_16636);
nand U19722 (N_19722,N_17096,N_17115);
nand U19723 (N_19723,N_17979,N_16719);
or U19724 (N_19724,N_17257,N_16837);
and U19725 (N_19725,N_16327,N_17823);
and U19726 (N_19726,N_17179,N_17346);
and U19727 (N_19727,N_16333,N_17746);
nand U19728 (N_19728,N_16867,N_16888);
or U19729 (N_19729,N_16376,N_17287);
nand U19730 (N_19730,N_17048,N_17960);
nor U19731 (N_19731,N_17873,N_16857);
xnor U19732 (N_19732,N_16534,N_17248);
and U19733 (N_19733,N_17906,N_16644);
or U19734 (N_19734,N_16080,N_17247);
nor U19735 (N_19735,N_16258,N_16577);
or U19736 (N_19736,N_17621,N_17623);
nand U19737 (N_19737,N_16624,N_16205);
or U19738 (N_19738,N_16276,N_16006);
or U19739 (N_19739,N_16398,N_17528);
or U19740 (N_19740,N_16787,N_17374);
or U19741 (N_19741,N_17307,N_16019);
or U19742 (N_19742,N_16225,N_17427);
and U19743 (N_19743,N_16807,N_17817);
and U19744 (N_19744,N_17280,N_17621);
or U19745 (N_19745,N_17406,N_16951);
and U19746 (N_19746,N_16817,N_17122);
and U19747 (N_19747,N_17977,N_16432);
nand U19748 (N_19748,N_17112,N_17803);
or U19749 (N_19749,N_17512,N_16332);
nor U19750 (N_19750,N_17982,N_17966);
nor U19751 (N_19751,N_17463,N_17743);
nor U19752 (N_19752,N_16090,N_16980);
nand U19753 (N_19753,N_17558,N_16359);
nand U19754 (N_19754,N_17660,N_17884);
nor U19755 (N_19755,N_16274,N_16021);
nand U19756 (N_19756,N_16492,N_16377);
nor U19757 (N_19757,N_16927,N_16752);
or U19758 (N_19758,N_16793,N_16924);
nand U19759 (N_19759,N_16894,N_16856);
nand U19760 (N_19760,N_16350,N_16896);
nor U19761 (N_19761,N_16875,N_16860);
or U19762 (N_19762,N_16898,N_16249);
nor U19763 (N_19763,N_17566,N_16139);
and U19764 (N_19764,N_17099,N_16095);
nor U19765 (N_19765,N_16792,N_17481);
or U19766 (N_19766,N_17433,N_17531);
nand U19767 (N_19767,N_17795,N_17872);
nand U19768 (N_19768,N_17901,N_17710);
or U19769 (N_19769,N_17423,N_17033);
or U19770 (N_19770,N_16049,N_16862);
or U19771 (N_19771,N_17559,N_16784);
nor U19772 (N_19772,N_16842,N_16229);
nor U19773 (N_19773,N_16349,N_17320);
nor U19774 (N_19774,N_16786,N_16315);
nand U19775 (N_19775,N_16841,N_17692);
nand U19776 (N_19776,N_16564,N_17185);
or U19777 (N_19777,N_16441,N_16252);
nand U19778 (N_19778,N_17524,N_16860);
or U19779 (N_19779,N_16026,N_16749);
or U19780 (N_19780,N_17165,N_16374);
and U19781 (N_19781,N_16007,N_17935);
or U19782 (N_19782,N_17960,N_16955);
nand U19783 (N_19783,N_17672,N_16062);
and U19784 (N_19784,N_16530,N_17821);
or U19785 (N_19785,N_16373,N_16841);
nand U19786 (N_19786,N_16097,N_16996);
or U19787 (N_19787,N_17837,N_16187);
nand U19788 (N_19788,N_16382,N_17314);
nand U19789 (N_19789,N_16343,N_17640);
and U19790 (N_19790,N_16779,N_17421);
nand U19791 (N_19791,N_17418,N_16170);
and U19792 (N_19792,N_16383,N_16988);
and U19793 (N_19793,N_17191,N_16540);
xor U19794 (N_19794,N_17390,N_17630);
nor U19795 (N_19795,N_16662,N_17128);
and U19796 (N_19796,N_16605,N_16820);
or U19797 (N_19797,N_17134,N_17420);
xnor U19798 (N_19798,N_17167,N_17747);
or U19799 (N_19799,N_17691,N_17710);
or U19800 (N_19800,N_16732,N_16084);
nand U19801 (N_19801,N_17003,N_16063);
nand U19802 (N_19802,N_17027,N_16143);
and U19803 (N_19803,N_17504,N_17296);
and U19804 (N_19804,N_17629,N_17557);
or U19805 (N_19805,N_16049,N_17023);
or U19806 (N_19806,N_16767,N_17417);
nand U19807 (N_19807,N_17988,N_16195);
and U19808 (N_19808,N_17791,N_16839);
and U19809 (N_19809,N_16187,N_17521);
nand U19810 (N_19810,N_16298,N_17041);
and U19811 (N_19811,N_17104,N_16361);
or U19812 (N_19812,N_16480,N_17236);
and U19813 (N_19813,N_16351,N_16592);
or U19814 (N_19814,N_17730,N_16732);
or U19815 (N_19815,N_16697,N_16934);
nor U19816 (N_19816,N_16731,N_17973);
nor U19817 (N_19817,N_17929,N_16055);
nand U19818 (N_19818,N_17231,N_17739);
nor U19819 (N_19819,N_16729,N_17761);
and U19820 (N_19820,N_17256,N_17239);
or U19821 (N_19821,N_17400,N_16191);
nor U19822 (N_19822,N_16557,N_17293);
or U19823 (N_19823,N_17966,N_16837);
nor U19824 (N_19824,N_16460,N_16005);
nor U19825 (N_19825,N_16385,N_17219);
and U19826 (N_19826,N_17762,N_17975);
nor U19827 (N_19827,N_17947,N_16134);
and U19828 (N_19828,N_17046,N_17144);
nand U19829 (N_19829,N_17382,N_16771);
or U19830 (N_19830,N_17518,N_16387);
or U19831 (N_19831,N_16081,N_16575);
or U19832 (N_19832,N_17810,N_17768);
or U19833 (N_19833,N_17711,N_17801);
nor U19834 (N_19834,N_16466,N_16573);
or U19835 (N_19835,N_16179,N_16096);
or U19836 (N_19836,N_17654,N_17409);
and U19837 (N_19837,N_16865,N_16973);
nor U19838 (N_19838,N_17563,N_17118);
nor U19839 (N_19839,N_16073,N_17974);
nor U19840 (N_19840,N_16453,N_17923);
or U19841 (N_19841,N_16450,N_17620);
or U19842 (N_19842,N_16074,N_16809);
nor U19843 (N_19843,N_17048,N_16992);
or U19844 (N_19844,N_17799,N_17503);
xor U19845 (N_19845,N_16021,N_17358);
nand U19846 (N_19846,N_16683,N_16474);
nand U19847 (N_19847,N_17524,N_16936);
and U19848 (N_19848,N_16658,N_16664);
nor U19849 (N_19849,N_16982,N_16882);
nor U19850 (N_19850,N_17088,N_17490);
nand U19851 (N_19851,N_17934,N_17146);
nor U19852 (N_19852,N_17400,N_17332);
or U19853 (N_19853,N_17672,N_16845);
or U19854 (N_19854,N_17146,N_17211);
and U19855 (N_19855,N_17843,N_17800);
nor U19856 (N_19856,N_16598,N_16158);
or U19857 (N_19857,N_17308,N_17561);
or U19858 (N_19858,N_16839,N_16049);
or U19859 (N_19859,N_16967,N_16439);
nand U19860 (N_19860,N_16525,N_16603);
or U19861 (N_19861,N_16739,N_16853);
nor U19862 (N_19862,N_17469,N_16027);
xor U19863 (N_19863,N_16308,N_17369);
and U19864 (N_19864,N_17773,N_16228);
nor U19865 (N_19865,N_16142,N_17947);
or U19866 (N_19866,N_16005,N_16986);
nand U19867 (N_19867,N_17318,N_16028);
nor U19868 (N_19868,N_16442,N_17572);
nand U19869 (N_19869,N_17182,N_17501);
and U19870 (N_19870,N_17075,N_16783);
nand U19871 (N_19871,N_17597,N_16793);
and U19872 (N_19872,N_16562,N_17491);
nor U19873 (N_19873,N_17993,N_16490);
or U19874 (N_19874,N_16412,N_16676);
xnor U19875 (N_19875,N_16545,N_17766);
or U19876 (N_19876,N_16380,N_16424);
or U19877 (N_19877,N_16189,N_17056);
or U19878 (N_19878,N_17936,N_17533);
or U19879 (N_19879,N_16704,N_16258);
nor U19880 (N_19880,N_17620,N_16169);
nand U19881 (N_19881,N_16767,N_17987);
or U19882 (N_19882,N_17482,N_16454);
and U19883 (N_19883,N_16717,N_17774);
or U19884 (N_19884,N_17982,N_17997);
nor U19885 (N_19885,N_17382,N_17178);
nor U19886 (N_19886,N_16580,N_16604);
nand U19887 (N_19887,N_17784,N_16111);
and U19888 (N_19888,N_17456,N_16992);
nand U19889 (N_19889,N_17105,N_17534);
nor U19890 (N_19890,N_17737,N_16088);
or U19891 (N_19891,N_17111,N_16594);
nand U19892 (N_19892,N_17309,N_17563);
or U19893 (N_19893,N_17980,N_16972);
nor U19894 (N_19894,N_16941,N_17853);
and U19895 (N_19895,N_16532,N_17435);
or U19896 (N_19896,N_17287,N_17676);
nor U19897 (N_19897,N_16685,N_16447);
nor U19898 (N_19898,N_16779,N_16413);
nand U19899 (N_19899,N_17705,N_16080);
nor U19900 (N_19900,N_16280,N_17819);
and U19901 (N_19901,N_17591,N_17798);
and U19902 (N_19902,N_16428,N_16371);
nand U19903 (N_19903,N_17869,N_16082);
nor U19904 (N_19904,N_17514,N_16495);
nor U19905 (N_19905,N_17963,N_16718);
and U19906 (N_19906,N_16099,N_16807);
and U19907 (N_19907,N_17451,N_16250);
nand U19908 (N_19908,N_16649,N_16441);
or U19909 (N_19909,N_16343,N_17363);
nand U19910 (N_19910,N_16270,N_17276);
nand U19911 (N_19911,N_17965,N_17652);
nor U19912 (N_19912,N_16802,N_17246);
nand U19913 (N_19913,N_17026,N_17381);
and U19914 (N_19914,N_17719,N_17099);
and U19915 (N_19915,N_17877,N_16050);
or U19916 (N_19916,N_16930,N_16849);
and U19917 (N_19917,N_16434,N_17089);
and U19918 (N_19918,N_17857,N_16659);
nand U19919 (N_19919,N_17191,N_16647);
nor U19920 (N_19920,N_16468,N_16006);
and U19921 (N_19921,N_16527,N_16019);
nand U19922 (N_19922,N_16422,N_16826);
nand U19923 (N_19923,N_17256,N_17995);
or U19924 (N_19924,N_17874,N_17047);
nor U19925 (N_19925,N_17910,N_17036);
nor U19926 (N_19926,N_17360,N_16301);
nand U19927 (N_19927,N_16920,N_16941);
and U19928 (N_19928,N_16479,N_16348);
or U19929 (N_19929,N_17609,N_17058);
nor U19930 (N_19930,N_17335,N_17337);
or U19931 (N_19931,N_16417,N_16392);
nand U19932 (N_19932,N_17831,N_16270);
nor U19933 (N_19933,N_17823,N_16766);
or U19934 (N_19934,N_16475,N_16246);
nand U19935 (N_19935,N_17566,N_17779);
nand U19936 (N_19936,N_17346,N_17196);
and U19937 (N_19937,N_17909,N_17046);
nand U19938 (N_19938,N_16531,N_17970);
nand U19939 (N_19939,N_16836,N_17061);
and U19940 (N_19940,N_16494,N_16223);
nor U19941 (N_19941,N_16828,N_16312);
nor U19942 (N_19942,N_16225,N_17265);
and U19943 (N_19943,N_17036,N_17690);
nor U19944 (N_19944,N_17793,N_16476);
nand U19945 (N_19945,N_17726,N_17237);
nand U19946 (N_19946,N_16458,N_16710);
nor U19947 (N_19947,N_17279,N_16524);
or U19948 (N_19948,N_16561,N_16735);
nand U19949 (N_19949,N_16484,N_16692);
nor U19950 (N_19950,N_16892,N_17375);
nor U19951 (N_19951,N_16085,N_17638);
or U19952 (N_19952,N_17009,N_16096);
and U19953 (N_19953,N_17944,N_17683);
and U19954 (N_19954,N_16844,N_17845);
or U19955 (N_19955,N_17533,N_16538);
nand U19956 (N_19956,N_17839,N_17824);
or U19957 (N_19957,N_17448,N_17923);
nand U19958 (N_19958,N_16024,N_16506);
nand U19959 (N_19959,N_17380,N_17576);
or U19960 (N_19960,N_16896,N_17411);
nand U19961 (N_19961,N_16663,N_16759);
nand U19962 (N_19962,N_16998,N_16331);
or U19963 (N_19963,N_16686,N_17970);
and U19964 (N_19964,N_17601,N_16749);
and U19965 (N_19965,N_17279,N_16012);
nor U19966 (N_19966,N_16569,N_17889);
or U19967 (N_19967,N_17540,N_17007);
or U19968 (N_19968,N_17825,N_16183);
nand U19969 (N_19969,N_16878,N_16485);
nor U19970 (N_19970,N_17762,N_16852);
and U19971 (N_19971,N_17656,N_17947);
and U19972 (N_19972,N_16741,N_16491);
or U19973 (N_19973,N_17418,N_17893);
or U19974 (N_19974,N_17560,N_17652);
or U19975 (N_19975,N_16184,N_16030);
or U19976 (N_19976,N_16215,N_16715);
nand U19977 (N_19977,N_16425,N_16076);
nor U19978 (N_19978,N_16679,N_16051);
nor U19979 (N_19979,N_17162,N_17632);
nor U19980 (N_19980,N_16778,N_16262);
or U19981 (N_19981,N_16653,N_16304);
and U19982 (N_19982,N_17210,N_17820);
or U19983 (N_19983,N_17171,N_17981);
and U19984 (N_19984,N_16950,N_16044);
and U19985 (N_19985,N_16008,N_16979);
nor U19986 (N_19986,N_17708,N_16081);
xnor U19987 (N_19987,N_16560,N_17280);
and U19988 (N_19988,N_17518,N_16050);
or U19989 (N_19989,N_16577,N_17543);
or U19990 (N_19990,N_16791,N_17656);
or U19991 (N_19991,N_16173,N_17210);
or U19992 (N_19992,N_16601,N_16537);
nand U19993 (N_19993,N_16076,N_17256);
and U19994 (N_19994,N_17199,N_17300);
and U19995 (N_19995,N_16739,N_16162);
or U19996 (N_19996,N_16400,N_16784);
nor U19997 (N_19997,N_16086,N_16942);
and U19998 (N_19998,N_16879,N_17037);
nor U19999 (N_19999,N_16698,N_17356);
or UO_0 (O_0,N_18220,N_18054);
nand UO_1 (O_1,N_19617,N_19260);
nand UO_2 (O_2,N_19993,N_18911);
nand UO_3 (O_3,N_18764,N_18274);
and UO_4 (O_4,N_19490,N_18730);
nand UO_5 (O_5,N_18494,N_18272);
or UO_6 (O_6,N_19436,N_19270);
nor UO_7 (O_7,N_19949,N_19195);
xor UO_8 (O_8,N_19284,N_19457);
and UO_9 (O_9,N_19155,N_18466);
nand UO_10 (O_10,N_19146,N_18292);
nor UO_11 (O_11,N_18543,N_18290);
nor UO_12 (O_12,N_18090,N_18035);
nand UO_13 (O_13,N_18161,N_19468);
and UO_14 (O_14,N_19899,N_18021);
or UO_15 (O_15,N_18676,N_19249);
nor UO_16 (O_16,N_18752,N_18571);
or UO_17 (O_17,N_19593,N_19778);
nor UO_18 (O_18,N_18209,N_19888);
and UO_19 (O_19,N_19362,N_18414);
nand UO_20 (O_20,N_18333,N_18694);
nor UO_21 (O_21,N_18348,N_18903);
or UO_22 (O_22,N_18082,N_19137);
or UO_23 (O_23,N_18648,N_18278);
and UO_24 (O_24,N_18187,N_18406);
nand UO_25 (O_25,N_19030,N_19838);
nand UO_26 (O_26,N_19883,N_19737);
nand UO_27 (O_27,N_19843,N_18975);
nor UO_28 (O_28,N_18664,N_18905);
nor UO_29 (O_29,N_19859,N_18792);
nand UO_30 (O_30,N_19753,N_18569);
xnor UO_31 (O_31,N_18644,N_19234);
nor UO_32 (O_32,N_19781,N_19629);
nor UO_33 (O_33,N_19412,N_19558);
or UO_34 (O_34,N_18800,N_19595);
nor UO_35 (O_35,N_18986,N_18769);
nand UO_36 (O_36,N_18554,N_19580);
nand UO_37 (O_37,N_19610,N_18103);
or UO_38 (O_38,N_19547,N_18207);
nor UO_39 (O_39,N_19369,N_19489);
nor UO_40 (O_40,N_18915,N_19719);
or UO_41 (O_41,N_18176,N_19214);
or UO_42 (O_42,N_18407,N_19563);
nor UO_43 (O_43,N_18255,N_18450);
or UO_44 (O_44,N_19349,N_19212);
or UO_45 (O_45,N_18024,N_19245);
nand UO_46 (O_46,N_18447,N_18020);
or UO_47 (O_47,N_19980,N_19114);
nor UO_48 (O_48,N_18839,N_18650);
or UO_49 (O_49,N_19674,N_19101);
nor UO_50 (O_50,N_19108,N_18072);
nor UO_51 (O_51,N_18258,N_18230);
nand UO_52 (O_52,N_18948,N_19743);
nand UO_53 (O_53,N_19879,N_18962);
nor UO_54 (O_54,N_18504,N_19091);
nand UO_55 (O_55,N_19045,N_18717);
nand UO_56 (O_56,N_18436,N_19426);
nor UO_57 (O_57,N_19598,N_19587);
nor UO_58 (O_58,N_18076,N_19764);
nor UO_59 (O_59,N_19543,N_18894);
or UO_60 (O_60,N_18555,N_18022);
or UO_61 (O_61,N_19707,N_18496);
and UO_62 (O_62,N_18749,N_18789);
nand UO_63 (O_63,N_18618,N_19898);
nand UO_64 (O_64,N_19196,N_19606);
nand UO_65 (O_65,N_19005,N_18095);
and UO_66 (O_66,N_18111,N_18830);
nand UO_67 (O_67,N_19867,N_19261);
or UO_68 (O_68,N_18308,N_18089);
and UO_69 (O_69,N_18900,N_18426);
or UO_70 (O_70,N_18475,N_19521);
or UO_71 (O_71,N_18287,N_18126);
nor UO_72 (O_72,N_19575,N_19130);
nor UO_73 (O_73,N_19067,N_18096);
and UO_74 (O_74,N_18509,N_18334);
nor UO_75 (O_75,N_18390,N_18378);
nand UO_76 (O_76,N_19433,N_19740);
nand UO_77 (O_77,N_19589,N_18886);
or UO_78 (O_78,N_18237,N_18429);
nand UO_79 (O_79,N_19493,N_19483);
or UO_80 (O_80,N_18271,N_19535);
nor UO_81 (O_81,N_18633,N_19300);
and UO_82 (O_82,N_18979,N_18640);
nor UO_83 (O_83,N_18027,N_18377);
nand UO_84 (O_84,N_18758,N_18615);
nor UO_85 (O_85,N_18007,N_18978);
and UO_86 (O_86,N_19806,N_18097);
and UO_87 (O_87,N_19757,N_19443);
or UO_88 (O_88,N_18208,N_19561);
nand UO_89 (O_89,N_18083,N_18533);
nor UO_90 (O_90,N_19076,N_19359);
or UO_91 (O_91,N_19789,N_18731);
and UO_92 (O_92,N_19160,N_19938);
nor UO_93 (O_93,N_19240,N_18195);
or UO_94 (O_94,N_18155,N_19276);
nand UO_95 (O_95,N_18701,N_18695);
and UO_96 (O_96,N_18798,N_19969);
and UO_97 (O_97,N_19511,N_18753);
and UO_98 (O_98,N_19275,N_19111);
or UO_99 (O_99,N_18037,N_18815);
nor UO_100 (O_100,N_19239,N_18924);
nor UO_101 (O_101,N_18844,N_19134);
nor UO_102 (O_102,N_18065,N_18771);
nand UO_103 (O_103,N_19669,N_19766);
nor UO_104 (O_104,N_18040,N_19927);
nor UO_105 (O_105,N_18128,N_19402);
nor UO_106 (O_106,N_19504,N_19001);
and UO_107 (O_107,N_18530,N_18358);
and UO_108 (O_108,N_18608,N_18046);
and UO_109 (O_109,N_19675,N_19180);
or UO_110 (O_110,N_18658,N_18060);
and UO_111 (O_111,N_19183,N_19166);
or UO_112 (O_112,N_19352,N_18478);
xnor UO_113 (O_113,N_18712,N_18225);
and UO_114 (O_114,N_19409,N_19152);
nand UO_115 (O_115,N_18952,N_19731);
and UO_116 (O_116,N_19250,N_18561);
nor UO_117 (O_117,N_19615,N_19386);
nand UO_118 (O_118,N_19653,N_19399);
nor UO_119 (O_119,N_18628,N_18235);
nor UO_120 (O_120,N_19200,N_18708);
nand UO_121 (O_121,N_18976,N_18122);
or UO_122 (O_122,N_19600,N_19799);
or UO_123 (O_123,N_18025,N_19122);
nor UO_124 (O_124,N_18394,N_19031);
nor UO_125 (O_125,N_19807,N_19325);
nand UO_126 (O_126,N_19253,N_19816);
nand UO_127 (O_127,N_18464,N_19159);
and UO_128 (O_128,N_18188,N_18245);
or UO_129 (O_129,N_19937,N_19657);
and UO_130 (O_130,N_19824,N_18068);
or UO_131 (O_131,N_19623,N_18073);
nand UO_132 (O_132,N_19424,N_19952);
and UO_133 (O_133,N_19024,N_18654);
and UO_134 (O_134,N_18874,N_18502);
nand UO_135 (O_135,N_19988,N_19312);
or UO_136 (O_136,N_18514,N_19939);
nor UO_137 (O_137,N_19501,N_18484);
nor UO_138 (O_138,N_19194,N_18688);
and UO_139 (O_139,N_18802,N_19099);
or UO_140 (O_140,N_19230,N_19186);
or UO_141 (O_141,N_18809,N_19765);
nor UO_142 (O_142,N_18148,N_19004);
nand UO_143 (O_143,N_18433,N_18101);
or UO_144 (O_144,N_18617,N_18227);
nand UO_145 (O_145,N_18768,N_18357);
and UO_146 (O_146,N_18444,N_19803);
nand UO_147 (O_147,N_18310,N_18567);
nor UO_148 (O_148,N_19118,N_19836);
and UO_149 (O_149,N_19225,N_18870);
or UO_150 (O_150,N_19204,N_18989);
or UO_151 (O_151,N_19699,N_19831);
and UO_152 (O_152,N_18120,N_19832);
or UO_153 (O_153,N_19692,N_19188);
and UO_154 (O_154,N_19073,N_18283);
or UO_155 (O_155,N_19301,N_19257);
nor UO_156 (O_156,N_18158,N_19112);
and UO_157 (O_157,N_18140,N_19242);
nand UO_158 (O_158,N_19711,N_19410);
or UO_159 (O_159,N_18596,N_19338);
and UO_160 (O_160,N_19631,N_18323);
or UO_161 (O_161,N_19648,N_18931);
xor UO_162 (O_162,N_18663,N_18277);
or UO_163 (O_163,N_19519,N_19174);
nand UO_164 (O_164,N_18189,N_18067);
and UO_165 (O_165,N_18675,N_18626);
and UO_166 (O_166,N_18636,N_18716);
nand UO_167 (O_167,N_18006,N_18869);
and UO_168 (O_168,N_18733,N_19794);
nor UO_169 (O_169,N_18198,N_19738);
nor UO_170 (O_170,N_18984,N_19599);
nand UO_171 (O_171,N_19448,N_18767);
and UO_172 (O_172,N_19259,N_19704);
xnor UO_173 (O_173,N_19298,N_18920);
and UO_174 (O_174,N_18536,N_18354);
and UO_175 (O_175,N_19425,N_19787);
or UO_176 (O_176,N_19470,N_19968);
nor UO_177 (O_177,N_19834,N_18346);
nand UO_178 (O_178,N_19583,N_19302);
or UO_179 (O_179,N_19461,N_19353);
nand UO_180 (O_180,N_19957,N_18091);
or UO_181 (O_181,N_19741,N_19213);
or UO_182 (O_182,N_19569,N_19100);
and UO_183 (O_183,N_18570,N_19603);
and UO_184 (O_184,N_19014,N_18835);
and UO_185 (O_185,N_19221,N_18385);
nor UO_186 (O_186,N_18641,N_18461);
nand UO_187 (O_187,N_19782,N_18216);
and UO_188 (O_188,N_19742,N_18755);
nand UO_189 (O_189,N_19286,N_19337);
and UO_190 (O_190,N_19248,N_18568);
or UO_191 (O_191,N_18019,N_18938);
nor UO_192 (O_192,N_18699,N_18481);
and UO_193 (O_193,N_19321,N_18551);
nor UO_194 (O_194,N_19280,N_19796);
and UO_195 (O_195,N_18489,N_18736);
nor UO_196 (O_196,N_18029,N_18453);
and UO_197 (O_197,N_18834,N_19320);
or UO_198 (O_198,N_18797,N_18234);
nand UO_199 (O_199,N_19793,N_18142);
or UO_200 (O_200,N_19418,N_18888);
nor UO_201 (O_201,N_18921,N_18412);
nor UO_202 (O_202,N_19153,N_18832);
nor UO_203 (O_203,N_19562,N_18868);
nand UO_204 (O_204,N_19560,N_19851);
or UO_205 (O_205,N_18030,N_19494);
nor UO_206 (O_206,N_18857,N_19954);
nand UO_207 (O_207,N_18313,N_18044);
or UO_208 (O_208,N_18579,N_19012);
nand UO_209 (O_209,N_18270,N_19528);
or UO_210 (O_210,N_18179,N_18949);
nand UO_211 (O_211,N_19708,N_19313);
nand UO_212 (O_212,N_19078,N_18693);
xor UO_213 (O_213,N_19517,N_19299);
and UO_214 (O_214,N_18192,N_19849);
and UO_215 (O_215,N_19278,N_19523);
or UO_216 (O_216,N_19139,N_19770);
and UO_217 (O_217,N_19785,N_18614);
and UO_218 (O_218,N_18885,N_19140);
nand UO_219 (O_219,N_19744,N_18325);
and UO_220 (O_220,N_18572,N_18933);
or UO_221 (O_221,N_19809,N_18154);
and UO_222 (O_222,N_18697,N_18244);
and UO_223 (O_223,N_19009,N_18837);
nor UO_224 (O_224,N_18167,N_18132);
or UO_225 (O_225,N_18081,N_19058);
nor UO_226 (O_226,N_18175,N_18350);
nand UO_227 (O_227,N_18670,N_19043);
nor UO_228 (O_228,N_18599,N_18214);
and UO_229 (O_229,N_19979,N_18652);
nand UO_230 (O_230,N_18744,N_18039);
nor UO_231 (O_231,N_18819,N_19181);
and UO_232 (O_232,N_19686,N_19752);
and UO_233 (O_233,N_19942,N_19021);
and UO_234 (O_234,N_18200,N_18770);
nand UO_235 (O_235,N_18973,N_18371);
and UO_236 (O_236,N_19854,N_19158);
and UO_237 (O_237,N_18144,N_19324);
nand UO_238 (O_238,N_19706,N_19419);
nor UO_239 (O_239,N_19071,N_19823);
nand UO_240 (O_240,N_19364,N_19978);
and UO_241 (O_241,N_18739,N_19668);
nand UO_242 (O_242,N_18413,N_18253);
or UO_243 (O_243,N_19694,N_19019);
or UO_244 (O_244,N_19633,N_19912);
nand UO_245 (O_245,N_18776,N_18704);
nor UO_246 (O_246,N_19946,N_19310);
and UO_247 (O_247,N_19437,N_19863);
nor UO_248 (O_248,N_19061,N_18314);
nor UO_249 (O_249,N_19087,N_18416);
or UO_250 (O_250,N_19034,N_18539);
nand UO_251 (O_251,N_18318,N_18910);
nand UO_252 (O_252,N_18965,N_18009);
or UO_253 (O_253,N_18129,N_19420);
or UO_254 (O_254,N_18836,N_19681);
nor UO_255 (O_255,N_19102,N_18124);
or UO_256 (O_256,N_19373,N_19844);
nand UO_257 (O_257,N_18164,N_19228);
or UO_258 (O_258,N_18026,N_18468);
or UO_259 (O_259,N_19607,N_19590);
or UO_260 (O_260,N_19294,N_18069);
and UO_261 (O_261,N_19372,N_18756);
or UO_262 (O_262,N_19736,N_19360);
and UO_263 (O_263,N_19878,N_19231);
and UO_264 (O_264,N_18174,N_18742);
nor UO_265 (O_265,N_18598,N_19588);
nor UO_266 (O_266,N_19476,N_18791);
nor UO_267 (O_267,N_18722,N_19289);
or UO_268 (O_268,N_19366,N_18880);
or UO_269 (O_269,N_18840,N_19222);
and UO_270 (O_270,N_19840,N_19281);
or UO_271 (O_271,N_18642,N_19170);
nand UO_272 (O_272,N_18719,N_19219);
nor UO_273 (O_273,N_18765,N_19572);
and UO_274 (O_274,N_18721,N_18172);
nand UO_275 (O_275,N_18462,N_19351);
and UO_276 (O_276,N_18557,N_19758);
nand UO_277 (O_277,N_19893,N_18532);
and UO_278 (O_278,N_18204,N_18223);
or UO_279 (O_279,N_19965,N_19077);
nor UO_280 (O_280,N_18391,N_19855);
and UO_281 (O_281,N_18517,N_18623);
and UO_282 (O_282,N_18259,N_19698);
nor UO_283 (O_283,N_19379,N_19406);
nor UO_284 (O_284,N_19304,N_18143);
nor UO_285 (O_285,N_19574,N_19747);
nor UO_286 (O_286,N_18224,N_18312);
nor UO_287 (O_287,N_19044,N_19544);
nand UO_288 (O_288,N_19917,N_18488);
nor UO_289 (O_289,N_18993,N_18233);
nand UO_290 (O_290,N_18330,N_18058);
nand UO_291 (O_291,N_18353,N_18610);
xnor UO_292 (O_292,N_18715,N_18469);
nand UO_293 (O_293,N_18268,N_19897);
nand UO_294 (O_294,N_18510,N_19396);
nor UO_295 (O_295,N_18594,N_19125);
nand UO_296 (O_296,N_18790,N_19862);
nor UO_297 (O_297,N_18275,N_19346);
nor UO_298 (O_298,N_19962,N_19924);
nor UO_299 (O_299,N_18612,N_18838);
nand UO_300 (O_300,N_19522,N_18783);
and UO_301 (O_301,N_19632,N_18854);
nand UO_302 (O_302,N_19955,N_18711);
and UO_303 (O_303,N_18041,N_18580);
nor UO_304 (O_304,N_19236,N_18092);
nand UO_305 (O_305,N_18045,N_18477);
nand UO_306 (O_306,N_18084,N_18063);
and UO_307 (O_307,N_19238,N_19546);
or UO_308 (O_308,N_19390,N_19693);
nor UO_309 (O_309,N_18546,N_19444);
nor UO_310 (O_310,N_18858,N_19217);
nor UO_311 (O_311,N_19171,N_18306);
and UO_312 (O_312,N_19054,N_18702);
or UO_313 (O_313,N_18607,N_18589);
and UO_314 (O_314,N_19847,N_19964);
or UO_315 (O_315,N_19833,N_19381);
nand UO_316 (O_316,N_19644,N_19918);
nor UO_317 (O_317,N_18899,N_18364);
or UO_318 (O_318,N_19496,N_18252);
nand UO_319 (O_319,N_19625,N_18898);
and UO_320 (O_320,N_18811,N_19997);
and UO_321 (O_321,N_19913,N_19143);
nand UO_322 (O_322,N_18941,N_19734);
and UO_323 (O_323,N_18890,N_19869);
or UO_324 (O_324,N_18162,N_19357);
nand UO_325 (O_325,N_18801,N_19901);
xor UO_326 (O_326,N_18653,N_18199);
nand UO_327 (O_327,N_18600,N_18743);
or UO_328 (O_328,N_18822,N_18309);
nand UO_329 (O_329,N_18232,N_19582);
nor UO_330 (O_330,N_18821,N_18945);
nor UO_331 (O_331,N_18028,N_18070);
nor UO_332 (O_332,N_19790,N_18947);
and UO_333 (O_333,N_18181,N_18635);
or UO_334 (O_334,N_18804,N_19876);
or UO_335 (O_335,N_19064,N_18441);
nor UO_336 (O_336,N_18262,N_19145);
nor UO_337 (O_337,N_18139,N_19010);
and UO_338 (O_338,N_19075,N_19920);
nor UO_339 (O_339,N_19841,N_19374);
or UO_340 (O_340,N_18171,N_19788);
and UO_341 (O_341,N_18341,N_19777);
or UO_342 (O_342,N_18520,N_19481);
and UO_343 (O_343,N_19113,N_18709);
nor UO_344 (O_344,N_18297,N_19646);
nor UO_345 (O_345,N_18566,N_18298);
and UO_346 (O_346,N_19350,N_19340);
or UO_347 (O_347,N_19970,N_18427);
and UO_348 (O_348,N_18643,N_18659);
nor UO_349 (O_349,N_19398,N_18231);
nor UO_350 (O_350,N_18656,N_18320);
or UO_351 (O_351,N_19786,N_19184);
or UO_352 (O_352,N_19571,N_19028);
nor UO_353 (O_353,N_18166,N_19342);
nor UO_354 (O_354,N_18891,N_19297);
and UO_355 (O_355,N_19126,N_19578);
nand UO_356 (O_356,N_18729,N_19116);
nor UO_357 (O_357,N_18328,N_19296);
nor UO_358 (O_358,N_18808,N_19667);
nor UO_359 (O_359,N_19601,N_19269);
nand UO_360 (O_360,N_19972,N_18690);
nor UO_361 (O_361,N_19209,N_19133);
or UO_362 (O_362,N_19232,N_18827);
and UO_363 (O_363,N_18226,N_19207);
nand UO_364 (O_364,N_19857,N_19515);
or UO_365 (O_365,N_18861,N_18928);
nand UO_366 (O_366,N_18786,N_18008);
and UO_367 (O_367,N_18707,N_19910);
nor UO_368 (O_368,N_19254,N_19464);
or UO_369 (O_369,N_18360,N_18877);
nand UO_370 (O_370,N_18518,N_19531);
nand UO_371 (O_371,N_18585,N_18700);
or UO_372 (O_372,N_19713,N_19439);
and UO_373 (O_373,N_19241,N_19775);
or UO_374 (O_374,N_18182,N_19487);
and UO_375 (O_375,N_18655,N_18398);
and UO_376 (O_376,N_19718,N_19192);
or UO_377 (O_377,N_18121,N_18823);
and UO_378 (O_378,N_19672,N_19772);
nor UO_379 (O_379,N_19035,N_19328);
nor UO_380 (O_380,N_19650,N_19554);
and UO_381 (O_381,N_18355,N_19107);
nand UO_382 (O_382,N_19990,N_19512);
nand UO_383 (O_383,N_18785,N_19908);
or UO_384 (O_384,N_19680,N_19656);
nand UO_385 (O_385,N_18105,N_18119);
nand UO_386 (O_386,N_19485,N_19976);
and UO_387 (O_387,N_19800,N_19482);
or UO_388 (O_388,N_19120,N_18556);
nor UO_389 (O_389,N_18750,N_18904);
or UO_390 (O_390,N_19921,N_18066);
nor UO_391 (O_391,N_18526,N_19048);
and UO_392 (O_392,N_19397,N_18490);
and UO_393 (O_393,N_19203,N_19144);
nor UO_394 (O_394,N_18582,N_19210);
and UO_395 (O_395,N_19268,N_19720);
or UO_396 (O_396,N_19592,N_18833);
nand UO_397 (O_397,N_19056,N_18423);
or UO_398 (O_398,N_19311,N_19709);
or UO_399 (O_399,N_19080,N_19760);
or UO_400 (O_400,N_18493,N_19380);
nand UO_401 (O_401,N_19916,N_19771);
and UO_402 (O_402,N_18500,N_19919);
nor UO_403 (O_403,N_18540,N_18956);
nand UO_404 (O_404,N_19395,N_18452);
nor UO_405 (O_405,N_19848,N_18524);
nor UO_406 (O_406,N_19597,N_19830);
and UO_407 (O_407,N_18738,N_19115);
nand UO_408 (O_408,N_18686,N_19127);
or UO_409 (O_409,N_18601,N_19336);
nand UO_410 (O_410,N_18110,N_19996);
nor UO_411 (O_411,N_19053,N_18813);
nor UO_412 (O_412,N_18828,N_19620);
and UO_413 (O_413,N_19341,N_19285);
nor UO_414 (O_414,N_19769,N_19432);
nor UO_415 (O_415,N_19252,N_19895);
nand UO_416 (O_416,N_18957,N_18657);
nor UO_417 (O_417,N_19040,N_18351);
nand UO_418 (O_418,N_19287,N_18997);
and UO_419 (O_419,N_18806,N_18296);
nand UO_420 (O_420,N_18408,N_18389);
or UO_421 (O_421,N_19948,N_18780);
nand UO_422 (O_422,N_18852,N_19573);
and UO_423 (O_423,N_19323,N_18146);
nand UO_424 (O_424,N_19052,N_19147);
and UO_425 (O_425,N_18817,N_18616);
xnor UO_426 (O_426,N_19027,N_19363);
nand UO_427 (O_427,N_18672,N_18471);
nor UO_428 (O_428,N_18332,N_19128);
or UO_429 (O_429,N_19923,N_18547);
nand UO_430 (O_430,N_18459,N_18677);
and UO_431 (O_431,N_18415,N_19393);
or UO_432 (O_432,N_18660,N_18953);
and UO_433 (O_433,N_18735,N_19084);
and UO_434 (O_434,N_19815,N_19002);
nand UO_435 (O_435,N_19985,N_18998);
nand UO_436 (O_436,N_19940,N_18882);
nand UO_437 (O_437,N_18723,N_18807);
nor UO_438 (O_438,N_18482,N_18562);
nand UO_439 (O_439,N_18191,N_18922);
nand UO_440 (O_440,N_18508,N_18432);
and UO_441 (O_441,N_18402,N_19375);
and UO_442 (O_442,N_18159,N_18917);
or UO_443 (O_443,N_19092,N_19331);
nor UO_444 (O_444,N_18160,N_18049);
nand UO_445 (O_445,N_18387,N_18681);
and UO_446 (O_446,N_19717,N_19703);
and UO_447 (O_447,N_19530,N_19157);
or UO_448 (O_448,N_19953,N_18212);
nor UO_449 (O_449,N_19628,N_18682);
nor UO_450 (O_450,N_19664,N_18734);
nor UO_451 (O_451,N_19688,N_18574);
nand UO_452 (O_452,N_18846,N_18291);
nand UO_453 (O_453,N_19036,N_19479);
nand UO_454 (O_454,N_19638,N_18609);
nor UO_455 (O_455,N_18583,N_19471);
nor UO_456 (O_456,N_19727,N_18971);
or UO_457 (O_457,N_19508,N_19626);
nor UO_458 (O_458,N_18288,N_18692);
or UO_459 (O_459,N_18392,N_18624);
nor UO_460 (O_460,N_18269,N_18201);
or UO_461 (O_461,N_19958,N_18247);
or UO_462 (O_462,N_18706,N_19665);
or UO_463 (O_463,N_19977,N_18909);
or UO_464 (O_464,N_19215,N_18362);
nor UO_465 (O_465,N_18077,N_18449);
nand UO_466 (O_466,N_18985,N_18714);
nor UO_467 (O_467,N_18679,N_19585);
nor UO_468 (O_468,N_18620,N_18629);
and UO_469 (O_469,N_19173,N_18125);
or UO_470 (O_470,N_19472,N_19509);
nand UO_471 (O_471,N_19000,N_18032);
nor UO_472 (O_472,N_19649,N_18982);
and UO_473 (O_473,N_18281,N_19728);
nor UO_474 (O_474,N_18958,N_19498);
and UO_475 (O_475,N_18454,N_18563);
nand UO_476 (O_476,N_19557,N_18969);
nor UO_477 (O_477,N_19208,N_19179);
nand UO_478 (O_478,N_19473,N_18505);
nor UO_479 (O_479,N_18728,N_19733);
nor UO_480 (O_480,N_18553,N_19712);
nand UO_481 (O_481,N_19885,N_19525);
or UO_482 (O_482,N_18936,N_18503);
nor UO_483 (O_483,N_19235,N_19550);
and UO_484 (O_484,N_18862,N_18180);
and UO_485 (O_485,N_19609,N_18229);
and UO_486 (O_486,N_18831,N_19982);
nand UO_487 (O_487,N_19466,N_19394);
nand UO_488 (O_488,N_18279,N_19037);
or UO_489 (O_489,N_18578,N_19696);
nand UO_490 (O_490,N_18380,N_19746);
or UO_491 (O_491,N_18375,N_19376);
nor UO_492 (O_492,N_18646,N_19683);
nor UO_493 (O_493,N_18919,N_19148);
nor UO_494 (O_494,N_19928,N_18523);
nor UO_495 (O_495,N_18254,N_18473);
or UO_496 (O_496,N_19066,N_18537);
nor UO_497 (O_497,N_18747,N_19416);
nand UO_498 (O_498,N_19507,N_18001);
nand UO_499 (O_499,N_18366,N_19678);
nand UO_500 (O_500,N_19537,N_19347);
and UO_501 (O_501,N_19400,N_18303);
nor UO_502 (O_502,N_18135,N_19538);
nor UO_503 (O_503,N_19427,N_19172);
and UO_504 (O_504,N_18050,N_18930);
nor UO_505 (O_505,N_18990,N_18376);
nor UO_506 (O_506,N_19630,N_18282);
or UO_507 (O_507,N_18052,N_19513);
nand UO_508 (O_508,N_18538,N_19199);
or UO_509 (O_509,N_18240,N_19821);
or UO_510 (O_510,N_18987,N_18873);
nand UO_511 (O_511,N_19552,N_19621);
nand UO_512 (O_512,N_19936,N_18343);
nand UO_513 (O_513,N_18038,N_18875);
nand UO_514 (O_514,N_19165,N_18053);
nand UO_515 (O_515,N_18178,N_18826);
nand UO_516 (O_516,N_18430,N_19011);
nor UO_517 (O_517,N_18942,N_19616);
nor UO_518 (O_518,N_19637,N_18867);
and UO_519 (O_519,N_18311,N_19963);
and UO_520 (O_520,N_18818,N_18528);
nand UO_521 (O_521,N_19845,N_18777);
nand UO_522 (O_522,N_18465,N_19032);
xnor UO_523 (O_523,N_19103,N_18929);
nor UO_524 (O_524,N_19860,N_19176);
and UO_525 (O_525,N_19059,N_19505);
nand UO_526 (O_526,N_19865,N_18703);
nor UO_527 (O_527,N_18883,N_19808);
nor UO_528 (O_528,N_18859,N_18411);
and UO_529 (O_529,N_18115,N_19246);
or UO_530 (O_530,N_19423,N_19907);
nor UO_531 (O_531,N_19542,N_19697);
or UO_532 (O_532,N_18264,N_19334);
and UO_533 (O_533,N_18943,N_18324);
and UO_534 (O_534,N_18944,N_18860);
and UO_535 (O_535,N_18959,N_19455);
nand UO_536 (O_536,N_18257,N_18338);
and UO_537 (O_537,N_19377,N_18327);
and UO_538 (O_538,N_18062,N_19008);
nand UO_539 (O_539,N_18866,N_19460);
nand UO_540 (O_540,N_19226,N_19877);
and UO_541 (O_541,N_19383,N_19541);
nand UO_542 (O_542,N_19905,N_18276);
nor UO_543 (O_543,N_18593,N_18141);
nor UO_544 (O_544,N_19817,N_18256);
or UO_545 (O_545,N_18273,N_19875);
nand UO_546 (O_546,N_18855,N_19023);
or UO_547 (O_547,N_19534,N_18535);
or UO_548 (O_548,N_18075,N_19013);
or UO_549 (O_549,N_19438,N_18645);
or UO_550 (O_550,N_19109,N_18955);
or UO_551 (O_551,N_19317,N_18145);
or UO_552 (O_552,N_18544,N_19434);
nand UO_553 (O_553,N_19654,N_19797);
or UO_554 (O_554,N_18960,N_19445);
and UO_555 (O_555,N_18856,N_19477);
and UO_556 (O_556,N_18964,N_18577);
or UO_557 (O_557,N_19567,N_18302);
nor UO_558 (O_558,N_19435,N_18410);
nand UO_559 (O_559,N_18995,N_19085);
nor UO_560 (O_560,N_18138,N_18051);
and UO_561 (O_561,N_19273,N_19882);
nand UO_562 (O_562,N_18991,N_18116);
or UO_563 (O_563,N_18285,N_18057);
nand UO_564 (O_564,N_18033,N_19887);
nand UO_565 (O_565,N_18590,N_18106);
and UO_566 (O_566,N_19858,N_18974);
or UO_567 (O_567,N_18056,N_19647);
or UO_568 (O_568,N_18250,N_19068);
and UO_569 (O_569,N_19072,N_19701);
and UO_570 (O_570,N_19062,N_19783);
or UO_571 (O_571,N_19943,N_19658);
nor UO_572 (O_572,N_19536,N_19033);
nor UO_573 (O_573,N_18206,N_19651);
nor UO_574 (O_574,N_19258,N_19662);
or UO_575 (O_575,N_19202,N_19442);
or UO_576 (O_576,N_19608,N_18136);
nand UO_577 (O_577,N_18887,N_19526);
nand UO_578 (O_578,N_18381,N_19614);
and UO_579 (O_579,N_19553,N_19729);
nor UO_580 (O_580,N_18017,N_18151);
xor UO_581 (O_581,N_18977,N_18434);
nor UO_582 (O_582,N_18266,N_19243);
and UO_583 (O_583,N_18102,N_18428);
nand UO_584 (O_584,N_18299,N_18242);
or UO_585 (O_585,N_18061,N_19057);
nor UO_586 (O_586,N_18527,N_18483);
or UO_587 (O_587,N_19149,N_18871);
nor UO_588 (O_588,N_18638,N_19828);
nor UO_589 (O_589,N_18671,N_19178);
or UO_590 (O_590,N_19763,N_18079);
and UO_591 (O_591,N_18451,N_19387);
or UO_592 (O_592,N_19211,N_18395);
nand UO_593 (O_593,N_18016,N_19762);
and UO_594 (O_594,N_19685,N_18374);
or UO_595 (O_595,N_18190,N_19135);
nor UO_596 (O_596,N_18901,N_18349);
nand UO_597 (O_597,N_18134,N_18668);
or UO_598 (O_598,N_18074,N_19999);
and UO_599 (O_599,N_19343,N_18511);
or UO_600 (O_600,N_19038,N_19779);
or UO_601 (O_601,N_18501,N_18994);
and UO_602 (O_602,N_19695,N_19655);
nor UO_603 (O_603,N_19306,N_18284);
and UO_604 (O_604,N_19190,N_18611);
or UO_605 (O_605,N_18368,N_19288);
nor UO_606 (O_606,N_19132,N_19813);
or UO_607 (O_607,N_19348,N_18713);
nand UO_608 (O_608,N_19974,N_18382);
and UO_609 (O_609,N_18521,N_19532);
xor UO_610 (O_610,N_18512,N_19322);
and UO_611 (O_611,N_19776,N_19440);
nand UO_612 (O_612,N_19539,N_18999);
nand UO_613 (O_613,N_19182,N_19689);
nor UO_614 (O_614,N_18211,N_18107);
and UO_615 (O_615,N_18267,N_18576);
or UO_616 (O_616,N_19429,N_19161);
xnor UO_617 (O_617,N_18361,N_19745);
nor UO_618 (O_618,N_18497,N_18961);
nor UO_619 (O_619,N_19710,N_19548);
or UO_620 (O_620,N_18741,N_18775);
nand UO_621 (O_621,N_18678,N_19835);
or UO_622 (O_622,N_18304,N_18621);
or UO_623 (O_623,N_19094,N_19335);
and UO_624 (O_624,N_19401,N_18499);
or UO_625 (O_625,N_19516,N_19079);
or UO_626 (O_626,N_18018,N_19431);
or UO_627 (O_627,N_18023,N_18761);
or UO_628 (O_628,N_18396,N_19206);
nand UO_629 (O_629,N_18445,N_19007);
or UO_630 (O_630,N_18215,N_19906);
or UO_631 (O_631,N_18996,N_18788);
or UO_632 (O_632,N_19355,N_19247);
nand UO_633 (O_633,N_18163,N_18926);
nand UO_634 (O_634,N_18100,N_18913);
and UO_635 (O_635,N_19846,N_19499);
nand UO_636 (O_636,N_19811,N_19518);
nand UO_637 (O_637,N_19852,N_18549);
and UO_638 (O_638,N_18003,N_18522);
nand UO_639 (O_639,N_18047,N_18665);
nand UO_640 (O_640,N_18841,N_19015);
or UO_641 (O_641,N_19929,N_18902);
and UO_642 (O_642,N_19715,N_18793);
nor UO_643 (O_643,N_18094,N_18864);
nand UO_644 (O_644,N_19909,N_18972);
nand UO_645 (O_645,N_19503,N_19827);
or UO_646 (O_646,N_19163,N_18968);
nor UO_647 (O_647,N_19935,N_18810);
nor UO_648 (O_648,N_19991,N_18093);
nand UO_649 (O_649,N_19088,N_19205);
nor UO_650 (O_650,N_18263,N_18674);
nand UO_651 (O_651,N_19659,N_18319);
xnor UO_652 (O_652,N_18923,N_18460);
nand UO_653 (O_653,N_19864,N_18295);
nand UO_654 (O_654,N_18757,N_18228);
nand UO_655 (O_655,N_18150,N_19660);
nor UO_656 (O_656,N_19488,N_19732);
or UO_657 (O_657,N_19365,N_19388);
nand UO_658 (O_658,N_19533,N_18177);
nor UO_659 (O_659,N_18002,N_19618);
nand UO_660 (O_660,N_19316,N_19998);
or UO_661 (O_661,N_19725,N_19791);
nand UO_662 (O_662,N_19989,N_19754);
or UO_663 (O_663,N_19403,N_18013);
and UO_664 (O_664,N_18662,N_18446);
nor UO_665 (O_665,N_18531,N_18000);
nand UO_666 (O_666,N_18326,N_18893);
or UO_667 (O_667,N_18219,N_19070);
nor UO_668 (O_668,N_19417,N_18850);
nor UO_669 (O_669,N_19081,N_19502);
nor UO_670 (O_670,N_19759,N_19082);
nand UO_671 (O_671,N_18365,N_19826);
and UO_672 (O_672,N_19295,N_18762);
nor UO_673 (O_673,N_19579,N_19006);
nand UO_674 (O_674,N_18104,N_19272);
and UO_675 (O_675,N_18363,N_18661);
nor UO_676 (O_676,N_19491,N_18156);
and UO_677 (O_677,N_18059,N_19124);
xnor UO_678 (O_678,N_19749,N_18080);
nand UO_679 (O_679,N_18906,N_18884);
or UO_680 (O_680,N_18602,N_19265);
nand UO_681 (O_681,N_19896,N_19814);
nand UO_682 (O_682,N_18085,N_19411);
nor UO_683 (O_683,N_19880,N_19110);
nor UO_684 (O_684,N_18004,N_19478);
nor UO_685 (O_685,N_18918,N_18667);
nor UO_686 (O_686,N_18260,N_19829);
or UO_687 (O_687,N_19700,N_18897);
and UO_688 (O_688,N_19046,N_18558);
nand UO_689 (O_689,N_18705,N_18908);
or UO_690 (O_690,N_19559,N_19151);
nor UO_691 (O_691,N_19750,N_19804);
nand UO_692 (O_692,N_19293,N_18519);
nand UO_693 (O_693,N_19096,N_18619);
nor UO_694 (O_694,N_18317,N_19389);
nor UO_695 (O_695,N_18595,N_18740);
or UO_696 (O_696,N_18940,N_19643);
nand UO_697 (O_697,N_18794,N_19549);
nor UO_698 (O_698,N_18896,N_18575);
nand UO_699 (O_699,N_18779,N_18631);
nor UO_700 (O_700,N_18404,N_19577);
nand UO_701 (O_701,N_18879,N_19812);
nor UO_702 (O_702,N_19474,N_19291);
or UO_703 (O_703,N_19627,N_18479);
and UO_704 (O_704,N_19086,N_18384);
or UO_705 (O_705,N_18814,N_19670);
and UO_706 (O_706,N_18463,N_19368);
or UO_707 (O_707,N_19422,N_19164);
or UO_708 (O_708,N_19624,N_19801);
and UO_709 (O_709,N_19837,N_19679);
nand UO_710 (O_710,N_18185,N_18417);
nand UO_711 (O_711,N_19105,N_18114);
nor UO_712 (O_712,N_18545,N_19748);
nand UO_713 (O_713,N_18980,N_19255);
and UO_714 (O_714,N_19279,N_19333);
or UO_715 (O_715,N_19452,N_19861);
nor UO_716 (O_716,N_19739,N_18746);
or UO_717 (O_717,N_18403,N_18967);
or UO_718 (O_718,N_19475,N_18153);
and UO_719 (O_719,N_18420,N_19721);
nor UO_720 (O_720,N_18573,N_19792);
nor UO_721 (O_721,N_19527,N_19271);
or UO_722 (O_722,N_19385,N_19795);
nand UO_723 (O_723,N_18950,N_18205);
nand UO_724 (O_724,N_18627,N_19613);
or UO_725 (O_725,N_19354,N_19095);
xor UO_726 (O_726,N_19818,N_19315);
and UO_727 (O_727,N_19881,N_19819);
nand UO_728 (O_728,N_18587,N_18431);
and UO_729 (O_729,N_19634,N_18359);
nor UO_730 (O_730,N_18766,N_18238);
and UO_731 (O_731,N_19332,N_18782);
and UO_732 (O_732,N_18043,N_19185);
and UO_733 (O_733,N_19303,N_19201);
and UO_734 (O_734,N_18812,N_18118);
nand UO_735 (O_735,N_19041,N_18937);
or UO_736 (O_736,N_19805,N_18865);
nand UO_737 (O_737,N_18300,N_18474);
nor UO_738 (O_738,N_19305,N_18286);
nand UO_739 (O_739,N_18034,N_19951);
and UO_740 (O_740,N_18213,N_18912);
and UO_741 (O_741,N_19619,N_18495);
and UO_742 (O_742,N_18946,N_19565);
nand UO_743 (O_743,N_19856,N_19356);
or UO_744 (O_744,N_18031,N_18344);
or UO_745 (O_745,N_18098,N_19193);
nor UO_746 (O_746,N_18516,N_19500);
and UO_747 (O_747,N_18246,N_19065);
nor UO_748 (O_748,N_19941,N_18889);
or UO_749 (O_749,N_19453,N_18386);
nand UO_750 (O_750,N_19220,N_18805);
or UO_751 (O_751,N_19802,N_18071);
or UO_752 (O_752,N_18925,N_18369);
nand UO_753 (O_753,N_18718,N_19673);
or UO_754 (O_754,N_19407,N_18824);
nor UO_755 (O_755,N_19641,N_18373);
nand UO_756 (O_756,N_19677,N_18687);
nand UO_757 (O_757,N_19063,N_18184);
or UO_758 (O_758,N_19900,N_19842);
nand UO_759 (O_759,N_18236,N_18487);
nand UO_760 (O_760,N_19361,N_19307);
and UO_761 (O_761,N_18117,N_19251);
nand UO_762 (O_762,N_19413,N_18724);
nand UO_763 (O_763,N_18078,N_18787);
or UO_764 (O_764,N_18981,N_18592);
nor UO_765 (O_765,N_19705,N_18625);
or UO_766 (O_766,N_19756,N_19129);
nand UO_767 (O_767,N_19216,N_18534);
nand UO_768 (O_768,N_18470,N_19378);
or UO_769 (O_769,N_19886,N_18895);
or UO_770 (O_770,N_19687,N_18112);
or UO_771 (O_771,N_18799,N_19469);
or UO_772 (O_772,N_18796,N_18480);
or UO_773 (O_773,N_18773,N_19973);
nand UO_774 (O_774,N_18603,N_19167);
or UO_775 (O_775,N_19576,N_18130);
nand UO_776 (O_776,N_18005,N_18507);
nor UO_777 (O_777,N_19150,N_18685);
or UO_778 (O_778,N_19932,N_19850);
or UO_779 (O_779,N_19414,N_19244);
nand UO_780 (O_780,N_19714,N_19684);
or UO_781 (O_781,N_19735,N_19405);
nand UO_782 (O_782,N_19131,N_19611);
and UO_783 (O_783,N_19604,N_18529);
or UO_784 (O_784,N_19961,N_19682);
or UO_785 (O_785,N_19168,N_19069);
or UO_786 (O_786,N_18845,N_18550);
and UO_787 (O_787,N_18892,N_18401);
nor UO_788 (O_788,N_19484,N_19454);
nor UO_789 (O_789,N_19138,N_19784);
and UO_790 (O_790,N_18680,N_19428);
or UO_791 (O_791,N_19981,N_18196);
and UO_792 (O_792,N_18165,N_19327);
and UO_793 (O_793,N_18419,N_18727);
and UO_794 (O_794,N_19971,N_18218);
and UO_795 (O_795,N_19050,N_19459);
nor UO_796 (O_796,N_18966,N_18131);
nand UO_797 (O_797,N_18356,N_18647);
and UO_798 (O_798,N_18683,N_18217);
nor UO_799 (O_799,N_19945,N_19510);
and UO_800 (O_800,N_19480,N_18347);
or UO_801 (O_801,N_18169,N_18383);
nand UO_802 (O_802,N_19117,N_19956);
and UO_803 (O_803,N_18525,N_19495);
nand UO_804 (O_804,N_19339,N_19944);
or UO_805 (O_805,N_18907,N_18605);
nor UO_806 (O_806,N_18748,N_18939);
nor UO_807 (O_807,N_19177,N_19556);
nand UO_808 (O_808,N_18515,N_19262);
nor UO_809 (O_809,N_18588,N_19911);
nand UO_810 (O_810,N_19524,N_19622);
nor UO_811 (O_811,N_19441,N_19274);
nor UO_812 (O_812,N_18565,N_19492);
and UO_813 (O_813,N_19890,N_19889);
nor UO_814 (O_814,N_19277,N_19702);
nand UO_815 (O_815,N_19097,N_19810);
nor UO_816 (O_816,N_18400,N_18560);
or UO_817 (O_817,N_18759,N_19197);
nand UO_818 (O_818,N_19645,N_18606);
nand UO_819 (O_819,N_18422,N_19224);
and UO_820 (O_820,N_18442,N_18335);
or UO_821 (O_821,N_19586,N_18173);
or UO_822 (O_822,N_19605,N_18379);
nand UO_823 (O_823,N_18418,N_18970);
or UO_824 (O_824,N_19514,N_19367);
nor UO_825 (O_825,N_18340,N_19894);
nor UO_826 (O_826,N_18878,N_18816);
or UO_827 (O_827,N_19671,N_18726);
nor UO_828 (O_828,N_19462,N_19773);
and UO_829 (O_829,N_19308,N_19903);
nor UO_830 (O_830,N_18249,N_19934);
nand UO_831 (O_831,N_18720,N_19467);
nand UO_832 (O_832,N_18293,N_18954);
or UO_833 (O_833,N_19768,N_18289);
nor UO_834 (O_834,N_18248,N_18604);
or UO_835 (O_835,N_19330,N_18584);
and UO_836 (O_836,N_19282,N_18440);
nand UO_837 (O_837,N_19925,N_18280);
and UO_838 (O_838,N_19992,N_19450);
and UO_839 (O_839,N_19871,N_18781);
nand UO_840 (O_840,N_19926,N_18559);
and UO_841 (O_841,N_19520,N_18221);
or UO_842 (O_842,N_19751,N_19175);
and UO_843 (O_843,N_18405,N_19825);
and UO_844 (O_844,N_19430,N_18763);
nand UO_845 (O_845,N_19870,N_18710);
and UO_846 (O_846,N_19584,N_18367);
or UO_847 (O_847,N_19642,N_19930);
or UO_848 (O_848,N_19123,N_19465);
nand UO_849 (O_849,N_19594,N_18669);
or UO_850 (O_850,N_19639,N_19136);
and UO_851 (O_851,N_19382,N_18443);
nor UO_852 (O_852,N_19904,N_19555);
or UO_853 (O_853,N_18486,N_18342);
nand UO_854 (O_854,N_19602,N_18935);
or UO_855 (O_855,N_19022,N_18760);
nand UO_856 (O_856,N_18458,N_19025);
nand UO_857 (O_857,N_18622,N_19640);
nand UO_858 (O_858,N_18754,N_19798);
nor UO_859 (O_859,N_19902,N_18498);
nor UO_860 (O_860,N_19020,N_18842);
nand UO_861 (O_861,N_19570,N_19506);
xor UO_862 (O_862,N_18696,N_19666);
and UO_863 (O_863,N_18261,N_19914);
nand UO_864 (O_864,N_19987,N_19415);
or UO_865 (O_865,N_19529,N_18113);
or UO_866 (O_866,N_19039,N_19017);
nand UO_867 (O_867,N_19292,N_19581);
nor UO_868 (O_868,N_18048,N_19098);
nor UO_869 (O_869,N_18435,N_19652);
or UO_870 (O_870,N_18372,N_18843);
and UO_871 (O_871,N_18222,N_19329);
xnor UO_872 (O_872,N_19093,N_18630);
or UO_873 (O_873,N_18513,N_19090);
nand UO_874 (O_874,N_19723,N_18149);
or UO_875 (O_875,N_18476,N_18634);
nor UO_876 (O_876,N_19822,N_18472);
and UO_877 (O_877,N_19891,N_19984);
nand UO_878 (O_878,N_18307,N_19966);
or UO_879 (O_879,N_19726,N_19026);
or UO_880 (O_880,N_18322,N_18666);
nor UO_881 (O_881,N_18872,N_19047);
nand UO_882 (O_882,N_18581,N_18983);
and UO_883 (O_883,N_19839,N_18457);
or UO_884 (O_884,N_18639,N_19545);
nor UO_885 (O_885,N_18202,N_19922);
or UO_886 (O_886,N_18152,N_18448);
or UO_887 (O_887,N_19029,N_19318);
and UO_888 (O_888,N_18691,N_18108);
nand UO_889 (O_889,N_18345,N_19089);
nand UO_890 (O_890,N_18137,N_18321);
nand UO_891 (O_891,N_18186,N_19767);
nand UO_892 (O_892,N_19960,N_19326);
nand UO_893 (O_893,N_19866,N_19568);
or UO_894 (O_894,N_18774,N_18591);
nor UO_895 (O_895,N_19915,N_18934);
or UO_896 (O_896,N_19635,N_18684);
and UO_897 (O_897,N_18455,N_19106);
nor UO_898 (O_898,N_18732,N_18689);
nor UO_899 (O_899,N_19358,N_19074);
nand UO_900 (O_900,N_18239,N_18491);
nor UO_901 (O_901,N_18829,N_19189);
or UO_902 (O_902,N_18010,N_18170);
and UO_903 (O_903,N_19959,N_19463);
nor UO_904 (O_904,N_19267,N_18087);
nor UO_905 (O_905,N_19141,N_18927);
and UO_906 (O_906,N_18014,N_18795);
nand UO_907 (O_907,N_18329,N_19853);
nor UO_908 (O_908,N_18265,N_18099);
and UO_909 (O_909,N_18881,N_18388);
nand UO_910 (O_910,N_18541,N_19119);
and UO_911 (O_911,N_18456,N_18393);
or UO_912 (O_912,N_18485,N_19223);
or UO_913 (O_913,N_19761,N_18863);
nor UO_914 (O_914,N_19421,N_18564);
nand UO_915 (O_915,N_18421,N_19967);
nor UO_916 (O_916,N_18597,N_18542);
nand UO_917 (O_917,N_18988,N_19187);
and UO_918 (O_918,N_18241,N_19218);
or UO_919 (O_919,N_18725,N_19169);
nand UO_920 (O_920,N_19596,N_19370);
nand UO_921 (O_921,N_19566,N_18737);
or UO_922 (O_922,N_19636,N_19042);
or UO_923 (O_923,N_18337,N_19691);
or UO_924 (O_924,N_18847,N_18305);
nor UO_925 (O_925,N_18168,N_19933);
or UO_926 (O_926,N_19309,N_19451);
and UO_927 (O_927,N_18951,N_18586);
or UO_928 (O_928,N_19391,N_18963);
and UO_929 (O_929,N_19564,N_18492);
nand UO_930 (O_930,N_19142,N_19121);
and UO_931 (O_931,N_18243,N_18745);
and UO_932 (O_932,N_18015,N_18064);
nor UO_933 (O_933,N_18548,N_19446);
nor UO_934 (O_934,N_19229,N_18336);
nand UO_935 (O_935,N_18637,N_19986);
nand UO_936 (O_936,N_18438,N_18203);
or UO_937 (O_937,N_18147,N_18123);
or UO_938 (O_938,N_18784,N_19456);
xnor UO_939 (O_939,N_18437,N_19227);
or UO_940 (O_940,N_19591,N_18127);
or UO_941 (O_941,N_18086,N_18012);
and UO_942 (O_942,N_18109,N_19676);
or UO_943 (O_943,N_18651,N_19884);
nor UO_944 (O_944,N_19873,N_18397);
and UO_945 (O_945,N_19314,N_18055);
or UO_946 (O_946,N_18751,N_18425);
nor UO_947 (O_947,N_19191,N_18772);
or UO_948 (O_948,N_18992,N_18399);
nand UO_949 (O_949,N_19690,N_18088);
nand UO_950 (O_950,N_18315,N_18194);
nor UO_951 (O_951,N_18409,N_18916);
or UO_952 (O_952,N_18932,N_18825);
or UO_953 (O_953,N_18613,N_19975);
nor UO_954 (O_954,N_19018,N_19449);
nand UO_955 (O_955,N_19104,N_19344);
nor UO_956 (O_956,N_19263,N_18876);
nand UO_957 (O_957,N_18506,N_19551);
or UO_958 (O_958,N_19266,N_19716);
nor UO_959 (O_959,N_19051,N_19283);
nand UO_960 (O_960,N_18294,N_19055);
xnor UO_961 (O_961,N_18649,N_19755);
xnor UO_962 (O_962,N_19931,N_19497);
or UO_963 (O_963,N_19408,N_19345);
or UO_964 (O_964,N_19264,N_19892);
and UO_965 (O_965,N_19237,N_19663);
and UO_966 (O_966,N_18778,N_18439);
and UO_967 (O_967,N_18851,N_19486);
and UO_968 (O_968,N_18632,N_19995);
or UO_969 (O_969,N_19083,N_19724);
or UO_970 (O_970,N_18467,N_19049);
nor UO_971 (O_971,N_19950,N_19661);
or UO_972 (O_972,N_18011,N_18157);
or UO_973 (O_973,N_18042,N_19003);
and UO_974 (O_974,N_19384,N_19774);
nor UO_975 (O_975,N_18251,N_18370);
and UO_976 (O_976,N_18673,N_19780);
nand UO_977 (O_977,N_19016,N_19868);
nor UO_978 (O_978,N_19994,N_18849);
nand UO_979 (O_979,N_19404,N_19162);
and UO_980 (O_980,N_18339,N_18698);
nor UO_981 (O_981,N_18183,N_18803);
nand UO_982 (O_982,N_19154,N_18133);
nand UO_983 (O_983,N_19447,N_18316);
xnor UO_984 (O_984,N_19872,N_19290);
nor UO_985 (O_985,N_19060,N_19820);
and UO_986 (O_986,N_19458,N_18914);
and UO_987 (O_987,N_19947,N_18036);
or UO_988 (O_988,N_18331,N_18848);
nand UO_989 (O_989,N_18301,N_19540);
nor UO_990 (O_990,N_19371,N_19730);
and UO_991 (O_991,N_19256,N_18552);
and UO_992 (O_992,N_18820,N_19156);
and UO_993 (O_993,N_19233,N_18853);
and UO_994 (O_994,N_18210,N_19983);
xnor UO_995 (O_995,N_18197,N_19198);
xnor UO_996 (O_996,N_19319,N_19612);
and UO_997 (O_997,N_19874,N_18424);
and UO_998 (O_998,N_19722,N_18193);
nor UO_999 (O_999,N_18352,N_19392);
nor UO_1000 (O_1000,N_19852,N_19360);
nand UO_1001 (O_1001,N_18467,N_19437);
and UO_1002 (O_1002,N_18560,N_18455);
or UO_1003 (O_1003,N_18528,N_18490);
xnor UO_1004 (O_1004,N_19221,N_18260);
nor UO_1005 (O_1005,N_18345,N_18289);
or UO_1006 (O_1006,N_18172,N_19242);
nand UO_1007 (O_1007,N_18684,N_19713);
and UO_1008 (O_1008,N_18284,N_18646);
nor UO_1009 (O_1009,N_19602,N_19467);
or UO_1010 (O_1010,N_19735,N_18611);
or UO_1011 (O_1011,N_19307,N_19257);
and UO_1012 (O_1012,N_19780,N_18774);
nand UO_1013 (O_1013,N_18094,N_18045);
or UO_1014 (O_1014,N_19582,N_19315);
nand UO_1015 (O_1015,N_19176,N_18539);
or UO_1016 (O_1016,N_19531,N_19707);
nand UO_1017 (O_1017,N_18449,N_19163);
nand UO_1018 (O_1018,N_18361,N_19935);
or UO_1019 (O_1019,N_19188,N_19186);
nand UO_1020 (O_1020,N_19025,N_18169);
and UO_1021 (O_1021,N_18793,N_18612);
nand UO_1022 (O_1022,N_18988,N_18850);
nand UO_1023 (O_1023,N_19684,N_19075);
and UO_1024 (O_1024,N_18702,N_19640);
nand UO_1025 (O_1025,N_19985,N_18276);
and UO_1026 (O_1026,N_19317,N_18171);
nand UO_1027 (O_1027,N_18251,N_18739);
nand UO_1028 (O_1028,N_18086,N_18935);
nor UO_1029 (O_1029,N_18616,N_18307);
or UO_1030 (O_1030,N_19555,N_18706);
xor UO_1031 (O_1031,N_19477,N_18261);
or UO_1032 (O_1032,N_19192,N_19077);
or UO_1033 (O_1033,N_18070,N_19598);
or UO_1034 (O_1034,N_18593,N_18319);
or UO_1035 (O_1035,N_19825,N_19538);
and UO_1036 (O_1036,N_18301,N_18191);
nand UO_1037 (O_1037,N_18871,N_18804);
nor UO_1038 (O_1038,N_19229,N_18148);
and UO_1039 (O_1039,N_18376,N_19373);
and UO_1040 (O_1040,N_18412,N_19332);
or UO_1041 (O_1041,N_18800,N_19917);
and UO_1042 (O_1042,N_18641,N_19209);
or UO_1043 (O_1043,N_19957,N_18847);
or UO_1044 (O_1044,N_18903,N_18053);
and UO_1045 (O_1045,N_19452,N_18580);
nor UO_1046 (O_1046,N_18854,N_19894);
or UO_1047 (O_1047,N_18789,N_18175);
nor UO_1048 (O_1048,N_18118,N_18726);
nor UO_1049 (O_1049,N_19727,N_18537);
and UO_1050 (O_1050,N_19125,N_18319);
and UO_1051 (O_1051,N_18896,N_18108);
nor UO_1052 (O_1052,N_18556,N_18558);
nor UO_1053 (O_1053,N_18924,N_18647);
xnor UO_1054 (O_1054,N_19682,N_19467);
nand UO_1055 (O_1055,N_19290,N_18458);
nor UO_1056 (O_1056,N_19328,N_19292);
and UO_1057 (O_1057,N_19161,N_19238);
or UO_1058 (O_1058,N_19711,N_18912);
nor UO_1059 (O_1059,N_18404,N_19666);
or UO_1060 (O_1060,N_18962,N_18501);
or UO_1061 (O_1061,N_18248,N_19171);
and UO_1062 (O_1062,N_19084,N_18090);
nor UO_1063 (O_1063,N_18911,N_18784);
nand UO_1064 (O_1064,N_19552,N_19968);
or UO_1065 (O_1065,N_18542,N_18684);
nand UO_1066 (O_1066,N_19215,N_18504);
and UO_1067 (O_1067,N_19135,N_18186);
and UO_1068 (O_1068,N_18113,N_19039);
nand UO_1069 (O_1069,N_18166,N_18032);
and UO_1070 (O_1070,N_19152,N_18393);
nor UO_1071 (O_1071,N_19106,N_18381);
and UO_1072 (O_1072,N_18993,N_18075);
or UO_1073 (O_1073,N_18760,N_18896);
nor UO_1074 (O_1074,N_19643,N_19465);
or UO_1075 (O_1075,N_18947,N_18658);
nand UO_1076 (O_1076,N_19576,N_19322);
and UO_1077 (O_1077,N_18496,N_19778);
xnor UO_1078 (O_1078,N_19253,N_18654);
nand UO_1079 (O_1079,N_19726,N_18676);
nor UO_1080 (O_1080,N_18135,N_18677);
and UO_1081 (O_1081,N_18134,N_18114);
xnor UO_1082 (O_1082,N_19754,N_19082);
or UO_1083 (O_1083,N_19008,N_18034);
nand UO_1084 (O_1084,N_18416,N_18341);
nand UO_1085 (O_1085,N_18645,N_18208);
nor UO_1086 (O_1086,N_18754,N_19339);
nor UO_1087 (O_1087,N_19457,N_18254);
or UO_1088 (O_1088,N_19563,N_18395);
nand UO_1089 (O_1089,N_19502,N_18116);
nor UO_1090 (O_1090,N_18758,N_19440);
xnor UO_1091 (O_1091,N_18544,N_19984);
nand UO_1092 (O_1092,N_19610,N_18840);
or UO_1093 (O_1093,N_18634,N_18084);
nor UO_1094 (O_1094,N_18729,N_19906);
nor UO_1095 (O_1095,N_18615,N_19840);
nand UO_1096 (O_1096,N_18676,N_18417);
or UO_1097 (O_1097,N_19888,N_19765);
and UO_1098 (O_1098,N_19137,N_19534);
or UO_1099 (O_1099,N_18216,N_18113);
and UO_1100 (O_1100,N_19144,N_19329);
nand UO_1101 (O_1101,N_19376,N_19246);
nand UO_1102 (O_1102,N_18065,N_19069);
nor UO_1103 (O_1103,N_19220,N_19608);
nand UO_1104 (O_1104,N_19244,N_19490);
or UO_1105 (O_1105,N_19652,N_18338);
and UO_1106 (O_1106,N_18764,N_19691);
nand UO_1107 (O_1107,N_19575,N_18312);
and UO_1108 (O_1108,N_18845,N_18619);
or UO_1109 (O_1109,N_18660,N_19397);
and UO_1110 (O_1110,N_18837,N_18204);
or UO_1111 (O_1111,N_18606,N_19351);
and UO_1112 (O_1112,N_19206,N_18430);
and UO_1113 (O_1113,N_18478,N_19439);
and UO_1114 (O_1114,N_18255,N_18666);
or UO_1115 (O_1115,N_18149,N_18419);
or UO_1116 (O_1116,N_19573,N_19852);
or UO_1117 (O_1117,N_19026,N_18078);
or UO_1118 (O_1118,N_19382,N_18574);
or UO_1119 (O_1119,N_18378,N_18884);
or UO_1120 (O_1120,N_19606,N_18917);
nor UO_1121 (O_1121,N_18125,N_18350);
and UO_1122 (O_1122,N_19517,N_18828);
or UO_1123 (O_1123,N_18272,N_19520);
or UO_1124 (O_1124,N_18579,N_19864);
nand UO_1125 (O_1125,N_19122,N_18937);
and UO_1126 (O_1126,N_19359,N_18263);
nor UO_1127 (O_1127,N_18478,N_18933);
nand UO_1128 (O_1128,N_19310,N_19737);
or UO_1129 (O_1129,N_19528,N_19617);
and UO_1130 (O_1130,N_18144,N_18826);
nor UO_1131 (O_1131,N_18245,N_19484);
or UO_1132 (O_1132,N_19149,N_18986);
nand UO_1133 (O_1133,N_19278,N_19822);
nand UO_1134 (O_1134,N_19172,N_18597);
nor UO_1135 (O_1135,N_18264,N_18572);
nor UO_1136 (O_1136,N_19348,N_18561);
and UO_1137 (O_1137,N_19061,N_18848);
and UO_1138 (O_1138,N_19184,N_19356);
and UO_1139 (O_1139,N_18500,N_19680);
and UO_1140 (O_1140,N_18352,N_18214);
or UO_1141 (O_1141,N_19728,N_18211);
or UO_1142 (O_1142,N_19273,N_19648);
nor UO_1143 (O_1143,N_19554,N_18683);
nand UO_1144 (O_1144,N_18279,N_18209);
or UO_1145 (O_1145,N_19590,N_19694);
nand UO_1146 (O_1146,N_18916,N_19749);
nand UO_1147 (O_1147,N_19949,N_18504);
nand UO_1148 (O_1148,N_18426,N_18610);
or UO_1149 (O_1149,N_18051,N_18033);
and UO_1150 (O_1150,N_19916,N_19870);
or UO_1151 (O_1151,N_18999,N_19238);
nor UO_1152 (O_1152,N_19500,N_18300);
nand UO_1153 (O_1153,N_18277,N_19824);
nand UO_1154 (O_1154,N_19219,N_18451);
and UO_1155 (O_1155,N_18266,N_18355);
or UO_1156 (O_1156,N_18173,N_18240);
or UO_1157 (O_1157,N_18845,N_19204);
and UO_1158 (O_1158,N_19588,N_18867);
nand UO_1159 (O_1159,N_19405,N_18674);
and UO_1160 (O_1160,N_18835,N_19171);
nand UO_1161 (O_1161,N_19364,N_18894);
nor UO_1162 (O_1162,N_18408,N_19920);
nand UO_1163 (O_1163,N_18736,N_18112);
nor UO_1164 (O_1164,N_19950,N_19768);
and UO_1165 (O_1165,N_19492,N_19350);
nor UO_1166 (O_1166,N_18177,N_18411);
nor UO_1167 (O_1167,N_18475,N_18106);
nor UO_1168 (O_1168,N_18442,N_19266);
nand UO_1169 (O_1169,N_19555,N_19779);
nand UO_1170 (O_1170,N_19587,N_19708);
nand UO_1171 (O_1171,N_18874,N_18492);
nor UO_1172 (O_1172,N_19076,N_18111);
nor UO_1173 (O_1173,N_19330,N_18610);
and UO_1174 (O_1174,N_19834,N_19536);
nor UO_1175 (O_1175,N_19607,N_18345);
nor UO_1176 (O_1176,N_19568,N_19507);
or UO_1177 (O_1177,N_18441,N_19456);
or UO_1178 (O_1178,N_19194,N_18472);
and UO_1179 (O_1179,N_19381,N_19569);
or UO_1180 (O_1180,N_19167,N_19431);
or UO_1181 (O_1181,N_19144,N_18820);
xor UO_1182 (O_1182,N_19856,N_19241);
nand UO_1183 (O_1183,N_19096,N_19661);
or UO_1184 (O_1184,N_19280,N_19661);
xnor UO_1185 (O_1185,N_18854,N_19172);
and UO_1186 (O_1186,N_18472,N_18100);
nand UO_1187 (O_1187,N_19797,N_19491);
and UO_1188 (O_1188,N_18449,N_18673);
nand UO_1189 (O_1189,N_18811,N_18993);
and UO_1190 (O_1190,N_18808,N_19606);
nor UO_1191 (O_1191,N_19790,N_19843);
or UO_1192 (O_1192,N_18208,N_19520);
nand UO_1193 (O_1193,N_18775,N_19568);
and UO_1194 (O_1194,N_18440,N_18743);
or UO_1195 (O_1195,N_19339,N_18510);
xor UO_1196 (O_1196,N_19012,N_19978);
and UO_1197 (O_1197,N_19376,N_19251);
nand UO_1198 (O_1198,N_19820,N_19698);
and UO_1199 (O_1199,N_19007,N_18367);
and UO_1200 (O_1200,N_18857,N_18806);
nor UO_1201 (O_1201,N_18179,N_18670);
and UO_1202 (O_1202,N_18803,N_19511);
nand UO_1203 (O_1203,N_19748,N_19608);
or UO_1204 (O_1204,N_19434,N_19488);
nand UO_1205 (O_1205,N_18279,N_18244);
and UO_1206 (O_1206,N_19842,N_19282);
nor UO_1207 (O_1207,N_19892,N_18795);
nor UO_1208 (O_1208,N_19901,N_18126);
and UO_1209 (O_1209,N_18560,N_19404);
or UO_1210 (O_1210,N_18450,N_18019);
or UO_1211 (O_1211,N_19646,N_18947);
nand UO_1212 (O_1212,N_19894,N_19178);
nand UO_1213 (O_1213,N_18695,N_19384);
or UO_1214 (O_1214,N_18963,N_18387);
nand UO_1215 (O_1215,N_19380,N_19932);
and UO_1216 (O_1216,N_18006,N_18620);
or UO_1217 (O_1217,N_19438,N_19575);
nor UO_1218 (O_1218,N_19013,N_18493);
and UO_1219 (O_1219,N_18463,N_19708);
or UO_1220 (O_1220,N_19174,N_18025);
nor UO_1221 (O_1221,N_18005,N_19318);
and UO_1222 (O_1222,N_18790,N_19315);
nand UO_1223 (O_1223,N_18706,N_19115);
or UO_1224 (O_1224,N_18851,N_19663);
and UO_1225 (O_1225,N_18183,N_19810);
nor UO_1226 (O_1226,N_18497,N_18080);
or UO_1227 (O_1227,N_19939,N_19831);
nor UO_1228 (O_1228,N_18334,N_19662);
nand UO_1229 (O_1229,N_18109,N_19803);
nor UO_1230 (O_1230,N_18709,N_18280);
nand UO_1231 (O_1231,N_18095,N_19106);
nor UO_1232 (O_1232,N_18209,N_18374);
nor UO_1233 (O_1233,N_19974,N_19414);
nor UO_1234 (O_1234,N_19384,N_19279);
or UO_1235 (O_1235,N_19828,N_19985);
or UO_1236 (O_1236,N_19296,N_19693);
and UO_1237 (O_1237,N_18719,N_18132);
nand UO_1238 (O_1238,N_18375,N_19610);
nor UO_1239 (O_1239,N_19325,N_19653);
nand UO_1240 (O_1240,N_18418,N_19341);
nand UO_1241 (O_1241,N_18269,N_19981);
nor UO_1242 (O_1242,N_19747,N_19133);
nand UO_1243 (O_1243,N_19755,N_19388);
nor UO_1244 (O_1244,N_19371,N_19490);
nor UO_1245 (O_1245,N_18283,N_18526);
nand UO_1246 (O_1246,N_19151,N_18821);
or UO_1247 (O_1247,N_19074,N_18428);
and UO_1248 (O_1248,N_19592,N_19549);
nand UO_1249 (O_1249,N_19129,N_18298);
nor UO_1250 (O_1250,N_19386,N_19878);
and UO_1251 (O_1251,N_18194,N_19751);
and UO_1252 (O_1252,N_19005,N_18888);
or UO_1253 (O_1253,N_19764,N_19754);
or UO_1254 (O_1254,N_19172,N_18523);
nand UO_1255 (O_1255,N_19840,N_18836);
or UO_1256 (O_1256,N_18478,N_19003);
nor UO_1257 (O_1257,N_19127,N_18929);
or UO_1258 (O_1258,N_18712,N_19666);
or UO_1259 (O_1259,N_18091,N_19387);
nand UO_1260 (O_1260,N_19231,N_19714);
and UO_1261 (O_1261,N_18527,N_18967);
and UO_1262 (O_1262,N_19375,N_18956);
nor UO_1263 (O_1263,N_18713,N_19106);
nand UO_1264 (O_1264,N_18184,N_18457);
or UO_1265 (O_1265,N_19284,N_19817);
and UO_1266 (O_1266,N_19666,N_19418);
or UO_1267 (O_1267,N_18677,N_19685);
nand UO_1268 (O_1268,N_19867,N_19231);
or UO_1269 (O_1269,N_19583,N_18511);
xnor UO_1270 (O_1270,N_19166,N_19086);
or UO_1271 (O_1271,N_19859,N_19395);
nand UO_1272 (O_1272,N_19846,N_18459);
and UO_1273 (O_1273,N_18101,N_18984);
nand UO_1274 (O_1274,N_19344,N_18656);
or UO_1275 (O_1275,N_19543,N_18113);
or UO_1276 (O_1276,N_18207,N_18021);
or UO_1277 (O_1277,N_18910,N_18803);
and UO_1278 (O_1278,N_18929,N_18956);
and UO_1279 (O_1279,N_19841,N_19468);
nor UO_1280 (O_1280,N_19669,N_18382);
or UO_1281 (O_1281,N_19634,N_18924);
or UO_1282 (O_1282,N_19417,N_19310);
and UO_1283 (O_1283,N_18605,N_18871);
nand UO_1284 (O_1284,N_18110,N_18323);
or UO_1285 (O_1285,N_18349,N_19709);
and UO_1286 (O_1286,N_18452,N_19656);
nor UO_1287 (O_1287,N_18896,N_18599);
and UO_1288 (O_1288,N_19297,N_19062);
or UO_1289 (O_1289,N_19423,N_18004);
or UO_1290 (O_1290,N_19581,N_19080);
nor UO_1291 (O_1291,N_19275,N_18339);
nand UO_1292 (O_1292,N_18912,N_18071);
and UO_1293 (O_1293,N_19786,N_19076);
nor UO_1294 (O_1294,N_19792,N_19539);
nand UO_1295 (O_1295,N_19680,N_19181);
nor UO_1296 (O_1296,N_18848,N_19230);
nor UO_1297 (O_1297,N_18719,N_19327);
or UO_1298 (O_1298,N_19492,N_19530);
nand UO_1299 (O_1299,N_19954,N_18518);
or UO_1300 (O_1300,N_19997,N_18286);
and UO_1301 (O_1301,N_19090,N_19921);
nor UO_1302 (O_1302,N_19868,N_18765);
nor UO_1303 (O_1303,N_18026,N_19920);
or UO_1304 (O_1304,N_18725,N_18973);
nor UO_1305 (O_1305,N_19786,N_19740);
nor UO_1306 (O_1306,N_19940,N_19802);
or UO_1307 (O_1307,N_19002,N_18611);
nor UO_1308 (O_1308,N_18827,N_18441);
nor UO_1309 (O_1309,N_19538,N_19970);
or UO_1310 (O_1310,N_18987,N_19112);
nand UO_1311 (O_1311,N_18468,N_18131);
nor UO_1312 (O_1312,N_19821,N_19422);
nand UO_1313 (O_1313,N_19713,N_18636);
nor UO_1314 (O_1314,N_18540,N_19818);
or UO_1315 (O_1315,N_18585,N_19322);
nand UO_1316 (O_1316,N_18777,N_18196);
nor UO_1317 (O_1317,N_19786,N_19104);
or UO_1318 (O_1318,N_19052,N_19043);
and UO_1319 (O_1319,N_18845,N_19274);
nand UO_1320 (O_1320,N_19141,N_19363);
and UO_1321 (O_1321,N_18684,N_18148);
nor UO_1322 (O_1322,N_19849,N_19834);
or UO_1323 (O_1323,N_19054,N_19013);
or UO_1324 (O_1324,N_18395,N_19069);
nand UO_1325 (O_1325,N_19857,N_19097);
and UO_1326 (O_1326,N_18281,N_19195);
or UO_1327 (O_1327,N_18158,N_19056);
nor UO_1328 (O_1328,N_18948,N_18747);
or UO_1329 (O_1329,N_19553,N_18683);
nand UO_1330 (O_1330,N_18233,N_19753);
or UO_1331 (O_1331,N_18188,N_19822);
nand UO_1332 (O_1332,N_18554,N_19687);
and UO_1333 (O_1333,N_19692,N_19337);
or UO_1334 (O_1334,N_19302,N_18833);
nand UO_1335 (O_1335,N_18505,N_18909);
nor UO_1336 (O_1336,N_19992,N_18620);
or UO_1337 (O_1337,N_18978,N_18582);
nor UO_1338 (O_1338,N_19004,N_18402);
or UO_1339 (O_1339,N_18984,N_19713);
nand UO_1340 (O_1340,N_18517,N_18280);
and UO_1341 (O_1341,N_18143,N_18548);
or UO_1342 (O_1342,N_19145,N_18135);
nand UO_1343 (O_1343,N_19703,N_18216);
or UO_1344 (O_1344,N_19338,N_19178);
nor UO_1345 (O_1345,N_18311,N_18948);
nor UO_1346 (O_1346,N_19697,N_18435);
nor UO_1347 (O_1347,N_18806,N_18092);
nor UO_1348 (O_1348,N_18439,N_18396);
or UO_1349 (O_1349,N_18134,N_19791);
and UO_1350 (O_1350,N_18167,N_18797);
or UO_1351 (O_1351,N_19160,N_19289);
and UO_1352 (O_1352,N_18889,N_19024);
nand UO_1353 (O_1353,N_19128,N_18415);
nor UO_1354 (O_1354,N_18663,N_18073);
and UO_1355 (O_1355,N_19513,N_18324);
and UO_1356 (O_1356,N_18945,N_18567);
or UO_1357 (O_1357,N_19530,N_19906);
nand UO_1358 (O_1358,N_19292,N_19514);
and UO_1359 (O_1359,N_19745,N_18260);
and UO_1360 (O_1360,N_18103,N_19770);
nor UO_1361 (O_1361,N_18013,N_19182);
nor UO_1362 (O_1362,N_18626,N_18260);
xor UO_1363 (O_1363,N_18004,N_19781);
and UO_1364 (O_1364,N_18406,N_19406);
nand UO_1365 (O_1365,N_19997,N_18973);
nor UO_1366 (O_1366,N_19437,N_19404);
nor UO_1367 (O_1367,N_18930,N_18427);
or UO_1368 (O_1368,N_19692,N_18251);
or UO_1369 (O_1369,N_18688,N_19251);
or UO_1370 (O_1370,N_18581,N_19580);
and UO_1371 (O_1371,N_19087,N_18543);
or UO_1372 (O_1372,N_18255,N_19236);
nand UO_1373 (O_1373,N_18751,N_18767);
or UO_1374 (O_1374,N_19987,N_19716);
nand UO_1375 (O_1375,N_19243,N_19282);
nand UO_1376 (O_1376,N_18982,N_18365);
and UO_1377 (O_1377,N_18923,N_19917);
or UO_1378 (O_1378,N_18343,N_18480);
nor UO_1379 (O_1379,N_19837,N_19552);
and UO_1380 (O_1380,N_19533,N_19045);
nor UO_1381 (O_1381,N_19253,N_18198);
nor UO_1382 (O_1382,N_19800,N_19035);
nand UO_1383 (O_1383,N_19582,N_18559);
and UO_1384 (O_1384,N_19950,N_19237);
nor UO_1385 (O_1385,N_18028,N_19682);
and UO_1386 (O_1386,N_19552,N_18884);
or UO_1387 (O_1387,N_18016,N_19499);
nor UO_1388 (O_1388,N_18310,N_18682);
or UO_1389 (O_1389,N_18146,N_19923);
nor UO_1390 (O_1390,N_18686,N_18308);
or UO_1391 (O_1391,N_18926,N_18173);
nand UO_1392 (O_1392,N_19765,N_19371);
and UO_1393 (O_1393,N_18411,N_19053);
or UO_1394 (O_1394,N_18286,N_19228);
or UO_1395 (O_1395,N_19435,N_19775);
nand UO_1396 (O_1396,N_19274,N_19155);
and UO_1397 (O_1397,N_18659,N_19663);
and UO_1398 (O_1398,N_19238,N_18357);
or UO_1399 (O_1399,N_18794,N_18003);
and UO_1400 (O_1400,N_18701,N_18409);
nor UO_1401 (O_1401,N_19079,N_18856);
and UO_1402 (O_1402,N_19667,N_19796);
and UO_1403 (O_1403,N_18018,N_19342);
nand UO_1404 (O_1404,N_18149,N_19579);
or UO_1405 (O_1405,N_19217,N_18302);
nand UO_1406 (O_1406,N_19404,N_18412);
nor UO_1407 (O_1407,N_18636,N_19864);
nand UO_1408 (O_1408,N_18084,N_19276);
or UO_1409 (O_1409,N_18747,N_19300);
or UO_1410 (O_1410,N_18542,N_18546);
and UO_1411 (O_1411,N_19383,N_19650);
or UO_1412 (O_1412,N_19300,N_19427);
nor UO_1413 (O_1413,N_18853,N_18124);
and UO_1414 (O_1414,N_18954,N_18401);
nor UO_1415 (O_1415,N_19548,N_19539);
or UO_1416 (O_1416,N_18126,N_18789);
nand UO_1417 (O_1417,N_18284,N_18203);
nand UO_1418 (O_1418,N_18275,N_19754);
nand UO_1419 (O_1419,N_18195,N_19394);
nor UO_1420 (O_1420,N_19848,N_19731);
and UO_1421 (O_1421,N_19345,N_19030);
nand UO_1422 (O_1422,N_19752,N_18308);
nand UO_1423 (O_1423,N_18386,N_18393);
or UO_1424 (O_1424,N_18146,N_18781);
nand UO_1425 (O_1425,N_19439,N_18819);
nor UO_1426 (O_1426,N_18131,N_18728);
nand UO_1427 (O_1427,N_18233,N_18594);
nand UO_1428 (O_1428,N_19783,N_19010);
and UO_1429 (O_1429,N_19718,N_18603);
nand UO_1430 (O_1430,N_18954,N_19192);
nor UO_1431 (O_1431,N_19635,N_18332);
nand UO_1432 (O_1432,N_18961,N_18594);
and UO_1433 (O_1433,N_19124,N_18132);
nand UO_1434 (O_1434,N_19616,N_18076);
or UO_1435 (O_1435,N_18075,N_19511);
or UO_1436 (O_1436,N_18650,N_18354);
nand UO_1437 (O_1437,N_19591,N_19572);
nand UO_1438 (O_1438,N_18898,N_19052);
nand UO_1439 (O_1439,N_18336,N_19054);
nand UO_1440 (O_1440,N_18545,N_19243);
nor UO_1441 (O_1441,N_19026,N_19062);
xnor UO_1442 (O_1442,N_19831,N_18150);
nor UO_1443 (O_1443,N_18254,N_19647);
nand UO_1444 (O_1444,N_18269,N_18325);
and UO_1445 (O_1445,N_18236,N_18540);
and UO_1446 (O_1446,N_18442,N_19029);
nand UO_1447 (O_1447,N_18154,N_18874);
nor UO_1448 (O_1448,N_18287,N_19503);
nand UO_1449 (O_1449,N_18387,N_19726);
nor UO_1450 (O_1450,N_19701,N_19590);
or UO_1451 (O_1451,N_18974,N_19692);
or UO_1452 (O_1452,N_18383,N_19117);
or UO_1453 (O_1453,N_18231,N_18775);
nand UO_1454 (O_1454,N_19000,N_19659);
nand UO_1455 (O_1455,N_18501,N_18292);
nor UO_1456 (O_1456,N_18384,N_19059);
nor UO_1457 (O_1457,N_18764,N_19141);
and UO_1458 (O_1458,N_19900,N_19742);
nor UO_1459 (O_1459,N_18284,N_19647);
and UO_1460 (O_1460,N_18984,N_18213);
or UO_1461 (O_1461,N_18027,N_18252);
or UO_1462 (O_1462,N_18865,N_19611);
and UO_1463 (O_1463,N_18593,N_19211);
nor UO_1464 (O_1464,N_19666,N_19644);
nor UO_1465 (O_1465,N_18390,N_18747);
or UO_1466 (O_1466,N_19693,N_18070);
or UO_1467 (O_1467,N_18211,N_19887);
and UO_1468 (O_1468,N_19082,N_19403);
or UO_1469 (O_1469,N_18835,N_19772);
and UO_1470 (O_1470,N_18253,N_19399);
and UO_1471 (O_1471,N_18951,N_18757);
or UO_1472 (O_1472,N_19624,N_18738);
or UO_1473 (O_1473,N_18559,N_19610);
nand UO_1474 (O_1474,N_19464,N_19267);
and UO_1475 (O_1475,N_18043,N_18837);
nand UO_1476 (O_1476,N_19286,N_19014);
nor UO_1477 (O_1477,N_18371,N_18319);
or UO_1478 (O_1478,N_18134,N_19143);
nand UO_1479 (O_1479,N_18075,N_19124);
nand UO_1480 (O_1480,N_18788,N_19947);
and UO_1481 (O_1481,N_19802,N_18560);
or UO_1482 (O_1482,N_18581,N_18342);
or UO_1483 (O_1483,N_18354,N_19507);
nor UO_1484 (O_1484,N_19340,N_19407);
nor UO_1485 (O_1485,N_18213,N_18992);
nor UO_1486 (O_1486,N_19854,N_18491);
nor UO_1487 (O_1487,N_18389,N_19565);
nor UO_1488 (O_1488,N_19966,N_19462);
and UO_1489 (O_1489,N_19723,N_19823);
or UO_1490 (O_1490,N_18498,N_18655);
and UO_1491 (O_1491,N_18027,N_18417);
and UO_1492 (O_1492,N_18797,N_18674);
nor UO_1493 (O_1493,N_19104,N_18781);
and UO_1494 (O_1494,N_18060,N_18401);
and UO_1495 (O_1495,N_19248,N_19714);
and UO_1496 (O_1496,N_18329,N_18910);
and UO_1497 (O_1497,N_19959,N_18050);
and UO_1498 (O_1498,N_18588,N_18445);
nand UO_1499 (O_1499,N_19589,N_19749);
or UO_1500 (O_1500,N_18778,N_19366);
xnor UO_1501 (O_1501,N_19063,N_18255);
and UO_1502 (O_1502,N_19610,N_19533);
nor UO_1503 (O_1503,N_18057,N_18958);
nand UO_1504 (O_1504,N_18657,N_18188);
and UO_1505 (O_1505,N_18441,N_19518);
and UO_1506 (O_1506,N_19061,N_19670);
or UO_1507 (O_1507,N_18028,N_18013);
and UO_1508 (O_1508,N_18311,N_18321);
and UO_1509 (O_1509,N_19415,N_18650);
and UO_1510 (O_1510,N_18270,N_19489);
or UO_1511 (O_1511,N_19763,N_19060);
nand UO_1512 (O_1512,N_18641,N_19339);
or UO_1513 (O_1513,N_18786,N_18518);
or UO_1514 (O_1514,N_19470,N_18516);
nor UO_1515 (O_1515,N_18919,N_18574);
nor UO_1516 (O_1516,N_18862,N_18020);
nor UO_1517 (O_1517,N_19771,N_19130);
and UO_1518 (O_1518,N_19361,N_19959);
nand UO_1519 (O_1519,N_18947,N_18185);
nand UO_1520 (O_1520,N_18295,N_18424);
nand UO_1521 (O_1521,N_18108,N_18592);
nand UO_1522 (O_1522,N_18070,N_18863);
nand UO_1523 (O_1523,N_19622,N_19299);
nor UO_1524 (O_1524,N_18431,N_18433);
or UO_1525 (O_1525,N_18952,N_18423);
and UO_1526 (O_1526,N_19475,N_19626);
or UO_1527 (O_1527,N_18619,N_18288);
and UO_1528 (O_1528,N_18715,N_19656);
nor UO_1529 (O_1529,N_19277,N_19544);
nand UO_1530 (O_1530,N_19231,N_19526);
or UO_1531 (O_1531,N_19963,N_19115);
and UO_1532 (O_1532,N_19785,N_19701);
nand UO_1533 (O_1533,N_18431,N_18764);
or UO_1534 (O_1534,N_19630,N_18878);
or UO_1535 (O_1535,N_18692,N_19846);
nand UO_1536 (O_1536,N_18251,N_18454);
nor UO_1537 (O_1537,N_18961,N_19367);
nor UO_1538 (O_1538,N_18026,N_18422);
and UO_1539 (O_1539,N_19447,N_18557);
nor UO_1540 (O_1540,N_19788,N_19330);
or UO_1541 (O_1541,N_19902,N_18060);
or UO_1542 (O_1542,N_18921,N_18919);
or UO_1543 (O_1543,N_18654,N_18348);
and UO_1544 (O_1544,N_19168,N_18588);
and UO_1545 (O_1545,N_19004,N_18202);
nor UO_1546 (O_1546,N_19230,N_18581);
and UO_1547 (O_1547,N_18015,N_18285);
nor UO_1548 (O_1548,N_19729,N_19488);
nand UO_1549 (O_1549,N_18067,N_18136);
or UO_1550 (O_1550,N_19166,N_18006);
nand UO_1551 (O_1551,N_19337,N_19327);
nand UO_1552 (O_1552,N_19731,N_18620);
or UO_1553 (O_1553,N_19191,N_18349);
nor UO_1554 (O_1554,N_18456,N_19956);
nand UO_1555 (O_1555,N_18661,N_19646);
nand UO_1556 (O_1556,N_18312,N_19864);
or UO_1557 (O_1557,N_19932,N_18717);
and UO_1558 (O_1558,N_18874,N_18160);
nor UO_1559 (O_1559,N_18402,N_18740);
and UO_1560 (O_1560,N_19033,N_18832);
nand UO_1561 (O_1561,N_18072,N_19974);
nand UO_1562 (O_1562,N_19822,N_18313);
or UO_1563 (O_1563,N_18053,N_18312);
nand UO_1564 (O_1564,N_18725,N_18379);
or UO_1565 (O_1565,N_18055,N_19477);
nand UO_1566 (O_1566,N_18989,N_18747);
or UO_1567 (O_1567,N_19576,N_19473);
and UO_1568 (O_1568,N_19423,N_18111);
and UO_1569 (O_1569,N_18401,N_18399);
or UO_1570 (O_1570,N_18830,N_19323);
nor UO_1571 (O_1571,N_18543,N_19332);
or UO_1572 (O_1572,N_19233,N_19783);
or UO_1573 (O_1573,N_18474,N_18495);
nand UO_1574 (O_1574,N_19340,N_19217);
and UO_1575 (O_1575,N_19096,N_18242);
and UO_1576 (O_1576,N_18162,N_18937);
nand UO_1577 (O_1577,N_18861,N_18429);
nand UO_1578 (O_1578,N_19047,N_19212);
nand UO_1579 (O_1579,N_18079,N_18962);
or UO_1580 (O_1580,N_18640,N_18370);
or UO_1581 (O_1581,N_19186,N_19778);
or UO_1582 (O_1582,N_19202,N_18055);
nand UO_1583 (O_1583,N_19149,N_19974);
nand UO_1584 (O_1584,N_19082,N_19191);
nand UO_1585 (O_1585,N_18255,N_18653);
and UO_1586 (O_1586,N_19758,N_18390);
or UO_1587 (O_1587,N_19833,N_18102);
or UO_1588 (O_1588,N_18091,N_19100);
nor UO_1589 (O_1589,N_18753,N_18621);
or UO_1590 (O_1590,N_19668,N_18553);
and UO_1591 (O_1591,N_18784,N_19876);
xnor UO_1592 (O_1592,N_19429,N_18043);
nand UO_1593 (O_1593,N_18996,N_19903);
nand UO_1594 (O_1594,N_18312,N_19291);
nor UO_1595 (O_1595,N_18494,N_18436);
nor UO_1596 (O_1596,N_19948,N_19960);
nor UO_1597 (O_1597,N_18079,N_19743);
or UO_1598 (O_1598,N_18828,N_18987);
nor UO_1599 (O_1599,N_18788,N_18285);
or UO_1600 (O_1600,N_18759,N_18625);
and UO_1601 (O_1601,N_19022,N_18641);
and UO_1602 (O_1602,N_19387,N_19393);
or UO_1603 (O_1603,N_19998,N_19128);
nor UO_1604 (O_1604,N_19907,N_19255);
nor UO_1605 (O_1605,N_19640,N_19898);
nor UO_1606 (O_1606,N_19975,N_19421);
nor UO_1607 (O_1607,N_18457,N_18705);
or UO_1608 (O_1608,N_19955,N_18504);
or UO_1609 (O_1609,N_19210,N_18593);
nand UO_1610 (O_1610,N_19179,N_19787);
nor UO_1611 (O_1611,N_18760,N_19276);
xnor UO_1612 (O_1612,N_19918,N_18644);
nand UO_1613 (O_1613,N_19734,N_18785);
or UO_1614 (O_1614,N_18077,N_19476);
or UO_1615 (O_1615,N_19846,N_18798);
nand UO_1616 (O_1616,N_19112,N_19614);
and UO_1617 (O_1617,N_19664,N_18407);
nor UO_1618 (O_1618,N_19526,N_19451);
and UO_1619 (O_1619,N_18401,N_18700);
or UO_1620 (O_1620,N_18800,N_18771);
nand UO_1621 (O_1621,N_18309,N_19278);
and UO_1622 (O_1622,N_19220,N_19259);
nor UO_1623 (O_1623,N_18372,N_19732);
and UO_1624 (O_1624,N_19172,N_19504);
and UO_1625 (O_1625,N_18201,N_19885);
nand UO_1626 (O_1626,N_19605,N_19881);
or UO_1627 (O_1627,N_19081,N_19082);
or UO_1628 (O_1628,N_19595,N_19816);
nor UO_1629 (O_1629,N_18343,N_18342);
nor UO_1630 (O_1630,N_18710,N_19504);
nand UO_1631 (O_1631,N_18173,N_19154);
and UO_1632 (O_1632,N_19892,N_18706);
and UO_1633 (O_1633,N_18237,N_19080);
and UO_1634 (O_1634,N_19572,N_19163);
and UO_1635 (O_1635,N_19395,N_19906);
nand UO_1636 (O_1636,N_19298,N_18537);
and UO_1637 (O_1637,N_18522,N_19505);
and UO_1638 (O_1638,N_18673,N_18727);
nand UO_1639 (O_1639,N_19018,N_18580);
or UO_1640 (O_1640,N_19954,N_18465);
or UO_1641 (O_1641,N_19489,N_18822);
nor UO_1642 (O_1642,N_18715,N_19645);
or UO_1643 (O_1643,N_19199,N_18829);
and UO_1644 (O_1644,N_18304,N_18547);
nor UO_1645 (O_1645,N_18078,N_19264);
nor UO_1646 (O_1646,N_18622,N_18408);
nand UO_1647 (O_1647,N_19897,N_18709);
or UO_1648 (O_1648,N_18638,N_19424);
or UO_1649 (O_1649,N_18066,N_18216);
nor UO_1650 (O_1650,N_18913,N_18292);
nor UO_1651 (O_1651,N_19508,N_18857);
and UO_1652 (O_1652,N_18043,N_19996);
nand UO_1653 (O_1653,N_19299,N_19014);
or UO_1654 (O_1654,N_18657,N_19406);
nand UO_1655 (O_1655,N_19198,N_19918);
nand UO_1656 (O_1656,N_18045,N_18135);
or UO_1657 (O_1657,N_18207,N_19649);
and UO_1658 (O_1658,N_18145,N_19496);
nand UO_1659 (O_1659,N_19295,N_18873);
or UO_1660 (O_1660,N_18845,N_18524);
or UO_1661 (O_1661,N_19730,N_19049);
or UO_1662 (O_1662,N_18982,N_19735);
and UO_1663 (O_1663,N_18784,N_19505);
or UO_1664 (O_1664,N_18501,N_19595);
nor UO_1665 (O_1665,N_19269,N_18216);
or UO_1666 (O_1666,N_18330,N_19720);
and UO_1667 (O_1667,N_19468,N_18281);
nand UO_1668 (O_1668,N_19317,N_19113);
and UO_1669 (O_1669,N_18749,N_19005);
and UO_1670 (O_1670,N_18668,N_19176);
and UO_1671 (O_1671,N_19145,N_18916);
and UO_1672 (O_1672,N_18246,N_19535);
or UO_1673 (O_1673,N_18536,N_19049);
or UO_1674 (O_1674,N_18378,N_19871);
xnor UO_1675 (O_1675,N_18802,N_18699);
and UO_1676 (O_1676,N_18621,N_19886);
or UO_1677 (O_1677,N_19170,N_19154);
or UO_1678 (O_1678,N_18724,N_18586);
nand UO_1679 (O_1679,N_18619,N_18376);
nand UO_1680 (O_1680,N_18179,N_19190);
and UO_1681 (O_1681,N_19603,N_18214);
nor UO_1682 (O_1682,N_19785,N_19890);
nor UO_1683 (O_1683,N_18796,N_18167);
nand UO_1684 (O_1684,N_18965,N_19734);
nand UO_1685 (O_1685,N_18668,N_19261);
nand UO_1686 (O_1686,N_19537,N_19569);
nor UO_1687 (O_1687,N_19425,N_19677);
or UO_1688 (O_1688,N_18863,N_18271);
or UO_1689 (O_1689,N_19058,N_18407);
nor UO_1690 (O_1690,N_19207,N_18710);
nand UO_1691 (O_1691,N_18539,N_19926);
nor UO_1692 (O_1692,N_19796,N_18164);
nand UO_1693 (O_1693,N_18038,N_18229);
or UO_1694 (O_1694,N_18644,N_18045);
nand UO_1695 (O_1695,N_19777,N_18795);
nand UO_1696 (O_1696,N_18101,N_18488);
and UO_1697 (O_1697,N_18982,N_18762);
nor UO_1698 (O_1698,N_19710,N_18930);
nand UO_1699 (O_1699,N_19863,N_18592);
nand UO_1700 (O_1700,N_18304,N_18092);
and UO_1701 (O_1701,N_19880,N_19196);
and UO_1702 (O_1702,N_18873,N_19585);
or UO_1703 (O_1703,N_19840,N_19690);
and UO_1704 (O_1704,N_19998,N_18534);
nor UO_1705 (O_1705,N_18948,N_19838);
and UO_1706 (O_1706,N_18348,N_19724);
nor UO_1707 (O_1707,N_19976,N_19445);
nor UO_1708 (O_1708,N_18844,N_18905);
nand UO_1709 (O_1709,N_18635,N_18515);
or UO_1710 (O_1710,N_19021,N_19412);
or UO_1711 (O_1711,N_19067,N_18550);
nand UO_1712 (O_1712,N_18614,N_18269);
and UO_1713 (O_1713,N_19368,N_18004);
and UO_1714 (O_1714,N_19999,N_19804);
or UO_1715 (O_1715,N_18868,N_18769);
or UO_1716 (O_1716,N_18400,N_18300);
and UO_1717 (O_1717,N_18852,N_19579);
nand UO_1718 (O_1718,N_19634,N_18533);
or UO_1719 (O_1719,N_18897,N_18636);
and UO_1720 (O_1720,N_18209,N_18621);
nand UO_1721 (O_1721,N_18367,N_19787);
nor UO_1722 (O_1722,N_18241,N_18373);
and UO_1723 (O_1723,N_18150,N_18015);
and UO_1724 (O_1724,N_19397,N_18623);
or UO_1725 (O_1725,N_18793,N_19782);
nand UO_1726 (O_1726,N_18620,N_18710);
nor UO_1727 (O_1727,N_18613,N_18853);
or UO_1728 (O_1728,N_19109,N_19489);
nand UO_1729 (O_1729,N_18941,N_18239);
nand UO_1730 (O_1730,N_18399,N_18587);
nor UO_1731 (O_1731,N_19022,N_18432);
nor UO_1732 (O_1732,N_18973,N_18317);
and UO_1733 (O_1733,N_19933,N_18522);
nor UO_1734 (O_1734,N_18851,N_19623);
nand UO_1735 (O_1735,N_18723,N_19124);
nor UO_1736 (O_1736,N_19663,N_18353);
nand UO_1737 (O_1737,N_19131,N_18975);
nor UO_1738 (O_1738,N_18082,N_18225);
and UO_1739 (O_1739,N_19428,N_18655);
and UO_1740 (O_1740,N_18521,N_19424);
or UO_1741 (O_1741,N_19678,N_18825);
or UO_1742 (O_1742,N_19655,N_18129);
and UO_1743 (O_1743,N_18775,N_19093);
xnor UO_1744 (O_1744,N_18870,N_18815);
nand UO_1745 (O_1745,N_18570,N_18042);
nand UO_1746 (O_1746,N_19944,N_18920);
nor UO_1747 (O_1747,N_19005,N_19927);
or UO_1748 (O_1748,N_19040,N_19740);
and UO_1749 (O_1749,N_18910,N_18135);
or UO_1750 (O_1750,N_19481,N_19104);
or UO_1751 (O_1751,N_18069,N_18352);
nor UO_1752 (O_1752,N_18916,N_18413);
nor UO_1753 (O_1753,N_19162,N_19256);
or UO_1754 (O_1754,N_19404,N_19230);
and UO_1755 (O_1755,N_18748,N_19244);
nand UO_1756 (O_1756,N_18821,N_19230);
and UO_1757 (O_1757,N_18469,N_19730);
and UO_1758 (O_1758,N_19818,N_19699);
nor UO_1759 (O_1759,N_18041,N_18363);
nor UO_1760 (O_1760,N_19010,N_19641);
or UO_1761 (O_1761,N_19860,N_18668);
or UO_1762 (O_1762,N_19450,N_18181);
nand UO_1763 (O_1763,N_18935,N_19582);
and UO_1764 (O_1764,N_18879,N_18498);
or UO_1765 (O_1765,N_18764,N_19314);
nand UO_1766 (O_1766,N_19239,N_18212);
and UO_1767 (O_1767,N_19185,N_19308);
nor UO_1768 (O_1768,N_19361,N_19631);
and UO_1769 (O_1769,N_19746,N_19700);
and UO_1770 (O_1770,N_18942,N_18284);
or UO_1771 (O_1771,N_19584,N_18127);
or UO_1772 (O_1772,N_19690,N_19616);
nand UO_1773 (O_1773,N_19376,N_19394);
or UO_1774 (O_1774,N_18164,N_19133);
or UO_1775 (O_1775,N_19539,N_19330);
and UO_1776 (O_1776,N_19615,N_19813);
nor UO_1777 (O_1777,N_19009,N_18816);
and UO_1778 (O_1778,N_19675,N_19007);
nor UO_1779 (O_1779,N_18154,N_18718);
nor UO_1780 (O_1780,N_19371,N_19900);
and UO_1781 (O_1781,N_18768,N_18478);
nand UO_1782 (O_1782,N_19615,N_19522);
nor UO_1783 (O_1783,N_18745,N_18294);
nand UO_1784 (O_1784,N_19379,N_19620);
nor UO_1785 (O_1785,N_18297,N_18607);
nor UO_1786 (O_1786,N_19439,N_19494);
or UO_1787 (O_1787,N_19294,N_19259);
nand UO_1788 (O_1788,N_19701,N_19186);
or UO_1789 (O_1789,N_19366,N_19936);
nand UO_1790 (O_1790,N_19215,N_19892);
or UO_1791 (O_1791,N_19822,N_18149);
and UO_1792 (O_1792,N_19665,N_19788);
and UO_1793 (O_1793,N_19061,N_18062);
nor UO_1794 (O_1794,N_18865,N_18008);
and UO_1795 (O_1795,N_19233,N_19968);
and UO_1796 (O_1796,N_18727,N_18468);
or UO_1797 (O_1797,N_19865,N_18455);
and UO_1798 (O_1798,N_18438,N_19776);
and UO_1799 (O_1799,N_18463,N_19794);
and UO_1800 (O_1800,N_19111,N_19670);
nor UO_1801 (O_1801,N_19480,N_19052);
nand UO_1802 (O_1802,N_19941,N_19859);
nand UO_1803 (O_1803,N_19510,N_18104);
and UO_1804 (O_1804,N_19852,N_18001);
or UO_1805 (O_1805,N_18294,N_18637);
and UO_1806 (O_1806,N_19398,N_19360);
and UO_1807 (O_1807,N_18395,N_18787);
nand UO_1808 (O_1808,N_18822,N_19165);
and UO_1809 (O_1809,N_19734,N_18228);
or UO_1810 (O_1810,N_19618,N_18773);
and UO_1811 (O_1811,N_18441,N_18615);
or UO_1812 (O_1812,N_19007,N_18796);
nor UO_1813 (O_1813,N_19634,N_19206);
nand UO_1814 (O_1814,N_18615,N_18085);
nor UO_1815 (O_1815,N_18059,N_18312);
or UO_1816 (O_1816,N_18824,N_18246);
nand UO_1817 (O_1817,N_19356,N_18887);
nand UO_1818 (O_1818,N_18547,N_18132);
or UO_1819 (O_1819,N_19867,N_19345);
nor UO_1820 (O_1820,N_19935,N_18386);
nand UO_1821 (O_1821,N_18661,N_18233);
nor UO_1822 (O_1822,N_18375,N_19088);
nor UO_1823 (O_1823,N_19528,N_18619);
and UO_1824 (O_1824,N_19680,N_18159);
and UO_1825 (O_1825,N_19255,N_19316);
nand UO_1826 (O_1826,N_19576,N_18279);
nor UO_1827 (O_1827,N_19975,N_18519);
and UO_1828 (O_1828,N_19285,N_18687);
or UO_1829 (O_1829,N_18471,N_19489);
nor UO_1830 (O_1830,N_18485,N_18273);
or UO_1831 (O_1831,N_19026,N_19319);
and UO_1832 (O_1832,N_18927,N_19651);
nor UO_1833 (O_1833,N_19074,N_18162);
or UO_1834 (O_1834,N_19859,N_19479);
nand UO_1835 (O_1835,N_18747,N_19880);
or UO_1836 (O_1836,N_18383,N_18139);
and UO_1837 (O_1837,N_18897,N_18834);
and UO_1838 (O_1838,N_18366,N_18044);
nand UO_1839 (O_1839,N_18641,N_18058);
or UO_1840 (O_1840,N_18509,N_18451);
and UO_1841 (O_1841,N_18254,N_18556);
nor UO_1842 (O_1842,N_19644,N_19533);
nor UO_1843 (O_1843,N_19413,N_18969);
and UO_1844 (O_1844,N_19853,N_18351);
nor UO_1845 (O_1845,N_19877,N_19797);
nand UO_1846 (O_1846,N_19481,N_18517);
and UO_1847 (O_1847,N_18822,N_18430);
nor UO_1848 (O_1848,N_18771,N_19541);
and UO_1849 (O_1849,N_18702,N_19584);
nor UO_1850 (O_1850,N_19174,N_18973);
nor UO_1851 (O_1851,N_19207,N_18495);
and UO_1852 (O_1852,N_19756,N_18538);
and UO_1853 (O_1853,N_19198,N_19701);
or UO_1854 (O_1854,N_19745,N_18280);
or UO_1855 (O_1855,N_18273,N_18449);
or UO_1856 (O_1856,N_18923,N_18529);
or UO_1857 (O_1857,N_19412,N_19117);
nor UO_1858 (O_1858,N_18213,N_18462);
or UO_1859 (O_1859,N_18640,N_18210);
nand UO_1860 (O_1860,N_19312,N_19219);
nand UO_1861 (O_1861,N_19008,N_18443);
and UO_1862 (O_1862,N_19018,N_18573);
nor UO_1863 (O_1863,N_19711,N_19463);
and UO_1864 (O_1864,N_18131,N_19521);
nor UO_1865 (O_1865,N_19702,N_18291);
nor UO_1866 (O_1866,N_19684,N_18042);
or UO_1867 (O_1867,N_19229,N_18392);
or UO_1868 (O_1868,N_19474,N_18930);
nand UO_1869 (O_1869,N_18443,N_18754);
nand UO_1870 (O_1870,N_19251,N_19195);
nor UO_1871 (O_1871,N_18523,N_18304);
nand UO_1872 (O_1872,N_19072,N_19877);
or UO_1873 (O_1873,N_18274,N_18170);
and UO_1874 (O_1874,N_19863,N_18808);
and UO_1875 (O_1875,N_19905,N_19718);
nand UO_1876 (O_1876,N_19447,N_19605);
or UO_1877 (O_1877,N_19586,N_18276);
nand UO_1878 (O_1878,N_18566,N_18479);
or UO_1879 (O_1879,N_19026,N_18326);
nor UO_1880 (O_1880,N_18045,N_19717);
or UO_1881 (O_1881,N_19598,N_18028);
and UO_1882 (O_1882,N_19508,N_19601);
or UO_1883 (O_1883,N_19669,N_18579);
and UO_1884 (O_1884,N_18899,N_19996);
and UO_1885 (O_1885,N_18475,N_18894);
and UO_1886 (O_1886,N_19379,N_18138);
or UO_1887 (O_1887,N_19595,N_18655);
nor UO_1888 (O_1888,N_19804,N_18012);
or UO_1889 (O_1889,N_18063,N_19306);
and UO_1890 (O_1890,N_19111,N_18041);
or UO_1891 (O_1891,N_18332,N_18508);
or UO_1892 (O_1892,N_19791,N_18364);
and UO_1893 (O_1893,N_19614,N_19434);
or UO_1894 (O_1894,N_19742,N_18119);
nand UO_1895 (O_1895,N_18435,N_18820);
nor UO_1896 (O_1896,N_19749,N_19322);
nor UO_1897 (O_1897,N_19328,N_19865);
and UO_1898 (O_1898,N_19601,N_19274);
nand UO_1899 (O_1899,N_19847,N_19067);
and UO_1900 (O_1900,N_19765,N_19894);
and UO_1901 (O_1901,N_19048,N_19880);
or UO_1902 (O_1902,N_19000,N_18750);
nor UO_1903 (O_1903,N_19993,N_18219);
and UO_1904 (O_1904,N_18380,N_19694);
nand UO_1905 (O_1905,N_19092,N_19602);
or UO_1906 (O_1906,N_19460,N_19827);
and UO_1907 (O_1907,N_18996,N_18377);
xnor UO_1908 (O_1908,N_18357,N_18235);
nor UO_1909 (O_1909,N_19616,N_19860);
nor UO_1910 (O_1910,N_19121,N_19832);
or UO_1911 (O_1911,N_19792,N_18557);
nor UO_1912 (O_1912,N_18736,N_19079);
nor UO_1913 (O_1913,N_19751,N_19019);
and UO_1914 (O_1914,N_18068,N_18843);
nor UO_1915 (O_1915,N_19174,N_19530);
nand UO_1916 (O_1916,N_19476,N_19432);
and UO_1917 (O_1917,N_18374,N_19258);
or UO_1918 (O_1918,N_19187,N_19138);
nor UO_1919 (O_1919,N_19057,N_18502);
and UO_1920 (O_1920,N_18401,N_19052);
nand UO_1921 (O_1921,N_19789,N_18898);
or UO_1922 (O_1922,N_18541,N_19479);
and UO_1923 (O_1923,N_18356,N_19416);
nand UO_1924 (O_1924,N_18623,N_19390);
and UO_1925 (O_1925,N_19715,N_19447);
or UO_1926 (O_1926,N_19404,N_19972);
and UO_1927 (O_1927,N_19655,N_18851);
nand UO_1928 (O_1928,N_18478,N_18764);
nand UO_1929 (O_1929,N_18038,N_18090);
nand UO_1930 (O_1930,N_18362,N_19913);
nor UO_1931 (O_1931,N_19361,N_18704);
or UO_1932 (O_1932,N_18247,N_19186);
and UO_1933 (O_1933,N_19013,N_19850);
nand UO_1934 (O_1934,N_19125,N_19414);
nand UO_1935 (O_1935,N_18176,N_18521);
xor UO_1936 (O_1936,N_19347,N_18702);
nor UO_1937 (O_1937,N_18547,N_19821);
and UO_1938 (O_1938,N_19615,N_19018);
or UO_1939 (O_1939,N_18911,N_19088);
or UO_1940 (O_1940,N_19987,N_18985);
and UO_1941 (O_1941,N_19149,N_19611);
nor UO_1942 (O_1942,N_18466,N_19996);
or UO_1943 (O_1943,N_18388,N_19033);
or UO_1944 (O_1944,N_18331,N_18673);
nor UO_1945 (O_1945,N_18457,N_19343);
and UO_1946 (O_1946,N_18172,N_18385);
nor UO_1947 (O_1947,N_19400,N_19765);
nand UO_1948 (O_1948,N_18881,N_18197);
nand UO_1949 (O_1949,N_19116,N_19537);
and UO_1950 (O_1950,N_19729,N_18590);
and UO_1951 (O_1951,N_18569,N_18886);
nor UO_1952 (O_1952,N_19522,N_18118);
nor UO_1953 (O_1953,N_18293,N_18160);
and UO_1954 (O_1954,N_18252,N_18696);
or UO_1955 (O_1955,N_18405,N_19566);
nand UO_1956 (O_1956,N_18223,N_18422);
xnor UO_1957 (O_1957,N_18442,N_19526);
nand UO_1958 (O_1958,N_19121,N_19421);
or UO_1959 (O_1959,N_19584,N_19579);
and UO_1960 (O_1960,N_19855,N_18187);
nor UO_1961 (O_1961,N_19623,N_19671);
nor UO_1962 (O_1962,N_18397,N_19302);
and UO_1963 (O_1963,N_18802,N_19567);
or UO_1964 (O_1964,N_19385,N_19045);
and UO_1965 (O_1965,N_18702,N_18809);
nor UO_1966 (O_1966,N_19964,N_18291);
or UO_1967 (O_1967,N_18056,N_19514);
nor UO_1968 (O_1968,N_19787,N_19570);
nor UO_1969 (O_1969,N_18338,N_19902);
and UO_1970 (O_1970,N_19439,N_19941);
nand UO_1971 (O_1971,N_19907,N_18662);
or UO_1972 (O_1972,N_19404,N_18965);
or UO_1973 (O_1973,N_18958,N_18279);
or UO_1974 (O_1974,N_19316,N_19413);
nor UO_1975 (O_1975,N_19285,N_19618);
nand UO_1976 (O_1976,N_19978,N_18858);
nand UO_1977 (O_1977,N_19820,N_19827);
nor UO_1978 (O_1978,N_19242,N_18606);
nor UO_1979 (O_1979,N_18141,N_19024);
and UO_1980 (O_1980,N_18819,N_18578);
and UO_1981 (O_1981,N_19532,N_18790);
or UO_1982 (O_1982,N_18841,N_18595);
nand UO_1983 (O_1983,N_18142,N_19332);
nor UO_1984 (O_1984,N_18677,N_19622);
or UO_1985 (O_1985,N_18130,N_19419);
nand UO_1986 (O_1986,N_18643,N_18981);
nor UO_1987 (O_1987,N_19760,N_19591);
nor UO_1988 (O_1988,N_18446,N_19693);
nor UO_1989 (O_1989,N_18681,N_18578);
or UO_1990 (O_1990,N_19239,N_18747);
nor UO_1991 (O_1991,N_18425,N_19876);
nand UO_1992 (O_1992,N_19601,N_18489);
or UO_1993 (O_1993,N_19351,N_19430);
nand UO_1994 (O_1994,N_19734,N_19492);
nand UO_1995 (O_1995,N_18267,N_18192);
and UO_1996 (O_1996,N_19134,N_19648);
nor UO_1997 (O_1997,N_18099,N_18360);
nand UO_1998 (O_1998,N_18128,N_19610);
nand UO_1999 (O_1999,N_19556,N_19910);
xor UO_2000 (O_2000,N_19019,N_19911);
nor UO_2001 (O_2001,N_18243,N_18898);
or UO_2002 (O_2002,N_18487,N_18627);
and UO_2003 (O_2003,N_19897,N_18938);
or UO_2004 (O_2004,N_19497,N_19390);
and UO_2005 (O_2005,N_18113,N_18293);
nand UO_2006 (O_2006,N_19688,N_19870);
and UO_2007 (O_2007,N_19028,N_19073);
and UO_2008 (O_2008,N_19451,N_18171);
and UO_2009 (O_2009,N_19564,N_18407);
nand UO_2010 (O_2010,N_19413,N_19444);
or UO_2011 (O_2011,N_18896,N_19586);
nor UO_2012 (O_2012,N_19705,N_18327);
xnor UO_2013 (O_2013,N_19935,N_19834);
and UO_2014 (O_2014,N_18010,N_18852);
nand UO_2015 (O_2015,N_19905,N_19850);
nor UO_2016 (O_2016,N_18014,N_18835);
nor UO_2017 (O_2017,N_19996,N_18915);
nor UO_2018 (O_2018,N_18113,N_18116);
or UO_2019 (O_2019,N_18752,N_19335);
and UO_2020 (O_2020,N_18212,N_19548);
nand UO_2021 (O_2021,N_18973,N_18250);
nand UO_2022 (O_2022,N_18059,N_19091);
or UO_2023 (O_2023,N_18989,N_18532);
nor UO_2024 (O_2024,N_19144,N_18560);
nand UO_2025 (O_2025,N_18423,N_19935);
nor UO_2026 (O_2026,N_18366,N_19265);
and UO_2027 (O_2027,N_18046,N_19812);
or UO_2028 (O_2028,N_18034,N_19999);
or UO_2029 (O_2029,N_19198,N_18068);
or UO_2030 (O_2030,N_18381,N_18290);
or UO_2031 (O_2031,N_18746,N_18631);
nor UO_2032 (O_2032,N_18873,N_19368);
nand UO_2033 (O_2033,N_18068,N_18367);
nor UO_2034 (O_2034,N_18544,N_18312);
and UO_2035 (O_2035,N_19090,N_18524);
nor UO_2036 (O_2036,N_19519,N_19389);
nand UO_2037 (O_2037,N_19761,N_19174);
and UO_2038 (O_2038,N_18744,N_18481);
and UO_2039 (O_2039,N_18484,N_19570);
nand UO_2040 (O_2040,N_19605,N_19649);
nor UO_2041 (O_2041,N_18885,N_19940);
and UO_2042 (O_2042,N_18047,N_18652);
nand UO_2043 (O_2043,N_19291,N_19518);
nor UO_2044 (O_2044,N_19991,N_18063);
and UO_2045 (O_2045,N_18704,N_18896);
nand UO_2046 (O_2046,N_18491,N_18577);
or UO_2047 (O_2047,N_19152,N_18015);
and UO_2048 (O_2048,N_18933,N_19649);
nand UO_2049 (O_2049,N_18559,N_19081);
and UO_2050 (O_2050,N_18975,N_18728);
and UO_2051 (O_2051,N_19038,N_18299);
and UO_2052 (O_2052,N_19359,N_18262);
nand UO_2053 (O_2053,N_18817,N_18351);
or UO_2054 (O_2054,N_19199,N_19030);
and UO_2055 (O_2055,N_19132,N_19764);
or UO_2056 (O_2056,N_18415,N_19825);
nand UO_2057 (O_2057,N_18124,N_18793);
nand UO_2058 (O_2058,N_18838,N_18590);
nand UO_2059 (O_2059,N_19822,N_19185);
and UO_2060 (O_2060,N_18848,N_18573);
and UO_2061 (O_2061,N_19991,N_19455);
or UO_2062 (O_2062,N_19152,N_19537);
nand UO_2063 (O_2063,N_18090,N_19633);
or UO_2064 (O_2064,N_19840,N_18894);
or UO_2065 (O_2065,N_18486,N_19921);
nand UO_2066 (O_2066,N_18485,N_19667);
and UO_2067 (O_2067,N_19635,N_19906);
or UO_2068 (O_2068,N_18554,N_19192);
or UO_2069 (O_2069,N_19506,N_18285);
and UO_2070 (O_2070,N_18026,N_18354);
and UO_2071 (O_2071,N_18153,N_19812);
nor UO_2072 (O_2072,N_19658,N_19839);
nand UO_2073 (O_2073,N_18953,N_18268);
nand UO_2074 (O_2074,N_19062,N_19247);
nor UO_2075 (O_2075,N_19922,N_18340);
or UO_2076 (O_2076,N_19486,N_19014);
or UO_2077 (O_2077,N_19319,N_18009);
and UO_2078 (O_2078,N_19634,N_18435);
nand UO_2079 (O_2079,N_19671,N_19480);
nand UO_2080 (O_2080,N_18667,N_18523);
nand UO_2081 (O_2081,N_19762,N_19883);
nor UO_2082 (O_2082,N_19850,N_19112);
nand UO_2083 (O_2083,N_18565,N_19184);
nor UO_2084 (O_2084,N_19501,N_18680);
nor UO_2085 (O_2085,N_19329,N_18149);
or UO_2086 (O_2086,N_19232,N_19383);
nand UO_2087 (O_2087,N_18264,N_19574);
nor UO_2088 (O_2088,N_19022,N_19628);
nor UO_2089 (O_2089,N_19191,N_18179);
or UO_2090 (O_2090,N_18885,N_19737);
xor UO_2091 (O_2091,N_19075,N_18009);
and UO_2092 (O_2092,N_18153,N_18277);
nor UO_2093 (O_2093,N_19644,N_19435);
nand UO_2094 (O_2094,N_19098,N_18686);
or UO_2095 (O_2095,N_19133,N_18191);
nand UO_2096 (O_2096,N_19494,N_18358);
or UO_2097 (O_2097,N_18318,N_19414);
or UO_2098 (O_2098,N_19477,N_18983);
and UO_2099 (O_2099,N_19188,N_18763);
nor UO_2100 (O_2100,N_18152,N_18582);
or UO_2101 (O_2101,N_19613,N_18966);
and UO_2102 (O_2102,N_18575,N_19365);
nor UO_2103 (O_2103,N_19605,N_18692);
nor UO_2104 (O_2104,N_19304,N_18739);
nor UO_2105 (O_2105,N_19073,N_18802);
nand UO_2106 (O_2106,N_18144,N_19508);
nand UO_2107 (O_2107,N_19079,N_19571);
nor UO_2108 (O_2108,N_18763,N_18072);
nand UO_2109 (O_2109,N_18378,N_18835);
nor UO_2110 (O_2110,N_18315,N_18336);
nor UO_2111 (O_2111,N_18800,N_18004);
or UO_2112 (O_2112,N_18319,N_18456);
nor UO_2113 (O_2113,N_18343,N_19514);
nand UO_2114 (O_2114,N_19279,N_19148);
and UO_2115 (O_2115,N_19917,N_18196);
nand UO_2116 (O_2116,N_19833,N_19180);
nand UO_2117 (O_2117,N_18529,N_18513);
nand UO_2118 (O_2118,N_18937,N_19573);
nor UO_2119 (O_2119,N_18171,N_19001);
and UO_2120 (O_2120,N_18651,N_19566);
nand UO_2121 (O_2121,N_19042,N_18541);
and UO_2122 (O_2122,N_18449,N_19362);
nor UO_2123 (O_2123,N_18539,N_18728);
or UO_2124 (O_2124,N_18927,N_18678);
nor UO_2125 (O_2125,N_19234,N_18264);
and UO_2126 (O_2126,N_19534,N_18322);
nor UO_2127 (O_2127,N_19096,N_19109);
nand UO_2128 (O_2128,N_19270,N_19602);
nor UO_2129 (O_2129,N_19528,N_18569);
nand UO_2130 (O_2130,N_18590,N_18367);
or UO_2131 (O_2131,N_18656,N_18806);
xnor UO_2132 (O_2132,N_18152,N_19741);
nand UO_2133 (O_2133,N_19484,N_19885);
or UO_2134 (O_2134,N_19458,N_19440);
nand UO_2135 (O_2135,N_19788,N_19447);
nand UO_2136 (O_2136,N_19727,N_19840);
or UO_2137 (O_2137,N_19284,N_18066);
nand UO_2138 (O_2138,N_18589,N_19034);
nand UO_2139 (O_2139,N_18092,N_18142);
nand UO_2140 (O_2140,N_18861,N_19869);
nor UO_2141 (O_2141,N_19334,N_18245);
or UO_2142 (O_2142,N_18730,N_19594);
nand UO_2143 (O_2143,N_19257,N_19668);
nor UO_2144 (O_2144,N_19119,N_19975);
nor UO_2145 (O_2145,N_18289,N_18930);
nor UO_2146 (O_2146,N_19477,N_18393);
and UO_2147 (O_2147,N_18207,N_19457);
or UO_2148 (O_2148,N_19090,N_19201);
and UO_2149 (O_2149,N_19305,N_18290);
or UO_2150 (O_2150,N_19694,N_18000);
nand UO_2151 (O_2151,N_19324,N_19454);
nor UO_2152 (O_2152,N_18945,N_19203);
nand UO_2153 (O_2153,N_18857,N_19779);
and UO_2154 (O_2154,N_18579,N_19872);
and UO_2155 (O_2155,N_18608,N_19441);
and UO_2156 (O_2156,N_18355,N_19075);
nand UO_2157 (O_2157,N_19536,N_19220);
or UO_2158 (O_2158,N_18533,N_18139);
nor UO_2159 (O_2159,N_18088,N_19512);
and UO_2160 (O_2160,N_19868,N_19983);
or UO_2161 (O_2161,N_19760,N_19372);
nand UO_2162 (O_2162,N_19517,N_19183);
nor UO_2163 (O_2163,N_19131,N_18655);
and UO_2164 (O_2164,N_19548,N_19462);
nor UO_2165 (O_2165,N_18850,N_19347);
nor UO_2166 (O_2166,N_19525,N_18366);
or UO_2167 (O_2167,N_19227,N_19094);
nand UO_2168 (O_2168,N_19196,N_18874);
nand UO_2169 (O_2169,N_19870,N_19395);
nor UO_2170 (O_2170,N_19004,N_18619);
or UO_2171 (O_2171,N_19639,N_19622);
or UO_2172 (O_2172,N_18855,N_18013);
or UO_2173 (O_2173,N_18805,N_19599);
nor UO_2174 (O_2174,N_18114,N_18255);
or UO_2175 (O_2175,N_18436,N_19522);
or UO_2176 (O_2176,N_19387,N_19025);
nand UO_2177 (O_2177,N_18187,N_19836);
or UO_2178 (O_2178,N_19168,N_18699);
and UO_2179 (O_2179,N_19510,N_18140);
and UO_2180 (O_2180,N_18065,N_19245);
nand UO_2181 (O_2181,N_18821,N_19518);
nand UO_2182 (O_2182,N_19137,N_18770);
or UO_2183 (O_2183,N_18792,N_19786);
and UO_2184 (O_2184,N_18285,N_18451);
nand UO_2185 (O_2185,N_19684,N_19201);
or UO_2186 (O_2186,N_18725,N_19782);
nand UO_2187 (O_2187,N_19961,N_18581);
and UO_2188 (O_2188,N_18915,N_19592);
nand UO_2189 (O_2189,N_19585,N_19365);
nand UO_2190 (O_2190,N_18808,N_18220);
or UO_2191 (O_2191,N_18878,N_18476);
and UO_2192 (O_2192,N_18886,N_18157);
nor UO_2193 (O_2193,N_19132,N_19088);
and UO_2194 (O_2194,N_19772,N_18715);
and UO_2195 (O_2195,N_18132,N_18376);
nand UO_2196 (O_2196,N_18012,N_19038);
and UO_2197 (O_2197,N_19891,N_18113);
nor UO_2198 (O_2198,N_18405,N_19549);
or UO_2199 (O_2199,N_18368,N_18105);
and UO_2200 (O_2200,N_18189,N_19598);
nor UO_2201 (O_2201,N_19853,N_18066);
nor UO_2202 (O_2202,N_18738,N_18534);
nand UO_2203 (O_2203,N_18791,N_19305);
and UO_2204 (O_2204,N_19449,N_18093);
nor UO_2205 (O_2205,N_19403,N_18019);
or UO_2206 (O_2206,N_19687,N_18519);
and UO_2207 (O_2207,N_19250,N_19895);
and UO_2208 (O_2208,N_19155,N_19857);
nand UO_2209 (O_2209,N_18715,N_19601);
or UO_2210 (O_2210,N_19256,N_19839);
or UO_2211 (O_2211,N_19648,N_18400);
or UO_2212 (O_2212,N_19689,N_18376);
or UO_2213 (O_2213,N_19832,N_19329);
nand UO_2214 (O_2214,N_18742,N_18633);
nor UO_2215 (O_2215,N_18350,N_19415);
or UO_2216 (O_2216,N_18844,N_18772);
nand UO_2217 (O_2217,N_19019,N_18964);
nor UO_2218 (O_2218,N_18700,N_19052);
or UO_2219 (O_2219,N_18337,N_18298);
and UO_2220 (O_2220,N_18502,N_19181);
nor UO_2221 (O_2221,N_19443,N_18115);
nand UO_2222 (O_2222,N_19984,N_19572);
xor UO_2223 (O_2223,N_19103,N_18297);
or UO_2224 (O_2224,N_19855,N_19552);
nor UO_2225 (O_2225,N_19626,N_18557);
or UO_2226 (O_2226,N_19982,N_19831);
or UO_2227 (O_2227,N_19528,N_19240);
nor UO_2228 (O_2228,N_18909,N_19715);
or UO_2229 (O_2229,N_19201,N_19239);
or UO_2230 (O_2230,N_19638,N_18974);
nor UO_2231 (O_2231,N_18106,N_18077);
or UO_2232 (O_2232,N_19113,N_18509);
nor UO_2233 (O_2233,N_19085,N_18286);
nand UO_2234 (O_2234,N_18110,N_19990);
or UO_2235 (O_2235,N_19707,N_18348);
nor UO_2236 (O_2236,N_18555,N_19829);
nand UO_2237 (O_2237,N_19544,N_19349);
and UO_2238 (O_2238,N_18781,N_18553);
nor UO_2239 (O_2239,N_19787,N_18515);
or UO_2240 (O_2240,N_18872,N_18890);
or UO_2241 (O_2241,N_19935,N_19009);
and UO_2242 (O_2242,N_18702,N_18952);
and UO_2243 (O_2243,N_19159,N_19921);
nor UO_2244 (O_2244,N_19669,N_19749);
and UO_2245 (O_2245,N_18585,N_18460);
nand UO_2246 (O_2246,N_18453,N_18006);
nand UO_2247 (O_2247,N_18758,N_18053);
nand UO_2248 (O_2248,N_19002,N_19870);
and UO_2249 (O_2249,N_18878,N_19324);
nor UO_2250 (O_2250,N_18436,N_19323);
nor UO_2251 (O_2251,N_18592,N_18320);
nand UO_2252 (O_2252,N_19472,N_19762);
nor UO_2253 (O_2253,N_19325,N_19611);
nor UO_2254 (O_2254,N_18511,N_18454);
or UO_2255 (O_2255,N_19327,N_19222);
or UO_2256 (O_2256,N_19300,N_19376);
and UO_2257 (O_2257,N_19099,N_19256);
and UO_2258 (O_2258,N_19521,N_18885);
nor UO_2259 (O_2259,N_18239,N_18298);
nand UO_2260 (O_2260,N_18293,N_18013);
nor UO_2261 (O_2261,N_18971,N_18004);
and UO_2262 (O_2262,N_19135,N_19948);
nand UO_2263 (O_2263,N_18068,N_18301);
or UO_2264 (O_2264,N_19054,N_18368);
nand UO_2265 (O_2265,N_18517,N_19370);
nor UO_2266 (O_2266,N_19229,N_18640);
and UO_2267 (O_2267,N_19957,N_18815);
or UO_2268 (O_2268,N_18924,N_19810);
nand UO_2269 (O_2269,N_19911,N_19575);
or UO_2270 (O_2270,N_18678,N_19776);
nor UO_2271 (O_2271,N_18167,N_19089);
and UO_2272 (O_2272,N_19511,N_18697);
nand UO_2273 (O_2273,N_18880,N_18892);
or UO_2274 (O_2274,N_19760,N_18357);
nor UO_2275 (O_2275,N_19725,N_19386);
nand UO_2276 (O_2276,N_19101,N_18271);
nor UO_2277 (O_2277,N_19448,N_19084);
or UO_2278 (O_2278,N_18674,N_18950);
nand UO_2279 (O_2279,N_18410,N_19433);
and UO_2280 (O_2280,N_19633,N_18242);
nor UO_2281 (O_2281,N_19600,N_19039);
or UO_2282 (O_2282,N_19093,N_18344);
nor UO_2283 (O_2283,N_19103,N_18923);
nand UO_2284 (O_2284,N_19959,N_19335);
nand UO_2285 (O_2285,N_19903,N_19204);
and UO_2286 (O_2286,N_18958,N_19383);
and UO_2287 (O_2287,N_18963,N_19859);
nor UO_2288 (O_2288,N_18953,N_19565);
and UO_2289 (O_2289,N_18611,N_18070);
and UO_2290 (O_2290,N_18534,N_18089);
and UO_2291 (O_2291,N_18181,N_18759);
or UO_2292 (O_2292,N_18602,N_18507);
nand UO_2293 (O_2293,N_19810,N_18661);
xnor UO_2294 (O_2294,N_18045,N_18803);
or UO_2295 (O_2295,N_18077,N_19102);
nor UO_2296 (O_2296,N_19744,N_19144);
and UO_2297 (O_2297,N_19612,N_18669);
and UO_2298 (O_2298,N_19563,N_19208);
or UO_2299 (O_2299,N_18211,N_18966);
nand UO_2300 (O_2300,N_18348,N_18325);
nor UO_2301 (O_2301,N_18621,N_18302);
and UO_2302 (O_2302,N_18297,N_18544);
nand UO_2303 (O_2303,N_18338,N_19477);
nand UO_2304 (O_2304,N_19517,N_19441);
or UO_2305 (O_2305,N_18011,N_18978);
or UO_2306 (O_2306,N_18520,N_18126);
nor UO_2307 (O_2307,N_19153,N_19087);
nand UO_2308 (O_2308,N_18482,N_18923);
nand UO_2309 (O_2309,N_18509,N_18405);
nand UO_2310 (O_2310,N_18962,N_18066);
or UO_2311 (O_2311,N_18294,N_18119);
or UO_2312 (O_2312,N_18540,N_19965);
xor UO_2313 (O_2313,N_18489,N_19596);
and UO_2314 (O_2314,N_18969,N_19199);
or UO_2315 (O_2315,N_18601,N_19751);
nand UO_2316 (O_2316,N_18819,N_18662);
nor UO_2317 (O_2317,N_18701,N_18783);
and UO_2318 (O_2318,N_19481,N_18240);
and UO_2319 (O_2319,N_18033,N_18508);
or UO_2320 (O_2320,N_18275,N_19540);
and UO_2321 (O_2321,N_19384,N_18627);
or UO_2322 (O_2322,N_19368,N_19122);
or UO_2323 (O_2323,N_18994,N_19861);
nor UO_2324 (O_2324,N_18659,N_19364);
nand UO_2325 (O_2325,N_19186,N_19986);
nor UO_2326 (O_2326,N_18766,N_19155);
or UO_2327 (O_2327,N_19661,N_18005);
nor UO_2328 (O_2328,N_19816,N_19946);
or UO_2329 (O_2329,N_18010,N_19717);
nand UO_2330 (O_2330,N_19810,N_19502);
and UO_2331 (O_2331,N_18900,N_19593);
nor UO_2332 (O_2332,N_19528,N_18075);
and UO_2333 (O_2333,N_18607,N_19442);
nand UO_2334 (O_2334,N_18101,N_19658);
and UO_2335 (O_2335,N_18034,N_19768);
nor UO_2336 (O_2336,N_18933,N_19577);
nor UO_2337 (O_2337,N_19956,N_18008);
or UO_2338 (O_2338,N_19356,N_18479);
nand UO_2339 (O_2339,N_18289,N_18550);
nand UO_2340 (O_2340,N_18595,N_19310);
or UO_2341 (O_2341,N_19788,N_18146);
nand UO_2342 (O_2342,N_18496,N_19701);
and UO_2343 (O_2343,N_19069,N_19952);
nand UO_2344 (O_2344,N_18772,N_19986);
nor UO_2345 (O_2345,N_18482,N_18500);
and UO_2346 (O_2346,N_19200,N_18999);
nand UO_2347 (O_2347,N_19197,N_19016);
nand UO_2348 (O_2348,N_19566,N_18283);
nor UO_2349 (O_2349,N_19058,N_18846);
nor UO_2350 (O_2350,N_18018,N_19315);
nor UO_2351 (O_2351,N_19960,N_19060);
or UO_2352 (O_2352,N_18358,N_19381);
nor UO_2353 (O_2353,N_19371,N_19460);
or UO_2354 (O_2354,N_18695,N_18020);
nor UO_2355 (O_2355,N_19353,N_19865);
or UO_2356 (O_2356,N_18079,N_18986);
and UO_2357 (O_2357,N_19650,N_19768);
nor UO_2358 (O_2358,N_19062,N_19120);
or UO_2359 (O_2359,N_19349,N_18723);
nor UO_2360 (O_2360,N_18954,N_18779);
nand UO_2361 (O_2361,N_18487,N_18849);
nand UO_2362 (O_2362,N_19274,N_19945);
nand UO_2363 (O_2363,N_18284,N_18781);
nor UO_2364 (O_2364,N_19236,N_19951);
and UO_2365 (O_2365,N_18694,N_19278);
and UO_2366 (O_2366,N_18586,N_19150);
nor UO_2367 (O_2367,N_19480,N_18812);
and UO_2368 (O_2368,N_19049,N_19437);
and UO_2369 (O_2369,N_19312,N_18867);
or UO_2370 (O_2370,N_19705,N_19906);
nand UO_2371 (O_2371,N_19509,N_18131);
and UO_2372 (O_2372,N_19620,N_19974);
nand UO_2373 (O_2373,N_19131,N_18365);
or UO_2374 (O_2374,N_19276,N_18857);
or UO_2375 (O_2375,N_19853,N_18185);
nand UO_2376 (O_2376,N_19373,N_19076);
nand UO_2377 (O_2377,N_19566,N_18524);
nand UO_2378 (O_2378,N_18103,N_18973);
nand UO_2379 (O_2379,N_18895,N_19685);
nand UO_2380 (O_2380,N_19146,N_19478);
or UO_2381 (O_2381,N_18636,N_18853);
nand UO_2382 (O_2382,N_19239,N_18935);
nor UO_2383 (O_2383,N_19515,N_19420);
and UO_2384 (O_2384,N_18017,N_18997);
or UO_2385 (O_2385,N_18119,N_19277);
xor UO_2386 (O_2386,N_18549,N_19351);
or UO_2387 (O_2387,N_19553,N_18309);
or UO_2388 (O_2388,N_18227,N_18043);
nor UO_2389 (O_2389,N_19239,N_19083);
and UO_2390 (O_2390,N_18654,N_18147);
or UO_2391 (O_2391,N_19119,N_18500);
and UO_2392 (O_2392,N_19551,N_18640);
nor UO_2393 (O_2393,N_19694,N_18152);
and UO_2394 (O_2394,N_18666,N_18585);
and UO_2395 (O_2395,N_18717,N_19069);
or UO_2396 (O_2396,N_18570,N_18815);
or UO_2397 (O_2397,N_18697,N_18765);
nand UO_2398 (O_2398,N_18135,N_19616);
nand UO_2399 (O_2399,N_18882,N_18353);
and UO_2400 (O_2400,N_19988,N_18867);
nor UO_2401 (O_2401,N_19380,N_19234);
nand UO_2402 (O_2402,N_19851,N_18150);
nand UO_2403 (O_2403,N_19309,N_18774);
or UO_2404 (O_2404,N_18271,N_18635);
nand UO_2405 (O_2405,N_18737,N_18264);
or UO_2406 (O_2406,N_18663,N_19757);
nor UO_2407 (O_2407,N_18562,N_18396);
or UO_2408 (O_2408,N_19369,N_18163);
or UO_2409 (O_2409,N_18010,N_19389);
and UO_2410 (O_2410,N_19242,N_19079);
nor UO_2411 (O_2411,N_18930,N_19130);
xor UO_2412 (O_2412,N_19505,N_19185);
or UO_2413 (O_2413,N_19586,N_18078);
nor UO_2414 (O_2414,N_18011,N_18973);
and UO_2415 (O_2415,N_19709,N_19786);
nor UO_2416 (O_2416,N_19067,N_18346);
nand UO_2417 (O_2417,N_18256,N_19570);
nand UO_2418 (O_2418,N_18150,N_18896);
or UO_2419 (O_2419,N_19539,N_18563);
nor UO_2420 (O_2420,N_18420,N_19951);
nand UO_2421 (O_2421,N_19562,N_18383);
or UO_2422 (O_2422,N_18992,N_19173);
or UO_2423 (O_2423,N_19412,N_19770);
nor UO_2424 (O_2424,N_19011,N_18018);
and UO_2425 (O_2425,N_19280,N_18957);
nand UO_2426 (O_2426,N_18923,N_19118);
or UO_2427 (O_2427,N_19075,N_18973);
and UO_2428 (O_2428,N_19740,N_18952);
nor UO_2429 (O_2429,N_19559,N_18655);
and UO_2430 (O_2430,N_19812,N_18054);
nor UO_2431 (O_2431,N_19263,N_19860);
nand UO_2432 (O_2432,N_18428,N_19770);
and UO_2433 (O_2433,N_18248,N_19696);
or UO_2434 (O_2434,N_19718,N_18714);
nand UO_2435 (O_2435,N_19899,N_19465);
nand UO_2436 (O_2436,N_19835,N_19633);
xnor UO_2437 (O_2437,N_18063,N_19088);
nand UO_2438 (O_2438,N_18777,N_18983);
nor UO_2439 (O_2439,N_18533,N_19656);
nor UO_2440 (O_2440,N_19128,N_19167);
and UO_2441 (O_2441,N_19719,N_18210);
or UO_2442 (O_2442,N_19731,N_19898);
or UO_2443 (O_2443,N_18229,N_19262);
or UO_2444 (O_2444,N_19277,N_18082);
and UO_2445 (O_2445,N_18470,N_19992);
or UO_2446 (O_2446,N_18661,N_19330);
or UO_2447 (O_2447,N_18714,N_18498);
nor UO_2448 (O_2448,N_19949,N_19505);
nor UO_2449 (O_2449,N_19707,N_19027);
and UO_2450 (O_2450,N_18867,N_19584);
nand UO_2451 (O_2451,N_18314,N_19890);
or UO_2452 (O_2452,N_18804,N_19331);
nor UO_2453 (O_2453,N_19988,N_19091);
or UO_2454 (O_2454,N_19112,N_19416);
and UO_2455 (O_2455,N_19334,N_18226);
and UO_2456 (O_2456,N_18140,N_19678);
nand UO_2457 (O_2457,N_19713,N_19466);
nor UO_2458 (O_2458,N_19574,N_18734);
and UO_2459 (O_2459,N_18186,N_18878);
nor UO_2460 (O_2460,N_19454,N_19143);
or UO_2461 (O_2461,N_18584,N_19108);
and UO_2462 (O_2462,N_18630,N_18095);
and UO_2463 (O_2463,N_18182,N_18407);
and UO_2464 (O_2464,N_18728,N_18008);
or UO_2465 (O_2465,N_19280,N_19046);
nand UO_2466 (O_2466,N_18818,N_19353);
nand UO_2467 (O_2467,N_19159,N_18691);
nand UO_2468 (O_2468,N_18180,N_19501);
xor UO_2469 (O_2469,N_18062,N_19887);
or UO_2470 (O_2470,N_18822,N_19001);
and UO_2471 (O_2471,N_19016,N_18917);
nor UO_2472 (O_2472,N_18001,N_18693);
nand UO_2473 (O_2473,N_19662,N_18783);
and UO_2474 (O_2474,N_18103,N_19982);
nand UO_2475 (O_2475,N_19548,N_18993);
or UO_2476 (O_2476,N_19474,N_18414);
nor UO_2477 (O_2477,N_18184,N_18797);
nand UO_2478 (O_2478,N_18386,N_19674);
and UO_2479 (O_2479,N_18290,N_19387);
and UO_2480 (O_2480,N_18167,N_18521);
nand UO_2481 (O_2481,N_19200,N_19187);
and UO_2482 (O_2482,N_19146,N_19090);
nor UO_2483 (O_2483,N_18981,N_18704);
and UO_2484 (O_2484,N_19279,N_19767);
and UO_2485 (O_2485,N_18607,N_19351);
nand UO_2486 (O_2486,N_18256,N_19812);
nand UO_2487 (O_2487,N_18165,N_18618);
or UO_2488 (O_2488,N_19284,N_18441);
nor UO_2489 (O_2489,N_19256,N_18055);
nand UO_2490 (O_2490,N_18746,N_18899);
and UO_2491 (O_2491,N_18824,N_18595);
and UO_2492 (O_2492,N_19375,N_19824);
or UO_2493 (O_2493,N_19349,N_19568);
or UO_2494 (O_2494,N_18689,N_18606);
nor UO_2495 (O_2495,N_19589,N_19552);
nor UO_2496 (O_2496,N_18416,N_19553);
nor UO_2497 (O_2497,N_18048,N_19184);
or UO_2498 (O_2498,N_18852,N_18505);
and UO_2499 (O_2499,N_19336,N_19976);
endmodule