module basic_2500_25000_3000_20_levels_10xor_3(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
or U0 (N_0,In_1803,In_467);
or U1 (N_1,In_275,In_752);
and U2 (N_2,In_2151,In_423);
xor U3 (N_3,In_1948,In_798);
nor U4 (N_4,In_806,In_702);
and U5 (N_5,In_136,In_1335);
nand U6 (N_6,In_776,In_2041);
xnor U7 (N_7,In_1665,In_677);
and U8 (N_8,In_1092,In_899);
nor U9 (N_9,In_2291,In_18);
or U10 (N_10,In_2468,In_430);
or U11 (N_11,In_2267,In_1025);
nor U12 (N_12,In_501,In_2422);
nor U13 (N_13,In_1498,In_2346);
nand U14 (N_14,In_838,In_2356);
xor U15 (N_15,In_1475,In_1462);
nor U16 (N_16,In_200,In_710);
xor U17 (N_17,In_134,In_810);
nor U18 (N_18,In_1779,In_586);
nand U19 (N_19,In_1552,In_2308);
nand U20 (N_20,In_732,In_2217);
nor U21 (N_21,In_2178,In_1773);
and U22 (N_22,In_1886,In_263);
nand U23 (N_23,In_1276,In_1627);
or U24 (N_24,In_853,In_1053);
nor U25 (N_25,In_1095,In_400);
nor U26 (N_26,In_2113,In_1590);
and U27 (N_27,In_966,In_1917);
nor U28 (N_28,In_1024,In_178);
and U29 (N_29,In_1302,In_2418);
or U30 (N_30,In_1546,In_1504);
xor U31 (N_31,In_609,In_2191);
nand U32 (N_32,In_1078,In_962);
and U33 (N_33,In_1018,In_886);
nor U34 (N_34,In_1481,In_1920);
or U35 (N_35,In_486,In_2248);
xnor U36 (N_36,In_1872,In_1512);
and U37 (N_37,In_1871,In_2097);
xor U38 (N_38,In_1457,In_2474);
or U39 (N_39,In_1807,In_2463);
xnor U40 (N_40,In_359,In_2261);
and U41 (N_41,In_2176,In_2358);
or U42 (N_42,In_22,In_1585);
xor U43 (N_43,In_866,In_2326);
or U44 (N_44,In_977,In_1305);
and U45 (N_45,In_1013,In_855);
nor U46 (N_46,In_1712,In_1353);
and U47 (N_47,In_790,In_2042);
or U48 (N_48,In_1572,In_1185);
nand U49 (N_49,In_690,In_2229);
and U50 (N_50,In_2200,In_2397);
xor U51 (N_51,In_1295,In_912);
or U52 (N_52,In_1605,In_2312);
nor U53 (N_53,In_982,In_1506);
and U54 (N_54,In_833,In_1369);
xor U55 (N_55,In_92,In_2034);
nor U56 (N_56,In_2426,In_640);
xor U57 (N_57,In_1818,In_662);
and U58 (N_58,In_28,In_203);
xor U59 (N_59,In_1775,In_1798);
nand U60 (N_60,In_2442,In_2439);
xnor U61 (N_61,In_137,In_2311);
nor U62 (N_62,In_462,In_1613);
nor U63 (N_63,In_1753,In_62);
nor U64 (N_64,In_1869,In_573);
nand U65 (N_65,In_1330,In_830);
xnor U66 (N_66,In_980,In_1242);
nand U67 (N_67,In_2466,In_2394);
xnor U68 (N_68,In_1780,In_1100);
and U69 (N_69,In_425,In_828);
nand U70 (N_70,In_708,In_2100);
xor U71 (N_71,In_1172,In_1105);
nand U72 (N_72,In_381,In_1350);
and U73 (N_73,In_2262,In_5);
nand U74 (N_74,In_71,In_441);
nand U75 (N_75,In_1183,In_252);
nor U76 (N_76,In_2232,In_1121);
nor U77 (N_77,In_685,In_1180);
nand U78 (N_78,In_1003,In_540);
and U79 (N_79,In_2082,In_1223);
or U80 (N_80,In_416,In_431);
nor U81 (N_81,In_1402,In_1472);
nor U82 (N_82,In_1165,In_1314);
or U83 (N_83,In_2373,In_459);
nor U84 (N_84,In_495,In_880);
and U85 (N_85,In_1301,In_588);
nor U86 (N_86,In_1876,In_754);
and U87 (N_87,In_1518,In_860);
or U88 (N_88,In_2121,In_572);
nand U89 (N_89,In_2378,In_1614);
and U90 (N_90,In_1226,In_676);
nand U91 (N_91,In_1254,In_13);
nand U92 (N_92,In_719,In_532);
nor U93 (N_93,In_2045,In_762);
and U94 (N_94,In_1080,In_1321);
and U95 (N_95,In_768,In_1111);
and U96 (N_96,In_668,In_1490);
nand U97 (N_97,In_2093,In_1919);
nand U98 (N_98,In_1714,In_1553);
nor U99 (N_99,In_353,In_1269);
xnor U100 (N_100,In_2103,In_1978);
or U101 (N_101,In_1908,In_1252);
xor U102 (N_102,In_665,In_240);
xor U103 (N_103,In_2107,In_1598);
xor U104 (N_104,In_642,In_1943);
nand U105 (N_105,In_2188,In_2456);
nor U106 (N_106,In_2416,In_43);
nor U107 (N_107,In_1249,In_2318);
xor U108 (N_108,In_1597,In_10);
nand U109 (N_109,In_1966,In_1157);
and U110 (N_110,In_1258,In_2381);
nor U111 (N_111,In_2197,In_1285);
and U112 (N_112,In_1713,In_1656);
xnor U113 (N_113,In_2390,In_308);
or U114 (N_114,In_273,In_904);
and U115 (N_115,In_700,In_96);
xor U116 (N_116,In_1804,In_1758);
or U117 (N_117,In_1926,In_923);
nand U118 (N_118,In_420,In_78);
or U119 (N_119,In_1397,In_1408);
and U120 (N_120,In_1678,In_835);
and U121 (N_121,In_785,In_1772);
nor U122 (N_122,In_248,In_819);
and U123 (N_123,In_2124,In_386);
or U124 (N_124,In_2167,In_2208);
nor U125 (N_125,In_298,In_1153);
nand U126 (N_126,In_120,In_505);
nor U127 (N_127,In_2013,In_352);
and U128 (N_128,In_1534,In_2379);
or U129 (N_129,In_219,In_2164);
nor U130 (N_130,In_1449,In_1097);
xor U131 (N_131,In_1759,In_2000);
and U132 (N_132,In_566,In_883);
or U133 (N_133,In_461,In_2295);
and U134 (N_134,In_1832,In_590);
nand U135 (N_135,In_1629,In_2289);
nand U136 (N_136,In_474,In_63);
xor U137 (N_137,In_543,In_2177);
and U138 (N_138,In_1407,In_1108);
and U139 (N_139,In_2410,In_872);
nand U140 (N_140,In_1448,In_3);
and U141 (N_141,In_1521,In_2206);
or U142 (N_142,In_2224,In_1533);
and U143 (N_143,In_2061,In_1272);
or U144 (N_144,In_321,In_816);
nor U145 (N_145,In_1833,In_1416);
nor U146 (N_146,In_1687,In_100);
xnor U147 (N_147,In_148,In_1983);
and U148 (N_148,In_1470,In_106);
xor U149 (N_149,In_341,In_2300);
xnor U150 (N_150,In_1455,In_832);
xnor U151 (N_151,In_322,In_1893);
xnor U152 (N_152,In_945,In_805);
xor U153 (N_153,In_2361,In_2196);
nor U154 (N_154,In_181,In_179);
nor U155 (N_155,In_1762,In_2084);
or U156 (N_156,In_1979,In_1537);
and U157 (N_157,In_2008,In_2328);
xor U158 (N_158,In_2486,In_1516);
xnor U159 (N_159,In_1756,In_207);
nor U160 (N_160,In_1539,In_1717);
and U161 (N_161,In_1428,In_1043);
xnor U162 (N_162,In_1998,In_215);
and U163 (N_163,In_2110,In_2115);
nand U164 (N_164,In_1234,In_1440);
and U165 (N_165,In_1468,In_1177);
nor U166 (N_166,In_670,In_2274);
or U167 (N_167,In_479,In_1137);
nor U168 (N_168,In_1733,In_1698);
nand U169 (N_169,In_1777,In_884);
nor U170 (N_170,In_715,In_163);
nand U171 (N_171,In_2341,In_1623);
or U172 (N_172,In_285,In_489);
and U173 (N_173,In_2004,In_1873);
nor U174 (N_174,In_382,In_1396);
and U175 (N_175,In_2117,In_651);
and U176 (N_176,In_1322,In_862);
nand U177 (N_177,In_463,In_879);
nand U178 (N_178,In_1076,In_1381);
and U179 (N_179,In_657,In_1438);
or U180 (N_180,In_39,In_1126);
or U181 (N_181,In_1661,In_885);
or U182 (N_182,In_1473,In_784);
and U183 (N_183,In_104,In_1827);
nor U184 (N_184,In_1579,In_2010);
and U185 (N_185,In_168,In_1471);
xor U186 (N_186,In_636,In_1805);
or U187 (N_187,In_2480,In_1030);
nor U188 (N_188,In_437,In_1587);
xnor U189 (N_189,In_786,In_2239);
nand U190 (N_190,In_242,In_1766);
nor U191 (N_191,In_1348,In_2259);
and U192 (N_192,In_758,In_477);
nand U193 (N_193,In_930,In_289);
nand U194 (N_194,In_2046,In_1128);
xor U195 (N_195,In_1958,In_31);
nand U196 (N_196,In_173,In_1515);
nand U197 (N_197,In_7,In_969);
or U198 (N_198,In_1461,In_2112);
nand U199 (N_199,In_1564,In_333);
xor U200 (N_200,In_2286,In_1328);
nor U201 (N_201,In_373,In_448);
nand U202 (N_202,In_1327,In_1159);
nand U203 (N_203,In_2080,In_396);
nand U204 (N_204,In_2174,In_473);
nand U205 (N_205,In_517,In_2050);
nor U206 (N_206,In_1543,In_926);
nor U207 (N_207,In_1808,In_189);
or U208 (N_208,In_541,In_1576);
nand U209 (N_209,In_648,In_531);
xor U210 (N_210,In_442,In_1158);
nor U211 (N_211,In_1316,In_1391);
nand U212 (N_212,In_1719,In_1768);
nor U213 (N_213,In_2019,In_983);
or U214 (N_214,In_1421,In_2420);
or U215 (N_215,In_2454,In_125);
and U216 (N_216,In_1433,In_1696);
and U217 (N_217,In_2132,In_1415);
or U218 (N_218,In_413,In_1835);
nand U219 (N_219,In_1615,In_344);
nand U220 (N_220,In_686,In_1778);
xor U221 (N_221,In_654,In_379);
and U222 (N_222,In_1846,In_2370);
nand U223 (N_223,In_1161,In_1822);
nand U224 (N_224,In_1444,In_1639);
and U225 (N_225,In_2471,In_1463);
xnor U226 (N_226,In_2056,In_155);
or U227 (N_227,In_2421,In_749);
nand U228 (N_228,In_2412,In_1437);
and U229 (N_229,In_2455,In_619);
and U230 (N_230,In_2225,In_2265);
or U231 (N_231,In_365,In_1082);
nor U232 (N_232,In_1439,In_2130);
nor U233 (N_233,In_206,In_380);
nand U234 (N_234,In_2448,In_1566);
and U235 (N_235,In_2281,In_2223);
or U236 (N_236,In_2302,In_2184);
or U237 (N_237,In_1371,In_1744);
nor U238 (N_238,In_124,In_274);
or U239 (N_239,In_1664,In_1582);
xor U240 (N_240,In_2487,In_1839);
nor U241 (N_241,In_658,In_21);
and U242 (N_242,In_457,In_1363);
or U243 (N_243,In_579,In_2205);
xnor U244 (N_244,In_388,In_484);
nor U245 (N_245,In_2494,In_2091);
nor U246 (N_246,In_653,In_2179);
nand U247 (N_247,In_1549,In_1797);
nor U248 (N_248,In_679,In_1251);
nor U249 (N_249,In_961,In_777);
and U250 (N_250,In_1862,In_1790);
or U251 (N_251,In_1284,In_1346);
xor U252 (N_252,In_89,In_1264);
and U253 (N_253,In_613,In_1253);
nand U254 (N_254,In_595,In_478);
xor U255 (N_255,In_2282,In_779);
xor U256 (N_256,In_1152,In_970);
or U257 (N_257,In_1352,In_1476);
or U258 (N_258,In_237,In_770);
nand U259 (N_259,In_1238,In_384);
and U260 (N_260,In_935,In_1200);
nand U261 (N_261,In_2193,In_615);
xor U262 (N_262,In_1483,In_2351);
and U263 (N_263,In_1046,In_1829);
nor U264 (N_264,In_2228,In_372);
xnor U265 (N_265,In_1334,In_364);
nor U266 (N_266,In_1509,In_597);
xnor U267 (N_267,In_127,In_2327);
and U268 (N_268,In_236,In_271);
nor U269 (N_269,In_792,In_184);
and U270 (N_270,In_946,In_351);
or U271 (N_271,In_1273,In_1729);
nor U272 (N_272,In_2280,In_1649);
nor U273 (N_273,In_497,In_1164);
and U274 (N_274,In_1116,In_852);
and U275 (N_275,In_1229,In_681);
and U276 (N_276,In_1634,In_1300);
and U277 (N_277,In_1250,In_447);
or U278 (N_278,In_2180,In_226);
and U279 (N_279,In_1500,In_2175);
and U280 (N_280,In_1842,In_1187);
nand U281 (N_281,In_1062,In_79);
xor U282 (N_282,In_2479,In_1606);
nand U283 (N_283,In_604,In_850);
xor U284 (N_284,In_2145,In_2297);
nor U285 (N_285,In_196,In_2192);
nor U286 (N_286,In_393,In_1542);
and U287 (N_287,In_1022,In_2018);
and U288 (N_288,In_2362,In_1995);
and U289 (N_289,In_2357,In_1697);
nand U290 (N_290,In_492,In_2033);
nand U291 (N_291,In_211,In_1558);
xnor U292 (N_292,In_458,In_210);
nor U293 (N_293,In_1163,In_1955);
xnor U294 (N_294,In_1771,In_756);
xor U295 (N_295,In_2380,In_1795);
and U296 (N_296,In_829,In_378);
and U297 (N_297,In_706,In_655);
nor U298 (N_298,In_453,In_2344);
nand U299 (N_299,In_2227,In_759);
or U300 (N_300,In_450,In_1118);
and U301 (N_301,In_1265,In_2059);
and U302 (N_302,In_1929,In_1290);
nand U303 (N_303,In_2491,In_1205);
or U304 (N_304,In_395,In_2347);
and U305 (N_305,In_842,In_1294);
nand U306 (N_306,In_1530,In_429);
nand U307 (N_307,In_800,In_464);
and U308 (N_308,In_160,In_327);
and U309 (N_309,In_1282,In_229);
or U310 (N_310,In_357,In_269);
or U311 (N_311,In_227,In_503);
xor U312 (N_312,In_797,In_897);
and U313 (N_313,In_1227,In_277);
xnor U314 (N_314,In_311,In_1347);
xnor U315 (N_315,In_722,In_72);
nand U316 (N_316,In_180,In_2382);
nor U317 (N_317,In_2398,In_731);
nor U318 (N_318,In_1067,In_527);
or U319 (N_319,In_48,In_2436);
and U320 (N_320,In_1341,In_304);
xor U321 (N_321,In_817,In_340);
nand U322 (N_322,In_799,In_950);
and U323 (N_323,In_139,In_1336);
nand U324 (N_324,In_1089,In_1898);
xnor U325 (N_325,In_2360,In_2148);
xnor U326 (N_326,In_214,In_331);
or U327 (N_327,In_2446,In_1378);
and U328 (N_328,In_2071,In_2186);
nor U329 (N_329,In_1856,In_1655);
nand U330 (N_330,In_2430,In_2141);
and U331 (N_331,In_262,In_1936);
and U332 (N_332,In_140,In_1141);
xor U333 (N_333,In_1370,In_235);
and U334 (N_334,In_1589,In_846);
or U335 (N_335,In_185,In_88);
nand U336 (N_336,In_2190,In_601);
xnor U337 (N_337,In_2079,In_2065);
or U338 (N_338,In_1642,In_2383);
xnor U339 (N_339,In_1073,In_1070);
xnor U340 (N_340,In_222,In_1213);
and U341 (N_341,In_1429,In_2472);
xor U342 (N_342,In_158,In_174);
nand U343 (N_343,In_2377,In_1474);
and U344 (N_344,In_2335,In_2022);
or U345 (N_345,In_1691,In_2083);
or U346 (N_346,In_631,In_1796);
or U347 (N_347,In_2162,In_2094);
or U348 (N_348,In_1975,In_494);
nand U349 (N_349,In_596,In_1890);
nor U350 (N_350,In_581,In_1666);
nand U351 (N_351,In_1855,In_2202);
and U352 (N_352,In_264,In_942);
xor U353 (N_353,In_2476,In_1909);
or U354 (N_354,In_1540,In_647);
nor U355 (N_355,In_2152,In_1166);
nor U356 (N_356,In_253,In_628);
and U357 (N_357,In_2102,In_2078);
xnor U358 (N_358,In_1863,In_1843);
and U359 (N_359,In_1460,In_1431);
and U360 (N_360,In_1736,In_827);
and U361 (N_361,In_1123,In_243);
nand U362 (N_362,In_803,In_175);
or U363 (N_363,In_1088,In_32);
and U364 (N_364,In_954,In_1545);
nand U365 (N_365,In_1033,In_730);
nor U366 (N_366,In_2234,In_1709);
or U367 (N_367,In_1907,In_2271);
or U368 (N_368,In_663,In_1311);
xnor U369 (N_369,In_576,In_1374);
nor U370 (N_370,In_1279,In_2369);
xnor U371 (N_371,In_326,In_1517);
or U372 (N_372,In_1257,In_2153);
xnor U373 (N_373,In_916,In_1299);
nor U374 (N_374,In_192,In_2220);
xnor U375 (N_375,In_671,In_1075);
nand U376 (N_376,In_394,In_144);
or U377 (N_377,In_1426,In_1551);
and U378 (N_378,In_1066,In_746);
nand U379 (N_379,In_482,In_117);
nand U380 (N_380,In_1609,In_528);
xnor U381 (N_381,In_301,In_84);
nand U382 (N_382,In_2150,In_1817);
nor U383 (N_383,In_498,In_2163);
xnor U384 (N_384,In_542,In_2047);
xnor U385 (N_385,In_1198,In_2105);
nand U386 (N_386,In_1529,In_398);
xnor U387 (N_387,In_1648,In_1349);
nor U388 (N_388,In_1487,In_2343);
nor U389 (N_389,In_65,In_1441);
nor U390 (N_390,In_2137,In_2146);
and U391 (N_391,In_2134,In_500);
nor U392 (N_392,In_2417,In_1464);
xor U393 (N_393,In_469,In_1212);
or U394 (N_394,In_1016,In_212);
nor U395 (N_395,In_2037,In_1939);
xor U396 (N_396,In_2183,In_774);
nand U397 (N_397,In_1323,In_2189);
or U398 (N_398,In_1868,In_919);
nor U399 (N_399,In_102,In_1644);
nand U400 (N_400,In_697,In_772);
nor U401 (N_401,In_1853,In_1256);
nand U402 (N_402,In_45,In_83);
or U403 (N_403,In_1959,In_1538);
nor U404 (N_404,In_2269,In_1662);
xor U405 (N_405,In_844,In_1565);
or U406 (N_406,In_2428,In_2388);
xnor U407 (N_407,In_512,In_1181);
xor U408 (N_408,In_551,In_2469);
and U409 (N_409,In_513,In_570);
xnor U410 (N_410,In_626,In_1726);
nand U411 (N_411,In_108,In_110);
nand U412 (N_412,In_1784,In_1864);
nor U413 (N_413,In_728,In_550);
xor U414 (N_414,In_981,In_796);
xnor U415 (N_415,In_455,In_112);
and U416 (N_416,In_856,In_1632);
nand U417 (N_417,In_1608,In_419);
and U418 (N_418,In_1313,In_217);
xnor U419 (N_419,In_1482,In_1637);
or U420 (N_420,In_948,In_228);
xnor U421 (N_421,In_1994,In_169);
xnor U422 (N_422,In_1554,In_667);
or U423 (N_423,In_361,In_2285);
and U424 (N_424,In_839,In_354);
nor U425 (N_425,In_1547,In_849);
and U426 (N_426,In_1233,In_592);
nand U427 (N_427,In_1973,In_154);
nor U428 (N_428,In_1297,In_2215);
and U429 (N_429,In_51,In_1786);
xnor U430 (N_430,In_1,In_422);
nor U431 (N_431,In_1283,In_1742);
nor U432 (N_432,In_1556,In_307);
xnor U433 (N_433,In_1686,In_1189);
or U434 (N_434,In_387,In_1934);
and U435 (N_435,In_2063,In_1711);
and U436 (N_436,In_1178,In_41);
xnor U437 (N_437,In_493,In_2185);
nand U438 (N_438,In_306,In_520);
or U439 (N_439,In_114,In_1899);
nand U440 (N_440,In_141,In_2154);
xnor U441 (N_441,In_721,In_1492);
or U442 (N_442,In_245,In_107);
nand U443 (N_443,In_2096,In_630);
or U444 (N_444,In_583,In_2389);
or U445 (N_445,In_1986,In_1010);
xor U446 (N_446,In_291,In_142);
xnor U447 (N_447,In_1902,In_2275);
xor U448 (N_448,In_1319,In_2201);
nand U449 (N_449,In_2074,In_2012);
nor U450 (N_450,In_2122,In_2114);
nor U451 (N_451,In_1049,In_766);
nor U452 (N_452,In_2324,In_1851);
nor U453 (N_453,In_119,In_221);
nor U454 (N_454,In_2230,In_2273);
xor U455 (N_455,In_1847,In_794);
xnor U456 (N_456,In_1124,In_1593);
nor U457 (N_457,In_958,In_1122);
and U458 (N_458,In_2098,In_76);
or U459 (N_459,In_995,In_1424);
nand U460 (N_460,In_131,In_392);
nor U461 (N_461,In_11,In_1601);
nor U462 (N_462,In_149,In_2195);
or U463 (N_463,In_1974,In_2235);
and U464 (N_464,In_733,In_1981);
and U465 (N_465,In_165,In_620);
xor U466 (N_466,In_1942,In_2073);
nor U467 (N_467,In_255,In_763);
or U468 (N_468,In_405,In_1896);
nor U469 (N_469,In_414,In_1800);
or U470 (N_470,In_2415,In_1887);
xnor U471 (N_471,In_2299,In_932);
or U472 (N_472,In_1217,In_661);
and U473 (N_473,In_523,In_404);
nand U474 (N_474,In_1247,In_1643);
xor U475 (N_475,In_1505,In_1479);
or U476 (N_476,In_1384,In_150);
xnor U477 (N_477,In_924,In_2258);
nand U478 (N_478,In_669,In_718);
nor U479 (N_479,In_1837,In_1625);
nor U480 (N_480,In_1340,In_281);
nand U481 (N_481,In_428,In_2256);
nand U482 (N_482,In_1581,In_741);
nand U483 (N_483,In_2473,In_220);
or U484 (N_484,In_1186,In_250);
and U485 (N_485,In_767,In_133);
nand U486 (N_486,In_553,In_2315);
and U487 (N_487,In_2488,In_2109);
nand U488 (N_488,In_2447,In_747);
nor U489 (N_489,In_764,In_2268);
or U490 (N_490,In_2287,In_1932);
nand U491 (N_491,In_1324,In_1970);
nand U492 (N_492,In_1764,In_113);
nor U493 (N_493,In_1931,In_1781);
and U494 (N_494,In_1560,In_2407);
xor U495 (N_495,In_845,In_1857);
or U496 (N_496,In_487,In_534);
xor U497 (N_497,In_612,In_1600);
and U498 (N_498,In_314,In_2449);
nand U499 (N_499,In_614,In_138);
nand U500 (N_500,In_1568,In_739);
nand U501 (N_501,In_2088,In_1592);
nor U502 (N_502,In_978,In_742);
xnor U503 (N_503,In_1865,In_868);
and U504 (N_504,In_2348,In_1513);
or U505 (N_505,In_2453,In_59);
xor U506 (N_506,In_703,In_913);
or U507 (N_507,In_1090,In_562);
xnor U508 (N_508,In_1069,In_1029);
and U509 (N_509,In_2116,In_2293);
xnor U510 (N_510,In_2264,In_1622);
nand U511 (N_511,In_1820,In_525);
nor U512 (N_512,In_1894,In_2160);
and U513 (N_513,In_1197,In_664);
xor U514 (N_514,In_2090,In_1596);
xor U515 (N_515,In_557,In_2495);
nor U516 (N_516,In_1425,In_1927);
nor U517 (N_517,In_826,In_802);
xnor U518 (N_518,In_336,In_1360);
nor U519 (N_519,In_2246,In_1459);
or U520 (N_520,In_2032,In_241);
or U521 (N_521,In_1039,In_1735);
nand U522 (N_522,In_2353,In_1617);
and U523 (N_523,In_1394,In_524);
nand U524 (N_524,In_2213,In_645);
or U525 (N_525,In_432,In_2016);
nand U526 (N_526,In_1211,In_1278);
and U527 (N_527,In_688,In_2372);
xnor U528 (N_528,In_1985,In_2218);
and U529 (N_529,In_616,In_2155);
xor U530 (N_530,In_564,In_675);
nand U531 (N_531,In_1501,In_1127);
xor U532 (N_532,In_476,In_24);
or U533 (N_533,In_1055,In_1971);
xor U534 (N_534,In_2067,In_1967);
nor U535 (N_535,In_1451,In_1281);
or U536 (N_536,In_452,In_1244);
xnor U537 (N_537,In_69,In_518);
or U538 (N_538,In_310,In_1716);
or U539 (N_539,In_1255,In_1338);
nand U540 (N_540,In_906,In_1002);
nor U541 (N_541,In_2493,In_66);
or U542 (N_542,In_905,In_2334);
or U543 (N_543,In_2391,In_258);
nor U544 (N_544,In_1236,In_1867);
or U545 (N_545,In_230,In_1823);
xnor U546 (N_546,In_75,In_1738);
and U547 (N_547,In_921,In_2029);
xor U548 (N_548,In_375,In_864);
or U549 (N_549,In_1103,In_2060);
xor U550 (N_550,In_2393,In_2255);
nor U551 (N_551,In_644,In_1412);
nor U552 (N_552,In_451,In_1237);
nor U553 (N_553,In_2009,In_1889);
nand U554 (N_554,In_1968,In_1280);
nor U555 (N_555,In_1184,In_2419);
nor U556 (N_556,In_329,In_330);
nand U557 (N_557,In_2433,In_2329);
nor U558 (N_558,In_1271,In_1571);
or U559 (N_559,In_376,In_521);
and U560 (N_560,In_1667,In_456);
nand U561 (N_561,In_496,In_1814);
xnor U562 (N_562,In_617,In_2349);
or U563 (N_563,In_684,In_743);
or U564 (N_564,In_788,In_313);
nand U565 (N_565,In_1012,In_1484);
nor U566 (N_566,In_834,In_2279);
and U567 (N_567,In_607,In_2290);
or U568 (N_568,In_287,In_40);
or U569 (N_569,In_471,In_2006);
nor U570 (N_570,In_406,In_1447);
nor U571 (N_571,In_1594,In_997);
nand U572 (N_572,In_268,In_317);
nand U573 (N_573,In_1417,In_1261);
nor U574 (N_574,In_1584,In_976);
and U575 (N_575,In_2440,In_943);
and U576 (N_576,In_190,In_836);
nor U577 (N_577,In_186,In_787);
and U578 (N_578,In_224,In_1139);
and U579 (N_579,In_1466,In_922);
nand U580 (N_580,In_2338,In_1631);
nand U581 (N_581,In_1120,In_1604);
xor U582 (N_582,In_941,In_2496);
nand U583 (N_583,In_937,In_1653);
and U584 (N_584,In_302,In_837);
nor U585 (N_585,In_705,In_594);
nand U586 (N_586,In_1423,In_1525);
nor U587 (N_587,In_591,In_1057);
or U588 (N_588,In_284,In_480);
nor U589 (N_589,In_2169,In_2076);
xnor U590 (N_590,In_418,In_811);
xnor U591 (N_591,In_901,In_247);
and U592 (N_592,In_1783,In_1945);
nor U593 (N_593,In_920,In_1355);
xor U594 (N_594,In_126,In_465);
xnor U595 (N_595,In_1386,In_223);
nand U596 (N_596,In_1050,In_621);
or U597 (N_597,In_1991,In_1883);
nand U598 (N_598,In_2366,In_2108);
nand U599 (N_599,In_1670,In_90);
nor U600 (N_600,In_890,In_239);
nand U601 (N_601,In_362,In_2464);
and U602 (N_602,In_346,In_1114);
or U603 (N_603,In_2461,In_1519);
nand U604 (N_604,In_1452,In_1502);
nor U605 (N_605,In_345,In_2431);
and U606 (N_606,In_544,In_1950);
xnor U607 (N_607,In_1432,In_2219);
nor U608 (N_608,In_748,In_1514);
nor U609 (N_609,In_1569,In_1951);
xnor U610 (N_610,In_533,In_729);
and U611 (N_611,In_587,In_1640);
nor U612 (N_612,In_618,In_130);
nand U613 (N_613,In_2371,In_91);
nand U614 (N_614,In_491,In_1776);
or U615 (N_615,In_2023,In_2209);
xnor U616 (N_616,In_1914,In_1398);
nor U617 (N_617,In_1916,In_652);
or U618 (N_618,In_1725,In_1510);
xnor U619 (N_619,In_911,In_1218);
and U620 (N_620,In_974,In_1913);
and U621 (N_621,In_964,In_182);
nand U622 (N_622,In_1112,In_2126);
xnor U623 (N_623,In_348,In_1792);
and U624 (N_624,In_1445,In_2399);
or U625 (N_625,In_2161,In_1176);
and U626 (N_626,In_1027,In_2020);
nand U627 (N_627,In_1750,In_2011);
nor U628 (N_628,In_128,In_488);
and U629 (N_629,In_1647,In_988);
or U630 (N_630,In_334,In_1739);
or U631 (N_631,In_558,In_1577);
nor U632 (N_632,In_1559,In_2323);
and U633 (N_633,In_1191,In_1052);
nor U634 (N_634,In_1787,In_1458);
and U635 (N_635,In_1684,In_183);
or U636 (N_636,In_143,In_843);
nand U637 (N_637,In_2238,In_1411);
nor U638 (N_638,In_1115,In_1390);
nand U639 (N_639,In_674,In_2171);
and U640 (N_640,In_1083,In_1129);
xor U641 (N_641,In_2147,In_103);
nand U642 (N_642,In_260,In_938);
or U643 (N_643,In_1150,In_1071);
nor U644 (N_644,In_1520,In_2104);
xnor U645 (N_645,In_1404,In_2272);
and U646 (N_646,In_2040,In_1826);
nand U647 (N_647,In_2408,In_1040);
nor U648 (N_648,In_472,In_1063);
and U649 (N_649,In_893,In_944);
nor U650 (N_650,In_2119,In_782);
or U651 (N_651,In_2445,In_1486);
xor U652 (N_652,In_1036,In_1102);
nand U653 (N_653,In_1304,In_2424);
and U654 (N_654,In_246,In_265);
nand U655 (N_655,In_870,In_1996);
xor U656 (N_656,In_1707,In_1673);
and U657 (N_657,In_1414,In_643);
nor U658 (N_658,In_1507,In_682);
nor U659 (N_659,In_809,In_2204);
or U660 (N_660,In_56,In_1267);
and U661 (N_661,In_1146,In_1875);
or U662 (N_662,In_1881,In_2136);
or U663 (N_663,In_385,In_771);
nand U664 (N_664,In_257,In_1791);
nand U665 (N_665,In_349,In_37);
and U666 (N_666,In_1044,In_793);
and U667 (N_667,In_1221,In_409);
xnor U668 (N_668,In_1992,In_38);
or U669 (N_669,In_6,In_1375);
or U670 (N_670,In_1203,In_2478);
xor U671 (N_671,In_1320,In_1834);
xor U672 (N_672,In_1045,In_468);
or U673 (N_673,In_443,In_2278);
and U674 (N_674,In_1326,In_251);
or U675 (N_675,In_2242,In_2296);
or U676 (N_676,In_1042,In_2435);
xor U677 (N_677,In_256,In_350);
nand U678 (N_678,In_44,In_1912);
nand U679 (N_679,In_1193,In_1870);
nand U680 (N_680,In_2156,In_773);
nand U681 (N_681,In_984,In_1658);
xnor U682 (N_682,In_1005,In_898);
and U683 (N_683,In_769,In_1028);
xor U684 (N_684,In_1020,In_1997);
xnor U685 (N_685,In_299,In_1984);
and U686 (N_686,In_582,In_1443);
or U687 (N_687,In_857,In_1954);
nor U688 (N_688,In_1065,In_1156);
xor U689 (N_689,In_1952,In_1925);
xor U690 (N_690,In_33,In_555);
and U691 (N_691,In_167,In_1387);
and U692 (N_692,In_2365,In_1357);
nand U693 (N_693,In_2005,In_358);
or U694 (N_694,In_483,In_1021);
nand U695 (N_695,In_656,In_1037);
xor U696 (N_696,In_187,In_266);
and U697 (N_697,In_1289,In_64);
nor U698 (N_698,In_1785,In_1924);
nand U699 (N_699,In_2173,In_1263);
xnor U700 (N_700,In_1173,In_1892);
nor U701 (N_701,In_672,In_2207);
nor U702 (N_702,In_1058,In_2036);
xnor U703 (N_703,In_1527,In_2035);
or U704 (N_704,In_1491,In_1006);
nor U705 (N_705,In_1532,In_454);
or U706 (N_706,In_891,In_1392);
nor U707 (N_707,In_2483,In_1214);
xnor U708 (N_708,In_1009,In_1293);
xor U709 (N_709,In_2484,In_356);
and U710 (N_710,In_2367,In_638);
or U711 (N_711,In_1143,In_634);
nand U712 (N_712,In_991,In_1017);
nor U713 (N_713,In_343,In_1859);
nor U714 (N_714,In_1160,In_996);
nor U715 (N_715,In_2120,In_2298);
nor U716 (N_716,In_927,In_2337);
nand U717 (N_717,In_1841,In_2460);
nor U718 (N_718,In_1171,In_545);
nor U719 (N_719,In_1325,In_261);
or U720 (N_720,In_1982,In_2497);
xnor U721 (N_721,In_1388,In_2194);
or U722 (N_722,In_694,In_8);
and U723 (N_723,In_509,In_377);
nand U724 (N_724,In_2423,In_2376);
and U725 (N_725,In_410,In_1094);
xor U726 (N_726,In_2432,In_650);
or U727 (N_727,In_1641,In_2352);
nand U728 (N_728,In_1413,In_701);
nand U729 (N_729,In_693,In_1201);
or U730 (N_730,In_814,In_1961);
and U731 (N_731,In_2165,In_1155);
xor U732 (N_732,In_2404,In_1232);
xor U733 (N_733,In_1848,In_1145);
xor U734 (N_734,In_205,In_234);
nor U735 (N_735,In_73,In_578);
nand U736 (N_736,In_2314,In_914);
xor U737 (N_737,In_1562,In_859);
or U738 (N_738,In_1701,In_1910);
xnor U739 (N_739,In_1162,In_1147);
or U740 (N_740,In_1573,In_153);
nand U741 (N_741,In_54,In_1495);
or U742 (N_742,In_1243,In_1099);
xnor U743 (N_743,In_1291,In_2026);
nand U744 (N_744,In_2007,In_67);
xor U745 (N_745,In_61,In_1224);
or U746 (N_746,In_1550,In_511);
or U747 (N_747,In_280,In_14);
nor U748 (N_748,In_1809,In_1700);
nand U749 (N_749,In_698,In_1493);
or U750 (N_750,In_439,In_2459);
nor U751 (N_751,In_267,In_426);
and U752 (N_752,In_1077,In_1765);
and U753 (N_753,In_1536,In_947);
nor U754 (N_754,In_1989,In_2221);
nand U755 (N_755,In_339,In_26);
and U756 (N_756,In_368,In_1574);
and U757 (N_757,In_87,In_1419);
nand U758 (N_758,In_1399,In_2305);
or U759 (N_759,In_1947,In_466);
nand U760 (N_760,In_724,In_1816);
or U761 (N_761,In_1689,In_1051);
nor U762 (N_762,In_1944,In_933);
xnor U763 (N_763,In_1953,In_1008);
nand U764 (N_764,In_318,In_1671);
and U765 (N_765,In_1059,In_360);
and U766 (N_766,In_2288,In_1651);
nand U767 (N_767,In_825,In_1119);
or U768 (N_768,In_1248,In_1900);
nand U769 (N_769,In_918,In_342);
nand U770 (N_770,In_691,In_1567);
nor U771 (N_771,In_2182,In_1204);
or U772 (N_772,In_1561,In_1794);
and U773 (N_773,In_696,In_225);
nor U774 (N_774,In_213,In_973);
and U775 (N_775,In_975,In_1903);
nor U776 (N_776,In_1400,In_1383);
nor U777 (N_777,In_369,In_775);
or U778 (N_778,In_402,In_2003);
and U779 (N_779,In_506,In_1720);
and U780 (N_780,In_1136,In_27);
xnor U781 (N_781,In_986,In_2270);
or U782 (N_782,In_1557,In_1362);
xnor U783 (N_783,In_2216,In_568);
or U784 (N_784,In_2072,In_1654);
nand U785 (N_785,In_389,In_780);
nand U786 (N_786,In_407,In_2025);
xor U787 (N_787,In_2322,In_1774);
nor U788 (N_788,In_1813,In_1544);
and U789 (N_789,In_109,In_1410);
nand U790 (N_790,In_1728,In_965);
nand U791 (N_791,In_446,In_370);
nor U792 (N_792,In_1946,In_565);
and U793 (N_793,In_1563,In_2342);
or U794 (N_794,In_1342,In_1752);
and U795 (N_795,In_1497,In_535);
nor U796 (N_796,In_1508,In_159);
nor U797 (N_797,In_2240,In_738);
and U798 (N_798,In_2490,In_1732);
xor U799 (N_799,In_1138,In_1599);
xor U800 (N_800,In_560,In_1084);
nor U801 (N_801,In_1332,In_2330);
and U802 (N_802,In_1578,In_1748);
nor U803 (N_803,In_2441,In_49);
and U804 (N_804,In_1339,In_1167);
nand U805 (N_805,In_1935,In_1937);
xnor U806 (N_806,In_323,In_680);
nor U807 (N_807,In_1406,In_2332);
and U808 (N_808,In_1526,In_519);
xor U809 (N_809,In_1047,In_1206);
and U810 (N_810,In_1072,In_254);
and U811 (N_811,In_1895,In_781);
nand U812 (N_812,In_1179,In_2363);
and U813 (N_813,In_1555,In_2048);
nand U814 (N_814,In_1618,In_1802);
xnor U815 (N_815,In_1048,In_1877);
and U816 (N_816,In_55,In_2139);
or U817 (N_817,In_2077,In_1845);
xor U818 (N_818,In_929,In_2170);
and U819 (N_819,In_1824,In_1131);
nor U820 (N_820,In_789,In_1174);
nand U821 (N_821,In_1677,In_97);
or U822 (N_822,In_2301,In_1923);
nor U823 (N_823,In_1395,In_1710);
nand U824 (N_824,In_320,In_1011);
or U825 (N_825,In_2499,In_2254);
or U826 (N_826,In_659,In_713);
nor U827 (N_827,In_1705,In_569);
xor U828 (N_828,In_637,In_2187);
and U829 (N_829,In_2368,In_2386);
nor U830 (N_830,In_421,In_999);
nand U831 (N_831,In_931,In_2172);
nand U832 (N_832,In_2294,In_968);
xor U833 (N_833,In_895,In_526);
nand U834 (N_834,In_559,In_122);
xnor U835 (N_835,In_2325,In_2292);
nand U836 (N_836,In_813,In_1969);
or U837 (N_837,In_2244,In_2212);
or U838 (N_838,In_1286,In_2354);
nand U839 (N_839,In_1635,In_305);
nand U840 (N_840,In_2414,In_972);
nor U841 (N_841,In_408,In_2157);
xor U842 (N_842,In_1246,In_1688);
nor U843 (N_843,In_1056,In_1734);
and U844 (N_844,In_1690,In_2333);
and U845 (N_845,In_1104,In_1382);
nand U846 (N_846,In_956,In_1318);
xnor U847 (N_847,In_1054,In_1963);
nand U848 (N_848,In_1453,In_2069);
or U849 (N_849,In_145,In_332);
or U850 (N_850,In_699,In_957);
nor U851 (N_851,In_1266,In_818);
and U852 (N_852,In_599,In_1422);
nand U853 (N_853,In_2064,In_1591);
nor U854 (N_854,In_1093,In_2401);
nand U855 (N_855,In_2236,In_622);
or U856 (N_856,In_1208,In_1081);
nor U857 (N_857,In_801,In_1828);
nor U858 (N_858,In_714,In_201);
and U859 (N_859,In_993,In_725);
nand U860 (N_860,In_1192,In_176);
xnor U861 (N_861,In_294,In_847);
xnor U862 (N_862,In_608,In_2092);
and U863 (N_863,In_1169,In_2053);
nand U864 (N_864,In_2345,In_172);
and U865 (N_865,In_171,In_15);
xor U866 (N_866,In_2477,In_2166);
nand U867 (N_867,In_1541,In_1675);
xor U868 (N_868,In_1356,In_1109);
nor U869 (N_869,In_765,In_309);
and U870 (N_870,In_2111,In_757);
or U871 (N_871,In_1801,In_2241);
nand U872 (N_872,In_295,In_199);
xor U873 (N_873,In_191,In_1418);
nand U874 (N_874,In_1888,In_1079);
nand U875 (N_875,In_12,In_709);
or U876 (N_876,In_2385,In_737);
and U877 (N_877,In_2142,In_29);
nor U878 (N_878,In_1523,In_403);
or U879 (N_879,In_98,In_16);
nor U880 (N_880,In_1879,In_2304);
and U881 (N_881,In_1064,In_1345);
xor U882 (N_882,In_1199,In_1906);
nand U883 (N_883,In_2211,In_1366);
or U884 (N_884,In_1806,In_23);
or U885 (N_885,In_1393,In_2359);
xnor U886 (N_886,In_712,In_0);
xnor U887 (N_887,In_2277,In_1674);
nor U888 (N_888,In_915,In_1724);
and U889 (N_889,In_1358,In_900);
nand U890 (N_890,In_2049,In_1019);
nor U891 (N_891,In_2475,In_1245);
nor U892 (N_892,In_1595,In_1531);
and U893 (N_893,In_760,In_723);
nor U894 (N_894,In_716,In_894);
nor U895 (N_895,In_908,In_873);
nor U896 (N_896,In_585,In_374);
and U897 (N_897,In_2149,In_1434);
xnor U898 (N_898,In_1993,In_1175);
nand U899 (N_899,In_1789,In_635);
or U900 (N_900,In_2252,In_2199);
nor U901 (N_901,In_435,In_936);
xor U902 (N_902,In_1494,In_539);
and U903 (N_903,In_2027,In_574);
nand U904 (N_904,In_1499,In_909);
or U905 (N_905,In_2044,In_971);
xor U906 (N_906,In_925,In_1041);
nor U907 (N_907,In_1086,In_1430);
or U908 (N_908,In_2135,In_778);
nor U909 (N_909,In_1240,In_1987);
nand U910 (N_910,In_1496,In_328);
and U911 (N_911,In_711,In_367);
nor U912 (N_912,In_639,In_2118);
nand U913 (N_913,In_869,In_952);
nor U914 (N_914,In_1586,In_1852);
xor U915 (N_915,In_627,In_1376);
or U916 (N_916,In_2321,In_147);
nand U917 (N_917,In_1747,In_2429);
xnor U918 (N_918,In_1610,In_990);
or U919 (N_919,In_867,In_60);
nand U920 (N_920,In_1303,In_9);
nand U921 (N_921,In_939,In_415);
xnor U922 (N_922,In_1607,In_2303);
nor U923 (N_923,In_2309,In_1405);
nand U924 (N_924,In_537,In_1068);
xor U925 (N_925,In_1210,In_2058);
or U926 (N_926,In_1511,In_1715);
nor U927 (N_927,In_740,In_2081);
xor U928 (N_928,In_695,In_750);
xor U929 (N_929,In_53,In_1860);
nand U930 (N_930,In_2129,In_485);
xnor U931 (N_931,In_475,In_874);
xnor U932 (N_932,In_1436,In_896);
or U933 (N_933,In_1231,In_994);
and U934 (N_934,In_2066,In_68);
xnor U935 (N_935,In_1706,In_1980);
xor U936 (N_936,In_1694,In_871);
nor U937 (N_937,In_2085,In_449);
or U938 (N_938,In_2467,In_2350);
and U939 (N_939,In_2133,In_2101);
xor U940 (N_940,In_1990,In_1815);
and U941 (N_941,In_151,In_1737);
nand U942 (N_942,In_1672,In_1659);
or U943 (N_943,In_2402,In_734);
nand U944 (N_944,In_25,In_1965);
or U945 (N_945,In_1761,In_1344);
and U946 (N_946,In_1988,In_481);
xor U947 (N_947,In_2427,In_1703);
nand U948 (N_948,In_967,In_391);
or U949 (N_949,In_1420,In_822);
and U950 (N_950,In_316,In_2457);
nand U951 (N_951,In_2250,In_1626);
xor U952 (N_952,In_1196,In_1548);
or U953 (N_953,In_2051,In_571);
or U954 (N_954,In_2014,In_861);
and U955 (N_955,In_812,In_2263);
and U956 (N_956,In_383,In_170);
xor U957 (N_957,In_1004,In_2425);
nand U958 (N_958,In_1580,In_1718);
nor U959 (N_959,In_166,In_1190);
nand U960 (N_960,In_1810,In_1957);
xnor U961 (N_961,In_678,In_1113);
and U962 (N_962,In_2017,In_1746);
or U963 (N_963,In_2168,In_1745);
and U964 (N_964,In_666,In_1854);
xor U965 (N_965,In_208,In_1722);
or U966 (N_966,In_1140,In_1524);
nor U967 (N_967,In_1657,In_1878);
nor U968 (N_968,In_1681,In_2310);
xor U969 (N_969,In_1570,In_1389);
xnor U970 (N_970,In_807,In_1669);
or U971 (N_971,In_552,In_123);
and U972 (N_972,In_216,In_2450);
or U973 (N_973,In_232,In_288);
and U974 (N_974,In_292,In_2222);
and U975 (N_975,In_1904,In_290);
nor U976 (N_976,In_2374,In_1901);
or U977 (N_977,In_1225,In_80);
or U978 (N_978,In_504,In_761);
or U979 (N_979,In_584,In_412);
xor U980 (N_980,In_1616,In_1838);
xor U981 (N_981,In_1891,In_1769);
xor U982 (N_982,In_1403,In_82);
nand U983 (N_983,In_1091,In_536);
xor U984 (N_984,In_1880,In_2226);
and U985 (N_985,In_507,In_4);
xor U986 (N_986,In_629,In_1454);
and U987 (N_987,In_2403,In_1361);
or U988 (N_988,In_2,In_1638);
nor U989 (N_989,In_278,In_1535);
or U990 (N_990,In_1149,In_99);
nor U991 (N_991,In_1142,In_1467);
and U992 (N_992,In_1693,In_17);
xor U993 (N_993,In_1442,In_1270);
nor U994 (N_994,In_397,In_194);
xnor U995 (N_995,In_2276,In_1074);
and U996 (N_996,In_77,In_959);
xnor U997 (N_997,In_1911,In_1630);
nor U998 (N_998,In_865,In_19);
and U999 (N_999,In_1619,In_1645);
and U1000 (N_1000,In_1292,In_2406);
nor U1001 (N_1001,In_2054,In_1222);
xnor U1002 (N_1002,In_2237,In_1819);
and U1003 (N_1003,In_902,In_1683);
nor U1004 (N_1004,In_624,In_470);
nor U1005 (N_1005,In_424,In_300);
nand U1006 (N_1006,In_2198,In_1209);
and U1007 (N_1007,In_1035,In_600);
nor U1008 (N_1008,In_1306,In_315);
nand U1009 (N_1009,In_2158,In_660);
or U1010 (N_1010,In_1151,In_434);
or U1011 (N_1011,In_101,In_538);
nor U1012 (N_1012,In_233,In_1977);
nor U1013 (N_1013,In_2492,In_411);
or U1014 (N_1014,In_1831,In_745);
or U1015 (N_1015,In_1359,In_1287);
nand U1016 (N_1016,In_2452,In_1195);
and U1017 (N_1017,In_2024,In_598);
xor U1018 (N_1018,In_683,In_249);
xnor U1019 (N_1019,In_132,In_707);
nand U1020 (N_1020,In_1821,In_1188);
nand U1021 (N_1021,In_1274,In_1897);
nor U1022 (N_1022,In_1962,In_105);
nor U1023 (N_1023,In_2214,In_2451);
xor U1024 (N_1024,In_2089,In_508);
or U1025 (N_1025,In_1026,In_1652);
nor U1026 (N_1026,In_1740,In_2257);
xnor U1027 (N_1027,In_1620,In_2481);
and U1028 (N_1028,In_1032,In_1364);
nor U1029 (N_1029,In_1373,In_1098);
xnor U1030 (N_1030,In_325,In_1478);
xnor U1031 (N_1031,In_804,In_726);
nand U1032 (N_1032,In_272,In_1110);
and U1033 (N_1033,In_1260,In_554);
nand U1034 (N_1034,In_1133,In_2317);
or U1035 (N_1035,In_202,In_198);
nand U1036 (N_1036,In_2411,In_2057);
and U1037 (N_1037,In_529,In_1938);
xor U1038 (N_1038,In_605,In_1446);
nand U1039 (N_1039,In_2039,In_1154);
nand U1040 (N_1040,In_81,In_1858);
nand U1041 (N_1041,In_2086,In_1182);
nor U1042 (N_1042,In_985,In_1874);
and U1043 (N_1043,In_673,In_460);
or U1044 (N_1044,In_2143,In_363);
and U1045 (N_1045,In_2444,In_2313);
xor U1046 (N_1046,In_1307,In_1107);
or U1047 (N_1047,In_2001,In_312);
or U1048 (N_1048,In_1000,In_2396);
nor U1049 (N_1049,In_1144,In_1317);
and U1050 (N_1050,In_875,In_2070);
or U1051 (N_1051,In_1296,In_2028);
nor U1052 (N_1052,In_197,In_1731);
nor U1053 (N_1053,In_1528,In_2485);
or U1054 (N_1054,In_1575,In_1014);
and U1055 (N_1055,In_1288,In_1215);
or U1056 (N_1056,In_1741,In_436);
nor U1057 (N_1057,In_390,In_1170);
nor U1058 (N_1058,In_878,In_892);
and U1059 (N_1059,In_1999,In_1930);
or U1060 (N_1060,In_1380,In_877);
or U1061 (N_1061,In_1235,In_1368);
nor U1062 (N_1062,In_1106,In_2320);
nor U1063 (N_1063,In_2144,In_283);
and U1064 (N_1064,In_30,In_689);
or U1065 (N_1065,In_1702,In_324);
or U1066 (N_1066,In_1602,In_1646);
nor U1067 (N_1067,In_1148,In_2031);
or U1068 (N_1068,In_848,In_1308);
or U1069 (N_1069,In_1915,In_2099);
xnor U1070 (N_1070,In_2307,In_2181);
nor U1071 (N_1071,In_2375,In_546);
nand U1072 (N_1072,In_1409,In_1450);
or U1073 (N_1073,In_522,In_889);
nor U1074 (N_1074,In_561,In_641);
nand U1075 (N_1075,In_987,In_1679);
nor U1076 (N_1076,In_1379,In_1668);
nand U1077 (N_1077,In_2243,In_1830);
and U1078 (N_1078,In_1699,In_1811);
and U1079 (N_1079,In_951,In_238);
xnor U1080 (N_1080,In_1135,In_502);
and U1081 (N_1081,In_417,In_2015);
and U1082 (N_1082,In_1770,In_335);
nor U1083 (N_1083,In_2087,In_783);
or U1084 (N_1084,In_2106,In_1168);
and U1085 (N_1085,In_687,In_2405);
xor U1086 (N_1086,In_858,In_1435);
xor U1087 (N_1087,In_282,In_162);
nor U1088 (N_1088,In_1101,In_593);
nand U1089 (N_1089,In_1277,In_1763);
or U1090 (N_1090,In_2260,In_2364);
nand U1091 (N_1091,In_2231,In_2434);
nor U1092 (N_1092,In_547,In_516);
xnor U1093 (N_1093,In_2055,In_876);
or U1094 (N_1094,In_1583,In_556);
xnor U1095 (N_1095,In_440,In_1207);
and U1096 (N_1096,In_2030,In_1007);
nor U1097 (N_1097,In_2283,In_46);
or U1098 (N_1098,In_2095,In_934);
or U1099 (N_1099,In_1488,In_646);
or U1100 (N_1100,In_74,In_1216);
or U1101 (N_1101,In_815,In_515);
and U1102 (N_1102,In_510,In_625);
or U1103 (N_1103,In_744,In_231);
and U1104 (N_1104,In_567,In_603);
nand U1105 (N_1105,In_2306,In_270);
or U1106 (N_1106,In_1134,In_1861);
xnor U1107 (N_1107,In_42,In_1401);
or U1108 (N_1108,In_960,In_1682);
nand U1109 (N_1109,In_1298,In_347);
nor U1110 (N_1110,In_47,In_1836);
and U1111 (N_1111,In_1960,In_720);
nand U1112 (N_1112,In_611,In_1202);
or U1113 (N_1113,In_1782,In_2062);
or U1114 (N_1114,In_1485,In_575);
or U1115 (N_1115,In_1940,In_649);
or U1116 (N_1116,In_1964,In_296);
nor U1117 (N_1117,In_1749,In_2438);
nand U1118 (N_1118,In_2038,In_2340);
nor U1119 (N_1119,In_824,In_1941);
nor U1120 (N_1120,In_34,In_2245);
xnor U1121 (N_1121,In_692,In_1588);
nor U1122 (N_1122,In_1612,In_1343);
xor U1123 (N_1123,In_337,In_1633);
xor U1124 (N_1124,In_606,In_118);
xor U1125 (N_1125,In_998,In_1918);
nand U1126 (N_1126,In_129,In_1866);
nor U1127 (N_1127,In_2355,In_1117);
and U1128 (N_1128,In_1268,In_1220);
xor U1129 (N_1129,In_955,In_1329);
or U1130 (N_1130,In_319,In_93);
or U1131 (N_1131,In_399,In_953);
or U1132 (N_1132,In_1034,In_499);
and U1133 (N_1133,In_2021,In_444);
and U1134 (N_1134,In_1385,In_121);
nor U1135 (N_1135,In_1767,In_580);
nand U1136 (N_1136,In_751,In_1228);
nand U1137 (N_1137,In_821,In_1351);
xor U1138 (N_1138,In_602,In_1333);
xnor U1139 (N_1139,In_50,In_193);
or U1140 (N_1140,In_135,In_563);
nand U1141 (N_1141,In_1850,In_1928);
xnor U1142 (N_1142,In_1132,In_1465);
and U1143 (N_1143,In_2443,In_52);
nand U1144 (N_1144,In_1760,In_161);
nand U1145 (N_1145,In_355,In_1312);
or U1146 (N_1146,In_704,In_1611);
or U1147 (N_1147,In_1469,In_2123);
xnor U1148 (N_1148,In_2462,In_1377);
and U1149 (N_1149,In_1905,In_514);
xnor U1150 (N_1150,In_979,In_2159);
nor U1151 (N_1151,In_1331,In_1663);
xnor U1152 (N_1152,In_907,In_1194);
nand U1153 (N_1153,In_1933,In_2409);
xor U1154 (N_1154,In_1976,In_94);
and U1155 (N_1155,In_1219,In_1522);
and U1156 (N_1156,In_1060,In_549);
and U1157 (N_1157,In_152,In_840);
or U1158 (N_1158,In_2400,In_854);
nand U1159 (N_1159,In_2392,In_820);
xnor U1160 (N_1160,In_2138,In_276);
or U1161 (N_1161,In_1624,In_1480);
nand U1162 (N_1162,In_1096,In_366);
nor U1163 (N_1163,In_949,In_1603);
or U1164 (N_1164,In_1799,In_1354);
nor U1165 (N_1165,In_1972,In_1949);
nand U1166 (N_1166,In_1038,In_823);
or U1167 (N_1167,In_1001,In_940);
nand U1168 (N_1168,In_989,In_1793);
and U1169 (N_1169,In_1636,In_2002);
nand U1170 (N_1170,In_992,In_2489);
or U1171 (N_1171,In_1704,In_2249);
and U1172 (N_1172,In_1755,In_85);
xnor U1173 (N_1173,In_1743,In_851);
or U1174 (N_1174,In_86,In_548);
and U1175 (N_1175,In_863,In_1685);
xor U1176 (N_1176,In_303,In_1621);
and U1177 (N_1177,In_753,In_1365);
nor U1178 (N_1178,In_157,In_2125);
nor U1179 (N_1179,In_1730,In_244);
nand U1180 (N_1180,In_1259,In_490);
or U1181 (N_1181,In_1310,In_1708);
nand U1182 (N_1182,In_1023,In_2437);
nand U1183 (N_1183,In_1489,In_2384);
and U1184 (N_1184,In_2316,In_2127);
and U1185 (N_1185,In_218,In_2458);
nor U1186 (N_1186,In_1650,In_36);
nand U1187 (N_1187,In_1087,In_433);
xnor U1188 (N_1188,In_2413,In_623);
or U1189 (N_1189,In_2470,In_401);
and U1190 (N_1190,In_1751,In_1885);
and U1191 (N_1191,In_156,In_1125);
xnor U1192 (N_1192,In_58,In_115);
nand U1193 (N_1193,In_831,In_727);
nand U1194 (N_1194,In_1825,In_2336);
nand U1195 (N_1195,In_1367,In_2068);
nor U1196 (N_1196,In_887,In_297);
or U1197 (N_1197,In_2253,In_2251);
nor U1198 (N_1198,In_2331,In_20);
nor U1199 (N_1199,In_1840,In_2131);
and U1200 (N_1200,In_57,In_2075);
xor U1201 (N_1201,In_1660,In_610);
or U1202 (N_1202,In_146,In_293);
nor U1203 (N_1203,In_1427,In_177);
or U1204 (N_1204,In_577,In_1921);
nor U1205 (N_1205,In_1844,In_35);
nor U1206 (N_1206,In_2140,In_791);
xor U1207 (N_1207,In_95,In_1754);
nand U1208 (N_1208,In_1882,In_1676);
nor U1209 (N_1209,In_755,In_2319);
xor U1210 (N_1210,In_1262,In_841);
xnor U1211 (N_1211,In_1956,In_259);
and U1212 (N_1212,In_2266,In_1315);
nor U1213 (N_1213,In_736,In_116);
and U1214 (N_1214,In_2498,In_1849);
xor U1215 (N_1215,In_1628,In_717);
nand U1216 (N_1216,In_530,In_2395);
and U1217 (N_1217,In_371,In_1884);
and U1218 (N_1218,In_1031,In_808);
or U1219 (N_1219,In_1015,In_1692);
nand U1220 (N_1220,In_2203,In_2043);
or U1221 (N_1221,In_2284,In_1788);
nor U1222 (N_1222,In_2247,In_438);
nor U1223 (N_1223,In_1085,In_1922);
xnor U1224 (N_1224,In_445,In_286);
nor U1225 (N_1225,In_1275,In_2339);
nor U1226 (N_1226,In_1680,In_1337);
and U1227 (N_1227,In_888,In_735);
and U1228 (N_1228,In_279,In_795);
nor U1229 (N_1229,In_427,In_1241);
and U1230 (N_1230,In_2052,In_164);
nor U1231 (N_1231,In_1503,In_1061);
or U1232 (N_1232,In_1372,In_1727);
nand U1233 (N_1233,In_928,In_632);
nand U1234 (N_1234,In_188,In_1723);
nor U1235 (N_1235,In_917,In_2482);
or U1236 (N_1236,In_195,In_633);
nand U1237 (N_1237,In_1477,In_1309);
and U1238 (N_1238,In_1695,In_2210);
nor U1239 (N_1239,In_2387,In_1239);
xor U1240 (N_1240,In_903,In_910);
xnor U1241 (N_1241,In_70,In_963);
nor U1242 (N_1242,In_111,In_1456);
or U1243 (N_1243,In_882,In_204);
xor U1244 (N_1244,In_2465,In_1721);
nand U1245 (N_1245,In_209,In_1130);
or U1246 (N_1246,In_2128,In_881);
or U1247 (N_1247,In_338,In_2233);
nand U1248 (N_1248,In_1812,In_1230);
nor U1249 (N_1249,In_1757,In_589);
and U1250 (N_1250,N_846,N_14);
xor U1251 (N_1251,N_377,N_6);
and U1252 (N_1252,N_1210,N_667);
or U1253 (N_1253,N_543,N_1061);
or U1254 (N_1254,N_727,N_291);
and U1255 (N_1255,N_1111,N_872);
or U1256 (N_1256,N_970,N_213);
xor U1257 (N_1257,N_295,N_535);
nor U1258 (N_1258,N_677,N_761);
or U1259 (N_1259,N_626,N_991);
and U1260 (N_1260,N_1010,N_865);
nor U1261 (N_1261,N_25,N_705);
nand U1262 (N_1262,N_262,N_431);
xor U1263 (N_1263,N_94,N_1161);
and U1264 (N_1264,N_1186,N_1194);
or U1265 (N_1265,N_985,N_1166);
or U1266 (N_1266,N_1027,N_160);
nand U1267 (N_1267,N_510,N_251);
xor U1268 (N_1268,N_249,N_828);
and U1269 (N_1269,N_695,N_1047);
or U1270 (N_1270,N_967,N_1172);
nand U1271 (N_1271,N_1245,N_495);
or U1272 (N_1272,N_1006,N_1115);
xnor U1273 (N_1273,N_276,N_185);
and U1274 (N_1274,N_379,N_837);
xor U1275 (N_1275,N_1135,N_747);
nor U1276 (N_1276,N_33,N_516);
and U1277 (N_1277,N_104,N_1171);
and U1278 (N_1278,N_390,N_1048);
and U1279 (N_1279,N_324,N_758);
or U1280 (N_1280,N_757,N_419);
nand U1281 (N_1281,N_915,N_1050);
xor U1282 (N_1282,N_42,N_670);
and U1283 (N_1283,N_69,N_898);
or U1284 (N_1284,N_437,N_129);
nor U1285 (N_1285,N_1080,N_341);
nor U1286 (N_1286,N_114,N_525);
and U1287 (N_1287,N_561,N_423);
and U1288 (N_1288,N_965,N_186);
or U1289 (N_1289,N_834,N_572);
nand U1290 (N_1290,N_247,N_123);
xor U1291 (N_1291,N_763,N_322);
or U1292 (N_1292,N_170,N_317);
or U1293 (N_1293,N_449,N_902);
or U1294 (N_1294,N_434,N_179);
xor U1295 (N_1295,N_564,N_149);
or U1296 (N_1296,N_63,N_1165);
and U1297 (N_1297,N_1244,N_526);
nand U1298 (N_1298,N_367,N_503);
xor U1299 (N_1299,N_1219,N_522);
nor U1300 (N_1300,N_190,N_376);
nand U1301 (N_1301,N_31,N_987);
nor U1302 (N_1302,N_1151,N_323);
or U1303 (N_1303,N_571,N_785);
nand U1304 (N_1304,N_1109,N_24);
and U1305 (N_1305,N_632,N_254);
nand U1306 (N_1306,N_1126,N_1018);
or U1307 (N_1307,N_118,N_821);
nor U1308 (N_1308,N_189,N_456);
nand U1309 (N_1309,N_82,N_614);
or U1310 (N_1310,N_120,N_820);
xnor U1311 (N_1311,N_781,N_91);
or U1312 (N_1312,N_601,N_471);
and U1313 (N_1313,N_266,N_839);
nand U1314 (N_1314,N_863,N_303);
or U1315 (N_1315,N_777,N_984);
or U1316 (N_1316,N_1236,N_11);
xor U1317 (N_1317,N_133,N_589);
xor U1318 (N_1318,N_1224,N_1076);
xor U1319 (N_1319,N_922,N_235);
or U1320 (N_1320,N_387,N_294);
or U1321 (N_1321,N_76,N_335);
or U1322 (N_1322,N_732,N_244);
xnor U1323 (N_1323,N_126,N_722);
or U1324 (N_1324,N_859,N_255);
nand U1325 (N_1325,N_893,N_829);
and U1326 (N_1326,N_48,N_443);
or U1327 (N_1327,N_1183,N_938);
and U1328 (N_1328,N_80,N_130);
nor U1329 (N_1329,N_708,N_1003);
and U1330 (N_1330,N_272,N_502);
and U1331 (N_1331,N_470,N_584);
xnor U1332 (N_1332,N_752,N_992);
xnor U1333 (N_1333,N_340,N_441);
or U1334 (N_1334,N_1130,N_674);
xor U1335 (N_1335,N_980,N_1137);
xnor U1336 (N_1336,N_982,N_227);
xnor U1337 (N_1337,N_765,N_813);
and U1338 (N_1338,N_39,N_201);
and U1339 (N_1339,N_1201,N_857);
nor U1340 (N_1340,N_814,N_1041);
or U1341 (N_1341,N_1203,N_351);
or U1342 (N_1342,N_690,N_246);
or U1343 (N_1343,N_669,N_110);
or U1344 (N_1344,N_523,N_689);
or U1345 (N_1345,N_337,N_856);
nand U1346 (N_1346,N_274,N_256);
xnor U1347 (N_1347,N_1097,N_299);
and U1348 (N_1348,N_326,N_1150);
xor U1349 (N_1349,N_1187,N_458);
and U1350 (N_1350,N_622,N_875);
xor U1351 (N_1351,N_306,N_477);
nand U1352 (N_1352,N_1182,N_993);
nand U1353 (N_1353,N_480,N_1146);
xnor U1354 (N_1354,N_701,N_579);
or U1355 (N_1355,N_278,N_842);
nand U1356 (N_1356,N_873,N_71);
nor U1357 (N_1357,N_840,N_888);
nor U1358 (N_1358,N_148,N_233);
and U1359 (N_1359,N_806,N_1051);
xnor U1360 (N_1360,N_529,N_412);
nand U1361 (N_1361,N_1237,N_1232);
and U1362 (N_1362,N_655,N_1230);
nand U1363 (N_1363,N_56,N_527);
nand U1364 (N_1364,N_35,N_457);
xnor U1365 (N_1365,N_767,N_729);
and U1366 (N_1366,N_287,N_958);
nor U1367 (N_1367,N_969,N_188);
nor U1368 (N_1368,N_800,N_75);
and U1369 (N_1369,N_688,N_1246);
and U1370 (N_1370,N_1247,N_772);
nand U1371 (N_1371,N_311,N_1148);
nor U1372 (N_1372,N_1113,N_1114);
or U1373 (N_1373,N_74,N_1024);
or U1374 (N_1374,N_560,N_325);
and U1375 (N_1375,N_230,N_264);
nand U1376 (N_1376,N_650,N_436);
nor U1377 (N_1377,N_21,N_1167);
or U1378 (N_1378,N_774,N_136);
xor U1379 (N_1379,N_803,N_496);
nor U1380 (N_1380,N_330,N_1086);
nand U1381 (N_1381,N_191,N_962);
or U1382 (N_1382,N_1128,N_103);
xor U1383 (N_1383,N_656,N_903);
nand U1384 (N_1384,N_716,N_858);
nor U1385 (N_1385,N_432,N_370);
xor U1386 (N_1386,N_1215,N_977);
xor U1387 (N_1387,N_548,N_55);
and U1388 (N_1388,N_1158,N_428);
xnor U1389 (N_1389,N_811,N_1168);
nand U1390 (N_1390,N_906,N_138);
xnor U1391 (N_1391,N_240,N_1071);
nand U1392 (N_1392,N_1191,N_223);
xor U1393 (N_1393,N_511,N_675);
nand U1394 (N_1394,N_666,N_485);
and U1395 (N_1395,N_259,N_745);
nor U1396 (N_1396,N_596,N_349);
nand U1397 (N_1397,N_651,N_680);
nand U1398 (N_1398,N_1132,N_1057);
xor U1399 (N_1399,N_155,N_146);
or U1400 (N_1400,N_1089,N_88);
or U1401 (N_1401,N_755,N_1004);
nand U1402 (N_1402,N_192,N_819);
xor U1403 (N_1403,N_196,N_494);
nor U1404 (N_1404,N_792,N_265);
xnor U1405 (N_1405,N_345,N_979);
or U1406 (N_1406,N_884,N_79);
and U1407 (N_1407,N_200,N_113);
xor U1408 (N_1408,N_162,N_1120);
xor U1409 (N_1409,N_1216,N_93);
xor U1410 (N_1410,N_288,N_253);
nand U1411 (N_1411,N_960,N_771);
nor U1412 (N_1412,N_8,N_1016);
and U1413 (N_1413,N_617,N_252);
xor U1414 (N_1414,N_1179,N_211);
nand U1415 (N_1415,N_1122,N_862);
nand U1416 (N_1416,N_1032,N_1222);
or U1417 (N_1417,N_112,N_1005);
and U1418 (N_1418,N_871,N_703);
nor U1419 (N_1419,N_1056,N_362);
nand U1420 (N_1420,N_1094,N_115);
nor U1421 (N_1421,N_1196,N_382);
nor U1422 (N_1422,N_352,N_60);
or U1423 (N_1423,N_229,N_1243);
and U1424 (N_1424,N_989,N_228);
nor U1425 (N_1425,N_484,N_887);
nor U1426 (N_1426,N_163,N_723);
nor U1427 (N_1427,N_1026,N_296);
or U1428 (N_1428,N_70,N_381);
and U1429 (N_1429,N_389,N_835);
or U1430 (N_1430,N_972,N_877);
nand U1431 (N_1431,N_861,N_649);
xor U1432 (N_1432,N_715,N_1);
or U1433 (N_1433,N_425,N_678);
nand U1434 (N_1434,N_1140,N_530);
xnor U1435 (N_1435,N_391,N_751);
nor U1436 (N_1436,N_445,N_1117);
nor U1437 (N_1437,N_718,N_316);
or U1438 (N_1438,N_927,N_911);
and U1439 (N_1439,N_99,N_409);
nand U1440 (N_1440,N_573,N_1031);
nand U1441 (N_1441,N_67,N_1014);
and U1442 (N_1442,N_929,N_217);
nor U1443 (N_1443,N_889,N_248);
nand U1444 (N_1444,N_706,N_999);
nor U1445 (N_1445,N_463,N_810);
nand U1446 (N_1446,N_1066,N_1133);
xor U1447 (N_1447,N_1233,N_838);
or U1448 (N_1448,N_1184,N_795);
nor U1449 (N_1449,N_1019,N_292);
or U1450 (N_1450,N_822,N_427);
or U1451 (N_1451,N_479,N_372);
nor U1452 (N_1452,N_194,N_77);
or U1453 (N_1453,N_284,N_68);
or U1454 (N_1454,N_426,N_446);
nand U1455 (N_1455,N_725,N_1157);
nor U1456 (N_1456,N_1017,N_654);
nor U1457 (N_1457,N_386,N_321);
nand U1458 (N_1458,N_1044,N_940);
and U1459 (N_1459,N_279,N_764);
xor U1460 (N_1460,N_853,N_1223);
nand U1461 (N_1461,N_1038,N_562);
or U1462 (N_1462,N_743,N_1144);
and U1463 (N_1463,N_38,N_275);
nand U1464 (N_1464,N_676,N_528);
nand U1465 (N_1465,N_894,N_1176);
and U1466 (N_1466,N_490,N_300);
xnor U1467 (N_1467,N_825,N_1107);
and U1468 (N_1468,N_717,N_1065);
nand U1469 (N_1469,N_2,N_553);
nand U1470 (N_1470,N_180,N_408);
and U1471 (N_1471,N_1073,N_12);
xor U1472 (N_1472,N_239,N_760);
and U1473 (N_1473,N_796,N_65);
xor U1474 (N_1474,N_257,N_1082);
and U1475 (N_1475,N_815,N_554);
and U1476 (N_1476,N_360,N_610);
and U1477 (N_1477,N_152,N_633);
nor U1478 (N_1478,N_241,N_1037);
xor U1479 (N_1479,N_867,N_195);
and U1480 (N_1480,N_1213,N_157);
and U1481 (N_1481,N_1204,N_687);
nor U1482 (N_1482,N_712,N_1081);
and U1483 (N_1483,N_413,N_1209);
nor U1484 (N_1484,N_164,N_890);
xnor U1485 (N_1485,N_250,N_1131);
xnor U1486 (N_1486,N_621,N_599);
and U1487 (N_1487,N_231,N_1054);
and U1488 (N_1488,N_559,N_462);
nand U1489 (N_1489,N_1202,N_1188);
or U1490 (N_1490,N_624,N_280);
and U1491 (N_1491,N_619,N_310);
nand U1492 (N_1492,N_547,N_424);
nand U1493 (N_1493,N_836,N_96);
nand U1494 (N_1494,N_396,N_62);
and U1495 (N_1495,N_684,N_245);
and U1496 (N_1496,N_101,N_492);
xor U1497 (N_1497,N_892,N_869);
and U1498 (N_1498,N_19,N_710);
xor U1499 (N_1499,N_134,N_711);
xnor U1500 (N_1500,N_730,N_1100);
nor U1501 (N_1501,N_841,N_378);
nor U1502 (N_1502,N_406,N_1022);
nand U1503 (N_1503,N_1160,N_883);
or U1504 (N_1504,N_896,N_878);
and U1505 (N_1505,N_639,N_150);
or U1506 (N_1506,N_879,N_974);
or U1507 (N_1507,N_779,N_145);
or U1508 (N_1508,N_585,N_786);
or U1509 (N_1509,N_482,N_753);
xnor U1510 (N_1510,N_519,N_84);
and U1511 (N_1511,N_583,N_53);
xnor U1512 (N_1512,N_1118,N_125);
nor U1513 (N_1513,N_997,N_1058);
and U1514 (N_1514,N_916,N_996);
xor U1515 (N_1515,N_580,N_305);
xor U1516 (N_1516,N_66,N_541);
nand U1517 (N_1517,N_491,N_1075);
or U1518 (N_1518,N_334,N_1012);
or U1519 (N_1519,N_85,N_1108);
and U1520 (N_1520,N_313,N_385);
nand U1521 (N_1521,N_224,N_147);
or U1522 (N_1522,N_269,N_661);
and U1523 (N_1523,N_595,N_221);
or U1524 (N_1524,N_934,N_348);
nor U1525 (N_1525,N_620,N_1025);
and U1526 (N_1526,N_364,N_1116);
xor U1527 (N_1527,N_986,N_741);
or U1528 (N_1528,N_100,N_1152);
and U1529 (N_1529,N_640,N_1242);
or U1530 (N_1530,N_860,N_225);
nor U1531 (N_1531,N_344,N_532);
nor U1532 (N_1532,N_176,N_536);
and U1533 (N_1533,N_631,N_108);
or U1534 (N_1534,N_812,N_435);
nor U1535 (N_1535,N_1072,N_117);
or U1536 (N_1536,N_1175,N_181);
and U1537 (N_1537,N_570,N_401);
or U1538 (N_1538,N_1154,N_628);
and U1539 (N_1539,N_173,N_606);
nand U1540 (N_1540,N_286,N_565);
or U1541 (N_1541,N_368,N_602);
nand U1542 (N_1542,N_816,N_801);
nor U1543 (N_1543,N_608,N_885);
xnor U1544 (N_1544,N_923,N_1009);
and U1545 (N_1545,N_618,N_928);
and U1546 (N_1546,N_951,N_954);
nand U1547 (N_1547,N_270,N_931);
or U1548 (N_1548,N_556,N_1207);
or U1549 (N_1549,N_144,N_833);
or U1550 (N_1550,N_913,N_558);
or U1551 (N_1551,N_478,N_302);
nand U1552 (N_1552,N_749,N_549);
or U1553 (N_1553,N_609,N_607);
nor U1554 (N_1554,N_486,N_216);
or U1555 (N_1555,N_307,N_23);
nor U1556 (N_1556,N_643,N_944);
xnor U1557 (N_1557,N_679,N_1226);
and U1558 (N_1558,N_460,N_98);
or U1559 (N_1559,N_37,N_778);
nand U1560 (N_1560,N_696,N_959);
nand U1561 (N_1561,N_1104,N_36);
nand U1562 (N_1562,N_327,N_92);
xor U1563 (N_1563,N_740,N_537);
nand U1564 (N_1564,N_612,N_346);
nor U1565 (N_1565,N_1069,N_1198);
nand U1566 (N_1566,N_210,N_475);
and U1567 (N_1567,N_489,N_122);
xnor U1568 (N_1568,N_673,N_635);
xor U1569 (N_1569,N_399,N_588);
xnor U1570 (N_1570,N_1021,N_693);
and U1571 (N_1571,N_581,N_1033);
or U1572 (N_1572,N_577,N_880);
xnor U1573 (N_1573,N_826,N_282);
nand U1574 (N_1574,N_668,N_868);
and U1575 (N_1575,N_440,N_1164);
and U1576 (N_1576,N_105,N_158);
xnor U1577 (N_1577,N_289,N_1229);
and U1578 (N_1578,N_1134,N_605);
nor U1579 (N_1579,N_16,N_59);
xnor U1580 (N_1580,N_51,N_339);
and U1581 (N_1581,N_1249,N_182);
and U1582 (N_1582,N_719,N_882);
and U1583 (N_1583,N_178,N_314);
nand U1584 (N_1584,N_512,N_402);
nand U1585 (N_1585,N_555,N_907);
nor U1586 (N_1586,N_756,N_15);
nand U1587 (N_1587,N_950,N_817);
nand U1588 (N_1588,N_488,N_198);
or U1589 (N_1589,N_942,N_333);
nand U1590 (N_1590,N_135,N_183);
or U1591 (N_1591,N_234,N_363);
nand U1592 (N_1592,N_636,N_964);
xor U1593 (N_1593,N_1199,N_226);
and U1594 (N_1594,N_790,N_121);
nand U1595 (N_1595,N_430,N_215);
nand U1596 (N_1596,N_78,N_1068);
or U1597 (N_1597,N_45,N_648);
and U1598 (N_1598,N_901,N_1074);
nand U1599 (N_1599,N_754,N_169);
nor U1600 (N_1600,N_976,N_943);
or U1601 (N_1601,N_593,N_1055);
and U1602 (N_1602,N_941,N_1177);
and U1603 (N_1603,N_27,N_634);
and U1604 (N_1604,N_805,N_769);
or U1605 (N_1605,N_1007,N_507);
or U1606 (N_1606,N_404,N_797);
xnor U1607 (N_1607,N_694,N_855);
nor U1608 (N_1608,N_1185,N_933);
nand U1609 (N_1609,N_193,N_1149);
nand U1610 (N_1610,N_874,N_140);
nand U1611 (N_1611,N_52,N_653);
nor U1612 (N_1612,N_768,N_1060);
nor U1613 (N_1613,N_920,N_737);
nor U1614 (N_1614,N_657,N_1178);
nor U1615 (N_1615,N_998,N_707);
or U1616 (N_1616,N_124,N_870);
nor U1617 (N_1617,N_83,N_736);
and U1618 (N_1618,N_469,N_864);
or U1619 (N_1619,N_1112,N_1241);
nor U1620 (N_1620,N_1101,N_1227);
xor U1621 (N_1621,N_414,N_539);
and U1622 (N_1622,N_319,N_338);
xnor U1623 (N_1623,N_1211,N_1091);
nand U1624 (N_1624,N_500,N_692);
nor U1625 (N_1625,N_107,N_205);
or U1626 (N_1626,N_646,N_538);
nor U1627 (N_1627,N_328,N_1136);
and U1628 (N_1628,N_935,N_791);
or U1629 (N_1629,N_1141,N_1052);
nand U1630 (N_1630,N_831,N_154);
nand U1631 (N_1631,N_1093,N_422);
nor U1632 (N_1632,N_468,N_297);
nor U1633 (N_1633,N_899,N_1142);
nor U1634 (N_1634,N_709,N_930);
nand U1635 (N_1635,N_798,N_905);
or U1636 (N_1636,N_904,N_1020);
nand U1637 (N_1637,N_29,N_637);
nor U1638 (N_1638,N_1067,N_397);
or U1639 (N_1639,N_347,N_968);
or U1640 (N_1640,N_127,N_1239);
nor U1641 (N_1641,N_283,N_1013);
nor U1642 (N_1642,N_652,N_1042);
nor U1643 (N_1643,N_383,N_542);
nor U1644 (N_1644,N_320,N_973);
nor U1645 (N_1645,N_481,N_533);
or U1646 (N_1646,N_474,N_1124);
nand U1647 (N_1647,N_442,N_735);
nand U1648 (N_1648,N_770,N_1192);
or U1649 (N_1649,N_983,N_551);
or U1650 (N_1650,N_848,N_243);
xor U1651 (N_1651,N_591,N_844);
nor U1652 (N_1652,N_220,N_128);
or U1653 (N_1653,N_616,N_452);
and U1654 (N_1654,N_809,N_1218);
nor U1655 (N_1655,N_197,N_594);
or U1656 (N_1656,N_876,N_260);
or U1657 (N_1657,N_659,N_28);
nor U1658 (N_1658,N_1087,N_937);
and U1659 (N_1659,N_361,N_1046);
nor U1660 (N_1660,N_611,N_517);
or U1661 (N_1661,N_881,N_665);
nand U1662 (N_1662,N_1214,N_132);
nand U1663 (N_1663,N_780,N_174);
nor U1664 (N_1664,N_1205,N_358);
xnor U1665 (N_1665,N_783,N_26);
nor U1666 (N_1666,N_209,N_1119);
xor U1667 (N_1667,N_411,N_1099);
nand U1668 (N_1668,N_20,N_949);
xor U1669 (N_1669,N_116,N_32);
and U1670 (N_1670,N_966,N_1153);
nand U1671 (N_1671,N_569,N_1079);
nand U1672 (N_1672,N_851,N_476);
or U1673 (N_1673,N_1083,N_331);
nor U1674 (N_1674,N_22,N_978);
and U1675 (N_1675,N_208,N_952);
nor U1676 (N_1676,N_1156,N_623);
xor U1677 (N_1677,N_1036,N_355);
or U1678 (N_1678,N_1039,N_308);
xor U1679 (N_1679,N_762,N_273);
nor U1680 (N_1680,N_945,N_1129);
or U1681 (N_1681,N_374,N_318);
xor U1682 (N_1682,N_461,N_604);
nor U1683 (N_1683,N_714,N_720);
or U1684 (N_1684,N_17,N_1001);
xnor U1685 (N_1685,N_1125,N_142);
nor U1686 (N_1686,N_237,N_849);
or U1687 (N_1687,N_172,N_955);
xnor U1688 (N_1688,N_567,N_336);
or U1689 (N_1689,N_369,N_702);
nand U1690 (N_1690,N_1174,N_137);
nor U1691 (N_1691,N_418,N_49);
and U1692 (N_1692,N_293,N_1049);
and U1693 (N_1693,N_151,N_451);
nor U1694 (N_1694,N_660,N_784);
or U1695 (N_1695,N_663,N_1085);
nand U1696 (N_1696,N_501,N_699);
xnor U1697 (N_1697,N_924,N_773);
xor U1698 (N_1698,N_1028,N_359);
and U1699 (N_1699,N_782,N_1139);
and U1700 (N_1700,N_615,N_932);
nand U1701 (N_1701,N_662,N_455);
xor U1702 (N_1702,N_546,N_373);
nor U1703 (N_1703,N_18,N_947);
nand U1704 (N_1704,N_9,N_1240);
and U1705 (N_1705,N_1189,N_281);
or U1706 (N_1706,N_177,N_214);
or U1707 (N_1707,N_854,N_592);
xor U1708 (N_1708,N_953,N_990);
and U1709 (N_1709,N_698,N_1059);
nand U1710 (N_1710,N_513,N_398);
nand U1711 (N_1711,N_41,N_384);
or U1712 (N_1712,N_1220,N_353);
nor U1713 (N_1713,N_356,N_1062);
or U1714 (N_1714,N_1238,N_354);
xnor U1715 (N_1715,N_392,N_776);
or U1716 (N_1716,N_166,N_312);
xnor U1717 (N_1717,N_212,N_102);
or U1718 (N_1718,N_832,N_645);
xor U1719 (N_1719,N_738,N_438);
nand U1720 (N_1720,N_1181,N_1180);
and U1721 (N_1721,N_1040,N_697);
nor U1722 (N_1722,N_1197,N_417);
or U1723 (N_1723,N_957,N_1231);
nor U1724 (N_1724,N_1088,N_498);
or U1725 (N_1725,N_429,N_165);
and U1726 (N_1726,N_808,N_199);
and U1727 (N_1727,N_590,N_380);
xor U1728 (N_1728,N_683,N_713);
and U1729 (N_1729,N_1173,N_202);
nor U1730 (N_1730,N_731,N_818);
nor U1731 (N_1731,N_388,N_603);
nor U1732 (N_1732,N_171,N_1015);
and U1733 (N_1733,N_975,N_444);
nand U1734 (N_1734,N_948,N_726);
nor U1735 (N_1735,N_242,N_1063);
nor U1736 (N_1736,N_671,N_748);
and U1737 (N_1737,N_421,N_95);
and U1738 (N_1738,N_206,N_578);
and U1739 (N_1739,N_161,N_824);
or U1740 (N_1740,N_1200,N_664);
and U1741 (N_1741,N_845,N_1206);
nand U1742 (N_1742,N_557,N_298);
or U1743 (N_1743,N_219,N_89);
nor U1744 (N_1744,N_682,N_46);
nand U1745 (N_1745,N_685,N_897);
nand U1746 (N_1746,N_375,N_1070);
and U1747 (N_1747,N_971,N_1162);
or U1748 (N_1748,N_919,N_90);
nor U1749 (N_1749,N_64,N_804);
xor U1750 (N_1750,N_0,N_420);
and U1751 (N_1751,N_97,N_742);
xnor U1752 (N_1752,N_153,N_823);
or U1753 (N_1753,N_400,N_1092);
or U1754 (N_1754,N_534,N_1084);
nor U1755 (N_1755,N_454,N_936);
xor U1756 (N_1756,N_1011,N_1155);
and U1757 (N_1757,N_5,N_544);
and U1758 (N_1758,N_540,N_1234);
and U1759 (N_1759,N_908,N_691);
nor U1760 (N_1760,N_733,N_439);
and U1761 (N_1761,N_1221,N_416);
or U1762 (N_1762,N_850,N_1110);
or U1763 (N_1763,N_1102,N_1127);
nor U1764 (N_1764,N_520,N_1235);
and U1765 (N_1765,N_600,N_1090);
xor U1766 (N_1766,N_61,N_766);
nand U1767 (N_1767,N_509,N_1002);
xor U1768 (N_1768,N_910,N_410);
or U1769 (N_1769,N_1123,N_141);
or U1770 (N_1770,N_582,N_263);
nand U1771 (N_1771,N_415,N_775);
or U1772 (N_1772,N_72,N_750);
nor U1773 (N_1773,N_939,N_506);
xnor U1774 (N_1774,N_487,N_946);
xor U1775 (N_1775,N_1143,N_1217);
nor U1776 (N_1776,N_1169,N_309);
and U1777 (N_1777,N_1208,N_1008);
nor U1778 (N_1778,N_448,N_552);
and U1779 (N_1779,N_86,N_568);
and U1780 (N_1780,N_1105,N_627);
nor U1781 (N_1781,N_143,N_566);
and U1782 (N_1782,N_357,N_799);
nand U1783 (N_1783,N_13,N_641);
and U1784 (N_1784,N_586,N_1023);
and U1785 (N_1785,N_638,N_258);
nand U1786 (N_1786,N_261,N_956);
and U1787 (N_1787,N_10,N_268);
nand U1788 (N_1788,N_43,N_493);
nand U1789 (N_1789,N_315,N_497);
xor U1790 (N_1790,N_73,N_472);
xnor U1791 (N_1791,N_734,N_483);
nand U1792 (N_1792,N_1121,N_587);
nand U1793 (N_1793,N_1193,N_1043);
nor U1794 (N_1794,N_746,N_508);
or U1795 (N_1795,N_290,N_332);
and U1796 (N_1796,N_914,N_304);
and U1797 (N_1797,N_886,N_788);
or U1798 (N_1798,N_629,N_111);
or U1799 (N_1799,N_681,N_630);
or U1800 (N_1800,N_827,N_613);
nor U1801 (N_1801,N_505,N_222);
xor U1802 (N_1802,N_1163,N_672);
xnor U1803 (N_1803,N_598,N_1248);
nor U1804 (N_1804,N_658,N_405);
and U1805 (N_1805,N_30,N_1053);
or U1806 (N_1806,N_891,N_184);
nand U1807 (N_1807,N_866,N_895);
nor U1808 (N_1808,N_1098,N_285);
or U1809 (N_1809,N_47,N_644);
xnor U1810 (N_1810,N_407,N_218);
nor U1811 (N_1811,N_504,N_329);
nand U1812 (N_1812,N_156,N_794);
nor U1813 (N_1813,N_515,N_203);
nand U1814 (N_1814,N_1064,N_433);
or U1815 (N_1815,N_807,N_57);
nor U1816 (N_1816,N_1029,N_518);
or U1817 (N_1817,N_106,N_550);
or U1818 (N_1818,N_464,N_1077);
nor U1819 (N_1819,N_925,N_917);
nor U1820 (N_1820,N_238,N_350);
nor U1821 (N_1821,N_395,N_1000);
and U1822 (N_1822,N_58,N_1145);
or U1823 (N_1823,N_759,N_54);
xor U1824 (N_1824,N_575,N_921);
or U1825 (N_1825,N_1228,N_342);
nand U1826 (N_1826,N_403,N_721);
nor U1827 (N_1827,N_207,N_447);
xor U1828 (N_1828,N_843,N_119);
xor U1829 (N_1829,N_465,N_1096);
and U1830 (N_1830,N_1035,N_187);
xor U1831 (N_1831,N_909,N_236);
xor U1832 (N_1832,N_686,N_40);
nor U1833 (N_1833,N_175,N_597);
xor U1834 (N_1834,N_1106,N_1078);
nor U1835 (N_1835,N_704,N_459);
nand U1836 (N_1836,N_301,N_34);
and U1837 (N_1837,N_830,N_109);
or U1838 (N_1838,N_728,N_576);
nand U1839 (N_1839,N_918,N_277);
nor U1840 (N_1840,N_524,N_744);
and U1841 (N_1841,N_521,N_3);
or U1842 (N_1842,N_981,N_563);
nor U1843 (N_1843,N_168,N_473);
xor U1844 (N_1844,N_994,N_139);
xnor U1845 (N_1845,N_204,N_724);
nand U1846 (N_1846,N_531,N_499);
nor U1847 (N_1847,N_271,N_1034);
xnor U1848 (N_1848,N_394,N_802);
nor U1849 (N_1849,N_466,N_1045);
or U1850 (N_1850,N_988,N_50);
nor U1851 (N_1851,N_467,N_1095);
or U1852 (N_1852,N_625,N_739);
nor U1853 (N_1853,N_545,N_1195);
nand U1854 (N_1854,N_232,N_453);
and U1855 (N_1855,N_1030,N_167);
and U1856 (N_1856,N_371,N_700);
xnor U1857 (N_1857,N_81,N_789);
nand U1858 (N_1858,N_7,N_574);
xor U1859 (N_1859,N_1170,N_963);
nor U1860 (N_1860,N_4,N_131);
nand U1861 (N_1861,N_1159,N_793);
nor U1862 (N_1862,N_1190,N_365);
or U1863 (N_1863,N_995,N_44);
and U1864 (N_1864,N_926,N_1103);
and U1865 (N_1865,N_87,N_852);
or U1866 (N_1866,N_900,N_1147);
nor U1867 (N_1867,N_393,N_514);
or U1868 (N_1868,N_647,N_642);
nand U1869 (N_1869,N_159,N_366);
or U1870 (N_1870,N_343,N_1138);
xnor U1871 (N_1871,N_961,N_1225);
xor U1872 (N_1872,N_267,N_1212);
and U1873 (N_1873,N_787,N_912);
nor U1874 (N_1874,N_847,N_450);
or U1875 (N_1875,N_753,N_356);
or U1876 (N_1876,N_893,N_359);
or U1877 (N_1877,N_280,N_1097);
xor U1878 (N_1878,N_1197,N_30);
and U1879 (N_1879,N_863,N_362);
nand U1880 (N_1880,N_958,N_508);
xor U1881 (N_1881,N_1181,N_128);
and U1882 (N_1882,N_115,N_1149);
and U1883 (N_1883,N_681,N_712);
or U1884 (N_1884,N_505,N_942);
nor U1885 (N_1885,N_1245,N_181);
nor U1886 (N_1886,N_463,N_918);
nor U1887 (N_1887,N_957,N_1248);
nand U1888 (N_1888,N_37,N_882);
and U1889 (N_1889,N_850,N_241);
and U1890 (N_1890,N_857,N_272);
nor U1891 (N_1891,N_393,N_96);
or U1892 (N_1892,N_1101,N_30);
or U1893 (N_1893,N_1024,N_224);
or U1894 (N_1894,N_307,N_857);
nand U1895 (N_1895,N_437,N_683);
xor U1896 (N_1896,N_747,N_498);
nand U1897 (N_1897,N_922,N_1157);
nor U1898 (N_1898,N_1102,N_153);
or U1899 (N_1899,N_1071,N_983);
xnor U1900 (N_1900,N_1239,N_107);
and U1901 (N_1901,N_851,N_1111);
xnor U1902 (N_1902,N_531,N_1117);
or U1903 (N_1903,N_354,N_480);
and U1904 (N_1904,N_909,N_1098);
xor U1905 (N_1905,N_385,N_415);
or U1906 (N_1906,N_1182,N_1049);
nor U1907 (N_1907,N_892,N_643);
xor U1908 (N_1908,N_86,N_401);
and U1909 (N_1909,N_1155,N_33);
and U1910 (N_1910,N_845,N_1227);
xnor U1911 (N_1911,N_964,N_429);
nand U1912 (N_1912,N_662,N_1104);
xnor U1913 (N_1913,N_1188,N_1100);
and U1914 (N_1914,N_514,N_381);
or U1915 (N_1915,N_1078,N_862);
or U1916 (N_1916,N_338,N_133);
nor U1917 (N_1917,N_241,N_822);
nand U1918 (N_1918,N_282,N_701);
nand U1919 (N_1919,N_1101,N_936);
xnor U1920 (N_1920,N_1035,N_203);
nand U1921 (N_1921,N_835,N_1011);
nor U1922 (N_1922,N_1110,N_802);
nor U1923 (N_1923,N_504,N_398);
nand U1924 (N_1924,N_341,N_256);
xor U1925 (N_1925,N_121,N_428);
xor U1926 (N_1926,N_1179,N_597);
nand U1927 (N_1927,N_634,N_493);
nor U1928 (N_1928,N_870,N_616);
nand U1929 (N_1929,N_246,N_977);
xor U1930 (N_1930,N_0,N_222);
nand U1931 (N_1931,N_20,N_512);
or U1932 (N_1932,N_629,N_710);
nor U1933 (N_1933,N_1178,N_1138);
nand U1934 (N_1934,N_1103,N_1216);
and U1935 (N_1935,N_345,N_34);
nand U1936 (N_1936,N_394,N_336);
xnor U1937 (N_1937,N_289,N_74);
nand U1938 (N_1938,N_199,N_740);
xnor U1939 (N_1939,N_743,N_475);
nand U1940 (N_1940,N_437,N_948);
nor U1941 (N_1941,N_752,N_1052);
nand U1942 (N_1942,N_227,N_756);
nor U1943 (N_1943,N_316,N_65);
or U1944 (N_1944,N_111,N_866);
nor U1945 (N_1945,N_595,N_422);
xor U1946 (N_1946,N_710,N_428);
xnor U1947 (N_1947,N_379,N_695);
nand U1948 (N_1948,N_887,N_1238);
and U1949 (N_1949,N_751,N_158);
nor U1950 (N_1950,N_798,N_154);
or U1951 (N_1951,N_668,N_864);
xor U1952 (N_1952,N_543,N_554);
nor U1953 (N_1953,N_102,N_730);
or U1954 (N_1954,N_196,N_441);
xnor U1955 (N_1955,N_920,N_438);
or U1956 (N_1956,N_67,N_605);
xnor U1957 (N_1957,N_244,N_449);
or U1958 (N_1958,N_55,N_896);
xor U1959 (N_1959,N_889,N_650);
or U1960 (N_1960,N_267,N_13);
nand U1961 (N_1961,N_144,N_37);
or U1962 (N_1962,N_280,N_639);
xnor U1963 (N_1963,N_164,N_741);
xor U1964 (N_1964,N_262,N_815);
nand U1965 (N_1965,N_867,N_158);
or U1966 (N_1966,N_664,N_1201);
nor U1967 (N_1967,N_963,N_1205);
nor U1968 (N_1968,N_1241,N_946);
or U1969 (N_1969,N_67,N_421);
xnor U1970 (N_1970,N_851,N_1001);
or U1971 (N_1971,N_696,N_1029);
xnor U1972 (N_1972,N_364,N_611);
and U1973 (N_1973,N_465,N_980);
or U1974 (N_1974,N_242,N_819);
nand U1975 (N_1975,N_1007,N_364);
nor U1976 (N_1976,N_519,N_1111);
xor U1977 (N_1977,N_849,N_590);
xor U1978 (N_1978,N_456,N_284);
and U1979 (N_1979,N_1219,N_231);
xnor U1980 (N_1980,N_978,N_874);
nand U1981 (N_1981,N_1075,N_709);
and U1982 (N_1982,N_603,N_1237);
nor U1983 (N_1983,N_1231,N_1159);
xor U1984 (N_1984,N_1174,N_718);
and U1985 (N_1985,N_962,N_243);
xnor U1986 (N_1986,N_242,N_143);
or U1987 (N_1987,N_601,N_1015);
or U1988 (N_1988,N_145,N_496);
nand U1989 (N_1989,N_1042,N_8);
xor U1990 (N_1990,N_626,N_810);
nor U1991 (N_1991,N_39,N_293);
nor U1992 (N_1992,N_553,N_811);
xor U1993 (N_1993,N_902,N_92);
and U1994 (N_1994,N_539,N_693);
or U1995 (N_1995,N_518,N_119);
xnor U1996 (N_1996,N_1086,N_1050);
and U1997 (N_1997,N_1108,N_444);
nand U1998 (N_1998,N_1106,N_139);
nor U1999 (N_1999,N_946,N_1062);
nand U2000 (N_2000,N_978,N_778);
nand U2001 (N_2001,N_565,N_607);
or U2002 (N_2002,N_835,N_495);
or U2003 (N_2003,N_120,N_252);
or U2004 (N_2004,N_531,N_172);
and U2005 (N_2005,N_200,N_1102);
xor U2006 (N_2006,N_364,N_619);
xor U2007 (N_2007,N_145,N_974);
nand U2008 (N_2008,N_61,N_934);
xor U2009 (N_2009,N_916,N_1115);
nor U2010 (N_2010,N_1051,N_154);
xor U2011 (N_2011,N_1095,N_1073);
nor U2012 (N_2012,N_318,N_125);
or U2013 (N_2013,N_700,N_579);
nor U2014 (N_2014,N_977,N_289);
xor U2015 (N_2015,N_892,N_1129);
and U2016 (N_2016,N_364,N_250);
nand U2017 (N_2017,N_709,N_881);
nand U2018 (N_2018,N_627,N_293);
or U2019 (N_2019,N_503,N_1235);
xnor U2020 (N_2020,N_48,N_1240);
nor U2021 (N_2021,N_974,N_1077);
or U2022 (N_2022,N_518,N_475);
xnor U2023 (N_2023,N_980,N_343);
and U2024 (N_2024,N_689,N_287);
or U2025 (N_2025,N_517,N_975);
xor U2026 (N_2026,N_888,N_1027);
nor U2027 (N_2027,N_205,N_21);
and U2028 (N_2028,N_465,N_678);
and U2029 (N_2029,N_1011,N_737);
nand U2030 (N_2030,N_915,N_734);
xnor U2031 (N_2031,N_456,N_651);
nand U2032 (N_2032,N_833,N_242);
xnor U2033 (N_2033,N_383,N_480);
nand U2034 (N_2034,N_763,N_279);
or U2035 (N_2035,N_484,N_746);
and U2036 (N_2036,N_420,N_1128);
xor U2037 (N_2037,N_87,N_1167);
nand U2038 (N_2038,N_714,N_448);
and U2039 (N_2039,N_866,N_617);
nor U2040 (N_2040,N_283,N_1155);
xnor U2041 (N_2041,N_962,N_1035);
and U2042 (N_2042,N_1114,N_69);
xor U2043 (N_2043,N_32,N_168);
and U2044 (N_2044,N_1066,N_176);
and U2045 (N_2045,N_293,N_907);
xor U2046 (N_2046,N_757,N_1051);
xnor U2047 (N_2047,N_1227,N_482);
xor U2048 (N_2048,N_711,N_526);
nor U2049 (N_2049,N_38,N_434);
or U2050 (N_2050,N_1214,N_322);
nor U2051 (N_2051,N_949,N_1040);
xnor U2052 (N_2052,N_1153,N_841);
and U2053 (N_2053,N_249,N_772);
and U2054 (N_2054,N_990,N_1005);
or U2055 (N_2055,N_246,N_802);
nand U2056 (N_2056,N_210,N_601);
or U2057 (N_2057,N_1027,N_1090);
nand U2058 (N_2058,N_667,N_521);
nand U2059 (N_2059,N_58,N_1185);
or U2060 (N_2060,N_678,N_206);
or U2061 (N_2061,N_660,N_337);
or U2062 (N_2062,N_1084,N_504);
nor U2063 (N_2063,N_494,N_1019);
or U2064 (N_2064,N_643,N_649);
or U2065 (N_2065,N_326,N_1131);
nor U2066 (N_2066,N_689,N_585);
xor U2067 (N_2067,N_581,N_108);
xnor U2068 (N_2068,N_351,N_1022);
nor U2069 (N_2069,N_1174,N_517);
or U2070 (N_2070,N_1139,N_1127);
or U2071 (N_2071,N_1242,N_613);
or U2072 (N_2072,N_989,N_524);
nor U2073 (N_2073,N_933,N_666);
nand U2074 (N_2074,N_973,N_521);
nor U2075 (N_2075,N_239,N_973);
xnor U2076 (N_2076,N_970,N_1219);
or U2077 (N_2077,N_463,N_779);
nor U2078 (N_2078,N_195,N_795);
nand U2079 (N_2079,N_905,N_133);
xnor U2080 (N_2080,N_1060,N_759);
and U2081 (N_2081,N_257,N_1150);
and U2082 (N_2082,N_1073,N_45);
nand U2083 (N_2083,N_547,N_1100);
nand U2084 (N_2084,N_723,N_642);
nand U2085 (N_2085,N_897,N_898);
nand U2086 (N_2086,N_678,N_1177);
xnor U2087 (N_2087,N_415,N_187);
nand U2088 (N_2088,N_500,N_137);
nor U2089 (N_2089,N_226,N_50);
nand U2090 (N_2090,N_904,N_245);
or U2091 (N_2091,N_160,N_181);
and U2092 (N_2092,N_812,N_379);
xor U2093 (N_2093,N_85,N_475);
xnor U2094 (N_2094,N_654,N_57);
or U2095 (N_2095,N_629,N_58);
nor U2096 (N_2096,N_1103,N_330);
nor U2097 (N_2097,N_787,N_1106);
or U2098 (N_2098,N_649,N_834);
and U2099 (N_2099,N_726,N_678);
or U2100 (N_2100,N_1202,N_1033);
xnor U2101 (N_2101,N_851,N_361);
or U2102 (N_2102,N_262,N_691);
and U2103 (N_2103,N_136,N_591);
nand U2104 (N_2104,N_127,N_25);
nor U2105 (N_2105,N_265,N_255);
nand U2106 (N_2106,N_756,N_760);
nor U2107 (N_2107,N_438,N_523);
xnor U2108 (N_2108,N_446,N_330);
xor U2109 (N_2109,N_1247,N_1136);
nor U2110 (N_2110,N_1201,N_1080);
xnor U2111 (N_2111,N_706,N_1132);
or U2112 (N_2112,N_391,N_989);
or U2113 (N_2113,N_322,N_292);
xnor U2114 (N_2114,N_1202,N_471);
and U2115 (N_2115,N_895,N_1129);
and U2116 (N_2116,N_665,N_926);
xnor U2117 (N_2117,N_421,N_159);
nor U2118 (N_2118,N_247,N_703);
nor U2119 (N_2119,N_672,N_1046);
nor U2120 (N_2120,N_1145,N_615);
xor U2121 (N_2121,N_1043,N_1129);
and U2122 (N_2122,N_1123,N_307);
xnor U2123 (N_2123,N_431,N_872);
nor U2124 (N_2124,N_359,N_212);
and U2125 (N_2125,N_209,N_582);
nand U2126 (N_2126,N_587,N_769);
nor U2127 (N_2127,N_87,N_591);
nor U2128 (N_2128,N_406,N_982);
nand U2129 (N_2129,N_726,N_35);
xnor U2130 (N_2130,N_816,N_946);
nor U2131 (N_2131,N_669,N_535);
nand U2132 (N_2132,N_309,N_254);
or U2133 (N_2133,N_236,N_755);
nor U2134 (N_2134,N_1120,N_1094);
nor U2135 (N_2135,N_34,N_1236);
and U2136 (N_2136,N_169,N_622);
or U2137 (N_2137,N_1217,N_316);
nor U2138 (N_2138,N_15,N_774);
xor U2139 (N_2139,N_504,N_581);
and U2140 (N_2140,N_595,N_332);
nand U2141 (N_2141,N_1163,N_1081);
nand U2142 (N_2142,N_638,N_409);
nand U2143 (N_2143,N_336,N_581);
and U2144 (N_2144,N_38,N_56);
nand U2145 (N_2145,N_664,N_804);
nor U2146 (N_2146,N_657,N_1193);
or U2147 (N_2147,N_327,N_892);
or U2148 (N_2148,N_1106,N_52);
and U2149 (N_2149,N_1152,N_26);
or U2150 (N_2150,N_735,N_587);
and U2151 (N_2151,N_165,N_980);
nand U2152 (N_2152,N_1064,N_14);
nand U2153 (N_2153,N_559,N_1047);
and U2154 (N_2154,N_640,N_1072);
xor U2155 (N_2155,N_901,N_926);
and U2156 (N_2156,N_969,N_777);
nor U2157 (N_2157,N_951,N_614);
and U2158 (N_2158,N_1233,N_1227);
nor U2159 (N_2159,N_531,N_1060);
or U2160 (N_2160,N_815,N_1194);
nor U2161 (N_2161,N_105,N_56);
or U2162 (N_2162,N_889,N_704);
nand U2163 (N_2163,N_488,N_187);
nor U2164 (N_2164,N_128,N_167);
nand U2165 (N_2165,N_1177,N_566);
and U2166 (N_2166,N_1151,N_226);
xnor U2167 (N_2167,N_832,N_29);
and U2168 (N_2168,N_1074,N_871);
and U2169 (N_2169,N_621,N_150);
nand U2170 (N_2170,N_251,N_867);
nor U2171 (N_2171,N_1126,N_1084);
and U2172 (N_2172,N_969,N_1201);
nand U2173 (N_2173,N_291,N_371);
and U2174 (N_2174,N_1013,N_1245);
nor U2175 (N_2175,N_279,N_216);
nand U2176 (N_2176,N_916,N_697);
xor U2177 (N_2177,N_59,N_1033);
and U2178 (N_2178,N_854,N_658);
nand U2179 (N_2179,N_645,N_471);
nor U2180 (N_2180,N_1174,N_280);
nor U2181 (N_2181,N_74,N_616);
and U2182 (N_2182,N_17,N_869);
nand U2183 (N_2183,N_76,N_767);
and U2184 (N_2184,N_48,N_637);
xnor U2185 (N_2185,N_22,N_113);
and U2186 (N_2186,N_1083,N_975);
or U2187 (N_2187,N_214,N_1075);
or U2188 (N_2188,N_986,N_1236);
xnor U2189 (N_2189,N_239,N_281);
nand U2190 (N_2190,N_639,N_680);
and U2191 (N_2191,N_480,N_536);
nand U2192 (N_2192,N_716,N_1011);
xnor U2193 (N_2193,N_86,N_452);
or U2194 (N_2194,N_762,N_1027);
nand U2195 (N_2195,N_1229,N_711);
xor U2196 (N_2196,N_856,N_12);
or U2197 (N_2197,N_267,N_858);
nor U2198 (N_2198,N_255,N_696);
nor U2199 (N_2199,N_201,N_918);
or U2200 (N_2200,N_693,N_189);
and U2201 (N_2201,N_851,N_855);
nor U2202 (N_2202,N_630,N_509);
nand U2203 (N_2203,N_1009,N_52);
nand U2204 (N_2204,N_553,N_785);
xor U2205 (N_2205,N_129,N_154);
nor U2206 (N_2206,N_45,N_1223);
or U2207 (N_2207,N_612,N_857);
xor U2208 (N_2208,N_1226,N_30);
or U2209 (N_2209,N_295,N_504);
xor U2210 (N_2210,N_1035,N_467);
nand U2211 (N_2211,N_250,N_594);
and U2212 (N_2212,N_690,N_687);
nor U2213 (N_2213,N_664,N_635);
or U2214 (N_2214,N_1110,N_28);
nor U2215 (N_2215,N_597,N_134);
xnor U2216 (N_2216,N_480,N_349);
or U2217 (N_2217,N_873,N_724);
nor U2218 (N_2218,N_219,N_430);
nor U2219 (N_2219,N_1055,N_350);
xor U2220 (N_2220,N_240,N_1121);
or U2221 (N_2221,N_466,N_995);
or U2222 (N_2222,N_307,N_514);
or U2223 (N_2223,N_1075,N_1202);
and U2224 (N_2224,N_362,N_782);
nor U2225 (N_2225,N_564,N_1036);
xnor U2226 (N_2226,N_121,N_189);
xnor U2227 (N_2227,N_356,N_377);
and U2228 (N_2228,N_1098,N_1241);
and U2229 (N_2229,N_1008,N_1218);
nor U2230 (N_2230,N_521,N_604);
and U2231 (N_2231,N_494,N_204);
nor U2232 (N_2232,N_432,N_681);
or U2233 (N_2233,N_1104,N_382);
xor U2234 (N_2234,N_683,N_689);
or U2235 (N_2235,N_662,N_1063);
nor U2236 (N_2236,N_564,N_483);
and U2237 (N_2237,N_1148,N_1045);
xor U2238 (N_2238,N_1198,N_562);
or U2239 (N_2239,N_187,N_453);
and U2240 (N_2240,N_981,N_627);
or U2241 (N_2241,N_1052,N_125);
nor U2242 (N_2242,N_386,N_1132);
nor U2243 (N_2243,N_874,N_618);
and U2244 (N_2244,N_1155,N_1118);
nor U2245 (N_2245,N_601,N_12);
and U2246 (N_2246,N_71,N_489);
and U2247 (N_2247,N_196,N_574);
nor U2248 (N_2248,N_114,N_761);
nor U2249 (N_2249,N_61,N_1171);
nor U2250 (N_2250,N_958,N_26);
xnor U2251 (N_2251,N_1189,N_1065);
or U2252 (N_2252,N_355,N_564);
nor U2253 (N_2253,N_176,N_287);
or U2254 (N_2254,N_3,N_1103);
or U2255 (N_2255,N_290,N_695);
and U2256 (N_2256,N_483,N_186);
or U2257 (N_2257,N_754,N_552);
or U2258 (N_2258,N_454,N_628);
or U2259 (N_2259,N_387,N_998);
xnor U2260 (N_2260,N_1069,N_945);
nand U2261 (N_2261,N_1158,N_963);
or U2262 (N_2262,N_1127,N_1075);
nand U2263 (N_2263,N_652,N_103);
or U2264 (N_2264,N_910,N_1037);
nor U2265 (N_2265,N_266,N_193);
nor U2266 (N_2266,N_995,N_691);
and U2267 (N_2267,N_965,N_330);
nand U2268 (N_2268,N_1093,N_144);
and U2269 (N_2269,N_486,N_117);
nand U2270 (N_2270,N_960,N_611);
and U2271 (N_2271,N_381,N_30);
and U2272 (N_2272,N_1022,N_1003);
or U2273 (N_2273,N_516,N_570);
and U2274 (N_2274,N_79,N_760);
nor U2275 (N_2275,N_167,N_557);
and U2276 (N_2276,N_90,N_201);
xor U2277 (N_2277,N_878,N_1077);
nand U2278 (N_2278,N_1106,N_987);
nand U2279 (N_2279,N_218,N_697);
nand U2280 (N_2280,N_811,N_271);
xor U2281 (N_2281,N_1186,N_252);
xnor U2282 (N_2282,N_697,N_191);
and U2283 (N_2283,N_1098,N_56);
xnor U2284 (N_2284,N_1163,N_481);
or U2285 (N_2285,N_739,N_522);
and U2286 (N_2286,N_937,N_929);
xor U2287 (N_2287,N_759,N_561);
or U2288 (N_2288,N_395,N_1198);
nand U2289 (N_2289,N_567,N_1106);
and U2290 (N_2290,N_1060,N_332);
or U2291 (N_2291,N_957,N_711);
nand U2292 (N_2292,N_747,N_403);
nand U2293 (N_2293,N_868,N_738);
or U2294 (N_2294,N_578,N_1134);
nor U2295 (N_2295,N_307,N_1171);
nand U2296 (N_2296,N_626,N_982);
and U2297 (N_2297,N_428,N_133);
nor U2298 (N_2298,N_690,N_946);
and U2299 (N_2299,N_177,N_898);
or U2300 (N_2300,N_496,N_139);
nor U2301 (N_2301,N_653,N_699);
or U2302 (N_2302,N_540,N_809);
and U2303 (N_2303,N_30,N_512);
xor U2304 (N_2304,N_554,N_1183);
and U2305 (N_2305,N_453,N_138);
nor U2306 (N_2306,N_347,N_928);
nor U2307 (N_2307,N_615,N_207);
nor U2308 (N_2308,N_784,N_651);
nand U2309 (N_2309,N_646,N_523);
or U2310 (N_2310,N_405,N_955);
nand U2311 (N_2311,N_695,N_1142);
or U2312 (N_2312,N_132,N_986);
and U2313 (N_2313,N_454,N_937);
or U2314 (N_2314,N_666,N_744);
and U2315 (N_2315,N_443,N_654);
or U2316 (N_2316,N_1017,N_602);
nand U2317 (N_2317,N_867,N_346);
and U2318 (N_2318,N_562,N_905);
or U2319 (N_2319,N_810,N_436);
nand U2320 (N_2320,N_19,N_893);
nand U2321 (N_2321,N_62,N_438);
xor U2322 (N_2322,N_445,N_1228);
and U2323 (N_2323,N_212,N_78);
nor U2324 (N_2324,N_690,N_893);
or U2325 (N_2325,N_688,N_718);
and U2326 (N_2326,N_248,N_451);
nor U2327 (N_2327,N_240,N_908);
or U2328 (N_2328,N_688,N_745);
nand U2329 (N_2329,N_1078,N_1180);
nor U2330 (N_2330,N_1062,N_742);
nor U2331 (N_2331,N_437,N_751);
or U2332 (N_2332,N_415,N_12);
xnor U2333 (N_2333,N_605,N_235);
or U2334 (N_2334,N_827,N_883);
or U2335 (N_2335,N_788,N_281);
and U2336 (N_2336,N_5,N_279);
or U2337 (N_2337,N_522,N_1135);
nor U2338 (N_2338,N_522,N_537);
and U2339 (N_2339,N_27,N_1003);
nor U2340 (N_2340,N_157,N_215);
or U2341 (N_2341,N_413,N_782);
and U2342 (N_2342,N_608,N_914);
and U2343 (N_2343,N_796,N_712);
xnor U2344 (N_2344,N_955,N_990);
nor U2345 (N_2345,N_688,N_748);
nor U2346 (N_2346,N_161,N_833);
nand U2347 (N_2347,N_1044,N_40);
or U2348 (N_2348,N_276,N_241);
or U2349 (N_2349,N_520,N_398);
or U2350 (N_2350,N_1058,N_424);
nand U2351 (N_2351,N_813,N_73);
and U2352 (N_2352,N_586,N_166);
and U2353 (N_2353,N_1098,N_57);
nor U2354 (N_2354,N_930,N_831);
nand U2355 (N_2355,N_741,N_67);
nor U2356 (N_2356,N_324,N_1120);
or U2357 (N_2357,N_1215,N_296);
nor U2358 (N_2358,N_111,N_1035);
nand U2359 (N_2359,N_337,N_842);
nand U2360 (N_2360,N_943,N_681);
or U2361 (N_2361,N_850,N_944);
nand U2362 (N_2362,N_383,N_1106);
and U2363 (N_2363,N_1032,N_249);
or U2364 (N_2364,N_235,N_419);
xor U2365 (N_2365,N_747,N_399);
and U2366 (N_2366,N_1000,N_521);
xnor U2367 (N_2367,N_119,N_573);
and U2368 (N_2368,N_10,N_304);
nand U2369 (N_2369,N_103,N_401);
and U2370 (N_2370,N_304,N_1006);
nor U2371 (N_2371,N_701,N_264);
or U2372 (N_2372,N_378,N_199);
xor U2373 (N_2373,N_580,N_388);
nand U2374 (N_2374,N_1243,N_639);
or U2375 (N_2375,N_674,N_1163);
xor U2376 (N_2376,N_939,N_825);
and U2377 (N_2377,N_910,N_1057);
nand U2378 (N_2378,N_893,N_110);
nand U2379 (N_2379,N_235,N_189);
nand U2380 (N_2380,N_385,N_130);
and U2381 (N_2381,N_1087,N_368);
and U2382 (N_2382,N_1042,N_512);
and U2383 (N_2383,N_1222,N_979);
nor U2384 (N_2384,N_561,N_1239);
xnor U2385 (N_2385,N_1089,N_371);
nand U2386 (N_2386,N_1233,N_40);
nand U2387 (N_2387,N_795,N_1113);
nand U2388 (N_2388,N_1059,N_1016);
nand U2389 (N_2389,N_785,N_1078);
or U2390 (N_2390,N_269,N_89);
xnor U2391 (N_2391,N_18,N_1034);
and U2392 (N_2392,N_608,N_105);
nor U2393 (N_2393,N_1138,N_771);
nor U2394 (N_2394,N_783,N_827);
nand U2395 (N_2395,N_369,N_918);
nand U2396 (N_2396,N_5,N_685);
and U2397 (N_2397,N_615,N_417);
or U2398 (N_2398,N_362,N_383);
or U2399 (N_2399,N_141,N_999);
and U2400 (N_2400,N_1021,N_855);
and U2401 (N_2401,N_552,N_1098);
xnor U2402 (N_2402,N_853,N_1249);
or U2403 (N_2403,N_839,N_298);
nand U2404 (N_2404,N_934,N_828);
and U2405 (N_2405,N_1060,N_835);
nor U2406 (N_2406,N_277,N_753);
and U2407 (N_2407,N_1161,N_132);
and U2408 (N_2408,N_492,N_853);
or U2409 (N_2409,N_642,N_558);
and U2410 (N_2410,N_587,N_1243);
or U2411 (N_2411,N_380,N_474);
or U2412 (N_2412,N_1124,N_65);
or U2413 (N_2413,N_1118,N_659);
nor U2414 (N_2414,N_1210,N_279);
nor U2415 (N_2415,N_182,N_1197);
nor U2416 (N_2416,N_563,N_1205);
nand U2417 (N_2417,N_354,N_279);
and U2418 (N_2418,N_1034,N_1116);
or U2419 (N_2419,N_354,N_790);
xnor U2420 (N_2420,N_327,N_149);
nand U2421 (N_2421,N_756,N_44);
and U2422 (N_2422,N_88,N_97);
nor U2423 (N_2423,N_885,N_896);
nand U2424 (N_2424,N_448,N_1177);
nand U2425 (N_2425,N_1199,N_856);
nor U2426 (N_2426,N_384,N_910);
nor U2427 (N_2427,N_745,N_601);
nand U2428 (N_2428,N_401,N_381);
nand U2429 (N_2429,N_95,N_29);
nand U2430 (N_2430,N_396,N_1035);
and U2431 (N_2431,N_408,N_609);
and U2432 (N_2432,N_408,N_694);
nand U2433 (N_2433,N_181,N_852);
nor U2434 (N_2434,N_894,N_838);
nor U2435 (N_2435,N_186,N_344);
or U2436 (N_2436,N_1202,N_633);
xor U2437 (N_2437,N_449,N_308);
nand U2438 (N_2438,N_74,N_405);
xor U2439 (N_2439,N_550,N_68);
or U2440 (N_2440,N_264,N_289);
or U2441 (N_2441,N_871,N_682);
nor U2442 (N_2442,N_193,N_60);
nor U2443 (N_2443,N_1197,N_453);
xnor U2444 (N_2444,N_179,N_22);
and U2445 (N_2445,N_281,N_887);
or U2446 (N_2446,N_896,N_219);
nand U2447 (N_2447,N_804,N_769);
nor U2448 (N_2448,N_982,N_68);
nand U2449 (N_2449,N_1,N_847);
and U2450 (N_2450,N_144,N_920);
or U2451 (N_2451,N_944,N_1042);
and U2452 (N_2452,N_240,N_43);
nor U2453 (N_2453,N_1125,N_281);
nor U2454 (N_2454,N_740,N_687);
nor U2455 (N_2455,N_1131,N_638);
and U2456 (N_2456,N_1092,N_896);
and U2457 (N_2457,N_1142,N_442);
nor U2458 (N_2458,N_349,N_720);
nor U2459 (N_2459,N_92,N_222);
and U2460 (N_2460,N_932,N_898);
nand U2461 (N_2461,N_290,N_515);
or U2462 (N_2462,N_1042,N_855);
nor U2463 (N_2463,N_449,N_1095);
or U2464 (N_2464,N_980,N_672);
and U2465 (N_2465,N_1185,N_81);
and U2466 (N_2466,N_311,N_998);
nand U2467 (N_2467,N_789,N_104);
nor U2468 (N_2468,N_556,N_18);
nand U2469 (N_2469,N_324,N_345);
nand U2470 (N_2470,N_391,N_828);
xor U2471 (N_2471,N_596,N_179);
or U2472 (N_2472,N_321,N_281);
and U2473 (N_2473,N_295,N_1162);
and U2474 (N_2474,N_714,N_328);
nand U2475 (N_2475,N_744,N_192);
and U2476 (N_2476,N_964,N_526);
or U2477 (N_2477,N_185,N_1231);
xor U2478 (N_2478,N_588,N_37);
or U2479 (N_2479,N_233,N_324);
nand U2480 (N_2480,N_70,N_585);
or U2481 (N_2481,N_226,N_7);
nand U2482 (N_2482,N_439,N_888);
xor U2483 (N_2483,N_216,N_371);
nand U2484 (N_2484,N_1081,N_880);
xnor U2485 (N_2485,N_345,N_1025);
nand U2486 (N_2486,N_380,N_993);
nand U2487 (N_2487,N_404,N_442);
nand U2488 (N_2488,N_235,N_351);
nand U2489 (N_2489,N_837,N_1034);
and U2490 (N_2490,N_1084,N_261);
nand U2491 (N_2491,N_634,N_192);
nor U2492 (N_2492,N_569,N_1118);
nor U2493 (N_2493,N_321,N_169);
xnor U2494 (N_2494,N_930,N_1081);
nand U2495 (N_2495,N_906,N_261);
nand U2496 (N_2496,N_857,N_1166);
nand U2497 (N_2497,N_717,N_601);
nor U2498 (N_2498,N_940,N_605);
nand U2499 (N_2499,N_401,N_4);
or U2500 (N_2500,N_1425,N_1912);
xor U2501 (N_2501,N_2120,N_2330);
and U2502 (N_2502,N_1937,N_1686);
and U2503 (N_2503,N_2492,N_2478);
xnor U2504 (N_2504,N_1824,N_1782);
nor U2505 (N_2505,N_1322,N_1476);
xor U2506 (N_2506,N_1525,N_1406);
and U2507 (N_2507,N_2374,N_1295);
and U2508 (N_2508,N_1332,N_1873);
nand U2509 (N_2509,N_1694,N_2017);
or U2510 (N_2510,N_1356,N_1656);
nor U2511 (N_2511,N_2367,N_1405);
or U2512 (N_2512,N_2240,N_2339);
or U2513 (N_2513,N_1521,N_1427);
nor U2514 (N_2514,N_1254,N_1276);
or U2515 (N_2515,N_1924,N_2485);
nand U2516 (N_2516,N_2475,N_2405);
xnor U2517 (N_2517,N_2165,N_1450);
or U2518 (N_2518,N_1714,N_1261);
xnor U2519 (N_2519,N_1371,N_1960);
or U2520 (N_2520,N_1372,N_1556);
xor U2521 (N_2521,N_1250,N_2122);
nor U2522 (N_2522,N_1483,N_2451);
nor U2523 (N_2523,N_2351,N_2385);
xnor U2524 (N_2524,N_2156,N_1411);
xnor U2525 (N_2525,N_2369,N_2084);
or U2526 (N_2526,N_1601,N_1514);
nor U2527 (N_2527,N_2461,N_2457);
and U2528 (N_2528,N_1424,N_2293);
nor U2529 (N_2529,N_2104,N_2440);
nor U2530 (N_2530,N_1401,N_1396);
and U2531 (N_2531,N_1610,N_2024);
xor U2532 (N_2532,N_1773,N_2463);
or U2533 (N_2533,N_2153,N_2264);
or U2534 (N_2534,N_2020,N_1669);
nor U2535 (N_2535,N_1699,N_1571);
nand U2536 (N_2536,N_1710,N_1992);
nand U2537 (N_2537,N_1465,N_1837);
nor U2538 (N_2538,N_1379,N_2487);
nand U2539 (N_2539,N_1552,N_1280);
xnor U2540 (N_2540,N_2035,N_2037);
nor U2541 (N_2541,N_2412,N_1900);
xnor U2542 (N_2542,N_1795,N_1765);
nand U2543 (N_2543,N_2381,N_2032);
nand U2544 (N_2544,N_2126,N_2443);
nand U2545 (N_2545,N_2252,N_2195);
nand U2546 (N_2546,N_2277,N_1857);
xor U2547 (N_2547,N_1586,N_1800);
nor U2548 (N_2548,N_2242,N_2263);
nor U2549 (N_2549,N_1292,N_2229);
nor U2550 (N_2550,N_2395,N_2481);
and U2551 (N_2551,N_1255,N_1839);
xnor U2552 (N_2552,N_2436,N_1670);
and U2553 (N_2553,N_2409,N_2149);
nor U2554 (N_2554,N_1343,N_1813);
or U2555 (N_2555,N_1784,N_1358);
xor U2556 (N_2556,N_2491,N_1646);
or U2557 (N_2557,N_1880,N_2125);
nand U2558 (N_2558,N_1385,N_1709);
nand U2559 (N_2559,N_1618,N_1602);
nor U2560 (N_2560,N_2352,N_2167);
and U2561 (N_2561,N_1897,N_1660);
xnor U2562 (N_2562,N_2151,N_1352);
and U2563 (N_2563,N_2201,N_1456);
and U2564 (N_2564,N_1755,N_1503);
and U2565 (N_2565,N_1805,N_1944);
xor U2566 (N_2566,N_2427,N_2011);
xor U2567 (N_2567,N_2426,N_1978);
nand U2568 (N_2568,N_1827,N_2190);
or U2569 (N_2569,N_1868,N_1852);
or U2570 (N_2570,N_2180,N_1417);
nand U2571 (N_2571,N_2086,N_2102);
xnor U2572 (N_2572,N_1674,N_2424);
or U2573 (N_2573,N_2007,N_1965);
nor U2574 (N_2574,N_1941,N_1722);
or U2575 (N_2575,N_1706,N_1653);
nor U2576 (N_2576,N_1329,N_1690);
nand U2577 (N_2577,N_1902,N_1467);
and U2578 (N_2578,N_1655,N_1613);
nor U2579 (N_2579,N_1855,N_1432);
nor U2580 (N_2580,N_1957,N_2444);
and U2581 (N_2581,N_2021,N_1468);
and U2582 (N_2582,N_1550,N_1374);
xnor U2583 (N_2583,N_1695,N_2009);
nor U2584 (N_2584,N_2121,N_1463);
nor U2585 (N_2585,N_2209,N_1859);
or U2586 (N_2586,N_2309,N_2090);
and U2587 (N_2587,N_2110,N_1736);
xor U2588 (N_2588,N_2148,N_2453);
xnor U2589 (N_2589,N_2313,N_2189);
or U2590 (N_2590,N_1812,N_2442);
and U2591 (N_2591,N_1335,N_2285);
or U2592 (N_2592,N_1604,N_2188);
nand U2593 (N_2593,N_1953,N_1664);
nor U2594 (N_2594,N_1445,N_1866);
xor U2595 (N_2595,N_2213,N_1461);
xnor U2596 (N_2596,N_2464,N_1717);
or U2597 (N_2597,N_2327,N_1841);
nand U2598 (N_2598,N_1407,N_1293);
xor U2599 (N_2599,N_1557,N_2376);
and U2600 (N_2600,N_2113,N_1661);
nor U2601 (N_2601,N_1310,N_1872);
xnor U2602 (N_2602,N_2298,N_1530);
or U2603 (N_2603,N_1451,N_2222);
or U2604 (N_2604,N_1938,N_1564);
nor U2605 (N_2605,N_1973,N_2085);
nor U2606 (N_2606,N_2158,N_1495);
nor U2607 (N_2607,N_1883,N_1911);
nand U2608 (N_2608,N_2407,N_1497);
and U2609 (N_2609,N_2228,N_2000);
xnor U2610 (N_2610,N_1752,N_1728);
and U2611 (N_2611,N_2254,N_1475);
nor U2612 (N_2612,N_1631,N_1625);
xnor U2613 (N_2613,N_2283,N_2386);
nand U2614 (N_2614,N_1575,N_2490);
nor U2615 (N_2615,N_2134,N_2029);
xor U2616 (N_2616,N_2109,N_2185);
xnor U2617 (N_2617,N_1548,N_1893);
nor U2618 (N_2618,N_2067,N_1865);
or U2619 (N_2619,N_2399,N_1500);
xor U2620 (N_2620,N_1394,N_2471);
and U2621 (N_2621,N_1366,N_2250);
xnor U2622 (N_2622,N_2336,N_2215);
nor U2623 (N_2623,N_1850,N_1914);
nor U2624 (N_2624,N_1623,N_1913);
nor U2625 (N_2625,N_1763,N_1729);
xor U2626 (N_2626,N_1315,N_2181);
nor U2627 (N_2627,N_2211,N_1415);
xnor U2628 (N_2628,N_2187,N_1616);
nor U2629 (N_2629,N_2382,N_1704);
nor U2630 (N_2630,N_1266,N_2324);
and U2631 (N_2631,N_2350,N_2059);
nor U2632 (N_2632,N_1447,N_1681);
and U2633 (N_2633,N_2160,N_1511);
xor U2634 (N_2634,N_2275,N_1317);
xor U2635 (N_2635,N_2145,N_2207);
nor U2636 (N_2636,N_1718,N_2301);
nand U2637 (N_2637,N_2019,N_1365);
and U2638 (N_2638,N_1864,N_2220);
and U2639 (N_2639,N_1874,N_1934);
nor U2640 (N_2640,N_1970,N_1323);
nand U2641 (N_2641,N_1448,N_1504);
or U2642 (N_2642,N_1481,N_1454);
xnor U2643 (N_2643,N_1338,N_1684);
and U2644 (N_2644,N_1825,N_1667);
nor U2645 (N_2645,N_2249,N_2458);
nor U2646 (N_2646,N_1522,N_1311);
xnor U2647 (N_2647,N_1357,N_1251);
xor U2648 (N_2648,N_1819,N_1856);
or U2649 (N_2649,N_1766,N_1532);
nor U2650 (N_2650,N_1940,N_1932);
nor U2651 (N_2651,N_1961,N_1489);
and U2652 (N_2652,N_2287,N_2439);
nand U2653 (N_2653,N_2403,N_2413);
xor U2654 (N_2654,N_1470,N_2251);
and U2655 (N_2655,N_1484,N_1834);
xnor U2656 (N_2656,N_1526,N_1933);
or U2657 (N_2657,N_2075,N_1288);
and U2658 (N_2658,N_1414,N_1318);
xor U2659 (N_2659,N_2018,N_1304);
nor U2660 (N_2660,N_1869,N_1927);
or U2661 (N_2661,N_1378,N_1362);
or U2662 (N_2662,N_2077,N_2438);
and U2663 (N_2663,N_1615,N_1359);
nor U2664 (N_2664,N_2166,N_2141);
nand U2665 (N_2665,N_1917,N_1705);
nand U2666 (N_2666,N_2106,N_1691);
and U2667 (N_2667,N_2095,N_2206);
or U2668 (N_2668,N_2172,N_1528);
nand U2669 (N_2669,N_2042,N_1723);
nand U2670 (N_2670,N_1386,N_1307);
nor U2671 (N_2671,N_1399,N_1324);
and U2672 (N_2672,N_1529,N_1888);
or U2673 (N_2673,N_1891,N_1585);
nor U2674 (N_2674,N_1693,N_1984);
or U2675 (N_2675,N_2061,N_1887);
nor U2676 (N_2676,N_1547,N_2316);
nor U2677 (N_2677,N_1517,N_1840);
xnor U2678 (N_2678,N_1423,N_2329);
nor U2679 (N_2679,N_1466,N_2100);
nand U2680 (N_2680,N_1297,N_2380);
nand U2681 (N_2681,N_1527,N_2318);
and U2682 (N_2682,N_2299,N_2331);
or U2683 (N_2683,N_1596,N_1999);
nand U2684 (N_2684,N_1789,N_2080);
and U2685 (N_2685,N_2346,N_1397);
and U2686 (N_2686,N_1867,N_2312);
xnor U2687 (N_2687,N_1491,N_2473);
and U2688 (N_2688,N_2493,N_2105);
and U2689 (N_2689,N_1457,N_2051);
nand U2690 (N_2690,N_1654,N_2448);
or U2691 (N_2691,N_1682,N_1726);
nand U2692 (N_2692,N_1898,N_1672);
nand U2693 (N_2693,N_1538,N_2495);
nor U2694 (N_2694,N_2014,N_2484);
and U2695 (N_2695,N_1929,N_1997);
and U2696 (N_2696,N_1761,N_1267);
or U2697 (N_2697,N_1790,N_2334);
or U2698 (N_2698,N_1712,N_1344);
and U2699 (N_2699,N_2154,N_1985);
and U2700 (N_2700,N_2361,N_1620);
or U2701 (N_2701,N_2226,N_2304);
and U2702 (N_2702,N_1435,N_1702);
nand U2703 (N_2703,N_1786,N_1942);
xor U2704 (N_2704,N_1871,N_2421);
nor U2705 (N_2705,N_1460,N_1707);
nand U2706 (N_2706,N_2199,N_1638);
nand U2707 (N_2707,N_2420,N_2150);
nand U2708 (N_2708,N_1634,N_2069);
nand U2709 (N_2709,N_2223,N_2186);
xor U2710 (N_2710,N_2040,N_2237);
nor U2711 (N_2711,N_2072,N_2370);
nor U2712 (N_2712,N_2398,N_2219);
nand U2713 (N_2713,N_2163,N_1594);
nand U2714 (N_2714,N_1862,N_1587);
xnor U2715 (N_2715,N_1746,N_2270);
and U2716 (N_2716,N_1713,N_1534);
nand U2717 (N_2717,N_1403,N_1779);
nand U2718 (N_2718,N_1796,N_2099);
nor U2719 (N_2719,N_2146,N_1648);
xor U2720 (N_2720,N_2498,N_2118);
nor U2721 (N_2721,N_1811,N_1611);
nand U2722 (N_2722,N_1993,N_1762);
xnor U2723 (N_2723,N_1303,N_2015);
xnor U2724 (N_2724,N_1679,N_2179);
nand U2725 (N_2725,N_1949,N_2247);
nor U2726 (N_2726,N_2288,N_2294);
xor U2727 (N_2727,N_1890,N_1482);
xnor U2728 (N_2728,N_1903,N_1732);
or U2729 (N_2729,N_1909,N_1991);
nand U2730 (N_2730,N_1260,N_2048);
or U2731 (N_2731,N_1389,N_2348);
nand U2732 (N_2732,N_2400,N_1472);
xnor U2733 (N_2733,N_1597,N_2266);
nor U2734 (N_2734,N_2447,N_2333);
or U2735 (N_2735,N_2202,N_1607);
nand U2736 (N_2736,N_2307,N_1633);
or U2737 (N_2737,N_1591,N_2469);
or U2738 (N_2738,N_2300,N_2483);
xor U2739 (N_2739,N_2353,N_1284);
xnor U2740 (N_2740,N_1543,N_1275);
xor U2741 (N_2741,N_1436,N_2114);
nand U2742 (N_2742,N_2383,N_1851);
and U2743 (N_2743,N_1719,N_1730);
or U2744 (N_2744,N_1747,N_1636);
xnor U2745 (N_2745,N_1383,N_1849);
and U2746 (N_2746,N_1540,N_2480);
nand U2747 (N_2747,N_1418,N_1531);
nor U2748 (N_2748,N_2183,N_1420);
and U2749 (N_2749,N_2107,N_1382);
and U2750 (N_2750,N_1926,N_2210);
nor U2751 (N_2751,N_2272,N_1626);
or U2752 (N_2752,N_1832,N_1496);
or U2753 (N_2753,N_1257,N_1823);
nand U2754 (N_2754,N_1627,N_1433);
nand U2755 (N_2755,N_1506,N_1434);
nor U2756 (N_2756,N_2235,N_1369);
and U2757 (N_2757,N_1922,N_2450);
or U2758 (N_2758,N_1889,N_2081);
or U2759 (N_2759,N_2452,N_1885);
and U2760 (N_2760,N_1325,N_1769);
nand U2761 (N_2761,N_1649,N_1774);
nor U2762 (N_2762,N_2174,N_2005);
or U2763 (N_2763,N_2119,N_1683);
xnor U2764 (N_2764,N_2083,N_1508);
xor U2765 (N_2765,N_2355,N_1921);
nand U2766 (N_2766,N_1925,N_2049);
nor U2767 (N_2767,N_1809,N_1858);
nor U2768 (N_2768,N_1493,N_2401);
nand U2769 (N_2769,N_2050,N_1593);
nand U2770 (N_2770,N_1665,N_1515);
and U2771 (N_2771,N_1539,N_2359);
xnor U2772 (N_2772,N_2038,N_1826);
nor U2773 (N_2773,N_2143,N_2257);
or U2774 (N_2774,N_2238,N_2064);
and U2775 (N_2775,N_1798,N_1689);
nand U2776 (N_2776,N_1563,N_1523);
and U2777 (N_2777,N_1551,N_2397);
or U2778 (N_2778,N_2454,N_2227);
nor U2779 (N_2779,N_1904,N_2411);
and U2780 (N_2780,N_2248,N_1252);
or U2781 (N_2781,N_2253,N_1737);
xnor U2782 (N_2782,N_1599,N_2071);
xnor U2783 (N_2783,N_2045,N_1640);
and U2784 (N_2784,N_1595,N_2030);
and U2785 (N_2785,N_1760,N_1348);
and U2786 (N_2786,N_2496,N_1884);
and U2787 (N_2787,N_1939,N_2203);
or U2788 (N_2788,N_1817,N_2332);
or U2789 (N_2789,N_1298,N_1963);
nand U2790 (N_2790,N_2244,N_1580);
or U2791 (N_2791,N_1629,N_1738);
nand U2792 (N_2792,N_2488,N_1845);
nand U2793 (N_2793,N_2322,N_1996);
nor U2794 (N_2794,N_1314,N_1637);
xor U2795 (N_2795,N_1576,N_2391);
and U2796 (N_2796,N_1778,N_1316);
nand U2797 (N_2797,N_1271,N_1931);
xnor U2798 (N_2798,N_1642,N_2023);
and U2799 (N_2799,N_2423,N_2265);
nand U2800 (N_2800,N_1802,N_1346);
or U2801 (N_2801,N_1969,N_2320);
nor U2802 (N_2802,N_1810,N_2344);
nand U2803 (N_2803,N_2378,N_1986);
and U2804 (N_2804,N_1264,N_2041);
nand U2805 (N_2805,N_1347,N_1886);
nand U2806 (N_2806,N_1748,N_2422);
or U2807 (N_2807,N_1830,N_2096);
xnor U2808 (N_2808,N_2073,N_2338);
and U2809 (N_2809,N_2261,N_1480);
nand U2810 (N_2810,N_1395,N_1512);
nor U2811 (N_2811,N_2255,N_1408);
or U2812 (N_2812,N_1505,N_2245);
xnor U2813 (N_2813,N_1390,N_1305);
nand U2814 (N_2814,N_2001,N_2328);
or U2815 (N_2815,N_1609,N_2124);
nor U2816 (N_2816,N_2295,N_2305);
nor U2817 (N_2817,N_2175,N_2177);
nor U2818 (N_2818,N_2441,N_1741);
nor U2819 (N_2819,N_2394,N_1647);
xnor U2820 (N_2820,N_2162,N_1946);
nor U2821 (N_2821,N_1474,N_2410);
nor U2822 (N_2822,N_1906,N_1750);
nor U2823 (N_2823,N_2058,N_1846);
nor U2824 (N_2824,N_1838,N_2357);
nand U2825 (N_2825,N_1377,N_2142);
and U2826 (N_2826,N_2326,N_2256);
xor U2827 (N_2827,N_2470,N_1589);
and U2828 (N_2828,N_1757,N_2499);
or U2829 (N_2829,N_2340,N_1402);
xnor U2830 (N_2830,N_1645,N_1605);
and U2831 (N_2831,N_1287,N_2170);
or U2832 (N_2832,N_1614,N_2204);
nand U2833 (N_2833,N_1549,N_1622);
or U2834 (N_2834,N_1892,N_2306);
nand U2835 (N_2835,N_1494,N_1606);
and U2836 (N_2836,N_2432,N_1847);
nand U2837 (N_2837,N_1799,N_2362);
xnor U2838 (N_2838,N_1662,N_1392);
nand U2839 (N_2839,N_2392,N_2097);
nand U2840 (N_2840,N_1536,N_2390);
xor U2841 (N_2841,N_2366,N_1915);
nand U2842 (N_2842,N_1772,N_1899);
nand U2843 (N_2843,N_1680,N_1313);
xnor U2844 (N_2844,N_1928,N_2089);
and U2845 (N_2845,N_2388,N_2416);
nor U2846 (N_2846,N_2200,N_1974);
or U2847 (N_2847,N_2321,N_1381);
nand U2848 (N_2848,N_1703,N_1603);
xnor U2849 (N_2849,N_2093,N_1833);
and U2850 (N_2850,N_1326,N_1485);
xor U2851 (N_2851,N_2062,N_1398);
and U2852 (N_2852,N_1650,N_2356);
xor U2853 (N_2853,N_1980,N_1624);
and U2854 (N_2854,N_1598,N_1330);
and U2855 (N_2855,N_2088,N_1351);
xor U2856 (N_2856,N_1520,N_1334);
nand U2857 (N_2857,N_1768,N_1464);
nand U2858 (N_2858,N_1780,N_1881);
nand U2859 (N_2859,N_1895,N_2196);
xnor U2860 (N_2860,N_2214,N_1806);
nand U2861 (N_2861,N_2433,N_1574);
and U2862 (N_2862,N_1278,N_2449);
nor U2863 (N_2863,N_2198,N_1458);
or U2864 (N_2864,N_1477,N_1579);
xnor U2865 (N_2865,N_1966,N_2466);
nor U2866 (N_2866,N_1367,N_1982);
or U2867 (N_2867,N_1989,N_1977);
nor U2868 (N_2868,N_2043,N_1758);
nand U2869 (N_2869,N_1578,N_2291);
or U2870 (N_2870,N_2002,N_1312);
or U2871 (N_2871,N_2087,N_1544);
nor U2872 (N_2872,N_1630,N_1339);
nand U2873 (N_2873,N_2415,N_1518);
or U2874 (N_2874,N_2360,N_1373);
and U2875 (N_2875,N_1308,N_1764);
nor U2876 (N_2876,N_1950,N_1328);
xnor U2877 (N_2877,N_1877,N_2130);
xnor U2878 (N_2878,N_1258,N_1854);
xor U2879 (N_2879,N_2091,N_1785);
or U2880 (N_2880,N_2078,N_2232);
or U2881 (N_2881,N_1767,N_1286);
nand U2882 (N_2882,N_1791,N_1588);
or U2883 (N_2883,N_2292,N_1268);
xnor U2884 (N_2884,N_2414,N_2065);
xor U2885 (N_2885,N_2406,N_2396);
nand U2886 (N_2886,N_1787,N_1289);
nand U2887 (N_2887,N_1701,N_2046);
xor U2888 (N_2888,N_2135,N_1443);
nand U2889 (N_2889,N_1582,N_2060);
xor U2890 (N_2890,N_2341,N_1509);
nand U2891 (N_2891,N_1519,N_2280);
or U2892 (N_2892,N_1513,N_2092);
nand U2893 (N_2893,N_1368,N_1901);
and U2894 (N_2894,N_1972,N_1797);
and U2895 (N_2895,N_2218,N_2236);
and U2896 (N_2896,N_2445,N_2116);
or U2897 (N_2897,N_2074,N_1777);
or U2898 (N_2898,N_2025,N_2027);
nand U2899 (N_2899,N_1641,N_2476);
or U2900 (N_2900,N_2314,N_2468);
or U2901 (N_2901,N_2022,N_2205);
xor U2902 (N_2902,N_1537,N_1444);
nor U2903 (N_2903,N_1816,N_1673);
and U2904 (N_2904,N_1498,N_2258);
xnor U2905 (N_2905,N_1400,N_1676);
xor U2906 (N_2906,N_1253,N_2171);
xnor U2907 (N_2907,N_1487,N_1793);
and U2908 (N_2908,N_2013,N_1727);
xor U2909 (N_2909,N_2197,N_1583);
nand U2910 (N_2910,N_1380,N_2034);
or U2911 (N_2911,N_1376,N_1700);
or U2912 (N_2912,N_2243,N_2082);
and U2913 (N_2913,N_2267,N_1745);
nand U2914 (N_2914,N_1370,N_1685);
or U2915 (N_2915,N_1724,N_1987);
or U2916 (N_2916,N_1256,N_2363);
xnor U2917 (N_2917,N_2225,N_1663);
xor U2918 (N_2918,N_2335,N_1262);
and U2919 (N_2919,N_1644,N_2435);
nand U2920 (N_2920,N_1945,N_1671);
nor U2921 (N_2921,N_2066,N_1783);
nor U2922 (N_2922,N_1716,N_1259);
or U2923 (N_2923,N_1959,N_2036);
or U2924 (N_2924,N_2325,N_1687);
xnor U2925 (N_2925,N_1958,N_1501);
or U2926 (N_2926,N_1265,N_2127);
or U2927 (N_2927,N_2479,N_1413);
nand U2928 (N_2928,N_2393,N_1441);
or U2929 (N_2929,N_2434,N_1320);
nand U2930 (N_2930,N_1964,N_2289);
nor U2931 (N_2931,N_2349,N_1421);
nor U2932 (N_2932,N_1341,N_1905);
nand U2933 (N_2933,N_2233,N_2234);
nand U2934 (N_2934,N_2379,N_1568);
nor U2935 (N_2935,N_2271,N_2133);
nand U2936 (N_2936,N_1462,N_1831);
or U2937 (N_2937,N_2460,N_1801);
or U2938 (N_2938,N_1279,N_1416);
or U2939 (N_2939,N_1870,N_2076);
nand U2940 (N_2940,N_2428,N_1302);
or U2941 (N_2941,N_1734,N_1566);
or U2942 (N_2942,N_2437,N_1876);
or U2943 (N_2943,N_1263,N_2310);
nand U2944 (N_2944,N_2159,N_1651);
nand U2945 (N_2945,N_2169,N_1269);
nand U2946 (N_2946,N_1469,N_1930);
nor U2947 (N_2947,N_1751,N_1422);
or U2948 (N_2948,N_2303,N_2052);
or U2949 (N_2949,N_2039,N_1842);
or U2950 (N_2950,N_2164,N_1455);
and U2951 (N_2951,N_1510,N_1569);
xnor U2952 (N_2952,N_2375,N_2274);
and U2953 (N_2953,N_1558,N_1355);
and U2954 (N_2954,N_1409,N_2108);
or U2955 (N_2955,N_1488,N_1619);
and U2956 (N_2956,N_2006,N_2230);
and U2957 (N_2957,N_1449,N_1731);
and U2958 (N_2958,N_1742,N_1822);
and U2959 (N_2959,N_1577,N_2026);
and U2960 (N_2960,N_1643,N_1565);
xor U2961 (N_2961,N_1971,N_2279);
and U2962 (N_2962,N_1273,N_1918);
nor U2963 (N_2963,N_2315,N_2284);
nand U2964 (N_2964,N_1688,N_2178);
and U2965 (N_2965,N_2486,N_2455);
nor U2966 (N_2966,N_2094,N_1894);
nand U2967 (N_2967,N_2033,N_2070);
nor U2968 (N_2968,N_1657,N_1471);
xnor U2969 (N_2969,N_2446,N_1749);
nand U2970 (N_2970,N_1967,N_1919);
nor U2971 (N_2971,N_1440,N_2389);
nand U2972 (N_2972,N_1535,N_1882);
or U2973 (N_2973,N_2139,N_1490);
nor U2974 (N_2974,N_1916,N_2137);
nor U2975 (N_2975,N_1896,N_1754);
or U2976 (N_2976,N_2372,N_1981);
and U2977 (N_2977,N_1479,N_1430);
nor U2978 (N_2978,N_1561,N_1794);
nor U2979 (N_2979,N_2068,N_1560);
and U2980 (N_2980,N_1920,N_1473);
and U2981 (N_2981,N_1282,N_2129);
nand U2982 (N_2982,N_1621,N_2281);
nor U2983 (N_2983,N_1478,N_1309);
or U2984 (N_2984,N_2117,N_2155);
nand U2985 (N_2985,N_1948,N_1725);
or U2986 (N_2986,N_2152,N_1628);
nor U2987 (N_2987,N_2138,N_1781);
xnor U2988 (N_2988,N_1590,N_2173);
xnor U2989 (N_2989,N_2157,N_2302);
nor U2990 (N_2990,N_2028,N_2269);
nand U2991 (N_2991,N_2132,N_1361);
xnor U2992 (N_2992,N_2364,N_1951);
or U2993 (N_2993,N_2342,N_1771);
or U2994 (N_2994,N_1828,N_1814);
or U2995 (N_2995,N_1281,N_1776);
or U2996 (N_2996,N_1438,N_2246);
nor U2997 (N_2997,N_1956,N_2128);
and U2998 (N_2998,N_1975,N_2354);
nor U2999 (N_2999,N_2311,N_1668);
nand U3000 (N_3000,N_1666,N_1533);
and U3001 (N_3001,N_1698,N_1943);
xnor U3002 (N_3002,N_2286,N_1733);
nor U3003 (N_3003,N_2221,N_1360);
or U3004 (N_3004,N_1721,N_2337);
or U3005 (N_3005,N_1639,N_1459);
and U3006 (N_3006,N_1290,N_2373);
nor U3007 (N_3007,N_1349,N_1696);
xnor U3008 (N_3008,N_1804,N_2047);
or U3009 (N_3009,N_2182,N_1820);
and U3010 (N_3010,N_1419,N_1301);
nor U3011 (N_3011,N_2192,N_1516);
or U3012 (N_3012,N_1848,N_1342);
nor U3013 (N_3013,N_2368,N_1553);
nor U3014 (N_3014,N_1954,N_1486);
nand U3015 (N_3015,N_1612,N_1492);
xnor U3016 (N_3016,N_2429,N_1502);
nand U3017 (N_3017,N_2347,N_1759);
and U3018 (N_3018,N_1907,N_1384);
nor U3019 (N_3019,N_2111,N_2377);
nor U3020 (N_3020,N_2297,N_1936);
and U3021 (N_3021,N_1744,N_2208);
nor U3022 (N_3022,N_1878,N_1935);
nand U3023 (N_3023,N_2489,N_2176);
and U3024 (N_3024,N_2123,N_2462);
and U3025 (N_3025,N_1283,N_2273);
or U3026 (N_3026,N_1545,N_2387);
nor U3027 (N_3027,N_1843,N_2497);
nand U3028 (N_3028,N_2268,N_1428);
xor U3029 (N_3029,N_1770,N_2343);
xnor U3030 (N_3030,N_1333,N_1983);
xor U3031 (N_3031,N_1998,N_2365);
xnor U3032 (N_3032,N_2319,N_1277);
nand U3033 (N_3033,N_2282,N_2371);
and U3034 (N_3034,N_1617,N_1375);
xnor U3035 (N_3035,N_1715,N_1995);
or U3036 (N_3036,N_2260,N_1844);
xnor U3037 (N_3037,N_1350,N_1429);
and U3038 (N_3038,N_2044,N_1572);
nand U3039 (N_3039,N_2482,N_2184);
nor U3040 (N_3040,N_2308,N_1567);
or U3041 (N_3041,N_2425,N_2003);
nor U3042 (N_3042,N_1337,N_1364);
nand U3043 (N_3043,N_2474,N_1404);
nand U3044 (N_3044,N_1439,N_1499);
or U3045 (N_3045,N_2057,N_1554);
and U3046 (N_3046,N_2259,N_1708);
nand U3047 (N_3047,N_1836,N_1678);
or U3048 (N_3048,N_2112,N_1285);
and U3049 (N_3049,N_2161,N_2217);
nor U3050 (N_3050,N_2402,N_1743);
xnor U3051 (N_3051,N_2239,N_1274);
nand U3052 (N_3052,N_1336,N_1573);
nor U3053 (N_3053,N_1412,N_2136);
xnor U3054 (N_3054,N_2276,N_1608);
and U3055 (N_3055,N_1976,N_1821);
nor U3056 (N_3056,N_1387,N_1792);
xnor U3057 (N_3057,N_2408,N_1340);
and U3058 (N_3058,N_1393,N_1835);
xor U3059 (N_3059,N_1677,N_1581);
or U3060 (N_3060,N_2216,N_1319);
and U3061 (N_3061,N_2467,N_2140);
and U3062 (N_3062,N_1345,N_1808);
or U3063 (N_3063,N_1299,N_1321);
nor U3064 (N_3064,N_1740,N_2456);
xnor U3065 (N_3065,N_2056,N_2010);
nand U3066 (N_3066,N_1853,N_1270);
nor U3067 (N_3067,N_1952,N_2008);
nand U3068 (N_3068,N_1524,N_2345);
nand U3069 (N_3069,N_1875,N_1659);
or U3070 (N_3070,N_1426,N_1453);
or U3071 (N_3071,N_1327,N_2101);
nand U3072 (N_3072,N_2323,N_1923);
nand U3073 (N_3073,N_1294,N_1863);
or U3074 (N_3074,N_2278,N_1753);
nor U3075 (N_3075,N_1739,N_2472);
nor U3076 (N_3076,N_2404,N_1584);
nand U3077 (N_3077,N_2063,N_1947);
or U3078 (N_3078,N_2296,N_2465);
nand U3079 (N_3079,N_1507,N_1815);
nand U3080 (N_3080,N_2317,N_2231);
nor U3081 (N_3081,N_1555,N_1711);
or U3082 (N_3082,N_1807,N_2004);
and U3083 (N_3083,N_1546,N_2194);
or U3084 (N_3084,N_1437,N_1720);
nor U3085 (N_3085,N_2262,N_2459);
nor U3086 (N_3086,N_1861,N_1541);
or U3087 (N_3087,N_1829,N_1962);
nor U3088 (N_3088,N_1272,N_2098);
and U3089 (N_3089,N_1994,N_1756);
and U3090 (N_3090,N_1592,N_2115);
nor U3091 (N_3091,N_1431,N_1300);
xnor U3092 (N_3092,N_2212,N_1446);
xor U3093 (N_3093,N_1542,N_1354);
nor U3094 (N_3094,N_1968,N_1652);
and U3095 (N_3095,N_1818,N_2417);
nor U3096 (N_3096,N_1955,N_1908);
or U3097 (N_3097,N_2054,N_2147);
nor U3098 (N_3098,N_2193,N_1775);
nor U3099 (N_3099,N_1658,N_2418);
nand U3100 (N_3100,N_2031,N_2103);
nand U3101 (N_3101,N_2419,N_2016);
or U3102 (N_3102,N_1692,N_1570);
nand U3103 (N_3103,N_1353,N_1391);
or U3104 (N_3104,N_2168,N_2384);
xnor U3105 (N_3105,N_1697,N_1410);
nand U3106 (N_3106,N_2012,N_1735);
and U3107 (N_3107,N_1632,N_2055);
nor U3108 (N_3108,N_1988,N_1306);
and U3109 (N_3109,N_1788,N_1559);
nor U3110 (N_3110,N_2494,N_1860);
or U3111 (N_3111,N_1442,N_1600);
nor U3112 (N_3112,N_2131,N_2079);
nand U3113 (N_3113,N_2290,N_2144);
xnor U3114 (N_3114,N_1979,N_2430);
nor U3115 (N_3115,N_2241,N_2191);
nand U3116 (N_3116,N_1879,N_2431);
or U3117 (N_3117,N_1675,N_1562);
and U3118 (N_3118,N_1388,N_1363);
xnor U3119 (N_3119,N_2053,N_2358);
and U3120 (N_3120,N_1990,N_1910);
xnor U3121 (N_3121,N_1331,N_1291);
nor U3122 (N_3122,N_1635,N_2477);
nand U3123 (N_3123,N_1803,N_1296);
nor U3124 (N_3124,N_1452,N_2224);
nand U3125 (N_3125,N_1385,N_2276);
and U3126 (N_3126,N_1602,N_1748);
and U3127 (N_3127,N_2397,N_1623);
or U3128 (N_3128,N_2044,N_1585);
nor U3129 (N_3129,N_2063,N_2381);
nand U3130 (N_3130,N_1706,N_1419);
nor U3131 (N_3131,N_2414,N_2316);
nor U3132 (N_3132,N_2284,N_1774);
nor U3133 (N_3133,N_1988,N_2071);
nand U3134 (N_3134,N_2399,N_1893);
nor U3135 (N_3135,N_2262,N_2016);
and U3136 (N_3136,N_1330,N_1368);
nor U3137 (N_3137,N_2197,N_1967);
nor U3138 (N_3138,N_1899,N_2199);
nor U3139 (N_3139,N_1359,N_1886);
nor U3140 (N_3140,N_2219,N_1532);
nand U3141 (N_3141,N_1775,N_1615);
xnor U3142 (N_3142,N_1473,N_1534);
nand U3143 (N_3143,N_1485,N_2156);
or U3144 (N_3144,N_1762,N_1753);
nand U3145 (N_3145,N_1541,N_2331);
or U3146 (N_3146,N_1635,N_2162);
nand U3147 (N_3147,N_2347,N_1904);
xor U3148 (N_3148,N_2392,N_1433);
nand U3149 (N_3149,N_2165,N_2257);
or U3150 (N_3150,N_2306,N_1774);
nor U3151 (N_3151,N_2394,N_2206);
xor U3152 (N_3152,N_2405,N_1285);
nand U3153 (N_3153,N_1658,N_2244);
and U3154 (N_3154,N_1656,N_2082);
nand U3155 (N_3155,N_1770,N_1706);
nand U3156 (N_3156,N_2075,N_1937);
nor U3157 (N_3157,N_2070,N_2349);
xnor U3158 (N_3158,N_1551,N_2072);
nand U3159 (N_3159,N_2186,N_1513);
nor U3160 (N_3160,N_2182,N_2330);
or U3161 (N_3161,N_2493,N_1399);
nor U3162 (N_3162,N_2445,N_1965);
nand U3163 (N_3163,N_1611,N_1716);
nand U3164 (N_3164,N_2183,N_1482);
xor U3165 (N_3165,N_1669,N_2060);
or U3166 (N_3166,N_1854,N_2179);
xor U3167 (N_3167,N_2148,N_1574);
and U3168 (N_3168,N_2293,N_1885);
xor U3169 (N_3169,N_2006,N_2397);
and U3170 (N_3170,N_1396,N_1695);
and U3171 (N_3171,N_1312,N_1569);
and U3172 (N_3172,N_1328,N_1312);
nor U3173 (N_3173,N_1493,N_2476);
and U3174 (N_3174,N_1804,N_2402);
xor U3175 (N_3175,N_1454,N_1708);
or U3176 (N_3176,N_2408,N_1813);
and U3177 (N_3177,N_1844,N_1793);
nand U3178 (N_3178,N_1512,N_1327);
or U3179 (N_3179,N_2087,N_1267);
or U3180 (N_3180,N_2444,N_1343);
nor U3181 (N_3181,N_2273,N_2100);
nand U3182 (N_3182,N_1348,N_2362);
or U3183 (N_3183,N_1755,N_1989);
xor U3184 (N_3184,N_1971,N_1528);
and U3185 (N_3185,N_2033,N_2446);
xor U3186 (N_3186,N_1323,N_1357);
and U3187 (N_3187,N_1747,N_2013);
nor U3188 (N_3188,N_2275,N_2329);
or U3189 (N_3189,N_1352,N_1859);
xnor U3190 (N_3190,N_1514,N_2129);
nor U3191 (N_3191,N_1921,N_1860);
xor U3192 (N_3192,N_1250,N_1817);
or U3193 (N_3193,N_1303,N_2326);
nor U3194 (N_3194,N_1982,N_2029);
nor U3195 (N_3195,N_2025,N_2376);
xnor U3196 (N_3196,N_2018,N_1872);
nor U3197 (N_3197,N_1586,N_1685);
or U3198 (N_3198,N_1487,N_1544);
xor U3199 (N_3199,N_2453,N_1718);
nand U3200 (N_3200,N_1845,N_2324);
nor U3201 (N_3201,N_1918,N_2140);
nor U3202 (N_3202,N_1661,N_2380);
nand U3203 (N_3203,N_1615,N_2022);
xnor U3204 (N_3204,N_1278,N_2078);
xnor U3205 (N_3205,N_1263,N_1412);
nand U3206 (N_3206,N_2410,N_1966);
or U3207 (N_3207,N_1993,N_1545);
xor U3208 (N_3208,N_1686,N_2359);
and U3209 (N_3209,N_1387,N_1767);
nand U3210 (N_3210,N_1676,N_1432);
or U3211 (N_3211,N_1698,N_2073);
or U3212 (N_3212,N_2054,N_2154);
and U3213 (N_3213,N_1685,N_2235);
nor U3214 (N_3214,N_1529,N_1619);
and U3215 (N_3215,N_1581,N_2052);
nor U3216 (N_3216,N_2396,N_2248);
nand U3217 (N_3217,N_2408,N_1727);
xor U3218 (N_3218,N_1345,N_1450);
nand U3219 (N_3219,N_2121,N_2211);
nor U3220 (N_3220,N_2446,N_2211);
xor U3221 (N_3221,N_1359,N_1960);
and U3222 (N_3222,N_1879,N_2021);
nor U3223 (N_3223,N_1743,N_1543);
and U3224 (N_3224,N_1274,N_1430);
xnor U3225 (N_3225,N_2464,N_2204);
xor U3226 (N_3226,N_1400,N_2266);
or U3227 (N_3227,N_1633,N_1729);
or U3228 (N_3228,N_1587,N_1574);
nand U3229 (N_3229,N_1677,N_1788);
and U3230 (N_3230,N_2427,N_2256);
nand U3231 (N_3231,N_1498,N_2160);
and U3232 (N_3232,N_2035,N_1994);
nand U3233 (N_3233,N_1619,N_1750);
or U3234 (N_3234,N_1841,N_2027);
and U3235 (N_3235,N_1671,N_1399);
or U3236 (N_3236,N_2258,N_2066);
xnor U3237 (N_3237,N_1507,N_2432);
or U3238 (N_3238,N_1468,N_2411);
xnor U3239 (N_3239,N_2149,N_1701);
nand U3240 (N_3240,N_2211,N_2325);
xnor U3241 (N_3241,N_1355,N_1957);
or U3242 (N_3242,N_2066,N_2184);
or U3243 (N_3243,N_2116,N_1678);
xor U3244 (N_3244,N_1312,N_1282);
nand U3245 (N_3245,N_2217,N_1386);
nand U3246 (N_3246,N_2198,N_2152);
or U3247 (N_3247,N_1303,N_2268);
and U3248 (N_3248,N_1665,N_2123);
nor U3249 (N_3249,N_2193,N_2187);
nor U3250 (N_3250,N_2284,N_2033);
nor U3251 (N_3251,N_1780,N_2104);
xor U3252 (N_3252,N_1982,N_1752);
xor U3253 (N_3253,N_1372,N_1620);
and U3254 (N_3254,N_1309,N_1271);
or U3255 (N_3255,N_2332,N_2406);
nor U3256 (N_3256,N_1817,N_2007);
nand U3257 (N_3257,N_2292,N_2458);
or U3258 (N_3258,N_2310,N_1698);
nor U3259 (N_3259,N_1252,N_2074);
nand U3260 (N_3260,N_1284,N_1872);
nor U3261 (N_3261,N_2078,N_1764);
nand U3262 (N_3262,N_1426,N_2314);
xnor U3263 (N_3263,N_1707,N_1369);
nor U3264 (N_3264,N_1923,N_1766);
xnor U3265 (N_3265,N_2052,N_1261);
and U3266 (N_3266,N_1974,N_1289);
nand U3267 (N_3267,N_1940,N_1797);
nand U3268 (N_3268,N_2143,N_1503);
nand U3269 (N_3269,N_1654,N_1259);
nand U3270 (N_3270,N_1809,N_1408);
xor U3271 (N_3271,N_2272,N_1326);
or U3272 (N_3272,N_1862,N_1496);
xnor U3273 (N_3273,N_2265,N_1294);
xnor U3274 (N_3274,N_2498,N_1835);
or U3275 (N_3275,N_1547,N_1341);
nor U3276 (N_3276,N_1993,N_2408);
and U3277 (N_3277,N_1538,N_1851);
or U3278 (N_3278,N_2247,N_1602);
and U3279 (N_3279,N_1568,N_1847);
nand U3280 (N_3280,N_1422,N_2196);
xor U3281 (N_3281,N_1287,N_2471);
xnor U3282 (N_3282,N_1987,N_2190);
or U3283 (N_3283,N_2368,N_2448);
or U3284 (N_3284,N_2041,N_1403);
nor U3285 (N_3285,N_2410,N_1555);
and U3286 (N_3286,N_2221,N_1473);
nor U3287 (N_3287,N_2477,N_2341);
xor U3288 (N_3288,N_1998,N_1774);
and U3289 (N_3289,N_1909,N_1611);
nor U3290 (N_3290,N_2288,N_2355);
and U3291 (N_3291,N_1648,N_2263);
xor U3292 (N_3292,N_2123,N_1542);
and U3293 (N_3293,N_1715,N_1366);
nand U3294 (N_3294,N_2163,N_1674);
and U3295 (N_3295,N_1364,N_2249);
nand U3296 (N_3296,N_2005,N_1502);
nor U3297 (N_3297,N_1357,N_2162);
nor U3298 (N_3298,N_2324,N_1557);
nand U3299 (N_3299,N_2002,N_1439);
nor U3300 (N_3300,N_2431,N_2210);
xor U3301 (N_3301,N_2019,N_1285);
xor U3302 (N_3302,N_2460,N_2238);
nand U3303 (N_3303,N_1575,N_1970);
and U3304 (N_3304,N_2199,N_1399);
and U3305 (N_3305,N_1367,N_1994);
nand U3306 (N_3306,N_1660,N_2278);
nand U3307 (N_3307,N_2216,N_1442);
nor U3308 (N_3308,N_1414,N_1719);
or U3309 (N_3309,N_2213,N_1720);
xnor U3310 (N_3310,N_2086,N_2053);
nor U3311 (N_3311,N_1616,N_1368);
nor U3312 (N_3312,N_2078,N_1576);
or U3313 (N_3313,N_2363,N_1330);
nand U3314 (N_3314,N_2059,N_2305);
or U3315 (N_3315,N_1994,N_1300);
xnor U3316 (N_3316,N_2039,N_1646);
and U3317 (N_3317,N_2331,N_2244);
or U3318 (N_3318,N_1934,N_2488);
and U3319 (N_3319,N_2472,N_1832);
and U3320 (N_3320,N_2092,N_1271);
nor U3321 (N_3321,N_1757,N_1536);
xnor U3322 (N_3322,N_2464,N_1543);
and U3323 (N_3323,N_1914,N_1388);
xnor U3324 (N_3324,N_1287,N_1493);
nor U3325 (N_3325,N_1251,N_2384);
or U3326 (N_3326,N_2215,N_1920);
and U3327 (N_3327,N_1651,N_2030);
and U3328 (N_3328,N_2168,N_2288);
or U3329 (N_3329,N_1620,N_2426);
xor U3330 (N_3330,N_1879,N_1346);
and U3331 (N_3331,N_1551,N_2478);
nand U3332 (N_3332,N_2382,N_2135);
xor U3333 (N_3333,N_2405,N_1959);
or U3334 (N_3334,N_1602,N_1991);
xnor U3335 (N_3335,N_1533,N_1925);
nor U3336 (N_3336,N_1526,N_1745);
and U3337 (N_3337,N_1965,N_1585);
or U3338 (N_3338,N_2397,N_1251);
nand U3339 (N_3339,N_2170,N_1848);
or U3340 (N_3340,N_1957,N_1474);
xnor U3341 (N_3341,N_1348,N_1488);
nor U3342 (N_3342,N_1468,N_1985);
and U3343 (N_3343,N_2148,N_2041);
nor U3344 (N_3344,N_1420,N_1996);
and U3345 (N_3345,N_1443,N_2003);
xor U3346 (N_3346,N_2468,N_1581);
or U3347 (N_3347,N_1464,N_1941);
nor U3348 (N_3348,N_2061,N_2391);
nand U3349 (N_3349,N_1372,N_2062);
or U3350 (N_3350,N_1713,N_1500);
or U3351 (N_3351,N_1368,N_2390);
or U3352 (N_3352,N_2202,N_2099);
xor U3353 (N_3353,N_2212,N_1992);
xor U3354 (N_3354,N_1282,N_1896);
xnor U3355 (N_3355,N_2095,N_2342);
or U3356 (N_3356,N_2069,N_1784);
or U3357 (N_3357,N_2488,N_1347);
xnor U3358 (N_3358,N_2085,N_1759);
nor U3359 (N_3359,N_2034,N_1522);
nor U3360 (N_3360,N_2479,N_2277);
xnor U3361 (N_3361,N_1497,N_2157);
nand U3362 (N_3362,N_1446,N_1274);
xor U3363 (N_3363,N_1470,N_1513);
nand U3364 (N_3364,N_1922,N_2038);
and U3365 (N_3365,N_1848,N_1829);
and U3366 (N_3366,N_1622,N_1811);
and U3367 (N_3367,N_1264,N_1352);
and U3368 (N_3368,N_2069,N_2028);
and U3369 (N_3369,N_1250,N_1668);
and U3370 (N_3370,N_1255,N_1623);
nand U3371 (N_3371,N_2257,N_1910);
or U3372 (N_3372,N_2005,N_1843);
and U3373 (N_3373,N_1534,N_1503);
or U3374 (N_3374,N_1980,N_1515);
or U3375 (N_3375,N_1333,N_1726);
or U3376 (N_3376,N_2477,N_2400);
xor U3377 (N_3377,N_2478,N_2191);
nand U3378 (N_3378,N_2060,N_1779);
nand U3379 (N_3379,N_2135,N_2284);
nor U3380 (N_3380,N_1651,N_2019);
or U3381 (N_3381,N_1410,N_2174);
or U3382 (N_3382,N_2440,N_1515);
and U3383 (N_3383,N_1275,N_1514);
xor U3384 (N_3384,N_1532,N_1274);
nand U3385 (N_3385,N_1638,N_1844);
xor U3386 (N_3386,N_2359,N_2301);
nor U3387 (N_3387,N_2059,N_2496);
and U3388 (N_3388,N_2139,N_1461);
nor U3389 (N_3389,N_1898,N_2482);
nor U3390 (N_3390,N_1982,N_1359);
nand U3391 (N_3391,N_1566,N_1696);
or U3392 (N_3392,N_1557,N_2033);
and U3393 (N_3393,N_2118,N_1822);
nand U3394 (N_3394,N_1309,N_1743);
nand U3395 (N_3395,N_2263,N_2097);
or U3396 (N_3396,N_2204,N_2055);
and U3397 (N_3397,N_1997,N_2440);
nand U3398 (N_3398,N_1698,N_2367);
xor U3399 (N_3399,N_2177,N_1937);
nand U3400 (N_3400,N_1717,N_2231);
nand U3401 (N_3401,N_1586,N_1725);
or U3402 (N_3402,N_1276,N_1853);
nor U3403 (N_3403,N_1415,N_1800);
nand U3404 (N_3404,N_1509,N_1590);
nor U3405 (N_3405,N_2186,N_2468);
or U3406 (N_3406,N_2464,N_2482);
or U3407 (N_3407,N_1423,N_1899);
nor U3408 (N_3408,N_1597,N_1761);
nand U3409 (N_3409,N_1305,N_2456);
or U3410 (N_3410,N_1722,N_1312);
nand U3411 (N_3411,N_2450,N_1824);
nor U3412 (N_3412,N_2322,N_2497);
and U3413 (N_3413,N_2235,N_1742);
nand U3414 (N_3414,N_1805,N_2140);
xor U3415 (N_3415,N_1963,N_2463);
and U3416 (N_3416,N_1281,N_1486);
or U3417 (N_3417,N_2211,N_2355);
or U3418 (N_3418,N_2374,N_2312);
and U3419 (N_3419,N_1404,N_1901);
xnor U3420 (N_3420,N_1596,N_2403);
xnor U3421 (N_3421,N_1412,N_2373);
nand U3422 (N_3422,N_2210,N_1988);
nor U3423 (N_3423,N_1672,N_1795);
nand U3424 (N_3424,N_2146,N_1903);
or U3425 (N_3425,N_1304,N_1843);
xnor U3426 (N_3426,N_1342,N_2181);
nor U3427 (N_3427,N_2412,N_1292);
and U3428 (N_3428,N_2277,N_2080);
xnor U3429 (N_3429,N_1412,N_1633);
xnor U3430 (N_3430,N_1603,N_1860);
nor U3431 (N_3431,N_1713,N_2169);
and U3432 (N_3432,N_1417,N_2297);
or U3433 (N_3433,N_1260,N_1413);
or U3434 (N_3434,N_2194,N_1590);
nand U3435 (N_3435,N_2173,N_2406);
nand U3436 (N_3436,N_1267,N_1874);
xor U3437 (N_3437,N_1490,N_2339);
or U3438 (N_3438,N_1792,N_2204);
xnor U3439 (N_3439,N_1979,N_1276);
nor U3440 (N_3440,N_1872,N_1619);
xnor U3441 (N_3441,N_2091,N_1619);
nand U3442 (N_3442,N_2224,N_1735);
xnor U3443 (N_3443,N_1973,N_1251);
and U3444 (N_3444,N_2392,N_2430);
xnor U3445 (N_3445,N_1854,N_1423);
xnor U3446 (N_3446,N_1497,N_1301);
nor U3447 (N_3447,N_1703,N_1456);
or U3448 (N_3448,N_1663,N_1539);
nand U3449 (N_3449,N_1425,N_2026);
and U3450 (N_3450,N_2181,N_1267);
xor U3451 (N_3451,N_2452,N_1792);
nand U3452 (N_3452,N_1782,N_2045);
xnor U3453 (N_3453,N_2302,N_1603);
nor U3454 (N_3454,N_2280,N_1845);
or U3455 (N_3455,N_2362,N_2341);
or U3456 (N_3456,N_1439,N_1772);
nor U3457 (N_3457,N_2085,N_2487);
xnor U3458 (N_3458,N_1749,N_1714);
nor U3459 (N_3459,N_1411,N_1859);
nand U3460 (N_3460,N_1953,N_2430);
and U3461 (N_3461,N_2249,N_1311);
and U3462 (N_3462,N_1459,N_1939);
or U3463 (N_3463,N_1921,N_2167);
or U3464 (N_3464,N_1251,N_1396);
nor U3465 (N_3465,N_1730,N_2314);
nand U3466 (N_3466,N_2068,N_2306);
nor U3467 (N_3467,N_2046,N_1643);
nor U3468 (N_3468,N_1807,N_2383);
nor U3469 (N_3469,N_1288,N_1388);
nor U3470 (N_3470,N_2017,N_1654);
and U3471 (N_3471,N_1833,N_2145);
nor U3472 (N_3472,N_2289,N_2094);
or U3473 (N_3473,N_1935,N_1909);
nor U3474 (N_3474,N_1759,N_2084);
xor U3475 (N_3475,N_1973,N_2072);
and U3476 (N_3476,N_1460,N_1948);
or U3477 (N_3477,N_1791,N_2363);
or U3478 (N_3478,N_1737,N_2393);
nand U3479 (N_3479,N_1732,N_1281);
nor U3480 (N_3480,N_2025,N_1433);
nor U3481 (N_3481,N_1964,N_2149);
and U3482 (N_3482,N_1797,N_1299);
xnor U3483 (N_3483,N_1731,N_1889);
nor U3484 (N_3484,N_2060,N_1287);
and U3485 (N_3485,N_1375,N_1751);
nor U3486 (N_3486,N_1533,N_1754);
and U3487 (N_3487,N_2386,N_1579);
nand U3488 (N_3488,N_2395,N_2322);
nor U3489 (N_3489,N_1919,N_1283);
or U3490 (N_3490,N_1769,N_1313);
xnor U3491 (N_3491,N_1267,N_2342);
xor U3492 (N_3492,N_1630,N_2351);
xor U3493 (N_3493,N_2455,N_1765);
and U3494 (N_3494,N_2443,N_1901);
nand U3495 (N_3495,N_1730,N_1950);
xor U3496 (N_3496,N_2390,N_1621);
xnor U3497 (N_3497,N_2106,N_1477);
nand U3498 (N_3498,N_1373,N_1332);
xor U3499 (N_3499,N_1312,N_1762);
and U3500 (N_3500,N_1441,N_2486);
or U3501 (N_3501,N_1894,N_1429);
xor U3502 (N_3502,N_2207,N_1411);
or U3503 (N_3503,N_2411,N_2028);
nand U3504 (N_3504,N_1542,N_1321);
or U3505 (N_3505,N_1568,N_2354);
or U3506 (N_3506,N_1696,N_1766);
nand U3507 (N_3507,N_2378,N_1981);
and U3508 (N_3508,N_1462,N_1262);
or U3509 (N_3509,N_1474,N_1380);
and U3510 (N_3510,N_1552,N_2006);
and U3511 (N_3511,N_1631,N_2329);
and U3512 (N_3512,N_2163,N_2363);
nand U3513 (N_3513,N_1745,N_2391);
and U3514 (N_3514,N_2315,N_2364);
and U3515 (N_3515,N_1415,N_2275);
or U3516 (N_3516,N_2128,N_1652);
nor U3517 (N_3517,N_1604,N_2431);
nand U3518 (N_3518,N_2065,N_1630);
nand U3519 (N_3519,N_2488,N_1563);
nor U3520 (N_3520,N_2042,N_2218);
nor U3521 (N_3521,N_1648,N_1649);
or U3522 (N_3522,N_2154,N_2373);
xnor U3523 (N_3523,N_2259,N_2066);
nand U3524 (N_3524,N_2292,N_1354);
or U3525 (N_3525,N_2161,N_2004);
xor U3526 (N_3526,N_1814,N_2158);
and U3527 (N_3527,N_1753,N_2220);
nor U3528 (N_3528,N_1377,N_2488);
and U3529 (N_3529,N_1856,N_2191);
nor U3530 (N_3530,N_1838,N_1474);
nor U3531 (N_3531,N_1510,N_1827);
nand U3532 (N_3532,N_1747,N_1964);
and U3533 (N_3533,N_1612,N_2189);
nand U3534 (N_3534,N_2029,N_1595);
and U3535 (N_3535,N_2313,N_1526);
xor U3536 (N_3536,N_2355,N_1648);
nand U3537 (N_3537,N_2381,N_1837);
nand U3538 (N_3538,N_1287,N_1608);
and U3539 (N_3539,N_1464,N_1473);
or U3540 (N_3540,N_1554,N_1783);
nor U3541 (N_3541,N_2458,N_1863);
nor U3542 (N_3542,N_1851,N_1426);
nand U3543 (N_3543,N_1369,N_1807);
nand U3544 (N_3544,N_1905,N_2134);
xor U3545 (N_3545,N_2270,N_1429);
and U3546 (N_3546,N_1387,N_2421);
nor U3547 (N_3547,N_2095,N_1462);
nor U3548 (N_3548,N_2042,N_1634);
nand U3549 (N_3549,N_1855,N_1856);
xnor U3550 (N_3550,N_1705,N_2403);
nor U3551 (N_3551,N_2406,N_1974);
or U3552 (N_3552,N_2473,N_1777);
nor U3553 (N_3553,N_2083,N_1343);
nand U3554 (N_3554,N_1860,N_1601);
nand U3555 (N_3555,N_1564,N_2188);
nor U3556 (N_3556,N_1619,N_2481);
nand U3557 (N_3557,N_1998,N_2263);
or U3558 (N_3558,N_2286,N_1903);
and U3559 (N_3559,N_2183,N_1616);
nand U3560 (N_3560,N_2438,N_2124);
xor U3561 (N_3561,N_2196,N_1255);
xnor U3562 (N_3562,N_2499,N_1964);
and U3563 (N_3563,N_1537,N_1341);
xnor U3564 (N_3564,N_2063,N_1668);
or U3565 (N_3565,N_1904,N_1649);
xnor U3566 (N_3566,N_1323,N_1452);
and U3567 (N_3567,N_2379,N_2023);
nor U3568 (N_3568,N_1544,N_1301);
or U3569 (N_3569,N_1940,N_2078);
or U3570 (N_3570,N_2220,N_2404);
or U3571 (N_3571,N_1994,N_1530);
and U3572 (N_3572,N_1905,N_1394);
or U3573 (N_3573,N_2252,N_1501);
xor U3574 (N_3574,N_2143,N_1960);
nand U3575 (N_3575,N_1906,N_1287);
and U3576 (N_3576,N_1847,N_1747);
and U3577 (N_3577,N_1836,N_2480);
and U3578 (N_3578,N_2381,N_2019);
nand U3579 (N_3579,N_1557,N_1491);
nor U3580 (N_3580,N_1296,N_2039);
or U3581 (N_3581,N_1300,N_1997);
nor U3582 (N_3582,N_2166,N_1343);
xnor U3583 (N_3583,N_2041,N_2213);
nand U3584 (N_3584,N_2143,N_1922);
and U3585 (N_3585,N_2362,N_1346);
nand U3586 (N_3586,N_1442,N_2057);
or U3587 (N_3587,N_1881,N_1932);
or U3588 (N_3588,N_1757,N_1764);
or U3589 (N_3589,N_2241,N_2384);
or U3590 (N_3590,N_1553,N_2025);
and U3591 (N_3591,N_1706,N_1561);
or U3592 (N_3592,N_1799,N_2276);
xor U3593 (N_3593,N_1800,N_2282);
nor U3594 (N_3594,N_2347,N_1919);
nand U3595 (N_3595,N_1828,N_1529);
nor U3596 (N_3596,N_1519,N_1293);
and U3597 (N_3597,N_1646,N_1395);
nor U3598 (N_3598,N_1926,N_2301);
or U3599 (N_3599,N_2241,N_2298);
xor U3600 (N_3600,N_1424,N_1574);
and U3601 (N_3601,N_2070,N_1375);
or U3602 (N_3602,N_1321,N_1362);
and U3603 (N_3603,N_2267,N_1974);
and U3604 (N_3604,N_1983,N_1683);
nor U3605 (N_3605,N_1286,N_1814);
and U3606 (N_3606,N_1256,N_1968);
or U3607 (N_3607,N_1943,N_1625);
nor U3608 (N_3608,N_1310,N_1565);
nand U3609 (N_3609,N_1450,N_2037);
and U3610 (N_3610,N_1946,N_2013);
xnor U3611 (N_3611,N_1697,N_1950);
xnor U3612 (N_3612,N_2082,N_1344);
or U3613 (N_3613,N_2474,N_1257);
nand U3614 (N_3614,N_2223,N_1802);
nand U3615 (N_3615,N_2139,N_1776);
and U3616 (N_3616,N_1264,N_1338);
xnor U3617 (N_3617,N_1835,N_2161);
and U3618 (N_3618,N_1889,N_2411);
and U3619 (N_3619,N_2132,N_1574);
or U3620 (N_3620,N_2255,N_1446);
nand U3621 (N_3621,N_2026,N_1592);
xnor U3622 (N_3622,N_2473,N_2202);
xnor U3623 (N_3623,N_1294,N_1984);
or U3624 (N_3624,N_1482,N_1401);
xor U3625 (N_3625,N_1509,N_1931);
nand U3626 (N_3626,N_1291,N_2388);
nor U3627 (N_3627,N_2129,N_2078);
and U3628 (N_3628,N_2417,N_2431);
or U3629 (N_3629,N_1909,N_2309);
or U3630 (N_3630,N_1841,N_2082);
xnor U3631 (N_3631,N_1606,N_2443);
and U3632 (N_3632,N_1830,N_2483);
nand U3633 (N_3633,N_2464,N_1603);
or U3634 (N_3634,N_2126,N_2210);
xnor U3635 (N_3635,N_2325,N_2326);
or U3636 (N_3636,N_1539,N_1766);
nor U3637 (N_3637,N_1934,N_1312);
xor U3638 (N_3638,N_1993,N_2268);
and U3639 (N_3639,N_2140,N_2105);
xnor U3640 (N_3640,N_1849,N_2264);
or U3641 (N_3641,N_1315,N_2066);
or U3642 (N_3642,N_1871,N_2054);
nor U3643 (N_3643,N_2045,N_1751);
or U3644 (N_3644,N_2180,N_1634);
nand U3645 (N_3645,N_1448,N_1487);
or U3646 (N_3646,N_1552,N_1985);
xnor U3647 (N_3647,N_1959,N_1951);
xor U3648 (N_3648,N_1607,N_2012);
and U3649 (N_3649,N_1966,N_1430);
xnor U3650 (N_3650,N_1666,N_2317);
nand U3651 (N_3651,N_2102,N_1828);
xor U3652 (N_3652,N_1477,N_1446);
xnor U3653 (N_3653,N_1666,N_1775);
nor U3654 (N_3654,N_1347,N_1655);
xor U3655 (N_3655,N_1504,N_1484);
or U3656 (N_3656,N_1331,N_2202);
nand U3657 (N_3657,N_2335,N_2322);
nand U3658 (N_3658,N_1667,N_2065);
or U3659 (N_3659,N_1414,N_1372);
and U3660 (N_3660,N_2470,N_2241);
and U3661 (N_3661,N_1331,N_1448);
nand U3662 (N_3662,N_1559,N_2345);
and U3663 (N_3663,N_1290,N_1547);
xnor U3664 (N_3664,N_2152,N_1780);
nand U3665 (N_3665,N_2193,N_1314);
and U3666 (N_3666,N_1568,N_1964);
nand U3667 (N_3667,N_1586,N_1627);
nor U3668 (N_3668,N_2074,N_1804);
and U3669 (N_3669,N_2295,N_1870);
nor U3670 (N_3670,N_2193,N_1677);
or U3671 (N_3671,N_2421,N_1630);
xor U3672 (N_3672,N_2368,N_1536);
xnor U3673 (N_3673,N_2138,N_2080);
and U3674 (N_3674,N_2356,N_1414);
nor U3675 (N_3675,N_2374,N_2171);
nor U3676 (N_3676,N_2044,N_1890);
xor U3677 (N_3677,N_1534,N_2343);
xor U3678 (N_3678,N_2374,N_2241);
and U3679 (N_3679,N_1527,N_1725);
or U3680 (N_3680,N_1360,N_1819);
xor U3681 (N_3681,N_1475,N_1252);
or U3682 (N_3682,N_2297,N_1283);
and U3683 (N_3683,N_1409,N_1512);
or U3684 (N_3684,N_1688,N_1978);
and U3685 (N_3685,N_1506,N_2137);
and U3686 (N_3686,N_2257,N_2304);
and U3687 (N_3687,N_1781,N_1959);
or U3688 (N_3688,N_1845,N_1398);
nand U3689 (N_3689,N_1877,N_1327);
xor U3690 (N_3690,N_1841,N_2370);
nor U3691 (N_3691,N_2056,N_1481);
nor U3692 (N_3692,N_1252,N_2019);
or U3693 (N_3693,N_2376,N_1744);
and U3694 (N_3694,N_2094,N_2335);
xnor U3695 (N_3695,N_2136,N_1625);
nand U3696 (N_3696,N_2494,N_1986);
nor U3697 (N_3697,N_1487,N_2011);
nor U3698 (N_3698,N_1583,N_1799);
and U3699 (N_3699,N_1789,N_1308);
or U3700 (N_3700,N_1914,N_1831);
xnor U3701 (N_3701,N_1946,N_1956);
nand U3702 (N_3702,N_2077,N_1533);
nand U3703 (N_3703,N_1989,N_1488);
nor U3704 (N_3704,N_1326,N_2121);
and U3705 (N_3705,N_1265,N_1895);
and U3706 (N_3706,N_1544,N_1594);
xor U3707 (N_3707,N_1683,N_2069);
nor U3708 (N_3708,N_1590,N_2277);
xor U3709 (N_3709,N_2427,N_2408);
xnor U3710 (N_3710,N_1944,N_1917);
nand U3711 (N_3711,N_2282,N_2002);
nand U3712 (N_3712,N_1818,N_2447);
or U3713 (N_3713,N_1576,N_2003);
nor U3714 (N_3714,N_1861,N_1828);
or U3715 (N_3715,N_1781,N_1725);
xnor U3716 (N_3716,N_2350,N_1792);
and U3717 (N_3717,N_2016,N_1589);
and U3718 (N_3718,N_1632,N_2271);
nor U3719 (N_3719,N_1488,N_1325);
and U3720 (N_3720,N_1678,N_2011);
nand U3721 (N_3721,N_2335,N_1440);
nand U3722 (N_3722,N_2148,N_1351);
xnor U3723 (N_3723,N_2400,N_1450);
nor U3724 (N_3724,N_1905,N_1264);
nand U3725 (N_3725,N_2395,N_1510);
and U3726 (N_3726,N_2441,N_1671);
nor U3727 (N_3727,N_1424,N_2191);
xnor U3728 (N_3728,N_1995,N_1368);
nand U3729 (N_3729,N_1997,N_2379);
nand U3730 (N_3730,N_2039,N_2196);
nand U3731 (N_3731,N_1781,N_1293);
or U3732 (N_3732,N_1778,N_1907);
and U3733 (N_3733,N_1922,N_2127);
nor U3734 (N_3734,N_1382,N_1704);
xnor U3735 (N_3735,N_1909,N_1688);
nor U3736 (N_3736,N_2152,N_2288);
nor U3737 (N_3737,N_2477,N_2435);
nor U3738 (N_3738,N_1751,N_1654);
or U3739 (N_3739,N_1511,N_1261);
and U3740 (N_3740,N_2143,N_2164);
nand U3741 (N_3741,N_1306,N_1942);
nor U3742 (N_3742,N_1293,N_1434);
xor U3743 (N_3743,N_1573,N_2218);
xnor U3744 (N_3744,N_1389,N_1994);
or U3745 (N_3745,N_1917,N_1345);
nand U3746 (N_3746,N_1276,N_1626);
or U3747 (N_3747,N_1619,N_2434);
nor U3748 (N_3748,N_1459,N_1796);
or U3749 (N_3749,N_2117,N_1812);
xor U3750 (N_3750,N_3124,N_3421);
xor U3751 (N_3751,N_3031,N_2998);
xor U3752 (N_3752,N_3548,N_3603);
nor U3753 (N_3753,N_3168,N_3176);
nor U3754 (N_3754,N_3268,N_3660);
nor U3755 (N_3755,N_3149,N_3221);
nand U3756 (N_3756,N_3534,N_2759);
or U3757 (N_3757,N_2797,N_2733);
xor U3758 (N_3758,N_3506,N_2635);
and U3759 (N_3759,N_3036,N_3111);
xnor U3760 (N_3760,N_2852,N_3059);
nor U3761 (N_3761,N_3055,N_3077);
or U3762 (N_3762,N_3669,N_2732);
nor U3763 (N_3763,N_2615,N_3143);
nor U3764 (N_3764,N_3401,N_2906);
or U3765 (N_3765,N_3248,N_3241);
or U3766 (N_3766,N_2815,N_3123);
and U3767 (N_3767,N_3576,N_2739);
nand U3768 (N_3768,N_2646,N_2853);
xor U3769 (N_3769,N_2749,N_3621);
xnor U3770 (N_3770,N_3452,N_3395);
xor U3771 (N_3771,N_2526,N_3704);
and U3772 (N_3772,N_3304,N_2654);
or U3773 (N_3773,N_3458,N_3240);
xor U3774 (N_3774,N_2531,N_3723);
and U3775 (N_3775,N_3447,N_3233);
xnor U3776 (N_3776,N_2968,N_2913);
or U3777 (N_3777,N_2620,N_3373);
nor U3778 (N_3778,N_3379,N_3449);
and U3779 (N_3779,N_3126,N_3601);
and U3780 (N_3780,N_2515,N_2680);
nor U3781 (N_3781,N_3525,N_3316);
nor U3782 (N_3782,N_3004,N_2831);
nand U3783 (N_3783,N_3728,N_3343);
and U3784 (N_3784,N_2929,N_3205);
xnor U3785 (N_3785,N_3035,N_3054);
xor U3786 (N_3786,N_2773,N_2737);
or U3787 (N_3787,N_3299,N_2803);
and U3788 (N_3788,N_3554,N_2835);
nand U3789 (N_3789,N_3220,N_2789);
nor U3790 (N_3790,N_3228,N_3308);
or U3791 (N_3791,N_2518,N_3387);
nand U3792 (N_3792,N_3399,N_2763);
or U3793 (N_3793,N_2708,N_3337);
nor U3794 (N_3794,N_3737,N_3436);
and U3795 (N_3795,N_3027,N_3462);
and U3796 (N_3796,N_3607,N_3612);
nor U3797 (N_3797,N_3635,N_2500);
and U3798 (N_3798,N_3008,N_3508);
nor U3799 (N_3799,N_3650,N_2900);
and U3800 (N_3800,N_2948,N_2878);
nor U3801 (N_3801,N_3046,N_2805);
xor U3802 (N_3802,N_3667,N_2694);
xnor U3803 (N_3803,N_2921,N_3466);
or U3804 (N_3804,N_2765,N_3375);
nor U3805 (N_3805,N_2838,N_3403);
nor U3806 (N_3806,N_3353,N_2910);
nor U3807 (N_3807,N_2967,N_3504);
or U3808 (N_3808,N_3202,N_3376);
xor U3809 (N_3809,N_3632,N_3719);
nor U3810 (N_3810,N_3072,N_2975);
nor U3811 (N_3811,N_3345,N_2858);
or U3812 (N_3812,N_3679,N_3408);
nor U3813 (N_3813,N_2501,N_2795);
or U3814 (N_3814,N_3544,N_2991);
or U3815 (N_3815,N_3386,N_3060);
and U3816 (N_3816,N_2653,N_2939);
or U3817 (N_3817,N_2586,N_2801);
nand U3818 (N_3818,N_3450,N_2816);
nand U3819 (N_3819,N_2548,N_2879);
nand U3820 (N_3820,N_3006,N_2582);
nand U3821 (N_3821,N_2774,N_2788);
nor U3822 (N_3822,N_3562,N_3453);
and U3823 (N_3823,N_3573,N_2981);
nor U3824 (N_3824,N_3608,N_3252);
and U3825 (N_3825,N_3493,N_3367);
nor U3826 (N_3826,N_2748,N_2516);
xor U3827 (N_3827,N_2828,N_3583);
xor U3828 (N_3828,N_3477,N_3690);
nand U3829 (N_3829,N_2886,N_3135);
nand U3830 (N_3830,N_2741,N_3182);
nand U3831 (N_3831,N_2812,N_2692);
or U3832 (N_3832,N_3747,N_3223);
nand U3833 (N_3833,N_2833,N_2872);
xnor U3834 (N_3834,N_3340,N_2866);
or U3835 (N_3835,N_2603,N_3334);
nor U3836 (N_3836,N_2710,N_3362);
xnor U3837 (N_3837,N_3226,N_3575);
nand U3838 (N_3838,N_2982,N_2513);
or U3839 (N_3839,N_3084,N_2829);
and U3840 (N_3840,N_2924,N_2770);
nor U3841 (N_3841,N_3480,N_2817);
nand U3842 (N_3842,N_3701,N_2587);
xnor U3843 (N_3843,N_2905,N_2623);
and U3844 (N_3844,N_3582,N_2810);
or U3845 (N_3845,N_3198,N_3336);
or U3846 (N_3846,N_2811,N_3194);
xor U3847 (N_3847,N_2895,N_3237);
or U3848 (N_3848,N_3263,N_2999);
and U3849 (N_3849,N_3646,N_3630);
and U3850 (N_3850,N_3645,N_3225);
and U3851 (N_3851,N_2786,N_3350);
nand U3852 (N_3852,N_3000,N_2706);
or U3853 (N_3853,N_3075,N_3680);
xnor U3854 (N_3854,N_2976,N_3571);
and U3855 (N_3855,N_2836,N_2647);
xor U3856 (N_3856,N_3191,N_3030);
nor U3857 (N_3857,N_2989,N_3025);
xnor U3858 (N_3858,N_2691,N_2678);
and U3859 (N_3859,N_2940,N_3214);
and U3860 (N_3860,N_3500,N_3593);
nand U3861 (N_3861,N_2699,N_2532);
nor U3862 (N_3862,N_3201,N_2934);
or U3863 (N_3863,N_3101,N_2639);
and U3864 (N_3864,N_3016,N_3509);
and U3865 (N_3865,N_2775,N_2777);
and U3866 (N_3866,N_2963,N_2882);
and U3867 (N_3867,N_3352,N_2645);
and U3868 (N_3868,N_3749,N_2863);
and U3869 (N_3869,N_2630,N_3076);
nor U3870 (N_3870,N_3653,N_3611);
nand U3871 (N_3871,N_2588,N_2550);
or U3872 (N_3872,N_3717,N_2958);
nor U3873 (N_3873,N_2605,N_3090);
or U3874 (N_3874,N_3192,N_2555);
and U3875 (N_3875,N_2755,N_2674);
nor U3876 (N_3876,N_3427,N_2747);
and U3877 (N_3877,N_3157,N_3163);
nand U3878 (N_3878,N_3020,N_2937);
and U3879 (N_3879,N_2622,N_3393);
nand U3880 (N_3880,N_2712,N_3254);
xnor U3881 (N_3881,N_3446,N_2718);
nand U3882 (N_3882,N_3244,N_3445);
and U3883 (N_3883,N_3307,N_2941);
or U3884 (N_3884,N_3580,N_2577);
nand U3885 (N_3885,N_3066,N_3280);
nand U3886 (N_3886,N_3581,N_2822);
and U3887 (N_3887,N_2977,N_3670);
nor U3888 (N_3888,N_3112,N_2693);
nor U3889 (N_3889,N_3563,N_2746);
and U3890 (N_3890,N_3037,N_2602);
nor U3891 (N_3891,N_3570,N_2648);
nor U3892 (N_3892,N_3127,N_3012);
nor U3893 (N_3893,N_3309,N_3166);
nor U3894 (N_3894,N_3113,N_3114);
nor U3895 (N_3895,N_2709,N_2926);
nor U3896 (N_3896,N_3663,N_3491);
nor U3897 (N_3897,N_2856,N_2945);
and U3898 (N_3898,N_3619,N_2619);
nand U3899 (N_3899,N_3195,N_3468);
nor U3900 (N_3900,N_2543,N_2517);
and U3901 (N_3901,N_3292,N_3433);
nand U3902 (N_3902,N_3415,N_2964);
xnor U3903 (N_3903,N_2771,N_2781);
and U3904 (N_3904,N_3715,N_3410);
nor U3905 (N_3905,N_3222,N_2553);
nor U3906 (N_3906,N_3599,N_3539);
and U3907 (N_3907,N_2799,N_3486);
nand U3908 (N_3908,N_3301,N_2849);
nor U3909 (N_3909,N_2506,N_2606);
nor U3910 (N_3910,N_2508,N_3472);
nand U3911 (N_3911,N_2804,N_2861);
nand U3912 (N_3912,N_2626,N_3426);
and U3913 (N_3913,N_3569,N_3564);
and U3914 (N_3914,N_3411,N_2867);
xnor U3915 (N_3915,N_3043,N_3147);
and U3916 (N_3916,N_2881,N_3041);
and U3917 (N_3917,N_2840,N_3366);
or U3918 (N_3918,N_2808,N_3588);
nand U3919 (N_3919,N_3530,N_3626);
or U3920 (N_3920,N_2965,N_3034);
nand U3921 (N_3921,N_3361,N_3174);
or U3922 (N_3922,N_3229,N_3718);
and U3923 (N_3923,N_3091,N_2807);
nand U3924 (N_3924,N_2627,N_3134);
xnor U3925 (N_3925,N_3473,N_2806);
nor U3926 (N_3926,N_3290,N_3722);
nand U3927 (N_3927,N_3407,N_3437);
or U3928 (N_3928,N_2688,N_3203);
and U3929 (N_3929,N_3400,N_3496);
or U3930 (N_3930,N_2621,N_3227);
nor U3931 (N_3931,N_3311,N_3412);
nor U3932 (N_3932,N_2633,N_2898);
nand U3933 (N_3933,N_3049,N_2675);
and U3934 (N_3934,N_3079,N_2698);
or U3935 (N_3935,N_2841,N_2679);
xor U3936 (N_3936,N_3274,N_3546);
nand U3937 (N_3937,N_3305,N_3706);
nand U3938 (N_3938,N_3398,N_2656);
or U3939 (N_3939,N_3584,N_3488);
nor U3940 (N_3940,N_3142,N_3618);
or U3941 (N_3941,N_3131,N_3199);
or U3942 (N_3942,N_2962,N_3070);
and U3943 (N_3943,N_3655,N_3098);
or U3944 (N_3944,N_2969,N_3594);
xnor U3945 (N_3945,N_2604,N_3555);
or U3946 (N_3946,N_2735,N_2883);
xor U3947 (N_3947,N_3711,N_2785);
and U3948 (N_3948,N_2721,N_3110);
nor U3949 (N_3949,N_3120,N_2961);
nor U3950 (N_3950,N_3677,N_3319);
and U3951 (N_3951,N_3703,N_2903);
nor U3952 (N_3952,N_2848,N_2752);
nor U3953 (N_3953,N_3118,N_2844);
or U3954 (N_3954,N_3325,N_3013);
nor U3955 (N_3955,N_2578,N_3743);
or U3956 (N_3956,N_3464,N_3108);
nor U3957 (N_3957,N_3193,N_3172);
nand U3958 (N_3958,N_3627,N_3115);
and U3959 (N_3959,N_3604,N_2936);
and U3960 (N_3960,N_3015,N_3092);
nor U3961 (N_3961,N_3324,N_3200);
xnor U3962 (N_3962,N_3636,N_2511);
nand U3963 (N_3963,N_3139,N_2819);
nor U3964 (N_3964,N_3140,N_3094);
xor U3965 (N_3965,N_3207,N_2927);
xnor U3966 (N_3966,N_2640,N_3681);
or U3967 (N_3967,N_2728,N_2845);
nand U3968 (N_3968,N_3086,N_3318);
nand U3969 (N_3969,N_2682,N_3536);
xor U3970 (N_3970,N_3259,N_3726);
xnor U3971 (N_3971,N_3678,N_3406);
xor U3972 (N_3972,N_2673,N_2711);
nand U3973 (N_3973,N_3338,N_3187);
or U3974 (N_3974,N_2512,N_3721);
and U3975 (N_3975,N_3328,N_2932);
xor U3976 (N_3976,N_3662,N_2832);
or U3977 (N_3977,N_3087,N_3017);
xnor U3978 (N_3978,N_3208,N_3355);
nand U3979 (N_3979,N_2760,N_2717);
xor U3980 (N_3980,N_3725,N_3740);
nor U3981 (N_3981,N_2909,N_3010);
nand U3982 (N_3982,N_3130,N_3005);
nor U3983 (N_3983,N_3026,N_3219);
and U3984 (N_3984,N_2534,N_2834);
or U3985 (N_3985,N_3665,N_3342);
and U3986 (N_3986,N_2670,N_3011);
nor U3987 (N_3987,N_3204,N_3730);
xnor U3988 (N_3988,N_2661,N_3556);
or U3989 (N_3989,N_2573,N_3093);
nor U3990 (N_3990,N_3152,N_3215);
nor U3991 (N_3991,N_2783,N_2876);
nor U3992 (N_3992,N_3652,N_3712);
nand U3993 (N_3993,N_2756,N_3489);
nand U3994 (N_3994,N_2618,N_2923);
and U3995 (N_3995,N_2689,N_3514);
xnor U3996 (N_3996,N_3184,N_2624);
or U3997 (N_3997,N_3674,N_3475);
nor U3998 (N_3998,N_2901,N_3413);
nor U3999 (N_3999,N_3592,N_3501);
nor U4000 (N_4000,N_3541,N_2649);
or U4001 (N_4001,N_3616,N_3145);
nand U4002 (N_4002,N_2970,N_3245);
or U4003 (N_4003,N_2600,N_3344);
or U4004 (N_4004,N_3298,N_2714);
xor U4005 (N_4005,N_2683,N_3171);
xor U4006 (N_4006,N_2850,N_3642);
xnor U4007 (N_4007,N_2652,N_3423);
nor U4008 (N_4008,N_2854,N_2769);
and U4009 (N_4009,N_3369,N_2597);
nor U4010 (N_4010,N_3380,N_3476);
or U4011 (N_4011,N_2601,N_2719);
and U4012 (N_4012,N_2542,N_3511);
nand U4013 (N_4013,N_3175,N_2942);
and U4014 (N_4014,N_3302,N_2726);
or U4015 (N_4015,N_3553,N_2571);
nor U4016 (N_4016,N_2520,N_3422);
and U4017 (N_4017,N_3467,N_2826);
nand U4018 (N_4018,N_2790,N_3161);
or U4019 (N_4019,N_2595,N_3064);
or U4020 (N_4020,N_3738,N_3210);
nand U4021 (N_4021,N_3474,N_2556);
and U4022 (N_4022,N_2920,N_3289);
and U4023 (N_4023,N_2946,N_2701);
and U4024 (N_4024,N_2902,N_3088);
nand U4025 (N_4025,N_3479,N_3609);
nand U4026 (N_4026,N_3080,N_3540);
nor U4027 (N_4027,N_3186,N_3656);
and U4028 (N_4028,N_3424,N_3409);
nand U4029 (N_4029,N_2782,N_2736);
xnor U4030 (N_4030,N_2592,N_3494);
nor U4031 (N_4031,N_2884,N_3487);
nand U4032 (N_4032,N_3552,N_2504);
or U4033 (N_4033,N_3365,N_2796);
xor U4034 (N_4034,N_2744,N_2598);
nand U4035 (N_4035,N_2957,N_2658);
nand U4036 (N_4036,N_2994,N_3471);
nand U4037 (N_4037,N_2643,N_3359);
and U4038 (N_4038,N_2824,N_2896);
and U4039 (N_4039,N_3668,N_3615);
nor U4040 (N_4040,N_3658,N_3062);
or U4041 (N_4041,N_2993,N_2912);
nand U4042 (N_4042,N_2891,N_3516);
and U4043 (N_4043,N_2702,N_2916);
nand U4044 (N_4044,N_3550,N_2537);
nor U4045 (N_4045,N_2549,N_2608);
nand U4046 (N_4046,N_3300,N_2636);
and U4047 (N_4047,N_3589,N_3264);
and U4048 (N_4048,N_3057,N_3461);
or U4049 (N_4049,N_3420,N_3105);
nand U4050 (N_4050,N_2557,N_3425);
and U4051 (N_4051,N_3047,N_3377);
nand U4052 (N_4052,N_2984,N_3524);
nand U4053 (N_4053,N_3051,N_3465);
and U4054 (N_4054,N_2935,N_2851);
or U4055 (N_4055,N_2651,N_3039);
xor U4056 (N_4056,N_3456,N_3396);
xor U4057 (N_4057,N_3158,N_3170);
or U4058 (N_4058,N_3330,N_2655);
and U4059 (N_4059,N_2928,N_3081);
and U4060 (N_4060,N_3694,N_3390);
or U4061 (N_4061,N_3598,N_2614);
xor U4062 (N_4062,N_3372,N_2596);
xnor U4063 (N_4063,N_3063,N_3071);
nor U4064 (N_4064,N_2566,N_2672);
nand U4065 (N_4065,N_3234,N_3572);
nor U4066 (N_4066,N_2669,N_3623);
and U4067 (N_4067,N_3748,N_3284);
xnor U4068 (N_4068,N_3526,N_3360);
xnor U4069 (N_4069,N_3083,N_2792);
nor U4070 (N_4070,N_2842,N_3249);
xor U4071 (N_4071,N_2581,N_2992);
xor U4072 (N_4072,N_3378,N_3414);
nor U4073 (N_4073,N_3082,N_3348);
nor U4074 (N_4074,N_3696,N_2869);
and U4075 (N_4075,N_3533,N_3085);
xor U4076 (N_4076,N_2611,N_3671);
xor U4077 (N_4077,N_3683,N_3247);
xor U4078 (N_4078,N_3442,N_2727);
nand U4079 (N_4079,N_3597,N_2880);
and U4080 (N_4080,N_3180,N_3699);
nor U4081 (N_4081,N_2973,N_2893);
or U4082 (N_4082,N_3351,N_2538);
and U4083 (N_4083,N_2870,N_3695);
and U4084 (N_4084,N_3121,N_3625);
nand U4085 (N_4085,N_3269,N_3547);
nand U4086 (N_4086,N_2864,N_2659);
or U4087 (N_4087,N_2885,N_2544);
nand U4088 (N_4088,N_2768,N_3022);
and U4089 (N_4089,N_3190,N_3255);
and U4090 (N_4090,N_3007,N_2628);
or U4091 (N_4091,N_3294,N_2529);
and U4092 (N_4092,N_2743,N_3457);
xor U4093 (N_4093,N_2971,N_3542);
xnor U4094 (N_4094,N_2540,N_3666);
xor U4095 (N_4095,N_3707,N_2952);
nand U4096 (N_4096,N_3392,N_3624);
nor U4097 (N_4097,N_3053,N_2997);
xor U4098 (N_4098,N_2938,N_2943);
xor U4099 (N_4099,N_3558,N_3661);
nand U4100 (N_4100,N_3382,N_2565);
nor U4101 (N_4101,N_3434,N_3038);
and U4102 (N_4102,N_3438,N_3067);
or U4103 (N_4103,N_3502,N_2818);
and U4104 (N_4104,N_2821,N_3160);
or U4105 (N_4105,N_3600,N_3567);
and U4106 (N_4106,N_3333,N_3326);
or U4107 (N_4107,N_2873,N_2641);
nor U4108 (N_4108,N_2889,N_3291);
nand U4109 (N_4109,N_2761,N_2705);
nand U4110 (N_4110,N_2892,N_3454);
nor U4111 (N_4111,N_3687,N_2584);
nor U4112 (N_4112,N_3439,N_2599);
nand U4113 (N_4113,N_3732,N_2564);
nand U4114 (N_4114,N_3744,N_2536);
xnor U4115 (N_4115,N_2613,N_3431);
nand U4116 (N_4116,N_3257,N_3528);
and U4117 (N_4117,N_3197,N_3078);
or U4118 (N_4118,N_3288,N_2990);
and U4119 (N_4119,N_2857,N_3512);
nand U4120 (N_4120,N_3238,N_3164);
nand U4121 (N_4121,N_3664,N_2987);
xor U4122 (N_4122,N_3578,N_3068);
xor U4123 (N_4123,N_2690,N_2874);
nand U4124 (N_4124,N_3106,N_2558);
and U4125 (N_4125,N_3050,N_3275);
nor U4126 (N_4126,N_3614,N_3014);
xnor U4127 (N_4127,N_2547,N_2843);
nor U4128 (N_4128,N_3102,N_2642);
and U4129 (N_4129,N_3745,N_3587);
or U4130 (N_4130,N_2585,N_3515);
or U4131 (N_4131,N_3560,N_3042);
xor U4132 (N_4132,N_3003,N_3224);
nor U4133 (N_4133,N_3416,N_3056);
xnor U4134 (N_4134,N_2569,N_3045);
nor U4135 (N_4135,N_2704,N_3383);
nand U4136 (N_4136,N_3739,N_3648);
nand U4137 (N_4137,N_3148,N_3672);
and U4138 (N_4138,N_2700,N_3103);
nand U4139 (N_4139,N_3384,N_3146);
nor U4140 (N_4140,N_2724,N_3040);
nand U4141 (N_4141,N_3295,N_3312);
xor U4142 (N_4142,N_3315,N_3048);
nand U4143 (N_4143,N_3507,N_2798);
and U4144 (N_4144,N_2996,N_3265);
nor U4145 (N_4145,N_2855,N_3286);
nor U4146 (N_4146,N_2667,N_2580);
and U4147 (N_4147,N_2610,N_3503);
and U4148 (N_4148,N_3485,N_2839);
nand U4149 (N_4149,N_2625,N_2551);
nand U4150 (N_4150,N_2570,N_2644);
nor U4151 (N_4151,N_2794,N_2949);
nor U4152 (N_4152,N_2980,N_3138);
nand U4153 (N_4153,N_3276,N_2955);
nor U4154 (N_4154,N_3287,N_2745);
and U4155 (N_4155,N_3676,N_3565);
nor U4156 (N_4156,N_2972,N_2888);
xnor U4157 (N_4157,N_3649,N_2772);
or U4158 (N_4158,N_2617,N_3230);
or U4159 (N_4159,N_2575,N_3385);
and U4160 (N_4160,N_3735,N_2533);
or U4161 (N_4161,N_3074,N_3402);
nor U4162 (N_4162,N_2507,N_2530);
or U4163 (N_4163,N_2931,N_2525);
and U4164 (N_4164,N_3451,N_2951);
nand U4165 (N_4165,N_2546,N_3685);
and U4166 (N_4166,N_3137,N_3370);
nand U4167 (N_4167,N_3313,N_3490);
nand U4168 (N_4168,N_3028,N_3235);
and U4169 (N_4169,N_2716,N_2730);
and U4170 (N_4170,N_3631,N_3132);
nand U4171 (N_4171,N_3151,N_3591);
nand U4172 (N_4172,N_2521,N_3418);
nand U4173 (N_4173,N_3156,N_3262);
and U4174 (N_4174,N_2830,N_2983);
nand U4175 (N_4175,N_2594,N_2665);
nor U4176 (N_4176,N_3709,N_3637);
nand U4177 (N_4177,N_3689,N_3271);
nand U4178 (N_4178,N_3073,N_3448);
and U4179 (N_4179,N_3272,N_3520);
or U4180 (N_4180,N_3178,N_3435);
nor U4181 (N_4181,N_3251,N_2681);
nor U4182 (N_4182,N_3577,N_3117);
or U4183 (N_4183,N_3720,N_3253);
nand U4184 (N_4184,N_3675,N_3358);
xor U4185 (N_4185,N_3432,N_3368);
or U4186 (N_4186,N_3256,N_2527);
nand U4187 (N_4187,N_3144,N_3519);
nor U4188 (N_4188,N_3443,N_2502);
nor U4189 (N_4189,N_2676,N_3498);
and U4190 (N_4190,N_3381,N_2576);
nor U4191 (N_4191,N_3129,N_2631);
and U4192 (N_4192,N_3150,N_2503);
and U4193 (N_4193,N_3212,N_3639);
and U4194 (N_4194,N_3613,N_3179);
xor U4195 (N_4195,N_3673,N_2753);
xor U4196 (N_4196,N_3742,N_3213);
xnor U4197 (N_4197,N_3239,N_2541);
nand U4198 (N_4198,N_2514,N_3497);
nor U4199 (N_4199,N_2930,N_2813);
and U4200 (N_4200,N_2590,N_3119);
or U4201 (N_4201,N_2925,N_3397);
and U4202 (N_4202,N_2915,N_2960);
or U4203 (N_4203,N_3189,N_2567);
xnor U4204 (N_4204,N_2684,N_2510);
nor U4205 (N_4205,N_2522,N_3141);
and U4206 (N_4206,N_2787,N_2959);
xnor U4207 (N_4207,N_3606,N_3586);
nor U4208 (N_4208,N_3492,N_2791);
or U4209 (N_4209,N_2560,N_2914);
and U4210 (N_4210,N_3517,N_3641);
nand U4211 (N_4211,N_3246,N_2995);
nor U4212 (N_4212,N_3331,N_2757);
nand U4213 (N_4213,N_3644,N_2634);
or U4214 (N_4214,N_2780,N_2956);
or U4215 (N_4215,N_2696,N_3159);
nor U4216 (N_4216,N_3527,N_2922);
xor U4217 (N_4217,N_2953,N_2988);
or U4218 (N_4218,N_3693,N_2809);
or U4219 (N_4219,N_3620,N_3216);
nand U4220 (N_4220,N_3460,N_2974);
and U4221 (N_4221,N_3686,N_2904);
and U4222 (N_4222,N_3716,N_2545);
xnor U4223 (N_4223,N_2766,N_3018);
and U4224 (N_4224,N_3167,N_2523);
nor U4225 (N_4225,N_3741,N_3521);
nor U4226 (N_4226,N_3270,N_3391);
xnor U4227 (N_4227,N_3329,N_2734);
or U4228 (N_4228,N_2837,N_3463);
or U4229 (N_4229,N_3746,N_2907);
xnor U4230 (N_4230,N_3339,N_2750);
nor U4231 (N_4231,N_2629,N_3363);
nor U4232 (N_4232,N_2589,N_2986);
nor U4233 (N_4233,N_2650,N_2793);
xnor U4234 (N_4234,N_3731,N_3107);
nand U4235 (N_4235,N_3185,N_2860);
or U4236 (N_4236,N_3133,N_3032);
xnor U4237 (N_4237,N_2660,N_3206);
xnor U4238 (N_4238,N_3128,N_2823);
and U4239 (N_4239,N_3688,N_2695);
nand U4240 (N_4240,N_3258,N_3455);
or U4241 (N_4241,N_3605,N_3596);
nand U4242 (N_4242,N_3069,N_3303);
and U4243 (N_4243,N_2800,N_3482);
xnor U4244 (N_4244,N_3566,N_3250);
xor U4245 (N_4245,N_2820,N_3549);
and U4246 (N_4246,N_2668,N_3096);
nor U4247 (N_4247,N_3267,N_3181);
and U4248 (N_4248,N_3634,N_3061);
nand U4249 (N_4249,N_3154,N_2591);
nand U4250 (N_4250,N_3697,N_2552);
or U4251 (N_4251,N_2762,N_2528);
nand U4252 (N_4252,N_3122,N_3388);
and U4253 (N_4253,N_3320,N_3684);
nor U4254 (N_4254,N_3002,N_3659);
or U4255 (N_4255,N_3231,N_3470);
nand U4256 (N_4256,N_3217,N_3109);
nand U4257 (N_4257,N_3095,N_3405);
nand U4258 (N_4258,N_3394,N_2919);
or U4259 (N_4259,N_3729,N_2950);
and U4260 (N_4260,N_3335,N_3651);
xnor U4261 (N_4261,N_2767,N_3293);
and U4262 (N_4262,N_2742,N_2583);
nor U4263 (N_4263,N_3529,N_2846);
nand U4264 (N_4264,N_3183,N_2751);
nor U4265 (N_4265,N_3211,N_3610);
nand U4266 (N_4266,N_2666,N_3579);
and U4267 (N_4267,N_3574,N_3236);
xor U4268 (N_4268,N_2687,N_3356);
or U4269 (N_4269,N_3551,N_2847);
nor U4270 (N_4270,N_2871,N_3724);
nand U4271 (N_4271,N_3513,N_2662);
or U4272 (N_4272,N_3306,N_2685);
and U4273 (N_4273,N_2509,N_3638);
nor U4274 (N_4274,N_2664,N_3389);
xor U4275 (N_4275,N_3535,N_3647);
or U4276 (N_4276,N_3242,N_3177);
and U4277 (N_4277,N_3602,N_2918);
nor U4278 (N_4278,N_2715,N_3510);
or U4279 (N_4279,N_2877,N_2758);
nor U4280 (N_4280,N_3296,N_3657);
nand U4281 (N_4281,N_3561,N_3617);
xnor U4282 (N_4282,N_2638,N_3021);
nor U4283 (N_4283,N_3100,N_3327);
xnor U4284 (N_4284,N_3273,N_3260);
or U4285 (N_4285,N_2954,N_2729);
and U4286 (N_4286,N_2609,N_3585);
nor U4287 (N_4287,N_2978,N_3266);
nand U4288 (N_4288,N_3505,N_2827);
xnor U4289 (N_4289,N_2933,N_3347);
and U4290 (N_4290,N_3595,N_3058);
or U4291 (N_4291,N_2539,N_3459);
xnor U4292 (N_4292,N_3733,N_3023);
nor U4293 (N_4293,N_2519,N_3702);
nand U4294 (N_4294,N_2616,N_3654);
or U4295 (N_4295,N_3691,N_3440);
xor U4296 (N_4296,N_3297,N_3430);
and U4297 (N_4297,N_2554,N_3044);
or U4298 (N_4298,N_3279,N_3033);
nand U4299 (N_4299,N_3495,N_3537);
nor U4300 (N_4300,N_3590,N_3089);
and U4301 (N_4301,N_3557,N_3518);
nand U4302 (N_4302,N_3349,N_3136);
nand U4303 (N_4303,N_2911,N_2572);
or U4304 (N_4304,N_3364,N_2713);
nor U4305 (N_4305,N_2908,N_3543);
or U4306 (N_4306,N_3209,N_3278);
nand U4307 (N_4307,N_2776,N_2859);
nor U4308 (N_4308,N_2784,N_3243);
xnor U4309 (N_4309,N_3322,N_2779);
nand U4310 (N_4310,N_3196,N_2723);
or U4311 (N_4311,N_3232,N_3404);
nor U4312 (N_4312,N_3341,N_3698);
nor U4313 (N_4313,N_2671,N_3165);
xnor U4314 (N_4314,N_3282,N_2720);
xnor U4315 (N_4315,N_3099,N_3622);
or U4316 (N_4316,N_2814,N_2632);
nor U4317 (N_4317,N_3419,N_3559);
or U4318 (N_4318,N_2725,N_3317);
nand U4319 (N_4319,N_3188,N_3314);
xor U4320 (N_4320,N_2561,N_3568);
xor U4321 (N_4321,N_3708,N_2966);
and U4322 (N_4322,N_2612,N_2559);
and U4323 (N_4323,N_3029,N_2574);
and U4324 (N_4324,N_2707,N_3710);
or U4325 (N_4325,N_3478,N_2764);
or U4326 (N_4326,N_3522,N_2754);
or U4327 (N_4327,N_3628,N_3346);
and U4328 (N_4328,N_3713,N_2868);
nor U4329 (N_4329,N_2568,N_3734);
and U4330 (N_4330,N_3640,N_3532);
nor U4331 (N_4331,N_2985,N_3283);
nand U4332 (N_4332,N_2703,N_2722);
and U4333 (N_4333,N_2875,N_2535);
nand U4334 (N_4334,N_2686,N_2731);
nor U4335 (N_4335,N_2979,N_2637);
nor U4336 (N_4336,N_2947,N_2740);
and U4337 (N_4337,N_2917,N_3277);
nand U4338 (N_4338,N_3001,N_3218);
and U4339 (N_4339,N_2899,N_3024);
xor U4340 (N_4340,N_2825,N_3484);
nor U4341 (N_4341,N_2563,N_2579);
nor U4342 (N_4342,N_2593,N_3444);
xnor U4343 (N_4343,N_3643,N_3441);
xnor U4344 (N_4344,N_3125,N_3310);
nor U4345 (N_4345,N_2607,N_3155);
nand U4346 (N_4346,N_3523,N_3323);
xnor U4347 (N_4347,N_3332,N_3281);
xor U4348 (N_4348,N_3065,N_2865);
xnor U4349 (N_4349,N_2562,N_3374);
or U4350 (N_4350,N_3469,N_2802);
and U4351 (N_4351,N_3429,N_3019);
xnor U4352 (N_4352,N_3483,N_3321);
nand U4353 (N_4353,N_3692,N_3052);
and U4354 (N_4354,N_3727,N_2505);
and U4355 (N_4355,N_3538,N_2862);
xor U4356 (N_4356,N_3261,N_3481);
or U4357 (N_4357,N_3705,N_3499);
or U4358 (N_4358,N_2663,N_3371);
nor U4359 (N_4359,N_3285,N_2778);
and U4360 (N_4360,N_3169,N_3633);
or U4361 (N_4361,N_3173,N_2897);
xor U4362 (N_4362,N_2697,N_3545);
and U4363 (N_4363,N_3682,N_2738);
and U4364 (N_4364,N_3736,N_3357);
or U4365 (N_4365,N_3162,N_3700);
xor U4366 (N_4366,N_3153,N_3354);
nor U4367 (N_4367,N_3116,N_2524);
and U4368 (N_4368,N_3714,N_3629);
nor U4369 (N_4369,N_3104,N_2677);
or U4370 (N_4370,N_3531,N_3428);
and U4371 (N_4371,N_3009,N_2944);
nand U4372 (N_4372,N_3097,N_3417);
and U4373 (N_4373,N_2894,N_2657);
or U4374 (N_4374,N_2887,N_2890);
xnor U4375 (N_4375,N_3483,N_2609);
and U4376 (N_4376,N_3016,N_3020);
nor U4377 (N_4377,N_3116,N_2568);
xor U4378 (N_4378,N_2716,N_3684);
and U4379 (N_4379,N_3286,N_2583);
xnor U4380 (N_4380,N_3644,N_3332);
nor U4381 (N_4381,N_2951,N_3679);
nor U4382 (N_4382,N_2638,N_2800);
xor U4383 (N_4383,N_3114,N_3367);
nand U4384 (N_4384,N_2996,N_2527);
xnor U4385 (N_4385,N_3603,N_2645);
nand U4386 (N_4386,N_3615,N_2741);
nor U4387 (N_4387,N_3736,N_2542);
xor U4388 (N_4388,N_2605,N_2998);
xnor U4389 (N_4389,N_3572,N_2897);
nand U4390 (N_4390,N_3099,N_3669);
nand U4391 (N_4391,N_3541,N_3041);
nor U4392 (N_4392,N_3383,N_3485);
or U4393 (N_4393,N_2949,N_3565);
xnor U4394 (N_4394,N_3730,N_2567);
or U4395 (N_4395,N_3698,N_3390);
or U4396 (N_4396,N_3552,N_2662);
nand U4397 (N_4397,N_3173,N_3340);
nand U4398 (N_4398,N_3472,N_3522);
xor U4399 (N_4399,N_3696,N_3242);
nor U4400 (N_4400,N_2615,N_3336);
and U4401 (N_4401,N_3169,N_3564);
xnor U4402 (N_4402,N_2881,N_3701);
nor U4403 (N_4403,N_2860,N_3200);
nand U4404 (N_4404,N_3646,N_3649);
nand U4405 (N_4405,N_2844,N_3391);
and U4406 (N_4406,N_3257,N_2741);
nand U4407 (N_4407,N_2717,N_3393);
nor U4408 (N_4408,N_3300,N_3150);
xor U4409 (N_4409,N_3399,N_3394);
nor U4410 (N_4410,N_3719,N_3241);
and U4411 (N_4411,N_2800,N_2801);
and U4412 (N_4412,N_2584,N_2995);
nor U4413 (N_4413,N_3631,N_2751);
and U4414 (N_4414,N_3379,N_2504);
nand U4415 (N_4415,N_3639,N_2593);
nor U4416 (N_4416,N_3016,N_3514);
nand U4417 (N_4417,N_3289,N_3587);
xnor U4418 (N_4418,N_3333,N_3299);
xor U4419 (N_4419,N_2751,N_3060);
nand U4420 (N_4420,N_3333,N_3108);
xnor U4421 (N_4421,N_3028,N_3166);
nor U4422 (N_4422,N_2685,N_2584);
xor U4423 (N_4423,N_3418,N_3269);
nand U4424 (N_4424,N_3527,N_2933);
and U4425 (N_4425,N_2891,N_3136);
xor U4426 (N_4426,N_3500,N_2683);
nor U4427 (N_4427,N_3179,N_3181);
and U4428 (N_4428,N_3181,N_3244);
or U4429 (N_4429,N_2585,N_3204);
nor U4430 (N_4430,N_2883,N_3089);
nor U4431 (N_4431,N_3332,N_3082);
xnor U4432 (N_4432,N_2565,N_3605);
and U4433 (N_4433,N_2556,N_3170);
or U4434 (N_4434,N_3132,N_2796);
xor U4435 (N_4435,N_3579,N_3165);
or U4436 (N_4436,N_2518,N_2946);
nand U4437 (N_4437,N_3704,N_3709);
xor U4438 (N_4438,N_3259,N_2733);
nand U4439 (N_4439,N_2623,N_3452);
nor U4440 (N_4440,N_2718,N_3621);
nand U4441 (N_4441,N_2543,N_3485);
or U4442 (N_4442,N_2604,N_2605);
nor U4443 (N_4443,N_2907,N_3284);
or U4444 (N_4444,N_3450,N_3367);
nand U4445 (N_4445,N_3231,N_3304);
xnor U4446 (N_4446,N_3236,N_2969);
nor U4447 (N_4447,N_2666,N_3663);
nand U4448 (N_4448,N_2584,N_3240);
or U4449 (N_4449,N_3312,N_3267);
xnor U4450 (N_4450,N_3661,N_3160);
nor U4451 (N_4451,N_2777,N_3518);
or U4452 (N_4452,N_2590,N_2607);
or U4453 (N_4453,N_2955,N_3341);
and U4454 (N_4454,N_3611,N_3190);
nor U4455 (N_4455,N_2996,N_3196);
nand U4456 (N_4456,N_2686,N_3691);
and U4457 (N_4457,N_3465,N_3683);
xor U4458 (N_4458,N_3330,N_3725);
xor U4459 (N_4459,N_3415,N_3339);
xnor U4460 (N_4460,N_2881,N_3505);
or U4461 (N_4461,N_2986,N_3356);
xnor U4462 (N_4462,N_3058,N_2535);
and U4463 (N_4463,N_3229,N_2727);
or U4464 (N_4464,N_2894,N_2622);
xnor U4465 (N_4465,N_3716,N_3436);
xnor U4466 (N_4466,N_2631,N_2573);
or U4467 (N_4467,N_3079,N_2767);
and U4468 (N_4468,N_3495,N_3619);
nand U4469 (N_4469,N_3292,N_3195);
nor U4470 (N_4470,N_2744,N_3243);
or U4471 (N_4471,N_3179,N_3048);
and U4472 (N_4472,N_3155,N_3084);
xnor U4473 (N_4473,N_3199,N_3612);
and U4474 (N_4474,N_3416,N_2744);
and U4475 (N_4475,N_3213,N_2548);
and U4476 (N_4476,N_2757,N_3430);
xor U4477 (N_4477,N_2568,N_2775);
or U4478 (N_4478,N_2898,N_3021);
or U4479 (N_4479,N_2693,N_3647);
or U4480 (N_4480,N_3504,N_3422);
xnor U4481 (N_4481,N_3296,N_3424);
nor U4482 (N_4482,N_3030,N_3335);
or U4483 (N_4483,N_3108,N_2515);
nand U4484 (N_4484,N_3101,N_2741);
or U4485 (N_4485,N_3713,N_2903);
xor U4486 (N_4486,N_3138,N_2860);
and U4487 (N_4487,N_2507,N_3420);
nor U4488 (N_4488,N_2662,N_2899);
xnor U4489 (N_4489,N_2922,N_3199);
and U4490 (N_4490,N_3417,N_2657);
nand U4491 (N_4491,N_3345,N_3318);
nor U4492 (N_4492,N_2682,N_2618);
or U4493 (N_4493,N_3478,N_3577);
nand U4494 (N_4494,N_3248,N_3731);
or U4495 (N_4495,N_3012,N_3196);
and U4496 (N_4496,N_3079,N_3158);
or U4497 (N_4497,N_3323,N_2720);
or U4498 (N_4498,N_3481,N_3404);
or U4499 (N_4499,N_3104,N_3352);
and U4500 (N_4500,N_3248,N_3524);
nand U4501 (N_4501,N_3181,N_2863);
nand U4502 (N_4502,N_2740,N_3676);
nor U4503 (N_4503,N_2870,N_3237);
nor U4504 (N_4504,N_2547,N_3630);
and U4505 (N_4505,N_2870,N_3103);
nand U4506 (N_4506,N_3707,N_3610);
nor U4507 (N_4507,N_3698,N_2687);
nand U4508 (N_4508,N_3465,N_3411);
xnor U4509 (N_4509,N_3028,N_3310);
and U4510 (N_4510,N_3431,N_2720);
and U4511 (N_4511,N_2550,N_2867);
or U4512 (N_4512,N_2718,N_3006);
nor U4513 (N_4513,N_3004,N_2977);
nand U4514 (N_4514,N_3309,N_3648);
nor U4515 (N_4515,N_3068,N_2679);
nor U4516 (N_4516,N_3543,N_2965);
xor U4517 (N_4517,N_3332,N_3155);
and U4518 (N_4518,N_3699,N_3134);
and U4519 (N_4519,N_3307,N_3627);
xor U4520 (N_4520,N_3666,N_2771);
and U4521 (N_4521,N_3669,N_2687);
xnor U4522 (N_4522,N_3480,N_2562);
nand U4523 (N_4523,N_3385,N_3429);
nand U4524 (N_4524,N_3564,N_3336);
nor U4525 (N_4525,N_3228,N_2985);
and U4526 (N_4526,N_3010,N_2923);
xnor U4527 (N_4527,N_3336,N_3152);
xnor U4528 (N_4528,N_3444,N_3294);
and U4529 (N_4529,N_3708,N_3497);
nand U4530 (N_4530,N_3150,N_3295);
xor U4531 (N_4531,N_2733,N_3583);
nand U4532 (N_4532,N_3177,N_2997);
xnor U4533 (N_4533,N_3211,N_3262);
xor U4534 (N_4534,N_2926,N_2511);
nand U4535 (N_4535,N_2723,N_3599);
or U4536 (N_4536,N_2700,N_3730);
or U4537 (N_4537,N_3248,N_3643);
and U4538 (N_4538,N_3714,N_3133);
or U4539 (N_4539,N_2606,N_2541);
and U4540 (N_4540,N_2558,N_3022);
and U4541 (N_4541,N_3141,N_3014);
nand U4542 (N_4542,N_3087,N_3328);
xor U4543 (N_4543,N_3063,N_3570);
or U4544 (N_4544,N_2898,N_3168);
nor U4545 (N_4545,N_3500,N_3270);
xnor U4546 (N_4546,N_3306,N_2859);
nand U4547 (N_4547,N_3080,N_2929);
and U4548 (N_4548,N_2607,N_3235);
or U4549 (N_4549,N_2955,N_3481);
and U4550 (N_4550,N_3176,N_3322);
and U4551 (N_4551,N_2532,N_2667);
xnor U4552 (N_4552,N_3696,N_2827);
nand U4553 (N_4553,N_3488,N_2672);
nor U4554 (N_4554,N_2871,N_3243);
and U4555 (N_4555,N_3015,N_3610);
nor U4556 (N_4556,N_3148,N_3135);
xnor U4557 (N_4557,N_3190,N_2558);
and U4558 (N_4558,N_3514,N_3367);
xor U4559 (N_4559,N_3327,N_3074);
and U4560 (N_4560,N_2756,N_2933);
nor U4561 (N_4561,N_3158,N_3265);
nor U4562 (N_4562,N_2726,N_2923);
nand U4563 (N_4563,N_3538,N_2978);
nor U4564 (N_4564,N_2792,N_3711);
nand U4565 (N_4565,N_2926,N_2647);
nand U4566 (N_4566,N_3215,N_2548);
xor U4567 (N_4567,N_2831,N_3245);
and U4568 (N_4568,N_2787,N_3715);
and U4569 (N_4569,N_2709,N_2956);
or U4570 (N_4570,N_3693,N_3748);
nor U4571 (N_4571,N_3327,N_3008);
xor U4572 (N_4572,N_3249,N_3257);
nor U4573 (N_4573,N_2933,N_3122);
and U4574 (N_4574,N_3565,N_2639);
nor U4575 (N_4575,N_2695,N_2597);
nor U4576 (N_4576,N_2576,N_2909);
nand U4577 (N_4577,N_3104,N_2920);
nor U4578 (N_4578,N_3533,N_2990);
nor U4579 (N_4579,N_2845,N_2680);
and U4580 (N_4580,N_3304,N_3356);
and U4581 (N_4581,N_3657,N_3142);
or U4582 (N_4582,N_3087,N_2889);
and U4583 (N_4583,N_2927,N_2551);
or U4584 (N_4584,N_2926,N_3375);
nor U4585 (N_4585,N_3481,N_2575);
and U4586 (N_4586,N_3196,N_3218);
or U4587 (N_4587,N_3154,N_2874);
nand U4588 (N_4588,N_2614,N_3381);
nand U4589 (N_4589,N_2616,N_2677);
nor U4590 (N_4590,N_3377,N_2964);
or U4591 (N_4591,N_3324,N_2803);
xnor U4592 (N_4592,N_3399,N_3544);
xor U4593 (N_4593,N_3319,N_3148);
xnor U4594 (N_4594,N_3168,N_3015);
nor U4595 (N_4595,N_2949,N_3556);
xnor U4596 (N_4596,N_3567,N_3250);
nand U4597 (N_4597,N_3663,N_3262);
xnor U4598 (N_4598,N_2621,N_2819);
xnor U4599 (N_4599,N_3345,N_3608);
and U4600 (N_4600,N_2785,N_3327);
or U4601 (N_4601,N_2968,N_3506);
or U4602 (N_4602,N_2966,N_2771);
or U4603 (N_4603,N_2693,N_3285);
nor U4604 (N_4604,N_2796,N_3412);
xnor U4605 (N_4605,N_3525,N_2802);
xor U4606 (N_4606,N_2630,N_3200);
nand U4607 (N_4607,N_2755,N_3084);
xor U4608 (N_4608,N_2849,N_2922);
and U4609 (N_4609,N_3540,N_2802);
and U4610 (N_4610,N_3681,N_3380);
and U4611 (N_4611,N_3099,N_2531);
or U4612 (N_4612,N_2905,N_2564);
nor U4613 (N_4613,N_2816,N_3246);
nor U4614 (N_4614,N_2954,N_3373);
xor U4615 (N_4615,N_2764,N_2731);
or U4616 (N_4616,N_2822,N_2592);
or U4617 (N_4617,N_2846,N_3339);
nor U4618 (N_4618,N_3226,N_2740);
or U4619 (N_4619,N_3142,N_3170);
nor U4620 (N_4620,N_3567,N_3615);
xnor U4621 (N_4621,N_2912,N_2772);
or U4622 (N_4622,N_3197,N_2500);
nand U4623 (N_4623,N_3221,N_3689);
xor U4624 (N_4624,N_3018,N_3561);
and U4625 (N_4625,N_3621,N_2751);
and U4626 (N_4626,N_3690,N_2798);
or U4627 (N_4627,N_3748,N_2757);
nor U4628 (N_4628,N_3276,N_3313);
nand U4629 (N_4629,N_3244,N_3121);
or U4630 (N_4630,N_3334,N_3681);
or U4631 (N_4631,N_3583,N_3542);
or U4632 (N_4632,N_3547,N_2823);
or U4633 (N_4633,N_2677,N_3089);
nand U4634 (N_4634,N_3617,N_2624);
or U4635 (N_4635,N_3492,N_3235);
xnor U4636 (N_4636,N_2598,N_3539);
nand U4637 (N_4637,N_3736,N_3356);
xor U4638 (N_4638,N_2722,N_3055);
or U4639 (N_4639,N_2752,N_3078);
xor U4640 (N_4640,N_3332,N_2773);
nand U4641 (N_4641,N_3240,N_2814);
nor U4642 (N_4642,N_3070,N_3028);
nor U4643 (N_4643,N_3103,N_3087);
nand U4644 (N_4644,N_3352,N_3603);
or U4645 (N_4645,N_3283,N_3110);
nor U4646 (N_4646,N_3698,N_3123);
or U4647 (N_4647,N_3065,N_3289);
nand U4648 (N_4648,N_3047,N_3562);
xnor U4649 (N_4649,N_2976,N_3728);
or U4650 (N_4650,N_3608,N_3213);
nor U4651 (N_4651,N_3300,N_3544);
and U4652 (N_4652,N_2899,N_3623);
and U4653 (N_4653,N_3625,N_3485);
or U4654 (N_4654,N_2559,N_3309);
or U4655 (N_4655,N_3657,N_2534);
and U4656 (N_4656,N_2742,N_2886);
nand U4657 (N_4657,N_3539,N_2974);
and U4658 (N_4658,N_3246,N_3586);
and U4659 (N_4659,N_3658,N_2981);
nand U4660 (N_4660,N_3017,N_2775);
nand U4661 (N_4661,N_2921,N_3215);
nor U4662 (N_4662,N_3488,N_3055);
xor U4663 (N_4663,N_3652,N_2692);
nand U4664 (N_4664,N_2979,N_3030);
xnor U4665 (N_4665,N_3402,N_2956);
nand U4666 (N_4666,N_2548,N_2592);
xor U4667 (N_4667,N_3176,N_2839);
and U4668 (N_4668,N_3682,N_2928);
nand U4669 (N_4669,N_3023,N_3028);
or U4670 (N_4670,N_3546,N_2869);
xnor U4671 (N_4671,N_2864,N_3642);
and U4672 (N_4672,N_3205,N_2554);
nand U4673 (N_4673,N_2968,N_3467);
and U4674 (N_4674,N_2954,N_2990);
or U4675 (N_4675,N_2892,N_2554);
xnor U4676 (N_4676,N_3158,N_2760);
and U4677 (N_4677,N_2926,N_2814);
nand U4678 (N_4678,N_2818,N_3363);
nor U4679 (N_4679,N_2550,N_2595);
nor U4680 (N_4680,N_2713,N_3018);
or U4681 (N_4681,N_2746,N_2657);
or U4682 (N_4682,N_2848,N_3500);
or U4683 (N_4683,N_3092,N_3000);
and U4684 (N_4684,N_2835,N_2509);
nand U4685 (N_4685,N_3494,N_2979);
nand U4686 (N_4686,N_3484,N_3431);
and U4687 (N_4687,N_2658,N_3718);
nand U4688 (N_4688,N_3429,N_2804);
nand U4689 (N_4689,N_3382,N_2742);
xor U4690 (N_4690,N_3276,N_2906);
xor U4691 (N_4691,N_3200,N_3703);
xnor U4692 (N_4692,N_2548,N_3720);
xnor U4693 (N_4693,N_2702,N_2848);
nor U4694 (N_4694,N_2594,N_2954);
nand U4695 (N_4695,N_2528,N_2744);
and U4696 (N_4696,N_3055,N_3515);
nand U4697 (N_4697,N_3445,N_2902);
or U4698 (N_4698,N_2871,N_2684);
or U4699 (N_4699,N_3218,N_2872);
xor U4700 (N_4700,N_2768,N_3107);
xor U4701 (N_4701,N_3279,N_3359);
nor U4702 (N_4702,N_3460,N_2810);
and U4703 (N_4703,N_3114,N_3282);
xor U4704 (N_4704,N_2801,N_2985);
or U4705 (N_4705,N_3679,N_2718);
xnor U4706 (N_4706,N_3566,N_2667);
xor U4707 (N_4707,N_3379,N_2913);
and U4708 (N_4708,N_2868,N_2748);
or U4709 (N_4709,N_2970,N_2746);
and U4710 (N_4710,N_2968,N_3731);
nor U4711 (N_4711,N_3678,N_3546);
or U4712 (N_4712,N_3224,N_3523);
nand U4713 (N_4713,N_3408,N_3027);
and U4714 (N_4714,N_3619,N_3009);
and U4715 (N_4715,N_3715,N_2740);
nand U4716 (N_4716,N_3403,N_3029);
or U4717 (N_4717,N_2739,N_3432);
xor U4718 (N_4718,N_3416,N_2635);
nor U4719 (N_4719,N_3600,N_2638);
nand U4720 (N_4720,N_2926,N_3298);
and U4721 (N_4721,N_2853,N_3326);
nor U4722 (N_4722,N_2877,N_3419);
and U4723 (N_4723,N_3537,N_2852);
or U4724 (N_4724,N_3550,N_3351);
nand U4725 (N_4725,N_2792,N_2966);
xor U4726 (N_4726,N_2876,N_2811);
and U4727 (N_4727,N_2663,N_3451);
nand U4728 (N_4728,N_2790,N_2957);
nand U4729 (N_4729,N_2931,N_2734);
nor U4730 (N_4730,N_3145,N_2887);
or U4731 (N_4731,N_3105,N_2991);
and U4732 (N_4732,N_2811,N_3228);
or U4733 (N_4733,N_3398,N_3700);
or U4734 (N_4734,N_3203,N_3610);
nand U4735 (N_4735,N_2588,N_3528);
and U4736 (N_4736,N_3508,N_2689);
and U4737 (N_4737,N_2808,N_2655);
xnor U4738 (N_4738,N_3281,N_3606);
xnor U4739 (N_4739,N_3171,N_2622);
xor U4740 (N_4740,N_2672,N_3710);
nand U4741 (N_4741,N_2534,N_3524);
xor U4742 (N_4742,N_3406,N_3076);
xor U4743 (N_4743,N_3358,N_3105);
and U4744 (N_4744,N_2506,N_3681);
xnor U4745 (N_4745,N_3581,N_3449);
nand U4746 (N_4746,N_3000,N_2910);
or U4747 (N_4747,N_2953,N_2923);
xor U4748 (N_4748,N_2856,N_3292);
or U4749 (N_4749,N_3323,N_2669);
and U4750 (N_4750,N_2539,N_2534);
nand U4751 (N_4751,N_2542,N_2962);
or U4752 (N_4752,N_3123,N_3070);
nand U4753 (N_4753,N_2568,N_3356);
nand U4754 (N_4754,N_3444,N_3011);
xnor U4755 (N_4755,N_3502,N_3673);
nand U4756 (N_4756,N_3480,N_2635);
nor U4757 (N_4757,N_3644,N_2685);
nor U4758 (N_4758,N_2769,N_3679);
and U4759 (N_4759,N_2854,N_3654);
xor U4760 (N_4760,N_3304,N_2675);
and U4761 (N_4761,N_3051,N_2748);
or U4762 (N_4762,N_3184,N_3223);
or U4763 (N_4763,N_3509,N_3332);
and U4764 (N_4764,N_2805,N_3363);
nor U4765 (N_4765,N_3044,N_2862);
or U4766 (N_4766,N_3345,N_2706);
nand U4767 (N_4767,N_3484,N_3553);
nor U4768 (N_4768,N_3591,N_2891);
nor U4769 (N_4769,N_2692,N_3574);
xor U4770 (N_4770,N_2592,N_3573);
and U4771 (N_4771,N_3057,N_3742);
or U4772 (N_4772,N_3728,N_3508);
nand U4773 (N_4773,N_2666,N_3587);
and U4774 (N_4774,N_3159,N_3252);
nand U4775 (N_4775,N_2912,N_3712);
and U4776 (N_4776,N_2674,N_3245);
nor U4777 (N_4777,N_3400,N_3472);
or U4778 (N_4778,N_2671,N_2674);
and U4779 (N_4779,N_3484,N_2774);
or U4780 (N_4780,N_3310,N_2579);
xnor U4781 (N_4781,N_3700,N_3432);
nor U4782 (N_4782,N_3460,N_2921);
nor U4783 (N_4783,N_3624,N_2957);
and U4784 (N_4784,N_3352,N_2740);
nor U4785 (N_4785,N_3452,N_3035);
nand U4786 (N_4786,N_2761,N_3284);
nor U4787 (N_4787,N_3671,N_3481);
or U4788 (N_4788,N_3634,N_3323);
and U4789 (N_4789,N_3612,N_3350);
xnor U4790 (N_4790,N_2773,N_2699);
xor U4791 (N_4791,N_3025,N_3628);
and U4792 (N_4792,N_3308,N_3050);
or U4793 (N_4793,N_3341,N_2844);
nor U4794 (N_4794,N_2676,N_3334);
and U4795 (N_4795,N_3327,N_3389);
nor U4796 (N_4796,N_2633,N_2648);
nand U4797 (N_4797,N_2848,N_2735);
and U4798 (N_4798,N_2857,N_3319);
xnor U4799 (N_4799,N_2893,N_3632);
nand U4800 (N_4800,N_2734,N_2872);
nand U4801 (N_4801,N_2793,N_3550);
nand U4802 (N_4802,N_2689,N_3264);
or U4803 (N_4803,N_2748,N_2546);
nor U4804 (N_4804,N_3509,N_2905);
nand U4805 (N_4805,N_2562,N_2720);
and U4806 (N_4806,N_2721,N_2549);
nand U4807 (N_4807,N_3072,N_3373);
nor U4808 (N_4808,N_2978,N_2589);
nand U4809 (N_4809,N_3042,N_2931);
or U4810 (N_4810,N_3136,N_2902);
and U4811 (N_4811,N_3200,N_3636);
xnor U4812 (N_4812,N_3525,N_3158);
and U4813 (N_4813,N_3383,N_2606);
xor U4814 (N_4814,N_3500,N_2588);
xor U4815 (N_4815,N_3240,N_3650);
xnor U4816 (N_4816,N_2515,N_2928);
or U4817 (N_4817,N_3357,N_2570);
nor U4818 (N_4818,N_3407,N_3288);
nand U4819 (N_4819,N_3514,N_3378);
or U4820 (N_4820,N_3309,N_3611);
and U4821 (N_4821,N_3598,N_3027);
nand U4822 (N_4822,N_2915,N_2914);
or U4823 (N_4823,N_3400,N_3471);
and U4824 (N_4824,N_2941,N_2880);
and U4825 (N_4825,N_3065,N_2629);
nor U4826 (N_4826,N_3709,N_2822);
nand U4827 (N_4827,N_3532,N_3572);
nand U4828 (N_4828,N_3529,N_2706);
or U4829 (N_4829,N_3333,N_2688);
nand U4830 (N_4830,N_2523,N_3016);
nand U4831 (N_4831,N_3098,N_3025);
xor U4832 (N_4832,N_3515,N_3080);
nand U4833 (N_4833,N_3388,N_3292);
nand U4834 (N_4834,N_3344,N_3239);
xor U4835 (N_4835,N_3637,N_2954);
nor U4836 (N_4836,N_2514,N_3089);
xnor U4837 (N_4837,N_3691,N_3369);
and U4838 (N_4838,N_2656,N_3521);
nand U4839 (N_4839,N_3137,N_3344);
nor U4840 (N_4840,N_3073,N_3236);
nand U4841 (N_4841,N_3683,N_3153);
nand U4842 (N_4842,N_2672,N_3697);
or U4843 (N_4843,N_2838,N_2630);
xor U4844 (N_4844,N_3560,N_3574);
or U4845 (N_4845,N_3601,N_3652);
nor U4846 (N_4846,N_3433,N_2546);
and U4847 (N_4847,N_2788,N_2566);
or U4848 (N_4848,N_2516,N_3415);
xnor U4849 (N_4849,N_3144,N_3304);
nor U4850 (N_4850,N_2593,N_3044);
nand U4851 (N_4851,N_3517,N_3185);
xor U4852 (N_4852,N_3546,N_3668);
or U4853 (N_4853,N_2612,N_2654);
xor U4854 (N_4854,N_2922,N_3233);
and U4855 (N_4855,N_3362,N_3358);
and U4856 (N_4856,N_3655,N_3249);
and U4857 (N_4857,N_3358,N_3258);
nor U4858 (N_4858,N_3035,N_2990);
nor U4859 (N_4859,N_3067,N_3599);
xor U4860 (N_4860,N_2614,N_3596);
xnor U4861 (N_4861,N_3457,N_3013);
nand U4862 (N_4862,N_3470,N_2503);
nand U4863 (N_4863,N_2696,N_2592);
or U4864 (N_4864,N_3408,N_3237);
and U4865 (N_4865,N_3020,N_3494);
or U4866 (N_4866,N_3636,N_3363);
or U4867 (N_4867,N_3728,N_2521);
and U4868 (N_4868,N_2722,N_3374);
nor U4869 (N_4869,N_3157,N_2725);
and U4870 (N_4870,N_2996,N_2995);
nand U4871 (N_4871,N_2992,N_2681);
nand U4872 (N_4872,N_3427,N_2548);
or U4873 (N_4873,N_3049,N_3625);
or U4874 (N_4874,N_3265,N_2625);
or U4875 (N_4875,N_2724,N_3412);
or U4876 (N_4876,N_2876,N_3370);
and U4877 (N_4877,N_2967,N_2940);
and U4878 (N_4878,N_3639,N_3555);
nor U4879 (N_4879,N_2865,N_3728);
and U4880 (N_4880,N_3687,N_3250);
nand U4881 (N_4881,N_3239,N_3685);
nand U4882 (N_4882,N_3265,N_2557);
and U4883 (N_4883,N_3448,N_2794);
nand U4884 (N_4884,N_3661,N_2555);
nor U4885 (N_4885,N_3422,N_3627);
and U4886 (N_4886,N_3353,N_2502);
or U4887 (N_4887,N_3285,N_3162);
and U4888 (N_4888,N_3719,N_3075);
and U4889 (N_4889,N_3735,N_2980);
xor U4890 (N_4890,N_3220,N_2742);
and U4891 (N_4891,N_3694,N_2975);
nand U4892 (N_4892,N_2947,N_3352);
nand U4893 (N_4893,N_2517,N_3526);
nor U4894 (N_4894,N_3679,N_2686);
xnor U4895 (N_4895,N_3021,N_3723);
nand U4896 (N_4896,N_2774,N_3513);
nor U4897 (N_4897,N_3579,N_3095);
xor U4898 (N_4898,N_3018,N_3486);
nand U4899 (N_4899,N_3737,N_3369);
or U4900 (N_4900,N_2859,N_3385);
nor U4901 (N_4901,N_2706,N_3110);
or U4902 (N_4902,N_3075,N_2972);
and U4903 (N_4903,N_2863,N_3072);
or U4904 (N_4904,N_3311,N_2583);
xnor U4905 (N_4905,N_3483,N_2709);
nand U4906 (N_4906,N_2576,N_3472);
and U4907 (N_4907,N_3021,N_3439);
or U4908 (N_4908,N_3166,N_3329);
and U4909 (N_4909,N_3671,N_2541);
nor U4910 (N_4910,N_3624,N_2514);
xnor U4911 (N_4911,N_3457,N_2760);
nand U4912 (N_4912,N_3165,N_3528);
nand U4913 (N_4913,N_3226,N_3526);
nand U4914 (N_4914,N_3291,N_3307);
nand U4915 (N_4915,N_2806,N_2586);
nor U4916 (N_4916,N_3049,N_3464);
xnor U4917 (N_4917,N_3235,N_3742);
nor U4918 (N_4918,N_3176,N_3414);
nand U4919 (N_4919,N_3504,N_3666);
xnor U4920 (N_4920,N_3079,N_2678);
nor U4921 (N_4921,N_2598,N_2697);
nand U4922 (N_4922,N_3144,N_3424);
xnor U4923 (N_4923,N_2930,N_2934);
or U4924 (N_4924,N_3547,N_3147);
nor U4925 (N_4925,N_3485,N_3134);
and U4926 (N_4926,N_2587,N_3163);
xor U4927 (N_4927,N_3084,N_3131);
and U4928 (N_4928,N_3251,N_2821);
and U4929 (N_4929,N_3476,N_3410);
xnor U4930 (N_4930,N_2513,N_2781);
and U4931 (N_4931,N_3737,N_3576);
nand U4932 (N_4932,N_3331,N_2720);
nand U4933 (N_4933,N_3625,N_2936);
nand U4934 (N_4934,N_2773,N_3263);
nor U4935 (N_4935,N_3058,N_2517);
nor U4936 (N_4936,N_3388,N_3082);
nand U4937 (N_4937,N_3290,N_3042);
or U4938 (N_4938,N_3474,N_3120);
nand U4939 (N_4939,N_3390,N_2611);
and U4940 (N_4940,N_3696,N_3039);
or U4941 (N_4941,N_2802,N_3740);
or U4942 (N_4942,N_3226,N_3453);
and U4943 (N_4943,N_3154,N_3549);
xnor U4944 (N_4944,N_2981,N_2559);
and U4945 (N_4945,N_3598,N_3224);
nand U4946 (N_4946,N_2907,N_3637);
and U4947 (N_4947,N_3508,N_2846);
or U4948 (N_4948,N_3317,N_3380);
or U4949 (N_4949,N_3550,N_3400);
xor U4950 (N_4950,N_2549,N_2651);
and U4951 (N_4951,N_2915,N_2838);
or U4952 (N_4952,N_3378,N_2966);
nor U4953 (N_4953,N_2618,N_2573);
nor U4954 (N_4954,N_3409,N_3334);
and U4955 (N_4955,N_3150,N_2731);
xnor U4956 (N_4956,N_2858,N_2506);
xor U4957 (N_4957,N_2719,N_2515);
or U4958 (N_4958,N_3204,N_2759);
and U4959 (N_4959,N_3523,N_3068);
and U4960 (N_4960,N_3027,N_3672);
nand U4961 (N_4961,N_2894,N_3082);
and U4962 (N_4962,N_3398,N_3110);
nand U4963 (N_4963,N_3117,N_2745);
xor U4964 (N_4964,N_2666,N_2978);
or U4965 (N_4965,N_3446,N_3138);
nand U4966 (N_4966,N_2737,N_3079);
and U4967 (N_4967,N_3608,N_3083);
or U4968 (N_4968,N_2968,N_2707);
and U4969 (N_4969,N_2509,N_3454);
and U4970 (N_4970,N_3192,N_2904);
nor U4971 (N_4971,N_3600,N_2749);
xnor U4972 (N_4972,N_2743,N_2910);
or U4973 (N_4973,N_3571,N_3067);
nor U4974 (N_4974,N_3402,N_3724);
xor U4975 (N_4975,N_3175,N_3304);
or U4976 (N_4976,N_3535,N_3676);
or U4977 (N_4977,N_3374,N_3574);
or U4978 (N_4978,N_3597,N_2620);
or U4979 (N_4979,N_3155,N_2960);
nor U4980 (N_4980,N_2607,N_3746);
nor U4981 (N_4981,N_3142,N_3183);
nor U4982 (N_4982,N_3028,N_2813);
nand U4983 (N_4983,N_2656,N_3133);
xor U4984 (N_4984,N_2877,N_3340);
nor U4985 (N_4985,N_3390,N_3482);
and U4986 (N_4986,N_2774,N_3219);
nand U4987 (N_4987,N_2526,N_3089);
and U4988 (N_4988,N_3398,N_2673);
and U4989 (N_4989,N_3495,N_3435);
nor U4990 (N_4990,N_2770,N_3076);
nand U4991 (N_4991,N_3535,N_3485);
xnor U4992 (N_4992,N_2823,N_2675);
xnor U4993 (N_4993,N_2882,N_3145);
nor U4994 (N_4994,N_3382,N_3624);
xnor U4995 (N_4995,N_3557,N_2660);
nand U4996 (N_4996,N_2573,N_2522);
nor U4997 (N_4997,N_3666,N_2886);
nor U4998 (N_4998,N_3393,N_3192);
xor U4999 (N_4999,N_3109,N_3654);
or U5000 (N_5000,N_3798,N_4607);
nor U5001 (N_5001,N_4597,N_4454);
and U5002 (N_5002,N_3985,N_4845);
xor U5003 (N_5003,N_4494,N_4295);
nand U5004 (N_5004,N_3992,N_4830);
nor U5005 (N_5005,N_4382,N_4620);
nor U5006 (N_5006,N_3811,N_4867);
nor U5007 (N_5007,N_4901,N_4157);
xnor U5008 (N_5008,N_3921,N_4812);
nor U5009 (N_5009,N_3754,N_4953);
nand U5010 (N_5010,N_3795,N_4720);
xor U5011 (N_5011,N_4371,N_4181);
xnor U5012 (N_5012,N_3865,N_4041);
nand U5013 (N_5013,N_4816,N_4155);
xor U5014 (N_5014,N_4228,N_4520);
or U5015 (N_5015,N_4869,N_4848);
nand U5016 (N_5016,N_4892,N_4207);
nand U5017 (N_5017,N_4459,N_4315);
or U5018 (N_5018,N_4254,N_4543);
nand U5019 (N_5019,N_4272,N_4193);
nor U5020 (N_5020,N_4870,N_4279);
nand U5021 (N_5021,N_4269,N_4137);
and U5022 (N_5022,N_4646,N_4366);
and U5023 (N_5023,N_4831,N_4813);
or U5024 (N_5024,N_4145,N_4495);
xnor U5025 (N_5025,N_4796,N_4426);
and U5026 (N_5026,N_4277,N_4955);
nand U5027 (N_5027,N_4350,N_4463);
and U5028 (N_5028,N_4839,N_4281);
xnor U5029 (N_5029,N_4648,N_4379);
and U5030 (N_5030,N_4466,N_4149);
or U5031 (N_5031,N_4310,N_4694);
nand U5032 (N_5032,N_4725,N_4726);
and U5033 (N_5033,N_4052,N_4227);
nand U5034 (N_5034,N_4095,N_4922);
or U5035 (N_5035,N_4417,N_3782);
nand U5036 (N_5036,N_4670,N_4067);
nand U5037 (N_5037,N_3825,N_4351);
nand U5038 (N_5038,N_3880,N_4159);
xor U5039 (N_5039,N_4802,N_4636);
nor U5040 (N_5040,N_3955,N_4630);
nand U5041 (N_5041,N_4151,N_4943);
nor U5042 (N_5042,N_4478,N_4480);
xor U5043 (N_5043,N_4788,N_3849);
nor U5044 (N_5044,N_4912,N_3853);
and U5045 (N_5045,N_4567,N_4642);
nor U5046 (N_5046,N_3889,N_4942);
and U5047 (N_5047,N_4563,N_3790);
or U5048 (N_5048,N_4069,N_3786);
nand U5049 (N_5049,N_4924,N_4045);
xor U5050 (N_5050,N_3924,N_3855);
nor U5051 (N_5051,N_4316,N_4001);
and U5052 (N_5052,N_4588,N_4732);
xor U5053 (N_5053,N_4217,N_4828);
xnor U5054 (N_5054,N_4598,N_4797);
and U5055 (N_5055,N_4715,N_4074);
and U5056 (N_5056,N_4457,N_4532);
nor U5057 (N_5057,N_4821,N_4283);
and U5058 (N_5058,N_4474,N_4589);
xor U5059 (N_5059,N_4171,N_3763);
nor U5060 (N_5060,N_3943,N_4215);
nor U5061 (N_5061,N_4083,N_3812);
or U5062 (N_5062,N_4179,N_4296);
nand U5063 (N_5063,N_4411,N_3820);
xor U5064 (N_5064,N_4496,N_3808);
or U5065 (N_5065,N_4147,N_4339);
xnor U5066 (N_5066,N_4110,N_3872);
nand U5067 (N_5067,N_4587,N_4262);
xor U5068 (N_5068,N_4218,N_3892);
or U5069 (N_5069,N_4745,N_4574);
nand U5070 (N_5070,N_4306,N_4618);
and U5071 (N_5071,N_4609,N_4432);
and U5072 (N_5072,N_4559,N_3902);
nor U5073 (N_5073,N_4723,N_4486);
and U5074 (N_5074,N_4195,N_3982);
or U5075 (N_5075,N_3996,N_4572);
or U5076 (N_5076,N_4801,N_4011);
xor U5077 (N_5077,N_4968,N_3914);
and U5078 (N_5078,N_4483,N_4441);
nand U5079 (N_5079,N_3874,N_4499);
or U5080 (N_5080,N_4319,N_3831);
nand U5081 (N_5081,N_4026,N_4043);
nor U5082 (N_5082,N_4142,N_4952);
nand U5083 (N_5083,N_4234,N_4687);
and U5084 (N_5084,N_4040,N_4448);
and U5085 (N_5085,N_4754,N_4513);
xor U5086 (N_5086,N_4073,N_4577);
and U5087 (N_5087,N_4396,N_4834);
nor U5088 (N_5088,N_4639,N_4487);
nand U5089 (N_5089,N_4879,N_3962);
xnor U5090 (N_5090,N_4717,N_4722);
and U5091 (N_5091,N_4086,N_4300);
xor U5092 (N_5092,N_4789,N_3884);
and U5093 (N_5093,N_4521,N_4603);
nand U5094 (N_5094,N_4772,N_4685);
and U5095 (N_5095,N_4003,N_3964);
or U5096 (N_5096,N_3823,N_4014);
or U5097 (N_5097,N_3922,N_3802);
nor U5098 (N_5098,N_3862,N_4158);
or U5099 (N_5099,N_4966,N_4187);
nand U5100 (N_5100,N_4427,N_4194);
and U5101 (N_5101,N_4883,N_4744);
xor U5102 (N_5102,N_4961,N_4735);
nor U5103 (N_5103,N_4767,N_4501);
nand U5104 (N_5104,N_4233,N_4053);
xnor U5105 (N_5105,N_3988,N_4653);
and U5106 (N_5106,N_4539,N_4492);
or U5107 (N_5107,N_3828,N_3885);
and U5108 (N_5108,N_4247,N_4177);
nor U5109 (N_5109,N_4707,N_3908);
xor U5110 (N_5110,N_4554,N_4519);
and U5111 (N_5111,N_4370,N_3761);
and U5112 (N_5112,N_3947,N_4470);
and U5113 (N_5113,N_4665,N_4399);
or U5114 (N_5114,N_4699,N_4032);
or U5115 (N_5115,N_4355,N_4395);
xor U5116 (N_5116,N_4547,N_4743);
and U5117 (N_5117,N_4645,N_4220);
xor U5118 (N_5118,N_4622,N_4993);
or U5119 (N_5119,N_3861,N_3838);
and U5120 (N_5120,N_4184,N_4757);
and U5121 (N_5121,N_4030,N_4855);
and U5122 (N_5122,N_4673,N_3777);
or U5123 (N_5123,N_3850,N_3762);
and U5124 (N_5124,N_4340,N_4736);
or U5125 (N_5125,N_3824,N_4376);
and U5126 (N_5126,N_4321,N_4654);
and U5127 (N_5127,N_4460,N_4777);
or U5128 (N_5128,N_4061,N_4275);
nand U5129 (N_5129,N_4063,N_4616);
and U5130 (N_5130,N_4257,N_4192);
nand U5131 (N_5131,N_4730,N_4581);
and U5132 (N_5132,N_4336,N_4889);
or U5133 (N_5133,N_4498,N_3806);
or U5134 (N_5134,N_4594,N_4927);
xnor U5135 (N_5135,N_4443,N_3876);
xnor U5136 (N_5136,N_4174,N_4141);
and U5137 (N_5137,N_3900,N_4239);
or U5138 (N_5138,N_4337,N_3839);
and U5139 (N_5139,N_4655,N_3793);
xnor U5140 (N_5140,N_4204,N_4437);
nor U5141 (N_5141,N_4982,N_4557);
nand U5142 (N_5142,N_4223,N_3863);
and U5143 (N_5143,N_4050,N_3773);
nand U5144 (N_5144,N_4225,N_4154);
nor U5145 (N_5145,N_4138,N_4540);
or U5146 (N_5146,N_4529,N_3909);
and U5147 (N_5147,N_4170,N_4168);
and U5148 (N_5148,N_4710,N_4768);
or U5149 (N_5149,N_4826,N_4209);
nand U5150 (N_5150,N_3835,N_4858);
nor U5151 (N_5151,N_4012,N_4515);
and U5152 (N_5152,N_4909,N_4385);
or U5153 (N_5153,N_4129,N_4760);
and U5154 (N_5154,N_4933,N_3784);
nand U5155 (N_5155,N_4114,N_4847);
nor U5156 (N_5156,N_4746,N_4614);
and U5157 (N_5157,N_4684,N_4438);
or U5158 (N_5158,N_4775,N_4886);
or U5159 (N_5159,N_4005,N_4527);
nor U5160 (N_5160,N_4271,N_3857);
nand U5161 (N_5161,N_4358,N_4903);
and U5162 (N_5162,N_4629,N_3851);
nor U5163 (N_5163,N_3774,N_4907);
nor U5164 (N_5164,N_3843,N_4156);
and U5165 (N_5165,N_3870,N_4435);
or U5166 (N_5166,N_4123,N_4373);
or U5167 (N_5167,N_4561,N_4851);
or U5168 (N_5168,N_3966,N_4708);
nor U5169 (N_5169,N_4844,N_4562);
nor U5170 (N_5170,N_3928,N_4335);
and U5171 (N_5171,N_4880,N_4731);
nor U5172 (N_5172,N_4128,N_4226);
nor U5173 (N_5173,N_4606,N_4660);
and U5174 (N_5174,N_3907,N_3965);
nor U5175 (N_5175,N_4028,N_4800);
xnor U5176 (N_5176,N_4268,N_4798);
nor U5177 (N_5177,N_3771,N_4442);
and U5178 (N_5178,N_4596,N_4795);
nor U5179 (N_5179,N_4092,N_4412);
and U5180 (N_5180,N_3933,N_3912);
nand U5181 (N_5181,N_4439,N_4163);
or U5182 (N_5182,N_3875,N_4444);
nor U5183 (N_5183,N_4747,N_4465);
or U5184 (N_5184,N_4238,N_4549);
nor U5185 (N_5185,N_4998,N_4729);
xor U5186 (N_5186,N_4160,N_4130);
nand U5187 (N_5187,N_4458,N_4065);
and U5188 (N_5188,N_4294,N_4688);
or U5189 (N_5189,N_3953,N_3967);
or U5190 (N_5190,N_3954,N_4936);
or U5191 (N_5191,N_4477,N_4348);
nand U5192 (N_5192,N_3856,N_4236);
nor U5193 (N_5193,N_4134,N_4692);
nor U5194 (N_5194,N_4786,N_4428);
nor U5195 (N_5195,N_4097,N_3958);
and U5196 (N_5196,N_4285,N_4049);
nand U5197 (N_5197,N_4656,N_4332);
or U5198 (N_5198,N_4910,N_4771);
or U5199 (N_5199,N_4921,N_4491);
or U5200 (N_5200,N_4183,N_4493);
nand U5201 (N_5201,N_4716,N_3877);
nor U5202 (N_5202,N_4817,N_4605);
nor U5203 (N_5203,N_3886,N_3927);
nand U5204 (N_5204,N_4000,N_3893);
or U5205 (N_5205,N_4558,N_3923);
xnor U5206 (N_5206,N_3829,N_3890);
or U5207 (N_5207,N_4996,N_4201);
or U5208 (N_5208,N_4017,N_4765);
or U5209 (N_5209,N_4770,N_4825);
nand U5210 (N_5210,N_4750,N_4256);
nand U5211 (N_5211,N_4278,N_4485);
xnor U5212 (N_5212,N_4693,N_4689);
xnor U5213 (N_5213,N_4308,N_4674);
or U5214 (N_5214,N_4132,N_4971);
nor U5215 (N_5215,N_4553,N_4956);
xnor U5216 (N_5216,N_4051,N_4713);
nor U5217 (N_5217,N_4579,N_4944);
nand U5218 (N_5218,N_4945,N_4230);
nor U5219 (N_5219,N_4785,N_4790);
xor U5220 (N_5220,N_4140,N_4829);
xor U5221 (N_5221,N_4117,N_4314);
xor U5222 (N_5222,N_4734,N_4251);
nand U5223 (N_5223,N_3977,N_4887);
xor U5224 (N_5224,N_3844,N_4102);
or U5225 (N_5225,N_4662,N_4222);
nor U5226 (N_5226,N_3887,N_4231);
and U5227 (N_5227,N_4377,N_3867);
nor U5228 (N_5228,N_4619,N_4364);
and U5229 (N_5229,N_4015,N_4506);
nand U5230 (N_5230,N_4946,N_3956);
nor U5231 (N_5231,N_4926,N_4803);
xnor U5232 (N_5232,N_4585,N_4988);
nor U5233 (N_5233,N_4891,N_4368);
nor U5234 (N_5234,N_4449,N_3792);
and U5235 (N_5235,N_4108,N_4995);
xor U5236 (N_5236,N_4914,N_4682);
nor U5237 (N_5237,N_4651,N_4447);
and U5238 (N_5238,N_4111,N_4404);
or U5239 (N_5239,N_3997,N_4677);
xnor U5240 (N_5240,N_4482,N_4548);
nor U5241 (N_5241,N_4416,N_4905);
nand U5242 (N_5242,N_3915,N_4071);
or U5243 (N_5243,N_4161,N_4057);
xnor U5244 (N_5244,N_3847,N_4804);
nand U5245 (N_5245,N_4556,N_4068);
and U5246 (N_5246,N_3934,N_4104);
xnor U5247 (N_5247,N_4512,N_4895);
nor U5248 (N_5248,N_4056,N_4490);
nor U5249 (N_5249,N_4591,N_4313);
and U5250 (N_5250,N_4617,N_4126);
nor U5251 (N_5251,N_4224,N_4873);
or U5252 (N_5252,N_4809,N_4343);
or U5253 (N_5253,N_4560,N_3832);
or U5254 (N_5254,N_3879,N_4601);
xnor U5255 (N_5255,N_4472,N_4590);
nand U5256 (N_5256,N_4211,N_4488);
nor U5257 (N_5257,N_3987,N_4253);
nand U5258 (N_5258,N_4143,N_3904);
nor U5259 (N_5259,N_4721,N_3791);
and U5260 (N_5260,N_4260,N_4626);
xnor U5261 (N_5261,N_4352,N_4446);
nand U5262 (N_5262,N_4349,N_4375);
xnor U5263 (N_5263,N_4960,N_4697);
and U5264 (N_5264,N_4182,N_4362);
or U5265 (N_5265,N_4538,N_4748);
nor U5266 (N_5266,N_4584,N_3895);
and U5267 (N_5267,N_4394,N_4451);
nand U5268 (N_5268,N_4706,N_4534);
nand U5269 (N_5269,N_4862,N_3899);
and U5270 (N_5270,N_4695,N_4401);
xor U5271 (N_5271,N_4365,N_3871);
nand U5272 (N_5272,N_4739,N_4380);
and U5273 (N_5273,N_4301,N_4890);
and U5274 (N_5274,N_4245,N_3752);
nand U5275 (N_5275,N_4672,N_3837);
nor U5276 (N_5276,N_3878,N_4628);
nand U5277 (N_5277,N_4980,N_4243);
and U5278 (N_5278,N_4810,N_4530);
or U5279 (N_5279,N_4633,N_3983);
nor U5280 (N_5280,N_4240,N_4038);
nor U5281 (N_5281,N_4523,N_4390);
nand U5282 (N_5282,N_4913,N_3750);
nor U5283 (N_5283,N_4386,N_4020);
xnor U5284 (N_5284,N_4302,N_4525);
or U5285 (N_5285,N_4611,N_4450);
nand U5286 (N_5286,N_4309,N_4324);
nand U5287 (N_5287,N_3926,N_4464);
or U5288 (N_5288,N_4524,N_4468);
and U5289 (N_5289,N_4080,N_4793);
or U5290 (N_5290,N_4019,N_4075);
xor U5291 (N_5291,N_4678,N_4081);
xor U5292 (N_5292,N_4929,N_4514);
xnor U5293 (N_5293,N_4774,N_4219);
xor U5294 (N_5294,N_3797,N_3801);
or U5295 (N_5295,N_4421,N_3898);
xnor U5296 (N_5296,N_4415,N_3783);
or U5297 (N_5297,N_4911,N_3767);
or U5298 (N_5298,N_3938,N_4778);
or U5299 (N_5299,N_4303,N_4393);
nor U5300 (N_5300,N_4334,N_4811);
xor U5301 (N_5301,N_4016,N_4361);
xnor U5302 (N_5302,N_4344,N_4904);
nand U5303 (N_5303,N_4144,N_4106);
and U5304 (N_5304,N_4461,N_4205);
or U5305 (N_5305,N_3920,N_4763);
xnor U5306 (N_5306,N_4741,N_4101);
xor U5307 (N_5307,N_4121,N_4383);
xor U5308 (N_5308,N_4923,N_4027);
xnor U5309 (N_5309,N_4791,N_4263);
nor U5310 (N_5310,N_4666,N_3971);
and U5311 (N_5311,N_4997,N_4479);
nand U5312 (N_5312,N_4249,N_3807);
or U5313 (N_5313,N_4103,N_4714);
nor U5314 (N_5314,N_3766,N_3978);
xor U5315 (N_5315,N_4954,N_4518);
nand U5316 (N_5316,N_4570,N_4854);
or U5317 (N_5317,N_4794,N_4055);
and U5318 (N_5318,N_4551,N_4510);
and U5319 (N_5319,N_4004,N_3776);
nor U5320 (N_5320,N_3990,N_3957);
xor U5321 (N_5321,N_3869,N_3960);
nand U5322 (N_5322,N_4719,N_4109);
and U5323 (N_5323,N_4152,N_4631);
nor U5324 (N_5324,N_4400,N_4162);
nand U5325 (N_5325,N_4190,N_4659);
and U5326 (N_5326,N_3975,N_4328);
nand U5327 (N_5327,N_4657,N_4838);
xnor U5328 (N_5328,N_4203,N_4273);
nand U5329 (N_5329,N_4987,N_4724);
nand U5330 (N_5330,N_4852,N_4761);
nand U5331 (N_5331,N_4918,N_4850);
xor U5332 (N_5332,N_4894,N_4031);
and U5333 (N_5333,N_4718,N_3854);
or U5334 (N_5334,N_3834,N_3950);
or U5335 (N_5335,N_4843,N_4976);
or U5336 (N_5336,N_4196,N_4388);
nand U5337 (N_5337,N_4330,N_3827);
nor U5338 (N_5338,N_4916,N_3944);
and U5339 (N_5339,N_3946,N_4503);
or U5340 (N_5340,N_4507,N_4359);
nand U5341 (N_5341,N_4089,N_4832);
or U5342 (N_5342,N_4007,N_4827);
xnor U5343 (N_5343,N_4882,N_4799);
nor U5344 (N_5344,N_3787,N_4116);
xor U5345 (N_5345,N_3785,N_4919);
and U5346 (N_5346,N_4042,N_4701);
xnor U5347 (N_5347,N_4807,N_4341);
nand U5348 (N_5348,N_3813,N_4469);
nor U5349 (N_5349,N_4649,N_4476);
nor U5350 (N_5350,N_4244,N_4978);
xnor U5351 (N_5351,N_3840,N_4002);
and U5352 (N_5352,N_4602,N_4599);
nor U5353 (N_5353,N_4897,N_3999);
nor U5354 (N_5354,N_4679,N_4902);
or U5355 (N_5355,N_4938,N_4197);
xnor U5356 (N_5356,N_4221,N_4769);
xor U5357 (N_5357,N_4752,N_4006);
xnor U5358 (N_5358,N_4727,N_3984);
or U5359 (N_5359,N_4323,N_4690);
nand U5360 (N_5360,N_4806,N_4608);
nor U5361 (N_5361,N_4571,N_4863);
and U5362 (N_5362,N_4917,N_4951);
or U5363 (N_5363,N_4835,N_4504);
and U5364 (N_5364,N_4984,N_4876);
nand U5365 (N_5365,N_4232,N_4868);
nand U5366 (N_5366,N_4210,N_4877);
xnor U5367 (N_5367,N_4823,N_4422);
xnor U5368 (N_5368,N_4173,N_4389);
xor U5369 (N_5369,N_3882,N_4787);
nand U5370 (N_5370,N_4311,N_4932);
or U5371 (N_5371,N_4737,N_4928);
xor U5372 (N_5372,N_4888,N_4583);
and U5373 (N_5373,N_4345,N_4985);
and U5374 (N_5374,N_3845,N_3976);
and U5375 (N_5375,N_4280,N_4105);
nor U5376 (N_5376,N_3918,N_3753);
nand U5377 (N_5377,N_4191,N_3910);
and U5378 (N_5378,N_4508,N_4047);
nand U5379 (N_5379,N_4299,N_4169);
nor U5380 (N_5380,N_4500,N_4833);
and U5381 (N_5381,N_4819,N_4044);
nand U5382 (N_5382,N_3816,N_4632);
nor U5383 (N_5383,N_4093,N_4267);
xor U5384 (N_5384,N_4934,N_4552);
xnor U5385 (N_5385,N_4096,N_4112);
nor U5386 (N_5386,N_3758,N_4118);
nand U5387 (N_5387,N_4008,N_4150);
nand U5388 (N_5388,N_4974,N_4975);
xor U5389 (N_5389,N_4545,N_4088);
xor U5390 (N_5390,N_4125,N_4317);
xor U5391 (N_5391,N_4291,N_4392);
nor U5392 (N_5392,N_4808,N_4431);
nor U5393 (N_5393,N_4270,N_4079);
nand U5394 (N_5394,N_4286,N_4255);
or U5395 (N_5395,N_3842,N_4756);
nor U5396 (N_5396,N_4024,N_4462);
or U5397 (N_5397,N_3822,N_4958);
nor U5398 (N_5398,N_3788,N_4409);
xor U5399 (N_5399,N_4066,N_4013);
and U5400 (N_5400,N_4592,N_3836);
nand U5401 (N_5401,N_4582,N_4347);
nand U5402 (N_5402,N_4555,N_3809);
xor U5403 (N_5403,N_4680,N_4021);
nor U5404 (N_5404,N_4683,N_4546);
nor U5405 (N_5405,N_4082,N_3780);
nor U5406 (N_5406,N_3841,N_4696);
or U5407 (N_5407,N_4039,N_4989);
or U5408 (N_5408,N_3751,N_4758);
and U5409 (N_5409,N_3852,N_4640);
and U5410 (N_5410,N_4070,N_3932);
or U5411 (N_5411,N_3858,N_3868);
nand U5412 (N_5412,N_3759,N_3757);
nand U5413 (N_5413,N_4010,N_4304);
nor U5414 (N_5414,N_4372,N_4935);
nor U5415 (N_5415,N_4456,N_4091);
or U5416 (N_5416,N_4864,N_3963);
xnor U5417 (N_5417,N_4189,N_4973);
nand U5418 (N_5418,N_4526,N_4658);
nand U5419 (N_5419,N_4290,N_3781);
nor U5420 (N_5420,N_3951,N_4397);
nor U5421 (N_5421,N_4753,N_3768);
nand U5422 (N_5422,N_4638,N_4733);
nor U5423 (N_5423,N_4516,N_3796);
or U5424 (N_5424,N_4094,N_4325);
and U5425 (N_5425,N_3859,N_4363);
nand U5426 (N_5426,N_4509,N_3937);
or U5427 (N_5427,N_4969,N_4078);
nor U5428 (N_5428,N_4113,N_4931);
and U5429 (N_5429,N_4610,N_4282);
and U5430 (N_5430,N_4025,N_3905);
nor U5431 (N_5431,N_4124,N_4398);
xor U5432 (N_5432,N_4505,N_4511);
nand U5433 (N_5433,N_4354,N_3848);
and U5434 (N_5434,N_4738,N_3939);
and U5435 (N_5435,N_4434,N_4625);
nor U5436 (N_5436,N_4836,N_4528);
or U5437 (N_5437,N_4406,N_4896);
or U5438 (N_5438,N_3952,N_3949);
nor U5439 (N_5439,N_4176,N_4235);
nand U5440 (N_5440,N_4849,N_4972);
nand U5441 (N_5441,N_4403,N_4861);
nand U5442 (N_5442,N_4535,N_4650);
xnor U5443 (N_5443,N_4261,N_4740);
and U5444 (N_5444,N_4467,N_4119);
xor U5445 (N_5445,N_4764,N_4357);
or U5446 (N_5446,N_4367,N_4623);
nand U5447 (N_5447,N_3998,N_4100);
nand U5448 (N_5448,N_4686,N_3896);
xnor U5449 (N_5449,N_4698,N_4425);
nand U5450 (N_5450,N_4214,N_4107);
xnor U5451 (N_5451,N_4172,N_4779);
or U5452 (N_5452,N_4387,N_3778);
xnor U5453 (N_5453,N_3959,N_3873);
or U5454 (N_5454,N_4120,N_4212);
and U5455 (N_5455,N_4898,N_4573);
xnor U5456 (N_5456,N_3931,N_4940);
nand U5457 (N_5457,N_3818,N_4115);
nor U5458 (N_5458,N_3911,N_4408);
nor U5459 (N_5459,N_4522,N_4815);
or U5460 (N_5460,N_4644,N_4994);
nor U5461 (N_5461,N_4578,N_4333);
nor U5462 (N_5462,N_4180,N_4676);
and U5463 (N_5463,N_4637,N_4568);
xnor U5464 (N_5464,N_4430,N_4884);
or U5465 (N_5465,N_3972,N_4615);
xor U5466 (N_5466,N_4949,N_3968);
nand U5467 (N_5467,N_4035,N_4292);
nand U5468 (N_5468,N_4153,N_3779);
nand U5469 (N_5469,N_4937,N_4675);
nand U5470 (N_5470,N_4920,N_4131);
and U5471 (N_5471,N_4705,N_4381);
or U5472 (N_5472,N_4178,N_4188);
or U5473 (N_5473,N_4139,N_4391);
xor U5474 (N_5474,N_4704,N_4420);
nand U5475 (N_5475,N_4959,N_4320);
nor U5476 (N_5476,N_4497,N_4840);
xor U5477 (N_5477,N_4353,N_4077);
nand U5478 (N_5478,N_4569,N_4908);
and U5479 (N_5479,N_4122,N_3945);
xnor U5480 (N_5480,N_4436,N_3770);
or U5481 (N_5481,N_4133,N_4700);
nand U5482 (N_5482,N_4580,N_3881);
or U5483 (N_5483,N_4058,N_4703);
nor U5484 (N_5484,N_4893,N_3929);
and U5485 (N_5485,N_4846,N_4652);
or U5486 (N_5486,N_4185,N_4085);
and U5487 (N_5487,N_3772,N_4762);
nand U5488 (N_5488,N_4208,N_4820);
nand U5489 (N_5489,N_4202,N_4517);
nor U5490 (N_5490,N_4647,N_4419);
nor U5491 (N_5491,N_4664,N_4950);
nand U5492 (N_5492,N_3980,N_4780);
or U5493 (N_5493,N_3940,N_3760);
and U5494 (N_5494,N_3969,N_4586);
and U5495 (N_5495,N_4537,N_4076);
nand U5496 (N_5496,N_4288,N_4668);
xor U5497 (N_5497,N_4979,N_3833);
xor U5498 (N_5498,N_3986,N_4440);
or U5499 (N_5499,N_4175,N_3989);
and U5500 (N_5500,N_4742,N_3866);
and U5501 (N_5501,N_4136,N_4248);
nor U5502 (N_5502,N_4087,N_4792);
xor U5503 (N_5503,N_4165,N_3846);
xor U5504 (N_5504,N_4252,N_4098);
xor U5505 (N_5505,N_3817,N_3799);
nand U5506 (N_5506,N_4776,N_4374);
nand U5507 (N_5507,N_4635,N_4681);
nand U5508 (N_5508,N_4413,N_4930);
nor U5509 (N_5509,N_3814,N_4072);
and U5510 (N_5510,N_4414,N_4298);
and U5511 (N_5511,N_4751,N_4595);
or U5512 (N_5512,N_4407,N_3883);
xor U5513 (N_5513,N_4022,N_4062);
and U5514 (N_5514,N_4213,N_4878);
nor U5515 (N_5515,N_3919,N_3803);
nand U5516 (N_5516,N_4604,N_4146);
and U5517 (N_5517,N_4613,N_4274);
and U5518 (N_5518,N_3815,N_3897);
and U5519 (N_5519,N_3804,N_4293);
or U5520 (N_5520,N_4037,N_4473);
nand U5521 (N_5521,N_4360,N_4977);
nand U5522 (N_5522,N_4541,N_4947);
or U5523 (N_5523,N_4818,N_4536);
and U5524 (N_5524,N_4663,N_3805);
and U5525 (N_5525,N_3981,N_4783);
and U5526 (N_5526,N_4900,N_4814);
nor U5527 (N_5527,N_3864,N_4957);
nor U5528 (N_5528,N_4452,N_3948);
and U5529 (N_5529,N_4433,N_4531);
nor U5530 (N_5530,N_3775,N_4064);
xnor U5531 (N_5531,N_4711,N_4054);
nor U5532 (N_5532,N_4962,N_3789);
nor U5533 (N_5533,N_4259,N_4964);
xnor U5534 (N_5534,N_4627,N_4805);
or U5535 (N_5535,N_4963,N_4661);
nand U5536 (N_5536,N_4265,N_4036);
or U5537 (N_5537,N_4643,N_4822);
and U5538 (N_5538,N_4941,N_4544);
xor U5539 (N_5539,N_4329,N_3917);
xor U5540 (N_5540,N_4593,N_3860);
nand U5541 (N_5541,N_4533,N_4346);
and U5542 (N_5542,N_4048,N_4009);
nand U5543 (N_5543,N_3973,N_4565);
nor U5544 (N_5544,N_4899,N_4502);
or U5545 (N_5545,N_4475,N_3993);
nor U5546 (N_5546,N_4773,N_4264);
or U5547 (N_5547,N_4099,N_4148);
or U5548 (N_5548,N_4881,N_4342);
nor U5549 (N_5549,N_4216,N_4489);
and U5550 (N_5550,N_4981,N_4824);
nand U5551 (N_5551,N_4241,N_4297);
nand U5552 (N_5552,N_4484,N_3930);
nand U5553 (N_5553,N_3935,N_3765);
xor U5554 (N_5554,N_4289,N_4853);
nand U5555 (N_5555,N_4229,N_4276);
and U5556 (N_5556,N_4023,N_3942);
xnor U5557 (N_5557,N_4948,N_4749);
or U5558 (N_5558,N_4135,N_4781);
xnor U5559 (N_5559,N_4318,N_4029);
nor U5560 (N_5560,N_4199,N_4621);
nor U5561 (N_5561,N_4865,N_4250);
nor U5562 (N_5562,N_3961,N_3830);
nor U5563 (N_5563,N_4127,N_3888);
and U5564 (N_5564,N_4576,N_4669);
nor U5565 (N_5565,N_4875,N_4034);
and U5566 (N_5566,N_4356,N_3756);
xor U5567 (N_5567,N_4200,N_3913);
and U5568 (N_5568,N_3755,N_4925);
nor U5569 (N_5569,N_4284,N_4566);
and U5570 (N_5570,N_4866,N_4564);
nor U5571 (N_5571,N_4766,N_4242);
xor U5572 (N_5572,N_4455,N_4471);
or U5573 (N_5573,N_4906,N_4237);
or U5574 (N_5574,N_3974,N_4327);
nor U5575 (N_5575,N_4258,N_4755);
nand U5576 (N_5576,N_3916,N_4837);
nor U5577 (N_5577,N_4542,N_4307);
nor U5578 (N_5578,N_4641,N_4481);
or U5579 (N_5579,N_4410,N_3764);
xor U5580 (N_5580,N_4198,N_4728);
or U5581 (N_5581,N_4322,N_4287);
and U5582 (N_5582,N_4429,N_4059);
nand U5583 (N_5583,N_4575,N_4305);
or U5584 (N_5584,N_4860,N_3821);
nand U5585 (N_5585,N_4266,N_4872);
xnor U5586 (N_5586,N_4018,N_4164);
xnor U5587 (N_5587,N_4369,N_4060);
nand U5588 (N_5588,N_4702,N_3991);
nand U5589 (N_5589,N_4634,N_3769);
nor U5590 (N_5590,N_4782,N_4671);
nor U5591 (N_5591,N_3901,N_4624);
or U5592 (N_5592,N_3995,N_4186);
and U5593 (N_5593,N_3810,N_4991);
nor U5594 (N_5594,N_4857,N_4967);
nor U5595 (N_5595,N_4709,N_4859);
xnor U5596 (N_5596,N_4206,N_4691);
or U5597 (N_5597,N_4033,N_3891);
and U5598 (N_5598,N_4915,N_4842);
or U5599 (N_5599,N_4166,N_4418);
or U5600 (N_5600,N_4090,N_3800);
or U5601 (N_5601,N_4965,N_3925);
xor U5602 (N_5602,N_4970,N_4856);
nand U5603 (N_5603,N_4999,N_4453);
or U5604 (N_5604,N_4046,N_4084);
or U5605 (N_5605,N_4424,N_4983);
and U5606 (N_5606,N_4338,N_4992);
xor U5607 (N_5607,N_4326,N_3903);
and U5608 (N_5608,N_4712,N_4445);
nand U5609 (N_5609,N_4312,N_4841);
or U5610 (N_5610,N_3941,N_3936);
nand U5611 (N_5611,N_4612,N_4331);
xor U5612 (N_5612,N_4246,N_3826);
or U5613 (N_5613,N_4402,N_3970);
and U5614 (N_5614,N_4759,N_4939);
nand U5615 (N_5615,N_3994,N_4990);
nand U5616 (N_5616,N_4874,N_3894);
xnor U5617 (N_5617,N_3819,N_4871);
xnor U5618 (N_5618,N_4423,N_3979);
and U5619 (N_5619,N_4784,N_4986);
nand U5620 (N_5620,N_4600,N_4405);
and U5621 (N_5621,N_3906,N_4167);
xor U5622 (N_5622,N_4550,N_4885);
or U5623 (N_5623,N_3794,N_4378);
and U5624 (N_5624,N_4384,N_4667);
or U5625 (N_5625,N_4847,N_4945);
nand U5626 (N_5626,N_4387,N_4121);
or U5627 (N_5627,N_4496,N_4591);
or U5628 (N_5628,N_4450,N_4427);
or U5629 (N_5629,N_4090,N_4864);
nor U5630 (N_5630,N_4981,N_4532);
xnor U5631 (N_5631,N_3960,N_3784);
nor U5632 (N_5632,N_3768,N_3809);
xor U5633 (N_5633,N_4973,N_4179);
and U5634 (N_5634,N_4269,N_4920);
and U5635 (N_5635,N_4891,N_4863);
nor U5636 (N_5636,N_4665,N_4458);
xnor U5637 (N_5637,N_3849,N_4694);
nor U5638 (N_5638,N_4428,N_4909);
and U5639 (N_5639,N_4359,N_3968);
nor U5640 (N_5640,N_4946,N_4205);
xnor U5641 (N_5641,N_4690,N_3826);
nor U5642 (N_5642,N_3837,N_4952);
and U5643 (N_5643,N_4108,N_4700);
nor U5644 (N_5644,N_4902,N_4010);
xnor U5645 (N_5645,N_4003,N_4881);
nor U5646 (N_5646,N_4922,N_4713);
xor U5647 (N_5647,N_4464,N_4570);
and U5648 (N_5648,N_4398,N_4531);
nor U5649 (N_5649,N_4754,N_4255);
and U5650 (N_5650,N_4237,N_4475);
nand U5651 (N_5651,N_4673,N_4419);
nor U5652 (N_5652,N_4404,N_4567);
xnor U5653 (N_5653,N_4470,N_4127);
xnor U5654 (N_5654,N_4964,N_4084);
nor U5655 (N_5655,N_4381,N_4918);
xnor U5656 (N_5656,N_4299,N_4981);
xor U5657 (N_5657,N_4283,N_4535);
and U5658 (N_5658,N_4594,N_4070);
nand U5659 (N_5659,N_4829,N_4035);
and U5660 (N_5660,N_4188,N_3838);
xor U5661 (N_5661,N_3962,N_3751);
nor U5662 (N_5662,N_4713,N_4898);
or U5663 (N_5663,N_4753,N_4423);
nor U5664 (N_5664,N_3963,N_3983);
and U5665 (N_5665,N_3979,N_4487);
and U5666 (N_5666,N_4355,N_3996);
xor U5667 (N_5667,N_4925,N_4999);
xor U5668 (N_5668,N_4820,N_3887);
xnor U5669 (N_5669,N_3761,N_4176);
and U5670 (N_5670,N_4390,N_4149);
xnor U5671 (N_5671,N_3847,N_4861);
xnor U5672 (N_5672,N_4326,N_4801);
xnor U5673 (N_5673,N_4273,N_4447);
nor U5674 (N_5674,N_3971,N_4248);
xnor U5675 (N_5675,N_4026,N_4884);
nor U5676 (N_5676,N_4084,N_4090);
or U5677 (N_5677,N_4294,N_4737);
xor U5678 (N_5678,N_4603,N_4309);
or U5679 (N_5679,N_4246,N_4420);
and U5680 (N_5680,N_4394,N_4852);
and U5681 (N_5681,N_4366,N_3914);
and U5682 (N_5682,N_3981,N_4226);
nand U5683 (N_5683,N_4145,N_4125);
and U5684 (N_5684,N_3753,N_4824);
nor U5685 (N_5685,N_3915,N_4875);
xnor U5686 (N_5686,N_4104,N_4505);
xor U5687 (N_5687,N_4746,N_4736);
xnor U5688 (N_5688,N_4979,N_4956);
nand U5689 (N_5689,N_3761,N_4073);
nand U5690 (N_5690,N_4032,N_4873);
and U5691 (N_5691,N_4799,N_4840);
nand U5692 (N_5692,N_4086,N_4379);
or U5693 (N_5693,N_4395,N_4213);
nor U5694 (N_5694,N_3779,N_4541);
nand U5695 (N_5695,N_3790,N_4072);
nor U5696 (N_5696,N_4199,N_4019);
or U5697 (N_5697,N_4767,N_4474);
xnor U5698 (N_5698,N_4442,N_4724);
nor U5699 (N_5699,N_4441,N_4075);
nor U5700 (N_5700,N_4230,N_4852);
nor U5701 (N_5701,N_4922,N_4184);
nand U5702 (N_5702,N_4290,N_4877);
nor U5703 (N_5703,N_3877,N_4419);
or U5704 (N_5704,N_3789,N_4063);
or U5705 (N_5705,N_3981,N_3941);
or U5706 (N_5706,N_4247,N_4758);
nor U5707 (N_5707,N_4005,N_4861);
or U5708 (N_5708,N_4140,N_3941);
xnor U5709 (N_5709,N_4362,N_4484);
nand U5710 (N_5710,N_4481,N_4455);
or U5711 (N_5711,N_4635,N_4158);
nor U5712 (N_5712,N_4963,N_4028);
and U5713 (N_5713,N_3886,N_3870);
and U5714 (N_5714,N_4077,N_4504);
xor U5715 (N_5715,N_4482,N_4111);
or U5716 (N_5716,N_4861,N_4036);
and U5717 (N_5717,N_4149,N_4513);
or U5718 (N_5718,N_3817,N_4266);
and U5719 (N_5719,N_4345,N_3838);
nand U5720 (N_5720,N_4602,N_4639);
nor U5721 (N_5721,N_4462,N_4674);
nor U5722 (N_5722,N_4711,N_4169);
nand U5723 (N_5723,N_4976,N_4693);
xor U5724 (N_5724,N_4612,N_4956);
xor U5725 (N_5725,N_4285,N_4263);
or U5726 (N_5726,N_4255,N_4324);
xor U5727 (N_5727,N_3928,N_3867);
nor U5728 (N_5728,N_4414,N_4826);
or U5729 (N_5729,N_3986,N_4205);
nor U5730 (N_5730,N_4525,N_4767);
nor U5731 (N_5731,N_4590,N_4906);
or U5732 (N_5732,N_3914,N_4510);
or U5733 (N_5733,N_4388,N_3942);
nand U5734 (N_5734,N_3859,N_4336);
or U5735 (N_5735,N_4133,N_4512);
and U5736 (N_5736,N_4170,N_4409);
xor U5737 (N_5737,N_4918,N_4318);
nor U5738 (N_5738,N_4883,N_3769);
nand U5739 (N_5739,N_4065,N_3880);
nand U5740 (N_5740,N_4517,N_3928);
and U5741 (N_5741,N_4372,N_4080);
or U5742 (N_5742,N_4913,N_4860);
and U5743 (N_5743,N_4358,N_4546);
and U5744 (N_5744,N_4041,N_4271);
or U5745 (N_5745,N_3902,N_4193);
xor U5746 (N_5746,N_4846,N_4001);
nand U5747 (N_5747,N_3832,N_4222);
and U5748 (N_5748,N_4234,N_4807);
nor U5749 (N_5749,N_4449,N_4704);
nand U5750 (N_5750,N_4003,N_3869);
nor U5751 (N_5751,N_4689,N_4650);
xnor U5752 (N_5752,N_4246,N_4392);
xnor U5753 (N_5753,N_4018,N_4820);
or U5754 (N_5754,N_4388,N_4395);
or U5755 (N_5755,N_4157,N_4234);
and U5756 (N_5756,N_3951,N_4155);
and U5757 (N_5757,N_3840,N_4531);
nor U5758 (N_5758,N_4238,N_4802);
nand U5759 (N_5759,N_4680,N_3788);
and U5760 (N_5760,N_4369,N_4508);
nand U5761 (N_5761,N_4479,N_4388);
and U5762 (N_5762,N_4652,N_4732);
or U5763 (N_5763,N_4118,N_4455);
nand U5764 (N_5764,N_4652,N_3960);
xor U5765 (N_5765,N_3984,N_4031);
and U5766 (N_5766,N_4986,N_4039);
and U5767 (N_5767,N_3948,N_4317);
nand U5768 (N_5768,N_3968,N_4321);
or U5769 (N_5769,N_4570,N_4688);
nor U5770 (N_5770,N_4952,N_4647);
nand U5771 (N_5771,N_3819,N_4298);
nand U5772 (N_5772,N_4713,N_4779);
or U5773 (N_5773,N_3953,N_4088);
and U5774 (N_5774,N_4004,N_4202);
nand U5775 (N_5775,N_4104,N_4739);
xnor U5776 (N_5776,N_4865,N_4014);
nand U5777 (N_5777,N_4868,N_3898);
nor U5778 (N_5778,N_4250,N_4399);
xnor U5779 (N_5779,N_3764,N_4949);
or U5780 (N_5780,N_4510,N_4827);
nand U5781 (N_5781,N_3755,N_3810);
or U5782 (N_5782,N_4520,N_4547);
nand U5783 (N_5783,N_4091,N_4215);
xnor U5784 (N_5784,N_4251,N_4446);
nor U5785 (N_5785,N_4448,N_4656);
or U5786 (N_5786,N_4798,N_4102);
xnor U5787 (N_5787,N_4946,N_4721);
nand U5788 (N_5788,N_4593,N_4117);
or U5789 (N_5789,N_4670,N_4933);
or U5790 (N_5790,N_4496,N_4275);
nand U5791 (N_5791,N_4422,N_4749);
nor U5792 (N_5792,N_4366,N_4639);
or U5793 (N_5793,N_4840,N_4185);
nand U5794 (N_5794,N_4079,N_4352);
and U5795 (N_5795,N_4267,N_4053);
or U5796 (N_5796,N_4278,N_4480);
or U5797 (N_5797,N_4691,N_4771);
nand U5798 (N_5798,N_4267,N_4440);
or U5799 (N_5799,N_4976,N_4908);
nand U5800 (N_5800,N_4910,N_4157);
or U5801 (N_5801,N_4645,N_4698);
or U5802 (N_5802,N_4117,N_4159);
and U5803 (N_5803,N_4923,N_4823);
and U5804 (N_5804,N_4647,N_3918);
or U5805 (N_5805,N_4401,N_3937);
or U5806 (N_5806,N_4424,N_4012);
nor U5807 (N_5807,N_4127,N_3812);
and U5808 (N_5808,N_4820,N_4229);
and U5809 (N_5809,N_4318,N_4771);
and U5810 (N_5810,N_4709,N_4011);
nand U5811 (N_5811,N_4494,N_4701);
nor U5812 (N_5812,N_4652,N_3803);
nor U5813 (N_5813,N_4903,N_4671);
nor U5814 (N_5814,N_4214,N_4966);
nand U5815 (N_5815,N_4476,N_4768);
or U5816 (N_5816,N_4046,N_4025);
nand U5817 (N_5817,N_4984,N_4734);
or U5818 (N_5818,N_3842,N_4824);
nand U5819 (N_5819,N_4093,N_4089);
or U5820 (N_5820,N_4642,N_4627);
nor U5821 (N_5821,N_4822,N_4932);
and U5822 (N_5822,N_4785,N_3787);
or U5823 (N_5823,N_4652,N_4413);
nand U5824 (N_5824,N_3892,N_4256);
xor U5825 (N_5825,N_4634,N_4970);
and U5826 (N_5826,N_4281,N_4283);
or U5827 (N_5827,N_3817,N_4894);
or U5828 (N_5828,N_4182,N_4364);
nand U5829 (N_5829,N_4196,N_4169);
or U5830 (N_5830,N_4117,N_3869);
or U5831 (N_5831,N_3880,N_4575);
or U5832 (N_5832,N_4252,N_3793);
or U5833 (N_5833,N_4508,N_3884);
and U5834 (N_5834,N_3788,N_4978);
or U5835 (N_5835,N_4373,N_4086);
xnor U5836 (N_5836,N_4186,N_4817);
and U5837 (N_5837,N_4131,N_4701);
and U5838 (N_5838,N_4393,N_4609);
and U5839 (N_5839,N_4117,N_4995);
xnor U5840 (N_5840,N_3946,N_3837);
xor U5841 (N_5841,N_4687,N_4425);
and U5842 (N_5842,N_4930,N_4943);
and U5843 (N_5843,N_4827,N_4799);
xor U5844 (N_5844,N_3784,N_4782);
nor U5845 (N_5845,N_4217,N_4794);
xor U5846 (N_5846,N_4773,N_4700);
and U5847 (N_5847,N_4431,N_4536);
xor U5848 (N_5848,N_4684,N_4527);
nor U5849 (N_5849,N_3948,N_4566);
xnor U5850 (N_5850,N_4175,N_4812);
nand U5851 (N_5851,N_4993,N_3911);
and U5852 (N_5852,N_4064,N_4009);
xnor U5853 (N_5853,N_4725,N_4571);
xnor U5854 (N_5854,N_4508,N_3985);
or U5855 (N_5855,N_4000,N_4405);
and U5856 (N_5856,N_4103,N_3775);
nand U5857 (N_5857,N_4480,N_4315);
and U5858 (N_5858,N_4927,N_4763);
and U5859 (N_5859,N_3973,N_4973);
and U5860 (N_5860,N_4126,N_4255);
xnor U5861 (N_5861,N_4613,N_4952);
or U5862 (N_5862,N_4387,N_4595);
nand U5863 (N_5863,N_4329,N_4986);
nand U5864 (N_5864,N_4578,N_4958);
xor U5865 (N_5865,N_4055,N_4860);
nor U5866 (N_5866,N_3863,N_4011);
nand U5867 (N_5867,N_4413,N_4667);
and U5868 (N_5868,N_3873,N_3760);
and U5869 (N_5869,N_4177,N_4747);
and U5870 (N_5870,N_3909,N_3865);
xnor U5871 (N_5871,N_3869,N_4076);
nand U5872 (N_5872,N_3859,N_4970);
xor U5873 (N_5873,N_4080,N_4754);
and U5874 (N_5874,N_4693,N_3998);
xor U5875 (N_5875,N_4272,N_4439);
nor U5876 (N_5876,N_4757,N_4801);
nor U5877 (N_5877,N_4937,N_4085);
nor U5878 (N_5878,N_3997,N_4922);
xnor U5879 (N_5879,N_3815,N_4163);
nor U5880 (N_5880,N_4576,N_4692);
xor U5881 (N_5881,N_4755,N_3986);
and U5882 (N_5882,N_4340,N_4316);
nor U5883 (N_5883,N_4346,N_3973);
nor U5884 (N_5884,N_4048,N_4031);
nand U5885 (N_5885,N_4487,N_4425);
nand U5886 (N_5886,N_4668,N_4466);
xnor U5887 (N_5887,N_4974,N_3975);
nor U5888 (N_5888,N_4971,N_4497);
and U5889 (N_5889,N_4383,N_4842);
xor U5890 (N_5890,N_4371,N_4694);
nor U5891 (N_5891,N_4685,N_4295);
and U5892 (N_5892,N_4946,N_3924);
and U5893 (N_5893,N_4392,N_4847);
xor U5894 (N_5894,N_4935,N_4645);
and U5895 (N_5895,N_4080,N_4172);
nor U5896 (N_5896,N_4940,N_3848);
nor U5897 (N_5897,N_4327,N_4755);
and U5898 (N_5898,N_4060,N_4493);
or U5899 (N_5899,N_3884,N_3954);
and U5900 (N_5900,N_4719,N_4692);
xnor U5901 (N_5901,N_4523,N_3766);
nor U5902 (N_5902,N_4886,N_4311);
nand U5903 (N_5903,N_4229,N_4463);
nor U5904 (N_5904,N_4274,N_4312);
xnor U5905 (N_5905,N_4752,N_3898);
and U5906 (N_5906,N_3782,N_4923);
xnor U5907 (N_5907,N_4498,N_3819);
nand U5908 (N_5908,N_4604,N_4774);
and U5909 (N_5909,N_4404,N_3885);
nor U5910 (N_5910,N_4241,N_4365);
xor U5911 (N_5911,N_4685,N_4801);
nor U5912 (N_5912,N_4890,N_4406);
nor U5913 (N_5913,N_4160,N_3988);
nand U5914 (N_5914,N_3922,N_4750);
xnor U5915 (N_5915,N_4977,N_4598);
or U5916 (N_5916,N_3964,N_4597);
nor U5917 (N_5917,N_4381,N_4775);
xor U5918 (N_5918,N_4848,N_4939);
or U5919 (N_5919,N_4787,N_3982);
nor U5920 (N_5920,N_4265,N_4253);
or U5921 (N_5921,N_4236,N_4121);
and U5922 (N_5922,N_4181,N_4319);
xor U5923 (N_5923,N_4094,N_4141);
nor U5924 (N_5924,N_4563,N_4437);
or U5925 (N_5925,N_4208,N_3978);
and U5926 (N_5926,N_4807,N_4464);
or U5927 (N_5927,N_4466,N_4123);
xor U5928 (N_5928,N_4301,N_4294);
xor U5929 (N_5929,N_4076,N_3998);
or U5930 (N_5930,N_3821,N_4230);
nand U5931 (N_5931,N_4289,N_4445);
or U5932 (N_5932,N_4158,N_4353);
xnor U5933 (N_5933,N_4622,N_4146);
or U5934 (N_5934,N_3751,N_4192);
nand U5935 (N_5935,N_3904,N_4500);
xnor U5936 (N_5936,N_4672,N_4729);
and U5937 (N_5937,N_3918,N_3970);
or U5938 (N_5938,N_4070,N_3993);
and U5939 (N_5939,N_4024,N_3802);
and U5940 (N_5940,N_3795,N_3853);
nor U5941 (N_5941,N_4929,N_4926);
xor U5942 (N_5942,N_4882,N_4782);
nand U5943 (N_5943,N_4747,N_4090);
nor U5944 (N_5944,N_4706,N_4912);
nor U5945 (N_5945,N_4298,N_4789);
or U5946 (N_5946,N_4861,N_4270);
xnor U5947 (N_5947,N_4372,N_4225);
nand U5948 (N_5948,N_4592,N_3841);
and U5949 (N_5949,N_4339,N_4949);
and U5950 (N_5950,N_3811,N_3818);
nand U5951 (N_5951,N_4211,N_4368);
or U5952 (N_5952,N_4310,N_4120);
and U5953 (N_5953,N_4002,N_4980);
nand U5954 (N_5954,N_4276,N_4961);
or U5955 (N_5955,N_4236,N_4162);
nand U5956 (N_5956,N_4435,N_4333);
xor U5957 (N_5957,N_4715,N_4554);
and U5958 (N_5958,N_3788,N_4073);
xnor U5959 (N_5959,N_4901,N_4517);
nand U5960 (N_5960,N_4406,N_4056);
nor U5961 (N_5961,N_4043,N_3971);
nand U5962 (N_5962,N_4522,N_4674);
and U5963 (N_5963,N_3955,N_4511);
and U5964 (N_5964,N_4808,N_4439);
nand U5965 (N_5965,N_4268,N_3987);
and U5966 (N_5966,N_4648,N_3968);
nor U5967 (N_5967,N_4074,N_4176);
or U5968 (N_5968,N_3896,N_4504);
nor U5969 (N_5969,N_3998,N_4665);
nand U5970 (N_5970,N_3942,N_4991);
and U5971 (N_5971,N_4009,N_3874);
nor U5972 (N_5972,N_4451,N_4012);
nor U5973 (N_5973,N_4270,N_4016);
and U5974 (N_5974,N_3847,N_4210);
xor U5975 (N_5975,N_4333,N_4703);
xnor U5976 (N_5976,N_4037,N_4326);
xor U5977 (N_5977,N_4859,N_4126);
xor U5978 (N_5978,N_4524,N_4444);
and U5979 (N_5979,N_4339,N_4533);
nor U5980 (N_5980,N_4491,N_4534);
nor U5981 (N_5981,N_4189,N_4845);
and U5982 (N_5982,N_4075,N_4144);
or U5983 (N_5983,N_4570,N_3979);
nor U5984 (N_5984,N_4097,N_4794);
or U5985 (N_5985,N_4052,N_4317);
nand U5986 (N_5986,N_4734,N_4570);
xor U5987 (N_5987,N_3954,N_4769);
and U5988 (N_5988,N_3863,N_4817);
nor U5989 (N_5989,N_4931,N_3983);
and U5990 (N_5990,N_4772,N_3932);
or U5991 (N_5991,N_4198,N_4832);
xnor U5992 (N_5992,N_4336,N_3769);
and U5993 (N_5993,N_4702,N_4621);
nor U5994 (N_5994,N_4163,N_4939);
xor U5995 (N_5995,N_4302,N_4194);
nand U5996 (N_5996,N_3795,N_4862);
nor U5997 (N_5997,N_4372,N_3933);
and U5998 (N_5998,N_4898,N_4959);
xnor U5999 (N_5999,N_4511,N_4921);
nor U6000 (N_6000,N_4676,N_4591);
and U6001 (N_6001,N_4792,N_4168);
nor U6002 (N_6002,N_4283,N_4362);
nand U6003 (N_6003,N_4325,N_3784);
and U6004 (N_6004,N_4234,N_4815);
and U6005 (N_6005,N_4668,N_3763);
and U6006 (N_6006,N_4336,N_4448);
nor U6007 (N_6007,N_4377,N_3782);
and U6008 (N_6008,N_4551,N_4267);
xnor U6009 (N_6009,N_4597,N_4517);
xnor U6010 (N_6010,N_4749,N_3837);
and U6011 (N_6011,N_3806,N_4948);
xor U6012 (N_6012,N_4017,N_4623);
xor U6013 (N_6013,N_3892,N_4980);
xnor U6014 (N_6014,N_4365,N_4281);
nor U6015 (N_6015,N_3905,N_4137);
nor U6016 (N_6016,N_4628,N_4747);
nand U6017 (N_6017,N_4384,N_4745);
and U6018 (N_6018,N_3778,N_4408);
nand U6019 (N_6019,N_4438,N_4709);
and U6020 (N_6020,N_4387,N_3842);
nor U6021 (N_6021,N_4473,N_4395);
nor U6022 (N_6022,N_4405,N_4841);
and U6023 (N_6023,N_3942,N_4419);
and U6024 (N_6024,N_3835,N_3985);
xor U6025 (N_6025,N_4350,N_4701);
or U6026 (N_6026,N_4913,N_3919);
or U6027 (N_6027,N_4381,N_4145);
xor U6028 (N_6028,N_4275,N_4091);
xor U6029 (N_6029,N_3892,N_4248);
xor U6030 (N_6030,N_4384,N_4181);
nor U6031 (N_6031,N_4905,N_4487);
nor U6032 (N_6032,N_3905,N_4764);
nor U6033 (N_6033,N_4628,N_4616);
nand U6034 (N_6034,N_3818,N_4493);
nor U6035 (N_6035,N_4267,N_4235);
nand U6036 (N_6036,N_4934,N_4800);
nor U6037 (N_6037,N_3992,N_4087);
and U6038 (N_6038,N_4029,N_4623);
xnor U6039 (N_6039,N_4904,N_4082);
and U6040 (N_6040,N_4658,N_3954);
nor U6041 (N_6041,N_4965,N_3936);
or U6042 (N_6042,N_3996,N_4822);
xor U6043 (N_6043,N_4231,N_3940);
nand U6044 (N_6044,N_4777,N_3930);
or U6045 (N_6045,N_4847,N_4178);
xor U6046 (N_6046,N_4379,N_4000);
and U6047 (N_6047,N_4968,N_3885);
nand U6048 (N_6048,N_4262,N_3823);
nor U6049 (N_6049,N_4028,N_3841);
xor U6050 (N_6050,N_4109,N_4131);
or U6051 (N_6051,N_4166,N_4788);
nand U6052 (N_6052,N_4043,N_4991);
and U6053 (N_6053,N_3995,N_4661);
xor U6054 (N_6054,N_3831,N_4791);
nor U6055 (N_6055,N_4439,N_4448);
nor U6056 (N_6056,N_4180,N_4296);
and U6057 (N_6057,N_4467,N_3938);
or U6058 (N_6058,N_4251,N_4286);
nor U6059 (N_6059,N_4746,N_4808);
and U6060 (N_6060,N_4707,N_3858);
nand U6061 (N_6061,N_4183,N_3940);
and U6062 (N_6062,N_3757,N_4600);
nand U6063 (N_6063,N_4842,N_3823);
xnor U6064 (N_6064,N_4749,N_4497);
nor U6065 (N_6065,N_4951,N_3888);
and U6066 (N_6066,N_4546,N_4239);
xnor U6067 (N_6067,N_4532,N_4036);
and U6068 (N_6068,N_4333,N_4724);
nand U6069 (N_6069,N_3797,N_4994);
or U6070 (N_6070,N_3756,N_4473);
or U6071 (N_6071,N_4586,N_3951);
and U6072 (N_6072,N_4458,N_4098);
nand U6073 (N_6073,N_4365,N_3867);
or U6074 (N_6074,N_4495,N_4746);
nor U6075 (N_6075,N_3947,N_4069);
nor U6076 (N_6076,N_3924,N_3900);
and U6077 (N_6077,N_4128,N_4428);
nor U6078 (N_6078,N_4146,N_4791);
nand U6079 (N_6079,N_3936,N_4081);
or U6080 (N_6080,N_4211,N_4987);
nor U6081 (N_6081,N_4144,N_4644);
nor U6082 (N_6082,N_4760,N_3941);
or U6083 (N_6083,N_4055,N_4251);
or U6084 (N_6084,N_4610,N_4143);
or U6085 (N_6085,N_3902,N_3890);
nand U6086 (N_6086,N_4502,N_4994);
xor U6087 (N_6087,N_3940,N_3801);
nor U6088 (N_6088,N_4324,N_3760);
xnor U6089 (N_6089,N_4231,N_4982);
or U6090 (N_6090,N_4437,N_4669);
nor U6091 (N_6091,N_4904,N_4070);
or U6092 (N_6092,N_4271,N_3961);
nor U6093 (N_6093,N_3995,N_4449);
xnor U6094 (N_6094,N_4970,N_4837);
or U6095 (N_6095,N_4184,N_4490);
nor U6096 (N_6096,N_4024,N_4026);
and U6097 (N_6097,N_4399,N_4654);
or U6098 (N_6098,N_4133,N_3798);
or U6099 (N_6099,N_4420,N_4098);
nor U6100 (N_6100,N_4473,N_4895);
xor U6101 (N_6101,N_4785,N_4610);
nand U6102 (N_6102,N_4711,N_3777);
and U6103 (N_6103,N_4801,N_4914);
xor U6104 (N_6104,N_4772,N_4550);
nor U6105 (N_6105,N_3890,N_4795);
xnor U6106 (N_6106,N_4636,N_4103);
xnor U6107 (N_6107,N_4119,N_3919);
nor U6108 (N_6108,N_4239,N_4744);
nor U6109 (N_6109,N_4406,N_4100);
nand U6110 (N_6110,N_4721,N_4421);
and U6111 (N_6111,N_4183,N_3920);
or U6112 (N_6112,N_4629,N_4952);
xor U6113 (N_6113,N_4594,N_4667);
nor U6114 (N_6114,N_4513,N_3876);
nand U6115 (N_6115,N_4621,N_4272);
xnor U6116 (N_6116,N_3941,N_4894);
nand U6117 (N_6117,N_3872,N_4460);
and U6118 (N_6118,N_3850,N_3862);
nor U6119 (N_6119,N_3754,N_4600);
nand U6120 (N_6120,N_4336,N_4970);
and U6121 (N_6121,N_4042,N_4244);
nand U6122 (N_6122,N_4469,N_4132);
nor U6123 (N_6123,N_4504,N_4319);
nor U6124 (N_6124,N_4959,N_4657);
or U6125 (N_6125,N_3834,N_4574);
and U6126 (N_6126,N_4455,N_3853);
xnor U6127 (N_6127,N_4763,N_3786);
nor U6128 (N_6128,N_4904,N_4804);
or U6129 (N_6129,N_4208,N_4329);
nor U6130 (N_6130,N_4897,N_4526);
xnor U6131 (N_6131,N_3812,N_3828);
or U6132 (N_6132,N_4498,N_3947);
nor U6133 (N_6133,N_3929,N_4355);
and U6134 (N_6134,N_4294,N_4839);
or U6135 (N_6135,N_3982,N_4894);
and U6136 (N_6136,N_4514,N_4312);
or U6137 (N_6137,N_4160,N_4859);
nand U6138 (N_6138,N_4473,N_4789);
xnor U6139 (N_6139,N_4655,N_4926);
or U6140 (N_6140,N_4415,N_4294);
and U6141 (N_6141,N_4783,N_3897);
nor U6142 (N_6142,N_4329,N_3783);
or U6143 (N_6143,N_4744,N_4220);
or U6144 (N_6144,N_4571,N_4788);
xor U6145 (N_6145,N_4408,N_4238);
xnor U6146 (N_6146,N_4846,N_4800);
xor U6147 (N_6147,N_3994,N_4678);
or U6148 (N_6148,N_4790,N_4199);
xor U6149 (N_6149,N_3791,N_4461);
or U6150 (N_6150,N_4206,N_4088);
nand U6151 (N_6151,N_3995,N_4802);
nand U6152 (N_6152,N_4899,N_4956);
nand U6153 (N_6153,N_4570,N_4455);
xor U6154 (N_6154,N_4856,N_4783);
and U6155 (N_6155,N_4284,N_4954);
or U6156 (N_6156,N_4570,N_3964);
nor U6157 (N_6157,N_4714,N_4474);
xor U6158 (N_6158,N_3976,N_4261);
nor U6159 (N_6159,N_4273,N_4253);
and U6160 (N_6160,N_3801,N_4461);
and U6161 (N_6161,N_4178,N_4042);
nand U6162 (N_6162,N_4649,N_4269);
or U6163 (N_6163,N_4642,N_4780);
xor U6164 (N_6164,N_4250,N_4862);
nand U6165 (N_6165,N_4029,N_4519);
nand U6166 (N_6166,N_4352,N_4156);
and U6167 (N_6167,N_4262,N_4830);
nand U6168 (N_6168,N_4278,N_4350);
nor U6169 (N_6169,N_4022,N_4471);
xor U6170 (N_6170,N_4751,N_4111);
and U6171 (N_6171,N_3869,N_4043);
xor U6172 (N_6172,N_4640,N_3955);
and U6173 (N_6173,N_4740,N_4448);
xnor U6174 (N_6174,N_3995,N_4809);
and U6175 (N_6175,N_4465,N_4410);
nand U6176 (N_6176,N_4358,N_4487);
nand U6177 (N_6177,N_4065,N_4428);
nor U6178 (N_6178,N_4415,N_4242);
or U6179 (N_6179,N_4193,N_3996);
and U6180 (N_6180,N_4437,N_4263);
nand U6181 (N_6181,N_4416,N_4863);
and U6182 (N_6182,N_3758,N_4960);
nor U6183 (N_6183,N_4479,N_4115);
and U6184 (N_6184,N_4380,N_3828);
nand U6185 (N_6185,N_3914,N_4067);
nor U6186 (N_6186,N_4704,N_4690);
or U6187 (N_6187,N_4460,N_4838);
and U6188 (N_6188,N_4031,N_4184);
xnor U6189 (N_6189,N_4830,N_3820);
nand U6190 (N_6190,N_4664,N_3815);
or U6191 (N_6191,N_4526,N_3902);
xor U6192 (N_6192,N_4878,N_3770);
nor U6193 (N_6193,N_3770,N_4961);
xor U6194 (N_6194,N_4613,N_4427);
or U6195 (N_6195,N_4613,N_4287);
nor U6196 (N_6196,N_4432,N_4002);
xor U6197 (N_6197,N_4860,N_4346);
or U6198 (N_6198,N_4019,N_4608);
nor U6199 (N_6199,N_4100,N_4010);
nand U6200 (N_6200,N_4591,N_4760);
nor U6201 (N_6201,N_4765,N_4496);
or U6202 (N_6202,N_3931,N_4761);
and U6203 (N_6203,N_4005,N_4077);
or U6204 (N_6204,N_3859,N_4249);
or U6205 (N_6205,N_4870,N_4017);
xnor U6206 (N_6206,N_4255,N_4066);
nor U6207 (N_6207,N_4182,N_4266);
and U6208 (N_6208,N_4346,N_4606);
xnor U6209 (N_6209,N_4274,N_4353);
or U6210 (N_6210,N_4716,N_4304);
and U6211 (N_6211,N_4129,N_4135);
nand U6212 (N_6212,N_3825,N_4107);
and U6213 (N_6213,N_4746,N_4628);
or U6214 (N_6214,N_3884,N_4020);
xnor U6215 (N_6215,N_4096,N_4626);
and U6216 (N_6216,N_4476,N_4465);
nor U6217 (N_6217,N_4388,N_4808);
xor U6218 (N_6218,N_4394,N_4826);
or U6219 (N_6219,N_4661,N_4063);
nand U6220 (N_6220,N_4673,N_4765);
nor U6221 (N_6221,N_4352,N_4517);
and U6222 (N_6222,N_4822,N_4090);
nor U6223 (N_6223,N_4473,N_4925);
xor U6224 (N_6224,N_4127,N_4531);
xnor U6225 (N_6225,N_4868,N_4002);
xnor U6226 (N_6226,N_4049,N_4212);
xor U6227 (N_6227,N_4437,N_4593);
or U6228 (N_6228,N_4820,N_4668);
xor U6229 (N_6229,N_4713,N_3904);
and U6230 (N_6230,N_4248,N_4806);
or U6231 (N_6231,N_4470,N_4988);
xor U6232 (N_6232,N_4397,N_4414);
nor U6233 (N_6233,N_3935,N_3766);
nand U6234 (N_6234,N_4537,N_4128);
nor U6235 (N_6235,N_4534,N_4507);
and U6236 (N_6236,N_4062,N_4702);
nand U6237 (N_6237,N_4270,N_4320);
or U6238 (N_6238,N_3945,N_4264);
nor U6239 (N_6239,N_4031,N_4052);
and U6240 (N_6240,N_4524,N_4128);
nand U6241 (N_6241,N_4485,N_3988);
and U6242 (N_6242,N_4788,N_4881);
xor U6243 (N_6243,N_4556,N_4335);
xnor U6244 (N_6244,N_4362,N_3839);
nor U6245 (N_6245,N_4283,N_3978);
xnor U6246 (N_6246,N_4284,N_4950);
or U6247 (N_6247,N_3905,N_4778);
or U6248 (N_6248,N_4543,N_4299);
nor U6249 (N_6249,N_4784,N_3828);
nor U6250 (N_6250,N_5318,N_5574);
nor U6251 (N_6251,N_5155,N_5973);
or U6252 (N_6252,N_5436,N_5621);
and U6253 (N_6253,N_5631,N_5791);
nand U6254 (N_6254,N_5729,N_5996);
or U6255 (N_6255,N_5448,N_5961);
nor U6256 (N_6256,N_6138,N_6242);
or U6257 (N_6257,N_5854,N_6063);
xnor U6258 (N_6258,N_5607,N_5223);
nand U6259 (N_6259,N_5648,N_5569);
nand U6260 (N_6260,N_5534,N_5234);
or U6261 (N_6261,N_5893,N_5117);
xnor U6262 (N_6262,N_5404,N_6245);
or U6263 (N_6263,N_5824,N_5734);
nor U6264 (N_6264,N_5027,N_5984);
xor U6265 (N_6265,N_5979,N_6064);
nor U6266 (N_6266,N_6163,N_5221);
nand U6267 (N_6267,N_5851,N_5685);
and U6268 (N_6268,N_5178,N_5711);
xor U6269 (N_6269,N_6041,N_5741);
nand U6270 (N_6270,N_6044,N_5236);
nand U6271 (N_6271,N_5058,N_5172);
or U6272 (N_6272,N_5186,N_5225);
nor U6273 (N_6273,N_5179,N_5232);
xor U6274 (N_6274,N_6034,N_6038);
nor U6275 (N_6275,N_5654,N_5006);
and U6276 (N_6276,N_5909,N_6093);
nor U6277 (N_6277,N_6082,N_6116);
xor U6278 (N_6278,N_5972,N_5086);
or U6279 (N_6279,N_5517,N_6211);
nand U6280 (N_6280,N_5633,N_5261);
nor U6281 (N_6281,N_5803,N_6095);
xor U6282 (N_6282,N_5920,N_5750);
xor U6283 (N_6283,N_6098,N_5901);
xnor U6284 (N_6284,N_5050,N_5153);
nand U6285 (N_6285,N_5556,N_5309);
nand U6286 (N_6286,N_5670,N_5481);
nand U6287 (N_6287,N_5363,N_5141);
or U6288 (N_6288,N_6222,N_5593);
xnor U6289 (N_6289,N_5806,N_5928);
and U6290 (N_6290,N_5558,N_5549);
or U6291 (N_6291,N_5280,N_5118);
nor U6292 (N_6292,N_6081,N_5564);
nand U6293 (N_6293,N_6100,N_5158);
or U6294 (N_6294,N_5169,N_6146);
nor U6295 (N_6295,N_5532,N_5813);
xnor U6296 (N_6296,N_5783,N_6090);
or U6297 (N_6297,N_5694,N_5079);
and U6298 (N_6298,N_5908,N_5781);
nand U6299 (N_6299,N_5195,N_5679);
xnor U6300 (N_6300,N_5568,N_5767);
nand U6301 (N_6301,N_5775,N_6059);
or U6302 (N_6302,N_5090,N_5342);
xnor U6303 (N_6303,N_5367,N_5745);
nand U6304 (N_6304,N_5146,N_5020);
xnor U6305 (N_6305,N_5978,N_5965);
or U6306 (N_6306,N_5277,N_6237);
or U6307 (N_6307,N_5562,N_5859);
or U6308 (N_6308,N_5473,N_5465);
and U6309 (N_6309,N_5337,N_5387);
xor U6310 (N_6310,N_5398,N_5474);
nand U6311 (N_6311,N_5926,N_5486);
xor U6312 (N_6312,N_5552,N_5187);
nand U6313 (N_6313,N_5077,N_5608);
and U6314 (N_6314,N_5735,N_5705);
nand U6315 (N_6315,N_5625,N_5494);
and U6316 (N_6316,N_5075,N_5270);
xor U6317 (N_6317,N_6129,N_6125);
nor U6318 (N_6318,N_5408,N_5106);
nor U6319 (N_6319,N_5850,N_5435);
or U6320 (N_6320,N_5639,N_5329);
and U6321 (N_6321,N_5524,N_5683);
and U6322 (N_6322,N_5561,N_5166);
xnor U6323 (N_6323,N_6122,N_6155);
nor U6324 (N_6324,N_5061,N_5930);
nand U6325 (N_6325,N_5864,N_5489);
or U6326 (N_6326,N_5637,N_6110);
xnor U6327 (N_6327,N_5801,N_5877);
nor U6328 (N_6328,N_6230,N_5403);
or U6329 (N_6329,N_5099,N_5272);
nand U6330 (N_6330,N_5753,N_5311);
nand U6331 (N_6331,N_5134,N_5067);
or U6332 (N_6332,N_6035,N_5906);
or U6333 (N_6333,N_5014,N_5487);
nor U6334 (N_6334,N_5416,N_5400);
xnor U6335 (N_6335,N_5033,N_6235);
and U6336 (N_6336,N_5617,N_5672);
and U6337 (N_6337,N_5848,N_5248);
nor U6338 (N_6338,N_5742,N_6067);
xor U6339 (N_6339,N_5511,N_5490);
and U6340 (N_6340,N_5888,N_5205);
nand U6341 (N_6341,N_5143,N_5827);
xnor U6342 (N_6342,N_5754,N_5314);
nor U6343 (N_6343,N_5656,N_5738);
nor U6344 (N_6344,N_5343,N_6198);
and U6345 (N_6345,N_5238,N_5054);
nand U6346 (N_6346,N_5084,N_6005);
nor U6347 (N_6347,N_5304,N_5194);
nand U6348 (N_6348,N_6241,N_6246);
nand U6349 (N_6349,N_5645,N_5540);
nand U6350 (N_6350,N_6128,N_5970);
xnor U6351 (N_6351,N_5525,N_5816);
and U6352 (N_6352,N_5392,N_5004);
nor U6353 (N_6353,N_5202,N_6200);
or U6354 (N_6354,N_5912,N_5339);
or U6355 (N_6355,N_5673,N_6065);
xnor U6356 (N_6356,N_5137,N_6088);
or U6357 (N_6357,N_5456,N_5044);
xnor U6358 (N_6358,N_6109,N_5140);
nor U6359 (N_6359,N_6040,N_6154);
and U6360 (N_6360,N_5998,N_6049);
and U6361 (N_6361,N_5442,N_5315);
nor U6362 (N_6362,N_6214,N_5276);
or U6363 (N_6363,N_5021,N_5989);
xnor U6364 (N_6364,N_5340,N_5449);
nor U6365 (N_6365,N_5862,N_6055);
and U6366 (N_6366,N_5797,N_5052);
nand U6367 (N_6367,N_5265,N_5183);
nor U6368 (N_6368,N_6012,N_5778);
and U6369 (N_6369,N_6073,N_5326);
and U6370 (N_6370,N_5706,N_6213);
and U6371 (N_6371,N_5838,N_6054);
and U6372 (N_6372,N_6182,N_5779);
nor U6373 (N_6373,N_5815,N_5284);
xnor U6374 (N_6374,N_5410,N_5165);
xor U6375 (N_6375,N_5530,N_6103);
nand U6376 (N_6376,N_5127,N_5676);
xor U6377 (N_6377,N_5010,N_5768);
or U6378 (N_6378,N_5262,N_5697);
nand U6379 (N_6379,N_5063,N_5509);
nand U6380 (N_6380,N_5590,N_5375);
and U6381 (N_6381,N_5758,N_5655);
or U6382 (N_6382,N_6231,N_5802);
nand U6383 (N_6383,N_5459,N_5942);
or U6384 (N_6384,N_6078,N_5413);
nor U6385 (N_6385,N_5437,N_5461);
and U6386 (N_6386,N_6018,N_5818);
nor U6387 (N_6387,N_5136,N_5759);
xnor U6388 (N_6388,N_5068,N_5477);
or U6389 (N_6389,N_5613,N_5857);
and U6390 (N_6390,N_5689,N_5418);
nand U6391 (N_6391,N_5414,N_5446);
xnor U6392 (N_6392,N_6210,N_5045);
nor U6393 (N_6393,N_5776,N_5531);
xor U6394 (N_6394,N_5120,N_5703);
xor U6395 (N_6395,N_5514,N_5856);
or U6396 (N_6396,N_5749,N_5661);
xnor U6397 (N_6397,N_5497,N_5298);
xnor U6398 (N_6398,N_5664,N_5871);
or U6399 (N_6399,N_5757,N_5982);
xor U6400 (N_6400,N_5081,N_5233);
or U6401 (N_6401,N_5949,N_5103);
nand U6402 (N_6402,N_5880,N_6037);
xnor U6403 (N_6403,N_5839,N_5722);
nand U6404 (N_6404,N_5089,N_6002);
nor U6405 (N_6405,N_5463,N_5668);
or U6406 (N_6406,N_5059,N_5171);
and U6407 (N_6407,N_6196,N_5377);
or U6408 (N_6408,N_5313,N_5629);
or U6409 (N_6409,N_5157,N_5836);
and U6410 (N_6410,N_5080,N_5635);
nor U6411 (N_6411,N_5515,N_5152);
or U6412 (N_6412,N_5282,N_5817);
and U6413 (N_6413,N_5420,N_6173);
and U6414 (N_6414,N_5290,N_5230);
or U6415 (N_6415,N_5736,N_5538);
xnor U6416 (N_6416,N_5162,N_5247);
nor U6417 (N_6417,N_6058,N_5878);
nor U6418 (N_6418,N_5724,N_6148);
nand U6419 (N_6419,N_5189,N_5896);
xnor U6420 (N_6420,N_5500,N_5325);
and U6421 (N_6421,N_5249,N_5364);
nor U6422 (N_6422,N_5929,N_5168);
nor U6423 (N_6423,N_5201,N_5419);
or U6424 (N_6424,N_5953,N_5874);
nor U6425 (N_6425,N_5185,N_6212);
or U6426 (N_6426,N_5601,N_6145);
or U6427 (N_6427,N_6030,N_6008);
and U6428 (N_6428,N_5330,N_5885);
and U6429 (N_6429,N_5782,N_6039);
nand U6430 (N_6430,N_5115,N_5296);
nor U6431 (N_6431,N_5373,N_6003);
nand U6432 (N_6432,N_5123,N_5522);
and U6433 (N_6433,N_5701,N_5107);
xor U6434 (N_6434,N_5472,N_5612);
nor U6435 (N_6435,N_5116,N_6136);
nand U6436 (N_6436,N_5658,N_6019);
nand U6437 (N_6437,N_5662,N_6130);
or U6438 (N_6438,N_5963,N_5840);
and U6439 (N_6439,N_6203,N_5482);
nor U6440 (N_6440,N_5647,N_5110);
nor U6441 (N_6441,N_5386,N_5206);
nor U6442 (N_6442,N_5085,N_5560);
nor U6443 (N_6443,N_5678,N_6015);
and U6444 (N_6444,N_5264,N_5671);
nand U6445 (N_6445,N_5269,N_5307);
nor U6446 (N_6446,N_5826,N_5721);
nand U6447 (N_6447,N_6089,N_5731);
nor U6448 (N_6448,N_5834,N_5097);
and U6449 (N_6449,N_5865,N_6244);
nor U6450 (N_6450,N_5426,N_5091);
xor U6451 (N_6451,N_5940,N_6115);
or U6452 (N_6452,N_5135,N_5932);
and U6453 (N_6453,N_6170,N_5312);
nand U6454 (N_6454,N_5521,N_5366);
nor U6455 (N_6455,N_5698,N_6068);
or U6456 (N_6456,N_5268,N_5102);
or U6457 (N_6457,N_6147,N_6105);
xor U6458 (N_6458,N_5792,N_5257);
xor U6459 (N_6459,N_5990,N_6119);
or U6460 (N_6460,N_5597,N_6046);
nand U6461 (N_6461,N_6106,N_6162);
nor U6462 (N_6462,N_5584,N_5526);
nor U6463 (N_6463,N_6118,N_5518);
xnor U6464 (N_6464,N_6205,N_6091);
nor U6465 (N_6465,N_5475,N_6004);
or U6466 (N_6466,N_6042,N_5293);
and U6467 (N_6467,N_5962,N_5921);
and U6468 (N_6468,N_5667,N_6234);
nand U6469 (N_6469,N_5899,N_5773);
xor U6470 (N_6470,N_5148,N_5933);
and U6471 (N_6471,N_5669,N_5001);
nor U6472 (N_6472,N_5174,N_5653);
and U6473 (N_6473,N_6032,N_5287);
nand U6474 (N_6474,N_5858,N_5348);
xor U6475 (N_6475,N_5592,N_5480);
nand U6476 (N_6476,N_5390,N_5231);
and U6477 (N_6477,N_5383,N_6248);
nor U6478 (N_6478,N_6180,N_5548);
nand U6479 (N_6479,N_5034,N_5139);
xor U6480 (N_6480,N_5379,N_5362);
nand U6481 (N_6481,N_5039,N_5048);
nor U6482 (N_6482,N_5046,N_5700);
and U6483 (N_6483,N_5628,N_5837);
or U6484 (N_6484,N_5554,N_5076);
xor U6485 (N_6485,N_5991,N_5915);
nand U6486 (N_6486,N_5830,N_5567);
xnor U6487 (N_6487,N_5447,N_5646);
and U6488 (N_6488,N_5130,N_5470);
xor U6489 (N_6489,N_5555,N_5934);
and U6490 (N_6490,N_6168,N_5692);
nand U6491 (N_6491,N_5104,N_5784);
nor U6492 (N_6492,N_5986,N_5725);
or U6493 (N_6493,N_5017,N_5660);
or U6494 (N_6494,N_6216,N_5780);
nand U6495 (N_6495,N_6202,N_5108);
nand U6496 (N_6496,N_6227,N_5259);
nor U6497 (N_6497,N_5144,N_5519);
nand U6498 (N_6498,N_5787,N_6104);
and U6499 (N_6499,N_5260,N_5317);
xnor U6500 (N_6500,N_5841,N_5935);
nor U6501 (N_6501,N_5409,N_5370);
or U6502 (N_6502,N_5863,N_5804);
nand U6503 (N_6503,N_6167,N_5897);
or U6504 (N_6504,N_5995,N_6204);
or U6505 (N_6505,N_6072,N_5715);
xnor U6506 (N_6506,N_5501,N_5177);
nor U6507 (N_6507,N_6141,N_5583);
xnor U6508 (N_6508,N_5113,N_5361);
and U6509 (N_6509,N_5121,N_5273);
or U6510 (N_6510,N_6243,N_5263);
and U6511 (N_6511,N_6111,N_6190);
xor U6512 (N_6512,N_6172,N_5709);
nand U6513 (N_6513,N_5512,N_6206);
nor U6514 (N_6514,N_5714,N_5611);
and U6515 (N_6515,N_5289,N_5354);
nor U6516 (N_6516,N_5299,N_5096);
and U6517 (N_6517,N_5536,N_5902);
or U6518 (N_6518,N_5212,N_5732);
xor U6519 (N_6519,N_5083,N_5029);
xor U6520 (N_6520,N_5977,N_5422);
or U6521 (N_6521,N_5433,N_6029);
or U6522 (N_6522,N_5682,N_5417);
and U6523 (N_6523,N_5886,N_6131);
and U6524 (N_6524,N_5832,N_5770);
and U6525 (N_6525,N_5923,N_5060);
nand U6526 (N_6526,N_5873,N_5271);
or U6527 (N_6527,N_5523,N_5030);
xor U6528 (N_6528,N_5712,N_5499);
xor U6529 (N_6529,N_5037,N_6142);
and U6530 (N_6530,N_6000,N_6149);
nor U6531 (N_6531,N_6077,N_5159);
xnor U6532 (N_6532,N_6074,N_5219);
nor U6533 (N_6533,N_5726,N_6171);
or U6534 (N_6534,N_5220,N_5295);
or U6535 (N_6535,N_5710,N_5203);
nor U6536 (N_6536,N_5719,N_5895);
xor U6537 (N_6537,N_5866,N_5596);
xor U6538 (N_6538,N_5038,N_5024);
or U6539 (N_6539,N_6158,N_6087);
nand U6540 (N_6540,N_6228,N_5603);
or U6541 (N_6541,N_5095,N_5746);
or U6542 (N_6542,N_5636,N_5495);
nand U6543 (N_6543,N_5959,N_5355);
nor U6544 (N_6544,N_5376,N_5844);
and U6545 (N_6545,N_5397,N_5003);
xor U6546 (N_6546,N_5427,N_5424);
and U6547 (N_6547,N_5253,N_6229);
nand U6548 (N_6548,N_5829,N_6166);
or U6549 (N_6549,N_5411,N_6051);
or U6550 (N_6550,N_5570,N_5087);
and U6551 (N_6551,N_6143,N_5520);
xnor U6552 (N_6552,N_5160,N_5618);
nand U6553 (N_6553,N_5306,N_6057);
nor U6554 (N_6554,N_5428,N_5215);
nand U6555 (N_6555,N_5308,N_5352);
nor U6556 (N_6556,N_5550,N_5351);
xnor U6557 (N_6557,N_5772,N_6027);
or U6558 (N_6558,N_5811,N_5035);
or U6559 (N_6559,N_5580,N_5008);
xnor U6560 (N_6560,N_5345,N_6208);
or U6561 (N_6561,N_5065,N_5423);
xor U6562 (N_6562,N_5774,N_5620);
and U6563 (N_6563,N_6183,N_5755);
nor U6564 (N_6564,N_6036,N_5161);
nor U6565 (N_6565,N_5241,N_5640);
and U6566 (N_6566,N_5142,N_6062);
xor U6567 (N_6567,N_5587,N_5200);
xor U6568 (N_6568,N_5328,N_6085);
xnor U6569 (N_6569,N_6238,N_6225);
nor U6570 (N_6570,N_5630,N_5336);
and U6571 (N_6571,N_5882,N_6031);
and U6572 (N_6572,N_5717,N_5810);
xor U6573 (N_6573,N_5957,N_5430);
nand U6574 (N_6574,N_5128,N_6249);
nand U6575 (N_6575,N_5733,N_5855);
or U6576 (N_6576,N_5980,N_6033);
xnor U6577 (N_6577,N_5847,N_5796);
xor U6578 (N_6578,N_6144,N_5266);
xor U6579 (N_6579,N_5150,N_5876);
nor U6580 (N_6580,N_5237,N_5057);
and U6581 (N_6581,N_5193,N_5393);
nand U6582 (N_6582,N_5022,N_5958);
xor U6583 (N_6583,N_5529,N_5327);
nand U6584 (N_6584,N_5610,N_5216);
nor U6585 (N_6585,N_5992,N_5192);
xnor U6586 (N_6586,N_5122,N_6226);
nand U6587 (N_6587,N_6094,N_6151);
and U6588 (N_6588,N_6193,N_5031);
or U6589 (N_6589,N_5846,N_5288);
and U6590 (N_6590,N_6117,N_5124);
nand U6591 (N_6591,N_5468,N_5156);
or U6592 (N_6592,N_5498,N_6133);
xnor U6593 (N_6593,N_5566,N_6160);
xnor U6594 (N_6594,N_6217,N_5632);
xor U6595 (N_6595,N_5074,N_5283);
xnor U6596 (N_6596,N_5066,N_5747);
nor U6597 (N_6597,N_5535,N_5819);
or U6598 (N_6598,N_5011,N_6124);
xor U6599 (N_6599,N_5279,N_5297);
and U6600 (N_6600,N_5394,N_6239);
xor U6601 (N_6601,N_5385,N_6188);
nand U6602 (N_6602,N_5278,N_5492);
nor U6603 (N_6603,N_5078,N_6157);
nand U6604 (N_6604,N_5861,N_5808);
nand U6605 (N_6605,N_6123,N_5559);
xor U6606 (N_6606,N_5028,N_6159);
nand U6607 (N_6607,N_6184,N_5814);
xnor U6608 (N_6608,N_5484,N_5182);
or U6609 (N_6609,N_5347,N_5537);
nor U6610 (N_6610,N_5365,N_5922);
or U6611 (N_6611,N_5372,N_6011);
nor U6612 (N_6612,N_5586,N_6023);
xor U6613 (N_6613,N_5209,N_5184);
and U6614 (N_6614,N_5582,N_5062);
nand U6615 (N_6615,N_5955,N_6134);
or U6616 (N_6616,N_5466,N_5769);
xor U6617 (N_6617,N_5546,N_5591);
or U6618 (N_6618,N_5360,N_6247);
nand U6619 (N_6619,N_5245,N_6020);
or U6620 (N_6620,N_5589,N_5619);
and U6621 (N_6621,N_5407,N_5267);
and U6622 (N_6622,N_5378,N_5258);
nor U6623 (N_6623,N_5002,N_5936);
xor U6624 (N_6624,N_5321,N_6108);
xnor U6625 (N_6625,N_6197,N_6061);
xnor U6626 (N_6626,N_6201,N_6112);
and U6627 (N_6627,N_5666,N_5576);
and U6628 (N_6628,N_5053,N_5565);
xor U6629 (N_6629,N_5975,N_5835);
or U6630 (N_6630,N_6096,N_6047);
or U6631 (N_6631,N_5323,N_5000);
nand U6632 (N_6632,N_5469,N_5381);
nor U6633 (N_6633,N_5795,N_5310);
nand U6634 (N_6634,N_5100,N_5910);
nor U6635 (N_6635,N_5944,N_5335);
xnor U6636 (N_6636,N_5686,N_5208);
nand U6637 (N_6637,N_5539,N_5842);
nor U6638 (N_6638,N_6215,N_5688);
and U6639 (N_6639,N_5577,N_5040);
or U6640 (N_6640,N_5598,N_5240);
nand U6641 (N_6641,N_5401,N_5485);
or U6642 (N_6642,N_5649,N_5527);
nor U6643 (N_6643,N_5828,N_5704);
or U6644 (N_6644,N_5444,N_5491);
nor U6645 (N_6645,N_6024,N_5579);
and U6646 (N_6646,N_5425,N_6194);
and U6647 (N_6647,N_5431,N_5204);
nand U6648 (N_6648,N_5274,N_5250);
nor U6649 (N_6649,N_5739,N_6221);
nand U6650 (N_6650,N_6092,N_6120);
and U6651 (N_6651,N_6048,N_5251);
nor U6652 (N_6652,N_6240,N_5406);
and U6653 (N_6653,N_5971,N_5905);
and U6654 (N_6654,N_5800,N_5049);
nor U6655 (N_6655,N_5879,N_5301);
nor U6656 (N_6656,N_5690,N_5764);
xor U6657 (N_6657,N_5916,N_5023);
nand U6658 (N_6658,N_5051,N_5082);
nor U6659 (N_6659,N_5164,N_5191);
or U6660 (N_6660,N_6174,N_6009);
nand U6661 (N_6661,N_5624,N_5019);
and U6662 (N_6662,N_5508,N_5785);
or U6663 (N_6663,N_5884,N_5228);
and U6664 (N_6664,N_5384,N_5890);
xnor U6665 (N_6665,N_5239,N_5956);
nand U6666 (N_6666,N_5357,N_5765);
or U6667 (N_6667,N_5380,N_6070);
or U6668 (N_6668,N_5762,N_5305);
nand U6669 (N_6669,N_6179,N_5748);
nand U6670 (N_6670,N_5402,N_5627);
nand U6671 (N_6671,N_5547,N_5198);
xor U6672 (N_6672,N_5479,N_5939);
nor U6673 (N_6673,N_5938,N_5695);
or U6674 (N_6674,N_6083,N_5918);
and U6675 (N_6675,N_6164,N_5903);
or U6676 (N_6676,N_5013,N_5496);
xnor U6677 (N_6677,N_5359,N_5443);
xor U6678 (N_6678,N_5396,N_6102);
and U6679 (N_6679,N_5513,N_5665);
and U6680 (N_6680,N_5615,N_5088);
nor U6681 (N_6681,N_5740,N_5476);
xor U6682 (N_6682,N_5788,N_5331);
nor U6683 (N_6683,N_5925,N_5650);
xnor U6684 (N_6684,N_5285,N_5616);
nor U6685 (N_6685,N_5173,N_5641);
or U6686 (N_6686,N_5875,N_5207);
nand U6687 (N_6687,N_6165,N_5129);
nand U6688 (N_6688,N_5941,N_5913);
or U6689 (N_6689,N_5016,N_6135);
xor U6690 (N_6690,N_6001,N_6156);
nand U6691 (N_6691,N_5892,N_5891);
and U6692 (N_6692,N_5983,N_6007);
and U6693 (N_6693,N_5244,N_6218);
or U6694 (N_6694,N_5976,N_5300);
nor U6695 (N_6695,N_5421,N_5588);
nand U6696 (N_6696,N_5723,N_6013);
or U6697 (N_6697,N_5213,N_5502);
xnor U6698 (N_6698,N_5506,N_5852);
or U6699 (N_6699,N_5793,N_5952);
nor U6700 (N_6700,N_5356,N_5071);
xor U6701 (N_6701,N_5946,N_5452);
and U6702 (N_6702,N_6195,N_5395);
nand U6703 (N_6703,N_6022,N_5720);
xnor U6704 (N_6704,N_5997,N_5771);
nand U6705 (N_6705,N_5510,N_5553);
nand U6706 (N_6706,N_5594,N_5981);
nand U6707 (N_6707,N_5849,N_5303);
xnor U6708 (N_6708,N_5415,N_5881);
nand U6709 (N_6709,N_5217,N_5438);
and U6710 (N_6710,N_5445,N_5214);
and U6711 (N_6711,N_5453,N_6114);
nand U6712 (N_6712,N_5581,N_5730);
xnor U6713 (N_6713,N_5825,N_6014);
nor U6714 (N_6714,N_5132,N_5737);
or U6715 (N_6715,N_5578,N_5786);
nor U6716 (N_6716,N_5349,N_5149);
or U6717 (N_6717,N_5807,N_5675);
nand U6718 (N_6718,N_5799,N_5708);
nor U6719 (N_6719,N_5987,N_5609);
and U6720 (N_6720,N_5954,N_5454);
xnor U6721 (N_6721,N_6017,N_6099);
nor U6722 (N_6722,N_5252,N_5041);
xor U6723 (N_6723,N_5138,N_6028);
or U6724 (N_6724,N_6137,N_5595);
or U6725 (N_6725,N_5889,N_5025);
nor U6726 (N_6726,N_5894,N_5105);
nor U6727 (N_6727,N_5218,N_5872);
and U6728 (N_6728,N_5763,N_5887);
or U6729 (N_6729,N_6052,N_6175);
and U6730 (N_6730,N_5320,N_6006);
xnor U6731 (N_6731,N_5119,N_5462);
xnor U6732 (N_6732,N_5728,N_5154);
and U6733 (N_6733,N_5677,N_6150);
or U6734 (N_6734,N_5036,N_5302);
or U6735 (N_6735,N_5812,N_5229);
or U6736 (N_6736,N_5012,N_5190);
nor U6737 (N_6737,N_5322,N_5391);
and U6738 (N_6738,N_5761,N_5516);
and U6739 (N_6739,N_5823,N_5716);
nand U6740 (N_6740,N_5007,N_5286);
or U6741 (N_6741,N_5602,N_5098);
nor U6742 (N_6742,N_5634,N_5180);
nand U6743 (N_6743,N_5070,N_5900);
nor U6744 (N_6744,N_5332,N_6010);
xnor U6745 (N_6745,N_6185,N_5211);
or U6746 (N_6746,N_5659,N_5911);
xnor U6747 (N_6747,N_6084,N_5188);
and U6748 (N_6748,N_5599,N_5943);
or U6749 (N_6749,N_5151,N_5114);
or U6750 (N_6750,N_5542,N_5663);
nor U6751 (N_6751,N_6189,N_5626);
nor U6752 (N_6752,N_5064,N_5693);
xnor U6753 (N_6753,N_5794,N_5696);
nand U6754 (N_6754,N_5450,N_6069);
nand U6755 (N_6755,N_5493,N_5805);
nor U6756 (N_6756,N_5533,N_5777);
nand U6757 (N_6757,N_5224,N_5126);
nor U6758 (N_6758,N_5073,N_5585);
xnor U6759 (N_6759,N_5604,N_5985);
or U6760 (N_6760,N_6153,N_5243);
xnor U6761 (N_6761,N_5324,N_5964);
xnor U6762 (N_6762,N_5072,N_5163);
xor U6763 (N_6763,N_5713,N_6161);
nand U6764 (N_6764,N_5101,N_5368);
or U6765 (N_6765,N_6050,N_5924);
and U6766 (N_6766,N_5358,N_5388);
or U6767 (N_6767,N_5572,N_5460);
nor U6768 (N_6768,N_6056,N_6192);
nor U6769 (N_6769,N_6026,N_5015);
and U6770 (N_6770,N_5528,N_5026);
xnor U6771 (N_6771,N_5919,N_5543);
xor U6772 (N_6772,N_5291,N_6016);
xor U6773 (N_6773,N_5809,N_5235);
or U6774 (N_6774,N_5766,N_5094);
or U6775 (N_6775,N_5969,N_5111);
or U6776 (N_6776,N_5718,N_5399);
xnor U6777 (N_6777,N_5557,N_5600);
xor U6778 (N_6778,N_6178,N_5055);
nor U6779 (N_6779,N_6140,N_5573);
nor U6780 (N_6780,N_5643,N_5281);
or U6781 (N_6781,N_5563,N_6075);
or U6782 (N_6782,N_5687,N_5222);
or U6783 (N_6783,N_6086,N_5575);
xor U6784 (N_6784,N_5369,N_5196);
or U6785 (N_6785,N_5457,N_5545);
or U6786 (N_6786,N_5464,N_6209);
xor U6787 (N_6787,N_6121,N_5032);
xnor U6788 (N_6788,N_6177,N_5382);
and U6789 (N_6789,N_6132,N_6207);
or U6790 (N_6790,N_5623,N_5005);
nor U6791 (N_6791,N_5948,N_5551);
xor U6792 (N_6792,N_5199,N_5853);
nor U6793 (N_6793,N_5968,N_5133);
and U6794 (N_6794,N_6076,N_5069);
and U6795 (N_6795,N_5255,N_6152);
xnor U6796 (N_6796,N_5167,N_5254);
nand U6797 (N_6797,N_5333,N_5951);
nand U6798 (N_6798,N_5727,N_5505);
or U6799 (N_6799,N_5353,N_6080);
nand U6800 (N_6800,N_5093,N_6021);
xor U6801 (N_6801,N_5507,N_6101);
or U6802 (N_6802,N_5242,N_6097);
or U6803 (N_6803,N_5432,N_5434);
or U6804 (N_6804,N_6232,N_5988);
xor U6805 (N_6805,N_5371,N_5467);
and U6806 (N_6806,N_5605,N_5743);
nand U6807 (N_6807,N_5544,N_5867);
nand U6808 (N_6808,N_5966,N_5652);
xnor U6809 (N_6809,N_5197,N_5042);
or U6810 (N_6810,N_5833,N_5109);
or U6811 (N_6811,N_5993,N_5831);
nor U6812 (N_6812,N_5458,N_5346);
nor U6813 (N_6813,N_6043,N_5503);
nand U6814 (N_6814,N_5960,N_6186);
xnor U6815 (N_6815,N_5439,N_5822);
xnor U6816 (N_6816,N_5292,N_5170);
or U6817 (N_6817,N_5870,N_5967);
nand U6818 (N_6818,N_5790,N_6236);
xnor U6819 (N_6819,N_6045,N_5478);
xor U6820 (N_6820,N_5056,N_5642);
and U6821 (N_6821,N_6053,N_5092);
or U6822 (N_6822,N_5914,N_5760);
nand U6823 (N_6823,N_5681,N_5756);
nor U6824 (N_6824,N_5606,N_5175);
xnor U6825 (N_6825,N_6191,N_5455);
nand U6826 (N_6826,N_5471,N_5702);
and U6827 (N_6827,N_5680,N_5350);
nand U6828 (N_6828,N_5451,N_6233);
nand U6829 (N_6829,N_6107,N_6176);
or U6830 (N_6830,N_5868,N_5674);
xnor U6831 (N_6831,N_6181,N_5047);
or U6832 (N_6832,N_5256,N_6220);
xnor U6833 (N_6833,N_5994,N_5752);
nor U6834 (N_6834,N_5483,N_5145);
or U6835 (N_6835,N_5845,N_5334);
or U6836 (N_6836,N_5917,N_5883);
nor U6837 (N_6837,N_5405,N_5691);
and U6838 (N_6838,N_5389,N_5644);
nand U6839 (N_6839,N_5707,N_5571);
nand U6840 (N_6840,N_6113,N_5820);
or U6841 (N_6841,N_5541,N_5950);
nand U6842 (N_6842,N_5945,N_6139);
and U6843 (N_6843,N_6071,N_5488);
nor U6844 (N_6844,N_5176,N_5999);
and U6845 (N_6845,N_5009,N_5344);
nor U6846 (N_6846,N_5316,N_5898);
or U6847 (N_6847,N_6187,N_5018);
and U6848 (N_6848,N_6066,N_5843);
nor U6849 (N_6849,N_5699,N_5412);
or U6850 (N_6850,N_6060,N_5751);
nor U6851 (N_6851,N_5860,N_6223);
xor U6852 (N_6852,N_5319,N_5341);
nand U6853 (N_6853,N_5684,N_5651);
xor U6854 (N_6854,N_5226,N_5821);
xor U6855 (N_6855,N_5937,N_5147);
or U6856 (N_6856,N_5210,N_5440);
xnor U6857 (N_6857,N_5338,N_5429);
or U6858 (N_6858,N_5125,N_5227);
nand U6859 (N_6859,N_5181,N_5614);
nand U6860 (N_6860,N_5931,N_5657);
nor U6861 (N_6861,N_5112,N_5907);
and U6862 (N_6862,N_5947,N_5904);
xor U6863 (N_6863,N_5798,N_5974);
or U6864 (N_6864,N_6126,N_5504);
xnor U6865 (N_6865,N_5043,N_5744);
or U6866 (N_6866,N_5246,N_5638);
and U6867 (N_6867,N_6079,N_5622);
and U6868 (N_6868,N_5927,N_6127);
nand U6869 (N_6869,N_5275,N_5294);
and U6870 (N_6870,N_6224,N_5789);
xor U6871 (N_6871,N_6219,N_6169);
nand U6872 (N_6872,N_5441,N_5869);
nand U6873 (N_6873,N_6025,N_5374);
and U6874 (N_6874,N_6199,N_5131);
nand U6875 (N_6875,N_5257,N_5463);
or U6876 (N_6876,N_6102,N_5584);
and U6877 (N_6877,N_5572,N_6232);
nor U6878 (N_6878,N_6225,N_5184);
nor U6879 (N_6879,N_5225,N_5752);
nand U6880 (N_6880,N_5551,N_5288);
nor U6881 (N_6881,N_5339,N_5249);
xnor U6882 (N_6882,N_5814,N_6052);
nor U6883 (N_6883,N_6221,N_6106);
xor U6884 (N_6884,N_5056,N_5866);
and U6885 (N_6885,N_5259,N_5841);
nor U6886 (N_6886,N_5952,N_5856);
or U6887 (N_6887,N_5067,N_5813);
xnor U6888 (N_6888,N_5082,N_5198);
or U6889 (N_6889,N_5934,N_5492);
xnor U6890 (N_6890,N_5033,N_5443);
and U6891 (N_6891,N_5834,N_5636);
nor U6892 (N_6892,N_5142,N_5945);
or U6893 (N_6893,N_5678,N_5121);
or U6894 (N_6894,N_5173,N_5347);
nor U6895 (N_6895,N_6042,N_5298);
nor U6896 (N_6896,N_5645,N_5357);
or U6897 (N_6897,N_5099,N_5875);
xor U6898 (N_6898,N_5534,N_5908);
xnor U6899 (N_6899,N_5608,N_5849);
xor U6900 (N_6900,N_5132,N_5144);
xnor U6901 (N_6901,N_5666,N_5406);
nand U6902 (N_6902,N_5105,N_5025);
or U6903 (N_6903,N_5458,N_5817);
or U6904 (N_6904,N_5386,N_5328);
nand U6905 (N_6905,N_5859,N_6233);
nor U6906 (N_6906,N_5250,N_5799);
and U6907 (N_6907,N_6231,N_5575);
and U6908 (N_6908,N_5608,N_5329);
nand U6909 (N_6909,N_5173,N_5969);
and U6910 (N_6910,N_6090,N_6063);
and U6911 (N_6911,N_5097,N_5905);
xor U6912 (N_6912,N_5906,N_5976);
nand U6913 (N_6913,N_5686,N_6101);
nand U6914 (N_6914,N_5858,N_5596);
nand U6915 (N_6915,N_5942,N_5592);
nand U6916 (N_6916,N_5321,N_5128);
xnor U6917 (N_6917,N_5200,N_5165);
xor U6918 (N_6918,N_5384,N_5900);
xnor U6919 (N_6919,N_5485,N_5738);
or U6920 (N_6920,N_5898,N_6030);
xor U6921 (N_6921,N_5805,N_5458);
nor U6922 (N_6922,N_6209,N_5637);
nand U6923 (N_6923,N_5164,N_5716);
xor U6924 (N_6924,N_5223,N_5414);
nand U6925 (N_6925,N_5313,N_5574);
nand U6926 (N_6926,N_5208,N_5062);
and U6927 (N_6927,N_5871,N_5620);
and U6928 (N_6928,N_5333,N_5709);
nand U6929 (N_6929,N_5328,N_5559);
and U6930 (N_6930,N_5652,N_6063);
nor U6931 (N_6931,N_6128,N_5951);
or U6932 (N_6932,N_5050,N_5109);
xnor U6933 (N_6933,N_5882,N_5448);
or U6934 (N_6934,N_5989,N_5322);
xnor U6935 (N_6935,N_5151,N_5474);
and U6936 (N_6936,N_5899,N_5780);
or U6937 (N_6937,N_5818,N_6121);
xnor U6938 (N_6938,N_5319,N_5014);
nand U6939 (N_6939,N_5019,N_5302);
nand U6940 (N_6940,N_5584,N_5702);
or U6941 (N_6941,N_5655,N_5312);
xor U6942 (N_6942,N_6073,N_6019);
xnor U6943 (N_6943,N_5031,N_5825);
nor U6944 (N_6944,N_5293,N_6105);
or U6945 (N_6945,N_6000,N_5812);
and U6946 (N_6946,N_5867,N_5235);
and U6947 (N_6947,N_5274,N_5008);
nor U6948 (N_6948,N_5419,N_5458);
xor U6949 (N_6949,N_5396,N_5599);
and U6950 (N_6950,N_5319,N_5730);
nand U6951 (N_6951,N_5256,N_5551);
and U6952 (N_6952,N_5688,N_5001);
and U6953 (N_6953,N_6063,N_5664);
nand U6954 (N_6954,N_5832,N_5007);
or U6955 (N_6955,N_5241,N_6096);
nor U6956 (N_6956,N_5203,N_5488);
nand U6957 (N_6957,N_6112,N_5630);
nand U6958 (N_6958,N_5556,N_5051);
nand U6959 (N_6959,N_5044,N_5100);
or U6960 (N_6960,N_5003,N_5355);
and U6961 (N_6961,N_5794,N_5214);
xnor U6962 (N_6962,N_5431,N_6090);
nor U6963 (N_6963,N_5519,N_5242);
or U6964 (N_6964,N_5966,N_5717);
or U6965 (N_6965,N_5226,N_5290);
nand U6966 (N_6966,N_5575,N_5067);
nand U6967 (N_6967,N_5162,N_5111);
nor U6968 (N_6968,N_5441,N_6055);
nor U6969 (N_6969,N_5299,N_5391);
or U6970 (N_6970,N_5760,N_6200);
xnor U6971 (N_6971,N_5307,N_5071);
or U6972 (N_6972,N_5122,N_5294);
or U6973 (N_6973,N_6146,N_5622);
nor U6974 (N_6974,N_5956,N_5415);
and U6975 (N_6975,N_5305,N_5593);
or U6976 (N_6976,N_6047,N_5734);
xnor U6977 (N_6977,N_5152,N_5178);
and U6978 (N_6978,N_5507,N_5386);
xnor U6979 (N_6979,N_5880,N_5077);
or U6980 (N_6980,N_5472,N_6011);
nor U6981 (N_6981,N_5829,N_5339);
nor U6982 (N_6982,N_5361,N_5951);
and U6983 (N_6983,N_5814,N_5832);
nand U6984 (N_6984,N_5891,N_5543);
nand U6985 (N_6985,N_5240,N_5571);
xor U6986 (N_6986,N_5094,N_5866);
nand U6987 (N_6987,N_6106,N_5220);
nand U6988 (N_6988,N_5266,N_5550);
nor U6989 (N_6989,N_5408,N_6066);
nor U6990 (N_6990,N_5766,N_5146);
and U6991 (N_6991,N_5250,N_5300);
or U6992 (N_6992,N_5625,N_5964);
nor U6993 (N_6993,N_5783,N_6151);
nor U6994 (N_6994,N_5748,N_5303);
xor U6995 (N_6995,N_5460,N_5439);
and U6996 (N_6996,N_5615,N_5995);
or U6997 (N_6997,N_5203,N_5550);
xnor U6998 (N_6998,N_5293,N_5411);
or U6999 (N_6999,N_5291,N_5755);
and U7000 (N_7000,N_5921,N_5752);
nor U7001 (N_7001,N_5301,N_5510);
or U7002 (N_7002,N_5156,N_6233);
or U7003 (N_7003,N_5558,N_5781);
nor U7004 (N_7004,N_5210,N_6117);
nor U7005 (N_7005,N_5263,N_5722);
nand U7006 (N_7006,N_5683,N_5123);
or U7007 (N_7007,N_5148,N_5769);
nor U7008 (N_7008,N_6054,N_5673);
nand U7009 (N_7009,N_5545,N_5989);
xor U7010 (N_7010,N_5265,N_5088);
or U7011 (N_7011,N_5253,N_5783);
xnor U7012 (N_7012,N_5067,N_5326);
nand U7013 (N_7013,N_6123,N_6046);
nand U7014 (N_7014,N_6093,N_6040);
nand U7015 (N_7015,N_5243,N_5800);
or U7016 (N_7016,N_5974,N_5384);
nand U7017 (N_7017,N_5473,N_5677);
nand U7018 (N_7018,N_5469,N_5699);
nor U7019 (N_7019,N_5467,N_5873);
and U7020 (N_7020,N_5802,N_6086);
xnor U7021 (N_7021,N_6123,N_5412);
xnor U7022 (N_7022,N_5277,N_5090);
xnor U7023 (N_7023,N_5895,N_5990);
xor U7024 (N_7024,N_5394,N_5460);
nand U7025 (N_7025,N_5173,N_5081);
or U7026 (N_7026,N_5124,N_5625);
or U7027 (N_7027,N_5346,N_5233);
and U7028 (N_7028,N_5524,N_6203);
or U7029 (N_7029,N_5629,N_6145);
nand U7030 (N_7030,N_5881,N_5494);
and U7031 (N_7031,N_5344,N_6123);
nor U7032 (N_7032,N_5079,N_6056);
and U7033 (N_7033,N_5425,N_5609);
and U7034 (N_7034,N_5120,N_5333);
xor U7035 (N_7035,N_5970,N_5841);
or U7036 (N_7036,N_6188,N_5491);
and U7037 (N_7037,N_6166,N_5219);
and U7038 (N_7038,N_6058,N_5631);
or U7039 (N_7039,N_5195,N_5505);
or U7040 (N_7040,N_5542,N_5813);
or U7041 (N_7041,N_5081,N_6001);
and U7042 (N_7042,N_6073,N_6228);
nor U7043 (N_7043,N_5047,N_5094);
or U7044 (N_7044,N_5478,N_5088);
nand U7045 (N_7045,N_5836,N_5173);
xor U7046 (N_7046,N_5237,N_5349);
or U7047 (N_7047,N_5168,N_5143);
nor U7048 (N_7048,N_5873,N_5697);
xnor U7049 (N_7049,N_5306,N_5659);
nand U7050 (N_7050,N_5795,N_5966);
and U7051 (N_7051,N_5593,N_5860);
or U7052 (N_7052,N_5355,N_5153);
or U7053 (N_7053,N_5075,N_5513);
xnor U7054 (N_7054,N_5999,N_5843);
or U7055 (N_7055,N_5538,N_5918);
xor U7056 (N_7056,N_5379,N_5018);
nor U7057 (N_7057,N_6159,N_5906);
or U7058 (N_7058,N_5989,N_6020);
and U7059 (N_7059,N_5595,N_5087);
or U7060 (N_7060,N_5518,N_5369);
nand U7061 (N_7061,N_6140,N_5327);
xnor U7062 (N_7062,N_5740,N_5915);
nor U7063 (N_7063,N_5463,N_5279);
and U7064 (N_7064,N_5233,N_5662);
nand U7065 (N_7065,N_5966,N_5353);
xor U7066 (N_7066,N_5448,N_6046);
nor U7067 (N_7067,N_5875,N_5462);
or U7068 (N_7068,N_6236,N_5000);
or U7069 (N_7069,N_6184,N_5502);
nor U7070 (N_7070,N_5868,N_6186);
xor U7071 (N_7071,N_5814,N_6002);
nor U7072 (N_7072,N_5253,N_5355);
and U7073 (N_7073,N_5230,N_5981);
or U7074 (N_7074,N_5250,N_5099);
or U7075 (N_7075,N_5721,N_5629);
or U7076 (N_7076,N_6184,N_6180);
or U7077 (N_7077,N_5691,N_5754);
nor U7078 (N_7078,N_5010,N_5360);
or U7079 (N_7079,N_5717,N_5972);
and U7080 (N_7080,N_5514,N_5116);
xnor U7081 (N_7081,N_6013,N_5463);
xnor U7082 (N_7082,N_5786,N_5525);
nor U7083 (N_7083,N_5758,N_5890);
nor U7084 (N_7084,N_5976,N_6156);
and U7085 (N_7085,N_6181,N_6203);
or U7086 (N_7086,N_5655,N_5054);
or U7087 (N_7087,N_6169,N_5685);
and U7088 (N_7088,N_5829,N_5895);
xor U7089 (N_7089,N_5384,N_6039);
nor U7090 (N_7090,N_5996,N_6127);
nand U7091 (N_7091,N_5987,N_6053);
and U7092 (N_7092,N_5644,N_5193);
nor U7093 (N_7093,N_5221,N_5724);
xor U7094 (N_7094,N_5561,N_6022);
or U7095 (N_7095,N_5781,N_5172);
nand U7096 (N_7096,N_6095,N_5021);
nor U7097 (N_7097,N_5538,N_6023);
xnor U7098 (N_7098,N_6182,N_5035);
xnor U7099 (N_7099,N_5310,N_5510);
xnor U7100 (N_7100,N_5048,N_5073);
nand U7101 (N_7101,N_5396,N_5186);
or U7102 (N_7102,N_5792,N_5190);
and U7103 (N_7103,N_5418,N_5414);
nor U7104 (N_7104,N_5060,N_5007);
nor U7105 (N_7105,N_5374,N_5707);
or U7106 (N_7106,N_5850,N_5255);
nor U7107 (N_7107,N_5383,N_5200);
or U7108 (N_7108,N_6101,N_6074);
xnor U7109 (N_7109,N_5556,N_5454);
nor U7110 (N_7110,N_5517,N_6056);
xor U7111 (N_7111,N_6164,N_5591);
nand U7112 (N_7112,N_5846,N_6053);
or U7113 (N_7113,N_6162,N_5855);
and U7114 (N_7114,N_6030,N_6183);
xor U7115 (N_7115,N_5285,N_5935);
xnor U7116 (N_7116,N_5554,N_5120);
xor U7117 (N_7117,N_5594,N_5361);
nor U7118 (N_7118,N_5283,N_6058);
or U7119 (N_7119,N_6205,N_5438);
nor U7120 (N_7120,N_5670,N_5394);
or U7121 (N_7121,N_5427,N_5092);
nand U7122 (N_7122,N_5183,N_5090);
and U7123 (N_7123,N_6183,N_5495);
nor U7124 (N_7124,N_6211,N_5428);
nand U7125 (N_7125,N_5283,N_5615);
nand U7126 (N_7126,N_5983,N_5954);
xnor U7127 (N_7127,N_5174,N_5611);
nand U7128 (N_7128,N_5027,N_5071);
nor U7129 (N_7129,N_5171,N_6056);
nor U7130 (N_7130,N_5992,N_5943);
nor U7131 (N_7131,N_5593,N_5040);
and U7132 (N_7132,N_5662,N_5294);
and U7133 (N_7133,N_5115,N_5515);
or U7134 (N_7134,N_5372,N_5396);
or U7135 (N_7135,N_5635,N_5538);
xor U7136 (N_7136,N_5903,N_5515);
xor U7137 (N_7137,N_6009,N_6106);
and U7138 (N_7138,N_6065,N_5956);
or U7139 (N_7139,N_6056,N_5984);
or U7140 (N_7140,N_5180,N_5297);
nor U7141 (N_7141,N_5191,N_5554);
xor U7142 (N_7142,N_5503,N_5427);
and U7143 (N_7143,N_5187,N_5331);
or U7144 (N_7144,N_5498,N_6170);
or U7145 (N_7145,N_5411,N_5831);
and U7146 (N_7146,N_5091,N_5561);
or U7147 (N_7147,N_5691,N_5482);
xor U7148 (N_7148,N_5324,N_5587);
nand U7149 (N_7149,N_5965,N_5199);
xnor U7150 (N_7150,N_5762,N_5907);
and U7151 (N_7151,N_5012,N_5215);
nand U7152 (N_7152,N_5920,N_6169);
xor U7153 (N_7153,N_5194,N_5708);
or U7154 (N_7154,N_6095,N_5195);
or U7155 (N_7155,N_5546,N_5203);
xnor U7156 (N_7156,N_5704,N_5057);
or U7157 (N_7157,N_5938,N_5244);
or U7158 (N_7158,N_5297,N_6149);
or U7159 (N_7159,N_5247,N_5367);
nand U7160 (N_7160,N_6208,N_5171);
xnor U7161 (N_7161,N_6217,N_5707);
or U7162 (N_7162,N_6074,N_5259);
xor U7163 (N_7163,N_6193,N_5687);
xnor U7164 (N_7164,N_5051,N_5950);
nor U7165 (N_7165,N_5643,N_5181);
and U7166 (N_7166,N_5175,N_5060);
or U7167 (N_7167,N_6052,N_5952);
nor U7168 (N_7168,N_5809,N_5670);
xor U7169 (N_7169,N_6152,N_5674);
nand U7170 (N_7170,N_5228,N_6122);
nor U7171 (N_7171,N_5891,N_5508);
nor U7172 (N_7172,N_5919,N_6004);
nor U7173 (N_7173,N_5670,N_5117);
or U7174 (N_7174,N_6230,N_6068);
nor U7175 (N_7175,N_5885,N_5221);
and U7176 (N_7176,N_6109,N_5167);
xor U7177 (N_7177,N_5183,N_5843);
xnor U7178 (N_7178,N_6113,N_6241);
nand U7179 (N_7179,N_6061,N_6032);
xnor U7180 (N_7180,N_5896,N_5874);
xnor U7181 (N_7181,N_5776,N_5639);
nor U7182 (N_7182,N_5248,N_5770);
or U7183 (N_7183,N_5944,N_5472);
nand U7184 (N_7184,N_5969,N_5424);
nand U7185 (N_7185,N_6091,N_5248);
nand U7186 (N_7186,N_5680,N_5693);
nand U7187 (N_7187,N_5022,N_5187);
xnor U7188 (N_7188,N_5195,N_6133);
and U7189 (N_7189,N_5585,N_5866);
and U7190 (N_7190,N_6016,N_5227);
or U7191 (N_7191,N_6225,N_5277);
or U7192 (N_7192,N_5294,N_6064);
or U7193 (N_7193,N_5181,N_5501);
nor U7194 (N_7194,N_6109,N_6037);
or U7195 (N_7195,N_5903,N_5143);
nor U7196 (N_7196,N_6053,N_5803);
nand U7197 (N_7197,N_5442,N_5363);
and U7198 (N_7198,N_5354,N_5800);
or U7199 (N_7199,N_6078,N_5611);
and U7200 (N_7200,N_5352,N_5426);
nand U7201 (N_7201,N_5041,N_5651);
nand U7202 (N_7202,N_5164,N_6201);
nor U7203 (N_7203,N_5189,N_5028);
nor U7204 (N_7204,N_5864,N_5942);
and U7205 (N_7205,N_5236,N_5693);
nand U7206 (N_7206,N_5354,N_5507);
and U7207 (N_7207,N_5819,N_5903);
xnor U7208 (N_7208,N_5011,N_5180);
and U7209 (N_7209,N_5923,N_5679);
nor U7210 (N_7210,N_5605,N_5515);
nand U7211 (N_7211,N_5005,N_5579);
xnor U7212 (N_7212,N_5608,N_5475);
and U7213 (N_7213,N_6041,N_5175);
nand U7214 (N_7214,N_5603,N_5558);
or U7215 (N_7215,N_6100,N_5052);
and U7216 (N_7216,N_5021,N_5319);
xor U7217 (N_7217,N_6034,N_5790);
or U7218 (N_7218,N_5939,N_5021);
nor U7219 (N_7219,N_5382,N_6063);
nor U7220 (N_7220,N_5785,N_5039);
and U7221 (N_7221,N_5868,N_5214);
and U7222 (N_7222,N_6214,N_5853);
and U7223 (N_7223,N_5728,N_5606);
nor U7224 (N_7224,N_5905,N_6162);
and U7225 (N_7225,N_5276,N_5979);
or U7226 (N_7226,N_5429,N_5079);
nand U7227 (N_7227,N_5186,N_5928);
nor U7228 (N_7228,N_5016,N_5072);
or U7229 (N_7229,N_5183,N_5635);
nand U7230 (N_7230,N_6215,N_5840);
xor U7231 (N_7231,N_5636,N_6035);
xnor U7232 (N_7232,N_5104,N_5089);
nand U7233 (N_7233,N_5686,N_5307);
xor U7234 (N_7234,N_5285,N_5642);
nand U7235 (N_7235,N_5958,N_5455);
xnor U7236 (N_7236,N_5178,N_5737);
nand U7237 (N_7237,N_5214,N_6080);
nand U7238 (N_7238,N_5829,N_5496);
nand U7239 (N_7239,N_5134,N_6116);
nor U7240 (N_7240,N_5045,N_6015);
and U7241 (N_7241,N_5227,N_5875);
nor U7242 (N_7242,N_5441,N_5726);
or U7243 (N_7243,N_5534,N_5213);
nand U7244 (N_7244,N_5237,N_5574);
nand U7245 (N_7245,N_5499,N_5143);
nor U7246 (N_7246,N_5714,N_5138);
or U7247 (N_7247,N_5716,N_5339);
nor U7248 (N_7248,N_5659,N_6203);
xor U7249 (N_7249,N_5591,N_5518);
and U7250 (N_7250,N_5550,N_6001);
xor U7251 (N_7251,N_6076,N_6112);
nor U7252 (N_7252,N_6082,N_5359);
nand U7253 (N_7253,N_5217,N_5960);
or U7254 (N_7254,N_5386,N_5809);
and U7255 (N_7255,N_5793,N_5751);
or U7256 (N_7256,N_5790,N_5439);
xor U7257 (N_7257,N_5541,N_5712);
or U7258 (N_7258,N_5979,N_5700);
and U7259 (N_7259,N_6246,N_5844);
and U7260 (N_7260,N_5659,N_5913);
and U7261 (N_7261,N_5381,N_5289);
nand U7262 (N_7262,N_5754,N_5683);
nor U7263 (N_7263,N_5742,N_5716);
xor U7264 (N_7264,N_5204,N_5732);
nor U7265 (N_7265,N_5498,N_5373);
nor U7266 (N_7266,N_5722,N_5961);
nand U7267 (N_7267,N_6042,N_5982);
or U7268 (N_7268,N_6156,N_5371);
nor U7269 (N_7269,N_5180,N_5878);
and U7270 (N_7270,N_5982,N_5155);
or U7271 (N_7271,N_5728,N_5364);
nor U7272 (N_7272,N_5909,N_5819);
or U7273 (N_7273,N_5885,N_5029);
and U7274 (N_7274,N_6174,N_5523);
xnor U7275 (N_7275,N_5073,N_6075);
nand U7276 (N_7276,N_5242,N_5629);
nand U7277 (N_7277,N_5837,N_5008);
or U7278 (N_7278,N_5175,N_5401);
and U7279 (N_7279,N_5458,N_5095);
nand U7280 (N_7280,N_5721,N_6038);
nand U7281 (N_7281,N_6057,N_5893);
and U7282 (N_7282,N_5566,N_6053);
xor U7283 (N_7283,N_5327,N_5055);
or U7284 (N_7284,N_5779,N_5801);
or U7285 (N_7285,N_6124,N_5892);
nor U7286 (N_7286,N_5565,N_5189);
nand U7287 (N_7287,N_5551,N_6248);
or U7288 (N_7288,N_5142,N_5689);
and U7289 (N_7289,N_5348,N_6104);
or U7290 (N_7290,N_5514,N_5710);
nand U7291 (N_7291,N_6049,N_5561);
nor U7292 (N_7292,N_5278,N_5095);
nand U7293 (N_7293,N_6166,N_5617);
nor U7294 (N_7294,N_5007,N_5880);
and U7295 (N_7295,N_5337,N_5799);
xor U7296 (N_7296,N_5430,N_6125);
or U7297 (N_7297,N_6012,N_5131);
and U7298 (N_7298,N_5720,N_5749);
nand U7299 (N_7299,N_5666,N_5307);
or U7300 (N_7300,N_5521,N_6064);
and U7301 (N_7301,N_5744,N_6205);
and U7302 (N_7302,N_5781,N_5550);
nor U7303 (N_7303,N_6218,N_5090);
nand U7304 (N_7304,N_5985,N_5021);
xor U7305 (N_7305,N_6202,N_5829);
xor U7306 (N_7306,N_5173,N_5046);
nor U7307 (N_7307,N_6115,N_5806);
nor U7308 (N_7308,N_5269,N_6206);
nand U7309 (N_7309,N_6138,N_5772);
or U7310 (N_7310,N_5989,N_5953);
or U7311 (N_7311,N_5591,N_5377);
nor U7312 (N_7312,N_5009,N_5124);
or U7313 (N_7313,N_6187,N_5518);
nor U7314 (N_7314,N_5098,N_5999);
nor U7315 (N_7315,N_6200,N_5867);
and U7316 (N_7316,N_5541,N_5228);
nand U7317 (N_7317,N_5232,N_5222);
and U7318 (N_7318,N_5675,N_5192);
nand U7319 (N_7319,N_5791,N_5666);
xnor U7320 (N_7320,N_6129,N_5762);
xor U7321 (N_7321,N_5909,N_5688);
or U7322 (N_7322,N_5170,N_6140);
and U7323 (N_7323,N_6142,N_5273);
and U7324 (N_7324,N_5147,N_6135);
nand U7325 (N_7325,N_5735,N_5437);
xor U7326 (N_7326,N_5748,N_5581);
nand U7327 (N_7327,N_5348,N_5557);
xnor U7328 (N_7328,N_6201,N_5239);
or U7329 (N_7329,N_5521,N_6161);
nand U7330 (N_7330,N_5847,N_5872);
or U7331 (N_7331,N_6003,N_5394);
and U7332 (N_7332,N_5026,N_5272);
or U7333 (N_7333,N_5327,N_5248);
and U7334 (N_7334,N_5724,N_6034);
nand U7335 (N_7335,N_5418,N_6222);
nand U7336 (N_7336,N_5438,N_5781);
and U7337 (N_7337,N_5385,N_6235);
and U7338 (N_7338,N_5664,N_5930);
nor U7339 (N_7339,N_5751,N_5035);
xor U7340 (N_7340,N_5570,N_5171);
nand U7341 (N_7341,N_5621,N_5701);
xnor U7342 (N_7342,N_5902,N_6238);
xnor U7343 (N_7343,N_5592,N_5822);
nor U7344 (N_7344,N_5292,N_5766);
or U7345 (N_7345,N_5467,N_6020);
nor U7346 (N_7346,N_6175,N_5479);
xnor U7347 (N_7347,N_5405,N_5006);
or U7348 (N_7348,N_5833,N_5068);
nor U7349 (N_7349,N_5949,N_5030);
or U7350 (N_7350,N_5510,N_5813);
and U7351 (N_7351,N_5675,N_6166);
nor U7352 (N_7352,N_5258,N_5896);
or U7353 (N_7353,N_5384,N_5110);
xor U7354 (N_7354,N_5168,N_5636);
and U7355 (N_7355,N_5802,N_6249);
or U7356 (N_7356,N_5546,N_6124);
or U7357 (N_7357,N_5821,N_5425);
and U7358 (N_7358,N_5811,N_5460);
and U7359 (N_7359,N_6188,N_6248);
xnor U7360 (N_7360,N_6240,N_5343);
or U7361 (N_7361,N_5008,N_5515);
or U7362 (N_7362,N_5173,N_5472);
nor U7363 (N_7363,N_5816,N_6237);
nand U7364 (N_7364,N_5039,N_5409);
xnor U7365 (N_7365,N_5974,N_5467);
xnor U7366 (N_7366,N_5235,N_5573);
or U7367 (N_7367,N_5490,N_5031);
xnor U7368 (N_7368,N_5418,N_5179);
and U7369 (N_7369,N_5706,N_5243);
xor U7370 (N_7370,N_5766,N_5633);
xor U7371 (N_7371,N_5659,N_5115);
or U7372 (N_7372,N_5063,N_5504);
and U7373 (N_7373,N_5679,N_5881);
and U7374 (N_7374,N_5606,N_5862);
and U7375 (N_7375,N_6064,N_6214);
or U7376 (N_7376,N_5658,N_5494);
nor U7377 (N_7377,N_5873,N_5874);
nor U7378 (N_7378,N_5718,N_5063);
and U7379 (N_7379,N_5189,N_5514);
or U7380 (N_7380,N_6227,N_5513);
and U7381 (N_7381,N_5426,N_5325);
xor U7382 (N_7382,N_5890,N_5505);
and U7383 (N_7383,N_5452,N_5297);
nor U7384 (N_7384,N_5959,N_6177);
or U7385 (N_7385,N_5352,N_5564);
xor U7386 (N_7386,N_5893,N_5824);
xnor U7387 (N_7387,N_5332,N_5744);
or U7388 (N_7388,N_5757,N_5093);
or U7389 (N_7389,N_5336,N_5903);
nand U7390 (N_7390,N_5532,N_5600);
xor U7391 (N_7391,N_5785,N_5388);
xnor U7392 (N_7392,N_5964,N_5928);
or U7393 (N_7393,N_6102,N_5152);
and U7394 (N_7394,N_5379,N_6108);
nand U7395 (N_7395,N_5164,N_5351);
or U7396 (N_7396,N_5041,N_6047);
nor U7397 (N_7397,N_5249,N_5039);
and U7398 (N_7398,N_5783,N_5405);
xnor U7399 (N_7399,N_6144,N_5992);
xnor U7400 (N_7400,N_5506,N_5703);
xor U7401 (N_7401,N_5792,N_5907);
or U7402 (N_7402,N_5412,N_5090);
xnor U7403 (N_7403,N_5599,N_5486);
nor U7404 (N_7404,N_5702,N_6121);
xor U7405 (N_7405,N_6010,N_5550);
xor U7406 (N_7406,N_5818,N_5659);
or U7407 (N_7407,N_5997,N_5396);
and U7408 (N_7408,N_5378,N_5606);
and U7409 (N_7409,N_6151,N_6079);
and U7410 (N_7410,N_5482,N_5392);
and U7411 (N_7411,N_5829,N_5762);
and U7412 (N_7412,N_6179,N_5817);
xnor U7413 (N_7413,N_6119,N_5244);
nand U7414 (N_7414,N_5716,N_5039);
or U7415 (N_7415,N_5492,N_6045);
and U7416 (N_7416,N_5127,N_5926);
or U7417 (N_7417,N_5819,N_5006);
and U7418 (N_7418,N_5239,N_5914);
nand U7419 (N_7419,N_6214,N_5500);
xor U7420 (N_7420,N_5375,N_5553);
or U7421 (N_7421,N_5907,N_5820);
nand U7422 (N_7422,N_5375,N_5126);
nand U7423 (N_7423,N_5130,N_5978);
nor U7424 (N_7424,N_5915,N_6214);
or U7425 (N_7425,N_5921,N_5227);
nor U7426 (N_7426,N_6115,N_5121);
xor U7427 (N_7427,N_5603,N_6110);
or U7428 (N_7428,N_5048,N_6092);
nor U7429 (N_7429,N_5009,N_5651);
or U7430 (N_7430,N_5027,N_6173);
and U7431 (N_7431,N_5856,N_5649);
xnor U7432 (N_7432,N_6187,N_5537);
nand U7433 (N_7433,N_5422,N_6208);
xor U7434 (N_7434,N_6011,N_5138);
and U7435 (N_7435,N_5885,N_5821);
and U7436 (N_7436,N_5628,N_5697);
nand U7437 (N_7437,N_6248,N_6124);
or U7438 (N_7438,N_5837,N_5055);
nor U7439 (N_7439,N_5758,N_5755);
and U7440 (N_7440,N_6233,N_5698);
or U7441 (N_7441,N_5800,N_5944);
xor U7442 (N_7442,N_5158,N_5808);
nor U7443 (N_7443,N_5047,N_5739);
xor U7444 (N_7444,N_5856,N_5965);
nand U7445 (N_7445,N_5292,N_5555);
xor U7446 (N_7446,N_5175,N_6241);
nor U7447 (N_7447,N_5310,N_5678);
nand U7448 (N_7448,N_5902,N_5935);
nor U7449 (N_7449,N_5631,N_5825);
nor U7450 (N_7450,N_6016,N_5092);
nand U7451 (N_7451,N_5795,N_5209);
nor U7452 (N_7452,N_5215,N_5869);
xor U7453 (N_7453,N_6222,N_5195);
and U7454 (N_7454,N_5284,N_5822);
xor U7455 (N_7455,N_5226,N_6150);
xor U7456 (N_7456,N_5988,N_5612);
xor U7457 (N_7457,N_5799,N_5394);
xor U7458 (N_7458,N_5301,N_5284);
nor U7459 (N_7459,N_5757,N_5900);
nand U7460 (N_7460,N_5070,N_5890);
xnor U7461 (N_7461,N_5923,N_6246);
or U7462 (N_7462,N_5674,N_5240);
xnor U7463 (N_7463,N_5709,N_5543);
or U7464 (N_7464,N_6013,N_6133);
nand U7465 (N_7465,N_5414,N_5728);
nand U7466 (N_7466,N_5820,N_5421);
and U7467 (N_7467,N_5112,N_5288);
nand U7468 (N_7468,N_6096,N_5588);
nor U7469 (N_7469,N_5481,N_5301);
nor U7470 (N_7470,N_5588,N_5067);
and U7471 (N_7471,N_6081,N_5107);
nand U7472 (N_7472,N_5134,N_5505);
xor U7473 (N_7473,N_6010,N_6006);
nand U7474 (N_7474,N_5515,N_5644);
nor U7475 (N_7475,N_6117,N_5725);
nand U7476 (N_7476,N_6096,N_5160);
xnor U7477 (N_7477,N_5458,N_6176);
and U7478 (N_7478,N_5059,N_5001);
nor U7479 (N_7479,N_5386,N_5497);
and U7480 (N_7480,N_5409,N_5757);
nor U7481 (N_7481,N_5557,N_5972);
nand U7482 (N_7482,N_6084,N_5272);
xnor U7483 (N_7483,N_5282,N_5155);
or U7484 (N_7484,N_5042,N_6154);
nand U7485 (N_7485,N_5723,N_5042);
and U7486 (N_7486,N_6182,N_5021);
nand U7487 (N_7487,N_5031,N_5964);
xor U7488 (N_7488,N_6214,N_5504);
and U7489 (N_7489,N_5909,N_5194);
nor U7490 (N_7490,N_5657,N_5493);
or U7491 (N_7491,N_5353,N_5357);
nand U7492 (N_7492,N_5868,N_6218);
nor U7493 (N_7493,N_5147,N_5003);
nand U7494 (N_7494,N_5994,N_5704);
and U7495 (N_7495,N_5420,N_6098);
xnor U7496 (N_7496,N_6117,N_5653);
xor U7497 (N_7497,N_5914,N_5365);
nand U7498 (N_7498,N_6038,N_5109);
nand U7499 (N_7499,N_5576,N_5328);
nand U7500 (N_7500,N_6448,N_7335);
and U7501 (N_7501,N_6833,N_6955);
nand U7502 (N_7502,N_6436,N_6495);
and U7503 (N_7503,N_7365,N_7491);
and U7504 (N_7504,N_6513,N_6980);
and U7505 (N_7505,N_7148,N_6873);
and U7506 (N_7506,N_6523,N_6874);
and U7507 (N_7507,N_7159,N_7102);
and U7508 (N_7508,N_6332,N_6838);
or U7509 (N_7509,N_7453,N_6530);
nor U7510 (N_7510,N_6649,N_6573);
xnor U7511 (N_7511,N_6345,N_6386);
or U7512 (N_7512,N_7441,N_6628);
or U7513 (N_7513,N_6420,N_7448);
nand U7514 (N_7514,N_6677,N_6443);
and U7515 (N_7515,N_6991,N_6477);
nand U7516 (N_7516,N_7112,N_7161);
or U7517 (N_7517,N_6293,N_7191);
and U7518 (N_7518,N_6383,N_7154);
nand U7519 (N_7519,N_6840,N_6913);
xor U7520 (N_7520,N_6887,N_6276);
nand U7521 (N_7521,N_7361,N_6426);
or U7522 (N_7522,N_6446,N_7036);
or U7523 (N_7523,N_6544,N_7027);
nand U7524 (N_7524,N_6532,N_7046);
nand U7525 (N_7525,N_7236,N_6300);
or U7526 (N_7526,N_6954,N_7196);
xnor U7527 (N_7527,N_6527,N_7095);
nor U7528 (N_7528,N_7397,N_6583);
or U7529 (N_7529,N_6503,N_7401);
or U7530 (N_7530,N_6995,N_7028);
xor U7531 (N_7531,N_6459,N_6491);
or U7532 (N_7532,N_7208,N_6964);
nand U7533 (N_7533,N_6558,N_6469);
or U7534 (N_7534,N_6851,N_6546);
xnor U7535 (N_7535,N_7319,N_6509);
or U7536 (N_7536,N_6591,N_6794);
or U7537 (N_7537,N_7187,N_6261);
nor U7538 (N_7538,N_6805,N_7143);
nor U7539 (N_7539,N_7141,N_7050);
xnor U7540 (N_7540,N_7293,N_6801);
xor U7541 (N_7541,N_7091,N_7416);
nor U7542 (N_7542,N_7472,N_6368);
xor U7543 (N_7543,N_6565,N_6941);
and U7544 (N_7544,N_6808,N_6882);
nand U7545 (N_7545,N_7287,N_6594);
or U7546 (N_7546,N_7254,N_6722);
nor U7547 (N_7547,N_6250,N_7226);
nor U7548 (N_7548,N_6827,N_6900);
nor U7549 (N_7549,N_7192,N_6639);
or U7550 (N_7550,N_7211,N_6770);
xnor U7551 (N_7551,N_6800,N_6487);
and U7552 (N_7552,N_6907,N_6608);
nor U7553 (N_7553,N_7151,N_6298);
and U7554 (N_7554,N_6986,N_6415);
or U7555 (N_7555,N_6408,N_6549);
xnor U7556 (N_7556,N_7436,N_7123);
xor U7557 (N_7557,N_6665,N_6783);
nand U7558 (N_7558,N_6971,N_7233);
xor U7559 (N_7559,N_7284,N_6668);
and U7560 (N_7560,N_6488,N_6835);
nand U7561 (N_7561,N_7173,N_7381);
and U7562 (N_7562,N_6437,N_7322);
nor U7563 (N_7563,N_6557,N_7043);
or U7564 (N_7564,N_6274,N_6921);
xor U7565 (N_7565,N_6550,N_6645);
xnor U7566 (N_7566,N_7337,N_6790);
and U7567 (N_7567,N_6650,N_7186);
xnor U7568 (N_7568,N_6708,N_7145);
and U7569 (N_7569,N_6581,N_6410);
and U7570 (N_7570,N_6864,N_7498);
or U7571 (N_7571,N_7304,N_6598);
or U7572 (N_7572,N_6881,N_7177);
and U7573 (N_7573,N_6868,N_6296);
nand U7574 (N_7574,N_6723,N_6924);
xor U7575 (N_7575,N_7008,N_6754);
nor U7576 (N_7576,N_6388,N_7240);
and U7577 (N_7577,N_7132,N_7446);
nand U7578 (N_7578,N_7331,N_7262);
and U7579 (N_7579,N_7190,N_6387);
nand U7580 (N_7580,N_7496,N_6475);
nand U7581 (N_7581,N_6484,N_7332);
xnor U7582 (N_7582,N_6958,N_7134);
xnor U7583 (N_7583,N_7185,N_7158);
xor U7584 (N_7584,N_7367,N_6713);
and U7585 (N_7585,N_6444,N_6641);
nand U7586 (N_7586,N_6592,N_7386);
nor U7587 (N_7587,N_6675,N_6901);
xnor U7588 (N_7588,N_6572,N_7355);
nand U7589 (N_7589,N_6452,N_6328);
nand U7590 (N_7590,N_6430,N_7181);
nand U7591 (N_7591,N_6866,N_7370);
xnor U7592 (N_7592,N_7379,N_7302);
nand U7593 (N_7593,N_6306,N_7020);
nand U7594 (N_7594,N_7189,N_7051);
or U7595 (N_7595,N_7395,N_6962);
and U7596 (N_7596,N_7022,N_7054);
xnor U7597 (N_7597,N_6998,N_6361);
and U7598 (N_7598,N_6372,N_7354);
xor U7599 (N_7599,N_7309,N_7307);
or U7600 (N_7600,N_6630,N_6703);
or U7601 (N_7601,N_7068,N_6680);
nand U7602 (N_7602,N_7471,N_7431);
nand U7603 (N_7603,N_6689,N_6334);
and U7604 (N_7604,N_7461,N_7258);
nand U7605 (N_7605,N_6876,N_7221);
nand U7606 (N_7606,N_6691,N_6462);
xor U7607 (N_7607,N_7423,N_7377);
or U7608 (N_7608,N_7251,N_7473);
and U7609 (N_7609,N_6619,N_6734);
xor U7610 (N_7610,N_6375,N_6685);
nand U7611 (N_7611,N_6762,N_6563);
xnor U7612 (N_7612,N_6416,N_6753);
or U7613 (N_7613,N_7040,N_6570);
or U7614 (N_7614,N_6682,N_7015);
nand U7615 (N_7615,N_7482,N_6423);
nand U7616 (N_7616,N_6845,N_6320);
nand U7617 (N_7617,N_6916,N_7497);
nor U7618 (N_7618,N_6862,N_6698);
xor U7619 (N_7619,N_6742,N_7353);
nand U7620 (N_7620,N_6347,N_7300);
xnor U7621 (N_7621,N_7247,N_6359);
xnor U7622 (N_7622,N_6857,N_6578);
nand U7623 (N_7623,N_7352,N_7212);
xnor U7624 (N_7624,N_7265,N_6611);
and U7625 (N_7625,N_7373,N_7444);
xnor U7626 (N_7626,N_6280,N_6409);
and U7627 (N_7627,N_6524,N_7375);
and U7628 (N_7628,N_7216,N_6362);
or U7629 (N_7629,N_7239,N_6582);
nor U7630 (N_7630,N_6366,N_7052);
nand U7631 (N_7631,N_6433,N_6910);
and U7632 (N_7632,N_6996,N_7316);
xor U7633 (N_7633,N_6759,N_6684);
xnor U7634 (N_7634,N_6351,N_6271);
and U7635 (N_7635,N_7308,N_6329);
nor U7636 (N_7636,N_7442,N_6621);
or U7637 (N_7637,N_7180,N_6538);
nor U7638 (N_7638,N_6839,N_6413);
and U7639 (N_7639,N_7103,N_7092);
or U7640 (N_7640,N_6837,N_6311);
xor U7641 (N_7641,N_6888,N_7421);
nand U7642 (N_7642,N_7034,N_6589);
or U7643 (N_7643,N_7345,N_6730);
nand U7644 (N_7644,N_6309,N_7256);
and U7645 (N_7645,N_7039,N_7255);
nand U7646 (N_7646,N_6674,N_7130);
xor U7647 (N_7647,N_7480,N_6391);
nand U7648 (N_7648,N_7172,N_6536);
or U7649 (N_7649,N_6406,N_6267);
nor U7650 (N_7650,N_7429,N_7317);
or U7651 (N_7651,N_7392,N_6404);
xnor U7652 (N_7652,N_7234,N_6919);
and U7653 (N_7653,N_6658,N_7273);
and U7654 (N_7654,N_7427,N_7244);
nor U7655 (N_7655,N_6405,N_6705);
xor U7656 (N_7656,N_6526,N_6449);
nand U7657 (N_7657,N_6385,N_6983);
and U7658 (N_7658,N_7351,N_6826);
nor U7659 (N_7659,N_6896,N_6953);
and U7660 (N_7660,N_7430,N_6467);
nor U7661 (N_7661,N_6584,N_6258);
nand U7662 (N_7662,N_6552,N_7435);
and U7663 (N_7663,N_6849,N_6319);
and U7664 (N_7664,N_7327,N_6468);
and U7665 (N_7665,N_6938,N_7334);
nor U7666 (N_7666,N_6771,N_7152);
nand U7667 (N_7667,N_6942,N_7452);
nand U7668 (N_7668,N_6364,N_6325);
xor U7669 (N_7669,N_7115,N_7023);
or U7670 (N_7670,N_6295,N_6884);
and U7671 (N_7671,N_7230,N_7396);
nor U7672 (N_7672,N_7065,N_7099);
xor U7673 (N_7673,N_6642,N_7175);
and U7674 (N_7674,N_6287,N_6317);
or U7675 (N_7675,N_6615,N_7467);
nor U7676 (N_7676,N_7021,N_6731);
and U7677 (N_7677,N_6804,N_6644);
or U7678 (N_7678,N_6828,N_6697);
and U7679 (N_7679,N_6496,N_7403);
xor U7680 (N_7680,N_6326,N_6715);
nor U7681 (N_7681,N_6392,N_6579);
or U7682 (N_7682,N_6307,N_6696);
nor U7683 (N_7683,N_7458,N_6612);
and U7684 (N_7684,N_6590,N_6920);
xor U7685 (N_7685,N_6714,N_7451);
and U7686 (N_7686,N_6330,N_7464);
xnor U7687 (N_7687,N_7113,N_6781);
nor U7688 (N_7688,N_6435,N_7104);
or U7689 (N_7689,N_6288,N_6451);
xor U7690 (N_7690,N_7166,N_7093);
nand U7691 (N_7691,N_6834,N_6871);
or U7692 (N_7692,N_7363,N_7083);
nand U7693 (N_7693,N_7098,N_6875);
nor U7694 (N_7694,N_6631,N_7409);
and U7695 (N_7695,N_7094,N_6848);
nor U7696 (N_7696,N_7275,N_6464);
xor U7697 (N_7697,N_6988,N_7076);
and U7698 (N_7698,N_6525,N_6323);
xor U7699 (N_7699,N_6507,N_6846);
nand U7700 (N_7700,N_7072,N_6403);
nor U7701 (N_7701,N_7232,N_6286);
xnor U7702 (N_7702,N_6706,N_7245);
xnor U7703 (N_7703,N_7126,N_6779);
and U7704 (N_7704,N_6729,N_6534);
nand U7705 (N_7705,N_7035,N_6663);
or U7706 (N_7706,N_6897,N_6376);
nand U7707 (N_7707,N_7356,N_6291);
nand U7708 (N_7708,N_7274,N_7231);
nor U7709 (N_7709,N_6441,N_6683);
xnor U7710 (N_7710,N_7106,N_6746);
nor U7711 (N_7711,N_7075,N_6627);
nor U7712 (N_7712,N_6502,N_6652);
nor U7713 (N_7713,N_6632,N_6735);
nor U7714 (N_7714,N_7378,N_6993);
nor U7715 (N_7715,N_7422,N_7405);
nor U7716 (N_7716,N_6548,N_7238);
nand U7717 (N_7717,N_6623,N_6763);
nor U7718 (N_7718,N_7449,N_6936);
or U7719 (N_7719,N_6820,N_7004);
nor U7720 (N_7720,N_6660,N_7417);
xnor U7721 (N_7721,N_6963,N_7457);
xnor U7722 (N_7722,N_6352,N_6314);
nand U7723 (N_7723,N_7100,N_6646);
nor U7724 (N_7724,N_6791,N_7385);
xnor U7725 (N_7725,N_7087,N_7026);
nand U7726 (N_7726,N_6363,N_7137);
and U7727 (N_7727,N_6447,N_7269);
xor U7728 (N_7728,N_7117,N_6516);
or U7729 (N_7729,N_6310,N_6407);
or U7730 (N_7730,N_7402,N_6694);
or U7731 (N_7731,N_7227,N_6348);
nand U7732 (N_7732,N_6847,N_7217);
and U7733 (N_7733,N_7299,N_6637);
and U7734 (N_7734,N_6973,N_6335);
nor U7735 (N_7735,N_7336,N_6456);
xnor U7736 (N_7736,N_6400,N_6795);
or U7737 (N_7737,N_7411,N_6737);
and U7738 (N_7738,N_7210,N_7082);
nor U7739 (N_7739,N_6890,N_7294);
nand U7740 (N_7740,N_6789,N_7318);
or U7741 (N_7741,N_7031,N_6629);
nor U7742 (N_7742,N_6990,N_7339);
xor U7743 (N_7743,N_7282,N_6471);
xnor U7744 (N_7744,N_7486,N_6662);
nor U7745 (N_7745,N_6282,N_6648);
or U7746 (N_7746,N_6470,N_7249);
and U7747 (N_7747,N_7489,N_7053);
nand U7748 (N_7748,N_6788,N_6785);
xnor U7749 (N_7749,N_7097,N_7248);
nand U7750 (N_7750,N_6542,N_7067);
nand U7751 (N_7751,N_6381,N_7271);
xnor U7752 (N_7752,N_6254,N_7179);
or U7753 (N_7753,N_6961,N_7218);
nand U7754 (N_7754,N_7153,N_7225);
nand U7755 (N_7755,N_6266,N_6595);
xnor U7756 (N_7756,N_6341,N_7295);
xnor U7757 (N_7757,N_7391,N_6798);
or U7758 (N_7758,N_6613,N_7481);
or U7759 (N_7759,N_6830,N_6365);
nor U7760 (N_7760,N_7463,N_6384);
xnor U7761 (N_7761,N_6543,N_7207);
nor U7762 (N_7762,N_6744,N_6643);
nor U7763 (N_7763,N_6500,N_7415);
or U7764 (N_7764,N_6688,N_6673);
or U7765 (N_7765,N_6279,N_6605);
or U7766 (N_7766,N_7183,N_6398);
or U7767 (N_7767,N_7278,N_7160);
nand U7768 (N_7768,N_6664,N_6893);
and U7769 (N_7769,N_7450,N_6636);
or U7770 (N_7770,N_6949,N_7492);
xnor U7771 (N_7771,N_6917,N_6299);
and U7772 (N_7772,N_6349,N_6976);
nand U7773 (N_7773,N_7133,N_7321);
xnor U7774 (N_7774,N_6902,N_7425);
or U7775 (N_7775,N_7199,N_6617);
nor U7776 (N_7776,N_7162,N_7206);
and U7777 (N_7777,N_6342,N_6360);
or U7778 (N_7778,N_6678,N_6289);
nand U7779 (N_7779,N_7338,N_7312);
or U7780 (N_7780,N_7038,N_7286);
nand U7781 (N_7781,N_6867,N_6262);
xor U7782 (N_7782,N_7017,N_7477);
nor U7783 (N_7783,N_6906,N_7488);
or U7784 (N_7784,N_6655,N_6518);
or U7785 (N_7785,N_7313,N_6556);
xor U7786 (N_7786,N_7016,N_7324);
and U7787 (N_7787,N_6784,N_7044);
xnor U7788 (N_7788,N_6721,N_6889);
nor U7789 (N_7789,N_6908,N_7303);
and U7790 (N_7790,N_6898,N_6429);
nor U7791 (N_7791,N_7086,N_6498);
nor U7792 (N_7792,N_7362,N_6895);
nor U7793 (N_7793,N_7292,N_6576);
nand U7794 (N_7794,N_6679,N_6959);
nand U7795 (N_7795,N_7494,N_7136);
nand U7796 (N_7796,N_6412,N_6305);
or U7797 (N_7797,N_7195,N_7326);
and U7798 (N_7798,N_6927,N_7155);
xor U7799 (N_7799,N_6728,N_6402);
xnor U7800 (N_7800,N_6894,N_6255);
nand U7801 (N_7801,N_6252,N_6760);
or U7802 (N_7802,N_6492,N_6493);
nand U7803 (N_7803,N_6350,N_7253);
xnor U7804 (N_7804,N_7445,N_6718);
nor U7805 (N_7805,N_7164,N_6600);
nor U7806 (N_7806,N_7368,N_7069);
xor U7807 (N_7807,N_7349,N_6782);
nor U7808 (N_7808,N_7285,N_7382);
nor U7809 (N_7809,N_7029,N_7495);
and U7810 (N_7810,N_6354,N_7209);
xor U7811 (N_7811,N_7005,N_6911);
nor U7812 (N_7812,N_6396,N_7090);
or U7813 (N_7813,N_6626,N_7364);
and U7814 (N_7814,N_6755,N_7298);
nand U7815 (N_7815,N_6585,N_7084);
or U7816 (N_7816,N_6659,N_6575);
nand U7817 (N_7817,N_7328,N_7456);
or U7818 (N_7818,N_7306,N_6390);
and U7819 (N_7819,N_6378,N_6440);
nand U7820 (N_7820,N_6654,N_7205);
nand U7821 (N_7821,N_6861,N_7242);
nor U7822 (N_7822,N_6514,N_6823);
xor U7823 (N_7823,N_6318,N_7150);
nand U7824 (N_7824,N_6302,N_6610);
xor U7825 (N_7825,N_7301,N_6599);
and U7826 (N_7826,N_6918,N_6399);
xor U7827 (N_7827,N_6251,N_7056);
xor U7828 (N_7828,N_6277,N_7414);
or U7829 (N_7829,N_6640,N_6473);
xnor U7830 (N_7830,N_6602,N_6950);
and U7831 (N_7831,N_7118,N_6340);
xnor U7832 (N_7832,N_6505,N_6256);
nor U7833 (N_7833,N_7165,N_6850);
xnor U7834 (N_7834,N_6923,N_6853);
nand U7835 (N_7835,N_6389,N_6977);
and U7836 (N_7836,N_7320,N_6494);
nand U7837 (N_7837,N_6499,N_6672);
xnor U7838 (N_7838,N_6686,N_7264);
and U7839 (N_7839,N_6695,N_7147);
nor U7840 (N_7840,N_6968,N_6947);
and U7841 (N_7841,N_7168,N_6315);
nand U7842 (N_7842,N_7131,N_6912);
nand U7843 (N_7843,N_6316,N_6308);
and U7844 (N_7844,N_6994,N_7057);
or U7845 (N_7845,N_6394,N_6356);
nor U7846 (N_7846,N_6922,N_6970);
xnor U7847 (N_7847,N_7438,N_7116);
xnor U7848 (N_7848,N_6490,N_7407);
nand U7849 (N_7849,N_6343,N_6374);
xnor U7850 (N_7850,N_7341,N_7260);
nand U7851 (N_7851,N_6461,N_6810);
or U7852 (N_7852,N_6987,N_6797);
xnor U7853 (N_7853,N_7447,N_6812);
or U7854 (N_7854,N_6768,N_7197);
or U7855 (N_7855,N_7174,N_6580);
nor U7856 (N_7856,N_7228,N_6635);
nor U7857 (N_7857,N_7111,N_6738);
or U7858 (N_7858,N_7156,N_7204);
xor U7859 (N_7859,N_6945,N_7184);
nor U7860 (N_7860,N_7012,N_6622);
and U7861 (N_7861,N_7214,N_7163);
and U7862 (N_7862,N_6418,N_7114);
or U7863 (N_7863,N_6438,N_6707);
nor U7864 (N_7864,N_6814,N_6285);
or U7865 (N_7865,N_7243,N_7019);
xnor U7866 (N_7866,N_6486,N_6339);
xor U7867 (N_7867,N_6786,N_7325);
and U7868 (N_7868,N_6442,N_6489);
xnor U7869 (N_7869,N_6531,N_6618);
and U7870 (N_7870,N_6792,N_7413);
nand U7871 (N_7871,N_7073,N_6860);
xor U7872 (N_7872,N_6353,N_7078);
or U7873 (N_7873,N_7394,N_6724);
and U7874 (N_7874,N_6869,N_6693);
or U7875 (N_7875,N_7418,N_7048);
nand U7876 (N_7876,N_6483,N_7045);
nor U7877 (N_7877,N_6829,N_6972);
or U7878 (N_7878,N_6880,N_7267);
nand U7879 (N_7879,N_7376,N_7224);
and U7880 (N_7880,N_6799,N_6268);
nor U7881 (N_7881,N_7235,N_6432);
nor U7882 (N_7882,N_6892,N_6304);
nor U7883 (N_7883,N_7041,N_7358);
and U7884 (N_7884,N_7074,N_6606);
nand U7885 (N_7885,N_7340,N_6275);
xor U7886 (N_7886,N_6609,N_6726);
nor U7887 (N_7887,N_7107,N_7109);
xor U7888 (N_7888,N_6460,N_6515);
xnor U7889 (N_7889,N_6292,N_6357);
nor U7890 (N_7890,N_7089,N_6369);
or U7891 (N_7891,N_6934,N_6944);
nand U7892 (N_7892,N_6832,N_7490);
nor U7893 (N_7893,N_7333,N_7101);
nand U7894 (N_7894,N_7433,N_6482);
or U7895 (N_7895,N_7010,N_7476);
or U7896 (N_7896,N_7060,N_6324);
nor U7897 (N_7897,N_6604,N_6511);
and U7898 (N_7898,N_7055,N_7003);
or U7899 (N_7899,N_6338,N_6508);
xor U7900 (N_7900,N_6748,N_7291);
or U7901 (N_7901,N_7009,N_6344);
nand U7902 (N_7902,N_7437,N_7121);
nand U7903 (N_7903,N_6769,N_6273);
and U7904 (N_7904,N_6725,N_6772);
xor U7905 (N_7905,N_6806,N_7280);
nand U7906 (N_7906,N_6588,N_6931);
xor U7907 (N_7907,N_6836,N_6653);
and U7908 (N_7908,N_6960,N_6747);
xor U7909 (N_7909,N_7266,N_6802);
or U7910 (N_7910,N_7139,N_6465);
nor U7911 (N_7911,N_6562,N_7419);
and U7912 (N_7912,N_6528,N_7263);
nor U7913 (N_7913,N_7261,N_6577);
nand U7914 (N_7914,N_7475,N_7032);
and U7915 (N_7915,N_6858,N_6634);
nor U7916 (N_7916,N_6380,N_6382);
xor U7917 (N_7917,N_7140,N_6535);
nand U7918 (N_7918,N_7011,N_6670);
and U7919 (N_7919,N_7281,N_6935);
nor U7920 (N_7920,N_7390,N_6926);
nand U7921 (N_7921,N_6774,N_6322);
nand U7922 (N_7922,N_6547,N_6752);
or U7923 (N_7923,N_7033,N_6967);
xnor U7924 (N_7924,N_6745,N_7215);
or U7925 (N_7925,N_6709,N_6943);
or U7926 (N_7926,N_7144,N_7079);
and U7927 (N_7927,N_6741,N_6520);
xor U7928 (N_7928,N_7323,N_6607);
and U7929 (N_7929,N_7459,N_6414);
and U7930 (N_7930,N_7167,N_6699);
nor U7931 (N_7931,N_6940,N_7096);
and U7932 (N_7932,N_6597,N_6620);
xnor U7933 (N_7933,N_6616,N_7443);
or U7934 (N_7934,N_6780,N_6909);
and U7935 (N_7935,N_6419,N_6567);
nor U7936 (N_7936,N_7454,N_6290);
or U7937 (N_7937,N_7188,N_6431);
nor U7938 (N_7938,N_6736,N_7315);
xor U7939 (N_7939,N_6816,N_7426);
nor U7940 (N_7940,N_6819,N_7289);
and U7941 (N_7941,N_6656,N_7222);
nand U7942 (N_7942,N_6601,N_6807);
xnor U7943 (N_7943,N_6756,N_7387);
xor U7944 (N_7944,N_6651,N_7124);
nand U7945 (N_7945,N_6716,N_6463);
nand U7946 (N_7946,N_6803,N_7420);
or U7947 (N_7947,N_7474,N_6966);
nor U7948 (N_7948,N_7479,N_6313);
xnor U7949 (N_7949,N_7290,N_6891);
and U7950 (N_7950,N_6504,N_7213);
and U7951 (N_7951,N_6455,N_6497);
xnor U7952 (N_7952,N_7372,N_6981);
nand U7953 (N_7953,N_7478,N_6818);
nor U7954 (N_7954,N_6373,N_7440);
nor U7955 (N_7955,N_6859,N_6787);
xnor U7956 (N_7956,N_7493,N_6270);
nand U7957 (N_7957,N_6586,N_7384);
or U7958 (N_7958,N_6914,N_7466);
xnor U7959 (N_7959,N_7178,N_6824);
xnor U7960 (N_7960,N_6560,N_6661);
nand U7961 (N_7961,N_6710,N_6476);
or U7962 (N_7962,N_7388,N_7393);
or U7963 (N_7963,N_6624,N_6681);
nor U7964 (N_7964,N_6263,N_7128);
nor U7965 (N_7965,N_6776,N_6928);
and U7966 (N_7966,N_6899,N_7194);
xor U7967 (N_7967,N_6903,N_6815);
or U7968 (N_7968,N_6427,N_6561);
and U7969 (N_7969,N_6568,N_6767);
and U7970 (N_7970,N_7272,N_6687);
xor U7971 (N_7971,N_7070,N_6480);
xnor U7972 (N_7972,N_6554,N_6666);
or U7973 (N_7973,N_6883,N_6457);
xor U7974 (N_7974,N_6522,N_6667);
and U7975 (N_7975,N_7277,N_6519);
or U7976 (N_7976,N_6740,N_7428);
xor U7977 (N_7977,N_6925,N_6625);
or U7978 (N_7978,N_7359,N_7059);
or U7979 (N_7979,N_6999,N_7469);
and U7980 (N_7980,N_6336,N_7202);
nor U7981 (N_7981,N_7343,N_7389);
and U7982 (N_7982,N_6411,N_6297);
nand U7983 (N_7983,N_6863,N_7071);
or U7984 (N_7984,N_6904,N_6395);
or U7985 (N_7985,N_7201,N_6766);
nand U7986 (N_7986,N_7383,N_6337);
or U7987 (N_7987,N_6793,N_7424);
and U7988 (N_7988,N_7025,N_7135);
and U7989 (N_7989,N_6956,N_7000);
xor U7990 (N_7990,N_7297,N_6647);
xor U7991 (N_7991,N_6555,N_7030);
or U7992 (N_7992,N_6401,N_7371);
nand U7993 (N_7993,N_7088,N_6957);
and U7994 (N_7994,N_7223,N_6603);
nand U7995 (N_7995,N_6870,N_6727);
and U7996 (N_7996,N_7037,N_6712);
and U7997 (N_7997,N_6501,N_6596);
nand U7998 (N_7998,N_7311,N_6951);
nand U7999 (N_7999,N_6379,N_6825);
and U8000 (N_8000,N_6571,N_6929);
and U8001 (N_8001,N_6852,N_6434);
xor U8002 (N_8002,N_7018,N_6424);
xor U8003 (N_8003,N_7346,N_6764);
or U8004 (N_8004,N_6811,N_7305);
xnor U8005 (N_8005,N_7085,N_7399);
nor U8006 (N_8006,N_7108,N_6265);
xor U8007 (N_8007,N_6478,N_6854);
nor U8008 (N_8008,N_7360,N_6842);
nor U8009 (N_8009,N_6711,N_6481);
xor U8010 (N_8010,N_7499,N_6506);
and U8011 (N_8011,N_6574,N_7105);
xnor U8012 (N_8012,N_7455,N_6346);
nor U8013 (N_8013,N_7348,N_6749);
nor U8014 (N_8014,N_7176,N_6331);
nor U8015 (N_8015,N_6377,N_6885);
xnor U8016 (N_8016,N_7229,N_6939);
nor U8017 (N_8017,N_6757,N_6458);
xor U8018 (N_8018,N_6856,N_6657);
nor U8019 (N_8019,N_7288,N_7268);
nand U8020 (N_8020,N_6321,N_6614);
nor U8021 (N_8021,N_7013,N_7049);
nor U8022 (N_8022,N_7330,N_6358);
nor U8023 (N_8023,N_6474,N_7171);
and U8024 (N_8024,N_6717,N_6593);
or U8025 (N_8025,N_6333,N_7406);
and U8026 (N_8026,N_6733,N_7250);
xor U8027 (N_8027,N_6633,N_6878);
nor U8028 (N_8028,N_6676,N_7182);
nand U8029 (N_8029,N_6743,N_6281);
xor U8030 (N_8030,N_6260,N_7483);
nor U8031 (N_8031,N_7398,N_6946);
xor U8032 (N_8032,N_6533,N_6843);
or U8033 (N_8033,N_6844,N_6992);
and U8034 (N_8034,N_6278,N_6371);
or U8035 (N_8035,N_7129,N_6969);
nand U8036 (N_8036,N_7080,N_6813);
and U8037 (N_8037,N_6777,N_6485);
xor U8038 (N_8038,N_6303,N_6417);
or U8039 (N_8039,N_7484,N_6948);
nor U8040 (N_8040,N_6539,N_6671);
or U8041 (N_8041,N_7241,N_7149);
xnor U8042 (N_8042,N_6453,N_6978);
nand U8043 (N_8043,N_6692,N_7252);
nand U8044 (N_8044,N_7061,N_6439);
nand U8045 (N_8045,N_6521,N_6669);
or U8046 (N_8046,N_7369,N_7468);
nor U8047 (N_8047,N_7006,N_6930);
and U8048 (N_8048,N_7257,N_7014);
nor U8049 (N_8049,N_7138,N_7200);
nand U8050 (N_8050,N_6831,N_6559);
or U8051 (N_8051,N_7062,N_7169);
or U8052 (N_8052,N_7310,N_7047);
nand U8053 (N_8053,N_7122,N_6872);
and U8054 (N_8054,N_7119,N_6510);
and U8055 (N_8055,N_6989,N_7347);
and U8056 (N_8056,N_6283,N_7276);
nor U8057 (N_8057,N_6269,N_7410);
nor U8058 (N_8058,N_6701,N_6975);
or U8059 (N_8059,N_7219,N_6879);
nand U8060 (N_8060,N_6690,N_7408);
nor U8061 (N_8061,N_6327,N_6355);
or U8062 (N_8062,N_6541,N_6720);
nand U8063 (N_8063,N_6719,N_6982);
and U8064 (N_8064,N_7063,N_7283);
xor U8065 (N_8065,N_6257,N_6773);
or U8066 (N_8066,N_7329,N_6965);
or U8067 (N_8067,N_6553,N_7434);
and U8068 (N_8068,N_7220,N_6809);
and U8069 (N_8069,N_6821,N_7001);
nand U8070 (N_8070,N_6479,N_6822);
xnor U8071 (N_8071,N_7259,N_6540);
xor U8072 (N_8072,N_6512,N_6952);
and U8073 (N_8073,N_6751,N_6454);
nand U8074 (N_8074,N_6700,N_6758);
xor U8075 (N_8075,N_7344,N_6569);
xnor U8076 (N_8076,N_6732,N_6932);
xor U8077 (N_8077,N_7064,N_7024);
and U8078 (N_8078,N_6425,N_7487);
nand U8079 (N_8079,N_6551,N_7342);
nand U8080 (N_8080,N_7270,N_7296);
and U8081 (N_8081,N_7432,N_7193);
and U8082 (N_8082,N_6259,N_6933);
or U8083 (N_8083,N_6750,N_7246);
xor U8084 (N_8084,N_7042,N_6886);
nor U8085 (N_8085,N_7237,N_7007);
xnor U8086 (N_8086,N_6397,N_7380);
xnor U8087 (N_8087,N_7081,N_7460);
nor U8088 (N_8088,N_6765,N_6817);
xor U8089 (N_8089,N_7439,N_6841);
nand U8090 (N_8090,N_7157,N_6421);
xor U8091 (N_8091,N_7374,N_6422);
nor U8092 (N_8092,N_7462,N_6997);
or U8093 (N_8093,N_6393,N_7350);
nor U8094 (N_8094,N_6855,N_7146);
nand U8095 (N_8095,N_7203,N_7485);
xor U8096 (N_8096,N_6796,N_6370);
and U8097 (N_8097,N_7412,N_7279);
nand U8098 (N_8098,N_6937,N_6472);
xor U8099 (N_8099,N_6974,N_7170);
nor U8100 (N_8100,N_6587,N_6778);
or U8101 (N_8101,N_6775,N_6566);
or U8102 (N_8102,N_6253,N_6517);
or U8103 (N_8103,N_6301,N_6877);
xor U8104 (N_8104,N_6428,N_7404);
nor U8105 (N_8105,N_6264,N_6564);
xnor U8106 (N_8106,N_7077,N_7142);
nand U8107 (N_8107,N_6445,N_7002);
or U8108 (N_8108,N_6761,N_6450);
and U8109 (N_8109,N_6984,N_7400);
xor U8110 (N_8110,N_6466,N_7465);
and U8111 (N_8111,N_7125,N_6272);
nor U8112 (N_8112,N_6985,N_6704);
xor U8113 (N_8113,N_7066,N_7314);
nand U8114 (N_8114,N_6638,N_6529);
and U8115 (N_8115,N_6312,N_7127);
or U8116 (N_8116,N_7120,N_6915);
and U8117 (N_8117,N_7357,N_6905);
xor U8118 (N_8118,N_6739,N_7110);
xor U8119 (N_8119,N_6367,N_6545);
xnor U8120 (N_8120,N_6294,N_7470);
and U8121 (N_8121,N_7058,N_6537);
nor U8122 (N_8122,N_7366,N_6702);
and U8123 (N_8123,N_7198,N_6284);
xor U8124 (N_8124,N_6865,N_6979);
nor U8125 (N_8125,N_6959,N_7243);
nand U8126 (N_8126,N_7288,N_7478);
xor U8127 (N_8127,N_7398,N_6589);
and U8128 (N_8128,N_7446,N_6522);
or U8129 (N_8129,N_7274,N_6833);
xnor U8130 (N_8130,N_7047,N_7163);
xnor U8131 (N_8131,N_6911,N_6726);
nand U8132 (N_8132,N_7417,N_7418);
and U8133 (N_8133,N_6960,N_6338);
nand U8134 (N_8134,N_7228,N_6730);
nor U8135 (N_8135,N_7394,N_7463);
xnor U8136 (N_8136,N_6934,N_6342);
and U8137 (N_8137,N_6882,N_6386);
or U8138 (N_8138,N_6855,N_7060);
xor U8139 (N_8139,N_7157,N_7025);
xnor U8140 (N_8140,N_7329,N_7497);
nand U8141 (N_8141,N_6521,N_6311);
nand U8142 (N_8142,N_6499,N_7219);
xor U8143 (N_8143,N_6974,N_6740);
and U8144 (N_8144,N_6806,N_7257);
and U8145 (N_8145,N_6707,N_7338);
nor U8146 (N_8146,N_7306,N_6660);
and U8147 (N_8147,N_6865,N_7463);
xor U8148 (N_8148,N_7139,N_6798);
nand U8149 (N_8149,N_7449,N_7070);
and U8150 (N_8150,N_6690,N_6745);
and U8151 (N_8151,N_7108,N_6414);
nor U8152 (N_8152,N_6478,N_7305);
or U8153 (N_8153,N_6277,N_6479);
xor U8154 (N_8154,N_7253,N_7268);
or U8155 (N_8155,N_6337,N_6445);
and U8156 (N_8156,N_6624,N_6657);
and U8157 (N_8157,N_7218,N_6584);
xor U8158 (N_8158,N_7483,N_7440);
nand U8159 (N_8159,N_6812,N_6251);
xor U8160 (N_8160,N_7295,N_6755);
nor U8161 (N_8161,N_7103,N_6741);
or U8162 (N_8162,N_6410,N_7079);
and U8163 (N_8163,N_7146,N_6926);
or U8164 (N_8164,N_6662,N_7272);
or U8165 (N_8165,N_7280,N_6562);
nor U8166 (N_8166,N_6575,N_7003);
nand U8167 (N_8167,N_7154,N_6491);
or U8168 (N_8168,N_7241,N_6640);
nor U8169 (N_8169,N_6709,N_6331);
nand U8170 (N_8170,N_7144,N_6672);
xor U8171 (N_8171,N_7245,N_7356);
or U8172 (N_8172,N_7098,N_7059);
or U8173 (N_8173,N_6937,N_7212);
or U8174 (N_8174,N_7210,N_7438);
xnor U8175 (N_8175,N_6810,N_6769);
xnor U8176 (N_8176,N_6502,N_7437);
and U8177 (N_8177,N_7013,N_7290);
or U8178 (N_8178,N_6633,N_6568);
nand U8179 (N_8179,N_6898,N_7198);
nand U8180 (N_8180,N_6649,N_7130);
and U8181 (N_8181,N_7180,N_6655);
nor U8182 (N_8182,N_6400,N_6778);
xor U8183 (N_8183,N_6313,N_6278);
or U8184 (N_8184,N_7261,N_6352);
nand U8185 (N_8185,N_7158,N_6767);
and U8186 (N_8186,N_7328,N_6283);
xor U8187 (N_8187,N_6936,N_6547);
xor U8188 (N_8188,N_6558,N_7249);
or U8189 (N_8189,N_6391,N_6781);
and U8190 (N_8190,N_6777,N_6342);
nand U8191 (N_8191,N_6948,N_7316);
or U8192 (N_8192,N_6277,N_6260);
nor U8193 (N_8193,N_6672,N_6641);
nand U8194 (N_8194,N_7439,N_7157);
nand U8195 (N_8195,N_7293,N_7306);
nand U8196 (N_8196,N_6276,N_7467);
or U8197 (N_8197,N_6624,N_7223);
xor U8198 (N_8198,N_6971,N_6743);
and U8199 (N_8199,N_7091,N_7205);
and U8200 (N_8200,N_6434,N_6262);
nor U8201 (N_8201,N_6897,N_7304);
nor U8202 (N_8202,N_7156,N_7291);
xnor U8203 (N_8203,N_7229,N_6295);
or U8204 (N_8204,N_7366,N_6500);
nor U8205 (N_8205,N_6967,N_6522);
and U8206 (N_8206,N_6871,N_7215);
and U8207 (N_8207,N_6306,N_7237);
xnor U8208 (N_8208,N_7056,N_6871);
and U8209 (N_8209,N_6561,N_6347);
and U8210 (N_8210,N_7175,N_6802);
nand U8211 (N_8211,N_7110,N_7265);
xor U8212 (N_8212,N_6636,N_7409);
or U8213 (N_8213,N_6781,N_6814);
nor U8214 (N_8214,N_7369,N_7394);
and U8215 (N_8215,N_7397,N_6857);
nand U8216 (N_8216,N_6948,N_7130);
and U8217 (N_8217,N_6480,N_7342);
nor U8218 (N_8218,N_7441,N_6884);
xor U8219 (N_8219,N_6416,N_7486);
nand U8220 (N_8220,N_7492,N_6373);
xor U8221 (N_8221,N_7320,N_7363);
nand U8222 (N_8222,N_7156,N_6269);
or U8223 (N_8223,N_6299,N_6907);
and U8224 (N_8224,N_7187,N_7394);
nor U8225 (N_8225,N_7321,N_7178);
nor U8226 (N_8226,N_7203,N_6958);
nor U8227 (N_8227,N_6634,N_6707);
or U8228 (N_8228,N_6841,N_6885);
nor U8229 (N_8229,N_6458,N_6715);
nor U8230 (N_8230,N_7444,N_6748);
nand U8231 (N_8231,N_6620,N_7218);
nor U8232 (N_8232,N_6450,N_6575);
nor U8233 (N_8233,N_7396,N_6371);
nand U8234 (N_8234,N_7148,N_6767);
xor U8235 (N_8235,N_6798,N_7320);
nand U8236 (N_8236,N_6648,N_6614);
or U8237 (N_8237,N_7337,N_6447);
xor U8238 (N_8238,N_6618,N_6268);
or U8239 (N_8239,N_7108,N_6405);
xnor U8240 (N_8240,N_6431,N_7377);
and U8241 (N_8241,N_6923,N_6386);
xor U8242 (N_8242,N_6553,N_7093);
xor U8243 (N_8243,N_6398,N_6898);
nand U8244 (N_8244,N_6336,N_7319);
xnor U8245 (N_8245,N_6299,N_6991);
xnor U8246 (N_8246,N_6627,N_6773);
xor U8247 (N_8247,N_6507,N_7044);
nor U8248 (N_8248,N_6278,N_6509);
nand U8249 (N_8249,N_6764,N_6376);
nor U8250 (N_8250,N_6767,N_6715);
or U8251 (N_8251,N_7373,N_6273);
or U8252 (N_8252,N_6405,N_7460);
and U8253 (N_8253,N_6433,N_7332);
nand U8254 (N_8254,N_7132,N_7255);
nand U8255 (N_8255,N_7473,N_7457);
nand U8256 (N_8256,N_7136,N_6346);
or U8257 (N_8257,N_7498,N_7404);
nor U8258 (N_8258,N_7241,N_6384);
or U8259 (N_8259,N_7045,N_6552);
nand U8260 (N_8260,N_7268,N_6655);
nor U8261 (N_8261,N_7281,N_6432);
nand U8262 (N_8262,N_7387,N_6472);
or U8263 (N_8263,N_6951,N_6602);
xor U8264 (N_8264,N_7212,N_7091);
nor U8265 (N_8265,N_7322,N_7167);
and U8266 (N_8266,N_7269,N_6260);
nor U8267 (N_8267,N_7054,N_6497);
nand U8268 (N_8268,N_7381,N_6755);
or U8269 (N_8269,N_7137,N_7408);
and U8270 (N_8270,N_7317,N_6595);
nor U8271 (N_8271,N_6749,N_7091);
nand U8272 (N_8272,N_7416,N_6905);
nand U8273 (N_8273,N_6413,N_6451);
nor U8274 (N_8274,N_7163,N_6685);
nand U8275 (N_8275,N_7151,N_7118);
nor U8276 (N_8276,N_6610,N_7296);
nor U8277 (N_8277,N_6395,N_6629);
or U8278 (N_8278,N_6920,N_6270);
nor U8279 (N_8279,N_7135,N_6642);
and U8280 (N_8280,N_6642,N_6536);
xnor U8281 (N_8281,N_7102,N_7386);
or U8282 (N_8282,N_7242,N_7397);
nand U8283 (N_8283,N_6463,N_6889);
or U8284 (N_8284,N_6299,N_6381);
or U8285 (N_8285,N_7427,N_7214);
nand U8286 (N_8286,N_6855,N_7357);
xor U8287 (N_8287,N_7428,N_7024);
nand U8288 (N_8288,N_6673,N_6747);
and U8289 (N_8289,N_7014,N_7339);
and U8290 (N_8290,N_7299,N_6823);
and U8291 (N_8291,N_6942,N_7006);
and U8292 (N_8292,N_6820,N_6740);
nand U8293 (N_8293,N_7382,N_6643);
nor U8294 (N_8294,N_6863,N_7010);
nor U8295 (N_8295,N_6747,N_6289);
nor U8296 (N_8296,N_6343,N_7140);
xor U8297 (N_8297,N_6576,N_7403);
xnor U8298 (N_8298,N_6452,N_7282);
and U8299 (N_8299,N_6551,N_7285);
or U8300 (N_8300,N_7469,N_7496);
xnor U8301 (N_8301,N_6567,N_6642);
xnor U8302 (N_8302,N_6968,N_7101);
or U8303 (N_8303,N_7069,N_6567);
xnor U8304 (N_8304,N_6667,N_6857);
and U8305 (N_8305,N_7017,N_6344);
or U8306 (N_8306,N_6762,N_7488);
and U8307 (N_8307,N_7226,N_7409);
nor U8308 (N_8308,N_6929,N_7058);
and U8309 (N_8309,N_6626,N_7042);
or U8310 (N_8310,N_6890,N_7213);
and U8311 (N_8311,N_7470,N_6582);
xnor U8312 (N_8312,N_6899,N_6793);
nor U8313 (N_8313,N_6814,N_6368);
or U8314 (N_8314,N_6423,N_7455);
or U8315 (N_8315,N_7190,N_7011);
xnor U8316 (N_8316,N_6290,N_6410);
nand U8317 (N_8317,N_6767,N_7285);
xnor U8318 (N_8318,N_6385,N_7242);
xnor U8319 (N_8319,N_6385,N_6723);
nor U8320 (N_8320,N_6927,N_6416);
nor U8321 (N_8321,N_6835,N_6690);
nor U8322 (N_8322,N_7187,N_6703);
nor U8323 (N_8323,N_6800,N_6525);
xnor U8324 (N_8324,N_6826,N_6678);
or U8325 (N_8325,N_6837,N_6714);
xnor U8326 (N_8326,N_7331,N_6357);
nor U8327 (N_8327,N_7070,N_7338);
xnor U8328 (N_8328,N_6651,N_7228);
nand U8329 (N_8329,N_6945,N_6727);
and U8330 (N_8330,N_7123,N_7163);
xnor U8331 (N_8331,N_6373,N_7334);
nand U8332 (N_8332,N_6425,N_6953);
nor U8333 (N_8333,N_7089,N_6876);
or U8334 (N_8334,N_7133,N_6779);
nand U8335 (N_8335,N_6609,N_6470);
nor U8336 (N_8336,N_6404,N_7350);
nand U8337 (N_8337,N_6681,N_6540);
and U8338 (N_8338,N_6955,N_7053);
and U8339 (N_8339,N_6778,N_7226);
or U8340 (N_8340,N_7259,N_7087);
xnor U8341 (N_8341,N_6645,N_6584);
nor U8342 (N_8342,N_6752,N_7109);
xnor U8343 (N_8343,N_6635,N_6850);
and U8344 (N_8344,N_6393,N_6826);
or U8345 (N_8345,N_6327,N_6947);
or U8346 (N_8346,N_6751,N_7383);
xor U8347 (N_8347,N_6490,N_7300);
nor U8348 (N_8348,N_6375,N_6396);
nand U8349 (N_8349,N_7375,N_7498);
or U8350 (N_8350,N_6522,N_7396);
xor U8351 (N_8351,N_6849,N_6962);
and U8352 (N_8352,N_6946,N_7197);
and U8353 (N_8353,N_7346,N_6266);
or U8354 (N_8354,N_7341,N_6597);
xnor U8355 (N_8355,N_7351,N_7353);
nor U8356 (N_8356,N_7402,N_6416);
nand U8357 (N_8357,N_6421,N_7132);
nand U8358 (N_8358,N_6449,N_6702);
and U8359 (N_8359,N_6743,N_6999);
and U8360 (N_8360,N_6728,N_7313);
nor U8361 (N_8361,N_7146,N_6485);
nor U8362 (N_8362,N_7162,N_6954);
or U8363 (N_8363,N_7324,N_6914);
nand U8364 (N_8364,N_7331,N_7339);
nand U8365 (N_8365,N_7171,N_6810);
nand U8366 (N_8366,N_6554,N_6590);
nor U8367 (N_8367,N_7426,N_7231);
xnor U8368 (N_8368,N_7172,N_7414);
and U8369 (N_8369,N_6738,N_6821);
and U8370 (N_8370,N_7281,N_6602);
nor U8371 (N_8371,N_7409,N_6854);
nand U8372 (N_8372,N_6266,N_6927);
nor U8373 (N_8373,N_6981,N_6928);
or U8374 (N_8374,N_7375,N_6555);
nand U8375 (N_8375,N_6791,N_7251);
or U8376 (N_8376,N_7476,N_7283);
nor U8377 (N_8377,N_7316,N_6750);
xnor U8378 (N_8378,N_6315,N_6278);
xnor U8379 (N_8379,N_6551,N_7298);
nor U8380 (N_8380,N_7269,N_7058);
and U8381 (N_8381,N_7111,N_7412);
nand U8382 (N_8382,N_7417,N_7372);
and U8383 (N_8383,N_7232,N_7006);
xor U8384 (N_8384,N_6979,N_6761);
xnor U8385 (N_8385,N_7043,N_6994);
nand U8386 (N_8386,N_6514,N_7039);
xor U8387 (N_8387,N_6993,N_7196);
and U8388 (N_8388,N_7079,N_7454);
nor U8389 (N_8389,N_7197,N_7234);
or U8390 (N_8390,N_6892,N_6950);
nand U8391 (N_8391,N_7323,N_7064);
xor U8392 (N_8392,N_7054,N_7091);
xnor U8393 (N_8393,N_7462,N_7352);
or U8394 (N_8394,N_6921,N_7314);
or U8395 (N_8395,N_6571,N_7182);
nand U8396 (N_8396,N_7405,N_6631);
xor U8397 (N_8397,N_7059,N_7396);
nor U8398 (N_8398,N_7231,N_6708);
nand U8399 (N_8399,N_6658,N_6603);
nand U8400 (N_8400,N_7470,N_6930);
or U8401 (N_8401,N_7076,N_7444);
and U8402 (N_8402,N_7462,N_6607);
nand U8403 (N_8403,N_7132,N_6823);
or U8404 (N_8404,N_7077,N_6803);
or U8405 (N_8405,N_7025,N_6850);
xnor U8406 (N_8406,N_6382,N_7081);
nand U8407 (N_8407,N_7169,N_7328);
xor U8408 (N_8408,N_7407,N_6604);
or U8409 (N_8409,N_7106,N_6427);
xnor U8410 (N_8410,N_7125,N_7339);
and U8411 (N_8411,N_7130,N_6562);
or U8412 (N_8412,N_6905,N_7239);
nor U8413 (N_8413,N_7114,N_6298);
nand U8414 (N_8414,N_6674,N_6428);
or U8415 (N_8415,N_6917,N_7069);
and U8416 (N_8416,N_7237,N_7413);
xnor U8417 (N_8417,N_6781,N_6255);
or U8418 (N_8418,N_6987,N_6748);
nor U8419 (N_8419,N_7223,N_6956);
nor U8420 (N_8420,N_6978,N_6484);
xnor U8421 (N_8421,N_6348,N_6401);
or U8422 (N_8422,N_6301,N_6367);
or U8423 (N_8423,N_7125,N_7157);
nor U8424 (N_8424,N_7437,N_6996);
nand U8425 (N_8425,N_6401,N_6912);
and U8426 (N_8426,N_6819,N_6845);
xnor U8427 (N_8427,N_6388,N_6327);
nor U8428 (N_8428,N_6917,N_6443);
or U8429 (N_8429,N_7247,N_7061);
and U8430 (N_8430,N_6564,N_7325);
and U8431 (N_8431,N_6604,N_6575);
and U8432 (N_8432,N_7309,N_6306);
nor U8433 (N_8433,N_6526,N_6565);
xor U8434 (N_8434,N_7286,N_6771);
xor U8435 (N_8435,N_6477,N_7429);
nor U8436 (N_8436,N_6559,N_6576);
and U8437 (N_8437,N_6658,N_7168);
xor U8438 (N_8438,N_6664,N_6632);
nor U8439 (N_8439,N_6742,N_6457);
and U8440 (N_8440,N_7273,N_7140);
xor U8441 (N_8441,N_7128,N_7330);
nand U8442 (N_8442,N_6772,N_6540);
nor U8443 (N_8443,N_7470,N_7126);
xnor U8444 (N_8444,N_6573,N_6622);
and U8445 (N_8445,N_7230,N_6691);
or U8446 (N_8446,N_6763,N_6536);
nand U8447 (N_8447,N_6669,N_6965);
nand U8448 (N_8448,N_6501,N_6633);
or U8449 (N_8449,N_6408,N_6781);
xor U8450 (N_8450,N_6730,N_6571);
or U8451 (N_8451,N_6848,N_7226);
or U8452 (N_8452,N_6425,N_7119);
xnor U8453 (N_8453,N_7239,N_6888);
and U8454 (N_8454,N_6547,N_6853);
and U8455 (N_8455,N_6312,N_6996);
or U8456 (N_8456,N_7333,N_6653);
nor U8457 (N_8457,N_6967,N_6720);
xnor U8458 (N_8458,N_7170,N_7059);
nand U8459 (N_8459,N_6557,N_7353);
and U8460 (N_8460,N_6791,N_6490);
nand U8461 (N_8461,N_7217,N_7461);
and U8462 (N_8462,N_6960,N_7082);
nand U8463 (N_8463,N_7337,N_7128);
or U8464 (N_8464,N_6774,N_7088);
nand U8465 (N_8465,N_7316,N_6535);
or U8466 (N_8466,N_7222,N_6592);
or U8467 (N_8467,N_6918,N_6543);
nand U8468 (N_8468,N_6827,N_7431);
nand U8469 (N_8469,N_6863,N_6380);
nor U8470 (N_8470,N_6986,N_7265);
and U8471 (N_8471,N_7013,N_6374);
nor U8472 (N_8472,N_6324,N_6638);
nand U8473 (N_8473,N_7267,N_6423);
nand U8474 (N_8474,N_6911,N_6257);
nor U8475 (N_8475,N_7223,N_6751);
xnor U8476 (N_8476,N_7124,N_7491);
xor U8477 (N_8477,N_6457,N_6301);
nor U8478 (N_8478,N_7254,N_7435);
or U8479 (N_8479,N_6535,N_7357);
xnor U8480 (N_8480,N_7024,N_6592);
nand U8481 (N_8481,N_7423,N_7453);
xnor U8482 (N_8482,N_6465,N_7153);
and U8483 (N_8483,N_7340,N_6483);
nor U8484 (N_8484,N_7247,N_6762);
and U8485 (N_8485,N_6548,N_6975);
nand U8486 (N_8486,N_6720,N_7111);
xor U8487 (N_8487,N_6906,N_7140);
and U8488 (N_8488,N_7314,N_6902);
nor U8489 (N_8489,N_6501,N_6901);
nand U8490 (N_8490,N_7001,N_6844);
nor U8491 (N_8491,N_6641,N_6684);
nand U8492 (N_8492,N_6839,N_6984);
nand U8493 (N_8493,N_7212,N_7415);
and U8494 (N_8494,N_6411,N_6898);
or U8495 (N_8495,N_6999,N_6614);
or U8496 (N_8496,N_6858,N_7262);
nor U8497 (N_8497,N_7059,N_6495);
nand U8498 (N_8498,N_7405,N_7072);
nand U8499 (N_8499,N_6355,N_6369);
nand U8500 (N_8500,N_7399,N_7275);
nor U8501 (N_8501,N_7160,N_6473);
nor U8502 (N_8502,N_7341,N_7258);
nand U8503 (N_8503,N_7477,N_6798);
xnor U8504 (N_8504,N_6289,N_7107);
nor U8505 (N_8505,N_7151,N_6468);
nand U8506 (N_8506,N_6385,N_6642);
and U8507 (N_8507,N_6361,N_6588);
and U8508 (N_8508,N_7275,N_7444);
nand U8509 (N_8509,N_6732,N_7386);
and U8510 (N_8510,N_7442,N_7058);
and U8511 (N_8511,N_6365,N_7468);
or U8512 (N_8512,N_6901,N_6350);
nor U8513 (N_8513,N_6614,N_7184);
nor U8514 (N_8514,N_6417,N_6457);
and U8515 (N_8515,N_6392,N_7031);
nor U8516 (N_8516,N_6787,N_6717);
and U8517 (N_8517,N_6674,N_7086);
nand U8518 (N_8518,N_7129,N_7162);
nand U8519 (N_8519,N_7283,N_7177);
or U8520 (N_8520,N_6638,N_6938);
or U8521 (N_8521,N_6799,N_7281);
and U8522 (N_8522,N_7069,N_7135);
or U8523 (N_8523,N_7215,N_6588);
nand U8524 (N_8524,N_6534,N_6351);
and U8525 (N_8525,N_6426,N_6494);
and U8526 (N_8526,N_6296,N_6823);
nand U8527 (N_8527,N_7014,N_7486);
nor U8528 (N_8528,N_6965,N_7086);
nand U8529 (N_8529,N_6557,N_6375);
nand U8530 (N_8530,N_7272,N_6255);
xnor U8531 (N_8531,N_7094,N_6353);
xor U8532 (N_8532,N_6514,N_6961);
xor U8533 (N_8533,N_6858,N_7132);
nor U8534 (N_8534,N_7322,N_7165);
xnor U8535 (N_8535,N_7480,N_6833);
nor U8536 (N_8536,N_6978,N_6503);
and U8537 (N_8537,N_6324,N_7476);
nor U8538 (N_8538,N_6687,N_6365);
nand U8539 (N_8539,N_7038,N_7202);
or U8540 (N_8540,N_6940,N_6710);
or U8541 (N_8541,N_6440,N_6781);
and U8542 (N_8542,N_7105,N_7142);
nor U8543 (N_8543,N_6597,N_7090);
nand U8544 (N_8544,N_6755,N_6735);
nand U8545 (N_8545,N_7391,N_6311);
nor U8546 (N_8546,N_6655,N_6463);
and U8547 (N_8547,N_6604,N_7353);
nand U8548 (N_8548,N_7259,N_7384);
or U8549 (N_8549,N_7245,N_7273);
or U8550 (N_8550,N_6759,N_7420);
nand U8551 (N_8551,N_6542,N_7398);
nand U8552 (N_8552,N_6735,N_6736);
nand U8553 (N_8553,N_6362,N_7225);
nand U8554 (N_8554,N_6484,N_6686);
nor U8555 (N_8555,N_7458,N_7385);
or U8556 (N_8556,N_6402,N_7296);
nand U8557 (N_8557,N_7455,N_7000);
xor U8558 (N_8558,N_6932,N_6738);
nor U8559 (N_8559,N_6929,N_6818);
xnor U8560 (N_8560,N_6649,N_7199);
or U8561 (N_8561,N_6492,N_6702);
xor U8562 (N_8562,N_7355,N_6772);
nor U8563 (N_8563,N_6475,N_6873);
nand U8564 (N_8564,N_7239,N_7277);
xnor U8565 (N_8565,N_7265,N_6750);
or U8566 (N_8566,N_6636,N_6534);
and U8567 (N_8567,N_6774,N_7089);
xor U8568 (N_8568,N_6547,N_7447);
and U8569 (N_8569,N_7048,N_6769);
or U8570 (N_8570,N_6818,N_6473);
xor U8571 (N_8571,N_6826,N_6623);
xnor U8572 (N_8572,N_7440,N_7491);
or U8573 (N_8573,N_7253,N_6907);
xnor U8574 (N_8574,N_7246,N_7404);
nor U8575 (N_8575,N_7444,N_7471);
xor U8576 (N_8576,N_7017,N_6591);
nand U8577 (N_8577,N_7083,N_6278);
and U8578 (N_8578,N_6400,N_7451);
nor U8579 (N_8579,N_6925,N_7116);
or U8580 (N_8580,N_6570,N_7265);
or U8581 (N_8581,N_6377,N_7014);
or U8582 (N_8582,N_6945,N_6961);
xor U8583 (N_8583,N_7432,N_6337);
xor U8584 (N_8584,N_6419,N_7029);
nor U8585 (N_8585,N_6413,N_6533);
or U8586 (N_8586,N_6270,N_6678);
or U8587 (N_8587,N_7014,N_6790);
nor U8588 (N_8588,N_6968,N_6596);
nor U8589 (N_8589,N_7437,N_7470);
and U8590 (N_8590,N_6787,N_6862);
or U8591 (N_8591,N_6550,N_7003);
nor U8592 (N_8592,N_6622,N_7293);
or U8593 (N_8593,N_7409,N_7100);
and U8594 (N_8594,N_6723,N_6967);
nor U8595 (N_8595,N_6626,N_7129);
and U8596 (N_8596,N_6741,N_7189);
or U8597 (N_8597,N_7013,N_7281);
and U8598 (N_8598,N_6589,N_6678);
nor U8599 (N_8599,N_6941,N_6830);
xor U8600 (N_8600,N_7044,N_7082);
and U8601 (N_8601,N_6613,N_7150);
and U8602 (N_8602,N_7180,N_6270);
nand U8603 (N_8603,N_6648,N_7323);
nor U8604 (N_8604,N_7102,N_7301);
nor U8605 (N_8605,N_7016,N_6820);
nor U8606 (N_8606,N_6438,N_6619);
nand U8607 (N_8607,N_6499,N_6865);
or U8608 (N_8608,N_6451,N_6997);
xor U8609 (N_8609,N_6516,N_6287);
or U8610 (N_8610,N_6277,N_6690);
nand U8611 (N_8611,N_6680,N_7202);
nor U8612 (N_8612,N_6749,N_6738);
nand U8613 (N_8613,N_7129,N_7216);
nor U8614 (N_8614,N_6489,N_6348);
nand U8615 (N_8615,N_6926,N_6602);
nor U8616 (N_8616,N_6812,N_6377);
nand U8617 (N_8617,N_6836,N_6297);
nor U8618 (N_8618,N_6616,N_6541);
xor U8619 (N_8619,N_7417,N_6713);
or U8620 (N_8620,N_6724,N_6912);
nand U8621 (N_8621,N_6697,N_6264);
nand U8622 (N_8622,N_7232,N_6641);
nand U8623 (N_8623,N_6905,N_7016);
or U8624 (N_8624,N_7296,N_7271);
nor U8625 (N_8625,N_6912,N_6422);
or U8626 (N_8626,N_7369,N_7423);
and U8627 (N_8627,N_6946,N_7302);
and U8628 (N_8628,N_6349,N_6597);
and U8629 (N_8629,N_7211,N_7178);
or U8630 (N_8630,N_6664,N_7337);
nor U8631 (N_8631,N_6909,N_6783);
or U8632 (N_8632,N_7415,N_6971);
or U8633 (N_8633,N_7039,N_7286);
nand U8634 (N_8634,N_6433,N_6904);
or U8635 (N_8635,N_7090,N_6310);
or U8636 (N_8636,N_6772,N_6724);
or U8637 (N_8637,N_6501,N_7204);
nand U8638 (N_8638,N_7018,N_6279);
and U8639 (N_8639,N_6684,N_7090);
or U8640 (N_8640,N_7258,N_7073);
or U8641 (N_8641,N_7165,N_7436);
xor U8642 (N_8642,N_7212,N_7100);
xnor U8643 (N_8643,N_6645,N_7031);
nand U8644 (N_8644,N_7118,N_6693);
and U8645 (N_8645,N_6997,N_6561);
and U8646 (N_8646,N_6821,N_6554);
or U8647 (N_8647,N_6682,N_6364);
nand U8648 (N_8648,N_6483,N_7433);
nand U8649 (N_8649,N_6636,N_6270);
xor U8650 (N_8650,N_6283,N_6531);
and U8651 (N_8651,N_7034,N_7490);
xor U8652 (N_8652,N_6998,N_6997);
xor U8653 (N_8653,N_6951,N_7400);
or U8654 (N_8654,N_6907,N_6338);
or U8655 (N_8655,N_6814,N_6801);
nand U8656 (N_8656,N_6814,N_6854);
nand U8657 (N_8657,N_6473,N_6541);
nand U8658 (N_8658,N_7371,N_6406);
xnor U8659 (N_8659,N_6430,N_7441);
or U8660 (N_8660,N_6854,N_6326);
or U8661 (N_8661,N_6484,N_7349);
and U8662 (N_8662,N_6537,N_7021);
and U8663 (N_8663,N_6650,N_6528);
or U8664 (N_8664,N_6772,N_6903);
or U8665 (N_8665,N_6681,N_6689);
or U8666 (N_8666,N_6899,N_7074);
nand U8667 (N_8667,N_7127,N_7403);
nor U8668 (N_8668,N_6298,N_7319);
or U8669 (N_8669,N_6868,N_6811);
or U8670 (N_8670,N_7399,N_7122);
nor U8671 (N_8671,N_7277,N_6736);
and U8672 (N_8672,N_6533,N_6308);
or U8673 (N_8673,N_7215,N_7449);
xor U8674 (N_8674,N_7199,N_7496);
nand U8675 (N_8675,N_7271,N_7157);
and U8676 (N_8676,N_7066,N_6271);
and U8677 (N_8677,N_7050,N_7213);
and U8678 (N_8678,N_7435,N_7146);
and U8679 (N_8679,N_7136,N_6265);
and U8680 (N_8680,N_7241,N_7256);
nand U8681 (N_8681,N_6599,N_6442);
nand U8682 (N_8682,N_7040,N_7337);
nand U8683 (N_8683,N_7231,N_6663);
or U8684 (N_8684,N_6596,N_7356);
nor U8685 (N_8685,N_7152,N_7493);
nor U8686 (N_8686,N_7073,N_6474);
nand U8687 (N_8687,N_7245,N_7220);
xnor U8688 (N_8688,N_6598,N_6450);
and U8689 (N_8689,N_6477,N_6863);
or U8690 (N_8690,N_6717,N_7418);
xor U8691 (N_8691,N_6675,N_6550);
or U8692 (N_8692,N_7206,N_6939);
or U8693 (N_8693,N_7264,N_6603);
nor U8694 (N_8694,N_7045,N_7276);
nor U8695 (N_8695,N_6710,N_7178);
xnor U8696 (N_8696,N_7059,N_6262);
and U8697 (N_8697,N_6871,N_7327);
nor U8698 (N_8698,N_6410,N_6505);
and U8699 (N_8699,N_6730,N_7313);
xnor U8700 (N_8700,N_6834,N_6591);
nor U8701 (N_8701,N_7028,N_7127);
and U8702 (N_8702,N_6434,N_6689);
and U8703 (N_8703,N_6851,N_6823);
or U8704 (N_8704,N_6351,N_7362);
and U8705 (N_8705,N_6906,N_7390);
nor U8706 (N_8706,N_6894,N_6456);
nand U8707 (N_8707,N_6959,N_6986);
nor U8708 (N_8708,N_6972,N_6663);
nand U8709 (N_8709,N_6611,N_7047);
nor U8710 (N_8710,N_6288,N_7335);
or U8711 (N_8711,N_7375,N_7176);
nand U8712 (N_8712,N_6915,N_6850);
and U8713 (N_8713,N_6278,N_6428);
or U8714 (N_8714,N_6417,N_7197);
nor U8715 (N_8715,N_6697,N_7206);
nor U8716 (N_8716,N_7364,N_7307);
or U8717 (N_8717,N_6736,N_7163);
nor U8718 (N_8718,N_6964,N_7231);
nand U8719 (N_8719,N_6439,N_6916);
nor U8720 (N_8720,N_6732,N_6347);
and U8721 (N_8721,N_6945,N_6704);
and U8722 (N_8722,N_7081,N_7188);
or U8723 (N_8723,N_6466,N_6887);
nor U8724 (N_8724,N_6819,N_6302);
and U8725 (N_8725,N_7263,N_6643);
xnor U8726 (N_8726,N_6680,N_7162);
xnor U8727 (N_8727,N_6295,N_6653);
xor U8728 (N_8728,N_6456,N_6466);
xnor U8729 (N_8729,N_7103,N_7428);
nor U8730 (N_8730,N_6432,N_6426);
or U8731 (N_8731,N_7316,N_6805);
and U8732 (N_8732,N_6761,N_6364);
nand U8733 (N_8733,N_6823,N_6860);
nand U8734 (N_8734,N_6252,N_7299);
xor U8735 (N_8735,N_6415,N_6406);
and U8736 (N_8736,N_7268,N_7421);
nor U8737 (N_8737,N_6255,N_7470);
or U8738 (N_8738,N_7042,N_7034);
xor U8739 (N_8739,N_7471,N_7267);
xor U8740 (N_8740,N_6603,N_6382);
and U8741 (N_8741,N_7343,N_7085);
nand U8742 (N_8742,N_6364,N_6634);
or U8743 (N_8743,N_6580,N_6785);
and U8744 (N_8744,N_7059,N_7128);
nor U8745 (N_8745,N_7416,N_6292);
xnor U8746 (N_8746,N_7283,N_7029);
or U8747 (N_8747,N_6793,N_7123);
xnor U8748 (N_8748,N_7173,N_6511);
or U8749 (N_8749,N_7004,N_6583);
nor U8750 (N_8750,N_8222,N_7767);
xor U8751 (N_8751,N_7636,N_7739);
xnor U8752 (N_8752,N_8198,N_7783);
and U8753 (N_8753,N_8283,N_8597);
and U8754 (N_8754,N_8266,N_7599);
nor U8755 (N_8755,N_8462,N_7754);
or U8756 (N_8756,N_7525,N_8588);
or U8757 (N_8757,N_8181,N_8669);
nor U8758 (N_8758,N_7878,N_7944);
or U8759 (N_8759,N_7942,N_8296);
nor U8760 (N_8760,N_7682,N_7723);
nand U8761 (N_8761,N_7912,N_7964);
nor U8762 (N_8762,N_7874,N_7749);
xnor U8763 (N_8763,N_7797,N_8385);
nor U8764 (N_8764,N_7616,N_8508);
nor U8765 (N_8765,N_8268,N_8446);
nand U8766 (N_8766,N_8285,N_8717);
xor U8767 (N_8767,N_7809,N_8312);
or U8768 (N_8768,N_7988,N_8425);
and U8769 (N_8769,N_8110,N_8005);
and U8770 (N_8770,N_8043,N_8246);
or U8771 (N_8771,N_8314,N_8592);
nor U8772 (N_8772,N_7715,N_8209);
or U8773 (N_8773,N_8474,N_8084);
nor U8774 (N_8774,N_8150,N_8599);
xor U8775 (N_8775,N_8131,N_7654);
or U8776 (N_8776,N_8277,N_7507);
nand U8777 (N_8777,N_8079,N_8227);
xnor U8778 (N_8778,N_8376,N_8306);
nand U8779 (N_8779,N_7983,N_7592);
nand U8780 (N_8780,N_7789,N_8677);
nor U8781 (N_8781,N_8457,N_8028);
nand U8782 (N_8782,N_8147,N_8031);
nor U8783 (N_8783,N_8279,N_7934);
nor U8784 (N_8784,N_8191,N_8322);
nand U8785 (N_8785,N_8078,N_8406);
xnor U8786 (N_8786,N_7518,N_8395);
nand U8787 (N_8787,N_8192,N_8284);
or U8788 (N_8788,N_8007,N_7824);
or U8789 (N_8789,N_7574,N_7893);
nand U8790 (N_8790,N_7710,N_8727);
or U8791 (N_8791,N_7625,N_8359);
and U8792 (N_8792,N_8747,N_8017);
xor U8793 (N_8793,N_7898,N_7872);
nor U8794 (N_8794,N_7840,N_8561);
xor U8795 (N_8795,N_8569,N_7848);
xor U8796 (N_8796,N_8418,N_8574);
nand U8797 (N_8797,N_8338,N_7502);
nand U8798 (N_8798,N_7930,N_8137);
and U8799 (N_8799,N_7564,N_8258);
nor U8800 (N_8800,N_7665,N_8094);
xnor U8801 (N_8801,N_7973,N_7796);
nand U8802 (N_8802,N_8009,N_7680);
or U8803 (N_8803,N_8026,N_8183);
xor U8804 (N_8804,N_8468,N_8030);
nor U8805 (N_8805,N_8719,N_8492);
nand U8806 (N_8806,N_7791,N_7613);
nor U8807 (N_8807,N_8441,N_7729);
xor U8808 (N_8808,N_8407,N_8722);
nor U8809 (N_8809,N_7867,N_8081);
xnor U8810 (N_8810,N_8257,N_8469);
nor U8811 (N_8811,N_8281,N_7588);
nor U8812 (N_8812,N_7871,N_8544);
and U8813 (N_8813,N_8251,N_7884);
or U8814 (N_8814,N_8336,N_8210);
nor U8815 (N_8815,N_7976,N_7632);
and U8816 (N_8816,N_7566,N_8313);
or U8817 (N_8817,N_7711,N_8220);
xnor U8818 (N_8818,N_8475,N_8151);
and U8819 (N_8819,N_8364,N_8311);
xnor U8820 (N_8820,N_8582,N_7825);
or U8821 (N_8821,N_8348,N_7559);
nand U8822 (N_8822,N_7759,N_8637);
and U8823 (N_8823,N_8627,N_8553);
xnor U8824 (N_8824,N_7788,N_8488);
nand U8825 (N_8825,N_7863,N_7556);
xnor U8826 (N_8826,N_7847,N_7583);
nor U8827 (N_8827,N_8093,N_7811);
nand U8828 (N_8828,N_7713,N_8608);
or U8829 (N_8829,N_8590,N_7902);
nand U8830 (N_8830,N_8269,N_8286);
and U8831 (N_8831,N_7883,N_8049);
nor U8832 (N_8832,N_8518,N_8309);
and U8833 (N_8833,N_8201,N_8153);
nor U8834 (N_8834,N_7866,N_8053);
nor U8835 (N_8835,N_7619,N_8485);
nand U8836 (N_8836,N_8214,N_8707);
or U8837 (N_8837,N_7508,N_7575);
or U8838 (N_8838,N_7536,N_7996);
or U8839 (N_8839,N_7717,N_8422);
nand U8840 (N_8840,N_8617,N_8231);
nand U8841 (N_8841,N_8662,N_7703);
and U8842 (N_8842,N_7532,N_7673);
nor U8843 (N_8843,N_8039,N_7937);
or U8844 (N_8844,N_8327,N_8540);
nand U8845 (N_8845,N_8687,N_7943);
and U8846 (N_8846,N_7600,N_7622);
and U8847 (N_8847,N_7845,N_8064);
and U8848 (N_8848,N_8352,N_8456);
xnor U8849 (N_8849,N_8573,N_8355);
or U8850 (N_8850,N_8448,N_8167);
or U8851 (N_8851,N_8433,N_7747);
xor U8852 (N_8852,N_8062,N_7728);
and U8853 (N_8853,N_8161,N_7774);
and U8854 (N_8854,N_7500,N_8700);
and U8855 (N_8855,N_8696,N_7869);
or U8856 (N_8856,N_8519,N_8480);
nor U8857 (N_8857,N_8587,N_8375);
or U8858 (N_8858,N_8447,N_8144);
xnor U8859 (N_8859,N_7799,N_8274);
xor U8860 (N_8860,N_7522,N_7980);
or U8861 (N_8861,N_7827,N_8333);
nand U8862 (N_8862,N_7505,N_8331);
nand U8863 (N_8863,N_8725,N_8729);
nor U8864 (N_8864,N_8550,N_8038);
and U8865 (N_8865,N_8105,N_8525);
nand U8866 (N_8866,N_7933,N_8136);
or U8867 (N_8867,N_8564,N_7699);
and U8868 (N_8868,N_7732,N_7766);
or U8869 (N_8869,N_8595,N_8109);
nor U8870 (N_8870,N_7537,N_7540);
nand U8871 (N_8871,N_8659,N_7635);
and U8872 (N_8872,N_8063,N_7877);
nor U8873 (N_8873,N_8413,N_8692);
or U8874 (N_8874,N_7590,N_7875);
nor U8875 (N_8875,N_7818,N_8168);
or U8876 (N_8876,N_8334,N_7610);
or U8877 (N_8877,N_8216,N_7596);
or U8878 (N_8878,N_8390,N_8373);
and U8879 (N_8879,N_7921,N_7515);
xor U8880 (N_8880,N_7666,N_7742);
nor U8881 (N_8881,N_8643,N_8559);
nor U8882 (N_8882,N_7951,N_7769);
nand U8883 (N_8883,N_8576,N_7855);
or U8884 (N_8884,N_8695,N_7862);
or U8885 (N_8885,N_7707,N_8675);
or U8886 (N_8886,N_8746,N_8232);
nand U8887 (N_8887,N_8353,N_7626);
nand U8888 (N_8888,N_7843,N_7519);
xnor U8889 (N_8889,N_7598,N_7568);
and U8890 (N_8890,N_7904,N_7770);
xor U8891 (N_8891,N_7919,N_8536);
and U8892 (N_8892,N_8575,N_8018);
nand U8893 (N_8893,N_8238,N_8683);
and U8894 (N_8894,N_8500,N_8023);
or U8895 (N_8895,N_8628,N_8521);
xnor U8896 (N_8896,N_8130,N_8688);
and U8897 (N_8897,N_7948,N_8638);
or U8898 (N_8898,N_8651,N_7648);
xor U8899 (N_8899,N_8034,N_7655);
nand U8900 (N_8900,N_8280,N_7593);
nor U8901 (N_8901,N_8567,N_8405);
or U8902 (N_8902,N_8021,N_8624);
and U8903 (N_8903,N_7523,N_8731);
nand U8904 (N_8904,N_8676,N_8234);
nand U8905 (N_8905,N_8491,N_7886);
and U8906 (N_8906,N_7755,N_7645);
nor U8907 (N_8907,N_7701,N_8530);
and U8908 (N_8908,N_7958,N_7546);
nand U8909 (N_8909,N_8744,N_7959);
and U8910 (N_8910,N_7837,N_7577);
nor U8911 (N_8911,N_7612,N_7631);
and U8912 (N_8912,N_8369,N_8495);
and U8913 (N_8913,N_8221,N_8732);
and U8914 (N_8914,N_7535,N_8558);
nand U8915 (N_8915,N_8660,N_7712);
nand U8916 (N_8916,N_7524,N_8070);
and U8917 (N_8917,N_7938,N_8261);
and U8918 (N_8918,N_7693,N_8438);
nor U8919 (N_8919,N_8092,N_8671);
xnor U8920 (N_8920,N_8114,N_8581);
nand U8921 (N_8921,N_8170,N_7910);
xnor U8922 (N_8922,N_7925,N_8149);
and U8923 (N_8923,N_8310,N_7646);
nand U8924 (N_8924,N_7814,N_8223);
nand U8925 (N_8925,N_7658,N_8159);
nor U8926 (N_8926,N_8562,N_8613);
nor U8927 (N_8927,N_8745,N_8726);
or U8928 (N_8928,N_7607,N_8256);
nor U8929 (N_8929,N_7901,N_7946);
and U8930 (N_8930,N_8354,N_7936);
nor U8931 (N_8931,N_7812,N_8622);
nand U8932 (N_8932,N_7589,N_7757);
or U8933 (N_8933,N_8211,N_8551);
nand U8934 (N_8934,N_8539,N_7700);
nand U8935 (N_8935,N_7801,N_7695);
and U8936 (N_8936,N_8351,N_7820);
nor U8937 (N_8937,N_7761,N_8012);
nand U8938 (N_8938,N_7614,N_7854);
nor U8939 (N_8939,N_8399,N_8734);
xnor U8940 (N_8940,N_7859,N_8097);
nand U8941 (N_8941,N_7989,N_8357);
xnor U8942 (N_8942,N_8206,N_8445);
xor U8943 (N_8943,N_8174,N_7579);
or U8944 (N_8944,N_8066,N_7621);
or U8945 (N_8945,N_8328,N_8027);
nand U8946 (N_8946,N_8554,N_7745);
or U8947 (N_8947,N_7852,N_8420);
nor U8948 (N_8948,N_7781,N_7580);
nor U8949 (N_8949,N_8000,N_8291);
xor U8950 (N_8950,N_8535,N_7851);
xor U8951 (N_8951,N_7746,N_8697);
xnor U8952 (N_8952,N_8089,N_7795);
nand U8953 (N_8953,N_8641,N_8188);
nand U8954 (N_8954,N_8400,N_7681);
and U8955 (N_8955,N_8004,N_8363);
or U8956 (N_8956,N_8102,N_7735);
or U8957 (N_8957,N_8247,N_8663);
nand U8958 (N_8958,N_8160,N_7653);
and U8959 (N_8959,N_8572,N_8640);
and U8960 (N_8960,N_7587,N_8449);
and U8961 (N_8961,N_7865,N_7839);
or U8962 (N_8962,N_7962,N_8496);
nor U8963 (N_8963,N_8712,N_8117);
and U8964 (N_8964,N_7963,N_8042);
and U8965 (N_8965,N_7652,N_7900);
and U8966 (N_8966,N_8403,N_7685);
xnor U8967 (N_8967,N_7690,N_8259);
nor U8968 (N_8968,N_8583,N_8740);
and U8969 (N_8969,N_8611,N_8245);
xnor U8970 (N_8970,N_8506,N_7618);
nor U8971 (N_8971,N_7911,N_7965);
and U8972 (N_8972,N_8557,N_8230);
or U8973 (N_8973,N_8386,N_7543);
or U8974 (N_8974,N_8080,N_8560);
nand U8975 (N_8975,N_8437,N_8233);
and U8976 (N_8976,N_7687,N_8527);
and U8977 (N_8977,N_7676,N_7941);
and U8978 (N_8978,N_7923,N_8370);
and U8979 (N_8979,N_8134,N_7932);
xnor U8980 (N_8980,N_8347,N_7786);
or U8981 (N_8981,N_8365,N_7914);
xnor U8982 (N_8982,N_8516,N_7803);
nand U8983 (N_8983,N_8204,N_7870);
xor U8984 (N_8984,N_8295,N_7952);
xnor U8985 (N_8985,N_8472,N_8463);
nor U8986 (N_8986,N_8392,N_7664);
or U8987 (N_8987,N_8749,N_8244);
xor U8988 (N_8988,N_8339,N_7947);
and U8989 (N_8989,N_8224,N_8393);
and U8990 (N_8990,N_8632,N_8631);
nand U8991 (N_8991,N_8476,N_7927);
nor U8992 (N_8992,N_8128,N_8185);
nand U8993 (N_8993,N_8195,N_8228);
nor U8994 (N_8994,N_7534,N_7576);
and U8995 (N_8995,N_7954,N_7503);
xor U8996 (N_8996,N_7853,N_7753);
nor U8997 (N_8997,N_8408,N_8529);
nor U8998 (N_8998,N_8095,N_8315);
nor U8999 (N_8999,N_8215,N_8654);
and U9000 (N_9000,N_7908,N_8022);
nor U9001 (N_9001,N_8416,N_8591);
nor U9002 (N_9002,N_7708,N_8265);
nor U9003 (N_9003,N_8158,N_8176);
nor U9004 (N_9004,N_7533,N_7868);
xor U9005 (N_9005,N_7586,N_7629);
and U9006 (N_9006,N_7716,N_7861);
nand U9007 (N_9007,N_7617,N_8694);
nor U9008 (N_9008,N_8415,N_7985);
nor U9009 (N_9009,N_7528,N_8250);
and U9010 (N_9010,N_7760,N_8524);
nand U9011 (N_9011,N_7724,N_8545);
nor U9012 (N_9012,N_8213,N_8497);
or U9013 (N_9013,N_8459,N_8388);
nand U9014 (N_9014,N_7808,N_8071);
xor U9015 (N_9015,N_7661,N_8479);
and U9016 (N_9016,N_7802,N_8240);
xnor U9017 (N_9017,N_8429,N_7987);
nand U9018 (N_9018,N_7800,N_8619);
xnor U9019 (N_9019,N_8596,N_7667);
or U9020 (N_9020,N_7916,N_8650);
and U9021 (N_9021,N_7897,N_7940);
nand U9022 (N_9022,N_7628,N_8145);
nand U9023 (N_9023,N_8050,N_8032);
xnor U9024 (N_9024,N_8382,N_8060);
or U9025 (N_9025,N_7705,N_8512);
and U9026 (N_9026,N_7553,N_8380);
nor U9027 (N_9027,N_8088,N_8625);
xnor U9028 (N_9028,N_8680,N_7644);
nor U9029 (N_9029,N_7999,N_8743);
or U9030 (N_9030,N_8054,N_8520);
or U9031 (N_9031,N_8024,N_7554);
nor U9032 (N_9032,N_8154,N_8267);
xnor U9033 (N_9033,N_8444,N_8200);
or U9034 (N_9034,N_8735,N_8389);
nor U9035 (N_9035,N_7756,N_7674);
or U9036 (N_9036,N_7634,N_8059);
xor U9037 (N_9037,N_8634,N_8297);
or U9038 (N_9038,N_8254,N_7849);
or U9039 (N_9039,N_8739,N_8642);
nand U9040 (N_9040,N_7513,N_7905);
and U9041 (N_9041,N_7822,N_7706);
xnor U9042 (N_9042,N_8040,N_8482);
nand U9043 (N_9043,N_8543,N_7961);
nand U9044 (N_9044,N_7858,N_7981);
xor U9045 (N_9045,N_7888,N_7955);
or U9046 (N_9046,N_8620,N_8452);
xor U9047 (N_9047,N_8427,N_7775);
xnor U9048 (N_9048,N_7581,N_8412);
nand U9049 (N_9049,N_8273,N_7890);
or U9050 (N_9050,N_8691,N_7597);
nand U9051 (N_9051,N_7828,N_8616);
and U9052 (N_9052,N_8604,N_7551);
nand U9053 (N_9053,N_7844,N_8718);
or U9054 (N_9054,N_7831,N_7967);
xor U9055 (N_9055,N_8451,N_8035);
xnor U9056 (N_9056,N_8271,N_8276);
nand U9057 (N_9057,N_8398,N_8686);
nor U9058 (N_9058,N_8523,N_8278);
nor U9059 (N_9059,N_8693,N_8229);
and U9060 (N_9060,N_8436,N_8293);
and U9061 (N_9061,N_8330,N_7887);
or U9062 (N_9062,N_8442,N_8318);
xor U9063 (N_9063,N_8504,N_8566);
or U9064 (N_9064,N_8001,N_7662);
and U9065 (N_9065,N_7529,N_7894);
or U9066 (N_9066,N_8402,N_7565);
nand U9067 (N_9067,N_7560,N_8341);
nor U9068 (N_9068,N_8493,N_8678);
or U9069 (N_9069,N_8419,N_8219);
nand U9070 (N_9070,N_8139,N_8517);
xnor U9071 (N_9071,N_8533,N_8260);
xnor U9072 (N_9072,N_8172,N_8454);
nor U9073 (N_9073,N_7856,N_8679);
and U9074 (N_9074,N_8720,N_8664);
or U9075 (N_9075,N_7702,N_8321);
xor U9076 (N_9076,N_8610,N_7917);
nand U9077 (N_9077,N_7918,N_8076);
and U9078 (N_9078,N_7798,N_7953);
and U9079 (N_9079,N_8723,N_8119);
or U9080 (N_9080,N_8371,N_7549);
and U9081 (N_9081,N_8367,N_8115);
nand U9082 (N_9082,N_8171,N_7578);
nand U9083 (N_9083,N_7939,N_8486);
nor U9084 (N_9084,N_8568,N_8455);
nand U9085 (N_9085,N_8409,N_8738);
or U9086 (N_9086,N_8248,N_8041);
xnor U9087 (N_9087,N_7928,N_7748);
or U9088 (N_9088,N_8253,N_7957);
nand U9089 (N_9089,N_8087,N_8118);
nand U9090 (N_9090,N_8629,N_7915);
or U9091 (N_9091,N_8262,N_8458);
or U9092 (N_9092,N_7733,N_7725);
and U9093 (N_9093,N_7823,N_7697);
and U9094 (N_9094,N_8316,N_8626);
nand U9095 (N_9095,N_8464,N_7741);
xnor U9096 (N_9096,N_8125,N_7516);
nor U9097 (N_9097,N_8074,N_7977);
and U9098 (N_9098,N_8381,N_7569);
xor U9099 (N_9099,N_7885,N_7738);
and U9100 (N_9100,N_8630,N_7704);
and U9101 (N_9101,N_8709,N_7696);
nand U9102 (N_9102,N_8414,N_7547);
or U9103 (N_9103,N_8397,N_7841);
or U9104 (N_9104,N_8166,N_7892);
nor U9105 (N_9105,N_8498,N_7765);
nor U9106 (N_9106,N_8202,N_8471);
nand U9107 (N_9107,N_8360,N_8708);
xor U9108 (N_9108,N_8470,N_8298);
nor U9109 (N_9109,N_8345,N_8661);
nor U9110 (N_9110,N_8699,N_7512);
xor U9111 (N_9111,N_7771,N_8716);
xnor U9112 (N_9112,N_8730,N_8647);
xnor U9113 (N_9113,N_7671,N_7567);
xnor U9114 (N_9114,N_8226,N_7677);
nand U9115 (N_9115,N_8346,N_8075);
nand U9116 (N_9116,N_8288,N_8391);
xor U9117 (N_9117,N_7604,N_8431);
or U9118 (N_9118,N_7743,N_7633);
nand U9119 (N_9119,N_7772,N_8721);
xnor U9120 (N_9120,N_8666,N_8607);
xnor U9121 (N_9121,N_8635,N_7530);
xnor U9122 (N_9122,N_7876,N_7995);
nor U9123 (N_9123,N_7584,N_7683);
xnor U9124 (N_9124,N_8072,N_8706);
nor U9125 (N_9125,N_7517,N_8531);
nand U9126 (N_9126,N_7881,N_7949);
xnor U9127 (N_9127,N_7538,N_7561);
nor U9128 (N_9128,N_7982,N_8547);
nor U9129 (N_9129,N_8335,N_8598);
and U9130 (N_9130,N_8439,N_8307);
nand U9131 (N_9131,N_8182,N_8065);
or U9132 (N_9132,N_7678,N_8173);
or U9133 (N_9133,N_7891,N_8636);
xor U9134 (N_9134,N_8156,N_8148);
or U9135 (N_9135,N_7555,N_7544);
nand U9136 (N_9136,N_8058,N_7929);
and U9137 (N_9137,N_8428,N_8673);
and U9138 (N_9138,N_7510,N_7882);
and U9139 (N_9139,N_8308,N_8112);
nand U9140 (N_9140,N_8421,N_8203);
nor U9141 (N_9141,N_8098,N_8129);
or U9142 (N_9142,N_8644,N_7926);
or U9143 (N_9143,N_8702,N_8401);
or U9144 (N_9144,N_7609,N_8655);
or U9145 (N_9145,N_7991,N_8703);
xnor U9146 (N_9146,N_7993,N_8342);
xor U9147 (N_9147,N_7968,N_7777);
nor U9148 (N_9148,N_8014,N_8249);
nor U9149 (N_9149,N_7650,N_7691);
and U9150 (N_9150,N_7520,N_8578);
and U9151 (N_9151,N_7986,N_7548);
xor U9152 (N_9152,N_8061,N_8478);
nand U9153 (N_9153,N_8711,N_8649);
or U9154 (N_9154,N_7806,N_8263);
nand U9155 (N_9155,N_8178,N_8349);
or U9156 (N_9156,N_8329,N_8239);
and U9157 (N_9157,N_7605,N_7785);
and U9158 (N_9158,N_7552,N_8733);
xnor U9159 (N_9159,N_8580,N_7778);
or U9160 (N_9160,N_7834,N_8272);
or U9161 (N_9161,N_7506,N_8101);
xor U9162 (N_9162,N_8618,N_8323);
nand U9163 (N_9163,N_8748,N_7889);
and U9164 (N_9164,N_7792,N_7850);
and U9165 (N_9165,N_8667,N_7714);
xnor U9166 (N_9166,N_8099,N_7838);
nand U9167 (N_9167,N_8264,N_8549);
and U9168 (N_9168,N_8621,N_8175);
nand U9169 (N_9169,N_8356,N_8255);
nor U9170 (N_9170,N_7864,N_7623);
nor U9171 (N_9171,N_7562,N_8140);
or U9172 (N_9172,N_8177,N_8411);
or U9173 (N_9173,N_8208,N_8690);
or U9174 (N_9174,N_8505,N_8473);
xor U9175 (N_9175,N_7571,N_8326);
and U9176 (N_9176,N_7641,N_7639);
xor U9177 (N_9177,N_7978,N_7601);
nor U9178 (N_9178,N_8197,N_8165);
and U9179 (N_9179,N_7582,N_8304);
nand U9180 (N_9180,N_8082,N_7920);
nand U9181 (N_9181,N_7793,N_8121);
and U9182 (N_9182,N_7573,N_8282);
xnor U9183 (N_9183,N_7880,N_8674);
nor U9184 (N_9184,N_8435,N_8374);
and U9185 (N_9185,N_8135,N_8502);
nor U9186 (N_9186,N_8522,N_8605);
nand U9187 (N_9187,N_8577,N_8685);
xor U9188 (N_9188,N_8100,N_7606);
nand U9189 (N_9189,N_8169,N_8410);
or U9190 (N_9190,N_8570,N_8483);
xor U9191 (N_9191,N_7620,N_8242);
xnor U9192 (N_9192,N_8019,N_8157);
or U9193 (N_9193,N_8120,N_8290);
nor U9194 (N_9194,N_8424,N_8737);
or U9195 (N_9195,N_8048,N_8275);
nand U9196 (N_9196,N_8510,N_8432);
nand U9197 (N_9197,N_7832,N_7935);
nor U9198 (N_9198,N_8689,N_8008);
and U9199 (N_9199,N_7787,N_7501);
and U9200 (N_9200,N_7764,N_7660);
xor U9201 (N_9201,N_8511,N_8537);
and U9202 (N_9202,N_7790,N_8187);
xnor U9203 (N_9203,N_8646,N_7627);
and U9204 (N_9204,N_7773,N_8507);
nand U9205 (N_9205,N_8325,N_7719);
and U9206 (N_9206,N_8085,N_8287);
xor U9207 (N_9207,N_8037,N_7721);
xor U9208 (N_9208,N_7649,N_8052);
xnor U9209 (N_9209,N_7572,N_7521);
xor U9210 (N_9210,N_7816,N_8434);
nor U9211 (N_9211,N_8713,N_7630);
or U9212 (N_9212,N_7509,N_7726);
nor U9213 (N_9213,N_8113,N_8585);
and U9214 (N_9214,N_7643,N_8565);
nor U9215 (N_9215,N_8542,N_7531);
and U9216 (N_9216,N_8029,N_7779);
or U9217 (N_9217,N_8602,N_8430);
xor U9218 (N_9218,N_8366,N_8036);
nand U9219 (N_9219,N_7813,N_7763);
nor U9220 (N_9220,N_8010,N_7722);
nand U9221 (N_9221,N_7611,N_7810);
and U9222 (N_9222,N_7737,N_7694);
or U9223 (N_9223,N_7857,N_7585);
and U9224 (N_9224,N_8377,N_7842);
and U9225 (N_9225,N_7836,N_8300);
nor U9226 (N_9226,N_7608,N_8704);
xnor U9227 (N_9227,N_8682,N_8742);
xor U9228 (N_9228,N_7570,N_8645);
and U9229 (N_9229,N_7846,N_8741);
nor U9230 (N_9230,N_8207,N_8011);
and U9231 (N_9231,N_7974,N_7768);
xor U9232 (N_9232,N_8555,N_8047);
and U9233 (N_9233,N_8091,N_8126);
and U9234 (N_9234,N_7720,N_7906);
xnor U9235 (N_9235,N_7591,N_8237);
and U9236 (N_9236,N_8609,N_7994);
nand U9237 (N_9237,N_7776,N_7689);
nor U9238 (N_9238,N_7971,N_7784);
and U9239 (N_9239,N_8243,N_8552);
xor U9240 (N_9240,N_8404,N_8241);
xnor U9241 (N_9241,N_7782,N_7913);
nor U9242 (N_9242,N_8106,N_8358);
xnor U9243 (N_9243,N_8684,N_8710);
nor U9244 (N_9244,N_8736,N_8073);
xnor U9245 (N_9245,N_8003,N_7931);
nand U9246 (N_9246,N_7998,N_7762);
or U9247 (N_9247,N_8648,N_8724);
or U9248 (N_9248,N_7752,N_8453);
nor U9249 (N_9249,N_8133,N_7970);
and U9250 (N_9250,N_8086,N_7990);
nor U9251 (N_9251,N_8189,N_8344);
xnor U9252 (N_9252,N_8394,N_7960);
xor U9253 (N_9253,N_8122,N_7603);
nand U9254 (N_9254,N_7675,N_7821);
xor U9255 (N_9255,N_7563,N_8236);
or U9256 (N_9256,N_7637,N_8612);
or U9257 (N_9257,N_8320,N_8513);
or U9258 (N_9258,N_7526,N_8440);
nor U9259 (N_9259,N_8218,N_8503);
and U9260 (N_9260,N_8090,N_7659);
and U9261 (N_9261,N_8450,N_7663);
and U9262 (N_9262,N_8652,N_8423);
and U9263 (N_9263,N_8138,N_8305);
and U9264 (N_9264,N_7615,N_8163);
nor U9265 (N_9265,N_7829,N_8235);
xor U9266 (N_9266,N_8601,N_8379);
nor U9267 (N_9267,N_8016,N_8199);
nand U9268 (N_9268,N_7826,N_7736);
nor U9269 (N_9269,N_7595,N_8292);
xor U9270 (N_9270,N_8103,N_7734);
nor U9271 (N_9271,N_8225,N_7642);
or U9272 (N_9272,N_8541,N_7751);
nor U9273 (N_9273,N_7879,N_7860);
and U9274 (N_9274,N_8299,N_8142);
xor U9275 (N_9275,N_8045,N_8051);
or U9276 (N_9276,N_8193,N_8584);
and U9277 (N_9277,N_8340,N_8623);
nand U9278 (N_9278,N_7727,N_8396);
nand U9279 (N_9279,N_8069,N_8656);
or U9280 (N_9280,N_7541,N_8603);
nor U9281 (N_9281,N_8294,N_8104);
xnor U9282 (N_9282,N_8487,N_7896);
nor U9283 (N_9283,N_7504,N_8481);
and U9284 (N_9284,N_8668,N_8467);
or U9285 (N_9285,N_8499,N_8461);
or U9286 (N_9286,N_8152,N_8417);
nand U9287 (N_9287,N_8658,N_8509);
xor U9288 (N_9288,N_7780,N_8368);
or U9289 (N_9289,N_7924,N_8528);
xnor U9290 (N_9290,N_7922,N_7997);
or U9291 (N_9291,N_8179,N_7514);
nor U9292 (N_9292,N_8196,N_8579);
nand U9293 (N_9293,N_7511,N_8015);
and U9294 (N_9294,N_8056,N_7545);
or U9295 (N_9295,N_7899,N_7815);
nand U9296 (N_9296,N_7830,N_8372);
nor U9297 (N_9297,N_7903,N_8002);
and U9298 (N_9298,N_7670,N_8107);
nand U9299 (N_9299,N_8701,N_7686);
or U9300 (N_9300,N_7817,N_8020);
and U9301 (N_9301,N_7972,N_8600);
xor U9302 (N_9302,N_8301,N_7819);
nor U9303 (N_9303,N_7718,N_8514);
or U9304 (N_9304,N_8146,N_7550);
nand U9305 (N_9305,N_8526,N_7647);
nand U9306 (N_9306,N_7672,N_7709);
nand U9307 (N_9307,N_8289,N_7950);
or U9308 (N_9308,N_8184,N_8343);
or U9309 (N_9309,N_7558,N_7669);
nand U9310 (N_9310,N_8657,N_8383);
and U9311 (N_9311,N_8466,N_7945);
xor U9312 (N_9312,N_8162,N_7794);
nand U9313 (N_9313,N_8698,N_8096);
and U9314 (N_9314,N_8155,N_7969);
nor U9315 (N_9315,N_8556,N_8594);
nor U9316 (N_9316,N_8270,N_8705);
nand U9317 (N_9317,N_8443,N_8068);
nand U9318 (N_9318,N_7679,N_8614);
xor U9319 (N_9319,N_8205,N_7873);
or U9320 (N_9320,N_8111,N_8046);
xor U9321 (N_9321,N_7966,N_8319);
and U9322 (N_9322,N_7804,N_8489);
nor U9323 (N_9323,N_8116,N_8633);
and U9324 (N_9324,N_7698,N_8317);
nor U9325 (N_9325,N_8077,N_8426);
and U9326 (N_9326,N_8563,N_8615);
xor U9327 (N_9327,N_8665,N_8127);
nor U9328 (N_9328,N_8672,N_8006);
xnor U9329 (N_9329,N_8534,N_7744);
nand U9330 (N_9330,N_8337,N_8546);
and U9331 (N_9331,N_7992,N_8532);
and U9332 (N_9332,N_7657,N_8639);
nor U9333 (N_9333,N_8494,N_8141);
and U9334 (N_9334,N_7594,N_8164);
nor U9335 (N_9335,N_7692,N_7835);
or U9336 (N_9336,N_7833,N_7557);
nand U9337 (N_9337,N_7895,N_8302);
and U9338 (N_9338,N_8123,N_7688);
nand U9339 (N_9339,N_8186,N_7956);
nor U9340 (N_9340,N_7750,N_8728);
xnor U9341 (N_9341,N_8361,N_7651);
nor U9342 (N_9342,N_8387,N_7527);
or U9343 (N_9343,N_8653,N_8013);
nor U9344 (N_9344,N_8055,N_8384);
nand U9345 (N_9345,N_8606,N_8715);
or U9346 (N_9346,N_8460,N_8465);
nor U9347 (N_9347,N_8593,N_8252);
xnor U9348 (N_9348,N_7975,N_7640);
or U9349 (N_9349,N_7909,N_7602);
or U9350 (N_9350,N_8571,N_8515);
nand U9351 (N_9351,N_7979,N_7668);
nand U9352 (N_9352,N_8033,N_7730);
and U9353 (N_9353,N_8378,N_7542);
and U9354 (N_9354,N_8194,N_8332);
nor U9355 (N_9355,N_7740,N_8670);
nand U9356 (N_9356,N_8589,N_8025);
nor U9357 (N_9357,N_8484,N_8044);
xor U9358 (N_9358,N_8324,N_8714);
and U9359 (N_9359,N_7656,N_8124);
or U9360 (N_9360,N_8108,N_8057);
or U9361 (N_9361,N_7731,N_8548);
xnor U9362 (N_9362,N_8501,N_8132);
nand U9363 (N_9363,N_7984,N_8362);
nand U9364 (N_9364,N_7907,N_8180);
nand U9365 (N_9365,N_7638,N_8477);
xnor U9366 (N_9366,N_7805,N_8067);
and U9367 (N_9367,N_8350,N_8190);
or U9368 (N_9368,N_8681,N_7539);
xnor U9369 (N_9369,N_8143,N_8083);
and U9370 (N_9370,N_8490,N_7807);
nand U9371 (N_9371,N_8538,N_8217);
nor U9372 (N_9372,N_7624,N_7758);
nor U9373 (N_9373,N_7684,N_8586);
nand U9374 (N_9374,N_8212,N_8303);
nand U9375 (N_9375,N_8276,N_8587);
nor U9376 (N_9376,N_8442,N_8590);
nor U9377 (N_9377,N_8735,N_8012);
xor U9378 (N_9378,N_7926,N_8673);
nor U9379 (N_9379,N_7729,N_8418);
nand U9380 (N_9380,N_7953,N_8178);
nor U9381 (N_9381,N_7568,N_7886);
nor U9382 (N_9382,N_8143,N_7996);
xnor U9383 (N_9383,N_7586,N_7887);
nor U9384 (N_9384,N_8704,N_8361);
xor U9385 (N_9385,N_7735,N_8066);
xnor U9386 (N_9386,N_7513,N_7963);
nor U9387 (N_9387,N_7669,N_8334);
and U9388 (N_9388,N_7551,N_7507);
or U9389 (N_9389,N_7526,N_8360);
nor U9390 (N_9390,N_8631,N_7836);
nor U9391 (N_9391,N_7764,N_7599);
or U9392 (N_9392,N_8502,N_8080);
xnor U9393 (N_9393,N_7836,N_8297);
nand U9394 (N_9394,N_7999,N_8062);
and U9395 (N_9395,N_8695,N_7693);
xor U9396 (N_9396,N_8146,N_8458);
nor U9397 (N_9397,N_8351,N_8154);
and U9398 (N_9398,N_7830,N_7812);
nor U9399 (N_9399,N_8333,N_7894);
nor U9400 (N_9400,N_7980,N_7616);
nand U9401 (N_9401,N_7729,N_7589);
xnor U9402 (N_9402,N_8127,N_8078);
nor U9403 (N_9403,N_8232,N_8557);
nand U9404 (N_9404,N_7621,N_8608);
and U9405 (N_9405,N_8727,N_7702);
nand U9406 (N_9406,N_7696,N_7656);
nand U9407 (N_9407,N_8086,N_7806);
and U9408 (N_9408,N_8706,N_7815);
nand U9409 (N_9409,N_8492,N_8616);
xnor U9410 (N_9410,N_7784,N_7871);
and U9411 (N_9411,N_8164,N_8039);
and U9412 (N_9412,N_8191,N_7717);
nor U9413 (N_9413,N_7683,N_7828);
or U9414 (N_9414,N_8124,N_8402);
and U9415 (N_9415,N_8300,N_7896);
xnor U9416 (N_9416,N_8157,N_8588);
and U9417 (N_9417,N_8226,N_7990);
and U9418 (N_9418,N_7714,N_7988);
or U9419 (N_9419,N_8439,N_8025);
xnor U9420 (N_9420,N_8590,N_7945);
or U9421 (N_9421,N_8259,N_7957);
nand U9422 (N_9422,N_8489,N_8259);
xnor U9423 (N_9423,N_8505,N_7559);
nand U9424 (N_9424,N_8559,N_8325);
nor U9425 (N_9425,N_7538,N_8426);
nand U9426 (N_9426,N_7609,N_7589);
nor U9427 (N_9427,N_7840,N_8567);
nand U9428 (N_9428,N_8230,N_8240);
and U9429 (N_9429,N_8231,N_8608);
or U9430 (N_9430,N_7540,N_7509);
nor U9431 (N_9431,N_7675,N_7867);
xnor U9432 (N_9432,N_8508,N_7968);
or U9433 (N_9433,N_7574,N_8052);
and U9434 (N_9434,N_8742,N_7549);
nor U9435 (N_9435,N_8667,N_8202);
xnor U9436 (N_9436,N_7747,N_8034);
xor U9437 (N_9437,N_7697,N_8557);
and U9438 (N_9438,N_7607,N_8621);
xnor U9439 (N_9439,N_8523,N_8134);
xnor U9440 (N_9440,N_8404,N_8612);
xnor U9441 (N_9441,N_8481,N_7562);
or U9442 (N_9442,N_8623,N_7723);
xnor U9443 (N_9443,N_7608,N_7862);
xor U9444 (N_9444,N_7849,N_8599);
or U9445 (N_9445,N_7932,N_7814);
nand U9446 (N_9446,N_7616,N_8404);
and U9447 (N_9447,N_7869,N_7528);
and U9448 (N_9448,N_7808,N_7949);
and U9449 (N_9449,N_7940,N_8344);
or U9450 (N_9450,N_8488,N_8238);
and U9451 (N_9451,N_8546,N_7985);
nand U9452 (N_9452,N_8425,N_8114);
or U9453 (N_9453,N_7766,N_8196);
xnor U9454 (N_9454,N_7551,N_8154);
nor U9455 (N_9455,N_8667,N_8427);
xnor U9456 (N_9456,N_8612,N_7959);
and U9457 (N_9457,N_8399,N_7668);
nand U9458 (N_9458,N_8508,N_8736);
nor U9459 (N_9459,N_8694,N_8326);
or U9460 (N_9460,N_8245,N_8304);
or U9461 (N_9461,N_7876,N_8034);
nor U9462 (N_9462,N_8296,N_8191);
xor U9463 (N_9463,N_8245,N_8081);
nand U9464 (N_9464,N_7938,N_7548);
nor U9465 (N_9465,N_8072,N_8533);
or U9466 (N_9466,N_8655,N_8336);
nor U9467 (N_9467,N_8068,N_8694);
and U9468 (N_9468,N_8358,N_8003);
nand U9469 (N_9469,N_7816,N_8412);
nand U9470 (N_9470,N_8191,N_8015);
and U9471 (N_9471,N_8566,N_8127);
xnor U9472 (N_9472,N_8275,N_7622);
xnor U9473 (N_9473,N_8260,N_7820);
and U9474 (N_9474,N_7883,N_7918);
xnor U9475 (N_9475,N_7824,N_8687);
nand U9476 (N_9476,N_7747,N_8102);
or U9477 (N_9477,N_7835,N_8507);
xnor U9478 (N_9478,N_7562,N_8391);
nor U9479 (N_9479,N_7545,N_8201);
nand U9480 (N_9480,N_8736,N_7506);
and U9481 (N_9481,N_8026,N_8068);
or U9482 (N_9482,N_7575,N_8232);
xnor U9483 (N_9483,N_7503,N_7968);
xnor U9484 (N_9484,N_8006,N_7998);
nand U9485 (N_9485,N_8192,N_8457);
and U9486 (N_9486,N_8018,N_8197);
xor U9487 (N_9487,N_8714,N_8669);
nor U9488 (N_9488,N_8653,N_8320);
or U9489 (N_9489,N_8008,N_7637);
or U9490 (N_9490,N_8149,N_7690);
nand U9491 (N_9491,N_8417,N_7689);
nand U9492 (N_9492,N_8106,N_7669);
or U9493 (N_9493,N_8444,N_7866);
nor U9494 (N_9494,N_7573,N_8292);
nor U9495 (N_9495,N_7721,N_8410);
nor U9496 (N_9496,N_7554,N_7836);
xnor U9497 (N_9497,N_7835,N_8492);
nand U9498 (N_9498,N_8107,N_8046);
and U9499 (N_9499,N_8204,N_8707);
nor U9500 (N_9500,N_8451,N_8455);
nand U9501 (N_9501,N_7610,N_8407);
and U9502 (N_9502,N_8413,N_8573);
or U9503 (N_9503,N_8520,N_7628);
xor U9504 (N_9504,N_7872,N_8253);
or U9505 (N_9505,N_8441,N_8370);
xor U9506 (N_9506,N_7628,N_8180);
xnor U9507 (N_9507,N_7593,N_8640);
and U9508 (N_9508,N_8239,N_7553);
nor U9509 (N_9509,N_8153,N_8697);
nand U9510 (N_9510,N_7569,N_7952);
xor U9511 (N_9511,N_8322,N_8666);
or U9512 (N_9512,N_7559,N_7629);
or U9513 (N_9513,N_7606,N_7769);
and U9514 (N_9514,N_8125,N_8397);
and U9515 (N_9515,N_8328,N_8072);
nor U9516 (N_9516,N_8284,N_7879);
and U9517 (N_9517,N_8207,N_7897);
nor U9518 (N_9518,N_8486,N_8745);
or U9519 (N_9519,N_7565,N_8491);
nand U9520 (N_9520,N_7664,N_8218);
and U9521 (N_9521,N_7728,N_7710);
nand U9522 (N_9522,N_8045,N_7548);
xnor U9523 (N_9523,N_8593,N_8109);
xor U9524 (N_9524,N_7823,N_8504);
or U9525 (N_9525,N_8381,N_7589);
nand U9526 (N_9526,N_8466,N_8378);
and U9527 (N_9527,N_8319,N_7515);
nor U9528 (N_9528,N_8101,N_8418);
nand U9529 (N_9529,N_8590,N_8594);
nand U9530 (N_9530,N_8524,N_8364);
nand U9531 (N_9531,N_7908,N_8324);
nand U9532 (N_9532,N_8279,N_7994);
xor U9533 (N_9533,N_8022,N_8743);
and U9534 (N_9534,N_8116,N_7635);
nand U9535 (N_9535,N_7947,N_8243);
nor U9536 (N_9536,N_8415,N_7749);
and U9537 (N_9537,N_8410,N_7864);
xnor U9538 (N_9538,N_7920,N_8450);
nand U9539 (N_9539,N_7958,N_7562);
xnor U9540 (N_9540,N_7938,N_8155);
nor U9541 (N_9541,N_8325,N_7837);
nor U9542 (N_9542,N_8486,N_8320);
nor U9543 (N_9543,N_7759,N_7641);
xor U9544 (N_9544,N_8109,N_7968);
and U9545 (N_9545,N_8105,N_8230);
or U9546 (N_9546,N_8435,N_8651);
nand U9547 (N_9547,N_8182,N_8615);
xor U9548 (N_9548,N_7697,N_8648);
and U9549 (N_9549,N_8541,N_8038);
or U9550 (N_9550,N_7903,N_8419);
nand U9551 (N_9551,N_8480,N_8203);
or U9552 (N_9552,N_7689,N_8144);
and U9553 (N_9553,N_8403,N_8722);
or U9554 (N_9554,N_7532,N_7675);
nor U9555 (N_9555,N_7640,N_7921);
xnor U9556 (N_9556,N_8720,N_8461);
or U9557 (N_9557,N_8163,N_7986);
xor U9558 (N_9558,N_8646,N_8699);
xor U9559 (N_9559,N_8714,N_7653);
and U9560 (N_9560,N_7961,N_7550);
nand U9561 (N_9561,N_8710,N_8592);
or U9562 (N_9562,N_8497,N_8565);
xnor U9563 (N_9563,N_8428,N_8423);
xnor U9564 (N_9564,N_8023,N_8630);
nand U9565 (N_9565,N_7934,N_8379);
and U9566 (N_9566,N_7710,N_7757);
nor U9567 (N_9567,N_7544,N_7839);
nand U9568 (N_9568,N_7991,N_8120);
nor U9569 (N_9569,N_7933,N_8344);
and U9570 (N_9570,N_7538,N_7503);
nor U9571 (N_9571,N_8042,N_7609);
or U9572 (N_9572,N_7733,N_7539);
nor U9573 (N_9573,N_8367,N_8428);
xor U9574 (N_9574,N_8729,N_8447);
xor U9575 (N_9575,N_8245,N_7514);
nor U9576 (N_9576,N_7610,N_8722);
xnor U9577 (N_9577,N_8174,N_7809);
or U9578 (N_9578,N_8689,N_8323);
nor U9579 (N_9579,N_8698,N_8263);
nor U9580 (N_9580,N_7773,N_7651);
and U9581 (N_9581,N_8402,N_7682);
or U9582 (N_9582,N_8222,N_7527);
nor U9583 (N_9583,N_7766,N_8339);
nor U9584 (N_9584,N_8168,N_7887);
or U9585 (N_9585,N_8435,N_8729);
nor U9586 (N_9586,N_8710,N_7982);
and U9587 (N_9587,N_8209,N_8078);
nand U9588 (N_9588,N_7887,N_7971);
and U9589 (N_9589,N_8419,N_8420);
nor U9590 (N_9590,N_8731,N_7871);
nand U9591 (N_9591,N_8096,N_8609);
nand U9592 (N_9592,N_7697,N_8257);
and U9593 (N_9593,N_7541,N_7752);
xor U9594 (N_9594,N_8190,N_8655);
nor U9595 (N_9595,N_7925,N_8523);
or U9596 (N_9596,N_8008,N_7838);
nor U9597 (N_9597,N_8128,N_8241);
nor U9598 (N_9598,N_8523,N_7637);
nand U9599 (N_9599,N_8019,N_7746);
nor U9600 (N_9600,N_7562,N_8081);
nor U9601 (N_9601,N_7620,N_7544);
or U9602 (N_9602,N_8508,N_7566);
xor U9603 (N_9603,N_7853,N_7637);
xnor U9604 (N_9604,N_8081,N_7999);
xor U9605 (N_9605,N_8449,N_8399);
xnor U9606 (N_9606,N_8238,N_8595);
nand U9607 (N_9607,N_8441,N_8363);
or U9608 (N_9608,N_8730,N_8743);
or U9609 (N_9609,N_8199,N_7536);
nor U9610 (N_9610,N_8680,N_7681);
or U9611 (N_9611,N_8315,N_8387);
and U9612 (N_9612,N_8661,N_8362);
or U9613 (N_9613,N_7556,N_8078);
and U9614 (N_9614,N_7528,N_8446);
and U9615 (N_9615,N_7969,N_7921);
nand U9616 (N_9616,N_8712,N_7904);
xnor U9617 (N_9617,N_7980,N_8743);
or U9618 (N_9618,N_7554,N_7953);
or U9619 (N_9619,N_8378,N_8488);
xor U9620 (N_9620,N_8282,N_8618);
or U9621 (N_9621,N_8315,N_7521);
or U9622 (N_9622,N_8065,N_7912);
nor U9623 (N_9623,N_8486,N_8548);
nand U9624 (N_9624,N_8635,N_8467);
nor U9625 (N_9625,N_8093,N_8031);
nor U9626 (N_9626,N_8267,N_7528);
nor U9627 (N_9627,N_7862,N_7847);
and U9628 (N_9628,N_7999,N_7862);
nand U9629 (N_9629,N_7509,N_8476);
or U9630 (N_9630,N_8073,N_8249);
or U9631 (N_9631,N_7587,N_7692);
and U9632 (N_9632,N_7688,N_7861);
nor U9633 (N_9633,N_8003,N_8420);
and U9634 (N_9634,N_7637,N_8056);
nor U9635 (N_9635,N_7665,N_7510);
and U9636 (N_9636,N_7822,N_7733);
nor U9637 (N_9637,N_7716,N_8080);
xnor U9638 (N_9638,N_8198,N_8137);
and U9639 (N_9639,N_7893,N_8205);
xor U9640 (N_9640,N_8663,N_8581);
or U9641 (N_9641,N_8156,N_7995);
nand U9642 (N_9642,N_7515,N_7540);
and U9643 (N_9643,N_7764,N_7623);
or U9644 (N_9644,N_8345,N_8446);
or U9645 (N_9645,N_8087,N_7916);
and U9646 (N_9646,N_8348,N_8400);
and U9647 (N_9647,N_7983,N_8147);
and U9648 (N_9648,N_8737,N_8252);
xor U9649 (N_9649,N_8118,N_7618);
nor U9650 (N_9650,N_8258,N_8209);
nand U9651 (N_9651,N_8058,N_8703);
and U9652 (N_9652,N_8355,N_8209);
and U9653 (N_9653,N_8593,N_8164);
or U9654 (N_9654,N_7676,N_7744);
or U9655 (N_9655,N_7947,N_7863);
nand U9656 (N_9656,N_8352,N_7959);
and U9657 (N_9657,N_8619,N_8126);
and U9658 (N_9658,N_8187,N_8281);
nand U9659 (N_9659,N_8689,N_8214);
nand U9660 (N_9660,N_7637,N_8352);
xnor U9661 (N_9661,N_7573,N_7652);
xor U9662 (N_9662,N_7733,N_7747);
nor U9663 (N_9663,N_8353,N_8403);
or U9664 (N_9664,N_8653,N_7953);
nor U9665 (N_9665,N_8308,N_7598);
or U9666 (N_9666,N_8481,N_8252);
xnor U9667 (N_9667,N_8387,N_8268);
nor U9668 (N_9668,N_8728,N_8558);
or U9669 (N_9669,N_7732,N_8584);
nor U9670 (N_9670,N_7993,N_7974);
nor U9671 (N_9671,N_8600,N_7944);
nor U9672 (N_9672,N_8565,N_8173);
or U9673 (N_9673,N_7567,N_8310);
or U9674 (N_9674,N_8593,N_8454);
and U9675 (N_9675,N_7516,N_8265);
and U9676 (N_9676,N_7715,N_8520);
xnor U9677 (N_9677,N_8229,N_8414);
nor U9678 (N_9678,N_7967,N_8150);
nand U9679 (N_9679,N_7930,N_8407);
or U9680 (N_9680,N_8350,N_8484);
nor U9681 (N_9681,N_8091,N_7864);
nand U9682 (N_9682,N_7590,N_7917);
nor U9683 (N_9683,N_8232,N_7999);
and U9684 (N_9684,N_7522,N_7563);
nor U9685 (N_9685,N_8323,N_8210);
or U9686 (N_9686,N_7643,N_8529);
nand U9687 (N_9687,N_7996,N_7822);
or U9688 (N_9688,N_7850,N_8097);
xnor U9689 (N_9689,N_7533,N_8307);
nand U9690 (N_9690,N_8400,N_8069);
nor U9691 (N_9691,N_8079,N_7758);
xor U9692 (N_9692,N_7586,N_8048);
or U9693 (N_9693,N_7787,N_8482);
and U9694 (N_9694,N_7728,N_8469);
nand U9695 (N_9695,N_7895,N_7766);
nand U9696 (N_9696,N_8255,N_8049);
and U9697 (N_9697,N_7872,N_8302);
nor U9698 (N_9698,N_8532,N_7636);
nor U9699 (N_9699,N_8404,N_7971);
nand U9700 (N_9700,N_8129,N_8393);
nor U9701 (N_9701,N_8005,N_7555);
nor U9702 (N_9702,N_8392,N_7511);
nand U9703 (N_9703,N_8264,N_7624);
and U9704 (N_9704,N_8740,N_8655);
or U9705 (N_9705,N_8518,N_8134);
nor U9706 (N_9706,N_8444,N_7591);
xor U9707 (N_9707,N_8453,N_7898);
or U9708 (N_9708,N_8019,N_7979);
and U9709 (N_9709,N_8381,N_8340);
or U9710 (N_9710,N_8016,N_8611);
nand U9711 (N_9711,N_8175,N_7502);
or U9712 (N_9712,N_8413,N_8583);
xnor U9713 (N_9713,N_7768,N_7868);
nand U9714 (N_9714,N_8543,N_7930);
nand U9715 (N_9715,N_7657,N_7648);
or U9716 (N_9716,N_7894,N_8437);
and U9717 (N_9717,N_8531,N_8534);
nand U9718 (N_9718,N_8056,N_7729);
or U9719 (N_9719,N_7796,N_8250);
nor U9720 (N_9720,N_8162,N_7864);
xnor U9721 (N_9721,N_8516,N_8078);
xor U9722 (N_9722,N_7755,N_8283);
nand U9723 (N_9723,N_7666,N_8049);
and U9724 (N_9724,N_8141,N_8215);
xor U9725 (N_9725,N_8435,N_8630);
or U9726 (N_9726,N_8078,N_7979);
xor U9727 (N_9727,N_8421,N_8028);
nand U9728 (N_9728,N_7582,N_8328);
nor U9729 (N_9729,N_7843,N_8374);
nor U9730 (N_9730,N_8626,N_8106);
and U9731 (N_9731,N_7681,N_8033);
or U9732 (N_9732,N_8472,N_7784);
or U9733 (N_9733,N_7556,N_8560);
and U9734 (N_9734,N_8072,N_8244);
or U9735 (N_9735,N_7915,N_8226);
nor U9736 (N_9736,N_8016,N_8405);
xnor U9737 (N_9737,N_8369,N_7667);
nand U9738 (N_9738,N_7724,N_8656);
and U9739 (N_9739,N_8229,N_8186);
nor U9740 (N_9740,N_7539,N_7606);
and U9741 (N_9741,N_8202,N_8081);
xor U9742 (N_9742,N_8265,N_7677);
nand U9743 (N_9743,N_7580,N_7535);
xnor U9744 (N_9744,N_7539,N_7886);
nor U9745 (N_9745,N_8547,N_7760);
nand U9746 (N_9746,N_7712,N_7949);
or U9747 (N_9747,N_7965,N_8038);
and U9748 (N_9748,N_8095,N_7717);
or U9749 (N_9749,N_8398,N_8311);
or U9750 (N_9750,N_7860,N_8559);
nor U9751 (N_9751,N_8039,N_8103);
nor U9752 (N_9752,N_8330,N_7778);
nor U9753 (N_9753,N_8247,N_8200);
xor U9754 (N_9754,N_8049,N_7733);
nand U9755 (N_9755,N_8462,N_8199);
xor U9756 (N_9756,N_8182,N_8511);
xor U9757 (N_9757,N_7729,N_8170);
xnor U9758 (N_9758,N_7510,N_7718);
nand U9759 (N_9759,N_7871,N_7669);
nand U9760 (N_9760,N_8460,N_8350);
nand U9761 (N_9761,N_8143,N_7843);
nor U9762 (N_9762,N_8729,N_8431);
and U9763 (N_9763,N_7761,N_8394);
and U9764 (N_9764,N_8550,N_7822);
and U9765 (N_9765,N_8704,N_8458);
xnor U9766 (N_9766,N_8314,N_7670);
xor U9767 (N_9767,N_7829,N_8616);
or U9768 (N_9768,N_8300,N_8384);
nand U9769 (N_9769,N_8378,N_8687);
nand U9770 (N_9770,N_8013,N_8146);
and U9771 (N_9771,N_7859,N_8415);
nor U9772 (N_9772,N_8730,N_8208);
and U9773 (N_9773,N_7632,N_8670);
or U9774 (N_9774,N_8105,N_7685);
nor U9775 (N_9775,N_7757,N_8079);
xnor U9776 (N_9776,N_7953,N_7536);
or U9777 (N_9777,N_8004,N_8483);
and U9778 (N_9778,N_8263,N_7864);
or U9779 (N_9779,N_8355,N_8415);
nand U9780 (N_9780,N_8237,N_8337);
and U9781 (N_9781,N_8419,N_7633);
and U9782 (N_9782,N_8415,N_8654);
and U9783 (N_9783,N_7511,N_8571);
nor U9784 (N_9784,N_8274,N_7907);
and U9785 (N_9785,N_8311,N_8661);
nor U9786 (N_9786,N_7538,N_8573);
or U9787 (N_9787,N_8635,N_8559);
nand U9788 (N_9788,N_7821,N_8744);
and U9789 (N_9789,N_7966,N_7862);
xnor U9790 (N_9790,N_8507,N_8387);
nand U9791 (N_9791,N_7755,N_8474);
xnor U9792 (N_9792,N_7765,N_7609);
and U9793 (N_9793,N_8029,N_7610);
nand U9794 (N_9794,N_7941,N_8256);
nor U9795 (N_9795,N_8742,N_7766);
and U9796 (N_9796,N_7928,N_8509);
and U9797 (N_9797,N_8554,N_7526);
nand U9798 (N_9798,N_8281,N_7855);
and U9799 (N_9799,N_7545,N_8739);
and U9800 (N_9800,N_8463,N_8338);
nor U9801 (N_9801,N_8498,N_7849);
and U9802 (N_9802,N_8535,N_8729);
nand U9803 (N_9803,N_7868,N_8076);
xor U9804 (N_9804,N_8385,N_7541);
and U9805 (N_9805,N_8490,N_7563);
nand U9806 (N_9806,N_8684,N_8419);
and U9807 (N_9807,N_8181,N_8480);
or U9808 (N_9808,N_8529,N_8565);
nand U9809 (N_9809,N_8479,N_8702);
xor U9810 (N_9810,N_8556,N_8090);
or U9811 (N_9811,N_8044,N_8586);
and U9812 (N_9812,N_8306,N_8589);
nor U9813 (N_9813,N_7570,N_8480);
or U9814 (N_9814,N_8717,N_7658);
xnor U9815 (N_9815,N_7764,N_8531);
nor U9816 (N_9816,N_7921,N_8192);
nand U9817 (N_9817,N_7947,N_7635);
nand U9818 (N_9818,N_7525,N_8663);
and U9819 (N_9819,N_8650,N_8311);
xor U9820 (N_9820,N_7730,N_8438);
nand U9821 (N_9821,N_8206,N_8080);
or U9822 (N_9822,N_8068,N_7789);
xnor U9823 (N_9823,N_8490,N_8567);
or U9824 (N_9824,N_7752,N_7744);
nor U9825 (N_9825,N_8246,N_8566);
xor U9826 (N_9826,N_8247,N_8033);
or U9827 (N_9827,N_8024,N_7509);
or U9828 (N_9828,N_8529,N_8089);
and U9829 (N_9829,N_8657,N_7808);
xnor U9830 (N_9830,N_7688,N_8747);
nand U9831 (N_9831,N_7749,N_7704);
and U9832 (N_9832,N_7776,N_7522);
or U9833 (N_9833,N_7929,N_8489);
or U9834 (N_9834,N_7833,N_8663);
or U9835 (N_9835,N_7941,N_8135);
nand U9836 (N_9836,N_8114,N_7950);
nor U9837 (N_9837,N_7784,N_7795);
or U9838 (N_9838,N_7691,N_8297);
nand U9839 (N_9839,N_8744,N_7806);
nor U9840 (N_9840,N_8066,N_8501);
nand U9841 (N_9841,N_8137,N_8031);
nand U9842 (N_9842,N_8402,N_8302);
and U9843 (N_9843,N_8451,N_8016);
nor U9844 (N_9844,N_7975,N_8465);
or U9845 (N_9845,N_8283,N_7698);
and U9846 (N_9846,N_7914,N_7869);
or U9847 (N_9847,N_8274,N_8077);
nor U9848 (N_9848,N_8459,N_8559);
and U9849 (N_9849,N_8306,N_8173);
or U9850 (N_9850,N_8382,N_7987);
xor U9851 (N_9851,N_8198,N_8681);
xor U9852 (N_9852,N_7718,N_7847);
xor U9853 (N_9853,N_7844,N_8613);
nand U9854 (N_9854,N_7992,N_8089);
or U9855 (N_9855,N_7955,N_8578);
nand U9856 (N_9856,N_8606,N_8161);
nor U9857 (N_9857,N_7906,N_8386);
and U9858 (N_9858,N_7903,N_7841);
or U9859 (N_9859,N_8550,N_7873);
xnor U9860 (N_9860,N_8258,N_7702);
nand U9861 (N_9861,N_7943,N_7704);
nand U9862 (N_9862,N_8711,N_8723);
and U9863 (N_9863,N_8647,N_8303);
nor U9864 (N_9864,N_7737,N_8357);
xnor U9865 (N_9865,N_7844,N_8379);
or U9866 (N_9866,N_8283,N_7593);
and U9867 (N_9867,N_8416,N_8722);
or U9868 (N_9868,N_7773,N_7980);
xor U9869 (N_9869,N_8224,N_8438);
nor U9870 (N_9870,N_8328,N_8344);
nor U9871 (N_9871,N_8389,N_7980);
nor U9872 (N_9872,N_8693,N_7626);
or U9873 (N_9873,N_7913,N_7691);
or U9874 (N_9874,N_8547,N_7781);
and U9875 (N_9875,N_8001,N_8075);
nand U9876 (N_9876,N_7893,N_8341);
nand U9877 (N_9877,N_8693,N_7793);
and U9878 (N_9878,N_8628,N_7991);
xor U9879 (N_9879,N_7858,N_8677);
and U9880 (N_9880,N_7735,N_7743);
xnor U9881 (N_9881,N_8012,N_7720);
nand U9882 (N_9882,N_8553,N_8599);
or U9883 (N_9883,N_7550,N_7763);
and U9884 (N_9884,N_7855,N_8545);
or U9885 (N_9885,N_8168,N_8475);
and U9886 (N_9886,N_8621,N_8410);
nand U9887 (N_9887,N_8261,N_7751);
nand U9888 (N_9888,N_8217,N_8215);
nand U9889 (N_9889,N_7865,N_7985);
xor U9890 (N_9890,N_8683,N_8705);
or U9891 (N_9891,N_8132,N_8148);
nand U9892 (N_9892,N_7579,N_7729);
nor U9893 (N_9893,N_8665,N_8644);
or U9894 (N_9894,N_8587,N_7612);
nor U9895 (N_9895,N_7782,N_8415);
nand U9896 (N_9896,N_7603,N_8431);
or U9897 (N_9897,N_8193,N_8137);
or U9898 (N_9898,N_8312,N_8475);
or U9899 (N_9899,N_8586,N_7603);
nand U9900 (N_9900,N_8695,N_7778);
and U9901 (N_9901,N_8608,N_8101);
nor U9902 (N_9902,N_8054,N_8055);
nand U9903 (N_9903,N_7984,N_8420);
nor U9904 (N_9904,N_8704,N_7615);
or U9905 (N_9905,N_7554,N_8418);
and U9906 (N_9906,N_8691,N_8092);
xnor U9907 (N_9907,N_8669,N_7688);
and U9908 (N_9908,N_7582,N_8550);
xor U9909 (N_9909,N_7817,N_7859);
xnor U9910 (N_9910,N_7991,N_8651);
nor U9911 (N_9911,N_7510,N_8208);
and U9912 (N_9912,N_7843,N_7939);
or U9913 (N_9913,N_8475,N_7762);
xor U9914 (N_9914,N_8280,N_8018);
and U9915 (N_9915,N_7956,N_7671);
nor U9916 (N_9916,N_7734,N_7773);
nand U9917 (N_9917,N_8482,N_8498);
xor U9918 (N_9918,N_8225,N_8507);
xor U9919 (N_9919,N_8647,N_7677);
xnor U9920 (N_9920,N_8144,N_8070);
or U9921 (N_9921,N_7622,N_8475);
and U9922 (N_9922,N_8378,N_8383);
xnor U9923 (N_9923,N_8608,N_8096);
or U9924 (N_9924,N_8197,N_7521);
nand U9925 (N_9925,N_8170,N_7561);
and U9926 (N_9926,N_7535,N_7528);
xor U9927 (N_9927,N_7993,N_8301);
or U9928 (N_9928,N_8584,N_7944);
xnor U9929 (N_9929,N_8423,N_7989);
and U9930 (N_9930,N_7941,N_8246);
nor U9931 (N_9931,N_8047,N_7831);
or U9932 (N_9932,N_7991,N_8680);
and U9933 (N_9933,N_8571,N_7788);
nor U9934 (N_9934,N_7571,N_7669);
xor U9935 (N_9935,N_8270,N_7500);
xor U9936 (N_9936,N_8440,N_8477);
and U9937 (N_9937,N_8656,N_7875);
or U9938 (N_9938,N_8182,N_8620);
xor U9939 (N_9939,N_7643,N_8326);
xnor U9940 (N_9940,N_7625,N_8344);
or U9941 (N_9941,N_8696,N_8254);
xnor U9942 (N_9942,N_8122,N_7803);
and U9943 (N_9943,N_8591,N_8559);
or U9944 (N_9944,N_7601,N_8462);
nor U9945 (N_9945,N_7987,N_8505);
nor U9946 (N_9946,N_8450,N_7515);
or U9947 (N_9947,N_7575,N_7526);
nand U9948 (N_9948,N_7521,N_8652);
nor U9949 (N_9949,N_7538,N_7774);
and U9950 (N_9950,N_8298,N_8016);
or U9951 (N_9951,N_8592,N_7590);
nand U9952 (N_9952,N_8586,N_8701);
nand U9953 (N_9953,N_7998,N_7637);
xor U9954 (N_9954,N_7794,N_8740);
xnor U9955 (N_9955,N_8029,N_8353);
nor U9956 (N_9956,N_7532,N_7521);
nor U9957 (N_9957,N_8564,N_8400);
nand U9958 (N_9958,N_8095,N_7667);
xnor U9959 (N_9959,N_8468,N_8272);
nand U9960 (N_9960,N_8463,N_8108);
and U9961 (N_9961,N_8477,N_7780);
and U9962 (N_9962,N_7883,N_7773);
and U9963 (N_9963,N_7894,N_8140);
nand U9964 (N_9964,N_8072,N_7794);
xor U9965 (N_9965,N_8415,N_7799);
nor U9966 (N_9966,N_8249,N_8681);
nand U9967 (N_9967,N_8701,N_7500);
nor U9968 (N_9968,N_7967,N_7541);
or U9969 (N_9969,N_7982,N_8421);
nor U9970 (N_9970,N_8552,N_8720);
nor U9971 (N_9971,N_8079,N_8388);
nand U9972 (N_9972,N_8183,N_7797);
nor U9973 (N_9973,N_8495,N_7532);
or U9974 (N_9974,N_8403,N_7597);
or U9975 (N_9975,N_8175,N_7767);
nor U9976 (N_9976,N_8117,N_8065);
nor U9977 (N_9977,N_7656,N_7801);
and U9978 (N_9978,N_8471,N_7659);
nor U9979 (N_9979,N_8541,N_7594);
or U9980 (N_9980,N_8176,N_8144);
or U9981 (N_9981,N_7919,N_7774);
or U9982 (N_9982,N_8196,N_8090);
xor U9983 (N_9983,N_7528,N_8022);
nor U9984 (N_9984,N_8169,N_8066);
or U9985 (N_9985,N_8742,N_7842);
or U9986 (N_9986,N_8308,N_8373);
and U9987 (N_9987,N_8230,N_7911);
nand U9988 (N_9988,N_8303,N_8552);
and U9989 (N_9989,N_7812,N_7560);
and U9990 (N_9990,N_7695,N_7523);
and U9991 (N_9991,N_8615,N_8099);
or U9992 (N_9992,N_7709,N_8400);
nor U9993 (N_9993,N_8608,N_7590);
and U9994 (N_9994,N_7760,N_7920);
nor U9995 (N_9995,N_7736,N_7687);
nor U9996 (N_9996,N_7779,N_8414);
or U9997 (N_9997,N_8253,N_8370);
nor U9998 (N_9998,N_7500,N_7596);
xnor U9999 (N_9999,N_7600,N_7526);
nand U10000 (N_10000,N_9623,N_9738);
nor U10001 (N_10001,N_9837,N_9242);
nor U10002 (N_10002,N_8864,N_9880);
and U10003 (N_10003,N_9686,N_9504);
nor U10004 (N_10004,N_9702,N_9443);
or U10005 (N_10005,N_9913,N_8976);
nand U10006 (N_10006,N_9775,N_9148);
nor U10007 (N_10007,N_9424,N_9706);
nor U10008 (N_10008,N_9399,N_9663);
xnor U10009 (N_10009,N_9402,N_8843);
xor U10010 (N_10010,N_9523,N_9867);
and U10011 (N_10011,N_9705,N_9013);
nand U10012 (N_10012,N_9394,N_8883);
or U10013 (N_10013,N_9754,N_8857);
nand U10014 (N_10014,N_9924,N_8850);
xnor U10015 (N_10015,N_8841,N_9935);
nor U10016 (N_10016,N_9547,N_9603);
nor U10017 (N_10017,N_9933,N_9866);
nand U10018 (N_10018,N_9747,N_9718);
nor U10019 (N_10019,N_9160,N_9561);
and U10020 (N_10020,N_9629,N_8980);
nand U10021 (N_10021,N_9959,N_9514);
or U10022 (N_10022,N_9423,N_9125);
and U10023 (N_10023,N_9591,N_9506);
or U10024 (N_10024,N_8760,N_8997);
xnor U10025 (N_10025,N_8984,N_9239);
nand U10026 (N_10026,N_9884,N_9051);
nand U10027 (N_10027,N_9908,N_9835);
nor U10028 (N_10028,N_9021,N_9109);
and U10029 (N_10029,N_9155,N_9627);
nor U10030 (N_10030,N_9464,N_9974);
and U10031 (N_10031,N_9293,N_8992);
xnor U10032 (N_10032,N_9206,N_8892);
xor U10033 (N_10033,N_9831,N_8898);
or U10034 (N_10034,N_9431,N_8855);
nand U10035 (N_10035,N_9784,N_9195);
and U10036 (N_10036,N_9819,N_8787);
nor U10037 (N_10037,N_9865,N_8777);
or U10038 (N_10038,N_9521,N_9066);
xor U10039 (N_10039,N_9720,N_9407);
and U10040 (N_10040,N_8758,N_9244);
nor U10041 (N_10041,N_9725,N_8948);
and U10042 (N_10042,N_8994,N_9951);
or U10043 (N_10043,N_9981,N_9681);
and U10044 (N_10044,N_9963,N_9077);
and U10045 (N_10045,N_9331,N_9224);
nand U10046 (N_10046,N_9783,N_9041);
or U10047 (N_10047,N_9765,N_9490);
or U10048 (N_10048,N_9961,N_9454);
nor U10049 (N_10049,N_9601,N_8937);
or U10050 (N_10050,N_8818,N_9126);
and U10051 (N_10051,N_9572,N_9220);
nand U10052 (N_10052,N_9513,N_9613);
nand U10053 (N_10053,N_8870,N_8869);
nor U10054 (N_10054,N_8830,N_8877);
xnor U10055 (N_10055,N_9232,N_9872);
nand U10056 (N_10056,N_8893,N_9903);
nor U10057 (N_10057,N_9914,N_9829);
nand U10058 (N_10058,N_9026,N_9893);
nor U10059 (N_10059,N_9729,N_9263);
and U10060 (N_10060,N_8833,N_8835);
and U10061 (N_10061,N_9216,N_9455);
or U10062 (N_10062,N_8968,N_9911);
nand U10063 (N_10063,N_9172,N_9578);
nor U10064 (N_10064,N_9215,N_8881);
xor U10065 (N_10065,N_9792,N_9577);
xor U10066 (N_10066,N_9973,N_9822);
nor U10067 (N_10067,N_9971,N_9522);
or U10068 (N_10068,N_9653,N_9201);
and U10069 (N_10069,N_9261,N_9171);
and U10070 (N_10070,N_9617,N_9833);
nor U10071 (N_10071,N_9698,N_9795);
nor U10072 (N_10072,N_9531,N_9062);
nand U10073 (N_10073,N_9248,N_9469);
nand U10074 (N_10074,N_9622,N_9839);
or U10075 (N_10075,N_9336,N_9417);
xor U10076 (N_10076,N_9061,N_9107);
and U10077 (N_10077,N_9344,N_9712);
nand U10078 (N_10078,N_9440,N_9910);
or U10079 (N_10079,N_9472,N_9983);
xnor U10080 (N_10080,N_9391,N_9587);
and U10081 (N_10081,N_9436,N_9868);
nand U10082 (N_10082,N_9310,N_8913);
and U10083 (N_10083,N_9750,N_9607);
and U10084 (N_10084,N_8813,N_9198);
xor U10085 (N_10085,N_9330,N_9323);
nand U10086 (N_10086,N_9058,N_9553);
nand U10087 (N_10087,N_9879,N_9213);
nor U10088 (N_10088,N_9098,N_9419);
and U10089 (N_10089,N_9921,N_9185);
or U10090 (N_10090,N_9102,N_9849);
nand U10091 (N_10091,N_8834,N_9088);
and U10092 (N_10092,N_9290,N_9429);
xor U10093 (N_10093,N_9453,N_9084);
and U10094 (N_10094,N_9002,N_9354);
xnor U10095 (N_10095,N_9489,N_9299);
or U10096 (N_10096,N_9709,N_9296);
nor U10097 (N_10097,N_9358,N_9333);
xnor U10098 (N_10098,N_9590,N_9116);
or U10099 (N_10099,N_9052,N_9965);
and U10100 (N_10100,N_9156,N_8908);
nor U10101 (N_10101,N_9138,N_9690);
nor U10102 (N_10102,N_9260,N_9448);
and U10103 (N_10103,N_9167,N_9934);
nor U10104 (N_10104,N_9928,N_9029);
xor U10105 (N_10105,N_9579,N_9497);
and U10106 (N_10106,N_9313,N_9281);
xnor U10107 (N_10107,N_9719,N_9063);
or U10108 (N_10108,N_9134,N_9153);
xor U10109 (N_10109,N_8923,N_9459);
xor U10110 (N_10110,N_9193,N_9863);
and U10111 (N_10111,N_9847,N_9298);
or U10112 (N_10112,N_8848,N_8823);
nor U10113 (N_10113,N_8921,N_9353);
xnor U10114 (N_10114,N_9977,N_9582);
xnor U10115 (N_10115,N_9007,N_8846);
and U10116 (N_10116,N_9673,N_9900);
xnor U10117 (N_10117,N_9962,N_8767);
and U10118 (N_10118,N_8889,N_9794);
nor U10119 (N_10119,N_9898,N_9165);
or U10120 (N_10120,N_9130,N_8924);
or U10121 (N_10121,N_9405,N_9787);
or U10122 (N_10122,N_9112,N_9069);
and U10123 (N_10123,N_9001,N_9192);
nand U10124 (N_10124,N_8847,N_9649);
nand U10125 (N_10125,N_9294,N_9487);
nand U10126 (N_10126,N_9095,N_9283);
and U10127 (N_10127,N_9647,N_9036);
xnor U10128 (N_10128,N_9003,N_9688);
or U10129 (N_10129,N_8915,N_8752);
nor U10130 (N_10130,N_9413,N_9624);
nor U10131 (N_10131,N_8790,N_9823);
nor U10132 (N_10132,N_9546,N_9289);
or U10133 (N_10133,N_9210,N_9039);
and U10134 (N_10134,N_9777,N_9078);
xor U10135 (N_10135,N_9748,N_8784);
or U10136 (N_10136,N_8819,N_9730);
nand U10137 (N_10137,N_9301,N_9105);
nor U10138 (N_10138,N_9997,N_8861);
or U10139 (N_10139,N_9483,N_9803);
or U10140 (N_10140,N_9559,N_9146);
and U10141 (N_10141,N_8868,N_9501);
xnor U10142 (N_10142,N_9231,N_8904);
xnor U10143 (N_10143,N_9179,N_9562);
nor U10144 (N_10144,N_9268,N_9945);
or U10145 (N_10145,N_9009,N_9498);
and U10146 (N_10146,N_9968,N_9732);
nand U10147 (N_10147,N_9957,N_9379);
and U10148 (N_10148,N_8955,N_9770);
xnor U10149 (N_10149,N_8945,N_9463);
and U10150 (N_10150,N_9687,N_8899);
xor U10151 (N_10151,N_9937,N_9357);
nor U10152 (N_10152,N_9633,N_9660);
or U10153 (N_10153,N_9876,N_9121);
and U10154 (N_10154,N_9269,N_8771);
and U10155 (N_10155,N_9644,N_9536);
nand U10156 (N_10156,N_9598,N_9801);
or U10157 (N_10157,N_9199,N_9420);
or U10158 (N_10158,N_9555,N_9986);
xnor U10159 (N_10159,N_8799,N_9466);
or U10160 (N_10160,N_9674,N_8990);
and U10161 (N_10161,N_8967,N_9669);
or U10162 (N_10162,N_8759,N_8845);
xor U10163 (N_10163,N_9131,N_9070);
nor U10164 (N_10164,N_8917,N_9438);
nand U10165 (N_10165,N_8936,N_9086);
and U10166 (N_10166,N_9626,N_8764);
nor U10167 (N_10167,N_8814,N_9312);
or U10168 (N_10168,N_9113,N_8981);
xor U10169 (N_10169,N_9948,N_9691);
nand U10170 (N_10170,N_9093,N_8977);
nand U10171 (N_10171,N_8878,N_9645);
nor U10172 (N_10172,N_8933,N_9122);
xor U10173 (N_10173,N_9208,N_9685);
nand U10174 (N_10174,N_9129,N_8902);
and U10175 (N_10175,N_8943,N_8789);
xor U10176 (N_10176,N_9592,N_8839);
nand U10177 (N_10177,N_9162,N_9790);
or U10178 (N_10178,N_9594,N_9442);
or U10179 (N_10179,N_8922,N_8803);
nand U10180 (N_10180,N_9573,N_9726);
nand U10181 (N_10181,N_9157,N_9650);
nand U10182 (N_10182,N_9169,N_9680);
nand U10183 (N_10183,N_9585,N_9264);
and U10184 (N_10184,N_9022,N_9288);
xnor U10185 (N_10185,N_9045,N_9796);
nand U10186 (N_10186,N_9306,N_9046);
or U10187 (N_10187,N_8912,N_8972);
nand U10188 (N_10188,N_9519,N_8873);
xor U10189 (N_10189,N_9825,N_9218);
nand U10190 (N_10190,N_9744,N_9178);
nor U10191 (N_10191,N_9307,N_9362);
and U10192 (N_10192,N_9348,N_9631);
and U10193 (N_10193,N_9300,N_8797);
nor U10194 (N_10194,N_9979,N_9988);
xnor U10195 (N_10195,N_9518,N_9999);
xnor U10196 (N_10196,N_9460,N_9050);
or U10197 (N_10197,N_9532,N_9858);
xor U10198 (N_10198,N_9495,N_8865);
or U10199 (N_10199,N_9017,N_9297);
nor U10200 (N_10200,N_9901,N_9196);
or U10201 (N_10201,N_9802,N_9895);
and U10202 (N_10202,N_8826,N_9149);
or U10203 (N_10203,N_9758,N_8811);
xor U10204 (N_10204,N_8932,N_9570);
nand U10205 (N_10205,N_9373,N_9387);
xor U10206 (N_10206,N_9856,N_9618);
nand U10207 (N_10207,N_8791,N_9241);
and U10208 (N_10208,N_9342,N_9485);
nand U10209 (N_10209,N_9068,N_9367);
or U10210 (N_10210,N_9860,N_9700);
xnor U10211 (N_10211,N_8775,N_9255);
or U10212 (N_10212,N_8754,N_9662);
or U10213 (N_10213,N_9378,N_9628);
nor U10214 (N_10214,N_9074,N_8989);
nor U10215 (N_10215,N_8930,N_9588);
nand U10216 (N_10216,N_9975,N_9275);
or U10217 (N_10217,N_9779,N_9119);
or U10218 (N_10218,N_9808,N_9509);
nor U10219 (N_10219,N_9083,N_9451);
nor U10220 (N_10220,N_8956,N_9966);
and U10221 (N_10221,N_9757,N_8970);
nor U10222 (N_10222,N_9987,N_8969);
or U10223 (N_10223,N_9304,N_8901);
and U10224 (N_10224,N_9564,N_9334);
nor U10225 (N_10225,N_9445,N_9818);
nor U10226 (N_10226,N_9541,N_9560);
and U10227 (N_10227,N_9529,N_8820);
nand U10228 (N_10228,N_9177,N_9717);
nor U10229 (N_10229,N_9780,N_8907);
or U10230 (N_10230,N_9551,N_8954);
or U10231 (N_10231,N_9549,N_9375);
nand U10232 (N_10232,N_9035,N_9788);
nand U10233 (N_10233,N_9222,N_9398);
xor U10234 (N_10234,N_8761,N_9659);
xor U10235 (N_10235,N_9094,N_9468);
and U10236 (N_10236,N_8838,N_9234);
nand U10237 (N_10237,N_9396,N_8974);
nor U10238 (N_10238,N_9535,N_9528);
and U10239 (N_10239,N_9851,N_8859);
or U10240 (N_10240,N_9651,N_9672);
and U10241 (N_10241,N_9015,N_9878);
nor U10242 (N_10242,N_9693,N_9595);
xnor U10243 (N_10243,N_9249,N_9484);
nand U10244 (N_10244,N_9597,N_9280);
nor U10245 (N_10245,N_9806,N_9363);
or U10246 (N_10246,N_8802,N_9891);
and U10247 (N_10247,N_8817,N_9144);
and U10248 (N_10248,N_9427,N_9871);
xor U10249 (N_10249,N_9145,N_9243);
and U10250 (N_10250,N_9655,N_9941);
xnor U10251 (N_10251,N_8996,N_9510);
nand U10252 (N_10252,N_9481,N_9656);
or U10253 (N_10253,N_9392,N_9376);
and U10254 (N_10254,N_9019,N_9616);
nor U10255 (N_10255,N_9230,N_8831);
xnor U10256 (N_10256,N_9952,N_9508);
or U10257 (N_10257,N_9332,N_9247);
nor U10258 (N_10258,N_9771,N_9727);
and U10259 (N_10259,N_9240,N_9110);
xnor U10260 (N_10260,N_9408,N_8858);
nor U10261 (N_10261,N_9733,N_9710);
nand U10262 (N_10262,N_9311,N_9273);
and U10263 (N_10263,N_9919,N_9677);
nor U10264 (N_10264,N_9768,N_9640);
or U10265 (N_10265,N_9414,N_9303);
nor U10266 (N_10266,N_9781,N_9400);
and U10267 (N_10267,N_9341,N_9814);
xor U10268 (N_10268,N_9743,N_9302);
xnor U10269 (N_10269,N_9187,N_8988);
nor U10270 (N_10270,N_8871,N_9173);
nand U10271 (N_10271,N_9204,N_9614);
or U10272 (N_10272,N_9772,N_8911);
nor U10273 (N_10273,N_9319,N_9740);
xnor U10274 (N_10274,N_9606,N_9071);
nand U10275 (N_10275,N_9619,N_9864);
nor U10276 (N_10276,N_9887,N_9734);
nand U10277 (N_10277,N_8934,N_9020);
xnor U10278 (N_10278,N_9569,N_9229);
or U10279 (N_10279,N_8832,N_8872);
nor U10280 (N_10280,N_9511,N_9761);
nand U10281 (N_10281,N_9753,N_9369);
nor U10282 (N_10282,N_8768,N_9478);
or U10283 (N_10283,N_9944,N_9888);
xor U10284 (N_10284,N_9128,N_9538);
nor U10285 (N_10285,N_9589,N_8903);
nor U10286 (N_10286,N_8900,N_8957);
and U10287 (N_10287,N_9393,N_9383);
or U10288 (N_10288,N_9540,N_9554);
and U10289 (N_10289,N_9949,N_9741);
and U10290 (N_10290,N_9221,N_9370);
nor U10291 (N_10291,N_9612,N_9256);
xor U10292 (N_10292,N_9175,N_8769);
and U10293 (N_10293,N_9776,N_9254);
nand U10294 (N_10294,N_8808,N_9972);
nor U10295 (N_10295,N_9053,N_9446);
or U10296 (N_10296,N_8800,N_9315);
or U10297 (N_10297,N_8765,N_9309);
or U10298 (N_10298,N_9024,N_9462);
and U10299 (N_10299,N_8793,N_9850);
nand U10300 (N_10300,N_9235,N_9181);
nand U10301 (N_10301,N_9998,N_9403);
nand U10302 (N_10302,N_9278,N_9339);
nand U10303 (N_10303,N_9343,N_9812);
nor U10304 (N_10304,N_9752,N_9883);
or U10305 (N_10305,N_9827,N_8876);
xor U10306 (N_10306,N_9324,N_9905);
or U10307 (N_10307,N_9166,N_9211);
or U10308 (N_10308,N_9286,N_9292);
nand U10309 (N_10309,N_9946,N_9507);
xnor U10310 (N_10310,N_9813,N_9412);
nand U10311 (N_10311,N_8986,N_8895);
nor U10312 (N_10312,N_9557,N_9409);
nand U10313 (N_10313,N_9896,N_9237);
xor U10314 (N_10314,N_9800,N_8897);
xor U10315 (N_10315,N_8905,N_9767);
nand U10316 (N_10316,N_9980,N_9090);
nand U10317 (N_10317,N_9075,N_9259);
nand U10318 (N_10318,N_9615,N_9713);
xor U10319 (N_10319,N_9347,N_8919);
nor U10320 (N_10320,N_8770,N_9525);
nand U10321 (N_10321,N_8983,N_8920);
and U10322 (N_10322,N_9586,N_8852);
or U10323 (N_10323,N_9227,N_9550);
nand U10324 (N_10324,N_9953,N_8815);
nand U10325 (N_10325,N_9843,N_8772);
nand U10326 (N_10326,N_9225,N_8860);
nand U10327 (N_10327,N_9217,N_8766);
and U10328 (N_10328,N_9205,N_9461);
and U10329 (N_10329,N_9912,N_9034);
and U10330 (N_10330,N_9543,N_9276);
nand U10331 (N_10331,N_8926,N_9202);
nand U10332 (N_10332,N_9524,N_9845);
xnor U10333 (N_10333,N_9262,N_9104);
and U10334 (N_10334,N_9253,N_9327);
nand U10335 (N_10335,N_8792,N_9599);
or U10336 (N_10336,N_9055,N_9415);
and U10337 (N_10337,N_9774,N_9141);
nand U10338 (N_10338,N_9721,N_9791);
nor U10339 (N_10339,N_9632,N_9158);
xor U10340 (N_10340,N_9188,N_9923);
xor U10341 (N_10341,N_9715,N_9915);
and U10342 (N_10342,N_9605,N_9683);
and U10343 (N_10343,N_9416,N_9724);
xor U10344 (N_10344,N_8995,N_9108);
and U10345 (N_10345,N_9625,N_9073);
nor U10346 (N_10346,N_9854,N_9374);
or U10347 (N_10347,N_9123,N_9545);
xnor U10348 (N_10348,N_9135,N_9992);
nand U10349 (N_10349,N_9811,N_9277);
xnor U10350 (N_10350,N_9096,N_8966);
and U10351 (N_10351,N_9170,N_9695);
or U10352 (N_10352,N_9372,N_9755);
and U10353 (N_10353,N_9954,N_8824);
nor U10354 (N_10354,N_9072,N_9516);
xnor U10355 (N_10355,N_9815,N_8890);
nor U10356 (N_10356,N_9749,N_9365);
nand U10357 (N_10357,N_9150,N_9892);
or U10358 (N_10358,N_8998,N_8875);
xor U10359 (N_10359,N_9190,N_8786);
nor U10360 (N_10360,N_9079,N_9922);
nand U10361 (N_10361,N_9346,N_9382);
or U10362 (N_10362,N_9982,N_9345);
or U10363 (N_10363,N_9920,N_9186);
and U10364 (N_10364,N_9101,N_9437);
and U10365 (N_10365,N_9566,N_9486);
and U10366 (N_10366,N_9164,N_9089);
and U10367 (N_10367,N_9384,N_9897);
nor U10368 (N_10368,N_9797,N_9236);
nand U10369 (N_10369,N_9246,N_9351);
nor U10370 (N_10370,N_8886,N_8781);
xor U10371 (N_10371,N_9793,N_8964);
nand U10372 (N_10372,N_8785,N_9401);
or U10373 (N_10373,N_9853,N_9025);
or U10374 (N_10374,N_9834,N_9799);
and U10375 (N_10375,N_9016,N_9023);
or U10376 (N_10376,N_9621,N_9657);
nand U10377 (N_10377,N_9060,N_9676);
or U10378 (N_10378,N_9708,N_9425);
or U10379 (N_10379,N_9159,N_8985);
nand U10380 (N_10380,N_8778,N_9735);
and U10381 (N_10381,N_9929,N_9696);
nor U10382 (N_10382,N_9918,N_9038);
nor U10383 (N_10383,N_9976,N_8941);
or U10384 (N_10384,N_9558,N_9426);
and U10385 (N_10385,N_9279,N_8805);
nand U10386 (N_10386,N_9778,N_9571);
nand U10387 (N_10387,N_9380,N_9287);
nor U10388 (N_10388,N_9641,N_9707);
and U10389 (N_10389,N_9000,N_9194);
and U10390 (N_10390,N_9238,N_9574);
and U10391 (N_10391,N_9421,N_9875);
and U10392 (N_10392,N_9366,N_9942);
nor U10393 (N_10393,N_9488,N_9943);
and U10394 (N_10394,N_9722,N_9450);
or U10395 (N_10395,N_9044,N_9267);
and U10396 (N_10396,N_8804,N_9984);
or U10397 (N_10397,N_9143,N_9634);
nand U10398 (N_10398,N_8909,N_8751);
xor U10399 (N_10399,N_9746,N_9909);
nand U10400 (N_10400,N_9652,N_8947);
nand U10401 (N_10401,N_9491,N_9881);
or U10402 (N_10402,N_9665,N_9010);
xnor U10403 (N_10403,N_9668,N_9386);
or U10404 (N_10404,N_9642,N_9028);
nand U10405 (N_10405,N_9926,N_9271);
or U10406 (N_10406,N_9120,N_8885);
nand U10407 (N_10407,N_9563,N_9515);
nand U10408 (N_10408,N_8801,N_9056);
nand U10409 (N_10409,N_8776,N_9906);
xor U10410 (N_10410,N_9004,N_9692);
or U10411 (N_10411,N_9932,N_9816);
nor U10412 (N_10412,N_9223,N_9356);
or U10413 (N_10413,N_9991,N_9841);
xor U10414 (N_10414,N_9274,N_8940);
xor U10415 (N_10415,N_8851,N_9639);
nand U10416 (N_10416,N_9678,N_9648);
or U10417 (N_10417,N_8798,N_8906);
xor U10418 (N_10418,N_9838,N_9970);
and U10419 (N_10419,N_8918,N_8795);
xnor U10420 (N_10420,N_8844,N_9505);
nand U10421 (N_10421,N_8916,N_9701);
xnor U10422 (N_10422,N_8806,N_9308);
and U10423 (N_10423,N_9361,N_9947);
nor U10424 (N_10424,N_8809,N_9861);
and U10425 (N_10425,N_9728,N_8783);
and U10426 (N_10426,N_9654,N_8829);
nor U10427 (N_10427,N_9465,N_9456);
xor U10428 (N_10428,N_9314,N_8828);
nor U10429 (N_10429,N_9184,N_9731);
nor U10430 (N_10430,N_8914,N_9467);
nor U10431 (N_10431,N_9043,N_9200);
nand U10432 (N_10432,N_8866,N_9596);
nor U10433 (N_10433,N_9539,N_9517);
and U10434 (N_10434,N_9661,N_9638);
nand U10435 (N_10435,N_9127,N_9844);
xnor U10436 (N_10436,N_9859,N_9183);
nor U10437 (N_10437,N_8987,N_9368);
and U10438 (N_10438,N_9114,N_8891);
or U10439 (N_10439,N_9492,N_9428);
or U10440 (N_10440,N_9682,N_9530);
xor U10441 (N_10441,N_9699,N_9272);
nor U10442 (N_10442,N_9228,N_9496);
xor U10443 (N_10443,N_9763,N_9785);
or U10444 (N_10444,N_9857,N_8821);
or U10445 (N_10445,N_9544,N_9349);
nand U10446 (N_10446,N_8991,N_9085);
or U10447 (N_10447,N_9012,N_9576);
nor U10448 (N_10448,N_9031,N_8763);
or U10449 (N_10449,N_9432,N_9786);
nand U10450 (N_10450,N_9994,N_9209);
or U10451 (N_10451,N_9671,N_9552);
nor U10452 (N_10452,N_9848,N_9477);
or U10453 (N_10453,N_8807,N_8836);
or U10454 (N_10454,N_8762,N_8973);
and U10455 (N_10455,N_9482,N_8812);
nor U10456 (N_10456,N_9385,N_9520);
and U10457 (N_10457,N_9667,N_9877);
nand U10458 (N_10458,N_9956,N_9435);
xnor U10459 (N_10459,N_9087,N_9940);
or U10460 (N_10460,N_8942,N_9140);
or U10461 (N_10461,N_9939,N_9282);
nand U10462 (N_10462,N_8952,N_9637);
nor U10463 (N_10463,N_8963,N_9320);
nor U10464 (N_10464,N_9161,N_9930);
xor U10465 (N_10465,N_9030,N_9359);
or U10466 (N_10466,N_8951,N_9575);
nand U10467 (N_10467,N_9397,N_9762);
nor U10468 (N_10468,N_8927,N_9534);
xnor U10469 (N_10469,N_9203,N_9630);
nand U10470 (N_10470,N_9014,N_9390);
nor U10471 (N_10471,N_9018,N_9789);
or U10472 (N_10472,N_8810,N_8816);
and U10473 (N_10473,N_8982,N_8978);
and U10474 (N_10474,N_9494,N_9008);
nor U10475 (N_10475,N_9580,N_9449);
xnor U10476 (N_10476,N_9042,N_9180);
or U10477 (N_10477,N_9291,N_9620);
nor U10478 (N_10478,N_9118,N_9608);
or U10479 (N_10479,N_9091,N_9646);
nand U10480 (N_10480,N_9742,N_9842);
nor U10481 (N_10481,N_9635,N_9360);
or U10482 (N_10482,N_9328,N_9411);
or U10483 (N_10483,N_9809,N_8935);
nand U10484 (N_10484,N_8884,N_9703);
nor U10485 (N_10485,N_9406,N_9852);
xnor U10486 (N_10486,N_9760,N_9147);
and U10487 (N_10487,N_9124,N_9936);
nor U10488 (N_10488,N_9139,N_9548);
xnor U10489 (N_10489,N_8788,N_9739);
xnor U10490 (N_10490,N_9207,N_9111);
xnor U10491 (N_10491,N_9723,N_9064);
nand U10492 (N_10492,N_9285,N_9870);
xnor U10493 (N_10493,N_9154,N_9080);
nor U10494 (N_10494,N_8750,N_9610);
xnor U10495 (N_10495,N_9978,N_9817);
nor U10496 (N_10496,N_9381,N_9894);
nand U10497 (N_10497,N_9985,N_8867);
and U10498 (N_10498,N_9902,N_9989);
and U10499 (N_10499,N_8910,N_8949);
and U10500 (N_10500,N_9950,N_9337);
nand U10501 (N_10501,N_9295,N_8925);
and U10502 (N_10502,N_9798,N_9364);
xor U10503 (N_10503,N_8780,N_9388);
or U10504 (N_10504,N_9054,N_9996);
and U10505 (N_10505,N_9136,N_9355);
nor U10506 (N_10506,N_9955,N_9889);
nor U10507 (N_10507,N_9751,N_8874);
or U10508 (N_10508,N_9137,N_9824);
nand U10509 (N_10509,N_9037,N_8880);
and U10510 (N_10510,N_9737,N_9318);
nor U10511 (N_10511,N_9828,N_9609);
nand U10512 (N_10512,N_9675,N_9142);
and U10513 (N_10513,N_9444,N_8856);
or U10514 (N_10514,N_9212,N_9335);
or U10515 (N_10515,N_9182,N_9745);
xor U10516 (N_10516,N_8979,N_9316);
nand U10517 (N_10517,N_9322,N_9704);
nor U10518 (N_10518,N_9890,N_9493);
nand U10519 (N_10519,N_9899,N_9658);
xor U10520 (N_10520,N_9476,N_9418);
nand U10521 (N_10521,N_9176,N_9115);
and U10522 (N_10522,N_9266,N_9471);
nand U10523 (N_10523,N_9502,N_9500);
nand U10524 (N_10524,N_9048,N_9995);
nor U10525 (N_10525,N_9756,N_8822);
or U10526 (N_10526,N_9377,N_9457);
and U10527 (N_10527,N_9604,N_9602);
nor U10528 (N_10528,N_9480,N_9470);
xnor U10529 (N_10529,N_9106,N_8840);
or U10530 (N_10530,N_9097,N_8794);
nor U10531 (N_10531,N_9475,N_9474);
nor U10532 (N_10532,N_8853,N_9352);
or U10533 (N_10533,N_8971,N_9100);
and U10534 (N_10534,N_9711,N_9820);
xnor U10535 (N_10535,N_9826,N_9197);
xnor U10536 (N_10536,N_9395,N_8888);
nand U10537 (N_10537,N_9714,N_8950);
and U10538 (N_10538,N_9168,N_9329);
nand U10539 (N_10539,N_9958,N_9321);
xnor U10540 (N_10540,N_9807,N_8961);
xor U10541 (N_10541,N_8837,N_9830);
and U10542 (N_10542,N_9133,N_9099);
xor U10543 (N_10543,N_9458,N_9410);
nor U10544 (N_10544,N_9151,N_9219);
xor U10545 (N_10545,N_9245,N_9214);
and U10546 (N_10546,N_9473,N_8939);
and U10547 (N_10547,N_8938,N_9766);
or U10548 (N_10548,N_9964,N_9103);
nand U10549 (N_10549,N_9057,N_9583);
nand U10550 (N_10550,N_9873,N_9993);
and U10551 (N_10551,N_9006,N_9033);
xor U10552 (N_10552,N_8965,N_9969);
nor U10553 (N_10553,N_9736,N_8999);
xnor U10554 (N_10554,N_9810,N_8774);
nand U10555 (N_10555,N_9542,N_8879);
nor U10556 (N_10556,N_8773,N_8928);
nand U10557 (N_10557,N_8755,N_8958);
xnor U10558 (N_10558,N_9759,N_9836);
or U10559 (N_10559,N_9931,N_9862);
nand U10560 (N_10560,N_9082,N_9593);
nor U10561 (N_10561,N_9027,N_9317);
nor U10562 (N_10562,N_9305,N_9773);
xnor U10563 (N_10563,N_8946,N_9251);
xnor U10564 (N_10564,N_9499,N_9081);
and U10565 (N_10565,N_9441,N_9643);
or U10566 (N_10566,N_9666,N_9040);
nand U10567 (N_10567,N_9556,N_9805);
nor U10568 (N_10568,N_9670,N_8993);
or U10569 (N_10569,N_9117,N_9389);
and U10570 (N_10570,N_9430,N_8960);
and U10571 (N_10571,N_9907,N_9694);
or U10572 (N_10572,N_9350,N_8753);
xnor U10573 (N_10573,N_9404,N_9325);
nand U10574 (N_10574,N_9568,N_9581);
xor U10575 (N_10575,N_9503,N_8894);
and U10576 (N_10576,N_8882,N_8862);
xor U10577 (N_10577,N_9371,N_9527);
nor U10578 (N_10578,N_8779,N_9917);
nand U10579 (N_10579,N_8782,N_9067);
nand U10580 (N_10580,N_8796,N_9567);
nor U10581 (N_10581,N_9537,N_9076);
and U10582 (N_10582,N_9132,N_9433);
and U10583 (N_10583,N_9270,N_9716);
nand U10584 (N_10584,N_9636,N_9005);
xnor U10585 (N_10585,N_9422,N_9439);
nand U10586 (N_10586,N_9584,N_9226);
nor U10587 (N_10587,N_9679,N_9174);
nand U10588 (N_10588,N_9874,N_9882);
and U10589 (N_10589,N_9047,N_9434);
xor U10590 (N_10590,N_9990,N_9152);
and U10591 (N_10591,N_8959,N_8757);
nand U10592 (N_10592,N_9925,N_9338);
xnor U10593 (N_10593,N_9764,N_9284);
nor U10594 (N_10594,N_9163,N_9846);
nand U10595 (N_10595,N_9804,N_9049);
or U10596 (N_10596,N_9252,N_9265);
nor U10597 (N_10597,N_9452,N_9533);
and U10598 (N_10598,N_9059,N_8962);
nand U10599 (N_10599,N_9886,N_9611);
nor U10600 (N_10600,N_9065,N_9257);
or U10601 (N_10601,N_8827,N_9855);
xnor U10602 (N_10602,N_8825,N_8929);
or U10603 (N_10603,N_8944,N_8854);
or U10604 (N_10604,N_9447,N_9967);
nand U10605 (N_10605,N_9885,N_9526);
nor U10606 (N_10606,N_9927,N_9032);
nand U10607 (N_10607,N_9250,N_9916);
nand U10608 (N_10608,N_8842,N_8931);
nor U10609 (N_10609,N_8756,N_9189);
nor U10610 (N_10610,N_9512,N_9769);
nand U10611 (N_10611,N_9233,N_8975);
or U10612 (N_10612,N_9479,N_9191);
nand U10613 (N_10613,N_9600,N_9092);
nand U10614 (N_10614,N_9258,N_8849);
nand U10615 (N_10615,N_9821,N_9326);
nand U10616 (N_10616,N_9340,N_9938);
and U10617 (N_10617,N_9840,N_9689);
and U10618 (N_10618,N_8863,N_8896);
xor U10619 (N_10619,N_9697,N_9782);
or U10620 (N_10620,N_9904,N_9832);
or U10621 (N_10621,N_8887,N_8953);
and U10622 (N_10622,N_9684,N_9960);
and U10623 (N_10623,N_9869,N_9565);
or U10624 (N_10624,N_9011,N_9664);
or U10625 (N_10625,N_9892,N_9492);
or U10626 (N_10626,N_9605,N_9696);
xor U10627 (N_10627,N_9500,N_9588);
xor U10628 (N_10628,N_9775,N_8974);
xor U10629 (N_10629,N_9873,N_9000);
nand U10630 (N_10630,N_9662,N_9989);
nand U10631 (N_10631,N_9635,N_9792);
xor U10632 (N_10632,N_9074,N_9387);
and U10633 (N_10633,N_9275,N_9214);
or U10634 (N_10634,N_9799,N_9440);
nand U10635 (N_10635,N_9413,N_9929);
nor U10636 (N_10636,N_9175,N_9727);
nor U10637 (N_10637,N_9928,N_9562);
nor U10638 (N_10638,N_9962,N_8794);
or U10639 (N_10639,N_9123,N_9919);
xnor U10640 (N_10640,N_9905,N_9912);
nand U10641 (N_10641,N_9818,N_9457);
and U10642 (N_10642,N_9756,N_9740);
nand U10643 (N_10643,N_9938,N_9554);
xor U10644 (N_10644,N_9506,N_9576);
nand U10645 (N_10645,N_9279,N_9658);
or U10646 (N_10646,N_9062,N_8765);
and U10647 (N_10647,N_9841,N_9780);
and U10648 (N_10648,N_9154,N_9001);
nor U10649 (N_10649,N_8975,N_9556);
nor U10650 (N_10650,N_9713,N_8786);
and U10651 (N_10651,N_9892,N_9110);
xnor U10652 (N_10652,N_9752,N_9514);
nor U10653 (N_10653,N_9885,N_9747);
and U10654 (N_10654,N_9007,N_9923);
and U10655 (N_10655,N_9725,N_9944);
nand U10656 (N_10656,N_9859,N_9596);
and U10657 (N_10657,N_9236,N_9456);
nor U10658 (N_10658,N_9446,N_9068);
and U10659 (N_10659,N_9236,N_9677);
nor U10660 (N_10660,N_8840,N_8802);
nor U10661 (N_10661,N_9625,N_9051);
xnor U10662 (N_10662,N_9242,N_9532);
nand U10663 (N_10663,N_9385,N_9991);
xnor U10664 (N_10664,N_9603,N_9806);
and U10665 (N_10665,N_8767,N_9216);
or U10666 (N_10666,N_9945,N_9977);
nor U10667 (N_10667,N_9632,N_9622);
or U10668 (N_10668,N_9531,N_9341);
nor U10669 (N_10669,N_8797,N_9145);
or U10670 (N_10670,N_9885,N_9558);
and U10671 (N_10671,N_9720,N_8929);
nor U10672 (N_10672,N_9433,N_8832);
xor U10673 (N_10673,N_9260,N_8986);
and U10674 (N_10674,N_9082,N_9181);
and U10675 (N_10675,N_9080,N_8934);
nand U10676 (N_10676,N_9743,N_9201);
xor U10677 (N_10677,N_9514,N_8928);
xnor U10678 (N_10678,N_9253,N_9966);
or U10679 (N_10679,N_9260,N_9749);
and U10680 (N_10680,N_9975,N_9144);
nor U10681 (N_10681,N_9307,N_9049);
nor U10682 (N_10682,N_8886,N_9003);
and U10683 (N_10683,N_9428,N_9067);
nand U10684 (N_10684,N_9295,N_8903);
or U10685 (N_10685,N_9474,N_8967);
or U10686 (N_10686,N_9574,N_9298);
and U10687 (N_10687,N_9736,N_9537);
nor U10688 (N_10688,N_9138,N_9788);
or U10689 (N_10689,N_9498,N_9681);
xnor U10690 (N_10690,N_8788,N_9904);
xor U10691 (N_10691,N_9730,N_9871);
xor U10692 (N_10692,N_9621,N_8812);
or U10693 (N_10693,N_9562,N_9946);
nand U10694 (N_10694,N_9258,N_9183);
nor U10695 (N_10695,N_9877,N_8833);
nand U10696 (N_10696,N_9110,N_8929);
or U10697 (N_10697,N_9596,N_8995);
nand U10698 (N_10698,N_9806,N_9376);
xnor U10699 (N_10699,N_9823,N_9867);
nand U10700 (N_10700,N_9913,N_9416);
xnor U10701 (N_10701,N_9654,N_9101);
nor U10702 (N_10702,N_9939,N_9975);
nor U10703 (N_10703,N_9495,N_9524);
nor U10704 (N_10704,N_9110,N_9009);
nor U10705 (N_10705,N_8910,N_9314);
nor U10706 (N_10706,N_9564,N_9525);
xor U10707 (N_10707,N_9189,N_8945);
or U10708 (N_10708,N_9448,N_9799);
nand U10709 (N_10709,N_9582,N_8927);
and U10710 (N_10710,N_8779,N_8934);
and U10711 (N_10711,N_8914,N_9760);
nand U10712 (N_10712,N_8920,N_8764);
or U10713 (N_10713,N_9698,N_8935);
nor U10714 (N_10714,N_9649,N_8890);
nor U10715 (N_10715,N_8811,N_9789);
nand U10716 (N_10716,N_9033,N_9485);
xnor U10717 (N_10717,N_8898,N_9615);
nand U10718 (N_10718,N_8940,N_9906);
or U10719 (N_10719,N_9636,N_9944);
and U10720 (N_10720,N_9899,N_9368);
and U10721 (N_10721,N_9003,N_9469);
or U10722 (N_10722,N_8832,N_9312);
and U10723 (N_10723,N_9538,N_8851);
and U10724 (N_10724,N_9611,N_9790);
xor U10725 (N_10725,N_9192,N_9695);
and U10726 (N_10726,N_9001,N_8929);
or U10727 (N_10727,N_9019,N_9128);
nand U10728 (N_10728,N_9516,N_9778);
nand U10729 (N_10729,N_9803,N_9004);
or U10730 (N_10730,N_9678,N_9223);
xor U10731 (N_10731,N_9673,N_9111);
nor U10732 (N_10732,N_8831,N_8951);
nor U10733 (N_10733,N_9765,N_9882);
or U10734 (N_10734,N_9340,N_9949);
xnor U10735 (N_10735,N_8958,N_8897);
and U10736 (N_10736,N_9829,N_8824);
xnor U10737 (N_10737,N_9975,N_9305);
or U10738 (N_10738,N_9560,N_8948);
and U10739 (N_10739,N_8910,N_9033);
nand U10740 (N_10740,N_9515,N_9550);
nor U10741 (N_10741,N_9090,N_9758);
or U10742 (N_10742,N_9349,N_9404);
or U10743 (N_10743,N_8914,N_9841);
nand U10744 (N_10744,N_8928,N_9230);
nand U10745 (N_10745,N_9349,N_9461);
nand U10746 (N_10746,N_9512,N_8928);
and U10747 (N_10747,N_9854,N_9685);
or U10748 (N_10748,N_9487,N_9212);
nor U10749 (N_10749,N_9134,N_9214);
xor U10750 (N_10750,N_9692,N_9212);
and U10751 (N_10751,N_9124,N_9040);
nand U10752 (N_10752,N_9966,N_8760);
or U10753 (N_10753,N_9756,N_9520);
and U10754 (N_10754,N_9188,N_9575);
nor U10755 (N_10755,N_9294,N_9302);
xnor U10756 (N_10756,N_9094,N_9003);
nand U10757 (N_10757,N_9123,N_9036);
nand U10758 (N_10758,N_9955,N_9572);
xnor U10759 (N_10759,N_9572,N_8862);
and U10760 (N_10760,N_9855,N_9044);
nor U10761 (N_10761,N_8860,N_8896);
and U10762 (N_10762,N_9478,N_9880);
xor U10763 (N_10763,N_9480,N_8831);
and U10764 (N_10764,N_9511,N_8877);
nand U10765 (N_10765,N_9382,N_8975);
or U10766 (N_10766,N_9777,N_9334);
xnor U10767 (N_10767,N_9118,N_9974);
xor U10768 (N_10768,N_9880,N_8884);
nand U10769 (N_10769,N_9058,N_9025);
and U10770 (N_10770,N_9625,N_9337);
nand U10771 (N_10771,N_9453,N_9726);
or U10772 (N_10772,N_9410,N_9397);
or U10773 (N_10773,N_9583,N_8812);
xnor U10774 (N_10774,N_8947,N_9607);
nor U10775 (N_10775,N_9027,N_9953);
or U10776 (N_10776,N_9950,N_9315);
xor U10777 (N_10777,N_8911,N_9256);
nor U10778 (N_10778,N_9521,N_9303);
nor U10779 (N_10779,N_9973,N_9126);
nand U10780 (N_10780,N_8759,N_9425);
and U10781 (N_10781,N_9666,N_9031);
xor U10782 (N_10782,N_9867,N_8754);
nand U10783 (N_10783,N_9326,N_9770);
xor U10784 (N_10784,N_9129,N_8769);
xnor U10785 (N_10785,N_8868,N_9905);
nand U10786 (N_10786,N_9056,N_9642);
or U10787 (N_10787,N_8795,N_9542);
xnor U10788 (N_10788,N_9761,N_8874);
nor U10789 (N_10789,N_9730,N_9239);
or U10790 (N_10790,N_9347,N_9045);
or U10791 (N_10791,N_9712,N_9122);
xnor U10792 (N_10792,N_9298,N_9008);
nor U10793 (N_10793,N_9425,N_9687);
or U10794 (N_10794,N_9036,N_9612);
or U10795 (N_10795,N_9571,N_9453);
nor U10796 (N_10796,N_9604,N_9460);
nand U10797 (N_10797,N_9265,N_9395);
nand U10798 (N_10798,N_9845,N_9046);
or U10799 (N_10799,N_8792,N_9952);
xnor U10800 (N_10800,N_9357,N_9754);
nor U10801 (N_10801,N_9497,N_9689);
nor U10802 (N_10802,N_9182,N_8947);
nor U10803 (N_10803,N_9491,N_9383);
and U10804 (N_10804,N_8800,N_8915);
and U10805 (N_10805,N_9978,N_9296);
xor U10806 (N_10806,N_9597,N_9460);
and U10807 (N_10807,N_9389,N_9753);
and U10808 (N_10808,N_9559,N_9915);
or U10809 (N_10809,N_9911,N_9377);
and U10810 (N_10810,N_9321,N_9649);
nand U10811 (N_10811,N_9472,N_9228);
nand U10812 (N_10812,N_9480,N_9486);
and U10813 (N_10813,N_9970,N_9878);
or U10814 (N_10814,N_9276,N_9609);
nand U10815 (N_10815,N_9497,N_9182);
nor U10816 (N_10816,N_9695,N_9620);
and U10817 (N_10817,N_9091,N_9469);
nand U10818 (N_10818,N_9666,N_8861);
nand U10819 (N_10819,N_9597,N_9108);
nand U10820 (N_10820,N_8886,N_9419);
and U10821 (N_10821,N_9476,N_9681);
and U10822 (N_10822,N_9108,N_8791);
nor U10823 (N_10823,N_9634,N_9757);
or U10824 (N_10824,N_9059,N_9555);
xor U10825 (N_10825,N_9226,N_9883);
and U10826 (N_10826,N_8928,N_9305);
and U10827 (N_10827,N_9165,N_9980);
or U10828 (N_10828,N_9255,N_8960);
nand U10829 (N_10829,N_8960,N_8801);
xnor U10830 (N_10830,N_9782,N_9456);
nor U10831 (N_10831,N_9177,N_9452);
or U10832 (N_10832,N_9687,N_9169);
and U10833 (N_10833,N_9260,N_9019);
nor U10834 (N_10834,N_9345,N_9715);
and U10835 (N_10835,N_9592,N_9676);
nand U10836 (N_10836,N_9832,N_9787);
and U10837 (N_10837,N_9840,N_9605);
or U10838 (N_10838,N_9757,N_8773);
and U10839 (N_10839,N_9302,N_9523);
and U10840 (N_10840,N_9669,N_8868);
nor U10841 (N_10841,N_9958,N_8887);
nand U10842 (N_10842,N_8826,N_9895);
nor U10843 (N_10843,N_8928,N_8987);
nor U10844 (N_10844,N_9780,N_9616);
or U10845 (N_10845,N_9114,N_9417);
nor U10846 (N_10846,N_9124,N_8898);
nand U10847 (N_10847,N_9463,N_8754);
and U10848 (N_10848,N_9652,N_9029);
nor U10849 (N_10849,N_8860,N_9072);
or U10850 (N_10850,N_9063,N_8973);
nor U10851 (N_10851,N_8889,N_9924);
nor U10852 (N_10852,N_9742,N_9610);
xor U10853 (N_10853,N_9698,N_9662);
nor U10854 (N_10854,N_9401,N_9281);
and U10855 (N_10855,N_9433,N_8927);
nand U10856 (N_10856,N_9158,N_9621);
xor U10857 (N_10857,N_9667,N_9743);
nor U10858 (N_10858,N_8819,N_8928);
and U10859 (N_10859,N_9989,N_8927);
xnor U10860 (N_10860,N_9879,N_9545);
and U10861 (N_10861,N_9745,N_9228);
and U10862 (N_10862,N_9792,N_9827);
or U10863 (N_10863,N_9199,N_9829);
or U10864 (N_10864,N_9152,N_9963);
or U10865 (N_10865,N_9713,N_9168);
or U10866 (N_10866,N_9221,N_9501);
xor U10867 (N_10867,N_9855,N_9367);
nor U10868 (N_10868,N_8852,N_9993);
xnor U10869 (N_10869,N_9796,N_8829);
and U10870 (N_10870,N_9647,N_8791);
or U10871 (N_10871,N_9745,N_9918);
nor U10872 (N_10872,N_8872,N_9844);
and U10873 (N_10873,N_9748,N_9535);
nor U10874 (N_10874,N_9594,N_8775);
or U10875 (N_10875,N_9680,N_8792);
or U10876 (N_10876,N_9399,N_8817);
and U10877 (N_10877,N_9479,N_9162);
nand U10878 (N_10878,N_9726,N_9552);
nor U10879 (N_10879,N_9181,N_9751);
nand U10880 (N_10880,N_9089,N_8957);
nor U10881 (N_10881,N_9447,N_9925);
xnor U10882 (N_10882,N_8961,N_9331);
and U10883 (N_10883,N_9596,N_8825);
nand U10884 (N_10884,N_9363,N_9125);
or U10885 (N_10885,N_9292,N_8945);
nor U10886 (N_10886,N_9554,N_9232);
or U10887 (N_10887,N_9586,N_9693);
or U10888 (N_10888,N_9445,N_9110);
nor U10889 (N_10889,N_9611,N_9432);
and U10890 (N_10890,N_9880,N_9457);
xor U10891 (N_10891,N_8904,N_8888);
and U10892 (N_10892,N_8845,N_8915);
nand U10893 (N_10893,N_9865,N_9333);
nand U10894 (N_10894,N_9772,N_9689);
or U10895 (N_10895,N_8994,N_9666);
or U10896 (N_10896,N_9912,N_9871);
and U10897 (N_10897,N_9341,N_9098);
nand U10898 (N_10898,N_9557,N_9118);
or U10899 (N_10899,N_9926,N_9879);
nand U10900 (N_10900,N_9593,N_8783);
or U10901 (N_10901,N_9068,N_9320);
nand U10902 (N_10902,N_9145,N_9899);
or U10903 (N_10903,N_9232,N_9435);
and U10904 (N_10904,N_8811,N_9350);
xor U10905 (N_10905,N_9029,N_8947);
xnor U10906 (N_10906,N_9812,N_9295);
nor U10907 (N_10907,N_8934,N_9211);
or U10908 (N_10908,N_9569,N_9422);
nor U10909 (N_10909,N_9731,N_9102);
and U10910 (N_10910,N_9747,N_9924);
xor U10911 (N_10911,N_9860,N_9171);
or U10912 (N_10912,N_9161,N_9222);
nor U10913 (N_10913,N_9382,N_8963);
xnor U10914 (N_10914,N_8933,N_9637);
xor U10915 (N_10915,N_9514,N_8760);
xnor U10916 (N_10916,N_9532,N_8927);
or U10917 (N_10917,N_8914,N_9850);
nand U10918 (N_10918,N_9700,N_8947);
xor U10919 (N_10919,N_9168,N_9553);
and U10920 (N_10920,N_8980,N_9395);
and U10921 (N_10921,N_9332,N_9354);
nor U10922 (N_10922,N_9352,N_9474);
xor U10923 (N_10923,N_9699,N_9960);
or U10924 (N_10924,N_9023,N_8839);
or U10925 (N_10925,N_9521,N_9366);
and U10926 (N_10926,N_8891,N_9190);
or U10927 (N_10927,N_9804,N_8884);
and U10928 (N_10928,N_9171,N_9755);
nor U10929 (N_10929,N_9233,N_9499);
or U10930 (N_10930,N_9485,N_8929);
nor U10931 (N_10931,N_9903,N_9731);
nor U10932 (N_10932,N_9912,N_9194);
nand U10933 (N_10933,N_9966,N_9150);
and U10934 (N_10934,N_9836,N_9655);
nand U10935 (N_10935,N_9251,N_9576);
nor U10936 (N_10936,N_9309,N_9367);
nor U10937 (N_10937,N_9717,N_9958);
xnor U10938 (N_10938,N_9312,N_9911);
and U10939 (N_10939,N_9347,N_9980);
nor U10940 (N_10940,N_8989,N_9464);
or U10941 (N_10941,N_9826,N_9836);
or U10942 (N_10942,N_9256,N_8859);
nor U10943 (N_10943,N_9401,N_8939);
nor U10944 (N_10944,N_9976,N_9863);
nor U10945 (N_10945,N_9951,N_9197);
nand U10946 (N_10946,N_9276,N_8857);
and U10947 (N_10947,N_9958,N_9829);
nor U10948 (N_10948,N_9307,N_8796);
nor U10949 (N_10949,N_9531,N_9009);
nand U10950 (N_10950,N_8939,N_9158);
nand U10951 (N_10951,N_9867,N_9932);
xnor U10952 (N_10952,N_9961,N_9983);
xnor U10953 (N_10953,N_9997,N_9100);
nand U10954 (N_10954,N_9831,N_9724);
and U10955 (N_10955,N_8796,N_9462);
nor U10956 (N_10956,N_9612,N_8788);
nor U10957 (N_10957,N_9626,N_9282);
or U10958 (N_10958,N_9998,N_9679);
and U10959 (N_10959,N_9561,N_9769);
xor U10960 (N_10960,N_8873,N_8840);
xnor U10961 (N_10961,N_9326,N_9679);
xnor U10962 (N_10962,N_9316,N_8851);
or U10963 (N_10963,N_8770,N_9797);
or U10964 (N_10964,N_9160,N_9101);
nand U10965 (N_10965,N_9182,N_9107);
xor U10966 (N_10966,N_8849,N_9451);
xor U10967 (N_10967,N_9452,N_9671);
and U10968 (N_10968,N_9955,N_8767);
or U10969 (N_10969,N_9437,N_9691);
nand U10970 (N_10970,N_9471,N_9097);
xor U10971 (N_10971,N_9264,N_9000);
and U10972 (N_10972,N_9415,N_9848);
and U10973 (N_10973,N_8837,N_8772);
nor U10974 (N_10974,N_9366,N_9468);
or U10975 (N_10975,N_9844,N_8965);
nand U10976 (N_10976,N_8787,N_9454);
or U10977 (N_10977,N_9000,N_9433);
nand U10978 (N_10978,N_9307,N_8996);
xnor U10979 (N_10979,N_9636,N_9537);
or U10980 (N_10980,N_9252,N_9269);
xnor U10981 (N_10981,N_8761,N_9815);
xor U10982 (N_10982,N_9412,N_9154);
xnor U10983 (N_10983,N_9551,N_9865);
xnor U10984 (N_10984,N_9749,N_9201);
and U10985 (N_10985,N_8994,N_9784);
nand U10986 (N_10986,N_9357,N_9682);
xor U10987 (N_10987,N_8815,N_8973);
or U10988 (N_10988,N_9471,N_9053);
nor U10989 (N_10989,N_9540,N_9504);
nor U10990 (N_10990,N_9996,N_9882);
nand U10991 (N_10991,N_8812,N_8938);
and U10992 (N_10992,N_8917,N_8830);
nand U10993 (N_10993,N_9209,N_9764);
nor U10994 (N_10994,N_9058,N_9055);
and U10995 (N_10995,N_9952,N_9583);
nor U10996 (N_10996,N_9939,N_9076);
xnor U10997 (N_10997,N_8873,N_9640);
nor U10998 (N_10998,N_9205,N_8932);
nor U10999 (N_10999,N_8898,N_9787);
nand U11000 (N_11000,N_9365,N_8998);
or U11001 (N_11001,N_9976,N_9754);
nand U11002 (N_11002,N_9471,N_8926);
nand U11003 (N_11003,N_9923,N_9612);
nand U11004 (N_11004,N_9009,N_9462);
or U11005 (N_11005,N_9954,N_8862);
nand U11006 (N_11006,N_9013,N_9838);
nand U11007 (N_11007,N_9341,N_8972);
and U11008 (N_11008,N_9655,N_9515);
or U11009 (N_11009,N_9647,N_9519);
nor U11010 (N_11010,N_9868,N_9864);
nor U11011 (N_11011,N_9599,N_9150);
xnor U11012 (N_11012,N_9472,N_9079);
nor U11013 (N_11013,N_9896,N_9614);
and U11014 (N_11014,N_9732,N_9226);
nand U11015 (N_11015,N_9833,N_9377);
xor U11016 (N_11016,N_9719,N_9861);
xnor U11017 (N_11017,N_9648,N_9936);
nand U11018 (N_11018,N_8978,N_9503);
xor U11019 (N_11019,N_8816,N_9723);
xnor U11020 (N_11020,N_8768,N_9928);
xnor U11021 (N_11021,N_9685,N_9993);
and U11022 (N_11022,N_9377,N_9017);
or U11023 (N_11023,N_8826,N_9408);
and U11024 (N_11024,N_8772,N_9307);
and U11025 (N_11025,N_9858,N_9671);
xor U11026 (N_11026,N_9191,N_9599);
nor U11027 (N_11027,N_8826,N_8975);
nand U11028 (N_11028,N_8763,N_9739);
or U11029 (N_11029,N_9144,N_8994);
or U11030 (N_11030,N_9669,N_8869);
or U11031 (N_11031,N_9142,N_9638);
nand U11032 (N_11032,N_9002,N_9454);
xnor U11033 (N_11033,N_8930,N_9656);
nor U11034 (N_11034,N_9583,N_8834);
xnor U11035 (N_11035,N_9002,N_9821);
xnor U11036 (N_11036,N_9466,N_9298);
nor U11037 (N_11037,N_9704,N_9438);
xor U11038 (N_11038,N_9799,N_8762);
nand U11039 (N_11039,N_9947,N_8846);
and U11040 (N_11040,N_9735,N_9831);
and U11041 (N_11041,N_9469,N_9676);
xor U11042 (N_11042,N_9692,N_9155);
and U11043 (N_11043,N_9500,N_9442);
or U11044 (N_11044,N_9954,N_9276);
xor U11045 (N_11045,N_9933,N_8987);
or U11046 (N_11046,N_9583,N_9219);
xnor U11047 (N_11047,N_9852,N_9252);
nor U11048 (N_11048,N_9013,N_9339);
nand U11049 (N_11049,N_9953,N_9607);
and U11050 (N_11050,N_9689,N_9147);
or U11051 (N_11051,N_9602,N_9479);
and U11052 (N_11052,N_9138,N_9602);
and U11053 (N_11053,N_9376,N_9121);
or U11054 (N_11054,N_9463,N_9487);
or U11055 (N_11055,N_9743,N_9405);
nand U11056 (N_11056,N_9013,N_9446);
xnor U11057 (N_11057,N_9115,N_9134);
nor U11058 (N_11058,N_9343,N_9842);
and U11059 (N_11059,N_9557,N_9069);
nand U11060 (N_11060,N_9617,N_9409);
nor U11061 (N_11061,N_8933,N_9567);
nand U11062 (N_11062,N_8761,N_9114);
and U11063 (N_11063,N_8954,N_9153);
nand U11064 (N_11064,N_8858,N_9397);
nor U11065 (N_11065,N_8937,N_9568);
and U11066 (N_11066,N_9410,N_8918);
and U11067 (N_11067,N_9255,N_9129);
and U11068 (N_11068,N_9469,N_9381);
xnor U11069 (N_11069,N_9659,N_9915);
and U11070 (N_11070,N_9273,N_9833);
or U11071 (N_11071,N_8984,N_8827);
nor U11072 (N_11072,N_9946,N_9871);
or U11073 (N_11073,N_9616,N_8896);
nor U11074 (N_11074,N_9696,N_9947);
nand U11075 (N_11075,N_9300,N_9432);
or U11076 (N_11076,N_9818,N_9841);
nor U11077 (N_11077,N_9824,N_8949);
nand U11078 (N_11078,N_8784,N_9687);
nor U11079 (N_11079,N_9746,N_9268);
or U11080 (N_11080,N_9591,N_8915);
and U11081 (N_11081,N_9524,N_9807);
xor U11082 (N_11082,N_9705,N_9084);
and U11083 (N_11083,N_9091,N_9598);
xor U11084 (N_11084,N_9496,N_9254);
xor U11085 (N_11085,N_8892,N_9733);
nand U11086 (N_11086,N_9469,N_9198);
and U11087 (N_11087,N_9629,N_8976);
and U11088 (N_11088,N_9151,N_8783);
xnor U11089 (N_11089,N_9089,N_9962);
xor U11090 (N_11090,N_8778,N_9972);
nor U11091 (N_11091,N_8762,N_9917);
and U11092 (N_11092,N_9349,N_9443);
xor U11093 (N_11093,N_9360,N_9512);
xor U11094 (N_11094,N_9036,N_8828);
or U11095 (N_11095,N_9739,N_9194);
and U11096 (N_11096,N_9983,N_8993);
xor U11097 (N_11097,N_8997,N_9416);
or U11098 (N_11098,N_9690,N_9158);
or U11099 (N_11099,N_9785,N_8813);
and U11100 (N_11100,N_9975,N_9815);
nand U11101 (N_11101,N_9307,N_9645);
nor U11102 (N_11102,N_9507,N_9025);
nand U11103 (N_11103,N_9568,N_9807);
or U11104 (N_11104,N_8776,N_8931);
nor U11105 (N_11105,N_9667,N_8909);
nor U11106 (N_11106,N_9321,N_9970);
nor U11107 (N_11107,N_9767,N_9390);
xnor U11108 (N_11108,N_9899,N_8836);
and U11109 (N_11109,N_9110,N_9691);
nand U11110 (N_11110,N_9829,N_8785);
and U11111 (N_11111,N_9544,N_9394);
xor U11112 (N_11112,N_9968,N_8980);
nand U11113 (N_11113,N_8935,N_8768);
or U11114 (N_11114,N_9375,N_9807);
or U11115 (N_11115,N_9042,N_8758);
and U11116 (N_11116,N_9265,N_9027);
nand U11117 (N_11117,N_9457,N_9503);
or U11118 (N_11118,N_8913,N_9885);
xnor U11119 (N_11119,N_9431,N_8931);
or U11120 (N_11120,N_9792,N_9057);
xnor U11121 (N_11121,N_8856,N_9841);
xor U11122 (N_11122,N_9272,N_9026);
nand U11123 (N_11123,N_8811,N_9587);
nor U11124 (N_11124,N_8885,N_9499);
nand U11125 (N_11125,N_9553,N_9285);
nor U11126 (N_11126,N_9365,N_9166);
nand U11127 (N_11127,N_9570,N_9944);
nor U11128 (N_11128,N_9845,N_9037);
and U11129 (N_11129,N_9239,N_9524);
xor U11130 (N_11130,N_9491,N_9747);
nor U11131 (N_11131,N_9853,N_9069);
xnor U11132 (N_11132,N_8785,N_9980);
or U11133 (N_11133,N_8813,N_9276);
and U11134 (N_11134,N_9076,N_9683);
and U11135 (N_11135,N_9827,N_9030);
xor U11136 (N_11136,N_9816,N_9956);
or U11137 (N_11137,N_8837,N_9061);
nor U11138 (N_11138,N_9442,N_8997);
and U11139 (N_11139,N_9174,N_9227);
and U11140 (N_11140,N_9639,N_8819);
nor U11141 (N_11141,N_9627,N_9408);
nor U11142 (N_11142,N_9714,N_9922);
nor U11143 (N_11143,N_9248,N_9899);
nand U11144 (N_11144,N_9478,N_9875);
nor U11145 (N_11145,N_9558,N_9006);
nand U11146 (N_11146,N_9009,N_9589);
and U11147 (N_11147,N_8875,N_8938);
and U11148 (N_11148,N_8964,N_9832);
nor U11149 (N_11149,N_9229,N_9232);
and U11150 (N_11150,N_9025,N_8754);
xnor U11151 (N_11151,N_9677,N_9061);
or U11152 (N_11152,N_9895,N_9293);
nor U11153 (N_11153,N_9992,N_9852);
xnor U11154 (N_11154,N_8998,N_9626);
or U11155 (N_11155,N_9109,N_9749);
nand U11156 (N_11156,N_9358,N_8970);
and U11157 (N_11157,N_9731,N_9290);
xor U11158 (N_11158,N_9062,N_9681);
nand U11159 (N_11159,N_9555,N_9424);
xnor U11160 (N_11160,N_9446,N_8855);
and U11161 (N_11161,N_9590,N_9515);
xnor U11162 (N_11162,N_9489,N_9658);
nand U11163 (N_11163,N_9551,N_9653);
nand U11164 (N_11164,N_8753,N_9589);
xnor U11165 (N_11165,N_9392,N_9187);
or U11166 (N_11166,N_9529,N_8873);
xnor U11167 (N_11167,N_9765,N_9912);
and U11168 (N_11168,N_9335,N_9038);
and U11169 (N_11169,N_9720,N_8863);
nor U11170 (N_11170,N_9642,N_9477);
or U11171 (N_11171,N_8848,N_9525);
and U11172 (N_11172,N_9703,N_9209);
xnor U11173 (N_11173,N_9951,N_9918);
or U11174 (N_11174,N_9282,N_9180);
and U11175 (N_11175,N_8976,N_9475);
nand U11176 (N_11176,N_9144,N_8782);
nor U11177 (N_11177,N_9734,N_9979);
nor U11178 (N_11178,N_9986,N_9275);
nand U11179 (N_11179,N_9153,N_9204);
or U11180 (N_11180,N_9925,N_9978);
or U11181 (N_11181,N_9903,N_8817);
and U11182 (N_11182,N_9744,N_9618);
nor U11183 (N_11183,N_9162,N_9887);
nor U11184 (N_11184,N_9902,N_8889);
xnor U11185 (N_11185,N_9602,N_9776);
xnor U11186 (N_11186,N_9471,N_8917);
nor U11187 (N_11187,N_9010,N_9221);
nor U11188 (N_11188,N_9315,N_9167);
and U11189 (N_11189,N_8877,N_9742);
xor U11190 (N_11190,N_9101,N_8989);
and U11191 (N_11191,N_9408,N_9270);
and U11192 (N_11192,N_9864,N_9824);
xnor U11193 (N_11193,N_9590,N_9014);
nand U11194 (N_11194,N_9521,N_8896);
and U11195 (N_11195,N_9666,N_9555);
nor U11196 (N_11196,N_9158,N_9047);
and U11197 (N_11197,N_9431,N_8997);
nor U11198 (N_11198,N_9981,N_9610);
xor U11199 (N_11199,N_9354,N_9152);
nand U11200 (N_11200,N_8926,N_9585);
nor U11201 (N_11201,N_9982,N_9277);
nor U11202 (N_11202,N_9235,N_9254);
xnor U11203 (N_11203,N_8896,N_9140);
nand U11204 (N_11204,N_9173,N_9965);
or U11205 (N_11205,N_9333,N_9762);
nand U11206 (N_11206,N_9405,N_9626);
and U11207 (N_11207,N_9019,N_9848);
nand U11208 (N_11208,N_8938,N_8929);
xnor U11209 (N_11209,N_9322,N_9117);
xnor U11210 (N_11210,N_9998,N_9788);
or U11211 (N_11211,N_9758,N_9670);
xor U11212 (N_11212,N_9172,N_9252);
nor U11213 (N_11213,N_9182,N_9671);
nor U11214 (N_11214,N_8966,N_9224);
nor U11215 (N_11215,N_9499,N_9822);
nand U11216 (N_11216,N_9919,N_9336);
xor U11217 (N_11217,N_9243,N_9215);
xor U11218 (N_11218,N_9474,N_9671);
or U11219 (N_11219,N_9065,N_9763);
nand U11220 (N_11220,N_9041,N_9572);
or U11221 (N_11221,N_8939,N_9862);
xor U11222 (N_11222,N_9444,N_9752);
xor U11223 (N_11223,N_9331,N_9821);
nor U11224 (N_11224,N_9281,N_9584);
nor U11225 (N_11225,N_9701,N_9606);
xnor U11226 (N_11226,N_8866,N_9228);
nand U11227 (N_11227,N_9961,N_9575);
or U11228 (N_11228,N_8800,N_9080);
xnor U11229 (N_11229,N_9824,N_8932);
or U11230 (N_11230,N_9244,N_9982);
and U11231 (N_11231,N_9399,N_9625);
or U11232 (N_11232,N_9956,N_9585);
nor U11233 (N_11233,N_9901,N_8867);
and U11234 (N_11234,N_9714,N_9463);
nand U11235 (N_11235,N_8889,N_9940);
nor U11236 (N_11236,N_8799,N_9021);
xnor U11237 (N_11237,N_8797,N_9478);
nor U11238 (N_11238,N_9274,N_9233);
and U11239 (N_11239,N_9060,N_9704);
nor U11240 (N_11240,N_9647,N_8929);
or U11241 (N_11241,N_9546,N_8775);
xnor U11242 (N_11242,N_8800,N_9515);
and U11243 (N_11243,N_9610,N_8992);
nand U11244 (N_11244,N_8751,N_8821);
nand U11245 (N_11245,N_8940,N_8857);
xnor U11246 (N_11246,N_9660,N_9618);
nand U11247 (N_11247,N_9089,N_9442);
and U11248 (N_11248,N_9859,N_9419);
or U11249 (N_11249,N_9681,N_8967);
and U11250 (N_11250,N_10188,N_10273);
nor U11251 (N_11251,N_10750,N_10746);
or U11252 (N_11252,N_10890,N_10315);
xor U11253 (N_11253,N_11071,N_10596);
nor U11254 (N_11254,N_10942,N_10901);
or U11255 (N_11255,N_11126,N_10154);
nor U11256 (N_11256,N_10199,N_10679);
nand U11257 (N_11257,N_10909,N_11150);
and U11258 (N_11258,N_10986,N_10364);
nand U11259 (N_11259,N_10248,N_10133);
or U11260 (N_11260,N_11127,N_10407);
or U11261 (N_11261,N_10039,N_11209);
nor U11262 (N_11262,N_10976,N_10705);
or U11263 (N_11263,N_11037,N_11055);
and U11264 (N_11264,N_10853,N_10802);
and U11265 (N_11265,N_10606,N_10061);
and U11266 (N_11266,N_10506,N_10049);
or U11267 (N_11267,N_10623,N_10322);
nand U11268 (N_11268,N_11121,N_10771);
nor U11269 (N_11269,N_11082,N_11035);
nand U11270 (N_11270,N_10877,N_10466);
xor U11271 (N_11271,N_10914,N_11145);
nor U11272 (N_11272,N_11222,N_10891);
xnor U11273 (N_11273,N_10689,N_10230);
and U11274 (N_11274,N_10932,N_10965);
xor U11275 (N_11275,N_10301,N_10622);
and U11276 (N_11276,N_10369,N_10565);
nor U11277 (N_11277,N_10189,N_10363);
and U11278 (N_11278,N_10751,N_10699);
or U11279 (N_11279,N_11208,N_10920);
xor U11280 (N_11280,N_10055,N_11128);
nor U11281 (N_11281,N_11031,N_10380);
and U11282 (N_11282,N_10324,N_10483);
nand U11283 (N_11283,N_11134,N_10422);
or U11284 (N_11284,N_10963,N_10334);
nor U11285 (N_11285,N_10654,N_10603);
or U11286 (N_11286,N_11234,N_10716);
xnor U11287 (N_11287,N_11003,N_10392);
xnor U11288 (N_11288,N_10217,N_10532);
and U11289 (N_11289,N_10872,N_10616);
nor U11290 (N_11290,N_10544,N_10703);
and U11291 (N_11291,N_10528,N_10101);
nand U11292 (N_11292,N_11096,N_11067);
or U11293 (N_11293,N_10631,N_10686);
xnor U11294 (N_11294,N_10576,N_10670);
xor U11295 (N_11295,N_10168,N_10029);
nand U11296 (N_11296,N_10768,N_11163);
nand U11297 (N_11297,N_10080,N_11075);
nor U11298 (N_11298,N_10685,N_10903);
or U11299 (N_11299,N_11142,N_10999);
and U11300 (N_11300,N_10897,N_10349);
nand U11301 (N_11301,N_10774,N_10103);
xor U11302 (N_11302,N_11132,N_10052);
or U11303 (N_11303,N_10373,N_10389);
nand U11304 (N_11304,N_10298,N_10737);
nand U11305 (N_11305,N_10045,N_10968);
nor U11306 (N_11306,N_10702,N_10321);
nand U11307 (N_11307,N_10573,N_10054);
nand U11308 (N_11308,N_10355,N_10869);
nand U11309 (N_11309,N_10658,N_10320);
nand U11310 (N_11310,N_10284,N_10379);
nand U11311 (N_11311,N_10038,N_10644);
or U11312 (N_11312,N_10536,N_10557);
and U11313 (N_11313,N_10667,N_10659);
nor U11314 (N_11314,N_11043,N_10031);
xnor U11315 (N_11315,N_10804,N_10717);
and U11316 (N_11316,N_10517,N_10312);
nand U11317 (N_11317,N_10933,N_10894);
and U11318 (N_11318,N_10310,N_10226);
xor U11319 (N_11319,N_11232,N_10181);
or U11320 (N_11320,N_10857,N_10791);
or U11321 (N_11321,N_10205,N_10251);
and U11322 (N_11322,N_11215,N_10594);
or U11323 (N_11323,N_10478,N_10192);
or U11324 (N_11324,N_10850,N_10957);
xor U11325 (N_11325,N_10775,N_10640);
nor U11326 (N_11326,N_10022,N_10912);
nand U11327 (N_11327,N_10091,N_11245);
or U11328 (N_11328,N_10607,N_10534);
nor U11329 (N_11329,N_10479,N_10260);
and U11330 (N_11330,N_10327,N_10161);
and U11331 (N_11331,N_11090,N_10065);
nand U11332 (N_11332,N_10155,N_10148);
nor U11333 (N_11333,N_11220,N_10524);
nand U11334 (N_11334,N_10359,N_10263);
or U11335 (N_11335,N_11064,N_11131);
xor U11336 (N_11336,N_11085,N_10278);
xor U11337 (N_11337,N_10639,N_11130);
nor U11338 (N_11338,N_10948,N_10035);
nand U11339 (N_11339,N_10243,N_10100);
nor U11340 (N_11340,N_10811,N_11025);
nor U11341 (N_11341,N_10842,N_10209);
nor U11342 (N_11342,N_10680,N_10428);
nor U11343 (N_11343,N_10739,N_10477);
or U11344 (N_11344,N_10258,N_11139);
nand U11345 (N_11345,N_10977,N_10391);
or U11346 (N_11346,N_10156,N_11249);
nand U11347 (N_11347,N_10120,N_11087);
and U11348 (N_11348,N_10564,N_10413);
nand U11349 (N_11349,N_10552,N_10515);
or U11350 (N_11350,N_10780,N_11048);
xnor U11351 (N_11351,N_10417,N_10086);
xor U11352 (N_11352,N_10332,N_10036);
nor U11353 (N_11353,N_10326,N_11189);
nor U11354 (N_11354,N_10374,N_11013);
and U11355 (N_11355,N_10475,N_10458);
xnor U11356 (N_11356,N_11103,N_10822);
and U11357 (N_11357,N_10924,N_10265);
nand U11358 (N_11358,N_11113,N_10510);
xnor U11359 (N_11359,N_10164,N_10106);
nor U11360 (N_11360,N_10668,N_11122);
nand U11361 (N_11361,N_10406,N_10462);
nand U11362 (N_11362,N_10190,N_10024);
nor U11363 (N_11363,N_10939,N_11235);
or U11364 (N_11364,N_10151,N_10443);
nand U11365 (N_11365,N_10711,N_10394);
nand U11366 (N_11366,N_10318,N_10064);
or U11367 (N_11367,N_11164,N_10809);
xor U11368 (N_11368,N_10601,N_10964);
and U11369 (N_11369,N_10004,N_10755);
nor U11370 (N_11370,N_10170,N_10366);
or U11371 (N_11371,N_11198,N_11180);
or U11372 (N_11372,N_10643,N_10937);
xnor U11373 (N_11373,N_10328,N_10222);
or U11374 (N_11374,N_10261,N_10114);
or U11375 (N_11375,N_10608,N_10858);
and U11376 (N_11376,N_10316,N_11138);
or U11377 (N_11377,N_10843,N_11050);
nor U11378 (N_11378,N_10076,N_10271);
nand U11379 (N_11379,N_11176,N_10602);
xor U11380 (N_11380,N_11211,N_11203);
nand U11381 (N_11381,N_10183,N_11034);
and U11382 (N_11382,N_10415,N_10730);
nor U11383 (N_11383,N_10219,N_10420);
nand U11384 (N_11384,N_10488,N_10581);
and U11385 (N_11385,N_10706,N_11162);
nand U11386 (N_11386,N_11206,N_10704);
or U11387 (N_11387,N_11144,N_10377);
or U11388 (N_11388,N_10911,N_10272);
and U11389 (N_11389,N_11086,N_10405);
nor U11390 (N_11390,N_10001,N_10830);
xnor U11391 (N_11391,N_11223,N_10424);
nand U11392 (N_11392,N_10208,N_10105);
xor U11393 (N_11393,N_10047,N_11136);
nand U11394 (N_11394,N_10958,N_10323);
nor U11395 (N_11395,N_10828,N_10354);
nor U11396 (N_11396,N_10815,N_10214);
or U11397 (N_11397,N_10126,N_10915);
xnor U11398 (N_11398,N_10060,N_10421);
xnor U11399 (N_11399,N_10425,N_10027);
nand U11400 (N_11400,N_11100,N_10441);
nor U11401 (N_11401,N_11158,N_11177);
and U11402 (N_11402,N_10728,N_11033);
xnor U11403 (N_11403,N_10966,N_10401);
and U11404 (N_11404,N_10378,N_10063);
nand U11405 (N_11405,N_10591,N_10457);
and U11406 (N_11406,N_10609,N_10729);
and U11407 (N_11407,N_10922,N_10333);
xor U11408 (N_11408,N_10671,N_10940);
nand U11409 (N_11409,N_10145,N_10788);
or U11410 (N_11410,N_10473,N_10783);
nor U11411 (N_11411,N_10393,N_10617);
nor U11412 (N_11412,N_10725,N_10396);
or U11413 (N_11413,N_10898,N_10980);
xor U11414 (N_11414,N_10635,N_10227);
or U11415 (N_11415,N_10246,N_10368);
or U11416 (N_11416,N_10496,N_10078);
xor U11417 (N_11417,N_10158,N_10094);
nor U11418 (N_11418,N_10043,N_10285);
xnor U11419 (N_11419,N_10874,N_10033);
and U11420 (N_11420,N_10371,N_10875);
nor U11421 (N_11421,N_10956,N_10876);
and U11422 (N_11422,N_10625,N_10143);
xor U11423 (N_11423,N_10849,N_11179);
nand U11424 (N_11424,N_10416,N_10302);
nand U11425 (N_11425,N_10878,N_10212);
or U11426 (N_11426,N_10715,N_10283);
and U11427 (N_11427,N_10134,N_10893);
nand U11428 (N_11428,N_10152,N_10972);
xnor U11429 (N_11429,N_10795,N_10238);
or U11430 (N_11430,N_10137,N_10837);
and U11431 (N_11431,N_10159,N_10993);
or U11432 (N_11432,N_10691,N_10513);
nor U11433 (N_11433,N_10628,N_10916);
or U11434 (N_11434,N_10068,N_10817);
and U11435 (N_11435,N_10868,N_10649);
and U11436 (N_11436,N_10587,N_11205);
and U11437 (N_11437,N_11023,N_11063);
xnor U11438 (N_11438,N_10382,N_11153);
or U11439 (N_11439,N_10203,N_10969);
or U11440 (N_11440,N_10995,N_11151);
or U11441 (N_11441,N_10376,N_10116);
xor U11442 (N_11442,N_11195,N_10867);
and U11443 (N_11443,N_10259,N_10262);
and U11444 (N_11444,N_10860,N_10089);
xnor U11445 (N_11445,N_10037,N_10147);
xnor U11446 (N_11446,N_11092,N_10132);
and U11447 (N_11447,N_10292,N_11202);
xor U11448 (N_11448,N_10941,N_10294);
nor U11449 (N_11449,N_10588,N_10032);
nand U11450 (N_11450,N_10432,N_11041);
and U11451 (N_11451,N_11143,N_10459);
nand U11452 (N_11452,N_10232,N_11088);
xnor U11453 (N_11453,N_10618,N_11006);
nand U11454 (N_11454,N_11230,N_10008);
nand U11455 (N_11455,N_10386,N_10339);
nor U11456 (N_11456,N_10082,N_10651);
nor U11457 (N_11457,N_10551,N_10991);
or U11458 (N_11458,N_10287,N_10648);
or U11459 (N_11459,N_10097,N_11160);
nor U11460 (N_11460,N_11196,N_11019);
xnor U11461 (N_11461,N_10288,N_10745);
nor U11462 (N_11462,N_10357,N_10303);
nor U11463 (N_11463,N_10166,N_10344);
and U11464 (N_11464,N_10683,N_10983);
nand U11465 (N_11465,N_10777,N_10854);
or U11466 (N_11466,N_10088,N_10529);
or U11467 (N_11467,N_10928,N_10257);
xnor U11468 (N_11468,N_10081,N_10062);
and U11469 (N_11469,N_11212,N_10182);
xor U11470 (N_11470,N_10930,N_10020);
nand U11471 (N_11471,N_11197,N_11089);
nand U11472 (N_11472,N_10215,N_10598);
nor U11473 (N_11473,N_11173,N_10550);
nor U11474 (N_11474,N_11133,N_10347);
or U11475 (N_11475,N_10994,N_10856);
nor U11476 (N_11476,N_10201,N_10652);
xor U11477 (N_11477,N_10638,N_10487);
or U11478 (N_11478,N_10010,N_10213);
nand U11479 (N_11479,N_11093,N_10484);
nand U11480 (N_11480,N_10676,N_10330);
and U11481 (N_11481,N_10423,N_10266);
nor U11482 (N_11482,N_10176,N_10071);
nand U11483 (N_11483,N_10697,N_10722);
and U11484 (N_11484,N_10887,N_10677);
nor U11485 (N_11485,N_11032,N_10153);
and U11486 (N_11486,N_10592,N_10814);
nand U11487 (N_11487,N_10992,N_10256);
nor U11488 (N_11488,N_10646,N_10350);
nand U11489 (N_11489,N_10838,N_10130);
and U11490 (N_11490,N_10974,N_10673);
nor U11491 (N_11491,N_10577,N_10526);
xnor U11492 (N_11492,N_10495,N_11115);
xor U11493 (N_11493,N_10489,N_11084);
and U11494 (N_11494,N_10899,N_10277);
or U11495 (N_11495,N_10763,N_10543);
nor U11496 (N_11496,N_11247,N_11001);
or U11497 (N_11497,N_10435,N_10178);
nand U11498 (N_11498,N_11059,N_10904);
nand U11499 (N_11499,N_11175,N_10463);
xnor U11500 (N_11500,N_10926,N_10426);
and U11501 (N_11501,N_10929,N_10007);
nand U11502 (N_11502,N_10018,N_10776);
nor U11503 (N_11503,N_10034,N_10343);
and U11504 (N_11504,N_11028,N_10952);
or U11505 (N_11505,N_10331,N_10707);
nand U11506 (N_11506,N_10485,N_10005);
and U11507 (N_11507,N_10753,N_10452);
nand U11508 (N_11508,N_10864,N_10681);
nand U11509 (N_11509,N_10090,N_10525);
nand U11510 (N_11510,N_10637,N_11024);
or U11511 (N_11511,N_11125,N_10665);
and U11512 (N_11512,N_10388,N_11178);
nand U11513 (N_11513,N_11194,N_10743);
and U11514 (N_11514,N_11004,N_10851);
nand U11515 (N_11515,N_10351,N_10537);
xor U11516 (N_11516,N_10279,N_10880);
nand U11517 (N_11517,N_10235,N_10925);
xnor U11518 (N_11518,N_10797,N_10656);
and U11519 (N_11519,N_10218,N_10056);
nand U11520 (N_11520,N_11040,N_10579);
or U11521 (N_11521,N_10862,N_11120);
and U11522 (N_11522,N_11233,N_10000);
xnor U11523 (N_11523,N_10863,N_11123);
xnor U11524 (N_11524,N_11237,N_11057);
or U11525 (N_11525,N_10778,N_10943);
and U11526 (N_11526,N_11052,N_11191);
and U11527 (N_11527,N_10437,N_10270);
nor U11528 (N_11528,N_11056,N_11137);
xnor U11529 (N_11529,N_10372,N_10570);
xnor U11530 (N_11530,N_10770,N_10852);
nand U11531 (N_11531,N_10571,N_10087);
nand U11532 (N_11532,N_10945,N_10693);
and U11533 (N_11533,N_11111,N_10954);
or U11534 (N_11534,N_10306,N_10732);
or U11535 (N_11535,N_10229,N_10070);
nor U11536 (N_11536,N_10023,N_10834);
nor U11537 (N_11537,N_10286,N_10522);
xnor U11538 (N_11538,N_10560,N_10695);
xnor U11539 (N_11539,N_10626,N_11114);
xor U11540 (N_11540,N_10512,N_10411);
nand U11541 (N_11541,N_10113,N_10855);
nor U11542 (N_11542,N_10497,N_10742);
nor U11543 (N_11543,N_11074,N_10664);
or U11544 (N_11544,N_10934,N_10160);
xnor U11545 (N_11545,N_11072,N_10779);
nand U11546 (N_11546,N_10481,N_11022);
nand U11547 (N_11547,N_10641,N_10311);
or U11548 (N_11548,N_11045,N_10122);
or U11549 (N_11549,N_10150,N_11070);
or U11550 (N_11550,N_11039,N_10655);
or U11551 (N_11551,N_10720,N_10900);
and U11552 (N_11552,N_10430,N_10498);
nand U11553 (N_11553,N_10998,N_10268);
or U11554 (N_11554,N_10600,N_10482);
or U11555 (N_11555,N_10210,N_10866);
nand U11556 (N_11556,N_10455,N_10634);
nor U11557 (N_11557,N_10092,N_11192);
xnor U11558 (N_11558,N_10519,N_10765);
and U11559 (N_11559,N_10696,N_10469);
and U11560 (N_11560,N_11054,N_10249);
xor U11561 (N_11561,N_10491,N_10494);
and U11562 (N_11562,N_10206,N_10612);
and U11563 (N_11563,N_10599,N_10580);
or U11564 (N_11564,N_11161,N_11030);
nand U11565 (N_11565,N_10724,N_10767);
or U11566 (N_11566,N_10040,N_11185);
xor U11567 (N_11567,N_10048,N_11224);
and U11568 (N_11568,N_10936,N_11012);
or U11569 (N_11569,N_10960,N_10666);
nor U11570 (N_11570,N_10395,N_10012);
nor U11571 (N_11571,N_10053,N_10541);
or U11572 (N_11572,N_10220,N_10823);
or U11573 (N_11573,N_10399,N_10381);
nand U11574 (N_11574,N_11236,N_11219);
xor U11575 (N_11575,N_10545,N_10169);
nor U11576 (N_11576,N_10955,N_10935);
xor U11577 (N_11577,N_10104,N_10449);
or U11578 (N_11578,N_10058,N_10030);
nand U11579 (N_11579,N_10810,N_10718);
xnor U11580 (N_11580,N_10953,N_11098);
xor U11581 (N_11581,N_10650,N_10236);
nand U11582 (N_11582,N_10848,N_10398);
nor U11583 (N_11583,N_10614,N_10508);
and U11584 (N_11584,N_10884,N_11017);
and U11585 (N_11585,N_10454,N_10444);
xor U11586 (N_11586,N_10172,N_11105);
nor U11587 (N_11587,N_10535,N_10889);
nor U11588 (N_11588,N_11021,N_10264);
nand U11589 (N_11589,N_10296,N_10710);
and U11590 (N_11590,N_10193,N_10511);
xor U11591 (N_11591,N_11106,N_10721);
and U11592 (N_11592,N_10784,N_10723);
or U11593 (N_11593,N_10672,N_11200);
or U11594 (N_11594,N_10412,N_10761);
xnor U11595 (N_11595,N_11020,N_10503);
and U11596 (N_11596,N_10507,N_10846);
and U11597 (N_11597,N_10562,N_10735);
nand U11598 (N_11598,N_10630,N_10548);
and U11599 (N_11599,N_11170,N_10317);
nand U11600 (N_11600,N_10233,N_11049);
and U11601 (N_11601,N_11009,N_11081);
or U11602 (N_11602,N_10984,N_10516);
and U11603 (N_11603,N_10520,N_10385);
nor U11604 (N_11604,N_11073,N_10253);
xnor U11605 (N_11605,N_10892,N_10613);
xor U11606 (N_11606,N_10445,N_10139);
and U11607 (N_11607,N_10549,N_10769);
or U11608 (N_11608,N_11169,N_10881);
nand U11609 (N_11609,N_10016,N_10051);
xnor U11610 (N_11610,N_10124,N_10300);
nor U11611 (N_11611,N_10727,N_11207);
nor U11612 (N_11612,N_10907,N_10174);
and U11613 (N_11613,N_11204,N_10514);
nor U11614 (N_11614,N_10223,N_10207);
xor U11615 (N_11615,N_10927,N_10346);
nor U11616 (N_11616,N_10772,N_10173);
nand U11617 (N_11617,N_10733,N_11181);
or U11618 (N_11618,N_10748,N_11068);
and U11619 (N_11619,N_10709,N_10404);
or U11620 (N_11620,N_10824,N_10414);
xor U11621 (N_11621,N_10067,N_10619);
and U11622 (N_11622,N_10293,N_10821);
nor U11623 (N_11623,N_10847,N_10237);
nand U11624 (N_11624,N_11110,N_10669);
and U11625 (N_11625,N_10859,N_10660);
or U11626 (N_11626,N_10611,N_11201);
and U11627 (N_11627,N_10074,N_10959);
nor U11628 (N_11628,N_11218,N_10231);
or U11629 (N_11629,N_10585,N_10179);
or U11630 (N_11630,N_10419,N_11117);
nor U11631 (N_11631,N_10017,N_10370);
and U11632 (N_11632,N_11129,N_10627);
xor U11633 (N_11633,N_11026,N_10605);
or U11634 (N_11634,N_11091,N_10636);
and U11635 (N_11635,N_11231,N_10621);
xnor U11636 (N_11636,N_11053,N_10938);
xnor U11637 (N_11637,N_10502,N_10861);
and U11638 (N_11638,N_10002,N_10692);
xnor U11639 (N_11639,N_10431,N_10115);
nor U11640 (N_11640,N_10028,N_10165);
nand U11641 (N_11641,N_11188,N_10624);
and U11642 (N_11642,N_10274,N_10708);
nor U11643 (N_11643,N_10865,N_10766);
nor U11644 (N_11644,N_10131,N_10314);
and U11645 (N_11645,N_10228,N_10329);
and U11646 (N_11646,N_10073,N_10845);
and U11647 (N_11647,N_10267,N_10194);
nand U11648 (N_11648,N_11156,N_10338);
nand U11649 (N_11649,N_11058,N_10099);
or U11650 (N_11650,N_10125,N_11016);
nand U11651 (N_11651,N_10888,N_10360);
xor U11652 (N_11652,N_10832,N_10798);
or U11653 (N_11653,N_10572,N_10353);
nor U11654 (N_11654,N_10447,N_10690);
xor U11655 (N_11655,N_10807,N_10275);
xor U11656 (N_11656,N_10474,N_11246);
nand U11657 (N_11657,N_10096,N_10409);
nand U11658 (N_11658,N_11042,N_10792);
xnor U11659 (N_11659,N_11069,N_10990);
nor U11660 (N_11660,N_10402,N_10460);
and U11661 (N_11661,N_10786,N_10662);
or U11662 (N_11662,N_10185,N_10533);
xnor U11663 (N_11663,N_10812,N_11243);
nand U11664 (N_11664,N_10918,N_10175);
and U11665 (N_11665,N_10509,N_10873);
or U11666 (N_11666,N_10006,N_11182);
nand U11667 (N_11667,N_10295,N_10245);
or U11668 (N_11668,N_11228,N_10818);
or U11669 (N_11669,N_10593,N_10714);
xor U11670 (N_11670,N_10141,N_11104);
or U11671 (N_11671,N_10400,N_10794);
or U11672 (N_11672,N_10712,N_10870);
nand U11673 (N_11673,N_10793,N_10997);
nand U11674 (N_11674,N_10642,N_11141);
or U11675 (N_11675,N_10200,N_10578);
nand U11676 (N_11676,N_10895,N_10467);
nand U11677 (N_11677,N_11029,N_10504);
and U11678 (N_11678,N_10661,N_10647);
and U11679 (N_11679,N_11061,N_11119);
and U11680 (N_11680,N_10569,N_10011);
and U11681 (N_11681,N_10352,N_10967);
and U11682 (N_11682,N_10072,N_10111);
or U11683 (N_11683,N_10254,N_11008);
and U11684 (N_11684,N_10657,N_10518);
xnor U11685 (N_11685,N_10586,N_10531);
and U11686 (N_11686,N_10461,N_10367);
xor U11687 (N_11687,N_10142,N_10910);
or U11688 (N_11688,N_11108,N_10726);
nor U11689 (N_11689,N_10325,N_10384);
nor U11690 (N_11690,N_10108,N_10184);
and U11691 (N_11691,N_11095,N_10003);
and U11692 (N_11692,N_10335,N_10615);
xor U11693 (N_11693,N_11097,N_10451);
and U11694 (N_11694,N_10568,N_10931);
nand U11695 (N_11695,N_10135,N_10800);
or U11696 (N_11696,N_10480,N_10244);
xnor U11697 (N_11697,N_10281,N_10553);
nand U11698 (N_11698,N_10902,N_10299);
nand U11699 (N_11699,N_10629,N_10799);
nand U11700 (N_11700,N_10046,N_10575);
nand U11701 (N_11701,N_10829,N_10136);
and U11702 (N_11702,N_10744,N_10981);
and U11703 (N_11703,N_10140,N_10803);
nand U11704 (N_11704,N_10687,N_11165);
or U11705 (N_11705,N_10996,N_10436);
xnor U11706 (N_11706,N_10840,N_10289);
nand U11707 (N_11707,N_10442,N_10951);
or U11708 (N_11708,N_10700,N_10042);
nand U11709 (N_11709,N_10950,N_10906);
xor U11710 (N_11710,N_10234,N_10202);
or U11711 (N_11711,N_11107,N_10149);
and U11712 (N_11712,N_10291,N_10163);
nand U11713 (N_11713,N_10808,N_11174);
nand U11714 (N_11714,N_10782,N_10678);
nor U11715 (N_11715,N_10741,N_10883);
nand U11716 (N_11716,N_11225,N_10758);
nand U11717 (N_11717,N_10556,N_10762);
nor U11718 (N_11718,N_10561,N_10408);
nor U11719 (N_11719,N_10736,N_10345);
nor U11720 (N_11720,N_10438,N_11241);
nand U11721 (N_11721,N_10186,N_11005);
or U11722 (N_11722,N_11217,N_10198);
nor U11723 (N_11723,N_10841,N_11186);
nand U11724 (N_11724,N_10180,N_10110);
nor U11725 (N_11725,N_11094,N_11083);
nor U11726 (N_11726,N_11227,N_11010);
and U11727 (N_11727,N_10781,N_10574);
nor U11728 (N_11728,N_10340,N_10610);
and U11729 (N_11729,N_10107,N_11240);
xor U11730 (N_11730,N_10913,N_10747);
or U11731 (N_11731,N_11065,N_10719);
nand U11732 (N_11732,N_10567,N_10684);
nand U11733 (N_11733,N_10144,N_10216);
or U11734 (N_11734,N_10985,N_11118);
nor U11735 (N_11735,N_10348,N_10632);
nand U11736 (N_11736,N_10688,N_10313);
and U11737 (N_11737,N_10127,N_10871);
nand U11738 (N_11738,N_11147,N_10464);
nand U11739 (N_11739,N_11216,N_10946);
nand U11740 (N_11740,N_10731,N_11027);
nand U11741 (N_11741,N_10013,N_10434);
or U11742 (N_11742,N_10453,N_10589);
nor U11743 (N_11743,N_10701,N_10456);
xnor U11744 (N_11744,N_10390,N_11000);
nor U11745 (N_11745,N_10439,N_11066);
nor U11746 (N_11746,N_10410,N_10342);
nand U11747 (N_11747,N_10558,N_11155);
and U11748 (N_11748,N_11051,N_10752);
xnor U11749 (N_11749,N_11183,N_11015);
or U11750 (N_11750,N_10337,N_10831);
and U11751 (N_11751,N_10276,N_10805);
and U11752 (N_11752,N_10117,N_10336);
nand U11753 (N_11753,N_10204,N_10129);
xor U11754 (N_11754,N_10523,N_10645);
xor U11755 (N_11755,N_10975,N_10083);
and U11756 (N_11756,N_10358,N_10988);
or U11757 (N_11757,N_10468,N_10050);
nor U11758 (N_11758,N_11244,N_10309);
and U11759 (N_11759,N_10123,N_11148);
or U11760 (N_11760,N_10225,N_10446);
nand U11761 (N_11761,N_11011,N_10566);
nor U11762 (N_11762,N_10280,N_11229);
xnor U11763 (N_11763,N_11214,N_10987);
and U11764 (N_11764,N_10713,N_10026);
and U11765 (N_11765,N_11112,N_10121);
nand U11766 (N_11766,N_11199,N_10500);
and U11767 (N_11767,N_10789,N_10538);
or U11768 (N_11768,N_11002,N_10240);
and U11769 (N_11769,N_10694,N_10282);
xnor U11770 (N_11770,N_11152,N_10604);
nand U11771 (N_11771,N_10825,N_11099);
or U11772 (N_11772,N_11018,N_10021);
xnor U11773 (N_11773,N_10433,N_11047);
nor U11774 (N_11774,N_10075,N_10896);
nor U11775 (N_11775,N_10128,N_10905);
xnor U11776 (N_11776,N_11116,N_10698);
and U11777 (N_11777,N_10663,N_10305);
nor U11778 (N_11778,N_10387,N_10015);
or U11779 (N_11779,N_10308,N_10836);
nand U11780 (N_11780,N_10675,N_11157);
or U11781 (N_11781,N_10440,N_10546);
nor U11782 (N_11782,N_10597,N_10383);
or U11783 (N_11783,N_10044,N_10429);
or U11784 (N_11784,N_10418,N_10095);
or U11785 (N_11785,N_10448,N_10989);
or U11786 (N_11786,N_10492,N_11190);
nor U11787 (N_11787,N_10109,N_11238);
nand U11788 (N_11788,N_10949,N_10749);
xor U11789 (N_11789,N_10540,N_10754);
or U11790 (N_11790,N_10486,N_10563);
nand U11791 (N_11791,N_11101,N_11226);
nand U11792 (N_11792,N_10839,N_10471);
xor U11793 (N_11793,N_11154,N_10269);
or U11794 (N_11794,N_10505,N_10472);
nor U11795 (N_11795,N_10738,N_10923);
and U11796 (N_11796,N_10138,N_11135);
nor U11797 (N_11797,N_10539,N_10908);
or U11798 (N_11798,N_10653,N_11014);
nand U11799 (N_11799,N_10191,N_10816);
xnor U11800 (N_11800,N_10361,N_11102);
or U11801 (N_11801,N_10157,N_11168);
nor U11802 (N_11802,N_10307,N_10973);
nor U11803 (N_11803,N_10247,N_10833);
or U11804 (N_11804,N_10242,N_11239);
nor U11805 (N_11805,N_10756,N_10921);
and U11806 (N_11806,N_10224,N_10944);
or U11807 (N_11807,N_10470,N_10098);
xor U11808 (N_11808,N_10403,N_11007);
or U11809 (N_11809,N_10554,N_10961);
nand U11810 (N_11810,N_10239,N_11079);
or U11811 (N_11811,N_11124,N_10947);
and U11812 (N_11812,N_10476,N_10465);
or U11813 (N_11813,N_10501,N_10555);
or U11814 (N_11814,N_10682,N_10069);
or U11815 (N_11815,N_10827,N_10085);
xnor U11816 (N_11816,N_10093,N_10757);
and U11817 (N_11817,N_11149,N_10844);
xor U11818 (N_11818,N_10499,N_10919);
xor U11819 (N_11819,N_10211,N_10801);
or U11820 (N_11820,N_11044,N_10527);
or U11821 (N_11821,N_10583,N_10250);
nor U11822 (N_11822,N_10057,N_10196);
xor U11823 (N_11823,N_10297,N_11172);
nand U11824 (N_11824,N_11167,N_10009);
nand U11825 (N_11825,N_10917,N_10365);
and U11826 (N_11826,N_10826,N_10582);
nor U11827 (N_11827,N_10787,N_10773);
nand U11828 (N_11828,N_10241,N_11248);
nand U11829 (N_11829,N_11076,N_10760);
xnor U11830 (N_11830,N_11077,N_10171);
and U11831 (N_11831,N_11221,N_10195);
or U11832 (N_11832,N_10397,N_10084);
or U11833 (N_11833,N_10559,N_10162);
nor U11834 (N_11834,N_10542,N_10785);
xnor U11835 (N_11835,N_10112,N_10493);
or U11836 (N_11836,N_10759,N_10620);
nor U11837 (N_11837,N_10362,N_10530);
xor U11838 (N_11838,N_10066,N_10025);
xor U11839 (N_11839,N_10820,N_10319);
nand U11840 (N_11840,N_11187,N_10197);
nand U11841 (N_11841,N_10740,N_10341);
nand U11842 (N_11842,N_11038,N_10187);
and U11843 (N_11843,N_10590,N_10979);
and U11844 (N_11844,N_10119,N_10102);
and U11845 (N_11845,N_10079,N_10427);
and U11846 (N_11846,N_11166,N_10595);
xnor U11847 (N_11847,N_10962,N_10885);
or U11848 (N_11848,N_10764,N_10255);
or U11849 (N_11849,N_10796,N_11046);
nor U11850 (N_11850,N_10041,N_10375);
nor U11851 (N_11851,N_11213,N_10290);
and U11852 (N_11852,N_10978,N_11171);
or U11853 (N_11853,N_10167,N_10971);
and U11854 (N_11854,N_10221,N_10019);
or U11855 (N_11855,N_10584,N_11078);
xor U11856 (N_11856,N_10252,N_10490);
or U11857 (N_11857,N_11060,N_11109);
xnor U11858 (N_11858,N_10806,N_10014);
and U11859 (N_11859,N_10879,N_10970);
xnor U11860 (N_11860,N_10177,N_11062);
nand U11861 (N_11861,N_11146,N_10790);
or U11862 (N_11862,N_10734,N_11193);
xor U11863 (N_11863,N_10356,N_10304);
and U11864 (N_11864,N_11159,N_10982);
nand U11865 (N_11865,N_10521,N_11242);
nor U11866 (N_11866,N_10813,N_11140);
and U11867 (N_11867,N_10118,N_10882);
xnor U11868 (N_11868,N_10835,N_10077);
or U11869 (N_11869,N_10819,N_11036);
nor U11870 (N_11870,N_10146,N_10059);
xnor U11871 (N_11871,N_11080,N_10674);
nand U11872 (N_11872,N_11210,N_10547);
xor U11873 (N_11873,N_11184,N_10633);
and U11874 (N_11874,N_10450,N_10886);
nand U11875 (N_11875,N_10578,N_10417);
or U11876 (N_11876,N_10877,N_10242);
nand U11877 (N_11877,N_11146,N_10978);
nand U11878 (N_11878,N_10520,N_10343);
xor U11879 (N_11879,N_10206,N_10078);
nor U11880 (N_11880,N_11043,N_10520);
nand U11881 (N_11881,N_10089,N_11036);
nand U11882 (N_11882,N_11129,N_10058);
or U11883 (N_11883,N_11002,N_10057);
and U11884 (N_11884,N_11205,N_10010);
and U11885 (N_11885,N_10906,N_10342);
and U11886 (N_11886,N_10620,N_10999);
xnor U11887 (N_11887,N_11021,N_10796);
xor U11888 (N_11888,N_10891,N_10839);
and U11889 (N_11889,N_10546,N_11193);
nand U11890 (N_11890,N_11214,N_11129);
and U11891 (N_11891,N_10067,N_10871);
xnor U11892 (N_11892,N_11167,N_10373);
nor U11893 (N_11893,N_10554,N_11165);
nand U11894 (N_11894,N_10789,N_11072);
xor U11895 (N_11895,N_10951,N_10612);
or U11896 (N_11896,N_10096,N_10964);
xnor U11897 (N_11897,N_10643,N_10277);
xnor U11898 (N_11898,N_10763,N_11078);
nor U11899 (N_11899,N_10683,N_11226);
xnor U11900 (N_11900,N_10590,N_10511);
nand U11901 (N_11901,N_10619,N_10608);
or U11902 (N_11902,N_10950,N_10614);
and U11903 (N_11903,N_10595,N_10614);
nand U11904 (N_11904,N_10973,N_10523);
nand U11905 (N_11905,N_10346,N_10480);
and U11906 (N_11906,N_10301,N_10837);
or U11907 (N_11907,N_10723,N_10775);
and U11908 (N_11908,N_10964,N_10818);
nand U11909 (N_11909,N_10679,N_11192);
xnor U11910 (N_11910,N_10448,N_10835);
nand U11911 (N_11911,N_10317,N_11116);
xor U11912 (N_11912,N_10150,N_10017);
nand U11913 (N_11913,N_10165,N_11177);
or U11914 (N_11914,N_11108,N_10793);
nor U11915 (N_11915,N_11098,N_11241);
or U11916 (N_11916,N_10711,N_10244);
or U11917 (N_11917,N_11024,N_11145);
and U11918 (N_11918,N_10682,N_10690);
or U11919 (N_11919,N_11086,N_10691);
and U11920 (N_11920,N_11096,N_10175);
nand U11921 (N_11921,N_10032,N_10508);
and U11922 (N_11922,N_10397,N_10354);
and U11923 (N_11923,N_10575,N_11236);
nor U11924 (N_11924,N_10026,N_10876);
and U11925 (N_11925,N_10772,N_10449);
xnor U11926 (N_11926,N_10536,N_10260);
or U11927 (N_11927,N_11006,N_10259);
xnor U11928 (N_11928,N_10519,N_10639);
nand U11929 (N_11929,N_11017,N_11199);
or U11930 (N_11930,N_10101,N_10309);
and U11931 (N_11931,N_11213,N_11069);
or U11932 (N_11932,N_10139,N_10271);
nor U11933 (N_11933,N_10633,N_10322);
or U11934 (N_11934,N_10227,N_11143);
or U11935 (N_11935,N_10053,N_10227);
nor U11936 (N_11936,N_10098,N_11139);
xnor U11937 (N_11937,N_10128,N_10056);
or U11938 (N_11938,N_11105,N_10224);
or U11939 (N_11939,N_10145,N_10278);
and U11940 (N_11940,N_10555,N_11000);
and U11941 (N_11941,N_10024,N_10963);
or U11942 (N_11942,N_10996,N_10679);
or U11943 (N_11943,N_10563,N_10564);
nand U11944 (N_11944,N_10842,N_10558);
and U11945 (N_11945,N_11064,N_10393);
and U11946 (N_11946,N_10861,N_11175);
or U11947 (N_11947,N_10458,N_10043);
and U11948 (N_11948,N_10750,N_10832);
and U11949 (N_11949,N_10776,N_10229);
xor U11950 (N_11950,N_10536,N_10986);
nand U11951 (N_11951,N_10545,N_10943);
nand U11952 (N_11952,N_10086,N_10160);
or U11953 (N_11953,N_10977,N_10795);
and U11954 (N_11954,N_11102,N_10544);
or U11955 (N_11955,N_10828,N_10948);
xnor U11956 (N_11956,N_10203,N_10041);
nor U11957 (N_11957,N_10712,N_10092);
or U11958 (N_11958,N_10549,N_10627);
or U11959 (N_11959,N_10660,N_10139);
and U11960 (N_11960,N_10023,N_10294);
and U11961 (N_11961,N_11241,N_10035);
nand U11962 (N_11962,N_10986,N_10034);
nand U11963 (N_11963,N_10942,N_11200);
or U11964 (N_11964,N_11056,N_10521);
nor U11965 (N_11965,N_10678,N_10229);
nor U11966 (N_11966,N_10661,N_10997);
or U11967 (N_11967,N_10216,N_10425);
xor U11968 (N_11968,N_10856,N_10770);
xnor U11969 (N_11969,N_10598,N_10661);
nand U11970 (N_11970,N_10858,N_10307);
or U11971 (N_11971,N_10455,N_11205);
nand U11972 (N_11972,N_10203,N_10611);
or U11973 (N_11973,N_11141,N_10142);
nand U11974 (N_11974,N_10245,N_10634);
nor U11975 (N_11975,N_10365,N_10005);
nand U11976 (N_11976,N_10477,N_10387);
xnor U11977 (N_11977,N_11129,N_11014);
and U11978 (N_11978,N_11187,N_10240);
or U11979 (N_11979,N_10842,N_10576);
nand U11980 (N_11980,N_10246,N_10449);
nor U11981 (N_11981,N_10629,N_10501);
nand U11982 (N_11982,N_10532,N_10612);
or U11983 (N_11983,N_10365,N_10023);
nor U11984 (N_11984,N_11039,N_11172);
nand U11985 (N_11985,N_10119,N_10318);
and U11986 (N_11986,N_10646,N_10286);
nand U11987 (N_11987,N_10488,N_10173);
or U11988 (N_11988,N_11065,N_10363);
xnor U11989 (N_11989,N_10646,N_10250);
nand U11990 (N_11990,N_10048,N_10029);
xnor U11991 (N_11991,N_10933,N_10968);
xnor U11992 (N_11992,N_10466,N_10689);
nand U11993 (N_11993,N_10328,N_10659);
or U11994 (N_11994,N_10638,N_10014);
and U11995 (N_11995,N_10272,N_10604);
nor U11996 (N_11996,N_10236,N_11161);
or U11997 (N_11997,N_10820,N_10980);
and U11998 (N_11998,N_11093,N_11115);
and U11999 (N_11999,N_11073,N_11179);
and U12000 (N_12000,N_11137,N_10592);
or U12001 (N_12001,N_10191,N_10001);
nor U12002 (N_12002,N_10301,N_11245);
xnor U12003 (N_12003,N_10280,N_10073);
and U12004 (N_12004,N_10230,N_10044);
and U12005 (N_12005,N_10231,N_10349);
nor U12006 (N_12006,N_10753,N_11145);
xor U12007 (N_12007,N_10921,N_10920);
and U12008 (N_12008,N_11199,N_10903);
nor U12009 (N_12009,N_11212,N_10886);
nor U12010 (N_12010,N_10216,N_10066);
and U12011 (N_12011,N_10045,N_10292);
nand U12012 (N_12012,N_10097,N_10936);
xnor U12013 (N_12013,N_11246,N_11165);
nand U12014 (N_12014,N_10677,N_10944);
nand U12015 (N_12015,N_10949,N_11028);
nor U12016 (N_12016,N_10835,N_10516);
nor U12017 (N_12017,N_10293,N_10823);
or U12018 (N_12018,N_10720,N_10217);
xor U12019 (N_12019,N_11033,N_11073);
and U12020 (N_12020,N_10060,N_10685);
or U12021 (N_12021,N_10496,N_10999);
or U12022 (N_12022,N_10028,N_10462);
or U12023 (N_12023,N_10879,N_10501);
nand U12024 (N_12024,N_10299,N_10691);
or U12025 (N_12025,N_10421,N_10101);
xor U12026 (N_12026,N_10759,N_10399);
and U12027 (N_12027,N_10475,N_10770);
and U12028 (N_12028,N_10402,N_10519);
nand U12029 (N_12029,N_11190,N_10560);
nor U12030 (N_12030,N_10924,N_10081);
nor U12031 (N_12031,N_10543,N_10734);
nand U12032 (N_12032,N_10440,N_10921);
and U12033 (N_12033,N_10314,N_10255);
and U12034 (N_12034,N_10683,N_11088);
xor U12035 (N_12035,N_10826,N_10747);
or U12036 (N_12036,N_10596,N_10752);
nand U12037 (N_12037,N_11228,N_10335);
xor U12038 (N_12038,N_10721,N_10438);
xor U12039 (N_12039,N_10491,N_10266);
or U12040 (N_12040,N_10426,N_10291);
or U12041 (N_12041,N_10304,N_11229);
xor U12042 (N_12042,N_10830,N_10764);
nand U12043 (N_12043,N_10972,N_10691);
and U12044 (N_12044,N_10879,N_10472);
xnor U12045 (N_12045,N_10764,N_10963);
or U12046 (N_12046,N_10714,N_11100);
or U12047 (N_12047,N_10047,N_10571);
or U12048 (N_12048,N_10376,N_10202);
nand U12049 (N_12049,N_11008,N_10314);
xnor U12050 (N_12050,N_10989,N_10286);
nor U12051 (N_12051,N_10107,N_10959);
nor U12052 (N_12052,N_10625,N_10887);
xor U12053 (N_12053,N_10447,N_10911);
nand U12054 (N_12054,N_10832,N_10243);
xnor U12055 (N_12055,N_10899,N_11033);
or U12056 (N_12056,N_10669,N_10749);
and U12057 (N_12057,N_10705,N_10429);
and U12058 (N_12058,N_10278,N_10365);
xor U12059 (N_12059,N_10298,N_10452);
nand U12060 (N_12060,N_11239,N_11113);
and U12061 (N_12061,N_10674,N_11032);
nor U12062 (N_12062,N_10531,N_10982);
nor U12063 (N_12063,N_10828,N_11176);
and U12064 (N_12064,N_11055,N_10086);
nor U12065 (N_12065,N_11137,N_11145);
nor U12066 (N_12066,N_11018,N_10183);
and U12067 (N_12067,N_10503,N_10905);
or U12068 (N_12068,N_10877,N_10418);
or U12069 (N_12069,N_11041,N_10844);
nand U12070 (N_12070,N_11213,N_11070);
nand U12071 (N_12071,N_10381,N_10828);
xor U12072 (N_12072,N_10484,N_11096);
nand U12073 (N_12073,N_10363,N_10569);
or U12074 (N_12074,N_10097,N_10719);
nor U12075 (N_12075,N_10288,N_11010);
or U12076 (N_12076,N_10491,N_10762);
xor U12077 (N_12077,N_10184,N_11035);
nand U12078 (N_12078,N_10325,N_10004);
nor U12079 (N_12079,N_10797,N_10554);
nand U12080 (N_12080,N_10160,N_10710);
and U12081 (N_12081,N_10844,N_10031);
and U12082 (N_12082,N_10967,N_11180);
or U12083 (N_12083,N_10123,N_11060);
nor U12084 (N_12084,N_10753,N_10484);
or U12085 (N_12085,N_10756,N_10336);
nand U12086 (N_12086,N_10778,N_10607);
nand U12087 (N_12087,N_10144,N_10244);
and U12088 (N_12088,N_10355,N_10058);
nand U12089 (N_12089,N_10779,N_11209);
and U12090 (N_12090,N_10363,N_10844);
nand U12091 (N_12091,N_11016,N_10607);
nand U12092 (N_12092,N_11167,N_10947);
nor U12093 (N_12093,N_10625,N_10508);
nand U12094 (N_12094,N_11101,N_10277);
or U12095 (N_12095,N_11120,N_10247);
nor U12096 (N_12096,N_10466,N_10037);
nor U12097 (N_12097,N_10488,N_10501);
nor U12098 (N_12098,N_10168,N_10272);
and U12099 (N_12099,N_10926,N_10610);
and U12100 (N_12100,N_10461,N_10702);
and U12101 (N_12101,N_10696,N_11103);
or U12102 (N_12102,N_10108,N_10626);
nand U12103 (N_12103,N_10984,N_10640);
and U12104 (N_12104,N_10316,N_11177);
or U12105 (N_12105,N_10723,N_10957);
and U12106 (N_12106,N_10391,N_10660);
nand U12107 (N_12107,N_10281,N_10527);
or U12108 (N_12108,N_10422,N_11172);
or U12109 (N_12109,N_11001,N_11225);
or U12110 (N_12110,N_10862,N_10476);
and U12111 (N_12111,N_10901,N_10829);
nand U12112 (N_12112,N_11005,N_10502);
and U12113 (N_12113,N_11110,N_10225);
nor U12114 (N_12114,N_10036,N_10745);
nor U12115 (N_12115,N_10143,N_10466);
xor U12116 (N_12116,N_10810,N_10534);
and U12117 (N_12117,N_11168,N_11126);
or U12118 (N_12118,N_11137,N_10871);
or U12119 (N_12119,N_10714,N_10370);
and U12120 (N_12120,N_10316,N_11208);
nand U12121 (N_12121,N_11194,N_10096);
and U12122 (N_12122,N_10496,N_11052);
nand U12123 (N_12123,N_10728,N_11221);
or U12124 (N_12124,N_10667,N_10850);
nand U12125 (N_12125,N_10492,N_10302);
nor U12126 (N_12126,N_11160,N_10458);
xnor U12127 (N_12127,N_10345,N_10351);
or U12128 (N_12128,N_10850,N_10732);
xnor U12129 (N_12129,N_10051,N_11035);
nand U12130 (N_12130,N_10106,N_10384);
or U12131 (N_12131,N_10587,N_10533);
nand U12132 (N_12132,N_10522,N_11177);
xnor U12133 (N_12133,N_10800,N_11053);
nand U12134 (N_12134,N_11153,N_10667);
nor U12135 (N_12135,N_11002,N_10486);
nand U12136 (N_12136,N_10571,N_10667);
and U12137 (N_12137,N_10362,N_11115);
nor U12138 (N_12138,N_11073,N_10848);
nor U12139 (N_12139,N_10278,N_10832);
or U12140 (N_12140,N_10032,N_10787);
nand U12141 (N_12141,N_10088,N_11047);
and U12142 (N_12142,N_10788,N_10314);
nand U12143 (N_12143,N_10390,N_10276);
xnor U12144 (N_12144,N_10658,N_11201);
nand U12145 (N_12145,N_10722,N_10820);
nor U12146 (N_12146,N_10002,N_11125);
xor U12147 (N_12147,N_10784,N_11025);
xnor U12148 (N_12148,N_10442,N_10529);
xor U12149 (N_12149,N_10969,N_10930);
nor U12150 (N_12150,N_10814,N_10199);
xnor U12151 (N_12151,N_10039,N_10239);
and U12152 (N_12152,N_10072,N_10359);
xor U12153 (N_12153,N_11130,N_10553);
or U12154 (N_12154,N_10968,N_11088);
xnor U12155 (N_12155,N_11060,N_10792);
nand U12156 (N_12156,N_10599,N_10726);
xor U12157 (N_12157,N_10830,N_11223);
nor U12158 (N_12158,N_11138,N_10831);
nor U12159 (N_12159,N_10015,N_11000);
or U12160 (N_12160,N_10639,N_10164);
nand U12161 (N_12161,N_10470,N_10411);
nor U12162 (N_12162,N_10584,N_10058);
and U12163 (N_12163,N_10902,N_10051);
nand U12164 (N_12164,N_10030,N_11003);
nand U12165 (N_12165,N_11238,N_11057);
nor U12166 (N_12166,N_10738,N_10518);
xor U12167 (N_12167,N_11173,N_10313);
or U12168 (N_12168,N_10462,N_11113);
nor U12169 (N_12169,N_10468,N_10298);
nor U12170 (N_12170,N_10968,N_10130);
nor U12171 (N_12171,N_10771,N_10541);
or U12172 (N_12172,N_10325,N_10406);
nor U12173 (N_12173,N_10859,N_10287);
or U12174 (N_12174,N_10771,N_10873);
nor U12175 (N_12175,N_10478,N_10094);
or U12176 (N_12176,N_10760,N_10873);
or U12177 (N_12177,N_10768,N_10181);
nor U12178 (N_12178,N_11079,N_10289);
xnor U12179 (N_12179,N_10801,N_10405);
nor U12180 (N_12180,N_10997,N_10248);
and U12181 (N_12181,N_10200,N_10516);
xnor U12182 (N_12182,N_10791,N_10776);
or U12183 (N_12183,N_10212,N_11204);
nor U12184 (N_12184,N_10339,N_10702);
xnor U12185 (N_12185,N_10038,N_10319);
or U12186 (N_12186,N_10968,N_10014);
xor U12187 (N_12187,N_11248,N_10482);
xor U12188 (N_12188,N_10897,N_11199);
and U12189 (N_12189,N_10343,N_11117);
xnor U12190 (N_12190,N_10001,N_10693);
and U12191 (N_12191,N_10913,N_10649);
nor U12192 (N_12192,N_10507,N_10078);
nand U12193 (N_12193,N_10779,N_10082);
nand U12194 (N_12194,N_11173,N_10718);
nor U12195 (N_12195,N_10417,N_10675);
nand U12196 (N_12196,N_11223,N_10102);
nor U12197 (N_12197,N_11053,N_10659);
xnor U12198 (N_12198,N_10855,N_10162);
or U12199 (N_12199,N_11083,N_10224);
xor U12200 (N_12200,N_10226,N_10690);
or U12201 (N_12201,N_10174,N_11190);
nor U12202 (N_12202,N_10684,N_11143);
xnor U12203 (N_12203,N_10124,N_11003);
xor U12204 (N_12204,N_10151,N_10510);
and U12205 (N_12205,N_10521,N_10663);
or U12206 (N_12206,N_11126,N_11103);
xor U12207 (N_12207,N_10412,N_10051);
nand U12208 (N_12208,N_10446,N_10358);
nand U12209 (N_12209,N_10904,N_10660);
and U12210 (N_12210,N_10799,N_10624);
xor U12211 (N_12211,N_10904,N_10467);
nand U12212 (N_12212,N_10800,N_10622);
and U12213 (N_12213,N_10880,N_10585);
xnor U12214 (N_12214,N_11143,N_10460);
xnor U12215 (N_12215,N_10139,N_11123);
nand U12216 (N_12216,N_10551,N_10737);
xor U12217 (N_12217,N_10929,N_10094);
and U12218 (N_12218,N_10803,N_10485);
nand U12219 (N_12219,N_10461,N_10268);
nand U12220 (N_12220,N_10714,N_10411);
nand U12221 (N_12221,N_10420,N_10013);
xor U12222 (N_12222,N_10967,N_10753);
nor U12223 (N_12223,N_11071,N_11092);
and U12224 (N_12224,N_10713,N_10851);
nor U12225 (N_12225,N_11228,N_11244);
xor U12226 (N_12226,N_10867,N_10202);
nor U12227 (N_12227,N_10200,N_10322);
nand U12228 (N_12228,N_10935,N_10140);
and U12229 (N_12229,N_10770,N_11038);
nand U12230 (N_12230,N_10617,N_10606);
nand U12231 (N_12231,N_11165,N_10187);
or U12232 (N_12232,N_10170,N_10848);
nor U12233 (N_12233,N_10945,N_10752);
nand U12234 (N_12234,N_11040,N_10080);
and U12235 (N_12235,N_10183,N_10703);
and U12236 (N_12236,N_10245,N_11137);
and U12237 (N_12237,N_10533,N_10089);
nor U12238 (N_12238,N_10860,N_10521);
nand U12239 (N_12239,N_10041,N_11123);
or U12240 (N_12240,N_10430,N_11241);
nand U12241 (N_12241,N_10996,N_10072);
xnor U12242 (N_12242,N_11095,N_10565);
and U12243 (N_12243,N_10497,N_10366);
nor U12244 (N_12244,N_10306,N_10343);
or U12245 (N_12245,N_10764,N_11151);
or U12246 (N_12246,N_10103,N_10213);
or U12247 (N_12247,N_10584,N_10582);
and U12248 (N_12248,N_10588,N_10405);
nand U12249 (N_12249,N_11184,N_10773);
nand U12250 (N_12250,N_11188,N_10541);
nor U12251 (N_12251,N_11003,N_10500);
nor U12252 (N_12252,N_10229,N_10536);
and U12253 (N_12253,N_10667,N_10171);
nand U12254 (N_12254,N_10936,N_11147);
nand U12255 (N_12255,N_11015,N_11108);
and U12256 (N_12256,N_11246,N_11121);
nor U12257 (N_12257,N_10693,N_10286);
nor U12258 (N_12258,N_10943,N_10779);
or U12259 (N_12259,N_10647,N_10358);
xnor U12260 (N_12260,N_11150,N_11248);
or U12261 (N_12261,N_11126,N_11237);
or U12262 (N_12262,N_10164,N_10274);
nor U12263 (N_12263,N_10344,N_10183);
and U12264 (N_12264,N_11050,N_10786);
and U12265 (N_12265,N_10093,N_10180);
xnor U12266 (N_12266,N_11181,N_10644);
or U12267 (N_12267,N_11124,N_10918);
xor U12268 (N_12268,N_10936,N_11032);
or U12269 (N_12269,N_11207,N_10733);
nand U12270 (N_12270,N_10179,N_10198);
nand U12271 (N_12271,N_10714,N_10081);
and U12272 (N_12272,N_10195,N_11192);
or U12273 (N_12273,N_10045,N_10731);
and U12274 (N_12274,N_10756,N_10127);
and U12275 (N_12275,N_11176,N_10570);
xor U12276 (N_12276,N_10066,N_10497);
and U12277 (N_12277,N_10366,N_10342);
nor U12278 (N_12278,N_10590,N_10081);
and U12279 (N_12279,N_10825,N_10084);
nor U12280 (N_12280,N_10929,N_10184);
or U12281 (N_12281,N_10331,N_11060);
and U12282 (N_12282,N_11161,N_10380);
nor U12283 (N_12283,N_11244,N_10837);
xnor U12284 (N_12284,N_10536,N_11190);
nor U12285 (N_12285,N_10462,N_10006);
xor U12286 (N_12286,N_10012,N_10017);
nor U12287 (N_12287,N_10295,N_10164);
nand U12288 (N_12288,N_10700,N_10208);
and U12289 (N_12289,N_11082,N_10678);
and U12290 (N_12290,N_10639,N_10631);
xor U12291 (N_12291,N_10342,N_11010);
xor U12292 (N_12292,N_10156,N_10816);
nor U12293 (N_12293,N_10221,N_11047);
nor U12294 (N_12294,N_10044,N_11122);
and U12295 (N_12295,N_11042,N_10594);
or U12296 (N_12296,N_10493,N_11239);
xor U12297 (N_12297,N_11196,N_10824);
or U12298 (N_12298,N_10924,N_10236);
xor U12299 (N_12299,N_11165,N_10586);
xnor U12300 (N_12300,N_10929,N_10328);
or U12301 (N_12301,N_11174,N_10390);
nand U12302 (N_12302,N_10364,N_10704);
nor U12303 (N_12303,N_10614,N_10745);
and U12304 (N_12304,N_10745,N_10404);
xor U12305 (N_12305,N_11075,N_11167);
nand U12306 (N_12306,N_11236,N_10595);
nand U12307 (N_12307,N_10315,N_10969);
or U12308 (N_12308,N_10937,N_10089);
xor U12309 (N_12309,N_10924,N_10193);
nor U12310 (N_12310,N_10157,N_10519);
nor U12311 (N_12311,N_10157,N_10769);
and U12312 (N_12312,N_10265,N_10030);
xor U12313 (N_12313,N_11124,N_11142);
xnor U12314 (N_12314,N_10693,N_11064);
xnor U12315 (N_12315,N_10364,N_10874);
nand U12316 (N_12316,N_10847,N_10471);
xor U12317 (N_12317,N_10711,N_11057);
xnor U12318 (N_12318,N_10081,N_10564);
nor U12319 (N_12319,N_10708,N_10353);
nand U12320 (N_12320,N_10460,N_10303);
nor U12321 (N_12321,N_10105,N_10737);
nor U12322 (N_12322,N_10737,N_10770);
xor U12323 (N_12323,N_10840,N_10212);
nand U12324 (N_12324,N_11215,N_10540);
nor U12325 (N_12325,N_11211,N_11065);
and U12326 (N_12326,N_10954,N_10436);
nor U12327 (N_12327,N_10460,N_11210);
or U12328 (N_12328,N_10500,N_11134);
and U12329 (N_12329,N_10054,N_10283);
and U12330 (N_12330,N_10119,N_11046);
xnor U12331 (N_12331,N_10935,N_10096);
or U12332 (N_12332,N_10011,N_11217);
nor U12333 (N_12333,N_10234,N_10905);
or U12334 (N_12334,N_10392,N_10364);
xor U12335 (N_12335,N_10412,N_11172);
nor U12336 (N_12336,N_10186,N_10138);
and U12337 (N_12337,N_11179,N_10817);
xor U12338 (N_12338,N_11036,N_10118);
nand U12339 (N_12339,N_10533,N_10813);
and U12340 (N_12340,N_10263,N_10821);
or U12341 (N_12341,N_10531,N_10901);
nand U12342 (N_12342,N_11163,N_10597);
nor U12343 (N_12343,N_10563,N_11008);
and U12344 (N_12344,N_11147,N_11213);
nor U12345 (N_12345,N_10407,N_11182);
and U12346 (N_12346,N_10149,N_11026);
xor U12347 (N_12347,N_10374,N_10547);
and U12348 (N_12348,N_10828,N_10902);
nor U12349 (N_12349,N_11154,N_10886);
nand U12350 (N_12350,N_10666,N_10971);
nor U12351 (N_12351,N_10878,N_11180);
xnor U12352 (N_12352,N_11136,N_11234);
nand U12353 (N_12353,N_10250,N_10432);
xor U12354 (N_12354,N_11082,N_10881);
xor U12355 (N_12355,N_11176,N_10288);
xnor U12356 (N_12356,N_10030,N_10833);
nor U12357 (N_12357,N_11099,N_10406);
nand U12358 (N_12358,N_11235,N_10800);
and U12359 (N_12359,N_10988,N_10619);
nand U12360 (N_12360,N_10100,N_10152);
and U12361 (N_12361,N_10526,N_10032);
or U12362 (N_12362,N_10616,N_10319);
or U12363 (N_12363,N_11192,N_11028);
or U12364 (N_12364,N_10299,N_10779);
and U12365 (N_12365,N_10150,N_10546);
and U12366 (N_12366,N_10240,N_10237);
or U12367 (N_12367,N_11030,N_10904);
nand U12368 (N_12368,N_10830,N_10481);
xnor U12369 (N_12369,N_10780,N_10389);
nor U12370 (N_12370,N_10182,N_10731);
or U12371 (N_12371,N_10402,N_11155);
or U12372 (N_12372,N_11116,N_10155);
or U12373 (N_12373,N_10742,N_10324);
and U12374 (N_12374,N_10239,N_10428);
or U12375 (N_12375,N_11116,N_10355);
nor U12376 (N_12376,N_10497,N_10135);
xor U12377 (N_12377,N_10852,N_10810);
or U12378 (N_12378,N_10135,N_10066);
xor U12379 (N_12379,N_10280,N_11079);
nand U12380 (N_12380,N_10311,N_10044);
or U12381 (N_12381,N_11129,N_11117);
or U12382 (N_12382,N_10745,N_10296);
and U12383 (N_12383,N_11184,N_10760);
xor U12384 (N_12384,N_10031,N_10731);
and U12385 (N_12385,N_10610,N_11057);
nand U12386 (N_12386,N_11060,N_11095);
and U12387 (N_12387,N_11128,N_10182);
nor U12388 (N_12388,N_10450,N_10125);
or U12389 (N_12389,N_11131,N_10237);
and U12390 (N_12390,N_10878,N_10964);
nor U12391 (N_12391,N_10464,N_10613);
or U12392 (N_12392,N_10032,N_10353);
xnor U12393 (N_12393,N_10858,N_11023);
nor U12394 (N_12394,N_10793,N_11153);
nand U12395 (N_12395,N_10106,N_11235);
and U12396 (N_12396,N_10306,N_10345);
nand U12397 (N_12397,N_10610,N_10438);
nor U12398 (N_12398,N_10714,N_10419);
nand U12399 (N_12399,N_10155,N_10349);
and U12400 (N_12400,N_11161,N_10949);
xor U12401 (N_12401,N_10264,N_10808);
xnor U12402 (N_12402,N_10232,N_10056);
nor U12403 (N_12403,N_10796,N_10280);
and U12404 (N_12404,N_10633,N_11047);
nand U12405 (N_12405,N_11096,N_11236);
and U12406 (N_12406,N_10167,N_11176);
nor U12407 (N_12407,N_10893,N_10843);
or U12408 (N_12408,N_10380,N_10444);
nand U12409 (N_12409,N_10381,N_10167);
or U12410 (N_12410,N_10838,N_10652);
or U12411 (N_12411,N_10160,N_10756);
nand U12412 (N_12412,N_10407,N_10398);
nand U12413 (N_12413,N_10948,N_11009);
nor U12414 (N_12414,N_10728,N_10508);
or U12415 (N_12415,N_10291,N_10289);
xnor U12416 (N_12416,N_10217,N_11059);
nor U12417 (N_12417,N_11085,N_10684);
and U12418 (N_12418,N_10768,N_10995);
nor U12419 (N_12419,N_11044,N_10689);
xnor U12420 (N_12420,N_10300,N_11129);
nand U12421 (N_12421,N_10217,N_10664);
nand U12422 (N_12422,N_10935,N_10828);
xor U12423 (N_12423,N_10900,N_10425);
nor U12424 (N_12424,N_10396,N_10724);
and U12425 (N_12425,N_10318,N_10745);
or U12426 (N_12426,N_11091,N_11228);
nand U12427 (N_12427,N_10342,N_10733);
and U12428 (N_12428,N_10331,N_10985);
xnor U12429 (N_12429,N_11137,N_10469);
nor U12430 (N_12430,N_10197,N_10350);
xnor U12431 (N_12431,N_10217,N_10695);
and U12432 (N_12432,N_10861,N_10438);
nand U12433 (N_12433,N_10286,N_10984);
nand U12434 (N_12434,N_10810,N_11063);
and U12435 (N_12435,N_10747,N_11040);
nand U12436 (N_12436,N_10567,N_11032);
nand U12437 (N_12437,N_10995,N_10392);
or U12438 (N_12438,N_11189,N_10312);
or U12439 (N_12439,N_11108,N_10316);
nand U12440 (N_12440,N_11015,N_11051);
and U12441 (N_12441,N_11218,N_10602);
xor U12442 (N_12442,N_10350,N_10477);
xnor U12443 (N_12443,N_10948,N_10515);
xnor U12444 (N_12444,N_10847,N_10318);
nand U12445 (N_12445,N_10069,N_10456);
or U12446 (N_12446,N_10196,N_10712);
nand U12447 (N_12447,N_11097,N_10751);
nand U12448 (N_12448,N_10566,N_10407);
nand U12449 (N_12449,N_10293,N_10562);
xnor U12450 (N_12450,N_10368,N_11167);
xnor U12451 (N_12451,N_10232,N_10736);
nor U12452 (N_12452,N_10527,N_10517);
nor U12453 (N_12453,N_10731,N_10662);
nand U12454 (N_12454,N_10488,N_10726);
xnor U12455 (N_12455,N_10108,N_10847);
or U12456 (N_12456,N_11232,N_10403);
xnor U12457 (N_12457,N_10964,N_10909);
or U12458 (N_12458,N_10690,N_11144);
nor U12459 (N_12459,N_10059,N_10907);
xnor U12460 (N_12460,N_10512,N_10991);
xnor U12461 (N_12461,N_10573,N_10960);
nand U12462 (N_12462,N_11019,N_11112);
and U12463 (N_12463,N_10704,N_10846);
and U12464 (N_12464,N_10461,N_10088);
and U12465 (N_12465,N_10122,N_10961);
xnor U12466 (N_12466,N_11079,N_10046);
or U12467 (N_12467,N_10859,N_10297);
nor U12468 (N_12468,N_10320,N_10159);
nor U12469 (N_12469,N_11099,N_10670);
or U12470 (N_12470,N_10977,N_10635);
nand U12471 (N_12471,N_10223,N_11139);
nand U12472 (N_12472,N_10976,N_10473);
nand U12473 (N_12473,N_10394,N_10963);
and U12474 (N_12474,N_10856,N_10043);
nor U12475 (N_12475,N_10986,N_10835);
nand U12476 (N_12476,N_10251,N_10893);
nor U12477 (N_12477,N_11127,N_10429);
xor U12478 (N_12478,N_10438,N_10912);
or U12479 (N_12479,N_10399,N_11082);
nor U12480 (N_12480,N_11102,N_11185);
or U12481 (N_12481,N_10701,N_10519);
xor U12482 (N_12482,N_11076,N_10553);
nor U12483 (N_12483,N_10619,N_10176);
nor U12484 (N_12484,N_11234,N_10362);
nand U12485 (N_12485,N_10512,N_10714);
xnor U12486 (N_12486,N_10221,N_10680);
or U12487 (N_12487,N_10015,N_10038);
nor U12488 (N_12488,N_10398,N_11096);
or U12489 (N_12489,N_10598,N_10476);
nand U12490 (N_12490,N_10258,N_10629);
and U12491 (N_12491,N_10688,N_11221);
or U12492 (N_12492,N_10246,N_10985);
or U12493 (N_12493,N_10105,N_11203);
and U12494 (N_12494,N_10287,N_10139);
and U12495 (N_12495,N_10943,N_11189);
or U12496 (N_12496,N_11105,N_11211);
nand U12497 (N_12497,N_10721,N_10382);
nand U12498 (N_12498,N_10334,N_10292);
nand U12499 (N_12499,N_10207,N_10839);
nand U12500 (N_12500,N_11607,N_12235);
nand U12501 (N_12501,N_11265,N_11819);
nand U12502 (N_12502,N_11801,N_12010);
or U12503 (N_12503,N_12207,N_12267);
and U12504 (N_12504,N_12009,N_11415);
and U12505 (N_12505,N_12290,N_12138);
xor U12506 (N_12506,N_11326,N_11650);
nand U12507 (N_12507,N_12310,N_11316);
nor U12508 (N_12508,N_11611,N_11598);
xnor U12509 (N_12509,N_12151,N_12278);
nor U12510 (N_12510,N_12470,N_11991);
nor U12511 (N_12511,N_11949,N_11412);
or U12512 (N_12512,N_12390,N_11643);
nor U12513 (N_12513,N_11642,N_12004);
xor U12514 (N_12514,N_11704,N_11581);
nand U12515 (N_12515,N_11453,N_12445);
and U12516 (N_12516,N_11505,N_12463);
or U12517 (N_12517,N_11706,N_12270);
or U12518 (N_12518,N_11295,N_12208);
xor U12519 (N_12519,N_11872,N_11448);
and U12520 (N_12520,N_11255,N_11383);
nand U12521 (N_12521,N_12354,N_12133);
nor U12522 (N_12522,N_11432,N_12141);
xnor U12523 (N_12523,N_11902,N_11683);
xor U12524 (N_12524,N_11889,N_12287);
nand U12525 (N_12525,N_11836,N_12122);
or U12526 (N_12526,N_12069,N_11495);
and U12527 (N_12527,N_12003,N_11551);
or U12528 (N_12528,N_11524,N_11945);
xor U12529 (N_12529,N_11484,N_11575);
nand U12530 (N_12530,N_11418,N_11437);
xor U12531 (N_12531,N_11943,N_11955);
or U12532 (N_12532,N_11413,N_11844);
or U12533 (N_12533,N_11997,N_12221);
nand U12534 (N_12534,N_12124,N_11275);
xnor U12535 (N_12535,N_11959,N_12274);
nor U12536 (N_12536,N_11749,N_11279);
nor U12537 (N_12537,N_11422,N_12259);
nand U12538 (N_12538,N_11885,N_12204);
nor U12539 (N_12539,N_11507,N_12461);
or U12540 (N_12540,N_12249,N_12349);
or U12541 (N_12541,N_11685,N_11263);
nor U12542 (N_12542,N_11332,N_12022);
nor U12543 (N_12543,N_11610,N_12321);
nor U12544 (N_12544,N_12469,N_12028);
nor U12545 (N_12545,N_11925,N_11877);
or U12546 (N_12546,N_11406,N_11501);
nor U12547 (N_12547,N_12484,N_11972);
nor U12548 (N_12548,N_12104,N_11766);
xor U12549 (N_12549,N_12228,N_11911);
xor U12550 (N_12550,N_11512,N_11975);
or U12551 (N_12551,N_12397,N_11274);
nand U12552 (N_12552,N_11591,N_11689);
and U12553 (N_12553,N_12455,N_11293);
or U12554 (N_12554,N_11903,N_12488);
xor U12555 (N_12555,N_11793,N_11761);
and U12556 (N_12556,N_12428,N_11330);
nor U12557 (N_12557,N_11417,N_11687);
nor U12558 (N_12558,N_11351,N_12113);
xor U12559 (N_12559,N_12260,N_12078);
nor U12560 (N_12560,N_11760,N_12144);
xnor U12561 (N_12561,N_11570,N_11763);
or U12562 (N_12562,N_11737,N_12370);
and U12563 (N_12563,N_12146,N_11257);
or U12564 (N_12564,N_12309,N_12190);
nor U12565 (N_12565,N_11476,N_12442);
xnor U12566 (N_12566,N_11751,N_12294);
and U12567 (N_12567,N_12498,N_11696);
nand U12568 (N_12568,N_12073,N_12376);
nor U12569 (N_12569,N_11810,N_11555);
and U12570 (N_12570,N_12191,N_11778);
nand U12571 (N_12571,N_12158,N_11800);
xnor U12572 (N_12572,N_11672,N_12060);
nand U12573 (N_12573,N_11479,N_12269);
nand U12574 (N_12574,N_12365,N_12211);
nor U12575 (N_12575,N_11654,N_12412);
nor U12576 (N_12576,N_11999,N_11742);
nand U12577 (N_12577,N_12014,N_12392);
nor U12578 (N_12578,N_12210,N_12007);
and U12579 (N_12579,N_11666,N_12074);
xnor U12580 (N_12580,N_11526,N_12458);
xor U12581 (N_12581,N_12468,N_12095);
nand U12582 (N_12582,N_11830,N_11525);
or U12583 (N_12583,N_11362,N_11770);
nand U12584 (N_12584,N_11985,N_11864);
nor U12585 (N_12585,N_11616,N_11593);
nand U12586 (N_12586,N_11335,N_12020);
nand U12587 (N_12587,N_12187,N_11967);
and U12588 (N_12588,N_12167,N_12033);
xor U12589 (N_12589,N_11857,N_11851);
or U12590 (N_12590,N_11559,N_11764);
nor U12591 (N_12591,N_12281,N_11963);
xor U12592 (N_12592,N_12040,N_11369);
and U12593 (N_12593,N_12029,N_11923);
nand U12594 (N_12594,N_12404,N_11636);
xor U12595 (N_12595,N_11807,N_11876);
xor U12596 (N_12596,N_12398,N_11387);
xnor U12597 (N_12597,N_11305,N_12465);
and U12598 (N_12598,N_11648,N_11832);
nand U12599 (N_12599,N_11269,N_11604);
and U12600 (N_12600,N_11659,N_12360);
or U12601 (N_12601,N_12177,N_11715);
nand U12602 (N_12602,N_11280,N_12082);
nor U12603 (N_12603,N_11663,N_11276);
nand U12604 (N_12604,N_11884,N_11940);
and U12605 (N_12605,N_12357,N_11894);
xnor U12606 (N_12606,N_12015,N_12233);
or U12607 (N_12607,N_11914,N_11409);
nand U12608 (N_12608,N_11865,N_11987);
nor U12609 (N_12609,N_11792,N_12178);
nand U12610 (N_12610,N_11966,N_11259);
nand U12611 (N_12611,N_12459,N_11986);
xnor U12612 (N_12612,N_12344,N_11671);
and U12613 (N_12613,N_12493,N_11717);
or U12614 (N_12614,N_12252,N_12006);
xnor U12615 (N_12615,N_12075,N_11652);
or U12616 (N_12616,N_11904,N_11386);
xnor U12617 (N_12617,N_12320,N_11932);
and U12618 (N_12618,N_11748,N_11441);
nor U12619 (N_12619,N_11818,N_11738);
xnor U12620 (N_12620,N_12254,N_11716);
and U12621 (N_12621,N_12284,N_12181);
or U12622 (N_12622,N_11374,N_11669);
nor U12623 (N_12623,N_12301,N_11393);
or U12624 (N_12624,N_11494,N_11730);
nand U12625 (N_12625,N_12486,N_11268);
and U12626 (N_12626,N_12225,N_12356);
and U12627 (N_12627,N_11912,N_12180);
and U12628 (N_12628,N_11929,N_11676);
nor U12629 (N_12629,N_12107,N_12064);
xor U12630 (N_12630,N_12044,N_12231);
nand U12631 (N_12631,N_11480,N_12026);
nor U12632 (N_12632,N_11947,N_11661);
nand U12633 (N_12633,N_11464,N_12467);
and U12634 (N_12634,N_12048,N_11303);
or U12635 (N_12635,N_11267,N_11626);
and U12636 (N_12636,N_11500,N_11796);
nor U12637 (N_12637,N_12092,N_11841);
nand U12638 (N_12638,N_11489,N_11782);
xor U12639 (N_12639,N_12099,N_11837);
nor U12640 (N_12640,N_11356,N_11511);
or U12641 (N_12641,N_11262,N_12197);
nand U12642 (N_12642,N_11371,N_11649);
and U12643 (N_12643,N_11250,N_11323);
nand U12644 (N_12644,N_11537,N_11336);
xnor U12645 (N_12645,N_11379,N_12382);
nor U12646 (N_12646,N_12426,N_12316);
xor U12647 (N_12647,N_12328,N_12169);
and U12648 (N_12648,N_12444,N_12000);
nor U12649 (N_12649,N_11514,N_12475);
nand U12650 (N_12650,N_11808,N_12080);
xor U12651 (N_12651,N_11445,N_11258);
or U12652 (N_12652,N_11523,N_11449);
nor U12653 (N_12653,N_11714,N_12372);
nor U12654 (N_12654,N_12434,N_11321);
xnor U12655 (N_12655,N_11655,N_12005);
nand U12656 (N_12656,N_12322,N_12430);
nand U12657 (N_12657,N_11868,N_11564);
or U12658 (N_12658,N_11419,N_12327);
nor U12659 (N_12659,N_11430,N_12253);
nand U12660 (N_12660,N_11855,N_12100);
nor U12661 (N_12661,N_12292,N_11314);
xor U12662 (N_12662,N_11266,N_12050);
nor U12663 (N_12663,N_11983,N_11567);
xnor U12664 (N_12664,N_11948,N_11522);
nor U12665 (N_12665,N_12352,N_12359);
nand U12666 (N_12666,N_11619,N_12237);
or U12667 (N_12667,N_11431,N_11467);
or U12668 (N_12668,N_12280,N_11623);
or U12669 (N_12669,N_12330,N_11317);
or U12670 (N_12670,N_11465,N_11497);
xor U12671 (N_12671,N_11842,N_11297);
or U12672 (N_12672,N_11906,N_11328);
nor U12673 (N_12673,N_11933,N_11550);
nor U12674 (N_12674,N_12499,N_12230);
nand U12675 (N_12675,N_11384,N_11402);
or U12676 (N_12676,N_11834,N_11828);
xnor U12677 (N_12677,N_12043,N_12325);
nor U12678 (N_12678,N_11756,N_11724);
xor U12679 (N_12679,N_12345,N_11377);
nand U12680 (N_12680,N_12192,N_11993);
or U12681 (N_12681,N_12018,N_11400);
nor U12682 (N_12682,N_11447,N_11583);
nor U12683 (N_12683,N_11839,N_11433);
or U12684 (N_12684,N_11887,N_12222);
nor U12685 (N_12685,N_11705,N_11961);
xor U12686 (N_12686,N_11558,N_12200);
xnor U12687 (N_12687,N_11814,N_11287);
xnor U12688 (N_12688,N_11915,N_11954);
and U12689 (N_12689,N_11566,N_12288);
or U12690 (N_12690,N_12418,N_11920);
xor U12691 (N_12691,N_12255,N_12019);
nor U12692 (N_12692,N_11746,N_12466);
or U12693 (N_12693,N_12102,N_11627);
or U12694 (N_12694,N_11310,N_11854);
xor U12695 (N_12695,N_11776,N_12049);
nor U12696 (N_12696,N_12205,N_12417);
xnor U12697 (N_12697,N_12199,N_11708);
and U12698 (N_12698,N_12313,N_11647);
nand U12699 (N_12699,N_12409,N_11773);
nand U12700 (N_12700,N_11937,N_11850);
or U12701 (N_12701,N_11290,N_12194);
xor U12702 (N_12702,N_11927,N_11859);
and U12703 (N_12703,N_12448,N_11428);
xnor U12704 (N_12704,N_11455,N_12385);
nand U12705 (N_12705,N_12227,N_12406);
nor U12706 (N_12706,N_12388,N_11879);
and U12707 (N_12707,N_12155,N_12185);
nor U12708 (N_12708,N_12411,N_11678);
or U12709 (N_12709,N_12241,N_11628);
or U12710 (N_12710,N_11935,N_12127);
or U12711 (N_12711,N_11600,N_11869);
and U12712 (N_12712,N_11488,N_11866);
nand U12713 (N_12713,N_12377,N_11907);
xnor U12714 (N_12714,N_12337,N_11404);
or U12715 (N_12715,N_11341,N_12156);
xor U12716 (N_12716,N_12054,N_12339);
and U12717 (N_12717,N_11534,N_12362);
nor U12718 (N_12718,N_12077,N_12195);
nand U12719 (N_12719,N_12381,N_11520);
and U12720 (N_12720,N_12196,N_11833);
nor U12721 (N_12721,N_12497,N_11973);
xor U12722 (N_12722,N_12214,N_11890);
nand U12723 (N_12723,N_11934,N_11521);
or U12724 (N_12724,N_11576,N_11893);
nor U12725 (N_12725,N_12447,N_12296);
nand U12726 (N_12726,N_12066,N_12478);
and U12727 (N_12727,N_11485,N_12016);
xor U12728 (N_12728,N_12424,N_12373);
nand U12729 (N_12729,N_11538,N_11586);
and U12730 (N_12730,N_12002,N_12164);
or U12731 (N_12731,N_11294,N_11641);
nand U12732 (N_12732,N_12450,N_12293);
or U12733 (N_12733,N_12175,N_12489);
or U12734 (N_12734,N_11965,N_11283);
nor U12735 (N_12735,N_11787,N_11840);
nand U12736 (N_12736,N_11998,N_11286);
nor U12737 (N_12737,N_11264,N_11530);
xor U12738 (N_12738,N_11322,N_12216);
nor U12739 (N_12739,N_11557,N_11815);
and U12740 (N_12740,N_12308,N_11364);
and U12741 (N_12741,N_11644,N_11783);
xor U12742 (N_12742,N_12242,N_12165);
nand U12743 (N_12743,N_12198,N_11498);
or U12744 (N_12744,N_11589,N_12304);
or U12745 (N_12745,N_12250,N_11366);
nand U12746 (N_12746,N_12336,N_12299);
or U12747 (N_12747,N_11813,N_11333);
nand U12748 (N_12748,N_12067,N_11896);
and U12749 (N_12749,N_11471,N_11824);
or U12750 (N_12750,N_12305,N_11443);
nand U12751 (N_12751,N_12268,N_12031);
and U12752 (N_12752,N_11976,N_11358);
xnor U12753 (N_12753,N_11539,N_11729);
xor U12754 (N_12754,N_12115,N_11506);
xnor U12755 (N_12755,N_12408,N_12474);
nor U12756 (N_12756,N_11681,N_11679);
xnor U12757 (N_12757,N_11981,N_11665);
and U12758 (N_12758,N_12298,N_11721);
and U12759 (N_12759,N_11860,N_12323);
and U12760 (N_12760,N_11779,N_12023);
and U12761 (N_12761,N_12369,N_11957);
or U12762 (N_12762,N_11552,N_11435);
and U12763 (N_12763,N_11345,N_12413);
and U12764 (N_12764,N_11962,N_12042);
and U12765 (N_12765,N_11759,N_11812);
or U12766 (N_12766,N_11385,N_12094);
and U12767 (N_12767,N_11434,N_11577);
xor U12768 (N_12768,N_12333,N_11995);
and U12769 (N_12769,N_12247,N_11261);
nand U12770 (N_12770,N_11795,N_11899);
and U12771 (N_12771,N_11414,N_11835);
nor U12772 (N_12772,N_12452,N_11282);
and U12773 (N_12773,N_12386,N_11592);
and U12774 (N_12774,N_12179,N_12343);
or U12775 (N_12775,N_12396,N_12446);
nand U12776 (N_12776,N_11281,N_12420);
xor U12777 (N_12777,N_11508,N_11612);
xor U12778 (N_12778,N_11582,N_11743);
or U12779 (N_12779,N_12024,N_11603);
nor U12780 (N_12780,N_11463,N_11784);
and U12781 (N_12781,N_11270,N_12081);
and U12782 (N_12782,N_12414,N_12279);
xor U12783 (N_12783,N_12093,N_11405);
nor U12784 (N_12784,N_11451,N_11673);
or U12785 (N_12785,N_12090,N_12402);
xor U12786 (N_12786,N_11692,N_11989);
xor U12787 (N_12787,N_11547,N_11517);
or U12788 (N_12788,N_11533,N_11472);
or U12789 (N_12789,N_11971,N_11950);
nand U12790 (N_12790,N_12248,N_12371);
xor U12791 (N_12791,N_12490,N_11769);
nor U12792 (N_12792,N_12213,N_11456);
or U12793 (N_12793,N_12462,N_11858);
nand U12794 (N_12794,N_12431,N_11910);
and U12795 (N_12795,N_11977,N_12273);
and U12796 (N_12796,N_11606,N_11426);
nor U12797 (N_12797,N_11953,N_11594);
xnor U12798 (N_12798,N_11767,N_11900);
nor U12799 (N_12799,N_11826,N_11599);
nand U12800 (N_12800,N_11919,N_11852);
nor U12801 (N_12801,N_11309,N_11367);
or U12802 (N_12802,N_12108,N_12262);
and U12803 (N_12803,N_11897,N_12217);
and U12804 (N_12804,N_12347,N_11313);
xor U12805 (N_12805,N_11510,N_12229);
xor U12806 (N_12806,N_11574,N_12189);
and U12807 (N_12807,N_11272,N_11470);
xnor U12808 (N_12808,N_12059,N_12340);
nand U12809 (N_12809,N_11768,N_12410);
nor U12810 (N_12810,N_11487,N_11390);
nor U12811 (N_12811,N_12130,N_11823);
nand U12812 (N_12812,N_12407,N_11605);
xnor U12813 (N_12813,N_11560,N_11822);
or U12814 (N_12814,N_12163,N_11693);
or U12815 (N_12815,N_11394,N_12283);
nor U12816 (N_12816,N_11970,N_11423);
xnor U12817 (N_12817,N_11601,N_12159);
nor U12818 (N_12818,N_11700,N_11597);
nand U12819 (N_12819,N_12206,N_11990);
nor U12820 (N_12820,N_11515,N_11349);
nand U12821 (N_12821,N_12387,N_11590);
xnor U12822 (N_12822,N_11639,N_11848);
or U12823 (N_12823,N_12209,N_11691);
and U12824 (N_12824,N_11300,N_11653);
nand U12825 (N_12825,N_12223,N_12171);
xnor U12826 (N_12826,N_11420,N_12232);
or U12827 (N_12827,N_12302,N_11454);
or U12828 (N_12828,N_11926,N_12312);
or U12829 (N_12829,N_12153,N_12261);
nand U12830 (N_12830,N_12129,N_11853);
xor U12831 (N_12831,N_11411,N_11735);
nand U12832 (N_12832,N_12495,N_12487);
or U12833 (N_12833,N_11765,N_11944);
or U12834 (N_12834,N_11278,N_12162);
nor U12835 (N_12835,N_12105,N_12072);
nor U12836 (N_12836,N_12496,N_12435);
and U12837 (N_12837,N_12338,N_11745);
and U12838 (N_12838,N_11509,N_12125);
or U12839 (N_12839,N_11785,N_11416);
and U12840 (N_12840,N_11573,N_11816);
nor U12841 (N_12841,N_11378,N_11450);
nor U12842 (N_12842,N_12244,N_12405);
nand U12843 (N_12843,N_11271,N_11634);
xor U12844 (N_12844,N_11338,N_11892);
nor U12845 (N_12845,N_12432,N_12368);
nor U12846 (N_12846,N_11924,N_11856);
or U12847 (N_12847,N_11916,N_12212);
nor U12848 (N_12848,N_12068,N_11452);
nand U12849 (N_12849,N_11645,N_11781);
or U12850 (N_12850,N_12172,N_12013);
nand U12851 (N_12851,N_11363,N_11625);
nand U12852 (N_12852,N_11786,N_11846);
nor U12853 (N_12853,N_11343,N_12135);
or U12854 (N_12854,N_12118,N_11381);
nand U12855 (N_12855,N_11389,N_11878);
xnor U12856 (N_12856,N_11803,N_12087);
nand U12857 (N_12857,N_11346,N_11862);
nand U12858 (N_12858,N_12291,N_11519);
nor U12859 (N_12859,N_12147,N_11516);
or U12860 (N_12860,N_11401,N_11331);
and U12861 (N_12861,N_11299,N_12186);
nor U12862 (N_12862,N_11662,N_11478);
or U12863 (N_12863,N_11365,N_11640);
xnor U12864 (N_12864,N_11752,N_12482);
xnor U12865 (N_12865,N_12326,N_11827);
nand U12866 (N_12866,N_12317,N_11825);
nor U12867 (N_12867,N_12139,N_11613);
or U12868 (N_12868,N_11838,N_11701);
xor U12869 (N_12869,N_11918,N_11888);
nand U12870 (N_12870,N_12355,N_12057);
xnor U12871 (N_12871,N_11368,N_11736);
nand U12872 (N_12872,N_11631,N_12300);
nor U12873 (N_12873,N_12275,N_11357);
xnor U12874 (N_12874,N_12348,N_11503);
nor U12875 (N_12875,N_11483,N_11388);
nor U12876 (N_12876,N_12439,N_11880);
xnor U12877 (N_12877,N_11324,N_11427);
or U12878 (N_12878,N_11609,N_11740);
nand U12879 (N_12879,N_12285,N_11499);
or U12880 (N_12880,N_11307,N_11579);
or U12881 (N_12881,N_11789,N_11289);
nand U12882 (N_12882,N_11325,N_11725);
xor U12883 (N_12883,N_11595,N_11355);
or U12884 (N_12884,N_12436,N_11458);
and U12885 (N_12885,N_11960,N_11811);
and U12886 (N_12886,N_12193,N_12297);
xor U12887 (N_12887,N_11475,N_11544);
and U12888 (N_12888,N_12065,N_11469);
nor U12889 (N_12889,N_11980,N_12342);
or U12890 (N_12890,N_12157,N_12101);
xnor U12891 (N_12891,N_12306,N_11298);
or U12892 (N_12892,N_11917,N_12236);
and U12893 (N_12893,N_11713,N_11477);
or U12894 (N_12894,N_11532,N_11491);
nor U12895 (N_12895,N_12041,N_11344);
nor U12896 (N_12896,N_11968,N_12136);
xnor U12897 (N_12897,N_11847,N_12047);
or U12898 (N_12898,N_12366,N_11474);
or U12899 (N_12899,N_11596,N_12378);
xor U12900 (N_12900,N_12085,N_11439);
xor U12901 (N_12901,N_12114,N_11462);
nor U12902 (N_12902,N_12176,N_11347);
and U12903 (N_12903,N_11429,N_12494);
and U12904 (N_12904,N_11291,N_12091);
xor U12905 (N_12905,N_12358,N_11668);
or U12906 (N_12906,N_11682,N_11712);
or U12907 (N_12907,N_12441,N_11315);
nand U12908 (N_12908,N_11535,N_11791);
and U12909 (N_12909,N_12419,N_12183);
or U12910 (N_12910,N_11938,N_11771);
or U12911 (N_12911,N_11350,N_11817);
or U12912 (N_12912,N_12464,N_11360);
nor U12913 (N_12913,N_12240,N_11622);
nand U12914 (N_12914,N_12036,N_11709);
xnor U12915 (N_12915,N_11905,N_11677);
nand U12916 (N_12916,N_11584,N_11277);
nand U12917 (N_12917,N_12238,N_11624);
nor U12918 (N_12918,N_12182,N_11956);
nor U12919 (N_12919,N_12480,N_11527);
xnor U12920 (N_12920,N_12140,N_11984);
and U12921 (N_12921,N_11946,N_11697);
xnor U12922 (N_12922,N_12361,N_11319);
nor U12923 (N_12923,N_12257,N_11799);
or U12924 (N_12924,N_11543,N_11632);
xor U12925 (N_12925,N_11482,N_11397);
and U12926 (N_12926,N_12226,N_11436);
and U12927 (N_12927,N_11901,N_12416);
nor U12928 (N_12928,N_11361,N_11722);
nor U12929 (N_12929,N_11440,N_11638);
and U12930 (N_12930,N_11790,N_11988);
nor U12931 (N_12931,N_12053,N_11540);
or U12932 (N_12932,N_12479,N_12170);
nor U12933 (N_12933,N_11380,N_11301);
nor U12934 (N_12934,N_11398,N_12303);
nor U12935 (N_12935,N_11461,N_12367);
or U12936 (N_12936,N_11849,N_12045);
and U12937 (N_12937,N_11621,N_12315);
and U12938 (N_12938,N_11306,N_12134);
nand U12939 (N_12939,N_11617,N_11553);
xnor U12940 (N_12940,N_11958,N_12295);
xor U12941 (N_12941,N_12403,N_12443);
or U12942 (N_12942,N_12335,N_12123);
or U12943 (N_12943,N_11667,N_11513);
xnor U12944 (N_12944,N_12460,N_12126);
xor U12945 (N_12945,N_11982,N_12039);
nor U12946 (N_12946,N_12389,N_12421);
nor U12947 (N_12947,N_11686,N_12266);
xor U12948 (N_12948,N_11320,N_11304);
and U12949 (N_12949,N_11861,N_11396);
nand U12950 (N_12950,N_12282,N_12307);
nand U12951 (N_12951,N_12384,N_11806);
nand U12952 (N_12952,N_12319,N_12451);
xor U12953 (N_12953,N_11774,N_11375);
nand U12954 (N_12954,N_11699,N_11758);
nand U12955 (N_12955,N_11909,N_12098);
xor U12956 (N_12956,N_11723,N_11720);
or U12957 (N_12957,N_12220,N_12399);
nor U12958 (N_12958,N_12109,N_12089);
xnor U12959 (N_12959,N_12056,N_12030);
nor U12960 (N_12960,N_12012,N_12400);
and U12961 (N_12961,N_11531,N_11754);
and U12962 (N_12962,N_12324,N_11941);
nor U12963 (N_12963,N_11656,N_11637);
xor U12964 (N_12964,N_11563,N_11542);
nor U12965 (N_12965,N_11254,N_11996);
or U12966 (N_12966,N_11794,N_11707);
xnor U12967 (N_12967,N_12160,N_11392);
or U12968 (N_12968,N_11546,N_12329);
nand U12969 (N_12969,N_12483,N_11568);
nand U12970 (N_12970,N_11536,N_11798);
nor U12971 (N_12971,N_11895,N_12492);
xnor U12972 (N_12972,N_11651,N_11425);
or U12973 (N_12973,N_11886,N_11353);
nor U12974 (N_12974,N_12096,N_11726);
nand U12975 (N_12975,N_11711,N_11408);
or U12976 (N_12976,N_11339,N_11549);
nand U12977 (N_12977,N_11493,N_11528);
nand U12978 (N_12978,N_11618,N_12245);
and U12979 (N_12979,N_11992,N_12456);
nor U12980 (N_12980,N_12256,N_11256);
or U12981 (N_12981,N_12481,N_11457);
and U12982 (N_12982,N_12174,N_11805);
and U12983 (N_12983,N_12393,N_11747);
xnor U12984 (N_12984,N_11602,N_12423);
or U12985 (N_12985,N_12145,N_11867);
and U12986 (N_12986,N_11898,N_12277);
xnor U12987 (N_12987,N_12415,N_11873);
and U12988 (N_12988,N_12243,N_12457);
nand U12989 (N_12989,N_11882,N_11399);
xnor U12990 (N_12990,N_11979,N_11780);
and U12991 (N_12991,N_11994,N_11845);
nor U12992 (N_12992,N_11804,N_11556);
nand U12993 (N_12993,N_11680,N_11629);
xor U12994 (N_12994,N_11670,N_11633);
xor U12995 (N_12995,N_12332,N_11391);
or U12996 (N_12996,N_11727,N_12425);
xnor U12997 (N_12997,N_12011,N_12017);
and U12998 (N_12998,N_11831,N_12070);
or U12999 (N_12999,N_12449,N_11585);
xnor U13000 (N_13000,N_11587,N_11870);
xor U13001 (N_13001,N_11718,N_12150);
or U13002 (N_13002,N_11424,N_11772);
and U13003 (N_13003,N_11753,N_11969);
nor U13004 (N_13004,N_12433,N_12422);
xor U13005 (N_13005,N_12061,N_12154);
nand U13006 (N_13006,N_11657,N_11410);
nand U13007 (N_13007,N_11658,N_12032);
nand U13008 (N_13008,N_12318,N_12276);
nor U13009 (N_13009,N_12440,N_11741);
nand U13010 (N_13010,N_11744,N_12314);
xor U13011 (N_13011,N_12331,N_11777);
nand U13012 (N_13012,N_12063,N_12188);
xnor U13013 (N_13013,N_12148,N_12055);
xnor U13014 (N_13014,N_12076,N_12473);
nand U13015 (N_13015,N_11529,N_11797);
nor U13016 (N_13016,N_11913,N_12363);
nor U13017 (N_13017,N_11710,N_11788);
xor U13018 (N_13018,N_11302,N_12471);
and U13019 (N_13019,N_11459,N_11373);
nand U13020 (N_13020,N_11951,N_11750);
or U13021 (N_13021,N_11874,N_11734);
or U13022 (N_13022,N_11646,N_11481);
nor U13023 (N_13023,N_11688,N_12173);
or U13024 (N_13024,N_12364,N_11492);
and U13025 (N_13025,N_12116,N_12341);
or U13026 (N_13026,N_11702,N_11561);
and U13027 (N_13027,N_11802,N_12027);
nor U13028 (N_13028,N_12097,N_11312);
or U13029 (N_13029,N_11311,N_11438);
nor U13030 (N_13030,N_11327,N_12103);
xor U13031 (N_13031,N_11496,N_12052);
and U13032 (N_13032,N_11260,N_11252);
nand U13033 (N_13033,N_11660,N_12035);
or U13034 (N_13034,N_12476,N_12351);
nand U13035 (N_13035,N_12251,N_11296);
or U13036 (N_13036,N_11308,N_12202);
or U13037 (N_13037,N_12117,N_12477);
and U13038 (N_13038,N_12395,N_11421);
xor U13039 (N_13039,N_12084,N_11978);
nor U13040 (N_13040,N_11936,N_11253);
nand U13041 (N_13041,N_12215,N_11251);
and U13042 (N_13042,N_11468,N_12168);
nand U13043 (N_13043,N_12454,N_12491);
and U13044 (N_13044,N_11775,N_12106);
or U13045 (N_13045,N_11821,N_11608);
and U13046 (N_13046,N_12037,N_11930);
and U13047 (N_13047,N_11329,N_11342);
nor U13048 (N_13048,N_12086,N_12137);
nor U13049 (N_13049,N_11545,N_12071);
nand U13050 (N_13050,N_12203,N_11466);
or U13051 (N_13051,N_12119,N_11952);
xor U13052 (N_13052,N_11733,N_11928);
nor U13053 (N_13053,N_12485,N_12021);
and U13054 (N_13054,N_11569,N_12429);
nand U13055 (N_13055,N_11554,N_12263);
and U13056 (N_13056,N_12111,N_12311);
xnor U13057 (N_13057,N_12427,N_11939);
nand U13058 (N_13058,N_11490,N_11502);
nor U13059 (N_13059,N_12149,N_12272);
and U13060 (N_13060,N_12286,N_11921);
nor U13061 (N_13061,N_12346,N_11376);
or U13062 (N_13062,N_12219,N_11562);
nor U13063 (N_13063,N_11407,N_11442);
xor U13064 (N_13064,N_12401,N_11630);
or U13065 (N_13065,N_11820,N_12394);
nor U13066 (N_13066,N_12143,N_11395);
xnor U13067 (N_13067,N_11284,N_11732);
nand U13068 (N_13068,N_12218,N_12201);
and U13069 (N_13069,N_12375,N_11863);
or U13070 (N_13070,N_11843,N_12008);
or U13071 (N_13071,N_12152,N_11891);
nand U13072 (N_13072,N_11664,N_12083);
and U13073 (N_13073,N_12334,N_12184);
nand U13074 (N_13074,N_11809,N_12038);
and U13075 (N_13075,N_12391,N_11580);
and U13076 (N_13076,N_11273,N_12289);
or U13077 (N_13077,N_12112,N_12374);
nor U13078 (N_13078,N_11285,N_12264);
nand U13079 (N_13079,N_12132,N_12161);
or U13080 (N_13080,N_11942,N_11731);
or U13081 (N_13081,N_11684,N_11974);
or U13082 (N_13082,N_12058,N_11340);
or U13083 (N_13083,N_12088,N_12234);
and U13084 (N_13084,N_11518,N_11318);
and U13085 (N_13085,N_12258,N_12472);
xor U13086 (N_13086,N_12246,N_11565);
and U13087 (N_13087,N_12001,N_11337);
xnor U13088 (N_13088,N_12453,N_11588);
or U13089 (N_13089,N_12379,N_11931);
or U13090 (N_13090,N_12142,N_11755);
nand U13091 (N_13091,N_11675,N_12034);
nor U13092 (N_13092,N_12239,N_11473);
nor U13093 (N_13093,N_11757,N_12131);
or U13094 (N_13094,N_11446,N_11674);
and U13095 (N_13095,N_11372,N_11382);
nand U13096 (N_13096,N_11703,N_11571);
nand U13097 (N_13097,N_11620,N_11908);
and U13098 (N_13098,N_11572,N_12062);
and U13099 (N_13099,N_12383,N_11614);
nor U13100 (N_13100,N_12120,N_12110);
xnor U13101 (N_13101,N_11548,N_11922);
and U13102 (N_13102,N_12046,N_11352);
nand U13103 (N_13103,N_11881,N_11444);
nand U13104 (N_13104,N_12128,N_11694);
and U13105 (N_13105,N_12353,N_12437);
nand U13106 (N_13106,N_11541,N_11875);
nand U13107 (N_13107,N_12350,N_11698);
xor U13108 (N_13108,N_12051,N_11460);
or U13109 (N_13109,N_11348,N_11690);
nand U13110 (N_13110,N_11829,N_11403);
or U13111 (N_13111,N_11359,N_11964);
and U13112 (N_13112,N_12271,N_11739);
and U13113 (N_13113,N_11292,N_11288);
nor U13114 (N_13114,N_12438,N_11719);
xnor U13115 (N_13115,N_11695,N_12224);
nand U13116 (N_13116,N_11486,N_11615);
nor U13117 (N_13117,N_12380,N_11883);
and U13118 (N_13118,N_11762,N_11370);
nor U13119 (N_13119,N_11334,N_11578);
and U13120 (N_13120,N_11635,N_11871);
or U13121 (N_13121,N_12025,N_11354);
nand U13122 (N_13122,N_11504,N_11728);
and U13123 (N_13123,N_12265,N_12121);
nor U13124 (N_13124,N_12166,N_12079);
nand U13125 (N_13125,N_12411,N_12380);
xor U13126 (N_13126,N_11793,N_11494);
and U13127 (N_13127,N_11440,N_12245);
nand U13128 (N_13128,N_11855,N_11352);
xnor U13129 (N_13129,N_11669,N_11404);
nand U13130 (N_13130,N_11841,N_12122);
nand U13131 (N_13131,N_11707,N_11893);
or U13132 (N_13132,N_11970,N_12358);
xor U13133 (N_13133,N_11454,N_11866);
and U13134 (N_13134,N_12499,N_12173);
or U13135 (N_13135,N_12156,N_11604);
nand U13136 (N_13136,N_12171,N_11414);
or U13137 (N_13137,N_11825,N_12045);
or U13138 (N_13138,N_11815,N_11579);
xor U13139 (N_13139,N_11494,N_12258);
or U13140 (N_13140,N_11771,N_11862);
nand U13141 (N_13141,N_12398,N_11723);
nand U13142 (N_13142,N_11633,N_12293);
or U13143 (N_13143,N_11404,N_11447);
and U13144 (N_13144,N_12300,N_11387);
nor U13145 (N_13145,N_12106,N_12249);
nor U13146 (N_13146,N_11286,N_12444);
or U13147 (N_13147,N_11525,N_11514);
xor U13148 (N_13148,N_12125,N_12213);
and U13149 (N_13149,N_11552,N_11363);
nand U13150 (N_13150,N_11677,N_11734);
and U13151 (N_13151,N_12002,N_11309);
or U13152 (N_13152,N_11489,N_12128);
nand U13153 (N_13153,N_12216,N_12172);
xnor U13154 (N_13154,N_11981,N_11276);
nor U13155 (N_13155,N_12466,N_11803);
and U13156 (N_13156,N_11297,N_12305);
xor U13157 (N_13157,N_11730,N_11880);
and U13158 (N_13158,N_12374,N_11968);
xor U13159 (N_13159,N_11531,N_11386);
xnor U13160 (N_13160,N_11400,N_11765);
xnor U13161 (N_13161,N_12136,N_11310);
xor U13162 (N_13162,N_11455,N_11353);
and U13163 (N_13163,N_11888,N_11295);
xor U13164 (N_13164,N_11949,N_11382);
xnor U13165 (N_13165,N_12378,N_11910);
nand U13166 (N_13166,N_12166,N_11341);
nor U13167 (N_13167,N_11625,N_12452);
and U13168 (N_13168,N_12131,N_12202);
or U13169 (N_13169,N_12462,N_12168);
xor U13170 (N_13170,N_11953,N_11326);
or U13171 (N_13171,N_11323,N_12059);
or U13172 (N_13172,N_11416,N_11274);
xor U13173 (N_13173,N_11365,N_11571);
or U13174 (N_13174,N_12348,N_12472);
and U13175 (N_13175,N_12432,N_11403);
or U13176 (N_13176,N_11547,N_11393);
nand U13177 (N_13177,N_12110,N_12202);
nor U13178 (N_13178,N_12357,N_12138);
or U13179 (N_13179,N_11916,N_11504);
nand U13180 (N_13180,N_11534,N_12149);
and U13181 (N_13181,N_12122,N_11283);
xnor U13182 (N_13182,N_12246,N_12138);
nand U13183 (N_13183,N_12406,N_11836);
and U13184 (N_13184,N_11643,N_11658);
nor U13185 (N_13185,N_11314,N_11875);
xor U13186 (N_13186,N_11463,N_11289);
nor U13187 (N_13187,N_12378,N_11786);
xnor U13188 (N_13188,N_11291,N_11579);
nor U13189 (N_13189,N_11493,N_11375);
nor U13190 (N_13190,N_12469,N_12223);
or U13191 (N_13191,N_11712,N_12017);
nor U13192 (N_13192,N_11979,N_12222);
and U13193 (N_13193,N_12143,N_11785);
nand U13194 (N_13194,N_11873,N_12087);
nand U13195 (N_13195,N_12343,N_11303);
or U13196 (N_13196,N_11708,N_12300);
or U13197 (N_13197,N_12171,N_11563);
or U13198 (N_13198,N_12370,N_11541);
nand U13199 (N_13199,N_11627,N_12230);
nor U13200 (N_13200,N_12423,N_11453);
nor U13201 (N_13201,N_12146,N_12316);
nor U13202 (N_13202,N_12301,N_11421);
xor U13203 (N_13203,N_11973,N_11943);
nand U13204 (N_13204,N_11725,N_11558);
or U13205 (N_13205,N_12302,N_11281);
and U13206 (N_13206,N_11641,N_11429);
or U13207 (N_13207,N_11800,N_12193);
nand U13208 (N_13208,N_11595,N_12331);
nand U13209 (N_13209,N_11571,N_12067);
or U13210 (N_13210,N_11824,N_12368);
or U13211 (N_13211,N_11311,N_11760);
or U13212 (N_13212,N_11694,N_11899);
nand U13213 (N_13213,N_11267,N_12210);
and U13214 (N_13214,N_11597,N_11583);
and U13215 (N_13215,N_11554,N_12411);
nor U13216 (N_13216,N_12352,N_11509);
nand U13217 (N_13217,N_12116,N_12181);
xor U13218 (N_13218,N_12318,N_11922);
xor U13219 (N_13219,N_11292,N_12455);
and U13220 (N_13220,N_11630,N_12255);
xnor U13221 (N_13221,N_11932,N_11496);
and U13222 (N_13222,N_12167,N_12016);
nor U13223 (N_13223,N_12496,N_11395);
and U13224 (N_13224,N_11878,N_12310);
or U13225 (N_13225,N_12064,N_12412);
or U13226 (N_13226,N_12128,N_12266);
xnor U13227 (N_13227,N_11860,N_11561);
or U13228 (N_13228,N_11393,N_11503);
nand U13229 (N_13229,N_11355,N_11673);
and U13230 (N_13230,N_11339,N_11787);
nor U13231 (N_13231,N_12494,N_11377);
nor U13232 (N_13232,N_11556,N_11368);
xor U13233 (N_13233,N_12403,N_11916);
nor U13234 (N_13234,N_11418,N_11741);
nand U13235 (N_13235,N_11257,N_11999);
and U13236 (N_13236,N_12436,N_11945);
xor U13237 (N_13237,N_11428,N_11485);
nor U13238 (N_13238,N_12376,N_12129);
xor U13239 (N_13239,N_12492,N_12359);
nand U13240 (N_13240,N_11550,N_11728);
nand U13241 (N_13241,N_12275,N_11690);
nand U13242 (N_13242,N_11316,N_12241);
and U13243 (N_13243,N_11408,N_12366);
xor U13244 (N_13244,N_12247,N_12091);
or U13245 (N_13245,N_12434,N_12111);
nand U13246 (N_13246,N_11515,N_12039);
nor U13247 (N_13247,N_12215,N_12126);
or U13248 (N_13248,N_11517,N_11919);
or U13249 (N_13249,N_11954,N_12097);
xor U13250 (N_13250,N_12008,N_11749);
nand U13251 (N_13251,N_11405,N_11797);
xnor U13252 (N_13252,N_12060,N_12181);
or U13253 (N_13253,N_12215,N_12453);
or U13254 (N_13254,N_12451,N_11308);
nor U13255 (N_13255,N_11291,N_11447);
xnor U13256 (N_13256,N_11620,N_12401);
or U13257 (N_13257,N_11402,N_11650);
nand U13258 (N_13258,N_11837,N_11927);
or U13259 (N_13259,N_12021,N_12213);
and U13260 (N_13260,N_12200,N_11911);
xor U13261 (N_13261,N_12435,N_11304);
xor U13262 (N_13262,N_11689,N_11352);
and U13263 (N_13263,N_11537,N_11944);
or U13264 (N_13264,N_11552,N_11871);
nor U13265 (N_13265,N_11259,N_11638);
and U13266 (N_13266,N_11599,N_11431);
nand U13267 (N_13267,N_12294,N_11602);
nand U13268 (N_13268,N_11903,N_11931);
nor U13269 (N_13269,N_11583,N_11352);
xnor U13270 (N_13270,N_11308,N_12164);
or U13271 (N_13271,N_11569,N_12189);
nand U13272 (N_13272,N_12347,N_11999);
or U13273 (N_13273,N_11486,N_11389);
xor U13274 (N_13274,N_12076,N_11954);
nor U13275 (N_13275,N_12067,N_11835);
xor U13276 (N_13276,N_11859,N_12248);
nor U13277 (N_13277,N_11325,N_11473);
xnor U13278 (N_13278,N_11967,N_11705);
nor U13279 (N_13279,N_11466,N_11901);
nand U13280 (N_13280,N_11702,N_11318);
or U13281 (N_13281,N_11655,N_12109);
xor U13282 (N_13282,N_12436,N_11578);
or U13283 (N_13283,N_11321,N_12144);
nand U13284 (N_13284,N_11965,N_12446);
and U13285 (N_13285,N_11979,N_11935);
or U13286 (N_13286,N_11955,N_11381);
nand U13287 (N_13287,N_11799,N_12231);
or U13288 (N_13288,N_12371,N_11852);
and U13289 (N_13289,N_11749,N_11409);
xor U13290 (N_13290,N_12166,N_12424);
nand U13291 (N_13291,N_11712,N_11838);
or U13292 (N_13292,N_11536,N_11335);
nor U13293 (N_13293,N_11769,N_12082);
and U13294 (N_13294,N_11686,N_12432);
or U13295 (N_13295,N_12394,N_12380);
or U13296 (N_13296,N_12031,N_12196);
nand U13297 (N_13297,N_11794,N_11291);
nand U13298 (N_13298,N_11615,N_11374);
nor U13299 (N_13299,N_12276,N_12372);
nor U13300 (N_13300,N_11943,N_11540);
nand U13301 (N_13301,N_12175,N_12479);
and U13302 (N_13302,N_11814,N_11350);
xnor U13303 (N_13303,N_11904,N_11374);
nand U13304 (N_13304,N_11860,N_11514);
xor U13305 (N_13305,N_11794,N_11523);
or U13306 (N_13306,N_12095,N_11306);
nand U13307 (N_13307,N_12236,N_11529);
nand U13308 (N_13308,N_12480,N_11325);
and U13309 (N_13309,N_11800,N_11843);
or U13310 (N_13310,N_12219,N_11494);
xnor U13311 (N_13311,N_12101,N_12295);
nor U13312 (N_13312,N_11673,N_12284);
and U13313 (N_13313,N_12285,N_12216);
xnor U13314 (N_13314,N_11709,N_12084);
and U13315 (N_13315,N_11950,N_11709);
nand U13316 (N_13316,N_12246,N_11707);
or U13317 (N_13317,N_12044,N_11869);
xor U13318 (N_13318,N_11346,N_11719);
and U13319 (N_13319,N_11598,N_12130);
and U13320 (N_13320,N_11647,N_12305);
xnor U13321 (N_13321,N_12317,N_11307);
nor U13322 (N_13322,N_11418,N_11422);
nor U13323 (N_13323,N_11904,N_11576);
nand U13324 (N_13324,N_12402,N_11899);
or U13325 (N_13325,N_12243,N_12207);
xor U13326 (N_13326,N_12180,N_12057);
or U13327 (N_13327,N_11408,N_11933);
nor U13328 (N_13328,N_11984,N_11949);
nand U13329 (N_13329,N_11500,N_11335);
and U13330 (N_13330,N_11979,N_12149);
or U13331 (N_13331,N_11342,N_12450);
or U13332 (N_13332,N_12068,N_12454);
or U13333 (N_13333,N_11827,N_11396);
nand U13334 (N_13334,N_11549,N_12367);
nor U13335 (N_13335,N_11800,N_11945);
and U13336 (N_13336,N_11353,N_11838);
nor U13337 (N_13337,N_12465,N_11991);
xnor U13338 (N_13338,N_11470,N_12258);
nand U13339 (N_13339,N_11727,N_11400);
and U13340 (N_13340,N_11756,N_11604);
and U13341 (N_13341,N_12300,N_11913);
nor U13342 (N_13342,N_11760,N_12001);
or U13343 (N_13343,N_12053,N_12101);
or U13344 (N_13344,N_12406,N_11381);
nand U13345 (N_13345,N_11712,N_11427);
or U13346 (N_13346,N_12337,N_12341);
xor U13347 (N_13347,N_11953,N_11404);
or U13348 (N_13348,N_12499,N_11805);
nor U13349 (N_13349,N_11256,N_11621);
xor U13350 (N_13350,N_12499,N_12120);
xor U13351 (N_13351,N_11882,N_11878);
nand U13352 (N_13352,N_11284,N_11907);
or U13353 (N_13353,N_11357,N_11602);
xnor U13354 (N_13354,N_11567,N_12369);
and U13355 (N_13355,N_11542,N_12256);
xor U13356 (N_13356,N_11838,N_12315);
xnor U13357 (N_13357,N_12258,N_12309);
nand U13358 (N_13358,N_12295,N_11311);
and U13359 (N_13359,N_11371,N_11343);
and U13360 (N_13360,N_12101,N_11492);
xnor U13361 (N_13361,N_12237,N_11944);
and U13362 (N_13362,N_12141,N_11926);
nand U13363 (N_13363,N_12447,N_11981);
and U13364 (N_13364,N_11801,N_12237);
xor U13365 (N_13365,N_11574,N_11355);
nor U13366 (N_13366,N_11594,N_11706);
or U13367 (N_13367,N_11790,N_12045);
nor U13368 (N_13368,N_11282,N_11886);
xnor U13369 (N_13369,N_12075,N_11674);
nor U13370 (N_13370,N_11499,N_11265);
nand U13371 (N_13371,N_11852,N_11830);
or U13372 (N_13372,N_12305,N_11680);
and U13373 (N_13373,N_11773,N_11572);
nand U13374 (N_13374,N_11251,N_11698);
nor U13375 (N_13375,N_12033,N_11795);
nand U13376 (N_13376,N_12143,N_12116);
nand U13377 (N_13377,N_11519,N_12304);
nand U13378 (N_13378,N_11693,N_12448);
or U13379 (N_13379,N_12097,N_11637);
nor U13380 (N_13380,N_12292,N_12370);
nand U13381 (N_13381,N_11303,N_11607);
nor U13382 (N_13382,N_11791,N_12219);
nand U13383 (N_13383,N_12085,N_12340);
nand U13384 (N_13384,N_12214,N_11915);
or U13385 (N_13385,N_12155,N_11715);
nor U13386 (N_13386,N_12302,N_11973);
nand U13387 (N_13387,N_11943,N_11645);
nor U13388 (N_13388,N_12115,N_11573);
and U13389 (N_13389,N_11303,N_12218);
xor U13390 (N_13390,N_11830,N_11427);
nand U13391 (N_13391,N_12425,N_11282);
or U13392 (N_13392,N_11640,N_11881);
nand U13393 (N_13393,N_12297,N_11741);
xnor U13394 (N_13394,N_11813,N_11698);
nor U13395 (N_13395,N_11959,N_12281);
and U13396 (N_13396,N_12096,N_12019);
or U13397 (N_13397,N_11558,N_11276);
nor U13398 (N_13398,N_12309,N_11571);
nor U13399 (N_13399,N_12376,N_11961);
xor U13400 (N_13400,N_11785,N_12470);
or U13401 (N_13401,N_11577,N_12037);
nor U13402 (N_13402,N_12263,N_11790);
nand U13403 (N_13403,N_11317,N_12464);
xnor U13404 (N_13404,N_11958,N_11907);
xnor U13405 (N_13405,N_12033,N_11773);
xor U13406 (N_13406,N_12461,N_11739);
and U13407 (N_13407,N_11251,N_11657);
nand U13408 (N_13408,N_12077,N_12471);
nor U13409 (N_13409,N_11876,N_11849);
xor U13410 (N_13410,N_12420,N_12229);
nor U13411 (N_13411,N_11339,N_11873);
and U13412 (N_13412,N_11467,N_12122);
nand U13413 (N_13413,N_12249,N_11847);
or U13414 (N_13414,N_11995,N_11414);
nor U13415 (N_13415,N_11324,N_11764);
or U13416 (N_13416,N_11384,N_11280);
or U13417 (N_13417,N_11680,N_11834);
xnor U13418 (N_13418,N_12220,N_11605);
xnor U13419 (N_13419,N_11823,N_11322);
xnor U13420 (N_13420,N_11384,N_12480);
xor U13421 (N_13421,N_11997,N_12409);
or U13422 (N_13422,N_11898,N_11589);
xor U13423 (N_13423,N_12344,N_12309);
xnor U13424 (N_13424,N_11400,N_12342);
or U13425 (N_13425,N_11839,N_12471);
or U13426 (N_13426,N_11403,N_12022);
nand U13427 (N_13427,N_11748,N_11573);
nor U13428 (N_13428,N_12363,N_11370);
or U13429 (N_13429,N_12082,N_12063);
nand U13430 (N_13430,N_12386,N_12098);
nor U13431 (N_13431,N_12156,N_12039);
nor U13432 (N_13432,N_12409,N_12135);
and U13433 (N_13433,N_12368,N_12090);
xor U13434 (N_13434,N_12123,N_11445);
xnor U13435 (N_13435,N_11314,N_12418);
and U13436 (N_13436,N_11345,N_11957);
nand U13437 (N_13437,N_11418,N_12153);
and U13438 (N_13438,N_12426,N_11613);
xnor U13439 (N_13439,N_11887,N_11372);
nand U13440 (N_13440,N_11425,N_11575);
and U13441 (N_13441,N_12205,N_12408);
or U13442 (N_13442,N_11810,N_12134);
nand U13443 (N_13443,N_12353,N_11678);
nor U13444 (N_13444,N_11933,N_12386);
nor U13445 (N_13445,N_11640,N_11868);
and U13446 (N_13446,N_12100,N_11968);
nor U13447 (N_13447,N_11375,N_11630);
nor U13448 (N_13448,N_11362,N_11366);
or U13449 (N_13449,N_11623,N_12076);
nand U13450 (N_13450,N_12134,N_11737);
nand U13451 (N_13451,N_11814,N_11942);
nand U13452 (N_13452,N_12181,N_11471);
nand U13453 (N_13453,N_11251,N_11705);
nor U13454 (N_13454,N_11958,N_11300);
nand U13455 (N_13455,N_11459,N_11771);
nand U13456 (N_13456,N_12092,N_11473);
or U13457 (N_13457,N_11938,N_11966);
nor U13458 (N_13458,N_12176,N_11392);
or U13459 (N_13459,N_12188,N_11680);
xor U13460 (N_13460,N_11861,N_12367);
or U13461 (N_13461,N_11411,N_12065);
xnor U13462 (N_13462,N_11810,N_11323);
and U13463 (N_13463,N_11309,N_12125);
xor U13464 (N_13464,N_11538,N_11759);
xor U13465 (N_13465,N_11317,N_12126);
and U13466 (N_13466,N_11304,N_12382);
nor U13467 (N_13467,N_11550,N_12112);
or U13468 (N_13468,N_12046,N_12190);
xor U13469 (N_13469,N_12002,N_12134);
nand U13470 (N_13470,N_11786,N_11896);
xor U13471 (N_13471,N_12400,N_11580);
nand U13472 (N_13472,N_12287,N_11696);
xor U13473 (N_13473,N_12356,N_12086);
xor U13474 (N_13474,N_12398,N_11323);
xor U13475 (N_13475,N_11441,N_11744);
xnor U13476 (N_13476,N_12139,N_11445);
nor U13477 (N_13477,N_11265,N_12187);
nand U13478 (N_13478,N_12354,N_11888);
or U13479 (N_13479,N_11944,N_12346);
nor U13480 (N_13480,N_11591,N_12490);
and U13481 (N_13481,N_11986,N_11281);
or U13482 (N_13482,N_11644,N_12059);
xor U13483 (N_13483,N_11406,N_12446);
nand U13484 (N_13484,N_11873,N_11315);
nand U13485 (N_13485,N_11449,N_12340);
nor U13486 (N_13486,N_11766,N_11547);
nor U13487 (N_13487,N_12188,N_12008);
xnor U13488 (N_13488,N_12047,N_11581);
and U13489 (N_13489,N_11531,N_11944);
nor U13490 (N_13490,N_11281,N_12188);
and U13491 (N_13491,N_11349,N_12032);
xnor U13492 (N_13492,N_12046,N_11999);
xnor U13493 (N_13493,N_11307,N_11922);
or U13494 (N_13494,N_11923,N_12196);
nand U13495 (N_13495,N_12191,N_12049);
or U13496 (N_13496,N_11872,N_12350);
or U13497 (N_13497,N_11277,N_12207);
nand U13498 (N_13498,N_12273,N_11985);
xor U13499 (N_13499,N_11884,N_11951);
nor U13500 (N_13500,N_12465,N_11637);
or U13501 (N_13501,N_12095,N_12307);
nand U13502 (N_13502,N_11568,N_11591);
xnor U13503 (N_13503,N_11586,N_12303);
xnor U13504 (N_13504,N_11551,N_11628);
nand U13505 (N_13505,N_11586,N_11753);
nor U13506 (N_13506,N_12446,N_11476);
and U13507 (N_13507,N_12280,N_11545);
or U13508 (N_13508,N_12239,N_11310);
xor U13509 (N_13509,N_11797,N_12477);
or U13510 (N_13510,N_11667,N_11906);
nor U13511 (N_13511,N_12483,N_12188);
and U13512 (N_13512,N_12355,N_12309);
xnor U13513 (N_13513,N_11594,N_11397);
or U13514 (N_13514,N_11767,N_11442);
or U13515 (N_13515,N_11450,N_11411);
or U13516 (N_13516,N_11525,N_11818);
nand U13517 (N_13517,N_12495,N_11832);
xor U13518 (N_13518,N_12094,N_11932);
xor U13519 (N_13519,N_11722,N_12340);
nand U13520 (N_13520,N_12093,N_11386);
nand U13521 (N_13521,N_11755,N_11988);
or U13522 (N_13522,N_11700,N_11464);
nor U13523 (N_13523,N_12175,N_11609);
nor U13524 (N_13524,N_11250,N_11446);
and U13525 (N_13525,N_11784,N_11250);
or U13526 (N_13526,N_11642,N_11939);
nor U13527 (N_13527,N_12269,N_11606);
nand U13528 (N_13528,N_11838,N_12077);
or U13529 (N_13529,N_11592,N_11341);
nand U13530 (N_13530,N_11300,N_11485);
nand U13531 (N_13531,N_12186,N_11988);
nor U13532 (N_13532,N_12085,N_12284);
nand U13533 (N_13533,N_11898,N_11971);
nor U13534 (N_13534,N_11703,N_11970);
and U13535 (N_13535,N_11342,N_11378);
xor U13536 (N_13536,N_12164,N_12416);
xnor U13537 (N_13537,N_12417,N_11468);
nand U13538 (N_13538,N_11501,N_11639);
or U13539 (N_13539,N_11880,N_11254);
nor U13540 (N_13540,N_11687,N_11752);
xor U13541 (N_13541,N_11554,N_11611);
or U13542 (N_13542,N_12299,N_11331);
and U13543 (N_13543,N_12037,N_11479);
xor U13544 (N_13544,N_12238,N_11430);
and U13545 (N_13545,N_11696,N_11733);
and U13546 (N_13546,N_12364,N_11784);
nor U13547 (N_13547,N_12058,N_12065);
xnor U13548 (N_13548,N_12371,N_11683);
and U13549 (N_13549,N_11613,N_11419);
nand U13550 (N_13550,N_11410,N_11792);
nor U13551 (N_13551,N_11624,N_11808);
and U13552 (N_13552,N_11415,N_12070);
and U13553 (N_13553,N_11774,N_11582);
nor U13554 (N_13554,N_12378,N_12266);
xor U13555 (N_13555,N_12038,N_12019);
xor U13556 (N_13556,N_11613,N_11546);
or U13557 (N_13557,N_11286,N_12215);
or U13558 (N_13558,N_11437,N_11422);
nand U13559 (N_13559,N_11479,N_12150);
or U13560 (N_13560,N_12289,N_11418);
and U13561 (N_13561,N_11845,N_11766);
or U13562 (N_13562,N_12081,N_12385);
nor U13563 (N_13563,N_11628,N_11489);
nor U13564 (N_13564,N_11631,N_11953);
xnor U13565 (N_13565,N_11923,N_12136);
xnor U13566 (N_13566,N_12044,N_11847);
xor U13567 (N_13567,N_11959,N_12080);
nor U13568 (N_13568,N_12118,N_11848);
nor U13569 (N_13569,N_12025,N_12012);
or U13570 (N_13570,N_11374,N_11935);
and U13571 (N_13571,N_12267,N_12260);
nor U13572 (N_13572,N_12319,N_12412);
nand U13573 (N_13573,N_12224,N_11982);
nor U13574 (N_13574,N_12442,N_11970);
or U13575 (N_13575,N_11337,N_11989);
or U13576 (N_13576,N_12423,N_11979);
nand U13577 (N_13577,N_12430,N_11533);
nor U13578 (N_13578,N_11354,N_12220);
and U13579 (N_13579,N_12382,N_12330);
xnor U13580 (N_13580,N_12291,N_11774);
xor U13581 (N_13581,N_11672,N_12311);
and U13582 (N_13582,N_12028,N_11679);
or U13583 (N_13583,N_12243,N_12399);
xnor U13584 (N_13584,N_11790,N_11776);
nor U13585 (N_13585,N_12201,N_11887);
nand U13586 (N_13586,N_11716,N_11484);
and U13587 (N_13587,N_11603,N_11902);
and U13588 (N_13588,N_11862,N_11837);
and U13589 (N_13589,N_11783,N_12427);
or U13590 (N_13590,N_11586,N_12061);
nor U13591 (N_13591,N_11886,N_11762);
nand U13592 (N_13592,N_11521,N_11915);
nor U13593 (N_13593,N_11619,N_11750);
or U13594 (N_13594,N_11515,N_11519);
xor U13595 (N_13595,N_12116,N_11370);
xnor U13596 (N_13596,N_11390,N_11617);
nor U13597 (N_13597,N_11284,N_11259);
and U13598 (N_13598,N_11596,N_11557);
nand U13599 (N_13599,N_12366,N_11459);
or U13600 (N_13600,N_11334,N_12414);
and U13601 (N_13601,N_11395,N_11687);
xnor U13602 (N_13602,N_11924,N_11761);
and U13603 (N_13603,N_12241,N_11496);
nor U13604 (N_13604,N_11814,N_11408);
nand U13605 (N_13605,N_11283,N_12239);
nand U13606 (N_13606,N_11366,N_12376);
nand U13607 (N_13607,N_12498,N_11960);
xor U13608 (N_13608,N_12214,N_12044);
and U13609 (N_13609,N_12465,N_11860);
xor U13610 (N_13610,N_12410,N_12428);
nor U13611 (N_13611,N_12020,N_11274);
and U13612 (N_13612,N_11936,N_12059);
xor U13613 (N_13613,N_11828,N_12205);
nand U13614 (N_13614,N_11612,N_12356);
and U13615 (N_13615,N_12476,N_12103);
xnor U13616 (N_13616,N_11753,N_11467);
xor U13617 (N_13617,N_11319,N_11992);
xor U13618 (N_13618,N_12231,N_11470);
or U13619 (N_13619,N_12324,N_11463);
xor U13620 (N_13620,N_11303,N_12181);
xnor U13621 (N_13621,N_11353,N_12417);
and U13622 (N_13622,N_11288,N_11713);
and U13623 (N_13623,N_11758,N_11724);
xnor U13624 (N_13624,N_12150,N_11614);
nand U13625 (N_13625,N_11894,N_12170);
and U13626 (N_13626,N_12204,N_11309);
and U13627 (N_13627,N_12017,N_11568);
nor U13628 (N_13628,N_11832,N_11337);
and U13629 (N_13629,N_11869,N_11644);
xnor U13630 (N_13630,N_11402,N_12243);
and U13631 (N_13631,N_12409,N_11410);
xnor U13632 (N_13632,N_11781,N_11434);
nor U13633 (N_13633,N_12299,N_11784);
and U13634 (N_13634,N_11503,N_11937);
and U13635 (N_13635,N_12400,N_11942);
nand U13636 (N_13636,N_12224,N_11392);
nor U13637 (N_13637,N_11301,N_11528);
and U13638 (N_13638,N_12358,N_11342);
xor U13639 (N_13639,N_12116,N_12281);
xnor U13640 (N_13640,N_12301,N_11872);
or U13641 (N_13641,N_11793,N_11625);
nand U13642 (N_13642,N_12124,N_11524);
nand U13643 (N_13643,N_11278,N_12423);
nand U13644 (N_13644,N_11329,N_11556);
nor U13645 (N_13645,N_12464,N_11797);
or U13646 (N_13646,N_11388,N_12402);
and U13647 (N_13647,N_11384,N_12172);
and U13648 (N_13648,N_12100,N_12252);
and U13649 (N_13649,N_12020,N_11738);
or U13650 (N_13650,N_12454,N_12172);
nor U13651 (N_13651,N_11401,N_12396);
and U13652 (N_13652,N_12232,N_12241);
xnor U13653 (N_13653,N_12411,N_12176);
and U13654 (N_13654,N_11992,N_12277);
nor U13655 (N_13655,N_11844,N_11313);
nor U13656 (N_13656,N_11933,N_11794);
xor U13657 (N_13657,N_12473,N_12116);
and U13658 (N_13658,N_12327,N_11955);
and U13659 (N_13659,N_12199,N_11897);
nor U13660 (N_13660,N_12195,N_11844);
xor U13661 (N_13661,N_12335,N_12344);
or U13662 (N_13662,N_11723,N_11975);
and U13663 (N_13663,N_12004,N_11555);
and U13664 (N_13664,N_12020,N_12466);
xor U13665 (N_13665,N_11772,N_12332);
or U13666 (N_13666,N_11892,N_11840);
nor U13667 (N_13667,N_11625,N_11519);
and U13668 (N_13668,N_11325,N_12277);
xnor U13669 (N_13669,N_12035,N_11349);
and U13670 (N_13670,N_12256,N_11311);
xnor U13671 (N_13671,N_12068,N_11586);
nor U13672 (N_13672,N_11693,N_11877);
or U13673 (N_13673,N_11425,N_11458);
xor U13674 (N_13674,N_11919,N_11298);
nor U13675 (N_13675,N_12490,N_12034);
xor U13676 (N_13676,N_11881,N_12393);
nor U13677 (N_13677,N_11864,N_11975);
nor U13678 (N_13678,N_12344,N_11875);
nor U13679 (N_13679,N_11429,N_12348);
nor U13680 (N_13680,N_11297,N_11629);
or U13681 (N_13681,N_11782,N_12366);
xnor U13682 (N_13682,N_11385,N_11598);
or U13683 (N_13683,N_11289,N_12444);
and U13684 (N_13684,N_12014,N_11598);
nor U13685 (N_13685,N_11979,N_11697);
or U13686 (N_13686,N_12016,N_11873);
xnor U13687 (N_13687,N_11949,N_12219);
xor U13688 (N_13688,N_12083,N_12001);
and U13689 (N_13689,N_12238,N_11883);
nor U13690 (N_13690,N_11461,N_11771);
xor U13691 (N_13691,N_12162,N_11358);
and U13692 (N_13692,N_12222,N_12471);
and U13693 (N_13693,N_12488,N_11848);
and U13694 (N_13694,N_11449,N_11504);
or U13695 (N_13695,N_11970,N_12371);
nand U13696 (N_13696,N_12092,N_11318);
and U13697 (N_13697,N_11579,N_12040);
nand U13698 (N_13698,N_11673,N_11497);
nor U13699 (N_13699,N_11299,N_12406);
and U13700 (N_13700,N_11481,N_12459);
xor U13701 (N_13701,N_11815,N_12137);
or U13702 (N_13702,N_11579,N_11508);
xnor U13703 (N_13703,N_11759,N_12173);
nand U13704 (N_13704,N_12340,N_11874);
nand U13705 (N_13705,N_11529,N_12289);
xnor U13706 (N_13706,N_11324,N_12063);
xnor U13707 (N_13707,N_11718,N_11997);
or U13708 (N_13708,N_12467,N_11440);
and U13709 (N_13709,N_11930,N_11679);
nor U13710 (N_13710,N_11677,N_11538);
or U13711 (N_13711,N_11566,N_12457);
nand U13712 (N_13712,N_11559,N_12091);
nor U13713 (N_13713,N_12298,N_12136);
nand U13714 (N_13714,N_12120,N_12181);
and U13715 (N_13715,N_11881,N_11357);
xnor U13716 (N_13716,N_12180,N_12019);
nor U13717 (N_13717,N_11793,N_11943);
nand U13718 (N_13718,N_11276,N_12191);
or U13719 (N_13719,N_11556,N_12023);
nand U13720 (N_13720,N_12222,N_11514);
nor U13721 (N_13721,N_12440,N_12162);
xor U13722 (N_13722,N_12103,N_12378);
or U13723 (N_13723,N_11479,N_12315);
nand U13724 (N_13724,N_11631,N_11397);
nand U13725 (N_13725,N_11797,N_11560);
or U13726 (N_13726,N_11504,N_12322);
nor U13727 (N_13727,N_12056,N_12262);
or U13728 (N_13728,N_12104,N_11749);
nand U13729 (N_13729,N_11467,N_11541);
xnor U13730 (N_13730,N_11749,N_12410);
and U13731 (N_13731,N_12117,N_11641);
nand U13732 (N_13732,N_11980,N_11543);
nand U13733 (N_13733,N_12297,N_11296);
or U13734 (N_13734,N_11844,N_11847);
nor U13735 (N_13735,N_11914,N_11869);
nor U13736 (N_13736,N_12342,N_11497);
and U13737 (N_13737,N_12413,N_11446);
xnor U13738 (N_13738,N_12057,N_12349);
xnor U13739 (N_13739,N_11678,N_11848);
nand U13740 (N_13740,N_11736,N_12466);
nand U13741 (N_13741,N_11377,N_12039);
nor U13742 (N_13742,N_12231,N_11905);
nor U13743 (N_13743,N_12117,N_11391);
and U13744 (N_13744,N_12114,N_12213);
and U13745 (N_13745,N_11556,N_11783);
nand U13746 (N_13746,N_11645,N_12303);
nor U13747 (N_13747,N_11677,N_11558);
and U13748 (N_13748,N_12025,N_12390);
nor U13749 (N_13749,N_11382,N_11422);
nor U13750 (N_13750,N_13279,N_12501);
and U13751 (N_13751,N_12730,N_12570);
xor U13752 (N_13752,N_13693,N_13244);
xnor U13753 (N_13753,N_13094,N_13123);
or U13754 (N_13754,N_13512,N_13377);
and U13755 (N_13755,N_13196,N_13487);
xor U13756 (N_13756,N_12644,N_13172);
or U13757 (N_13757,N_13453,N_13410);
xnor U13758 (N_13758,N_12913,N_13673);
xnor U13759 (N_13759,N_13523,N_13606);
nor U13760 (N_13760,N_12524,N_12582);
and U13761 (N_13761,N_13238,N_13021);
nand U13762 (N_13762,N_12540,N_12867);
xor U13763 (N_13763,N_12507,N_13239);
and U13764 (N_13764,N_13653,N_12775);
and U13765 (N_13765,N_13563,N_12684);
and U13766 (N_13766,N_13597,N_13380);
nor U13767 (N_13767,N_13630,N_13403);
xnor U13768 (N_13768,N_13249,N_13148);
nand U13769 (N_13769,N_13546,N_13030);
xnor U13770 (N_13770,N_12958,N_13068);
xnor U13771 (N_13771,N_12639,N_12990);
nand U13772 (N_13772,N_13526,N_13460);
or U13773 (N_13773,N_12973,N_13588);
or U13774 (N_13774,N_13703,N_13026);
or U13775 (N_13775,N_12919,N_13311);
and U13776 (N_13776,N_12549,N_12715);
nor U13777 (N_13777,N_13137,N_13428);
or U13778 (N_13778,N_12793,N_13086);
or U13779 (N_13779,N_13330,N_13479);
and U13780 (N_13780,N_13285,N_12536);
or U13781 (N_13781,N_13534,N_13560);
nor U13782 (N_13782,N_12643,N_12771);
or U13783 (N_13783,N_13045,N_12912);
xor U13784 (N_13784,N_13580,N_13223);
xnor U13785 (N_13785,N_13013,N_13685);
nand U13786 (N_13786,N_12816,N_13495);
xor U13787 (N_13787,N_12803,N_13491);
or U13788 (N_13788,N_13120,N_13423);
nor U13789 (N_13789,N_13517,N_13500);
or U13790 (N_13790,N_12889,N_13215);
nand U13791 (N_13791,N_13351,N_13452);
xor U13792 (N_13792,N_13054,N_13686);
or U13793 (N_13793,N_12817,N_13722);
nand U13794 (N_13794,N_13486,N_13401);
and U13795 (N_13795,N_12970,N_12753);
xnor U13796 (N_13796,N_13218,N_12598);
and U13797 (N_13797,N_13710,N_13438);
nand U13798 (N_13798,N_13352,N_13095);
xor U13799 (N_13799,N_13023,N_13040);
xnor U13800 (N_13800,N_13129,N_13724);
xnor U13801 (N_13801,N_12949,N_13419);
and U13802 (N_13802,N_13248,N_13125);
and U13803 (N_13803,N_12593,N_12967);
or U13804 (N_13804,N_13701,N_13201);
xor U13805 (N_13805,N_13658,N_12806);
or U13806 (N_13806,N_12691,N_13250);
and U13807 (N_13807,N_13187,N_13038);
nand U13808 (N_13808,N_12752,N_13144);
nor U13809 (N_13809,N_12703,N_12587);
nor U13810 (N_13810,N_12802,N_12899);
nor U13811 (N_13811,N_12689,N_12930);
nor U13812 (N_13812,N_13576,N_12845);
nor U13813 (N_13813,N_13212,N_12682);
or U13814 (N_13814,N_12884,N_13532);
and U13815 (N_13815,N_12903,N_13198);
xor U13816 (N_13816,N_13078,N_13474);
and U13817 (N_13817,N_13104,N_13591);
nand U13818 (N_13818,N_13374,N_13001);
xnor U13819 (N_13819,N_12736,N_12768);
xnor U13820 (N_13820,N_12788,N_13700);
and U13821 (N_13821,N_13189,N_12944);
nand U13822 (N_13822,N_13269,N_13458);
or U13823 (N_13823,N_12774,N_13048);
xor U13824 (N_13824,N_13052,N_13340);
xor U13825 (N_13825,N_13370,N_12995);
nand U13826 (N_13826,N_13375,N_13584);
or U13827 (N_13827,N_12947,N_13463);
and U13828 (N_13828,N_13719,N_13267);
xnor U13829 (N_13829,N_12993,N_13284);
and U13830 (N_13830,N_13437,N_12764);
and U13831 (N_13831,N_12792,N_13574);
and U13832 (N_13832,N_13390,N_13521);
nor U13833 (N_13833,N_13009,N_13691);
and U13834 (N_13834,N_13675,N_12581);
nand U13835 (N_13835,N_12698,N_12881);
xor U13836 (N_13836,N_12565,N_12592);
and U13837 (N_13837,N_12807,N_13613);
nand U13838 (N_13838,N_12572,N_12971);
or U13839 (N_13839,N_12800,N_13169);
and U13840 (N_13840,N_13501,N_13671);
nand U13841 (N_13841,N_12522,N_13631);
nor U13842 (N_13842,N_12630,N_13502);
nand U13843 (N_13843,N_12925,N_12789);
nor U13844 (N_13844,N_13348,N_12966);
xnor U13845 (N_13845,N_12586,N_12527);
xnor U13846 (N_13846,N_12997,N_13126);
and U13847 (N_13847,N_12762,N_12596);
or U13848 (N_13848,N_13027,N_12737);
xor U13849 (N_13849,N_13434,N_13720);
and U13850 (N_13850,N_13077,N_12657);
nand U13851 (N_13851,N_12875,N_13639);
nand U13852 (N_13852,N_12878,N_12887);
nand U13853 (N_13853,N_12797,N_12589);
or U13854 (N_13854,N_13273,N_13076);
nor U13855 (N_13855,N_12963,N_12917);
nand U13856 (N_13856,N_12674,N_12590);
or U13857 (N_13857,N_12526,N_13538);
nand U13858 (N_13858,N_13306,N_13436);
or U13859 (N_13859,N_13373,N_12724);
xor U13860 (N_13860,N_13002,N_13356);
nor U13861 (N_13861,N_12982,N_13413);
or U13862 (N_13862,N_13718,N_13012);
and U13863 (N_13863,N_12848,N_13282);
and U13864 (N_13864,N_12991,N_13733);
nor U13865 (N_13865,N_13025,N_12977);
nor U13866 (N_13866,N_13092,N_12563);
xor U13867 (N_13867,N_12514,N_13206);
and U13868 (N_13868,N_13432,N_13667);
nor U13869 (N_13869,N_12683,N_13657);
xor U13870 (N_13870,N_12740,N_13213);
xnor U13871 (N_13871,N_13583,N_13229);
nor U13872 (N_13872,N_13305,N_12650);
and U13873 (N_13873,N_12820,N_12861);
nand U13874 (N_13874,N_13354,N_13214);
or U13875 (N_13875,N_13032,N_13530);
or U13876 (N_13876,N_12760,N_13477);
or U13877 (N_13877,N_13661,N_13732);
xor U13878 (N_13878,N_13096,N_12747);
xor U13879 (N_13879,N_13743,N_13738);
nand U13880 (N_13880,N_13561,N_12904);
or U13881 (N_13881,N_12945,N_13222);
nor U13882 (N_13882,N_13531,N_12621);
xor U13883 (N_13883,N_12994,N_13258);
and U13884 (N_13884,N_12758,N_12710);
and U13885 (N_13885,N_12761,N_13283);
nand U13886 (N_13886,N_13292,N_13084);
nor U13887 (N_13887,N_12948,N_13513);
or U13888 (N_13888,N_13676,N_13360);
nor U13889 (N_13889,N_12687,N_12855);
nor U13890 (N_13890,N_12850,N_13665);
xnor U13891 (N_13891,N_12559,N_13582);
nor U13892 (N_13892,N_12525,N_13100);
nor U13893 (N_13893,N_13117,N_13216);
nor U13894 (N_13894,N_13058,N_13256);
and U13895 (N_13895,N_12599,N_13016);
and U13896 (N_13896,N_13579,N_13062);
and U13897 (N_13897,N_12631,N_13439);
nand U13898 (N_13898,N_12924,N_13539);
or U13899 (N_13899,N_13556,N_13227);
or U13900 (N_13900,N_12863,N_12645);
xnor U13901 (N_13901,N_13168,N_12574);
and U13902 (N_13902,N_12825,N_12809);
or U13903 (N_13903,N_12604,N_12942);
or U13904 (N_13904,N_12591,N_13492);
nor U13905 (N_13905,N_12634,N_12794);
and U13906 (N_13906,N_12512,N_13252);
or U13907 (N_13907,N_13398,N_13565);
or U13908 (N_13908,N_12838,N_13225);
or U13909 (N_13909,N_13527,N_13695);
xor U13910 (N_13910,N_13276,N_13644);
and U13911 (N_13911,N_13047,N_13571);
xnor U13912 (N_13912,N_12892,N_13660);
and U13913 (N_13913,N_12777,N_12579);
nand U13914 (N_13914,N_12923,N_13181);
nand U13915 (N_13915,N_12726,N_13368);
or U13916 (N_13916,N_12503,N_13620);
nand U13917 (N_13917,N_13072,N_13594);
or U13918 (N_13918,N_13601,N_12561);
nor U13919 (N_13919,N_13000,N_12988);
nor U13920 (N_13920,N_13706,N_12876);
or U13921 (N_13921,N_12989,N_12606);
nor U13922 (N_13922,N_13431,N_13290);
xnor U13923 (N_13923,N_12811,N_13666);
xnor U13924 (N_13924,N_12516,N_13656);
and U13925 (N_13925,N_12541,N_13024);
xnor U13926 (N_13926,N_12661,N_13589);
nor U13927 (N_13927,N_12801,N_12957);
nand U13928 (N_13928,N_13635,N_12713);
nand U13929 (N_13929,N_13332,N_13747);
nor U13930 (N_13930,N_13274,N_12712);
xnor U13931 (N_13931,N_13506,N_12840);
nor U13932 (N_13932,N_13060,N_13465);
or U13933 (N_13933,N_13412,N_12571);
or U13934 (N_13934,N_13327,N_12986);
xnor U13935 (N_13935,N_12920,N_13197);
nand U13936 (N_13936,N_13134,N_13698);
nor U13937 (N_13937,N_12669,N_13070);
nand U13938 (N_13938,N_13379,N_12699);
or U13939 (N_13939,N_13383,N_13010);
nor U13940 (N_13940,N_13586,N_13268);
nor U13941 (N_13941,N_13384,N_12984);
nor U13942 (N_13942,N_13299,N_13191);
and U13943 (N_13943,N_13240,N_13254);
nand U13944 (N_13944,N_13497,N_13572);
or U13945 (N_13945,N_12539,N_12719);
nand U13946 (N_13946,N_13643,N_12795);
nor U13947 (N_13947,N_12695,N_13610);
and U13948 (N_13948,N_12622,N_13470);
and U13949 (N_13949,N_13446,N_12672);
nor U13950 (N_13950,N_13320,N_12612);
nand U13951 (N_13951,N_12615,N_13081);
or U13952 (N_13952,N_12521,N_12562);
or U13953 (N_13953,N_13551,N_13464);
xor U13954 (N_13954,N_13646,N_12616);
and U13955 (N_13955,N_13199,N_12844);
or U13956 (N_13956,N_13259,N_13541);
or U13957 (N_13957,N_12696,N_12833);
xnor U13958 (N_13958,N_13457,N_13746);
nand U13959 (N_13959,N_13385,N_12856);
nor U13960 (N_13960,N_13429,N_13344);
xor U13961 (N_13961,N_13489,N_13114);
nor U13962 (N_13962,N_13231,N_13549);
or U13963 (N_13963,N_12648,N_13298);
or U13964 (N_13964,N_13696,N_13478);
xor U13965 (N_13965,N_12759,N_13494);
nor U13966 (N_13966,N_13272,N_13251);
and U13967 (N_13967,N_13550,N_12655);
xnor U13968 (N_13968,N_12603,N_12573);
nand U13969 (N_13969,N_13294,N_12564);
xnor U13970 (N_13970,N_13113,N_13605);
xor U13971 (N_13971,N_13087,N_12814);
or U13972 (N_13972,N_12767,N_13185);
xor U13973 (N_13973,N_12609,N_12731);
nand U13974 (N_13974,N_12543,N_13418);
xor U13975 (N_13975,N_12865,N_12854);
or U13976 (N_13976,N_12810,N_13558);
nand U13977 (N_13977,N_12992,N_12705);
or U13978 (N_13978,N_12721,N_12637);
xnor U13979 (N_13979,N_13246,N_12868);
nor U13980 (N_13980,N_13308,N_12941);
xor U13981 (N_13981,N_13573,N_12504);
nand U13982 (N_13982,N_13466,N_13587);
and U13983 (N_13983,N_13405,N_13441);
or U13984 (N_13984,N_13303,N_12769);
and U13985 (N_13985,N_12534,N_13603);
or U13986 (N_13986,N_13074,N_13049);
nor U13987 (N_13987,N_12813,N_12776);
and U13988 (N_13988,N_12659,N_13386);
nand U13989 (N_13989,N_12542,N_13101);
and U13990 (N_13990,N_13005,N_12658);
xor U13991 (N_13991,N_13055,N_12836);
nand U13992 (N_13992,N_12987,N_13515);
nand U13993 (N_13993,N_13493,N_13712);
nor U13994 (N_13994,N_13145,N_12723);
or U13995 (N_13995,N_13624,N_13670);
nand U13996 (N_13996,N_13545,N_12638);
and U13997 (N_13997,N_13618,N_12773);
and U13998 (N_13998,N_13063,N_12891);
or U13999 (N_13999,N_12938,N_13627);
and U14000 (N_14000,N_12931,N_13548);
or U14001 (N_14001,N_12700,N_12784);
nor U14002 (N_14002,N_13008,N_13116);
or U14003 (N_14003,N_12766,N_12937);
nor U14004 (N_14004,N_12751,N_12826);
or U14005 (N_14005,N_12842,N_12972);
and U14006 (N_14006,N_13683,N_13593);
or U14007 (N_14007,N_13397,N_13536);
nand U14008 (N_14008,N_13544,N_13173);
nor U14009 (N_14009,N_12859,N_13388);
nor U14010 (N_14010,N_12535,N_13018);
xnor U14011 (N_14011,N_12716,N_12894);
nor U14012 (N_14012,N_13089,N_13361);
nand U14013 (N_14013,N_13727,N_13190);
nor U14014 (N_14014,N_13233,N_13577);
or U14015 (N_14015,N_12862,N_13468);
nand U14016 (N_14016,N_13162,N_13209);
and U14017 (N_14017,N_12544,N_13031);
and U14018 (N_14018,N_13296,N_13245);
xnor U14019 (N_14019,N_13369,N_12694);
xnor U14020 (N_14020,N_13357,N_13518);
or U14021 (N_14021,N_12714,N_13358);
xor U14022 (N_14022,N_12821,N_13443);
or U14023 (N_14023,N_12602,N_13057);
nor U14024 (N_14024,N_12607,N_12569);
or U14025 (N_14025,N_12595,N_13219);
xor U14026 (N_14026,N_12664,N_12511);
nand U14027 (N_14027,N_12757,N_12896);
and U14028 (N_14028,N_13147,N_13575);
or U14029 (N_14029,N_12594,N_13614);
xnor U14030 (N_14030,N_13681,N_12837);
nor U14031 (N_14031,N_13456,N_12934);
or U14032 (N_14032,N_12585,N_12929);
nand U14033 (N_14033,N_13490,N_13247);
and U14034 (N_14034,N_13080,N_13371);
nor U14035 (N_14035,N_12677,N_12866);
nand U14036 (N_14036,N_12915,N_13473);
or U14037 (N_14037,N_13694,N_13411);
xnor U14038 (N_14038,N_13488,N_12629);
nand U14039 (N_14039,N_12831,N_13485);
xor U14040 (N_14040,N_13180,N_12545);
and U14041 (N_14041,N_12628,N_13736);
nand U14042 (N_14042,N_13406,N_13142);
xnor U14043 (N_14043,N_13399,N_13085);
nor U14044 (N_14044,N_13596,N_12567);
nor U14045 (N_14045,N_13499,N_13158);
xor U14046 (N_14046,N_13409,N_12897);
or U14047 (N_14047,N_13537,N_13297);
xor U14048 (N_14048,N_13309,N_12728);
nor U14049 (N_14049,N_12576,N_12560);
nor U14050 (N_14050,N_13365,N_12676);
or U14051 (N_14051,N_12588,N_12927);
or U14052 (N_14052,N_13564,N_12907);
or U14053 (N_14053,N_13083,N_13342);
nor U14054 (N_14054,N_13175,N_13204);
nand U14055 (N_14055,N_12508,N_13160);
or U14056 (N_14056,N_12790,N_12783);
nand U14057 (N_14057,N_13280,N_12605);
nor U14058 (N_14058,N_12946,N_13152);
nand U14059 (N_14059,N_13514,N_12523);
nor U14060 (N_14060,N_13133,N_13567);
nand U14061 (N_14061,N_13524,N_13715);
xnor U14062 (N_14062,N_13607,N_12553);
nand U14063 (N_14063,N_12787,N_13636);
xnor U14064 (N_14064,N_13394,N_12781);
nor U14065 (N_14065,N_12706,N_13061);
or U14066 (N_14066,N_12532,N_13236);
nand U14067 (N_14067,N_13598,N_12953);
nand U14068 (N_14068,N_13498,N_13393);
nor U14069 (N_14069,N_13228,N_13350);
or U14070 (N_14070,N_12968,N_13265);
nand U14071 (N_14071,N_12601,N_12746);
xnor U14072 (N_14072,N_13149,N_12969);
nand U14073 (N_14073,N_13726,N_12951);
and U14074 (N_14074,N_13600,N_12555);
nand U14075 (N_14075,N_13623,N_13260);
and U14076 (N_14076,N_12979,N_13407);
or U14077 (N_14077,N_12786,N_12898);
xor U14078 (N_14078,N_13243,N_13402);
xor U14079 (N_14079,N_13091,N_12575);
nand U14080 (N_14080,N_12685,N_13723);
nor U14081 (N_14081,N_13562,N_12708);
xor U14082 (N_14082,N_13680,N_13697);
nor U14083 (N_14083,N_13037,N_12743);
xor U14084 (N_14084,N_12597,N_13131);
or U14085 (N_14085,N_13621,N_13682);
nand U14086 (N_14086,N_12909,N_12846);
xnor U14087 (N_14087,N_13102,N_13638);
and U14088 (N_14088,N_12910,N_13034);
or U14089 (N_14089,N_12886,N_13122);
or U14090 (N_14090,N_12675,N_12882);
or U14091 (N_14091,N_12885,N_12557);
xnor U14092 (N_14092,N_13640,N_12611);
and U14093 (N_14093,N_12780,N_12707);
or U14094 (N_14094,N_12600,N_12617);
and U14095 (N_14095,N_12939,N_12546);
xnor U14096 (N_14096,N_13135,N_13017);
and U14097 (N_14097,N_13511,N_13569);
nand U14098 (N_14098,N_12916,N_13184);
xnor U14099 (N_14099,N_13318,N_13046);
and U14100 (N_14100,N_13232,N_13312);
nand U14101 (N_14101,N_13608,N_12921);
and U14102 (N_14102,N_12734,N_13166);
nor U14103 (N_14103,N_12952,N_12651);
xnor U14104 (N_14104,N_12547,N_13349);
or U14105 (N_14105,N_13645,N_12872);
and U14106 (N_14106,N_12652,N_13264);
nand U14107 (N_14107,N_12502,N_13447);
and U14108 (N_14108,N_13655,N_12940);
or U14109 (N_14109,N_12829,N_13036);
xnor U14110 (N_14110,N_13304,N_12890);
or U14111 (N_14111,N_13263,N_12956);
nor U14112 (N_14112,N_12819,N_13672);
or U14113 (N_14113,N_12619,N_13075);
or U14114 (N_14114,N_13554,N_12667);
nor U14115 (N_14115,N_13469,N_13699);
xor U14116 (N_14116,N_12692,N_13455);
and U14117 (N_14117,N_13302,N_13178);
or U14118 (N_14118,N_13728,N_13186);
and U14119 (N_14119,N_12818,N_12580);
xnor U14120 (N_14120,N_12983,N_12960);
or U14121 (N_14121,N_12640,N_13028);
xnor U14122 (N_14122,N_13689,N_12738);
nand U14123 (N_14123,N_13073,N_13355);
nand U14124 (N_14124,N_13004,N_13731);
and U14125 (N_14125,N_13041,N_12873);
or U14126 (N_14126,N_13353,N_13200);
nor U14127 (N_14127,N_13713,N_13748);
or U14128 (N_14128,N_12770,N_13414);
xor U14129 (N_14129,N_13420,N_13165);
nand U14130 (N_14130,N_12900,N_12888);
nor U14131 (N_14131,N_12624,N_12625);
or U14132 (N_14132,N_13121,N_13343);
or U14133 (N_14133,N_13341,N_13484);
xnor U14134 (N_14134,N_13053,N_12928);
and U14135 (N_14135,N_13103,N_13221);
xnor U14136 (N_14136,N_13064,N_13167);
and U14137 (N_14137,N_13734,N_12893);
nor U14138 (N_14138,N_13275,N_12725);
xor U14139 (N_14139,N_12517,N_13421);
or U14140 (N_14140,N_13338,N_12955);
xor U14141 (N_14141,N_12828,N_13615);
and U14142 (N_14142,N_13079,N_12779);
or U14143 (N_14143,N_13331,N_13171);
xor U14144 (N_14144,N_13188,N_12849);
nor U14145 (N_14145,N_13124,N_13744);
and U14146 (N_14146,N_12870,N_13322);
nand U14147 (N_14147,N_13444,N_12902);
and U14148 (N_14148,N_12618,N_13115);
xor U14149 (N_14149,N_13570,N_13157);
nand U14150 (N_14150,N_13707,N_13616);
nand U14151 (N_14151,N_12641,N_12911);
nand U14152 (N_14152,N_12702,N_12530);
xor U14153 (N_14153,N_13389,N_13067);
xnor U14154 (N_14154,N_13262,N_13301);
or U14155 (N_14155,N_13424,N_13329);
xnor U14156 (N_14156,N_13179,N_12805);
nor U14157 (N_14157,N_13449,N_12879);
nor U14158 (N_14158,N_13020,N_13622);
or U14159 (N_14159,N_13395,N_13519);
nand U14160 (N_14160,N_13730,N_12733);
or U14161 (N_14161,N_13663,N_12975);
and U14162 (N_14162,N_13011,N_13504);
and U14163 (N_14163,N_13033,N_12681);
xnor U14164 (N_14164,N_13347,N_13326);
xor U14165 (N_14165,N_12626,N_13345);
and U14166 (N_14166,N_13195,N_13234);
xnor U14167 (N_14167,N_13333,N_13430);
or U14168 (N_14168,N_13739,N_13459);
or U14169 (N_14169,N_13300,N_13127);
nor U14170 (N_14170,N_12799,N_13611);
nor U14171 (N_14171,N_13174,N_13679);
nor U14172 (N_14172,N_12670,N_12671);
or U14173 (N_14173,N_13372,N_12510);
nand U14174 (N_14174,N_12785,N_13128);
and U14175 (N_14175,N_12744,N_13328);
nor U14176 (N_14176,N_13266,N_13684);
and U14177 (N_14177,N_13362,N_13146);
nand U14178 (N_14178,N_13105,N_13462);
or U14179 (N_14179,N_13111,N_12750);
nand U14180 (N_14180,N_12922,N_12688);
and U14181 (N_14181,N_12509,N_12505);
xor U14182 (N_14182,N_12642,N_13692);
nor U14183 (N_14183,N_13217,N_13648);
nand U14184 (N_14184,N_13110,N_13293);
or U14185 (N_14185,N_12851,N_13286);
nand U14186 (N_14186,N_13056,N_13193);
and U14187 (N_14187,N_13566,N_13346);
or U14188 (N_14188,N_12627,N_13737);
and U14189 (N_14189,N_13677,N_13050);
nand U14190 (N_14190,N_13735,N_13609);
nand U14191 (N_14191,N_13650,N_13749);
or U14192 (N_14192,N_13578,N_13288);
nand U14193 (N_14193,N_13043,N_13604);
nand U14194 (N_14194,N_13107,N_13364);
nor U14195 (N_14195,N_12823,N_13687);
nand U14196 (N_14196,N_12964,N_13632);
nand U14197 (N_14197,N_12722,N_13535);
or U14198 (N_14198,N_13321,N_13422);
nor U14199 (N_14199,N_12690,N_13471);
and U14200 (N_14200,N_13003,N_13448);
nand U14201 (N_14201,N_13547,N_12739);
or U14202 (N_14202,N_12778,N_13163);
xor U14203 (N_14203,N_13503,N_13281);
or U14204 (N_14204,N_13617,N_13295);
nand U14205 (N_14205,N_12701,N_13323);
or U14206 (N_14206,N_13192,N_13704);
xor U14207 (N_14207,N_12880,N_13022);
or U14208 (N_14208,N_13654,N_12772);
nand U14209 (N_14209,N_12528,N_13130);
or U14210 (N_14210,N_13709,N_13143);
or U14211 (N_14211,N_13427,N_13161);
nand U14212 (N_14212,N_12735,N_12976);
xor U14213 (N_14213,N_12709,N_13602);
or U14214 (N_14214,N_13059,N_12860);
nor U14215 (N_14215,N_12832,N_12858);
or U14216 (N_14216,N_13315,N_12558);
or U14217 (N_14217,N_12720,N_12693);
nand U14218 (N_14218,N_13678,N_13674);
xor U14219 (N_14219,N_13480,N_12662);
and U14220 (N_14220,N_12798,N_12815);
nand U14221 (N_14221,N_12841,N_12538);
xor U14222 (N_14222,N_12895,N_13641);
nand U14223 (N_14223,N_12847,N_13220);
nand U14224 (N_14224,N_13664,N_13278);
and U14225 (N_14225,N_13118,N_13106);
nor U14226 (N_14226,N_13376,N_13261);
xnor U14227 (N_14227,N_13253,N_12636);
nand U14228 (N_14228,N_13559,N_13387);
nor U14229 (N_14229,N_13625,N_13093);
xor U14230 (N_14230,N_12548,N_12839);
nor U14231 (N_14231,N_12834,N_13150);
and U14232 (N_14232,N_13339,N_12943);
nand U14233 (N_14233,N_13426,N_13507);
or U14234 (N_14234,N_12623,N_12857);
and U14235 (N_14235,N_12804,N_12756);
or U14236 (N_14236,N_12635,N_12877);
or U14237 (N_14237,N_13391,N_12974);
xor U14238 (N_14238,N_12745,N_12749);
and U14239 (N_14239,N_13029,N_13416);
nand U14240 (N_14240,N_12936,N_12653);
xnor U14241 (N_14241,N_12978,N_13109);
nor U14242 (N_14242,N_13177,N_13467);
and U14243 (N_14243,N_13226,N_13359);
nand U14244 (N_14244,N_13065,N_13334);
nand U14245 (N_14245,N_12568,N_13505);
nand U14246 (N_14246,N_13522,N_13612);
nand U14247 (N_14247,N_12985,N_13740);
nor U14248 (N_14248,N_12914,N_13182);
and U14249 (N_14249,N_12727,N_13141);
nand U14250 (N_14250,N_13151,N_12717);
nor U14251 (N_14251,N_13289,N_13090);
xor U14252 (N_14252,N_13337,N_12665);
or U14253 (N_14253,N_12551,N_12999);
or U14254 (N_14254,N_13649,N_12763);
nor U14255 (N_14255,N_13019,N_12537);
nand U14256 (N_14256,N_12554,N_13496);
nand U14257 (N_14257,N_12577,N_13533);
and U14258 (N_14258,N_12908,N_13367);
xor U14259 (N_14259,N_12808,N_13400);
nand U14260 (N_14260,N_13408,N_12610);
nor U14261 (N_14261,N_12578,N_13378);
or U14262 (N_14262,N_13159,N_13741);
xnor U14263 (N_14263,N_13015,N_13335);
xnor U14264 (N_14264,N_12646,N_12741);
xnor U14265 (N_14265,N_12883,N_12932);
nor U14266 (N_14266,N_13205,N_13014);
nand U14267 (N_14267,N_13557,N_13425);
nor U14268 (N_14268,N_12673,N_13599);
xnor U14269 (N_14269,N_13417,N_13585);
nand U14270 (N_14270,N_12647,N_13714);
nor U14271 (N_14271,N_13396,N_12679);
nand U14272 (N_14272,N_13183,N_12566);
xnor U14273 (N_14273,N_13381,N_13555);
nand U14274 (N_14274,N_13237,N_13257);
xnor U14275 (N_14275,N_12918,N_13508);
nor U14276 (N_14276,N_13669,N_12620);
or U14277 (N_14277,N_12822,N_12748);
or U14278 (N_14278,N_13202,N_13450);
xor U14279 (N_14279,N_12998,N_13039);
xor U14280 (N_14280,N_13433,N_13528);
xor U14281 (N_14281,N_13721,N_13224);
or U14282 (N_14282,N_12906,N_13164);
xnor U14283 (N_14283,N_13442,N_12765);
or U14284 (N_14284,N_13155,N_13277);
and U14285 (N_14285,N_13088,N_13472);
xor U14286 (N_14286,N_13176,N_13454);
xor U14287 (N_14287,N_13042,N_12632);
nor U14288 (N_14288,N_13153,N_13287);
nand U14289 (N_14289,N_12959,N_13651);
or U14290 (N_14290,N_13170,N_13516);
nor U14291 (N_14291,N_13140,N_12519);
nor U14292 (N_14292,N_13235,N_13363);
nor U14293 (N_14293,N_13540,N_12901);
nand U14294 (N_14294,N_13210,N_13510);
nor U14295 (N_14295,N_12871,N_13581);
and U14296 (N_14296,N_12961,N_13404);
xor U14297 (N_14297,N_13336,N_13659);
nor U14298 (N_14298,N_13702,N_12518);
xnor U14299 (N_14299,N_12686,N_12660);
and U14300 (N_14300,N_12980,N_13119);
xnor U14301 (N_14301,N_12830,N_12529);
nand U14302 (N_14302,N_13194,N_12663);
and U14303 (N_14303,N_13319,N_13435);
or U14304 (N_14304,N_12556,N_13207);
xnor U14305 (N_14305,N_13668,N_13525);
nand U14306 (N_14306,N_13662,N_12926);
nand U14307 (N_14307,N_13520,N_12812);
nand U14308 (N_14308,N_13069,N_13270);
and U14309 (N_14309,N_12824,N_13392);
and U14310 (N_14310,N_13325,N_13112);
nor U14311 (N_14311,N_13482,N_13642);
nand U14312 (N_14312,N_13097,N_13099);
xnor U14313 (N_14313,N_13139,N_13382);
or U14314 (N_14314,N_13291,N_12933);
or U14315 (N_14315,N_13006,N_13366);
or U14316 (N_14316,N_13742,N_12649);
xnor U14317 (N_14317,N_12656,N_13690);
xor U14318 (N_14318,N_12755,N_12791);
or U14319 (N_14319,N_13035,N_12550);
nor U14320 (N_14320,N_12533,N_13051);
nand U14321 (N_14321,N_12874,N_13628);
nand U14322 (N_14322,N_12584,N_12633);
xor U14323 (N_14323,N_13461,N_13066);
nor U14324 (N_14324,N_13590,N_13688);
or U14325 (N_14325,N_13717,N_12853);
and U14326 (N_14326,N_12864,N_12668);
nor U14327 (N_14327,N_13241,N_13729);
nand U14328 (N_14328,N_13619,N_12500);
or U14329 (N_14329,N_13745,N_13633);
and U14330 (N_14330,N_13313,N_13595);
nor U14331 (N_14331,N_13705,N_13509);
nor U14332 (N_14332,N_12965,N_12729);
xnor U14333 (N_14333,N_13132,N_13637);
xor U14334 (N_14334,N_12935,N_13647);
and U14335 (N_14335,N_13136,N_13483);
xor U14336 (N_14336,N_12654,N_13314);
or U14337 (N_14337,N_12742,N_13307);
and U14338 (N_14338,N_13716,N_13629);
nor U14339 (N_14339,N_12796,N_12962);
nand U14340 (N_14340,N_13552,N_12513);
nor U14341 (N_14341,N_12608,N_13476);
nor U14342 (N_14342,N_12531,N_13543);
nand U14343 (N_14343,N_13451,N_12996);
nor U14344 (N_14344,N_13317,N_13529);
xor U14345 (N_14345,N_13568,N_12583);
and U14346 (N_14346,N_12981,N_13242);
and U14347 (N_14347,N_13440,N_12711);
nor U14348 (N_14348,N_13542,N_13138);
nand U14349 (N_14349,N_12782,N_12506);
nor U14350 (N_14350,N_12552,N_13708);
nand U14351 (N_14351,N_12954,N_13208);
nand U14352 (N_14352,N_12697,N_12704);
and U14353 (N_14353,N_13108,N_12732);
xor U14354 (N_14354,N_13230,N_13324);
and U14355 (N_14355,N_13082,N_12680);
or U14356 (N_14356,N_13481,N_13255);
and U14357 (N_14357,N_13203,N_13592);
xor U14358 (N_14358,N_13154,N_12852);
nand U14359 (N_14359,N_13044,N_12754);
nor U14360 (N_14360,N_12950,N_13415);
xnor U14361 (N_14361,N_12718,N_13316);
nor U14362 (N_14362,N_13711,N_13007);
xnor U14363 (N_14363,N_13553,N_13098);
nand U14364 (N_14364,N_13626,N_12905);
nor U14365 (N_14365,N_13725,N_13211);
nor U14366 (N_14366,N_13271,N_12614);
xnor U14367 (N_14367,N_13445,N_13652);
nand U14368 (N_14368,N_12666,N_12515);
or U14369 (N_14369,N_13475,N_12678);
and U14370 (N_14370,N_12869,N_12827);
or U14371 (N_14371,N_13634,N_13310);
or U14372 (N_14372,N_12613,N_13071);
and U14373 (N_14373,N_12835,N_13156);
or U14374 (N_14374,N_12843,N_12520);
or U14375 (N_14375,N_12530,N_12543);
nor U14376 (N_14376,N_13373,N_12840);
nand U14377 (N_14377,N_12503,N_13142);
xnor U14378 (N_14378,N_13356,N_12754);
nor U14379 (N_14379,N_13163,N_13197);
or U14380 (N_14380,N_12816,N_12561);
xor U14381 (N_14381,N_13136,N_13644);
and U14382 (N_14382,N_13674,N_13419);
and U14383 (N_14383,N_12506,N_13177);
or U14384 (N_14384,N_12633,N_12763);
xor U14385 (N_14385,N_13664,N_13647);
nor U14386 (N_14386,N_13004,N_12867);
or U14387 (N_14387,N_13114,N_12792);
xor U14388 (N_14388,N_12748,N_13640);
xor U14389 (N_14389,N_13488,N_12743);
xor U14390 (N_14390,N_13175,N_12968);
nor U14391 (N_14391,N_13208,N_13479);
nor U14392 (N_14392,N_12902,N_12958);
nor U14393 (N_14393,N_12725,N_12885);
nand U14394 (N_14394,N_13457,N_12642);
xnor U14395 (N_14395,N_13188,N_12700);
xor U14396 (N_14396,N_13644,N_12515);
xor U14397 (N_14397,N_13539,N_13453);
nand U14398 (N_14398,N_13343,N_12697);
and U14399 (N_14399,N_12732,N_12863);
and U14400 (N_14400,N_12778,N_12824);
and U14401 (N_14401,N_13673,N_13021);
nor U14402 (N_14402,N_13342,N_12815);
xor U14403 (N_14403,N_12704,N_13654);
nor U14404 (N_14404,N_13437,N_13612);
nor U14405 (N_14405,N_12886,N_13063);
nor U14406 (N_14406,N_13384,N_13005);
xnor U14407 (N_14407,N_12577,N_12506);
nand U14408 (N_14408,N_12538,N_13061);
xor U14409 (N_14409,N_13336,N_13504);
and U14410 (N_14410,N_13419,N_12563);
and U14411 (N_14411,N_12913,N_13325);
xnor U14412 (N_14412,N_13342,N_12980);
nand U14413 (N_14413,N_13240,N_13451);
and U14414 (N_14414,N_13422,N_12975);
or U14415 (N_14415,N_13013,N_13659);
xnor U14416 (N_14416,N_13067,N_13343);
and U14417 (N_14417,N_12598,N_13226);
or U14418 (N_14418,N_12793,N_12837);
or U14419 (N_14419,N_13157,N_13163);
nand U14420 (N_14420,N_13689,N_12762);
nor U14421 (N_14421,N_12668,N_12929);
nor U14422 (N_14422,N_13565,N_12824);
and U14423 (N_14423,N_13070,N_12730);
xor U14424 (N_14424,N_12718,N_13679);
nand U14425 (N_14425,N_12974,N_13711);
nand U14426 (N_14426,N_13497,N_12534);
nor U14427 (N_14427,N_13024,N_13036);
and U14428 (N_14428,N_13516,N_12720);
nor U14429 (N_14429,N_13408,N_13043);
and U14430 (N_14430,N_13186,N_13377);
xor U14431 (N_14431,N_13635,N_12548);
nand U14432 (N_14432,N_13396,N_13210);
xnor U14433 (N_14433,N_13353,N_12736);
nand U14434 (N_14434,N_13155,N_13696);
nand U14435 (N_14435,N_13410,N_13250);
nor U14436 (N_14436,N_13060,N_13209);
nand U14437 (N_14437,N_13538,N_13740);
nand U14438 (N_14438,N_12629,N_13322);
nor U14439 (N_14439,N_13194,N_12753);
or U14440 (N_14440,N_13292,N_13341);
or U14441 (N_14441,N_13549,N_12559);
and U14442 (N_14442,N_13530,N_13327);
and U14443 (N_14443,N_12582,N_13006);
xnor U14444 (N_14444,N_12768,N_13349);
nand U14445 (N_14445,N_13060,N_12912);
and U14446 (N_14446,N_13524,N_12986);
nor U14447 (N_14447,N_12503,N_12718);
or U14448 (N_14448,N_12575,N_12628);
xor U14449 (N_14449,N_13732,N_13272);
nor U14450 (N_14450,N_13159,N_12631);
nand U14451 (N_14451,N_13721,N_12597);
nor U14452 (N_14452,N_12770,N_13219);
or U14453 (N_14453,N_13544,N_13697);
xor U14454 (N_14454,N_13250,N_12569);
xor U14455 (N_14455,N_13494,N_12651);
nand U14456 (N_14456,N_13316,N_13572);
nor U14457 (N_14457,N_13202,N_12669);
nand U14458 (N_14458,N_13666,N_12724);
nand U14459 (N_14459,N_12556,N_13363);
or U14460 (N_14460,N_13305,N_12735);
nand U14461 (N_14461,N_12604,N_13709);
nand U14462 (N_14462,N_13381,N_13394);
nor U14463 (N_14463,N_13350,N_13517);
nor U14464 (N_14464,N_13026,N_13478);
xnor U14465 (N_14465,N_13401,N_13366);
nand U14466 (N_14466,N_13059,N_13339);
or U14467 (N_14467,N_13409,N_12917);
nor U14468 (N_14468,N_12715,N_13104);
and U14469 (N_14469,N_13561,N_12773);
and U14470 (N_14470,N_13377,N_12660);
or U14471 (N_14471,N_12653,N_13743);
nor U14472 (N_14472,N_12722,N_13530);
or U14473 (N_14473,N_13361,N_13049);
xnor U14474 (N_14474,N_13726,N_12549);
nor U14475 (N_14475,N_13615,N_13131);
or U14476 (N_14476,N_13091,N_12767);
nor U14477 (N_14477,N_13149,N_13151);
nand U14478 (N_14478,N_13480,N_13699);
or U14479 (N_14479,N_12926,N_13294);
nand U14480 (N_14480,N_13235,N_13561);
xnor U14481 (N_14481,N_12800,N_12742);
xnor U14482 (N_14482,N_13040,N_13132);
nand U14483 (N_14483,N_13399,N_12914);
nor U14484 (N_14484,N_12633,N_13262);
nor U14485 (N_14485,N_12696,N_13687);
and U14486 (N_14486,N_12618,N_13211);
nand U14487 (N_14487,N_13072,N_12554);
and U14488 (N_14488,N_12559,N_12536);
and U14489 (N_14489,N_13671,N_12511);
and U14490 (N_14490,N_13723,N_12758);
xor U14491 (N_14491,N_13436,N_12761);
or U14492 (N_14492,N_13697,N_13464);
nand U14493 (N_14493,N_13704,N_13582);
or U14494 (N_14494,N_13197,N_12889);
xnor U14495 (N_14495,N_12789,N_13051);
nor U14496 (N_14496,N_13022,N_12927);
xnor U14497 (N_14497,N_13306,N_13317);
nand U14498 (N_14498,N_12662,N_13727);
or U14499 (N_14499,N_13243,N_12679);
xor U14500 (N_14500,N_13074,N_13614);
nand U14501 (N_14501,N_13740,N_13335);
and U14502 (N_14502,N_13341,N_12666);
or U14503 (N_14503,N_13142,N_13638);
nor U14504 (N_14504,N_13412,N_12606);
or U14505 (N_14505,N_13744,N_13055);
or U14506 (N_14506,N_13178,N_13003);
or U14507 (N_14507,N_12516,N_13076);
xnor U14508 (N_14508,N_13144,N_13055);
xnor U14509 (N_14509,N_13440,N_13481);
xnor U14510 (N_14510,N_12645,N_13195);
or U14511 (N_14511,N_13110,N_13647);
nand U14512 (N_14512,N_12658,N_13137);
xnor U14513 (N_14513,N_12623,N_12987);
and U14514 (N_14514,N_13725,N_12833);
or U14515 (N_14515,N_13019,N_12740);
xnor U14516 (N_14516,N_13688,N_12501);
and U14517 (N_14517,N_13585,N_12523);
nor U14518 (N_14518,N_12868,N_13062);
nor U14519 (N_14519,N_13378,N_13180);
or U14520 (N_14520,N_12851,N_13128);
nor U14521 (N_14521,N_12699,N_12984);
and U14522 (N_14522,N_13478,N_13689);
and U14523 (N_14523,N_12747,N_13253);
nor U14524 (N_14524,N_13271,N_13350);
nand U14525 (N_14525,N_13020,N_13003);
nand U14526 (N_14526,N_13735,N_13305);
and U14527 (N_14527,N_13192,N_13237);
nand U14528 (N_14528,N_13211,N_13128);
or U14529 (N_14529,N_13335,N_13112);
or U14530 (N_14530,N_12539,N_13047);
nor U14531 (N_14531,N_13315,N_13531);
and U14532 (N_14532,N_13434,N_13397);
nor U14533 (N_14533,N_12894,N_13469);
xnor U14534 (N_14534,N_13073,N_13337);
nor U14535 (N_14535,N_12676,N_13110);
or U14536 (N_14536,N_12936,N_13167);
and U14537 (N_14537,N_12548,N_13139);
nor U14538 (N_14538,N_12946,N_13113);
xnor U14539 (N_14539,N_12855,N_13690);
nor U14540 (N_14540,N_13364,N_12901);
and U14541 (N_14541,N_12841,N_13496);
or U14542 (N_14542,N_12837,N_13218);
nor U14543 (N_14543,N_12870,N_12595);
xnor U14544 (N_14544,N_13395,N_12800);
or U14545 (N_14545,N_13575,N_12910);
nor U14546 (N_14546,N_13268,N_12935);
xnor U14547 (N_14547,N_13313,N_13526);
xor U14548 (N_14548,N_13017,N_13036);
and U14549 (N_14549,N_12639,N_12615);
nand U14550 (N_14550,N_13020,N_13696);
or U14551 (N_14551,N_13505,N_12985);
nand U14552 (N_14552,N_13428,N_12546);
nor U14553 (N_14553,N_12556,N_13111);
nand U14554 (N_14554,N_13237,N_13096);
nor U14555 (N_14555,N_13244,N_13360);
nand U14556 (N_14556,N_13268,N_13578);
and U14557 (N_14557,N_12997,N_13213);
and U14558 (N_14558,N_13588,N_13274);
xnor U14559 (N_14559,N_12631,N_12892);
xor U14560 (N_14560,N_13498,N_12760);
nand U14561 (N_14561,N_12692,N_13100);
nor U14562 (N_14562,N_13577,N_12611);
or U14563 (N_14563,N_12863,N_13504);
and U14564 (N_14564,N_12794,N_13543);
nand U14565 (N_14565,N_13547,N_13599);
xor U14566 (N_14566,N_12973,N_13434);
nor U14567 (N_14567,N_12541,N_12769);
nand U14568 (N_14568,N_12566,N_13169);
nor U14569 (N_14569,N_13594,N_13477);
and U14570 (N_14570,N_13480,N_13064);
nor U14571 (N_14571,N_13030,N_13516);
nand U14572 (N_14572,N_13548,N_13597);
nand U14573 (N_14573,N_12549,N_12971);
xor U14574 (N_14574,N_12788,N_12701);
or U14575 (N_14575,N_12963,N_13420);
or U14576 (N_14576,N_12908,N_13079);
xnor U14577 (N_14577,N_12671,N_12878);
xor U14578 (N_14578,N_13430,N_13018);
nor U14579 (N_14579,N_13044,N_13049);
nor U14580 (N_14580,N_13258,N_12956);
nand U14581 (N_14581,N_13421,N_12777);
xor U14582 (N_14582,N_13314,N_12513);
xnor U14583 (N_14583,N_13581,N_12615);
and U14584 (N_14584,N_12573,N_12972);
nand U14585 (N_14585,N_12990,N_13730);
or U14586 (N_14586,N_13124,N_12699);
nor U14587 (N_14587,N_12972,N_13524);
xor U14588 (N_14588,N_12999,N_12880);
or U14589 (N_14589,N_12787,N_13120);
nor U14590 (N_14590,N_12993,N_13078);
or U14591 (N_14591,N_13447,N_13680);
nor U14592 (N_14592,N_12995,N_12700);
xor U14593 (N_14593,N_13470,N_13051);
xor U14594 (N_14594,N_12757,N_13480);
nand U14595 (N_14595,N_13707,N_12830);
or U14596 (N_14596,N_12855,N_13495);
nor U14597 (N_14597,N_12846,N_13108);
xor U14598 (N_14598,N_13678,N_12772);
and U14599 (N_14599,N_12551,N_12784);
nor U14600 (N_14600,N_13730,N_13330);
or U14601 (N_14601,N_13718,N_13547);
nand U14602 (N_14602,N_13618,N_12738);
nand U14603 (N_14603,N_13380,N_12960);
xnor U14604 (N_14604,N_13123,N_12894);
and U14605 (N_14605,N_12750,N_12843);
nor U14606 (N_14606,N_13503,N_12950);
xor U14607 (N_14607,N_13744,N_13700);
and U14608 (N_14608,N_13565,N_12992);
or U14609 (N_14609,N_13095,N_13059);
nor U14610 (N_14610,N_12982,N_13101);
xnor U14611 (N_14611,N_12815,N_12835);
nand U14612 (N_14612,N_13128,N_13122);
xor U14613 (N_14613,N_12680,N_12671);
and U14614 (N_14614,N_12936,N_13227);
xor U14615 (N_14615,N_13608,N_13522);
or U14616 (N_14616,N_13517,N_13373);
or U14617 (N_14617,N_12720,N_13036);
xnor U14618 (N_14618,N_13445,N_13113);
nand U14619 (N_14619,N_12708,N_13628);
and U14620 (N_14620,N_13610,N_12957);
nor U14621 (N_14621,N_13244,N_13134);
xor U14622 (N_14622,N_13390,N_12539);
or U14623 (N_14623,N_13516,N_12845);
xnor U14624 (N_14624,N_13008,N_12758);
nor U14625 (N_14625,N_13560,N_13015);
xor U14626 (N_14626,N_12515,N_12837);
xnor U14627 (N_14627,N_13181,N_12652);
or U14628 (N_14628,N_13282,N_13126);
and U14629 (N_14629,N_13016,N_13066);
or U14630 (N_14630,N_12717,N_12872);
or U14631 (N_14631,N_13448,N_13045);
xnor U14632 (N_14632,N_13438,N_13386);
and U14633 (N_14633,N_13487,N_13369);
nor U14634 (N_14634,N_12807,N_13718);
and U14635 (N_14635,N_12902,N_13615);
xnor U14636 (N_14636,N_13175,N_13205);
and U14637 (N_14637,N_12606,N_13565);
nand U14638 (N_14638,N_13724,N_13351);
nand U14639 (N_14639,N_13186,N_12942);
and U14640 (N_14640,N_13239,N_13129);
xnor U14641 (N_14641,N_13159,N_13566);
xor U14642 (N_14642,N_13543,N_12949);
xor U14643 (N_14643,N_13583,N_12544);
nand U14644 (N_14644,N_12761,N_12887);
xnor U14645 (N_14645,N_13560,N_13040);
or U14646 (N_14646,N_13425,N_13410);
xnor U14647 (N_14647,N_12861,N_13605);
nand U14648 (N_14648,N_12879,N_12732);
and U14649 (N_14649,N_12842,N_13016);
xnor U14650 (N_14650,N_13555,N_12517);
nor U14651 (N_14651,N_12932,N_12579);
or U14652 (N_14652,N_13549,N_13290);
nor U14653 (N_14653,N_12725,N_13639);
nor U14654 (N_14654,N_13424,N_12781);
and U14655 (N_14655,N_13369,N_13546);
nand U14656 (N_14656,N_13655,N_13241);
nor U14657 (N_14657,N_13574,N_12535);
or U14658 (N_14658,N_12605,N_13540);
and U14659 (N_14659,N_12959,N_13469);
or U14660 (N_14660,N_12710,N_13626);
nor U14661 (N_14661,N_12877,N_12687);
xor U14662 (N_14662,N_13341,N_12696);
and U14663 (N_14663,N_12869,N_12625);
xor U14664 (N_14664,N_12830,N_13073);
nor U14665 (N_14665,N_12652,N_13061);
and U14666 (N_14666,N_12740,N_13276);
xnor U14667 (N_14667,N_12744,N_13631);
and U14668 (N_14668,N_13242,N_12775);
and U14669 (N_14669,N_13574,N_13385);
nand U14670 (N_14670,N_13363,N_12643);
nand U14671 (N_14671,N_12721,N_13441);
and U14672 (N_14672,N_13528,N_13536);
or U14673 (N_14673,N_12727,N_13364);
and U14674 (N_14674,N_12764,N_12845);
nand U14675 (N_14675,N_12967,N_13185);
or U14676 (N_14676,N_12872,N_13241);
nor U14677 (N_14677,N_12793,N_13464);
and U14678 (N_14678,N_13611,N_12761);
xnor U14679 (N_14679,N_12890,N_13635);
or U14680 (N_14680,N_12789,N_12888);
or U14681 (N_14681,N_12969,N_13547);
nor U14682 (N_14682,N_13702,N_13006);
xor U14683 (N_14683,N_12846,N_13306);
and U14684 (N_14684,N_13559,N_12601);
nand U14685 (N_14685,N_12822,N_12846);
or U14686 (N_14686,N_12703,N_13028);
xor U14687 (N_14687,N_13644,N_13238);
xnor U14688 (N_14688,N_12805,N_13148);
nand U14689 (N_14689,N_13450,N_13130);
xnor U14690 (N_14690,N_13647,N_13004);
nor U14691 (N_14691,N_12724,N_13396);
nand U14692 (N_14692,N_13191,N_12506);
or U14693 (N_14693,N_12561,N_12742);
and U14694 (N_14694,N_12638,N_12719);
or U14695 (N_14695,N_12512,N_13101);
or U14696 (N_14696,N_12873,N_13679);
nor U14697 (N_14697,N_12647,N_13449);
or U14698 (N_14698,N_12523,N_13299);
or U14699 (N_14699,N_13542,N_12907);
nand U14700 (N_14700,N_12994,N_13287);
nand U14701 (N_14701,N_13340,N_13443);
nor U14702 (N_14702,N_13463,N_13627);
or U14703 (N_14703,N_12698,N_13500);
or U14704 (N_14704,N_12592,N_12582);
nor U14705 (N_14705,N_13486,N_12681);
or U14706 (N_14706,N_13739,N_13482);
nand U14707 (N_14707,N_13063,N_13252);
xnor U14708 (N_14708,N_12844,N_13004);
nor U14709 (N_14709,N_13322,N_12910);
nor U14710 (N_14710,N_12561,N_12544);
xor U14711 (N_14711,N_13737,N_13247);
xor U14712 (N_14712,N_13232,N_13519);
xor U14713 (N_14713,N_13633,N_12909);
xnor U14714 (N_14714,N_13441,N_12625);
and U14715 (N_14715,N_12598,N_13005);
nor U14716 (N_14716,N_12890,N_12631);
nor U14717 (N_14717,N_13596,N_13168);
and U14718 (N_14718,N_13120,N_12567);
and U14719 (N_14719,N_13363,N_12590);
nor U14720 (N_14720,N_13572,N_12988);
nor U14721 (N_14721,N_13083,N_13090);
nor U14722 (N_14722,N_12520,N_12756);
or U14723 (N_14723,N_13426,N_13714);
xnor U14724 (N_14724,N_13354,N_12809);
nor U14725 (N_14725,N_13524,N_12559);
or U14726 (N_14726,N_13138,N_12681);
nor U14727 (N_14727,N_12738,N_13702);
xnor U14728 (N_14728,N_13396,N_12619);
or U14729 (N_14729,N_12679,N_12567);
and U14730 (N_14730,N_12630,N_13290);
xor U14731 (N_14731,N_13163,N_13139);
nand U14732 (N_14732,N_12852,N_12764);
or U14733 (N_14733,N_13693,N_12573);
xnor U14734 (N_14734,N_12882,N_13404);
or U14735 (N_14735,N_13507,N_12590);
nand U14736 (N_14736,N_13495,N_12663);
nand U14737 (N_14737,N_13597,N_13088);
and U14738 (N_14738,N_12664,N_13151);
xor U14739 (N_14739,N_12525,N_12781);
nand U14740 (N_14740,N_13373,N_13111);
xor U14741 (N_14741,N_12524,N_12594);
xnor U14742 (N_14742,N_13030,N_12708);
nand U14743 (N_14743,N_13624,N_13425);
nor U14744 (N_14744,N_13601,N_12547);
or U14745 (N_14745,N_13534,N_13717);
nor U14746 (N_14746,N_13444,N_12893);
or U14747 (N_14747,N_12875,N_12977);
xor U14748 (N_14748,N_12879,N_12691);
and U14749 (N_14749,N_12957,N_13354);
xor U14750 (N_14750,N_12700,N_13650);
xor U14751 (N_14751,N_13383,N_13645);
or U14752 (N_14752,N_12721,N_13045);
nor U14753 (N_14753,N_13533,N_13636);
xor U14754 (N_14754,N_12674,N_13363);
or U14755 (N_14755,N_12568,N_12785);
nor U14756 (N_14756,N_12635,N_13464);
nor U14757 (N_14757,N_13512,N_12648);
nand U14758 (N_14758,N_12849,N_13682);
or U14759 (N_14759,N_12551,N_13602);
nor U14760 (N_14760,N_13440,N_13176);
nand U14761 (N_14761,N_12912,N_13740);
nor U14762 (N_14762,N_13573,N_12508);
nand U14763 (N_14763,N_12650,N_13119);
nor U14764 (N_14764,N_13240,N_12528);
nor U14765 (N_14765,N_12547,N_12525);
or U14766 (N_14766,N_12759,N_12512);
and U14767 (N_14767,N_13049,N_12917);
and U14768 (N_14768,N_13396,N_12921);
nand U14769 (N_14769,N_13252,N_12585);
nand U14770 (N_14770,N_13210,N_12898);
nor U14771 (N_14771,N_12632,N_13724);
nor U14772 (N_14772,N_13170,N_13454);
xor U14773 (N_14773,N_13068,N_12578);
xor U14774 (N_14774,N_12916,N_13553);
or U14775 (N_14775,N_13691,N_13021);
or U14776 (N_14776,N_13555,N_12808);
nand U14777 (N_14777,N_13270,N_13684);
xnor U14778 (N_14778,N_13379,N_13632);
xor U14779 (N_14779,N_12554,N_12727);
nor U14780 (N_14780,N_13037,N_13599);
nand U14781 (N_14781,N_13710,N_12648);
nand U14782 (N_14782,N_12656,N_13015);
xnor U14783 (N_14783,N_12796,N_13609);
nor U14784 (N_14784,N_12690,N_12875);
xor U14785 (N_14785,N_13347,N_13010);
and U14786 (N_14786,N_13637,N_13022);
nor U14787 (N_14787,N_12671,N_12504);
and U14788 (N_14788,N_13561,N_13363);
or U14789 (N_14789,N_13340,N_12530);
or U14790 (N_14790,N_13470,N_12523);
and U14791 (N_14791,N_13366,N_12895);
and U14792 (N_14792,N_13083,N_13086);
or U14793 (N_14793,N_13475,N_13630);
and U14794 (N_14794,N_12821,N_13583);
xnor U14795 (N_14795,N_12534,N_13375);
xor U14796 (N_14796,N_12586,N_13686);
nand U14797 (N_14797,N_12748,N_12828);
and U14798 (N_14798,N_12992,N_13622);
and U14799 (N_14799,N_12829,N_13070);
xor U14800 (N_14800,N_13283,N_13303);
xnor U14801 (N_14801,N_13541,N_13694);
and U14802 (N_14802,N_13411,N_12880);
nand U14803 (N_14803,N_13362,N_13204);
or U14804 (N_14804,N_12890,N_13155);
nor U14805 (N_14805,N_12767,N_12641);
nand U14806 (N_14806,N_12678,N_13234);
and U14807 (N_14807,N_12708,N_13580);
xor U14808 (N_14808,N_13332,N_13715);
and U14809 (N_14809,N_13721,N_13718);
and U14810 (N_14810,N_13640,N_13148);
or U14811 (N_14811,N_13539,N_13588);
or U14812 (N_14812,N_12965,N_12653);
nor U14813 (N_14813,N_12671,N_12771);
nand U14814 (N_14814,N_13051,N_12783);
nor U14815 (N_14815,N_12574,N_13580);
nand U14816 (N_14816,N_12557,N_12828);
or U14817 (N_14817,N_13539,N_13673);
or U14818 (N_14818,N_12839,N_12942);
and U14819 (N_14819,N_13035,N_13707);
and U14820 (N_14820,N_13241,N_13405);
nor U14821 (N_14821,N_13206,N_13708);
nor U14822 (N_14822,N_12907,N_12741);
nor U14823 (N_14823,N_13721,N_12789);
nor U14824 (N_14824,N_13506,N_12512);
nor U14825 (N_14825,N_12933,N_12626);
or U14826 (N_14826,N_13502,N_13555);
and U14827 (N_14827,N_13132,N_13147);
or U14828 (N_14828,N_13437,N_13281);
nand U14829 (N_14829,N_13536,N_12832);
xnor U14830 (N_14830,N_13551,N_13146);
and U14831 (N_14831,N_13095,N_12679);
nand U14832 (N_14832,N_12941,N_13225);
and U14833 (N_14833,N_12745,N_13178);
and U14834 (N_14834,N_13434,N_12820);
nor U14835 (N_14835,N_12871,N_13211);
and U14836 (N_14836,N_13510,N_12686);
or U14837 (N_14837,N_12540,N_13109);
nand U14838 (N_14838,N_12529,N_13052);
xnor U14839 (N_14839,N_13536,N_13435);
nor U14840 (N_14840,N_12645,N_12747);
and U14841 (N_14841,N_13154,N_13193);
and U14842 (N_14842,N_12916,N_13678);
and U14843 (N_14843,N_13425,N_12937);
xnor U14844 (N_14844,N_12921,N_12788);
xnor U14845 (N_14845,N_12859,N_13145);
nor U14846 (N_14846,N_13176,N_12983);
xnor U14847 (N_14847,N_12709,N_13101);
nand U14848 (N_14848,N_12521,N_13121);
nand U14849 (N_14849,N_13734,N_13334);
nor U14850 (N_14850,N_13605,N_12770);
nor U14851 (N_14851,N_12800,N_12712);
or U14852 (N_14852,N_13212,N_12909);
nand U14853 (N_14853,N_13025,N_13111);
and U14854 (N_14854,N_12704,N_12658);
or U14855 (N_14855,N_13592,N_13566);
nand U14856 (N_14856,N_13167,N_12708);
and U14857 (N_14857,N_13059,N_12912);
or U14858 (N_14858,N_13543,N_13602);
and U14859 (N_14859,N_13055,N_13280);
nand U14860 (N_14860,N_13335,N_12895);
nor U14861 (N_14861,N_13275,N_13597);
or U14862 (N_14862,N_13554,N_13234);
and U14863 (N_14863,N_13433,N_13336);
or U14864 (N_14864,N_13212,N_13337);
or U14865 (N_14865,N_12521,N_12989);
or U14866 (N_14866,N_13100,N_13531);
and U14867 (N_14867,N_12584,N_12941);
and U14868 (N_14868,N_13362,N_13523);
and U14869 (N_14869,N_13180,N_12521);
and U14870 (N_14870,N_12888,N_13562);
and U14871 (N_14871,N_12793,N_13216);
xnor U14872 (N_14872,N_13438,N_12570);
and U14873 (N_14873,N_12867,N_13647);
nor U14874 (N_14874,N_13170,N_13648);
xor U14875 (N_14875,N_13411,N_12647);
or U14876 (N_14876,N_13658,N_12565);
xor U14877 (N_14877,N_13208,N_12709);
xnor U14878 (N_14878,N_12729,N_12832);
nor U14879 (N_14879,N_12892,N_12650);
nand U14880 (N_14880,N_13005,N_13562);
and U14881 (N_14881,N_13731,N_13733);
nor U14882 (N_14882,N_13487,N_12998);
and U14883 (N_14883,N_13562,N_13206);
or U14884 (N_14884,N_13209,N_13199);
nand U14885 (N_14885,N_13326,N_12599);
and U14886 (N_14886,N_12837,N_12562);
xor U14887 (N_14887,N_13183,N_12717);
nand U14888 (N_14888,N_12733,N_13298);
nor U14889 (N_14889,N_12637,N_13215);
xor U14890 (N_14890,N_12696,N_13387);
or U14891 (N_14891,N_13595,N_13573);
xor U14892 (N_14892,N_12781,N_12714);
xor U14893 (N_14893,N_13263,N_13195);
nand U14894 (N_14894,N_12762,N_13509);
nand U14895 (N_14895,N_13657,N_13642);
nor U14896 (N_14896,N_12670,N_13642);
or U14897 (N_14897,N_13680,N_12554);
nor U14898 (N_14898,N_12961,N_13347);
xnor U14899 (N_14899,N_12589,N_12891);
and U14900 (N_14900,N_12720,N_12809);
xor U14901 (N_14901,N_13608,N_13729);
and U14902 (N_14902,N_13312,N_13297);
or U14903 (N_14903,N_13454,N_13225);
nand U14904 (N_14904,N_13206,N_13339);
and U14905 (N_14905,N_12597,N_13082);
nor U14906 (N_14906,N_12580,N_13542);
or U14907 (N_14907,N_12561,N_13055);
or U14908 (N_14908,N_13023,N_13710);
and U14909 (N_14909,N_13359,N_12618);
xnor U14910 (N_14910,N_13167,N_12861);
or U14911 (N_14911,N_13265,N_13430);
nand U14912 (N_14912,N_13667,N_13225);
or U14913 (N_14913,N_13448,N_13659);
nor U14914 (N_14914,N_12572,N_12986);
nand U14915 (N_14915,N_12870,N_12548);
or U14916 (N_14916,N_12801,N_12645);
nand U14917 (N_14917,N_13416,N_12588);
and U14918 (N_14918,N_13416,N_12558);
xor U14919 (N_14919,N_12865,N_12556);
xor U14920 (N_14920,N_12844,N_12914);
nor U14921 (N_14921,N_12528,N_13267);
nand U14922 (N_14922,N_12602,N_12560);
nand U14923 (N_14923,N_13551,N_13555);
and U14924 (N_14924,N_13241,N_12791);
or U14925 (N_14925,N_13087,N_12501);
nand U14926 (N_14926,N_12832,N_12894);
or U14927 (N_14927,N_13239,N_12952);
nand U14928 (N_14928,N_12844,N_13313);
and U14929 (N_14929,N_13513,N_13012);
nand U14930 (N_14930,N_13085,N_13135);
nor U14931 (N_14931,N_12993,N_13076);
nand U14932 (N_14932,N_13731,N_13038);
and U14933 (N_14933,N_13692,N_12794);
nor U14934 (N_14934,N_13085,N_13498);
nor U14935 (N_14935,N_13698,N_13238);
and U14936 (N_14936,N_13192,N_12810);
or U14937 (N_14937,N_12524,N_13490);
nand U14938 (N_14938,N_13447,N_12591);
xor U14939 (N_14939,N_13424,N_13527);
nor U14940 (N_14940,N_13075,N_13031);
xor U14941 (N_14941,N_12722,N_12655);
or U14942 (N_14942,N_13735,N_13403);
nor U14943 (N_14943,N_13297,N_13281);
xnor U14944 (N_14944,N_12628,N_13740);
or U14945 (N_14945,N_13305,N_13558);
and U14946 (N_14946,N_12714,N_12630);
and U14947 (N_14947,N_12588,N_12928);
and U14948 (N_14948,N_12807,N_13676);
xor U14949 (N_14949,N_13542,N_13431);
nor U14950 (N_14950,N_13249,N_13124);
nor U14951 (N_14951,N_13260,N_12533);
nand U14952 (N_14952,N_13624,N_12850);
or U14953 (N_14953,N_13404,N_12509);
nand U14954 (N_14954,N_12580,N_13641);
nand U14955 (N_14955,N_12806,N_13622);
nand U14956 (N_14956,N_12561,N_12737);
xnor U14957 (N_14957,N_13430,N_13233);
nor U14958 (N_14958,N_13326,N_13461);
nor U14959 (N_14959,N_13253,N_12930);
and U14960 (N_14960,N_13551,N_12842);
or U14961 (N_14961,N_13732,N_13747);
or U14962 (N_14962,N_13290,N_12796);
and U14963 (N_14963,N_13496,N_13417);
or U14964 (N_14964,N_13518,N_12655);
and U14965 (N_14965,N_13703,N_13518);
and U14966 (N_14966,N_12969,N_13045);
and U14967 (N_14967,N_13225,N_13546);
and U14968 (N_14968,N_13148,N_12507);
nand U14969 (N_14969,N_13275,N_13481);
nor U14970 (N_14970,N_13154,N_12976);
and U14971 (N_14971,N_13554,N_12998);
xor U14972 (N_14972,N_13435,N_13184);
xnor U14973 (N_14973,N_13277,N_13545);
nor U14974 (N_14974,N_13716,N_12700);
nand U14975 (N_14975,N_13112,N_12937);
and U14976 (N_14976,N_13111,N_12837);
or U14977 (N_14977,N_12778,N_13541);
and U14978 (N_14978,N_12757,N_13710);
nand U14979 (N_14979,N_12918,N_13070);
or U14980 (N_14980,N_13408,N_12888);
or U14981 (N_14981,N_12519,N_12552);
and U14982 (N_14982,N_13679,N_13054);
and U14983 (N_14983,N_12999,N_12623);
and U14984 (N_14984,N_13553,N_12632);
nand U14985 (N_14985,N_13508,N_13193);
nor U14986 (N_14986,N_12941,N_13429);
xnor U14987 (N_14987,N_13486,N_13199);
and U14988 (N_14988,N_12755,N_12691);
nor U14989 (N_14989,N_13070,N_12711);
nand U14990 (N_14990,N_13540,N_13132);
or U14991 (N_14991,N_13072,N_13447);
nand U14992 (N_14992,N_13079,N_12959);
or U14993 (N_14993,N_12703,N_12680);
nor U14994 (N_14994,N_12852,N_13384);
nor U14995 (N_14995,N_12776,N_13336);
nor U14996 (N_14996,N_12951,N_13634);
or U14997 (N_14997,N_13327,N_13156);
xnor U14998 (N_14998,N_13468,N_13408);
nand U14999 (N_14999,N_12795,N_12763);
xor U15000 (N_15000,N_14728,N_14120);
nor U15001 (N_15001,N_14347,N_14431);
xnor U15002 (N_15002,N_14534,N_14752);
nand U15003 (N_15003,N_14593,N_14675);
xnor U15004 (N_15004,N_14931,N_14296);
or U15005 (N_15005,N_14771,N_13928);
and U15006 (N_15006,N_14326,N_14208);
xnor U15007 (N_15007,N_14690,N_14730);
nor U15008 (N_15008,N_14579,N_14928);
nand U15009 (N_15009,N_14516,N_14169);
and U15010 (N_15010,N_14736,N_14681);
nor U15011 (N_15011,N_14100,N_14842);
and U15012 (N_15012,N_14787,N_14987);
or U15013 (N_15013,N_14857,N_14570);
xor U15014 (N_15014,N_14606,N_13945);
or U15015 (N_15015,N_14267,N_14035);
and U15016 (N_15016,N_13785,N_13895);
xnor U15017 (N_15017,N_14163,N_14676);
nand U15018 (N_15018,N_14007,N_14332);
nor U15019 (N_15019,N_14656,N_14571);
xor U15020 (N_15020,N_13993,N_14995);
or U15021 (N_15021,N_14459,N_14301);
or U15022 (N_15022,N_13869,N_13891);
and U15023 (N_15023,N_14381,N_14474);
and U15024 (N_15024,N_14444,N_14637);
or U15025 (N_15025,N_14945,N_14879);
nand U15026 (N_15026,N_14909,N_14456);
xor U15027 (N_15027,N_14652,N_14303);
xnor U15028 (N_15028,N_13797,N_14461);
nand U15029 (N_15029,N_14822,N_14940);
or U15030 (N_15030,N_14698,N_14045);
xnor U15031 (N_15031,N_14733,N_14290);
nand U15032 (N_15032,N_14544,N_14358);
and U15033 (N_15033,N_14337,N_14318);
nor U15034 (N_15034,N_14229,N_14595);
nand U15035 (N_15035,N_14075,N_14311);
or U15036 (N_15036,N_14006,N_14111);
xor U15037 (N_15037,N_14071,N_13990);
nor U15038 (N_15038,N_14869,N_14629);
or U15039 (N_15039,N_14216,N_14789);
xnor U15040 (N_15040,N_14126,N_14648);
nor U15041 (N_15041,N_14955,N_14322);
nand U15042 (N_15042,N_14307,N_13949);
and U15043 (N_15043,N_14333,N_14014);
and U15044 (N_15044,N_13953,N_14785);
nor U15045 (N_15045,N_14118,N_13817);
and U15046 (N_15046,N_14882,N_13936);
xnor U15047 (N_15047,N_14486,N_14349);
xnor U15048 (N_15048,N_13824,N_14466);
and U15049 (N_15049,N_14195,N_14555);
or U15050 (N_15050,N_14625,N_14884);
or U15051 (N_15051,N_14027,N_14259);
xnor U15052 (N_15052,N_14268,N_14241);
and U15053 (N_15053,N_14697,N_14427);
xnor U15054 (N_15054,N_13951,N_14012);
nand U15055 (N_15055,N_13792,N_14578);
xnor U15056 (N_15056,N_14392,N_13809);
and U15057 (N_15057,N_14297,N_13777);
or U15058 (N_15058,N_14335,N_14385);
nand U15059 (N_15059,N_14946,N_13909);
or U15060 (N_15060,N_14407,N_13944);
or U15061 (N_15061,N_13986,N_14061);
xor U15062 (N_15062,N_14867,N_14680);
nand U15063 (N_15063,N_14896,N_14808);
nor U15064 (N_15064,N_13985,N_14149);
xor U15065 (N_15065,N_13873,N_14091);
nand U15066 (N_15066,N_14031,N_14125);
nor U15067 (N_15067,N_14905,N_14965);
xnor U15068 (N_15068,N_14141,N_13798);
xnor U15069 (N_15069,N_14541,N_13967);
or U15070 (N_15070,N_13803,N_14339);
xnor U15071 (N_15071,N_14168,N_14959);
or U15072 (N_15072,N_14877,N_14596);
and U15073 (N_15073,N_14806,N_14791);
or U15074 (N_15074,N_13889,N_13752);
or U15075 (N_15075,N_14671,N_14384);
nand U15076 (N_15076,N_14131,N_13979);
nand U15077 (N_15077,N_14066,N_13906);
nor U15078 (N_15078,N_14522,N_14503);
nor U15079 (N_15079,N_13841,N_13907);
nor U15080 (N_15080,N_14559,N_14258);
and U15081 (N_15081,N_13815,N_14623);
nand U15082 (N_15082,N_13919,N_13755);
or U15083 (N_15083,N_14792,N_13876);
nor U15084 (N_15084,N_14451,N_13789);
or U15085 (N_15085,N_13839,N_13956);
and U15086 (N_15086,N_13939,N_13870);
nor U15087 (N_15087,N_14479,N_14353);
and U15088 (N_15088,N_14925,N_14133);
and U15089 (N_15089,N_14527,N_14532);
or U15090 (N_15090,N_13925,N_13838);
xnor U15091 (N_15091,N_14183,N_14722);
and U15092 (N_15092,N_14394,N_13753);
and U15093 (N_15093,N_14432,N_14615);
xnor U15094 (N_15094,N_14600,N_14719);
nor U15095 (N_15095,N_14247,N_14288);
nand U15096 (N_15096,N_13998,N_14452);
nand U15097 (N_15097,N_14420,N_14199);
nor U15098 (N_15098,N_13900,N_13999);
or U15099 (N_15099,N_14849,N_14561);
nor U15100 (N_15100,N_13854,N_14017);
nor U15101 (N_15101,N_14670,N_14812);
and U15102 (N_15102,N_13968,N_14000);
nand U15103 (N_15103,N_14374,N_14298);
or U15104 (N_15104,N_14363,N_14252);
nor U15105 (N_15105,N_14814,N_14881);
and U15106 (N_15106,N_14110,N_14783);
nand U15107 (N_15107,N_14362,N_14661);
or U15108 (N_15108,N_14412,N_14552);
xnor U15109 (N_15109,N_14684,N_14211);
nor U15110 (N_15110,N_14630,N_14469);
xor U15111 (N_15111,N_13970,N_13862);
and U15112 (N_15112,N_14817,N_14351);
and U15113 (N_15113,N_14210,N_14793);
nor U15114 (N_15114,N_14261,N_14878);
nor U15115 (N_15115,N_14009,N_14321);
nand U15116 (N_15116,N_14341,N_14725);
and U15117 (N_15117,N_14497,N_14203);
and U15118 (N_15118,N_14748,N_14060);
or U15119 (N_15119,N_13856,N_14860);
nand U15120 (N_15120,N_14189,N_14607);
nor U15121 (N_15121,N_14373,N_14865);
nor U15122 (N_15122,N_14836,N_14313);
nand U15123 (N_15123,N_14440,N_13959);
and U15124 (N_15124,N_13762,N_14610);
nor U15125 (N_15125,N_13886,N_14853);
nor U15126 (N_15126,N_14778,N_14482);
nor U15127 (N_15127,N_14892,N_14749);
or U15128 (N_15128,N_14651,N_14434);
or U15129 (N_15129,N_14284,N_14171);
nand U15130 (N_15130,N_14591,N_14868);
and U15131 (N_15131,N_14426,N_14634);
and U15132 (N_15132,N_13989,N_14939);
nand U15133 (N_15133,N_14696,N_14077);
and U15134 (N_15134,N_14574,N_14714);
and U15135 (N_15135,N_14985,N_14597);
nor U15136 (N_15136,N_14174,N_14370);
xor U15137 (N_15137,N_13830,N_14535);
nand U15138 (N_15138,N_14057,N_14908);
and U15139 (N_15139,N_14643,N_14694);
or U15140 (N_15140,N_14734,N_14958);
nand U15141 (N_15141,N_14888,N_13950);
nor U15142 (N_15142,N_14399,N_14847);
and U15143 (N_15143,N_14155,N_14864);
or U15144 (N_15144,N_14705,N_14269);
xnor U15145 (N_15145,N_14816,N_14530);
nor U15146 (N_15146,N_13831,N_14108);
xnor U15147 (N_15147,N_13794,N_14492);
xor U15148 (N_15148,N_14220,N_14685);
or U15149 (N_15149,N_14813,N_14973);
nand U15150 (N_15150,N_14720,N_14902);
xor U15151 (N_15151,N_14213,N_14447);
xor U15152 (N_15152,N_13784,N_13877);
nor U15153 (N_15153,N_14123,N_14344);
or U15154 (N_15154,N_14646,N_14274);
xnor U15155 (N_15155,N_14202,N_13757);
and U15156 (N_15156,N_13751,N_14718);
and U15157 (N_15157,N_14617,N_14078);
or U15158 (N_15158,N_14821,N_14063);
nor U15159 (N_15159,N_13810,N_14033);
nor U15160 (N_15160,N_14312,N_14846);
xnor U15161 (N_15161,N_14895,N_14546);
xnor U15162 (N_15162,N_14343,N_14134);
or U15163 (N_15163,N_13901,N_14473);
nor U15164 (N_15164,N_13811,N_13954);
nand U15165 (N_15165,N_14419,N_14716);
and U15166 (N_15166,N_14488,N_14914);
or U15167 (N_15167,N_14186,N_13804);
nand U15168 (N_15168,N_14660,N_14390);
xor U15169 (N_15169,N_13855,N_13992);
or U15170 (N_15170,N_14624,N_14010);
nand U15171 (N_15171,N_14135,N_14187);
nand U15172 (N_15172,N_13997,N_14599);
nand U15173 (N_15173,N_14081,N_14139);
nand U15174 (N_15174,N_14166,N_14413);
xnor U15175 (N_15175,N_14543,N_14568);
xnor U15176 (N_15176,N_14467,N_14885);
nor U15177 (N_15177,N_13933,N_14383);
xnor U15178 (N_15178,N_14132,N_13756);
xnor U15179 (N_15179,N_14891,N_14701);
xnor U15180 (N_15180,N_13969,N_14319);
nor U15181 (N_15181,N_14105,N_14635);
and U15182 (N_15182,N_14359,N_14201);
xnor U15183 (N_15183,N_14244,N_14436);
xnor U15184 (N_15184,N_14899,N_14365);
xor U15185 (N_15185,N_14641,N_14861);
and U15186 (N_15186,N_14415,N_14683);
or U15187 (N_15187,N_13917,N_14445);
nor U15188 (N_15188,N_13929,N_14198);
nor U15189 (N_15189,N_14471,N_14936);
xnor U15190 (N_15190,N_14996,N_14128);
xnor U15191 (N_15191,N_13942,N_14160);
nor U15192 (N_15192,N_14382,N_13973);
or U15193 (N_15193,N_14205,N_14871);
nor U15194 (N_15194,N_14421,N_13828);
and U15195 (N_15195,N_14018,N_14124);
nor U15196 (N_15196,N_13982,N_13975);
xnor U15197 (N_15197,N_14011,N_14904);
or U15198 (N_15198,N_13972,N_13832);
and U15199 (N_15199,N_14372,N_13938);
and U15200 (N_15200,N_13913,N_13890);
nor U15201 (N_15201,N_14355,N_14352);
nor U15202 (N_15202,N_14642,N_13754);
and U15203 (N_15203,N_14517,N_13984);
xor U15204 (N_15204,N_13914,N_13920);
xnor U15205 (N_15205,N_14872,N_14059);
nor U15206 (N_15206,N_14531,N_14260);
or U15207 (N_15207,N_13868,N_13885);
nor U15208 (N_15208,N_14622,N_14336);
and U15209 (N_15209,N_14450,N_14754);
xnor U15210 (N_15210,N_13981,N_14502);
nand U15211 (N_15211,N_14234,N_14453);
and U15212 (N_15212,N_14549,N_14655);
xor U15213 (N_15213,N_14550,N_14056);
and U15214 (N_15214,N_13960,N_13971);
or U15215 (N_15215,N_13910,N_14978);
xnor U15216 (N_15216,N_14414,N_14324);
nand U15217 (N_15217,N_14115,N_14947);
and U15218 (N_15218,N_14994,N_13926);
nor U15219 (N_15219,N_14150,N_13996);
nor U15220 (N_15220,N_14524,N_14140);
and U15221 (N_15221,N_14691,N_13922);
and U15222 (N_15222,N_14569,N_14442);
xnor U15223 (N_15223,N_13905,N_14961);
nand U15224 (N_15224,N_14092,N_14292);
xor U15225 (N_15225,N_14233,N_14929);
xnor U15226 (N_15226,N_13871,N_14026);
nor U15227 (N_15227,N_14299,N_14911);
nor U15228 (N_15228,N_14796,N_14693);
nand U15229 (N_15229,N_13779,N_14251);
nor U15230 (N_15230,N_14536,N_14040);
or U15231 (N_15231,N_14448,N_14400);
nor U15232 (N_15232,N_14048,N_14393);
nand U15233 (N_15233,N_13816,N_14470);
and U15234 (N_15234,N_14455,N_14493);
and U15235 (N_15235,N_14594,N_14300);
xor U15236 (N_15236,N_14927,N_14844);
nand U15237 (N_15237,N_14880,N_14176);
nor U15238 (N_15238,N_14246,N_14222);
nand U15239 (N_15239,N_14551,N_13976);
nand U15240 (N_15240,N_13836,N_14036);
and U15241 (N_15241,N_14560,N_14523);
xnor U15242 (N_15242,N_14030,N_14308);
and U15243 (N_15243,N_14807,N_14788);
or U15244 (N_15244,N_14766,N_14511);
nand U15245 (N_15245,N_13850,N_14510);
nor U15246 (N_15246,N_14922,N_14538);
xnor U15247 (N_15247,N_14238,N_14484);
nor U15248 (N_15248,N_13835,N_14547);
and U15249 (N_15249,N_13892,N_14378);
or U15250 (N_15250,N_13758,N_13820);
nor U15251 (N_15251,N_14981,N_14285);
nand U15252 (N_15252,N_14874,N_14741);
xnor U15253 (N_15253,N_14514,N_14627);
xor U15254 (N_15254,N_13995,N_14264);
xnor U15255 (N_15255,N_13894,N_13888);
xnor U15256 (N_15256,N_14818,N_13823);
or U15257 (N_15257,N_14856,N_14245);
xnor U15258 (N_15258,N_14657,N_14567);
nor U15259 (N_15259,N_14515,N_14411);
and U15260 (N_15260,N_13875,N_13987);
nor U15261 (N_15261,N_13843,N_14416);
nor U15262 (N_15262,N_13897,N_14287);
and U15263 (N_15263,N_13874,N_13916);
xnor U15264 (N_15264,N_14329,N_14013);
nor U15265 (N_15265,N_14525,N_14257);
and U15266 (N_15266,N_14016,N_14106);
xnor U15267 (N_15267,N_14395,N_13883);
and U15268 (N_15268,N_14553,N_14673);
or U15269 (N_15269,N_14920,N_14932);
and U15270 (N_15270,N_13872,N_14197);
or U15271 (N_15271,N_14540,N_14859);
nor U15272 (N_15272,N_14829,N_14811);
xor U15273 (N_15273,N_14957,N_14357);
nand U15274 (N_15274,N_13833,N_14430);
nand U15275 (N_15275,N_13902,N_14023);
and U15276 (N_15276,N_14726,N_13851);
xor U15277 (N_15277,N_14249,N_14750);
or U15278 (N_15278,N_14963,N_14636);
xnor U15279 (N_15279,N_13846,N_13799);
xnor U15280 (N_15280,N_14645,N_14763);
nand U15281 (N_15281,N_14397,N_14401);
xnor U15282 (N_15282,N_13860,N_14790);
nand U15283 (N_15283,N_14585,N_14121);
xor U15284 (N_15284,N_14855,N_14103);
xnor U15285 (N_15285,N_14387,N_14148);
or U15286 (N_15286,N_14196,N_14388);
or U15287 (N_15287,N_14944,N_14602);
nor U15288 (N_15288,N_14433,N_14508);
nand U15289 (N_15289,N_14147,N_14991);
and U15290 (N_15290,N_14699,N_14500);
nor U15291 (N_15291,N_14153,N_14917);
xnor U15292 (N_15292,N_14085,N_13840);
nand U15293 (N_15293,N_13826,N_14679);
and U15294 (N_15294,N_14028,N_13988);
xor U15295 (N_15295,N_14731,N_14145);
nand U15296 (N_15296,N_14239,N_13834);
nand U15297 (N_15297,N_14406,N_14338);
or U15298 (N_15298,N_14949,N_14727);
nand U15299 (N_15299,N_14224,N_14327);
and U15300 (N_15300,N_14494,N_14611);
nor U15301 (N_15301,N_13930,N_14175);
nor U15302 (N_15302,N_14226,N_14744);
nor U15303 (N_15303,N_14770,N_14889);
and U15304 (N_15304,N_14590,N_13941);
nor U15305 (N_15305,N_14154,N_14747);
and U15306 (N_15306,N_14248,N_14490);
and U15307 (N_15307,N_14631,N_14505);
and U15308 (N_15308,N_14437,N_14890);
nand U15309 (N_15309,N_14886,N_14639);
or U15310 (N_15310,N_14152,N_14528);
or U15311 (N_15311,N_14087,N_14460);
xnor U15312 (N_15312,N_14737,N_14852);
and U15313 (N_15313,N_13781,N_14938);
nand U15314 (N_15314,N_14518,N_14612);
nor U15315 (N_15315,N_14604,N_14782);
and U15316 (N_15316,N_14403,N_14255);
nand U15317 (N_15317,N_14758,N_14073);
nor U15318 (N_15318,N_13852,N_14263);
and U15319 (N_15319,N_13788,N_14423);
nor U15320 (N_15320,N_14043,N_14498);
nand U15321 (N_15321,N_14640,N_14775);
or U15322 (N_15322,N_14526,N_14361);
or U15323 (N_15323,N_13859,N_14454);
and U15324 (N_15324,N_13946,N_13863);
or U15325 (N_15325,N_14784,N_14046);
or U15326 (N_15326,N_14702,N_14369);
or U15327 (N_15327,N_13927,N_14519);
or U15328 (N_15328,N_14193,N_14227);
and U15329 (N_15329,N_13775,N_14843);
xor U15330 (N_15330,N_14653,N_14465);
xnor U15331 (N_15331,N_14130,N_14107);
nor U15332 (N_15332,N_14709,N_14117);
and U15333 (N_15333,N_14165,N_14286);
nor U15334 (N_15334,N_14707,N_14875);
and U15335 (N_15335,N_14280,N_14826);
or U15336 (N_15336,N_14837,N_14746);
nor U15337 (N_15337,N_14968,N_14356);
xor U15338 (N_15338,N_14751,N_14765);
nand U15339 (N_15339,N_14666,N_14489);
nand U15340 (N_15340,N_14659,N_14941);
nand U15341 (N_15341,N_14088,N_14906);
nand U15342 (N_15342,N_14278,N_14094);
xnor U15343 (N_15343,N_14180,N_14930);
xor U15344 (N_15344,N_13924,N_13790);
nor U15345 (N_15345,N_14854,N_13842);
nand U15346 (N_15346,N_14710,N_14743);
or U15347 (N_15347,N_14887,N_14240);
or U15348 (N_15348,N_14367,N_14986);
nor U15349 (N_15349,N_14554,N_14368);
xor U15350 (N_15350,N_13808,N_14964);
or U15351 (N_15351,N_14977,N_14019);
and U15352 (N_15352,N_14218,N_14232);
nor U15353 (N_15353,N_14769,N_14797);
nand U15354 (N_15354,N_14177,N_14619);
nand U15355 (N_15355,N_13849,N_14638);
xor U15356 (N_15356,N_14700,N_13837);
xnor U15357 (N_15357,N_14563,N_14162);
and U15358 (N_15358,N_14223,N_14034);
or U15359 (N_15359,N_14058,N_14776);
xnor U15360 (N_15360,N_14819,N_13964);
xnor U15361 (N_15361,N_14052,N_14950);
nor U15362 (N_15362,N_14032,N_14104);
xnor U15363 (N_15363,N_14802,N_14620);
xor U15364 (N_15364,N_14663,N_13763);
xor U15365 (N_15365,N_14001,N_13819);
nor U15366 (N_15366,N_14587,N_14144);
nand U15367 (N_15367,N_13825,N_14309);
nor U15368 (N_15368,N_14824,N_14200);
nor U15369 (N_15369,N_13812,N_14832);
xnor U15370 (N_15370,N_14348,N_14316);
and U15371 (N_15371,N_13899,N_14158);
xor U15372 (N_15372,N_13937,N_13965);
and U15373 (N_15373,N_14037,N_14015);
or U15374 (N_15374,N_14558,N_14988);
nor U15375 (N_15375,N_14050,N_14074);
or U15376 (N_15376,N_14926,N_14161);
and U15377 (N_15377,N_14167,N_14557);
and U15378 (N_15378,N_13764,N_14476);
nand U15379 (N_15379,N_13921,N_13795);
nor U15380 (N_15380,N_14935,N_14398);
nand U15381 (N_15381,N_14225,N_14678);
xnor U15382 (N_15382,N_14136,N_14883);
or U15383 (N_15383,N_14601,N_14067);
xnor U15384 (N_15384,N_14417,N_14649);
xnor U15385 (N_15385,N_14458,N_14375);
or U15386 (N_15386,N_14182,N_14281);
or U15387 (N_15387,N_14242,N_14967);
or U15388 (N_15388,N_14025,N_14256);
and U15389 (N_15389,N_14980,N_14366);
nor U15390 (N_15390,N_14848,N_14004);
nor U15391 (N_15391,N_14098,N_13991);
or U15392 (N_15392,N_14575,N_14761);
or U15393 (N_15393,N_14116,N_14439);
xnor U15394 (N_15394,N_14389,N_14667);
nand U15395 (N_15395,N_14151,N_14112);
nand U15396 (N_15396,N_14674,N_13782);
nor U15397 (N_15397,N_14485,N_14633);
or U15398 (N_15398,N_13770,N_14827);
nand U15399 (N_15399,N_14084,N_14055);
xor U15400 (N_15400,N_14330,N_14371);
nor U15401 (N_15401,N_14539,N_14672);
and U15402 (N_15402,N_14418,N_14275);
and U15403 (N_15403,N_13952,N_14794);
xnor U15404 (N_15404,N_14501,N_14632);
xor U15405 (N_15405,N_14320,N_14194);
or U15406 (N_15406,N_13776,N_14065);
and U15407 (N_15407,N_14190,N_14801);
or U15408 (N_15408,N_13881,N_14901);
xnor U15409 (N_15409,N_14212,N_14713);
xnor U15410 (N_15410,N_14086,N_13974);
nor U15411 (N_15411,N_13821,N_13923);
or U15412 (N_15412,N_13766,N_14157);
or U15413 (N_15413,N_14265,N_14496);
and U15414 (N_15414,N_13857,N_14952);
or U15415 (N_15415,N_14404,N_14068);
and U15416 (N_15416,N_13767,N_14305);
nand U15417 (N_15417,N_13772,N_13858);
and U15418 (N_15418,N_14833,N_14076);
and U15419 (N_15419,N_14923,N_13878);
nor U15420 (N_15420,N_14047,N_14894);
and U15421 (N_15421,N_14295,N_14215);
nand U15422 (N_15422,N_14277,N_14306);
or U15423 (N_15423,N_14270,N_14310);
and U15424 (N_15424,N_14834,N_13769);
xnor U15425 (N_15425,N_14304,N_14438);
or U15426 (N_15426,N_14317,N_14664);
nand U15427 (N_15427,N_14689,N_13961);
and U15428 (N_15428,N_14231,N_14828);
nand U15429 (N_15429,N_14520,N_14090);
xnor U15430 (N_15430,N_14109,N_13983);
xnor U15431 (N_15431,N_14283,N_14723);
and U15432 (N_15432,N_13771,N_13829);
or U15433 (N_15433,N_13908,N_14129);
nand U15434 (N_15434,N_14990,N_14703);
nand U15435 (N_15435,N_14051,N_13940);
or U15436 (N_15436,N_14509,N_14457);
nand U15437 (N_15437,N_14008,N_14603);
nor U15438 (N_15438,N_14402,N_14137);
nor U15439 (N_15439,N_14279,N_14768);
and U15440 (N_15440,N_14478,N_13866);
and U15441 (N_15441,N_14712,N_13867);
nand U15442 (N_15442,N_14815,N_14462);
nor U15443 (N_15443,N_14753,N_14943);
or U15444 (N_15444,N_14686,N_13818);
nand U15445 (N_15445,N_14805,N_14545);
nand U15446 (N_15446,N_14779,N_14410);
and U15447 (N_15447,N_14029,N_14647);
nand U15448 (N_15448,N_14823,N_13805);
and U15449 (N_15449,N_14795,N_14276);
nor U15450 (N_15450,N_14221,N_14767);
nand U15451 (N_15451,N_14706,N_13935);
and U15452 (N_15452,N_14206,N_14379);
and U15453 (N_15453,N_13932,N_14391);
nand U15454 (N_15454,N_14219,N_14425);
nor U15455 (N_15455,N_14992,N_14038);
or U15456 (N_15456,N_14858,N_14942);
nor U15457 (N_15457,N_14266,N_14507);
xnor U15458 (N_15458,N_14443,N_14506);
or U15459 (N_15459,N_14463,N_14735);
nor U15460 (N_15460,N_14122,N_14291);
and U15461 (N_15461,N_14272,N_14207);
or U15462 (N_15462,N_14188,N_14893);
xnor U15463 (N_15463,N_14159,N_14605);
or U15464 (N_15464,N_14898,N_14170);
nor U15465 (N_15465,N_14658,N_14039);
xnor U15466 (N_15466,N_14975,N_14529);
nor U15467 (N_15467,N_14984,N_13787);
xor U15468 (N_15468,N_14962,N_14504);
nand U15469 (N_15469,N_14042,N_13978);
and U15470 (N_15470,N_14429,N_13813);
nand U15471 (N_15471,N_14237,N_14780);
and U15472 (N_15472,N_14096,N_14960);
nor U15473 (N_15473,N_13943,N_14692);
xor U15474 (N_15474,N_14003,N_14838);
xnor U15475 (N_15475,N_14480,N_13912);
nand U15476 (N_15476,N_14799,N_14989);
nand U15477 (N_15477,N_14956,N_14628);
or U15478 (N_15478,N_13861,N_13773);
nand U15479 (N_15479,N_14993,N_14072);
xor U15480 (N_15480,N_14717,N_14650);
xnor U15481 (N_15481,N_14178,N_14209);
xnor U15482 (N_15482,N_14583,N_14093);
or U15483 (N_15483,N_13887,N_13994);
and U15484 (N_15484,N_14293,N_14774);
or U15485 (N_15485,N_13918,N_14910);
and U15486 (N_15486,N_14850,N_13904);
xor U15487 (N_15487,N_14971,N_14876);
xnor U15488 (N_15488,N_14863,N_14851);
xor U15489 (N_15489,N_14273,N_14127);
nor U15490 (N_15490,N_14933,N_14364);
and U15491 (N_15491,N_14953,N_13931);
or U15492 (N_15492,N_13774,N_14997);
nand U15493 (N_15493,N_14919,N_14830);
xnor U15494 (N_15494,N_13896,N_13864);
nand U15495 (N_15495,N_14119,N_14921);
nand U15496 (N_15496,N_14577,N_14054);
xor U15497 (N_15497,N_14786,N_14424);
and U15498 (N_15498,N_14253,N_14873);
xnor U15499 (N_15499,N_13898,N_14435);
nor U15500 (N_15500,N_13915,N_14831);
or U15501 (N_15501,N_13882,N_14820);
nor U15502 (N_15502,N_13948,N_14588);
xnor U15503 (N_15503,N_14446,N_14613);
xnor U15504 (N_15504,N_13958,N_14024);
or U15505 (N_15505,N_14951,N_13963);
and U15506 (N_15506,N_14998,N_14669);
or U15507 (N_15507,N_13947,N_13957);
nor U15508 (N_15508,N_14101,N_14070);
nand U15509 (N_15509,N_14662,N_14204);
xnor U15510 (N_15510,N_14764,N_13934);
and U15511 (N_15511,N_14315,N_14665);
nand U15512 (N_15512,N_14983,N_14715);
nand U15513 (N_15513,N_14621,N_14825);
xnor U15514 (N_15514,N_14191,N_14773);
xor U15515 (N_15515,N_14214,N_14079);
xor U15516 (N_15516,N_13791,N_14254);
or U15517 (N_15517,N_14083,N_14739);
and U15518 (N_15518,N_14449,N_14156);
nor U15519 (N_15519,N_14724,N_14704);
or U15520 (N_15520,N_14138,N_14721);
or U15521 (N_15521,N_14302,N_14080);
xor U15522 (N_15522,N_13750,N_14475);
or U15523 (N_15523,N_14668,N_14062);
nor U15524 (N_15524,N_13760,N_13893);
nand U15525 (N_15525,N_14262,N_14682);
or U15526 (N_15526,N_14113,N_14755);
and U15527 (N_15527,N_14334,N_14907);
nand U15528 (N_15528,N_13783,N_14616);
nand U15529 (N_15529,N_14803,N_14483);
nand U15530 (N_15530,N_13853,N_14835);
or U15531 (N_15531,N_13980,N_14934);
xor U15532 (N_15532,N_14082,N_14688);
nand U15533 (N_15533,N_14566,N_14740);
nand U15534 (N_15534,N_13814,N_14491);
xnor U15535 (N_15535,N_14772,N_14582);
and U15536 (N_15536,N_14377,N_13793);
xor U15537 (N_15537,N_13765,N_14331);
nand U15538 (N_15538,N_14114,N_14562);
xor U15539 (N_15539,N_14542,N_14781);
or U15540 (N_15540,N_13903,N_14937);
or U15541 (N_15541,N_14798,N_14513);
or U15542 (N_15542,N_14576,N_14172);
and U15543 (N_15543,N_14862,N_14102);
nor U15544 (N_15544,N_14687,N_14477);
or U15545 (N_15545,N_14271,N_14228);
nand U15546 (N_15546,N_14405,N_14708);
and U15547 (N_15547,N_14342,N_13884);
and U15548 (N_15548,N_14380,N_14760);
nor U15549 (N_15549,N_14573,N_14592);
nand U15550 (N_15550,N_14396,N_14839);
or U15551 (N_15551,N_14729,N_14745);
or U15552 (N_15552,N_14537,N_14900);
xor U15553 (N_15553,N_14325,N_13827);
nand U15554 (N_15554,N_14915,N_14608);
nor U15555 (N_15555,N_14564,N_14468);
nand U15556 (N_15556,N_13845,N_14143);
and U15557 (N_15557,N_14282,N_14142);
nand U15558 (N_15558,N_14345,N_14512);
nand U15559 (N_15559,N_14584,N_14386);
and U15560 (N_15560,N_13801,N_13847);
nor U15561 (N_15561,N_13822,N_14548);
nand U15562 (N_15562,N_14732,N_14314);
xnor U15563 (N_15563,N_14044,N_13880);
xnor U15564 (N_15564,N_14618,N_13977);
nor U15565 (N_15565,N_14217,N_14360);
nand U15566 (N_15566,N_14021,N_14376);
and U15567 (N_15567,N_14924,N_14097);
or U15568 (N_15568,N_14185,N_13778);
xnor U15569 (N_15569,N_14572,N_14845);
or U15570 (N_15570,N_14409,N_14236);
and U15571 (N_15571,N_14069,N_14005);
or U15572 (N_15572,N_13780,N_14626);
and U15573 (N_15573,N_13802,N_13865);
nor U15574 (N_15574,N_14866,N_14614);
nand U15575 (N_15575,N_14422,N_14979);
and U15576 (N_15576,N_14840,N_14580);
or U15577 (N_15577,N_14870,N_13768);
and U15578 (N_15578,N_13807,N_14999);
xor U15579 (N_15579,N_14969,N_14742);
xnor U15580 (N_15580,N_14762,N_14521);
or U15581 (N_15581,N_14230,N_14913);
or U15582 (N_15582,N_14472,N_14982);
or U15583 (N_15583,N_13966,N_14757);
nand U15584 (N_15584,N_14049,N_14565);
nor U15585 (N_15585,N_13962,N_14020);
nor U15586 (N_15586,N_14738,N_14695);
or U15587 (N_15587,N_14918,N_14609);
and U15588 (N_15588,N_14181,N_14581);
nand U15589 (N_15589,N_14346,N_14897);
xor U15590 (N_15590,N_14323,N_14064);
xor U15591 (N_15591,N_14099,N_14192);
xnor U15592 (N_15592,N_14235,N_14041);
nand U15593 (N_15593,N_13759,N_14022);
nor U15594 (N_15594,N_14146,N_13796);
or U15595 (N_15595,N_14966,N_14328);
xor U15596 (N_15596,N_14598,N_13800);
nand U15597 (N_15597,N_13879,N_14586);
and U15598 (N_15598,N_14804,N_14970);
nor U15599 (N_15599,N_14179,N_14777);
xnor U15600 (N_15600,N_14644,N_14556);
or U15601 (N_15601,N_14841,N_14800);
nand U15602 (N_15602,N_14350,N_14289);
or U15603 (N_15603,N_14976,N_14441);
or U15604 (N_15604,N_13806,N_13911);
and U15605 (N_15605,N_14654,N_14677);
nand U15606 (N_15606,N_14250,N_13761);
or U15607 (N_15607,N_14164,N_14974);
nand U15608 (N_15608,N_13844,N_14408);
and U15609 (N_15609,N_14089,N_13848);
and U15610 (N_15610,N_14903,N_14756);
and U15611 (N_15611,N_13955,N_13786);
and U15612 (N_15612,N_14173,N_14810);
and U15613 (N_15613,N_14354,N_14095);
xor U15614 (N_15614,N_14294,N_14916);
and U15615 (N_15615,N_14184,N_14487);
and U15616 (N_15616,N_14481,N_14711);
nand U15617 (N_15617,N_14243,N_14340);
and U15618 (N_15618,N_14759,N_14912);
xor U15619 (N_15619,N_14972,N_14499);
nand U15620 (N_15620,N_14428,N_14589);
nand U15621 (N_15621,N_14495,N_14464);
nand U15622 (N_15622,N_14053,N_14002);
or U15623 (N_15623,N_14948,N_14954);
and U15624 (N_15624,N_14809,N_14533);
or U15625 (N_15625,N_14447,N_14751);
and U15626 (N_15626,N_14293,N_14958);
and U15627 (N_15627,N_14506,N_14617);
xnor U15628 (N_15628,N_14714,N_14822);
xnor U15629 (N_15629,N_14723,N_14807);
nand U15630 (N_15630,N_14123,N_14735);
and U15631 (N_15631,N_14073,N_14502);
nand U15632 (N_15632,N_14889,N_14016);
and U15633 (N_15633,N_14965,N_13878);
or U15634 (N_15634,N_14727,N_14299);
xor U15635 (N_15635,N_14274,N_14577);
nand U15636 (N_15636,N_14108,N_14152);
or U15637 (N_15637,N_13961,N_14718);
xor U15638 (N_15638,N_14362,N_14791);
nor U15639 (N_15639,N_14741,N_14102);
nand U15640 (N_15640,N_14242,N_14394);
and U15641 (N_15641,N_14371,N_14229);
xor U15642 (N_15642,N_13874,N_14163);
xor U15643 (N_15643,N_14515,N_13859);
nor U15644 (N_15644,N_13985,N_14589);
nor U15645 (N_15645,N_14699,N_14577);
xor U15646 (N_15646,N_13912,N_14157);
nand U15647 (N_15647,N_14027,N_14654);
nor U15648 (N_15648,N_14653,N_14228);
or U15649 (N_15649,N_14072,N_14021);
or U15650 (N_15650,N_13927,N_14059);
or U15651 (N_15651,N_13821,N_13838);
nand U15652 (N_15652,N_14449,N_14732);
or U15653 (N_15653,N_13824,N_14677);
xnor U15654 (N_15654,N_13946,N_14322);
or U15655 (N_15655,N_14903,N_14437);
and U15656 (N_15656,N_14683,N_14649);
nand U15657 (N_15657,N_14309,N_14639);
xnor U15658 (N_15658,N_14915,N_14600);
nor U15659 (N_15659,N_14209,N_14083);
nand U15660 (N_15660,N_13890,N_14633);
nand U15661 (N_15661,N_14787,N_14166);
xnor U15662 (N_15662,N_14011,N_14057);
and U15663 (N_15663,N_14205,N_14039);
and U15664 (N_15664,N_14200,N_14873);
nor U15665 (N_15665,N_14646,N_14407);
xor U15666 (N_15666,N_14338,N_14824);
nand U15667 (N_15667,N_14593,N_13767);
nand U15668 (N_15668,N_13935,N_14378);
nor U15669 (N_15669,N_14082,N_14077);
and U15670 (N_15670,N_14795,N_13940);
or U15671 (N_15671,N_14506,N_14955);
or U15672 (N_15672,N_14466,N_14354);
xor U15673 (N_15673,N_14434,N_14616);
xnor U15674 (N_15674,N_14461,N_14573);
and U15675 (N_15675,N_14322,N_14258);
nand U15676 (N_15676,N_14326,N_14402);
and U15677 (N_15677,N_14578,N_14424);
nand U15678 (N_15678,N_14935,N_14567);
and U15679 (N_15679,N_14391,N_13907);
and U15680 (N_15680,N_14365,N_14954);
and U15681 (N_15681,N_14603,N_14325);
and U15682 (N_15682,N_14367,N_14875);
and U15683 (N_15683,N_13871,N_14839);
and U15684 (N_15684,N_14862,N_14242);
or U15685 (N_15685,N_14719,N_14761);
and U15686 (N_15686,N_14192,N_14309);
and U15687 (N_15687,N_14522,N_13765);
and U15688 (N_15688,N_14206,N_13818);
nand U15689 (N_15689,N_14388,N_14679);
xor U15690 (N_15690,N_14764,N_14830);
nor U15691 (N_15691,N_14655,N_14752);
and U15692 (N_15692,N_14176,N_14533);
nor U15693 (N_15693,N_14308,N_14807);
xnor U15694 (N_15694,N_13979,N_14364);
or U15695 (N_15695,N_14550,N_14315);
or U15696 (N_15696,N_14560,N_14647);
nor U15697 (N_15697,N_14893,N_14510);
or U15698 (N_15698,N_14778,N_13908);
and U15699 (N_15699,N_14577,N_13770);
or U15700 (N_15700,N_14271,N_14810);
nand U15701 (N_15701,N_14255,N_14851);
or U15702 (N_15702,N_14921,N_14774);
or U15703 (N_15703,N_14209,N_14650);
and U15704 (N_15704,N_14153,N_13988);
and U15705 (N_15705,N_13806,N_14209);
nand U15706 (N_15706,N_13793,N_14825);
nand U15707 (N_15707,N_13927,N_14022);
nand U15708 (N_15708,N_14041,N_14307);
or U15709 (N_15709,N_14879,N_13882);
nor U15710 (N_15710,N_14589,N_14572);
xnor U15711 (N_15711,N_14614,N_14607);
nor U15712 (N_15712,N_14481,N_14065);
or U15713 (N_15713,N_14534,N_14066);
xor U15714 (N_15714,N_14048,N_13941);
nand U15715 (N_15715,N_14059,N_13916);
nand U15716 (N_15716,N_13912,N_14169);
or U15717 (N_15717,N_14424,N_14004);
and U15718 (N_15718,N_14551,N_14848);
nand U15719 (N_15719,N_14044,N_14219);
and U15720 (N_15720,N_14851,N_14090);
or U15721 (N_15721,N_14416,N_14636);
xor U15722 (N_15722,N_14304,N_14892);
nand U15723 (N_15723,N_14172,N_14443);
xnor U15724 (N_15724,N_14232,N_14906);
nor U15725 (N_15725,N_13813,N_14784);
or U15726 (N_15726,N_14648,N_14206);
xnor U15727 (N_15727,N_14931,N_14079);
and U15728 (N_15728,N_14614,N_14413);
nor U15729 (N_15729,N_14505,N_14381);
xnor U15730 (N_15730,N_14153,N_14527);
nor U15731 (N_15731,N_14020,N_14764);
and U15732 (N_15732,N_14909,N_14583);
xnor U15733 (N_15733,N_14093,N_14783);
or U15734 (N_15734,N_14152,N_14300);
or U15735 (N_15735,N_14765,N_14381);
nor U15736 (N_15736,N_14336,N_14409);
and U15737 (N_15737,N_14478,N_14520);
or U15738 (N_15738,N_14381,N_14955);
and U15739 (N_15739,N_14299,N_13955);
xor U15740 (N_15740,N_14130,N_14359);
and U15741 (N_15741,N_14868,N_14221);
nor U15742 (N_15742,N_14186,N_14035);
nand U15743 (N_15743,N_14505,N_13862);
nand U15744 (N_15744,N_14100,N_14732);
nor U15745 (N_15745,N_14732,N_14844);
nor U15746 (N_15746,N_14619,N_14373);
xnor U15747 (N_15747,N_14861,N_13898);
nor U15748 (N_15748,N_14572,N_13791);
xnor U15749 (N_15749,N_13845,N_14610);
nand U15750 (N_15750,N_14441,N_14526);
and U15751 (N_15751,N_13954,N_14778);
and U15752 (N_15752,N_13978,N_14610);
nand U15753 (N_15753,N_14568,N_14661);
nand U15754 (N_15754,N_14211,N_14108);
nor U15755 (N_15755,N_13993,N_14011);
nor U15756 (N_15756,N_14947,N_14836);
and U15757 (N_15757,N_14564,N_14347);
or U15758 (N_15758,N_14832,N_14718);
nor U15759 (N_15759,N_14849,N_13907);
nand U15760 (N_15760,N_13774,N_14489);
xor U15761 (N_15761,N_13777,N_13893);
nor U15762 (N_15762,N_13850,N_13804);
xnor U15763 (N_15763,N_13899,N_14781);
or U15764 (N_15764,N_14381,N_14400);
nand U15765 (N_15765,N_14629,N_14930);
xor U15766 (N_15766,N_14673,N_13943);
or U15767 (N_15767,N_14338,N_14538);
xor U15768 (N_15768,N_14391,N_13984);
or U15769 (N_15769,N_14633,N_14601);
xor U15770 (N_15770,N_14037,N_14095);
nor U15771 (N_15771,N_14806,N_13941);
xnor U15772 (N_15772,N_14822,N_13930);
or U15773 (N_15773,N_13780,N_14323);
and U15774 (N_15774,N_14381,N_14624);
nor U15775 (N_15775,N_14957,N_14109);
xor U15776 (N_15776,N_13816,N_14757);
and U15777 (N_15777,N_14645,N_14320);
nand U15778 (N_15778,N_14240,N_14985);
nor U15779 (N_15779,N_14242,N_14218);
or U15780 (N_15780,N_13953,N_14097);
xor U15781 (N_15781,N_13925,N_14695);
xnor U15782 (N_15782,N_14596,N_14526);
xor U15783 (N_15783,N_14380,N_14059);
or U15784 (N_15784,N_14594,N_14966);
xnor U15785 (N_15785,N_14106,N_14472);
xnor U15786 (N_15786,N_14531,N_14366);
nand U15787 (N_15787,N_14887,N_14354);
nor U15788 (N_15788,N_14122,N_14499);
and U15789 (N_15789,N_14614,N_13867);
nand U15790 (N_15790,N_14526,N_14284);
and U15791 (N_15791,N_14747,N_13757);
xnor U15792 (N_15792,N_13829,N_14645);
nor U15793 (N_15793,N_13962,N_14848);
xor U15794 (N_15794,N_13829,N_14416);
or U15795 (N_15795,N_14436,N_14743);
and U15796 (N_15796,N_13898,N_13855);
xnor U15797 (N_15797,N_14582,N_13804);
nand U15798 (N_15798,N_13995,N_14964);
nand U15799 (N_15799,N_13783,N_14248);
and U15800 (N_15800,N_14223,N_14619);
or U15801 (N_15801,N_14235,N_14557);
or U15802 (N_15802,N_14067,N_13870);
and U15803 (N_15803,N_14630,N_14749);
or U15804 (N_15804,N_13989,N_14806);
nor U15805 (N_15805,N_14757,N_14878);
nand U15806 (N_15806,N_14272,N_14364);
nand U15807 (N_15807,N_13854,N_14515);
nand U15808 (N_15808,N_14155,N_14572);
and U15809 (N_15809,N_14660,N_14823);
or U15810 (N_15810,N_14641,N_14851);
xnor U15811 (N_15811,N_13873,N_13972);
nor U15812 (N_15812,N_13979,N_14834);
and U15813 (N_15813,N_14406,N_14525);
xor U15814 (N_15814,N_13854,N_14757);
nand U15815 (N_15815,N_13897,N_13910);
xnor U15816 (N_15816,N_14742,N_13799);
nor U15817 (N_15817,N_13870,N_14788);
nand U15818 (N_15818,N_14381,N_14617);
or U15819 (N_15819,N_13807,N_14934);
and U15820 (N_15820,N_14144,N_14020);
nand U15821 (N_15821,N_14717,N_14413);
nand U15822 (N_15822,N_14814,N_14759);
nor U15823 (N_15823,N_14251,N_14587);
nand U15824 (N_15824,N_14455,N_14177);
nor U15825 (N_15825,N_14024,N_14772);
xnor U15826 (N_15826,N_14746,N_14221);
nand U15827 (N_15827,N_14953,N_14558);
nor U15828 (N_15828,N_14511,N_14977);
or U15829 (N_15829,N_14511,N_14502);
nor U15830 (N_15830,N_14995,N_14657);
and U15831 (N_15831,N_14465,N_14831);
or U15832 (N_15832,N_14308,N_14350);
and U15833 (N_15833,N_13981,N_14571);
xor U15834 (N_15834,N_14010,N_14118);
xnor U15835 (N_15835,N_13977,N_14887);
xnor U15836 (N_15836,N_14677,N_14499);
xor U15837 (N_15837,N_14457,N_14093);
nand U15838 (N_15838,N_14504,N_13944);
nand U15839 (N_15839,N_14854,N_14282);
xnor U15840 (N_15840,N_13845,N_14795);
nor U15841 (N_15841,N_14122,N_14892);
nand U15842 (N_15842,N_14529,N_14983);
and U15843 (N_15843,N_13962,N_14898);
or U15844 (N_15844,N_14430,N_14118);
xnor U15845 (N_15845,N_13924,N_14905);
or U15846 (N_15846,N_14983,N_14212);
nor U15847 (N_15847,N_13928,N_14531);
and U15848 (N_15848,N_14043,N_14917);
or U15849 (N_15849,N_13754,N_13856);
and U15850 (N_15850,N_14414,N_13929);
nand U15851 (N_15851,N_14684,N_14162);
nand U15852 (N_15852,N_14169,N_14811);
nor U15853 (N_15853,N_14674,N_14654);
xor U15854 (N_15854,N_13817,N_13916);
nor U15855 (N_15855,N_14252,N_13911);
nor U15856 (N_15856,N_13880,N_14917);
nor U15857 (N_15857,N_14048,N_14228);
nand U15858 (N_15858,N_14164,N_14896);
nor U15859 (N_15859,N_14191,N_14733);
nor U15860 (N_15860,N_13827,N_14163);
or U15861 (N_15861,N_14002,N_14948);
nor U15862 (N_15862,N_14777,N_14626);
or U15863 (N_15863,N_14999,N_14613);
xnor U15864 (N_15864,N_13922,N_14268);
nand U15865 (N_15865,N_14194,N_13905);
and U15866 (N_15866,N_14726,N_13823);
nand U15867 (N_15867,N_14889,N_14287);
or U15868 (N_15868,N_14943,N_14642);
and U15869 (N_15869,N_13854,N_14256);
nor U15870 (N_15870,N_13791,N_14205);
nand U15871 (N_15871,N_14044,N_14707);
nor U15872 (N_15872,N_14235,N_14591);
or U15873 (N_15873,N_14122,N_14317);
xor U15874 (N_15874,N_14802,N_13878);
nand U15875 (N_15875,N_14123,N_14243);
or U15876 (N_15876,N_14644,N_14961);
nand U15877 (N_15877,N_13802,N_14832);
or U15878 (N_15878,N_13826,N_14716);
and U15879 (N_15879,N_13901,N_14309);
and U15880 (N_15880,N_14153,N_14978);
or U15881 (N_15881,N_13970,N_14422);
or U15882 (N_15882,N_14373,N_14534);
xor U15883 (N_15883,N_13840,N_14229);
nand U15884 (N_15884,N_14292,N_14164);
nand U15885 (N_15885,N_14643,N_14381);
nor U15886 (N_15886,N_14582,N_14558);
xnor U15887 (N_15887,N_14759,N_14935);
xnor U15888 (N_15888,N_14171,N_14999);
and U15889 (N_15889,N_14037,N_14918);
nor U15890 (N_15890,N_14905,N_14619);
or U15891 (N_15891,N_14272,N_14210);
nand U15892 (N_15892,N_14110,N_14957);
nand U15893 (N_15893,N_13837,N_14724);
nand U15894 (N_15894,N_13990,N_14910);
nand U15895 (N_15895,N_14555,N_13898);
xnor U15896 (N_15896,N_13769,N_14047);
and U15897 (N_15897,N_14748,N_14274);
nand U15898 (N_15898,N_14213,N_14124);
xor U15899 (N_15899,N_14378,N_13802);
and U15900 (N_15900,N_14101,N_14376);
nor U15901 (N_15901,N_14596,N_14018);
nand U15902 (N_15902,N_14129,N_14960);
nor U15903 (N_15903,N_14392,N_14509);
xnor U15904 (N_15904,N_14666,N_14598);
or U15905 (N_15905,N_14695,N_14816);
nor U15906 (N_15906,N_14709,N_13869);
and U15907 (N_15907,N_14460,N_14528);
nor U15908 (N_15908,N_14460,N_14424);
and U15909 (N_15909,N_14462,N_14977);
nor U15910 (N_15910,N_14286,N_14313);
or U15911 (N_15911,N_14179,N_14106);
and U15912 (N_15912,N_14910,N_14427);
and U15913 (N_15913,N_14608,N_13843);
nand U15914 (N_15914,N_14937,N_14352);
and U15915 (N_15915,N_14038,N_14545);
nand U15916 (N_15916,N_13847,N_14242);
and U15917 (N_15917,N_14787,N_14089);
nand U15918 (N_15918,N_13904,N_14098);
and U15919 (N_15919,N_14253,N_14146);
nand U15920 (N_15920,N_14653,N_13863);
nand U15921 (N_15921,N_14873,N_14912);
nor U15922 (N_15922,N_13982,N_14023);
or U15923 (N_15923,N_13893,N_14855);
nand U15924 (N_15924,N_14694,N_14781);
xnor U15925 (N_15925,N_14975,N_14979);
or U15926 (N_15926,N_13997,N_13938);
or U15927 (N_15927,N_14074,N_14334);
nor U15928 (N_15928,N_14973,N_13816);
and U15929 (N_15929,N_14143,N_13965);
xnor U15930 (N_15930,N_14035,N_14522);
nor U15931 (N_15931,N_14049,N_14478);
or U15932 (N_15932,N_14749,N_13755);
and U15933 (N_15933,N_14408,N_14709);
xor U15934 (N_15934,N_13839,N_14372);
and U15935 (N_15935,N_14398,N_14415);
or U15936 (N_15936,N_14956,N_14915);
nor U15937 (N_15937,N_14697,N_14388);
nand U15938 (N_15938,N_14828,N_14454);
and U15939 (N_15939,N_13962,N_14002);
xor U15940 (N_15940,N_14300,N_14493);
nor U15941 (N_15941,N_13824,N_14661);
nand U15942 (N_15942,N_14659,N_13861);
xnor U15943 (N_15943,N_14681,N_14156);
xnor U15944 (N_15944,N_13782,N_14666);
or U15945 (N_15945,N_14126,N_14210);
xnor U15946 (N_15946,N_13757,N_14391);
xor U15947 (N_15947,N_14179,N_14933);
nand U15948 (N_15948,N_14519,N_14692);
or U15949 (N_15949,N_14131,N_14565);
xnor U15950 (N_15950,N_14676,N_13827);
nor U15951 (N_15951,N_14899,N_14556);
or U15952 (N_15952,N_14951,N_14829);
or U15953 (N_15953,N_14753,N_14320);
nor U15954 (N_15954,N_14787,N_13930);
nand U15955 (N_15955,N_14105,N_13936);
or U15956 (N_15956,N_14237,N_13980);
nor U15957 (N_15957,N_13831,N_14298);
nand U15958 (N_15958,N_14679,N_14851);
and U15959 (N_15959,N_13753,N_13795);
nor U15960 (N_15960,N_14920,N_14993);
nor U15961 (N_15961,N_14688,N_14049);
nor U15962 (N_15962,N_13989,N_14781);
or U15963 (N_15963,N_14586,N_14205);
and U15964 (N_15964,N_14570,N_13952);
xor U15965 (N_15965,N_13890,N_14673);
nor U15966 (N_15966,N_14179,N_14006);
nand U15967 (N_15967,N_14989,N_14734);
or U15968 (N_15968,N_14476,N_14941);
nor U15969 (N_15969,N_14839,N_14562);
and U15970 (N_15970,N_14955,N_13904);
and U15971 (N_15971,N_14940,N_14107);
nor U15972 (N_15972,N_13899,N_14223);
or U15973 (N_15973,N_14648,N_13997);
nor U15974 (N_15974,N_14627,N_14719);
xnor U15975 (N_15975,N_14731,N_13845);
nor U15976 (N_15976,N_14183,N_13931);
nand U15977 (N_15977,N_13753,N_14398);
or U15978 (N_15978,N_14796,N_14369);
xnor U15979 (N_15979,N_14174,N_13987);
or U15980 (N_15980,N_14822,N_14674);
and U15981 (N_15981,N_14694,N_14851);
nor U15982 (N_15982,N_14240,N_14069);
xnor U15983 (N_15983,N_14204,N_14153);
and U15984 (N_15984,N_14694,N_14795);
or U15985 (N_15985,N_14040,N_14737);
nand U15986 (N_15986,N_14577,N_14434);
and U15987 (N_15987,N_14870,N_14584);
nand U15988 (N_15988,N_14779,N_14706);
or U15989 (N_15989,N_14523,N_14071);
nand U15990 (N_15990,N_14851,N_13993);
and U15991 (N_15991,N_14325,N_14979);
xnor U15992 (N_15992,N_13835,N_14689);
and U15993 (N_15993,N_14815,N_14077);
nand U15994 (N_15994,N_13962,N_14488);
or U15995 (N_15995,N_14241,N_14152);
and U15996 (N_15996,N_14810,N_14635);
nor U15997 (N_15997,N_14927,N_14659);
nor U15998 (N_15998,N_13811,N_14686);
or U15999 (N_15999,N_14959,N_14142);
nand U16000 (N_16000,N_14502,N_14596);
nor U16001 (N_16001,N_14000,N_14219);
or U16002 (N_16002,N_14711,N_13765);
nor U16003 (N_16003,N_14602,N_14368);
xor U16004 (N_16004,N_14016,N_14002);
and U16005 (N_16005,N_14371,N_13975);
nand U16006 (N_16006,N_14125,N_13897);
xnor U16007 (N_16007,N_14656,N_14460);
nor U16008 (N_16008,N_14716,N_13872);
and U16009 (N_16009,N_13873,N_14823);
nand U16010 (N_16010,N_13826,N_14278);
nor U16011 (N_16011,N_14235,N_14694);
xnor U16012 (N_16012,N_13766,N_14464);
and U16013 (N_16013,N_14197,N_13972);
xor U16014 (N_16014,N_14400,N_14260);
nor U16015 (N_16015,N_14563,N_14650);
or U16016 (N_16016,N_14609,N_14262);
or U16017 (N_16017,N_14057,N_14117);
nand U16018 (N_16018,N_14490,N_14815);
or U16019 (N_16019,N_14545,N_14885);
nand U16020 (N_16020,N_14544,N_14591);
and U16021 (N_16021,N_14615,N_14158);
xnor U16022 (N_16022,N_14810,N_14291);
and U16023 (N_16023,N_14332,N_14226);
nor U16024 (N_16024,N_14847,N_14917);
and U16025 (N_16025,N_13807,N_13987);
xor U16026 (N_16026,N_13860,N_14625);
or U16027 (N_16027,N_13813,N_14761);
xor U16028 (N_16028,N_14182,N_14747);
nor U16029 (N_16029,N_13900,N_13955);
and U16030 (N_16030,N_13988,N_14530);
nand U16031 (N_16031,N_14356,N_14485);
or U16032 (N_16032,N_14981,N_14248);
or U16033 (N_16033,N_14724,N_14885);
xnor U16034 (N_16034,N_14987,N_14677);
and U16035 (N_16035,N_14826,N_14078);
or U16036 (N_16036,N_14963,N_14116);
xor U16037 (N_16037,N_14657,N_14359);
xnor U16038 (N_16038,N_14319,N_14951);
nor U16039 (N_16039,N_14292,N_14050);
nor U16040 (N_16040,N_14351,N_13918);
or U16041 (N_16041,N_13901,N_14219);
nand U16042 (N_16042,N_14878,N_13985);
xnor U16043 (N_16043,N_14636,N_14706);
nor U16044 (N_16044,N_14923,N_14847);
or U16045 (N_16045,N_13871,N_14537);
nand U16046 (N_16046,N_14992,N_14563);
or U16047 (N_16047,N_14608,N_13831);
nand U16048 (N_16048,N_14365,N_13812);
or U16049 (N_16049,N_14277,N_14246);
nor U16050 (N_16050,N_14972,N_14593);
nor U16051 (N_16051,N_14608,N_14536);
or U16052 (N_16052,N_14743,N_13831);
xnor U16053 (N_16053,N_13894,N_14497);
xor U16054 (N_16054,N_14469,N_14017);
and U16055 (N_16055,N_14911,N_14255);
or U16056 (N_16056,N_14921,N_14952);
nand U16057 (N_16057,N_14893,N_14628);
nand U16058 (N_16058,N_14081,N_14676);
and U16059 (N_16059,N_13942,N_14841);
or U16060 (N_16060,N_14498,N_13755);
nand U16061 (N_16061,N_14058,N_14668);
nand U16062 (N_16062,N_14316,N_14261);
nand U16063 (N_16063,N_13883,N_14247);
and U16064 (N_16064,N_14595,N_14264);
nor U16065 (N_16065,N_14096,N_14074);
nand U16066 (N_16066,N_14888,N_14903);
and U16067 (N_16067,N_14977,N_14221);
nand U16068 (N_16068,N_14142,N_14104);
and U16069 (N_16069,N_14645,N_14440);
nand U16070 (N_16070,N_14118,N_14319);
or U16071 (N_16071,N_14116,N_14859);
nor U16072 (N_16072,N_14208,N_14385);
nand U16073 (N_16073,N_14701,N_13994);
or U16074 (N_16074,N_14288,N_14129);
nor U16075 (N_16075,N_14742,N_14210);
or U16076 (N_16076,N_14760,N_14097);
nand U16077 (N_16077,N_14800,N_13798);
nor U16078 (N_16078,N_13979,N_14286);
xor U16079 (N_16079,N_13886,N_14096);
and U16080 (N_16080,N_14310,N_14518);
nor U16081 (N_16081,N_14613,N_14108);
nand U16082 (N_16082,N_14130,N_14218);
or U16083 (N_16083,N_14888,N_14441);
nor U16084 (N_16084,N_13783,N_14020);
xnor U16085 (N_16085,N_14953,N_14189);
nand U16086 (N_16086,N_14003,N_13791);
or U16087 (N_16087,N_13897,N_14102);
and U16088 (N_16088,N_14268,N_14381);
and U16089 (N_16089,N_14830,N_14940);
nand U16090 (N_16090,N_13826,N_14295);
or U16091 (N_16091,N_14917,N_14126);
nor U16092 (N_16092,N_13868,N_14294);
nand U16093 (N_16093,N_14622,N_14370);
nand U16094 (N_16094,N_13754,N_14924);
and U16095 (N_16095,N_13825,N_14544);
and U16096 (N_16096,N_14671,N_13759);
nand U16097 (N_16097,N_14285,N_14859);
nand U16098 (N_16098,N_14596,N_14036);
nor U16099 (N_16099,N_14342,N_14571);
nor U16100 (N_16100,N_14170,N_14607);
and U16101 (N_16101,N_14484,N_14990);
xor U16102 (N_16102,N_14836,N_14610);
xnor U16103 (N_16103,N_14615,N_14144);
and U16104 (N_16104,N_13816,N_14763);
nor U16105 (N_16105,N_14775,N_14680);
and U16106 (N_16106,N_14001,N_14814);
or U16107 (N_16107,N_14590,N_14129);
nor U16108 (N_16108,N_14546,N_14146);
and U16109 (N_16109,N_14218,N_14608);
and U16110 (N_16110,N_14741,N_14987);
xnor U16111 (N_16111,N_14285,N_14019);
nand U16112 (N_16112,N_14721,N_13860);
xnor U16113 (N_16113,N_14886,N_14122);
xnor U16114 (N_16114,N_14080,N_13880);
nor U16115 (N_16115,N_14657,N_14894);
xor U16116 (N_16116,N_14201,N_14653);
nor U16117 (N_16117,N_14977,N_14072);
or U16118 (N_16118,N_14096,N_14720);
nor U16119 (N_16119,N_14290,N_14829);
xnor U16120 (N_16120,N_14168,N_13985);
and U16121 (N_16121,N_14456,N_13918);
xor U16122 (N_16122,N_13977,N_14373);
xnor U16123 (N_16123,N_14605,N_14737);
or U16124 (N_16124,N_14256,N_14888);
xnor U16125 (N_16125,N_14872,N_14108);
nand U16126 (N_16126,N_14132,N_14978);
xor U16127 (N_16127,N_14705,N_14089);
xor U16128 (N_16128,N_13878,N_14524);
or U16129 (N_16129,N_14282,N_13809);
xor U16130 (N_16130,N_14350,N_14270);
xnor U16131 (N_16131,N_13811,N_14371);
or U16132 (N_16132,N_14865,N_14543);
or U16133 (N_16133,N_14472,N_14414);
xnor U16134 (N_16134,N_14210,N_14761);
or U16135 (N_16135,N_14646,N_13958);
nor U16136 (N_16136,N_14907,N_14011);
and U16137 (N_16137,N_14429,N_14357);
nor U16138 (N_16138,N_14435,N_14499);
xor U16139 (N_16139,N_14268,N_14004);
nand U16140 (N_16140,N_14907,N_14290);
nor U16141 (N_16141,N_14523,N_14719);
or U16142 (N_16142,N_14270,N_14502);
or U16143 (N_16143,N_13814,N_14831);
nand U16144 (N_16144,N_13818,N_14825);
or U16145 (N_16145,N_13832,N_13800);
nand U16146 (N_16146,N_13826,N_13937);
and U16147 (N_16147,N_14818,N_14946);
or U16148 (N_16148,N_13919,N_14211);
or U16149 (N_16149,N_14160,N_14055);
nand U16150 (N_16150,N_14839,N_14823);
nand U16151 (N_16151,N_14541,N_14575);
or U16152 (N_16152,N_14757,N_14402);
nor U16153 (N_16153,N_14433,N_14862);
nor U16154 (N_16154,N_14765,N_14998);
or U16155 (N_16155,N_13838,N_13940);
nor U16156 (N_16156,N_14044,N_14171);
xnor U16157 (N_16157,N_14883,N_14091);
xnor U16158 (N_16158,N_14868,N_14325);
nand U16159 (N_16159,N_14828,N_14378);
or U16160 (N_16160,N_14876,N_13917);
nand U16161 (N_16161,N_14908,N_13840);
or U16162 (N_16162,N_13840,N_13921);
or U16163 (N_16163,N_14377,N_13983);
and U16164 (N_16164,N_14351,N_13857);
nand U16165 (N_16165,N_14912,N_13871);
xor U16166 (N_16166,N_14803,N_13865);
and U16167 (N_16167,N_14961,N_14251);
or U16168 (N_16168,N_13854,N_13755);
xnor U16169 (N_16169,N_14389,N_14677);
and U16170 (N_16170,N_14109,N_14885);
nor U16171 (N_16171,N_14916,N_14204);
nor U16172 (N_16172,N_14375,N_14394);
xor U16173 (N_16173,N_14230,N_14596);
nand U16174 (N_16174,N_14704,N_14707);
or U16175 (N_16175,N_14460,N_13839);
nand U16176 (N_16176,N_14664,N_14014);
or U16177 (N_16177,N_14104,N_14929);
nand U16178 (N_16178,N_14379,N_14293);
or U16179 (N_16179,N_14903,N_14067);
nor U16180 (N_16180,N_14486,N_14389);
nor U16181 (N_16181,N_14624,N_14574);
nand U16182 (N_16182,N_14293,N_14690);
xor U16183 (N_16183,N_13919,N_14353);
nor U16184 (N_16184,N_14833,N_14366);
or U16185 (N_16185,N_14281,N_14097);
nand U16186 (N_16186,N_14026,N_13806);
and U16187 (N_16187,N_14211,N_13927);
nand U16188 (N_16188,N_14190,N_14422);
and U16189 (N_16189,N_13779,N_14368);
xor U16190 (N_16190,N_14450,N_14339);
xor U16191 (N_16191,N_14112,N_14770);
nor U16192 (N_16192,N_14723,N_14095);
nand U16193 (N_16193,N_13768,N_14749);
or U16194 (N_16194,N_14272,N_14751);
nand U16195 (N_16195,N_14995,N_14745);
nand U16196 (N_16196,N_14854,N_14547);
nand U16197 (N_16197,N_14295,N_14898);
nor U16198 (N_16198,N_14375,N_14853);
xor U16199 (N_16199,N_14299,N_14528);
nand U16200 (N_16200,N_13925,N_14562);
nor U16201 (N_16201,N_14267,N_14375);
xnor U16202 (N_16202,N_14479,N_14066);
and U16203 (N_16203,N_14643,N_13832);
nand U16204 (N_16204,N_14759,N_14355);
nor U16205 (N_16205,N_14739,N_14815);
nor U16206 (N_16206,N_14539,N_14465);
xor U16207 (N_16207,N_13840,N_13872);
nor U16208 (N_16208,N_13787,N_14641);
xnor U16209 (N_16209,N_14056,N_14209);
nor U16210 (N_16210,N_13797,N_13823);
xnor U16211 (N_16211,N_14403,N_13985);
or U16212 (N_16212,N_14303,N_14347);
xnor U16213 (N_16213,N_14487,N_14027);
nand U16214 (N_16214,N_14814,N_14614);
or U16215 (N_16215,N_14749,N_13926);
nor U16216 (N_16216,N_14193,N_14548);
xor U16217 (N_16217,N_14785,N_14091);
nand U16218 (N_16218,N_14855,N_14703);
and U16219 (N_16219,N_14124,N_14669);
xor U16220 (N_16220,N_14272,N_14939);
and U16221 (N_16221,N_14800,N_14566);
nand U16222 (N_16222,N_14369,N_14091);
or U16223 (N_16223,N_14000,N_13786);
or U16224 (N_16224,N_14500,N_14436);
xnor U16225 (N_16225,N_14986,N_14857);
nor U16226 (N_16226,N_14672,N_14408);
xnor U16227 (N_16227,N_14420,N_13841);
xnor U16228 (N_16228,N_14645,N_14463);
xnor U16229 (N_16229,N_13787,N_14334);
and U16230 (N_16230,N_14314,N_14832);
xor U16231 (N_16231,N_14980,N_14720);
or U16232 (N_16232,N_14292,N_14461);
nor U16233 (N_16233,N_14336,N_14909);
xor U16234 (N_16234,N_14747,N_13804);
nor U16235 (N_16235,N_14137,N_13918);
or U16236 (N_16236,N_13864,N_14405);
nor U16237 (N_16237,N_14178,N_14232);
or U16238 (N_16238,N_14809,N_14450);
xor U16239 (N_16239,N_14240,N_14758);
nor U16240 (N_16240,N_14345,N_14001);
xor U16241 (N_16241,N_14686,N_14585);
nor U16242 (N_16242,N_14008,N_14345);
nand U16243 (N_16243,N_14637,N_14359);
nor U16244 (N_16244,N_14529,N_14422);
nor U16245 (N_16245,N_13795,N_14522);
or U16246 (N_16246,N_14620,N_14919);
nor U16247 (N_16247,N_14585,N_14133);
and U16248 (N_16248,N_13871,N_13779);
or U16249 (N_16249,N_14164,N_14140);
or U16250 (N_16250,N_15766,N_15357);
or U16251 (N_16251,N_15488,N_16160);
and U16252 (N_16252,N_15566,N_15169);
and U16253 (N_16253,N_16159,N_15468);
nand U16254 (N_16254,N_16097,N_16030);
xor U16255 (N_16255,N_15992,N_15844);
nand U16256 (N_16256,N_15818,N_15881);
and U16257 (N_16257,N_15816,N_15453);
nor U16258 (N_16258,N_15591,N_15230);
or U16259 (N_16259,N_15295,N_16164);
or U16260 (N_16260,N_16178,N_16080);
and U16261 (N_16261,N_15895,N_15864);
or U16262 (N_16262,N_15142,N_15603);
xor U16263 (N_16263,N_16041,N_15671);
and U16264 (N_16264,N_15751,N_15224);
nor U16265 (N_16265,N_15989,N_15189);
nor U16266 (N_16266,N_16013,N_16121);
or U16267 (N_16267,N_15791,N_15977);
or U16268 (N_16268,N_16083,N_15660);
nor U16269 (N_16269,N_15546,N_15690);
or U16270 (N_16270,N_15408,N_15059);
nand U16271 (N_16271,N_15374,N_15839);
nor U16272 (N_16272,N_15858,N_16082);
xor U16273 (N_16273,N_15054,N_15787);
nor U16274 (N_16274,N_15903,N_15642);
nor U16275 (N_16275,N_15337,N_15849);
and U16276 (N_16276,N_15792,N_15820);
and U16277 (N_16277,N_15372,N_15819);
and U16278 (N_16278,N_15076,N_15853);
nand U16279 (N_16279,N_16109,N_15950);
or U16280 (N_16280,N_15099,N_15214);
and U16281 (N_16281,N_15795,N_15510);
nand U16282 (N_16282,N_15416,N_15156);
nor U16283 (N_16283,N_15356,N_15748);
xor U16284 (N_16284,N_15843,N_15559);
xnor U16285 (N_16285,N_15410,N_16192);
nor U16286 (N_16286,N_15427,N_15702);
nor U16287 (N_16287,N_15002,N_15062);
nor U16288 (N_16288,N_16107,N_15639);
nand U16289 (N_16289,N_15432,N_16103);
and U16290 (N_16290,N_15784,N_15531);
nand U16291 (N_16291,N_15562,N_15484);
xnor U16292 (N_16292,N_15392,N_16173);
or U16293 (N_16293,N_15759,N_15580);
nand U16294 (N_16294,N_15153,N_16196);
and U16295 (N_16295,N_16072,N_15921);
xnor U16296 (N_16296,N_15065,N_15840);
or U16297 (N_16297,N_15343,N_16248);
nand U16298 (N_16298,N_16119,N_15871);
nor U16299 (N_16299,N_15389,N_15877);
xor U16300 (N_16300,N_15037,N_15708);
and U16301 (N_16301,N_15874,N_15404);
nand U16302 (N_16302,N_15483,N_15164);
and U16303 (N_16303,N_16106,N_15929);
nand U16304 (N_16304,N_15873,N_15543);
or U16305 (N_16305,N_15683,N_15016);
or U16306 (N_16306,N_15685,N_15129);
and U16307 (N_16307,N_15362,N_15331);
nand U16308 (N_16308,N_15833,N_15000);
nand U16309 (N_16309,N_15563,N_15560);
and U16310 (N_16310,N_15346,N_15493);
nor U16311 (N_16311,N_15110,N_15624);
nor U16312 (N_16312,N_15090,N_15472);
or U16313 (N_16313,N_15712,N_15737);
xor U16314 (N_16314,N_15569,N_15042);
and U16315 (N_16315,N_15181,N_15567);
nand U16316 (N_16316,N_16139,N_15985);
nor U16317 (N_16317,N_16091,N_15750);
nand U16318 (N_16318,N_15834,N_15268);
or U16319 (N_16319,N_15278,N_15023);
nand U16320 (N_16320,N_15261,N_16057);
and U16321 (N_16321,N_15707,N_15595);
nand U16322 (N_16322,N_15915,N_15947);
and U16323 (N_16323,N_15383,N_15956);
nand U16324 (N_16324,N_15705,N_15553);
or U16325 (N_16325,N_16108,N_15315);
xor U16326 (N_16326,N_15237,N_15443);
and U16327 (N_16327,N_16169,N_15323);
nor U16328 (N_16328,N_15353,N_15241);
or U16329 (N_16329,N_15201,N_15260);
and U16330 (N_16330,N_15263,N_15980);
nand U16331 (N_16331,N_15288,N_15084);
nor U16332 (N_16332,N_16226,N_16092);
nand U16333 (N_16333,N_15534,N_15186);
nor U16334 (N_16334,N_15758,N_16074);
nand U16335 (N_16335,N_15347,N_15266);
nor U16336 (N_16336,N_15361,N_15991);
xnor U16337 (N_16337,N_15137,N_15893);
and U16338 (N_16338,N_15317,N_16238);
and U16339 (N_16339,N_15338,N_15857);
nand U16340 (N_16340,N_16149,N_15293);
xnor U16341 (N_16341,N_15909,N_15025);
nor U16342 (N_16342,N_16128,N_15598);
xnor U16343 (N_16343,N_15637,N_15774);
and U16344 (N_16344,N_15222,N_15327);
xnor U16345 (N_16345,N_15652,N_16167);
nand U16346 (N_16346,N_15092,N_15300);
or U16347 (N_16347,N_15400,N_15437);
nor U16348 (N_16348,N_15967,N_15131);
nor U16349 (N_16349,N_15718,N_16059);
nor U16350 (N_16350,N_15280,N_15005);
xor U16351 (N_16351,N_15243,N_15157);
nor U16352 (N_16352,N_15020,N_15206);
nor U16353 (N_16353,N_15987,N_16098);
xor U16354 (N_16354,N_15140,N_15739);
xor U16355 (N_16355,N_15093,N_15942);
and U16356 (N_16356,N_15611,N_15878);
or U16357 (N_16357,N_15167,N_15255);
xnor U16358 (N_16358,N_15886,N_15756);
xnor U16359 (N_16359,N_15572,N_15355);
or U16360 (N_16360,N_15015,N_16202);
or U16361 (N_16361,N_16158,N_15066);
nor U16362 (N_16362,N_15182,N_15281);
or U16363 (N_16363,N_15662,N_15141);
xor U16364 (N_16364,N_15646,N_15163);
nand U16365 (N_16365,N_15876,N_15313);
or U16366 (N_16366,N_16211,N_16034);
nand U16367 (N_16367,N_15934,N_16145);
and U16368 (N_16368,N_15173,N_15018);
and U16369 (N_16369,N_16191,N_15533);
xor U16370 (N_16370,N_15183,N_15749);
xor U16371 (N_16371,N_15095,N_15729);
nand U16372 (N_16372,N_15867,N_15863);
or U16373 (N_16373,N_15862,N_15574);
xnor U16374 (N_16374,N_15064,N_15291);
nand U16375 (N_16375,N_15767,N_15826);
and U16376 (N_16376,N_16125,N_15407);
nand U16377 (N_16377,N_15974,N_16155);
or U16378 (N_16378,N_15587,N_15134);
xor U16379 (N_16379,N_15375,N_15350);
and U16380 (N_16380,N_15755,N_15412);
nand U16381 (N_16381,N_15068,N_15390);
nor U16382 (N_16382,N_15511,N_15161);
nor U16383 (N_16383,N_15986,N_16180);
nand U16384 (N_16384,N_16079,N_15231);
nand U16385 (N_16385,N_15512,N_15663);
xor U16386 (N_16386,N_15846,N_15556);
and U16387 (N_16387,N_15938,N_15664);
nand U16388 (N_16388,N_15673,N_15732);
nand U16389 (N_16389,N_15925,N_15936);
xnor U16390 (N_16390,N_15087,N_15686);
nor U16391 (N_16391,N_15238,N_15244);
nor U16392 (N_16392,N_15223,N_15406);
xnor U16393 (N_16393,N_15115,N_15401);
and U16394 (N_16394,N_15778,N_15848);
nor U16395 (N_16395,N_16064,N_15379);
or U16396 (N_16396,N_15460,N_15117);
xor U16397 (N_16397,N_15860,N_15462);
nand U16398 (N_16398,N_16242,N_15882);
xnor U16399 (N_16399,N_15588,N_15594);
xnor U16400 (N_16400,N_15202,N_15612);
xnor U16401 (N_16401,N_15668,N_15684);
nand U16402 (N_16402,N_15490,N_15417);
xor U16403 (N_16403,N_15665,N_15184);
xor U16404 (N_16404,N_15190,N_16019);
and U16405 (N_16405,N_15289,N_15828);
nand U16406 (N_16406,N_16100,N_16234);
nand U16407 (N_16407,N_15108,N_15122);
nor U16408 (N_16408,N_15249,N_15529);
or U16409 (N_16409,N_15616,N_15258);
and U16410 (N_16410,N_15645,N_15609);
or U16411 (N_16411,N_15365,N_15627);
xnor U16412 (N_16412,N_16210,N_16136);
or U16413 (N_16413,N_15957,N_15101);
xnor U16414 (N_16414,N_15763,N_15388);
nor U16415 (N_16415,N_15777,N_15040);
and U16416 (N_16416,N_16032,N_16183);
nor U16417 (N_16417,N_16005,N_15058);
and U16418 (N_16418,N_15709,N_16081);
and U16419 (N_16419,N_15172,N_15855);
nor U16420 (N_16420,N_15815,N_15807);
xnor U16421 (N_16421,N_15333,N_15923);
nand U16422 (N_16422,N_15803,N_15381);
nand U16423 (N_16423,N_15813,N_15414);
and U16424 (N_16424,N_16049,N_15455);
xor U16425 (N_16425,N_15901,N_15177);
nand U16426 (N_16426,N_15339,N_16201);
and U16427 (N_16427,N_15364,N_15378);
and U16428 (N_16428,N_15396,N_15586);
nand U16429 (N_16429,N_15485,N_15297);
or U16430 (N_16430,N_15780,N_15074);
nand U16431 (N_16431,N_15139,N_15854);
nand U16432 (N_16432,N_15608,N_15838);
nor U16433 (N_16433,N_15688,N_15622);
nor U16434 (N_16434,N_15109,N_15366);
xor U16435 (N_16435,N_16245,N_15711);
and U16436 (N_16436,N_16231,N_16190);
and U16437 (N_16437,N_15461,N_15118);
or U16438 (N_16438,N_15158,N_15841);
nand U16439 (N_16439,N_15382,N_15552);
nor U16440 (N_16440,N_15677,N_15007);
nor U16441 (N_16441,N_15091,N_15228);
or U16442 (N_16442,N_15527,N_15304);
xor U16443 (N_16443,N_15330,N_15779);
xnor U16444 (N_16444,N_16235,N_15053);
and U16445 (N_16445,N_16162,N_15935);
nand U16446 (N_16446,N_16143,N_15889);
and U16447 (N_16447,N_15028,N_15088);
xnor U16448 (N_16448,N_15457,N_15963);
nand U16449 (N_16449,N_15875,N_15227);
nand U16450 (N_16450,N_15080,N_16138);
or U16451 (N_16451,N_15786,N_15928);
nor U16452 (N_16452,N_16070,N_15997);
nand U16453 (N_16453,N_16084,N_15638);
or U16454 (N_16454,N_15789,N_15910);
nand U16455 (N_16455,N_15530,N_15212);
xor U16456 (N_16456,N_16176,N_16221);
nor U16457 (N_16457,N_15340,N_15648);
nor U16458 (N_16458,N_16227,N_15395);
xor U16459 (N_16459,N_15229,N_16040);
and U16460 (N_16460,N_15623,N_15976);
and U16461 (N_16461,N_15273,N_15049);
nor U16462 (N_16462,N_15719,N_15575);
xnor U16463 (N_16463,N_15504,N_15644);
and U16464 (N_16464,N_15336,N_16104);
and U16465 (N_16465,N_15880,N_15904);
and U16466 (N_16466,N_15341,N_15680);
xnor U16467 (N_16467,N_15983,N_15492);
and U16468 (N_16468,N_15681,N_15405);
nand U16469 (N_16469,N_15618,N_15576);
xor U16470 (N_16470,N_15692,N_16111);
nor U16471 (N_16471,N_15011,N_15620);
nor U16472 (N_16472,N_15104,N_15344);
or U16473 (N_16473,N_16193,N_15275);
nor U16474 (N_16474,N_15017,N_16152);
and U16475 (N_16475,N_16053,N_15165);
xor U16476 (N_16476,N_16045,N_16020);
xnor U16477 (N_16477,N_15498,N_16050);
or U16478 (N_16478,N_15348,N_16007);
or U16479 (N_16479,N_15103,N_16224);
xnor U16480 (N_16480,N_15445,N_15292);
nor U16481 (N_16481,N_15653,N_15486);
nor U16482 (N_16482,N_15305,N_15981);
nor U16483 (N_16483,N_15192,N_16011);
or U16484 (N_16484,N_15402,N_15319);
and U16485 (N_16485,N_15812,N_16117);
nand U16486 (N_16486,N_15440,N_15502);
and U16487 (N_16487,N_15359,N_15666);
nand U16488 (N_16488,N_15600,N_15953);
or U16489 (N_16489,N_16179,N_15822);
xor U16490 (N_16490,N_15334,N_16120);
or U16491 (N_16491,N_15418,N_15265);
xor U16492 (N_16492,N_15994,N_15727);
xnor U16493 (N_16493,N_15513,N_16156);
or U16494 (N_16494,N_15937,N_15496);
nand U16495 (N_16495,N_15900,N_15403);
and U16496 (N_16496,N_15741,N_15473);
nor U16497 (N_16497,N_16177,N_15162);
xnor U16498 (N_16498,N_15969,N_15450);
xnor U16499 (N_16499,N_15063,N_15428);
nor U16500 (N_16500,N_15318,N_15593);
nand U16501 (N_16501,N_16229,N_15931);
nand U16502 (N_16502,N_15776,N_15503);
and U16503 (N_16503,N_16067,N_15806);
or U16504 (N_16504,N_15917,N_15036);
nor U16505 (N_16505,N_15125,N_15501);
nand U16506 (N_16506,N_15415,N_15276);
xnor U16507 (N_16507,N_15831,N_15655);
or U16508 (N_16508,N_15973,N_15602);
nor U16509 (N_16509,N_15479,N_15596);
or U16510 (N_16510,N_15772,N_15670);
and U16511 (N_16511,N_16187,N_15470);
nor U16512 (N_16512,N_15207,N_15194);
nor U16513 (N_16513,N_15233,N_15522);
or U16514 (N_16514,N_15674,N_15810);
or U16515 (N_16515,N_15733,N_15247);
nor U16516 (N_16516,N_15892,N_15649);
or U16517 (N_16517,N_15217,N_15286);
xor U16518 (N_16518,N_15085,N_15218);
or U16519 (N_16519,N_15285,N_16068);
xnor U16520 (N_16520,N_15151,N_15883);
and U16521 (N_16521,N_15466,N_15940);
and U16522 (N_16522,N_15647,N_15597);
nand U16523 (N_16523,N_15782,N_15640);
nor U16524 (N_16524,N_16220,N_15146);
nand U16525 (N_16525,N_16085,N_15689);
nand U16526 (N_16526,N_15982,N_15545);
or U16527 (N_16527,N_15185,N_16036);
and U16528 (N_16528,N_15113,N_15475);
nand U16529 (N_16529,N_16142,N_15918);
nand U16530 (N_16530,N_15430,N_15061);
nand U16531 (N_16531,N_16124,N_15298);
xnor U16532 (N_16532,N_16056,N_15254);
and U16533 (N_16533,N_15879,N_16209);
nand U16534 (N_16534,N_16203,N_15262);
xor U16535 (N_16535,N_15480,N_16060);
or U16536 (N_16536,N_15138,N_15724);
nor U16537 (N_16537,N_15342,N_15271);
or U16538 (N_16538,N_16008,N_15436);
or U16539 (N_16539,N_15006,N_15377);
and U16540 (N_16540,N_15558,N_16218);
xnor U16541 (N_16541,N_15523,N_15145);
xor U16542 (N_16542,N_15519,N_15927);
or U16543 (N_16543,N_15120,N_15500);
and U16544 (N_16544,N_15474,N_15220);
and U16545 (N_16545,N_15625,N_15868);
or U16546 (N_16546,N_15538,N_15924);
nor U16547 (N_16547,N_16055,N_16004);
and U16548 (N_16548,N_15012,N_16246);
nand U16549 (N_16549,N_15824,N_15544);
xor U16550 (N_16550,N_15451,N_15526);
nand U16551 (N_16551,N_15078,N_15897);
xnor U16552 (N_16552,N_15699,N_16010);
nor U16553 (N_16553,N_15199,N_15585);
nand U16554 (N_16554,N_15630,N_15615);
xor U16555 (N_16555,N_16094,N_15111);
nor U16556 (N_16556,N_15055,N_16236);
and U16557 (N_16557,N_15010,N_15213);
nand U16558 (N_16558,N_15399,N_16182);
xor U16559 (N_16559,N_15105,N_15852);
nor U16560 (N_16560,N_15469,N_15635);
and U16561 (N_16561,N_15208,N_15550);
nand U16562 (N_16562,N_15850,N_15051);
and U16563 (N_16563,N_15659,N_16163);
or U16564 (N_16564,N_15713,N_15761);
or U16565 (N_16565,N_16243,N_15565);
or U16566 (N_16566,N_15887,N_15604);
xnor U16567 (N_16567,N_16022,N_15069);
nand U16568 (N_16568,N_16043,N_15861);
nor U16569 (N_16569,N_16207,N_15539);
and U16570 (N_16570,N_15832,N_15335);
nand U16571 (N_16571,N_16017,N_15962);
nor U16572 (N_16572,N_15497,N_16071);
xor U16573 (N_16573,N_16112,N_16223);
nor U16574 (N_16574,N_15411,N_16029);
and U16575 (N_16575,N_15248,N_15482);
xor U16576 (N_16576,N_15606,N_16174);
nand U16577 (N_16577,N_15817,N_15004);
nor U16578 (N_16578,N_15132,N_15001);
xnor U16579 (N_16579,N_16077,N_15380);
nand U16580 (N_16580,N_15715,N_16087);
xnor U16581 (N_16581,N_16054,N_15203);
or U16582 (N_16582,N_15768,N_15035);
or U16583 (N_16583,N_16214,N_15592);
nor U16584 (N_16584,N_15371,N_15256);
nor U16585 (N_16585,N_15252,N_15210);
and U16586 (N_16586,N_15632,N_15573);
or U16587 (N_16587,N_15701,N_16239);
nor U16588 (N_16588,N_16023,N_15204);
nand U16589 (N_16589,N_16151,N_16063);
nand U16590 (N_16590,N_15176,N_15532);
or U16591 (N_16591,N_15413,N_15021);
nand U16592 (N_16592,N_15106,N_15481);
and U16593 (N_16593,N_15825,N_15170);
or U16594 (N_16594,N_15514,N_15471);
xor U16595 (N_16595,N_16096,N_15913);
xnor U16596 (N_16596,N_15730,N_16137);
or U16597 (N_16597,N_16047,N_15933);
nor U16598 (N_16598,N_15746,N_15654);
and U16599 (N_16599,N_15870,N_15083);
xor U16600 (N_16600,N_16146,N_15975);
xor U16601 (N_16601,N_16184,N_15706);
or U16602 (N_16602,N_15384,N_15769);
nand U16603 (N_16603,N_15765,N_15740);
or U16604 (N_16604,N_16009,N_15147);
nor U16605 (N_16605,N_15951,N_15507);
xor U16606 (N_16606,N_16212,N_16101);
xnor U16607 (N_16607,N_15958,N_16076);
nor U16608 (N_16608,N_15166,N_15738);
nand U16609 (N_16609,N_15253,N_15926);
nor U16610 (N_16610,N_16026,N_15008);
nor U16611 (N_16611,N_15859,N_15964);
and U16612 (N_16612,N_16147,N_15128);
or U16613 (N_16613,N_16127,N_15272);
and U16614 (N_16614,N_15454,N_15676);
nand U16615 (N_16615,N_15143,N_15745);
and U16616 (N_16616,N_15024,N_15310);
or U16617 (N_16617,N_15056,N_15150);
or U16618 (N_16618,N_16217,N_15041);
or U16619 (N_16619,N_16206,N_15352);
or U16620 (N_16620,N_15643,N_15578);
and U16621 (N_16621,N_15014,N_15726);
or U16622 (N_16622,N_15089,N_16105);
nor U16623 (N_16623,N_15823,N_15376);
and U16624 (N_16624,N_16044,N_15720);
and U16625 (N_16625,N_16200,N_15112);
xnor U16626 (N_16626,N_15785,N_15155);
nor U16627 (N_16627,N_15836,N_15495);
xor U16628 (N_16628,N_15039,N_15013);
xor U16629 (N_16629,N_15235,N_15325);
xnor U16630 (N_16630,N_15747,N_15731);
nand U16631 (N_16631,N_16126,N_15219);
or U16632 (N_16632,N_16150,N_15703);
or U16633 (N_16633,N_16129,N_15775);
nor U16634 (N_16634,N_16058,N_15048);
and U16635 (N_16635,N_15193,N_15809);
xor U16636 (N_16636,N_15232,N_15521);
or U16637 (N_16637,N_15905,N_15439);
xnor U16638 (N_16638,N_16195,N_15075);
and U16639 (N_16639,N_15762,N_16073);
xor U16640 (N_16640,N_15046,N_15296);
or U16641 (N_16641,N_15050,N_15830);
xnor U16642 (N_16642,N_15988,N_15571);
nor U16643 (N_16643,N_15517,N_15043);
nor U16644 (N_16644,N_15299,N_15851);
nor U16645 (N_16645,N_15052,N_15796);
or U16646 (N_16646,N_15661,N_15302);
and U16647 (N_16647,N_15409,N_15136);
xor U16648 (N_16648,N_15242,N_15245);
nor U16649 (N_16649,N_16170,N_15047);
and U16650 (N_16650,N_15160,N_15094);
nor U16651 (N_16651,N_15426,N_15790);
xnor U16652 (N_16652,N_15393,N_15736);
nor U16653 (N_16653,N_15998,N_15941);
xnor U16654 (N_16654,N_15865,N_15696);
or U16655 (N_16655,N_15697,N_15633);
nor U16656 (N_16656,N_15067,N_15996);
or U16657 (N_16657,N_16115,N_16133);
or U16658 (N_16658,N_16153,N_15525);
or U16659 (N_16659,N_15277,N_16095);
xnor U16660 (N_16660,N_15954,N_15629);
and U16661 (N_16661,N_15345,N_15060);
or U16662 (N_16662,N_15943,N_15351);
or U16663 (N_16663,N_15397,N_15970);
nand U16664 (N_16664,N_15524,N_15551);
xnor U16665 (N_16665,N_15695,N_15902);
or U16666 (N_16666,N_16233,N_15124);
nor U16667 (N_16667,N_16186,N_16228);
nor U16668 (N_16668,N_15171,N_15282);
nand U16669 (N_16669,N_15694,N_15442);
and U16670 (N_16670,N_15456,N_15209);
xor U16671 (N_16671,N_16213,N_15234);
nand U16672 (N_16672,N_15385,N_16021);
or U16673 (N_16673,N_16114,N_15528);
nand U16674 (N_16674,N_15329,N_15205);
and U16675 (N_16675,N_15847,N_15211);
and U16676 (N_16676,N_15743,N_15081);
nand U16677 (N_16677,N_16006,N_16189);
or U16678 (N_16678,N_16215,N_16172);
nor U16679 (N_16679,N_15914,N_15434);
nor U16680 (N_16680,N_16130,N_16157);
or U16681 (N_16681,N_15126,N_15425);
and U16682 (N_16682,N_16046,N_15387);
nor U16683 (N_16683,N_15518,N_15908);
xor U16684 (N_16684,N_16185,N_15581);
nor U16685 (N_16685,N_15890,N_15650);
nand U16686 (N_16686,N_15033,N_16140);
and U16687 (N_16687,N_15599,N_16000);
nand U16688 (N_16688,N_15423,N_15239);
xor U16689 (N_16689,N_15722,N_15130);
and U16690 (N_16690,N_15554,N_15894);
and U16691 (N_16691,N_15959,N_15752);
and U16692 (N_16692,N_16089,N_15948);
and U16693 (N_16693,N_15320,N_15398);
or U16694 (N_16694,N_15770,N_16219);
or U16695 (N_16695,N_15449,N_15601);
or U16696 (N_16696,N_15386,N_15179);
nor U16697 (N_16697,N_16237,N_15829);
and U16698 (N_16698,N_15907,N_15360);
xor U16699 (N_16699,N_16099,N_15491);
or U16700 (N_16700,N_16171,N_15788);
xnor U16701 (N_16701,N_15658,N_15760);
nor U16702 (N_16702,N_15174,N_15773);
and U16703 (N_16703,N_15031,N_16018);
or U16704 (N_16704,N_16027,N_16241);
nor U16705 (N_16705,N_15509,N_16052);
and U16706 (N_16706,N_15734,N_15999);
nand U16707 (N_16707,N_16116,N_16118);
or U16708 (N_16708,N_15783,N_15236);
or U16709 (N_16709,N_15148,N_16135);
nor U16710 (N_16710,N_15930,N_15717);
xor U16711 (N_16711,N_15872,N_15949);
or U16712 (N_16712,N_16197,N_15541);
nand U16713 (N_16713,N_15102,N_15979);
nand U16714 (N_16714,N_16154,N_16166);
xor U16715 (N_16715,N_15358,N_15187);
and U16716 (N_16716,N_15429,N_15274);
and U16717 (N_16717,N_15570,N_15431);
xor U16718 (N_16718,N_16065,N_15944);
xnor U16719 (N_16719,N_15693,N_15435);
and U16720 (N_16720,N_15764,N_16038);
xnor U16721 (N_16721,N_16198,N_15314);
or U16722 (N_16722,N_15306,N_15096);
nor U16723 (N_16723,N_15899,N_15520);
xnor U16724 (N_16724,N_15499,N_15422);
xnor U16725 (N_16725,N_16122,N_15798);
nor U16726 (N_16726,N_16039,N_15463);
nand U16727 (N_16727,N_15607,N_15621);
xnor U16728 (N_16728,N_15257,N_15771);
xor U16729 (N_16729,N_16225,N_16086);
nand U16730 (N_16730,N_15716,N_15188);
nand U16731 (N_16731,N_15960,N_15373);
nand U16732 (N_16732,N_15515,N_15728);
nor U16733 (N_16733,N_15154,N_16208);
xor U16734 (N_16734,N_15003,N_16240);
nor U16735 (N_16735,N_15896,N_15919);
nor U16736 (N_16736,N_15993,N_16247);
xnor U16737 (N_16737,N_15478,N_15367);
and U16738 (N_16738,N_15626,N_15477);
nor U16739 (N_16739,N_15856,N_15200);
xor U16740 (N_16740,N_15577,N_15446);
xnor U16741 (N_16741,N_15196,N_15097);
and U16742 (N_16742,N_16199,N_16204);
nand U16743 (N_16743,N_15885,N_15547);
nand U16744 (N_16744,N_15579,N_16148);
nor U16745 (N_16745,N_15634,N_15489);
nor U16746 (N_16746,N_15197,N_16012);
or U16747 (N_16747,N_15326,N_15116);
nor U16748 (N_16748,N_15121,N_15191);
nand U16749 (N_16749,N_15029,N_15700);
nand U16750 (N_16750,N_16222,N_15516);
nand U16751 (N_16751,N_15019,N_15582);
and U16752 (N_16752,N_15267,N_16134);
nand U16753 (N_16753,N_16069,N_16035);
xnor U16754 (N_16754,N_15100,N_16088);
nor U16755 (N_16755,N_16033,N_15656);
xor U16756 (N_16756,N_15250,N_15424);
nor U16757 (N_16757,N_16031,N_15419);
or U16758 (N_16758,N_15114,N_15869);
or U16759 (N_16759,N_15610,N_16181);
nand U16760 (N_16760,N_16062,N_16144);
xnor U16761 (N_16761,N_15557,N_15968);
nand U16762 (N_16762,N_15368,N_15613);
and U16763 (N_16763,N_15672,N_15631);
and U16764 (N_16764,N_16075,N_15687);
or U16765 (N_16765,N_15691,N_15704);
and U16766 (N_16766,N_15866,N_15322);
nand U16767 (N_16767,N_16113,N_15133);
and U16768 (N_16768,N_15195,N_15321);
nand U16769 (N_16769,N_16216,N_16002);
nand U16770 (N_16770,N_15744,N_16037);
nand U16771 (N_16771,N_15564,N_15438);
and U16772 (N_16772,N_15804,N_16205);
and U16773 (N_16773,N_15583,N_15045);
or U16774 (N_16774,N_15269,N_15781);
xor U16775 (N_16775,N_15605,N_16093);
nor U16776 (N_16776,N_15026,N_15754);
nand U16777 (N_16777,N_15178,N_15906);
nor U16778 (N_16778,N_16131,N_15303);
and U16779 (N_16779,N_15536,N_15952);
or U16780 (N_16780,N_15226,N_15971);
xnor U16781 (N_16781,N_15535,N_16194);
nor U16782 (N_16782,N_15284,N_15753);
nand U16783 (N_16783,N_15082,N_15038);
nand U16784 (N_16784,N_15316,N_15444);
nor U16785 (N_16785,N_15290,N_15240);
nor U16786 (N_16786,N_15127,N_15441);
nor U16787 (N_16787,N_16051,N_15742);
nand U16788 (N_16788,N_15287,N_15542);
nor U16789 (N_16789,N_15467,N_15448);
xnor U16790 (N_16790,N_16015,N_16003);
xor U16791 (N_16791,N_15590,N_15458);
and U16792 (N_16792,N_15487,N_15678);
and U16793 (N_16793,N_15794,N_16110);
xnor U16794 (N_16794,N_15301,N_15667);
xnor U16795 (N_16795,N_15168,N_15433);
and U16796 (N_16796,N_15932,N_15135);
xnor U16797 (N_16797,N_15452,N_15294);
nor U16798 (N_16798,N_15152,N_16141);
xnor U16799 (N_16799,N_15086,N_15675);
nor U16800 (N_16800,N_15175,N_16249);
nor U16801 (N_16801,N_15476,N_15030);
xor U16802 (N_16802,N_15619,N_15636);
nand U16803 (N_16803,N_16078,N_15363);
xor U16804 (N_16804,N_15978,N_16165);
or U16805 (N_16805,N_15800,N_15328);
or U16806 (N_16806,N_15072,N_15369);
nand U16807 (N_16807,N_16232,N_16014);
or U16808 (N_16808,N_15714,N_15568);
nor U16809 (N_16809,N_15679,N_15898);
nor U16810 (N_16810,N_15641,N_15027);
and U16811 (N_16811,N_15922,N_15447);
or U16812 (N_16812,N_15332,N_16123);
or U16813 (N_16813,N_16102,N_15561);
xor U16814 (N_16814,N_15682,N_15808);
nand U16815 (N_16815,N_15888,N_15032);
xor U16816 (N_16816,N_15802,N_15721);
xnor U16817 (N_16817,N_15628,N_16028);
and U16818 (N_16818,N_15349,N_15073);
xor U16819 (N_16819,N_15119,N_15669);
nor U16820 (N_16820,N_16161,N_15814);
and U16821 (N_16821,N_15549,N_15354);
xnor U16822 (N_16822,N_16025,N_15805);
nand U16823 (N_16823,N_15494,N_15797);
or U16824 (N_16824,N_15057,N_15657);
or U16825 (N_16825,N_15801,N_15098);
or U16826 (N_16826,N_15984,N_16244);
nand U16827 (N_16827,N_15077,N_15842);
and U16828 (N_16828,N_15149,N_15916);
and U16829 (N_16829,N_15939,N_15246);
nor U16830 (N_16830,N_15555,N_15022);
nand U16831 (N_16831,N_15465,N_16042);
and U16832 (N_16832,N_15966,N_15537);
xnor U16833 (N_16833,N_15180,N_15107);
nand U16834 (N_16834,N_15835,N_15216);
xor U16835 (N_16835,N_15505,N_15589);
nand U16836 (N_16836,N_16024,N_15912);
or U16837 (N_16837,N_15225,N_15370);
nand U16838 (N_16838,N_15123,N_15459);
nor U16839 (N_16839,N_15614,N_16230);
nand U16840 (N_16840,N_15221,N_15995);
or U16841 (N_16841,N_16175,N_15420);
nor U16842 (N_16842,N_15710,N_15799);
xor U16843 (N_16843,N_15540,N_15961);
nand U16844 (N_16844,N_15651,N_16090);
nor U16845 (N_16845,N_15159,N_15215);
xor U16846 (N_16846,N_15827,N_15884);
nor U16847 (N_16847,N_15845,N_15394);
or U16848 (N_16848,N_15309,N_15421);
or U16849 (N_16849,N_15821,N_16001);
xor U16850 (N_16850,N_15548,N_15617);
and U16851 (N_16851,N_15312,N_15071);
xnor U16852 (N_16852,N_15391,N_15009);
nor U16853 (N_16853,N_15034,N_15837);
and U16854 (N_16854,N_16066,N_16132);
nand U16855 (N_16855,N_15308,N_15920);
and U16856 (N_16856,N_15891,N_15044);
and U16857 (N_16857,N_15793,N_15270);
and U16858 (N_16858,N_16061,N_15946);
and U16859 (N_16859,N_15070,N_15324);
nand U16860 (N_16860,N_15283,N_15264);
nor U16861 (N_16861,N_15251,N_15945);
nand U16862 (N_16862,N_15198,N_15965);
and U16863 (N_16863,N_15990,N_15279);
xnor U16864 (N_16864,N_15911,N_15698);
and U16865 (N_16865,N_16188,N_15144);
or U16866 (N_16866,N_15311,N_15506);
xnor U16867 (N_16867,N_15259,N_16016);
nor U16868 (N_16868,N_16168,N_15464);
and U16869 (N_16869,N_15079,N_15955);
and U16870 (N_16870,N_15307,N_15811);
and U16871 (N_16871,N_15508,N_15972);
nand U16872 (N_16872,N_16048,N_15723);
or U16873 (N_16873,N_15584,N_15725);
or U16874 (N_16874,N_15735,N_15757);
nand U16875 (N_16875,N_15821,N_16236);
nor U16876 (N_16876,N_15145,N_15309);
or U16877 (N_16877,N_15045,N_15506);
xor U16878 (N_16878,N_15486,N_15731);
and U16879 (N_16879,N_15869,N_15536);
xnor U16880 (N_16880,N_15817,N_15993);
nand U16881 (N_16881,N_15005,N_15525);
and U16882 (N_16882,N_15364,N_15536);
or U16883 (N_16883,N_16126,N_16012);
or U16884 (N_16884,N_15879,N_15333);
nor U16885 (N_16885,N_15050,N_16100);
and U16886 (N_16886,N_15453,N_15327);
or U16887 (N_16887,N_16165,N_15429);
nor U16888 (N_16888,N_15638,N_15680);
nor U16889 (N_16889,N_15331,N_15808);
or U16890 (N_16890,N_15885,N_15681);
xnor U16891 (N_16891,N_15587,N_15044);
nor U16892 (N_16892,N_15808,N_15707);
or U16893 (N_16893,N_15113,N_15980);
nor U16894 (N_16894,N_16210,N_15647);
and U16895 (N_16895,N_15866,N_15879);
xor U16896 (N_16896,N_16173,N_15399);
nor U16897 (N_16897,N_15876,N_16036);
nor U16898 (N_16898,N_15840,N_15332);
nand U16899 (N_16899,N_15154,N_16136);
nand U16900 (N_16900,N_16071,N_15578);
or U16901 (N_16901,N_16161,N_15523);
and U16902 (N_16902,N_16081,N_15272);
and U16903 (N_16903,N_15075,N_15875);
or U16904 (N_16904,N_15362,N_15189);
nor U16905 (N_16905,N_15003,N_16029);
nor U16906 (N_16906,N_16014,N_15591);
and U16907 (N_16907,N_16100,N_15003);
nand U16908 (N_16908,N_15061,N_16116);
nor U16909 (N_16909,N_15942,N_15973);
or U16910 (N_16910,N_15764,N_15519);
and U16911 (N_16911,N_15372,N_15390);
xor U16912 (N_16912,N_15948,N_15773);
nand U16913 (N_16913,N_15618,N_15455);
xor U16914 (N_16914,N_15471,N_15391);
nand U16915 (N_16915,N_16084,N_16190);
and U16916 (N_16916,N_15464,N_16136);
or U16917 (N_16917,N_16093,N_15512);
or U16918 (N_16918,N_15252,N_15015);
xnor U16919 (N_16919,N_15677,N_15700);
and U16920 (N_16920,N_15990,N_15790);
and U16921 (N_16921,N_16015,N_16056);
nand U16922 (N_16922,N_15784,N_15936);
nand U16923 (N_16923,N_15907,N_16140);
nand U16924 (N_16924,N_15843,N_15441);
nand U16925 (N_16925,N_16153,N_15543);
or U16926 (N_16926,N_15444,N_15544);
xor U16927 (N_16927,N_16045,N_15959);
xor U16928 (N_16928,N_15035,N_15992);
xnor U16929 (N_16929,N_15730,N_15841);
xnor U16930 (N_16930,N_16026,N_15089);
xor U16931 (N_16931,N_15223,N_15697);
or U16932 (N_16932,N_15614,N_15705);
xor U16933 (N_16933,N_15120,N_15854);
and U16934 (N_16934,N_15265,N_16062);
or U16935 (N_16935,N_15044,N_15516);
nand U16936 (N_16936,N_16083,N_15730);
nor U16937 (N_16937,N_16157,N_15956);
and U16938 (N_16938,N_15925,N_16144);
or U16939 (N_16939,N_15233,N_15436);
nor U16940 (N_16940,N_15870,N_16092);
or U16941 (N_16941,N_15875,N_15128);
nor U16942 (N_16942,N_15268,N_15945);
xor U16943 (N_16943,N_15987,N_15346);
nor U16944 (N_16944,N_16027,N_15515);
nand U16945 (N_16945,N_16191,N_15827);
nor U16946 (N_16946,N_15327,N_15928);
or U16947 (N_16947,N_15831,N_16134);
xnor U16948 (N_16948,N_15255,N_15770);
and U16949 (N_16949,N_15410,N_15004);
or U16950 (N_16950,N_15297,N_15108);
nand U16951 (N_16951,N_15216,N_16024);
and U16952 (N_16952,N_15052,N_15054);
nand U16953 (N_16953,N_16249,N_15122);
and U16954 (N_16954,N_15321,N_15989);
or U16955 (N_16955,N_15658,N_15009);
or U16956 (N_16956,N_15178,N_15799);
nor U16957 (N_16957,N_15027,N_16227);
nor U16958 (N_16958,N_15415,N_15965);
or U16959 (N_16959,N_16178,N_16223);
xnor U16960 (N_16960,N_15028,N_15533);
nand U16961 (N_16961,N_15763,N_16020);
nor U16962 (N_16962,N_15142,N_15454);
and U16963 (N_16963,N_15759,N_15549);
xor U16964 (N_16964,N_16239,N_15162);
nor U16965 (N_16965,N_15987,N_15942);
nor U16966 (N_16966,N_15368,N_15230);
nor U16967 (N_16967,N_15242,N_15445);
nand U16968 (N_16968,N_16112,N_16198);
nor U16969 (N_16969,N_15212,N_15345);
or U16970 (N_16970,N_15721,N_16242);
xor U16971 (N_16971,N_15729,N_15509);
nor U16972 (N_16972,N_15798,N_15334);
and U16973 (N_16973,N_15783,N_16172);
nand U16974 (N_16974,N_16170,N_15757);
nand U16975 (N_16975,N_15084,N_15362);
nand U16976 (N_16976,N_15847,N_15136);
nand U16977 (N_16977,N_15106,N_15589);
xor U16978 (N_16978,N_15180,N_16003);
nand U16979 (N_16979,N_15176,N_15581);
and U16980 (N_16980,N_15842,N_15585);
xor U16981 (N_16981,N_15383,N_16094);
or U16982 (N_16982,N_15236,N_15109);
or U16983 (N_16983,N_16111,N_15799);
nand U16984 (N_16984,N_15126,N_15818);
and U16985 (N_16985,N_16215,N_15646);
nor U16986 (N_16986,N_15236,N_15426);
and U16987 (N_16987,N_16193,N_16209);
nand U16988 (N_16988,N_15346,N_16056);
nand U16989 (N_16989,N_15708,N_15485);
and U16990 (N_16990,N_15092,N_15623);
and U16991 (N_16991,N_16165,N_16228);
nand U16992 (N_16992,N_15832,N_15650);
xnor U16993 (N_16993,N_16138,N_15042);
and U16994 (N_16994,N_15842,N_15736);
nor U16995 (N_16995,N_15973,N_16010);
or U16996 (N_16996,N_16156,N_15500);
nand U16997 (N_16997,N_15634,N_15220);
nor U16998 (N_16998,N_15050,N_15133);
nand U16999 (N_16999,N_15207,N_16095);
nor U17000 (N_17000,N_15261,N_16247);
nand U17001 (N_17001,N_15644,N_16049);
nand U17002 (N_17002,N_15649,N_15983);
or U17003 (N_17003,N_15159,N_15330);
or U17004 (N_17004,N_16023,N_15193);
nor U17005 (N_17005,N_15582,N_15075);
nand U17006 (N_17006,N_15244,N_16060);
nand U17007 (N_17007,N_15866,N_15777);
xor U17008 (N_17008,N_15545,N_15270);
nor U17009 (N_17009,N_16108,N_15540);
xnor U17010 (N_17010,N_15326,N_15631);
nor U17011 (N_17011,N_15831,N_15880);
nand U17012 (N_17012,N_15482,N_15179);
or U17013 (N_17013,N_15375,N_15294);
nand U17014 (N_17014,N_15364,N_16238);
nor U17015 (N_17015,N_16134,N_15213);
or U17016 (N_17016,N_15414,N_15638);
nand U17017 (N_17017,N_15037,N_15250);
or U17018 (N_17018,N_16246,N_15242);
xor U17019 (N_17019,N_15187,N_15840);
or U17020 (N_17020,N_15266,N_15793);
and U17021 (N_17021,N_16034,N_15736);
xor U17022 (N_17022,N_15008,N_16117);
xnor U17023 (N_17023,N_15493,N_15726);
xor U17024 (N_17024,N_15495,N_15358);
and U17025 (N_17025,N_15686,N_15355);
and U17026 (N_17026,N_15868,N_15242);
or U17027 (N_17027,N_15143,N_15181);
nand U17028 (N_17028,N_15460,N_15602);
xor U17029 (N_17029,N_15395,N_15847);
nor U17030 (N_17030,N_15794,N_15053);
nor U17031 (N_17031,N_15525,N_16238);
or U17032 (N_17032,N_15197,N_15112);
nor U17033 (N_17033,N_15940,N_15063);
xor U17034 (N_17034,N_15613,N_15478);
and U17035 (N_17035,N_15195,N_15783);
nand U17036 (N_17036,N_15526,N_15357);
nand U17037 (N_17037,N_15456,N_16202);
nand U17038 (N_17038,N_15800,N_16064);
and U17039 (N_17039,N_15791,N_15865);
or U17040 (N_17040,N_15130,N_15535);
nand U17041 (N_17041,N_15065,N_15911);
or U17042 (N_17042,N_15302,N_15688);
nor U17043 (N_17043,N_15815,N_15916);
and U17044 (N_17044,N_15938,N_15370);
nor U17045 (N_17045,N_15099,N_15930);
nand U17046 (N_17046,N_15989,N_16126);
or U17047 (N_17047,N_15624,N_15690);
or U17048 (N_17048,N_15602,N_16184);
xnor U17049 (N_17049,N_16036,N_16007);
nand U17050 (N_17050,N_15525,N_16149);
nor U17051 (N_17051,N_15556,N_15409);
nor U17052 (N_17052,N_15764,N_15040);
xnor U17053 (N_17053,N_15302,N_15648);
nor U17054 (N_17054,N_15694,N_15517);
nor U17055 (N_17055,N_15952,N_15217);
and U17056 (N_17056,N_16208,N_15280);
nand U17057 (N_17057,N_15120,N_15455);
xor U17058 (N_17058,N_15390,N_15221);
or U17059 (N_17059,N_16028,N_15457);
nand U17060 (N_17060,N_16065,N_15318);
xnor U17061 (N_17061,N_15231,N_15086);
and U17062 (N_17062,N_15859,N_15933);
and U17063 (N_17063,N_15458,N_16065);
and U17064 (N_17064,N_16167,N_15309);
or U17065 (N_17065,N_15196,N_16101);
xor U17066 (N_17066,N_15225,N_16160);
xnor U17067 (N_17067,N_16132,N_16098);
and U17068 (N_17068,N_15137,N_16192);
or U17069 (N_17069,N_15215,N_15417);
xor U17070 (N_17070,N_15883,N_15073);
and U17071 (N_17071,N_16228,N_15048);
xor U17072 (N_17072,N_15924,N_15383);
nand U17073 (N_17073,N_16025,N_15388);
nand U17074 (N_17074,N_16053,N_15849);
nor U17075 (N_17075,N_15129,N_15710);
nand U17076 (N_17076,N_15723,N_15963);
and U17077 (N_17077,N_15025,N_15322);
xor U17078 (N_17078,N_15058,N_16202);
nand U17079 (N_17079,N_15989,N_16167);
nand U17080 (N_17080,N_15086,N_16014);
or U17081 (N_17081,N_15151,N_15285);
nor U17082 (N_17082,N_16050,N_16107);
nand U17083 (N_17083,N_16115,N_16063);
or U17084 (N_17084,N_15420,N_15371);
or U17085 (N_17085,N_15208,N_15529);
and U17086 (N_17086,N_16212,N_15504);
or U17087 (N_17087,N_15065,N_16144);
xnor U17088 (N_17088,N_15262,N_16149);
or U17089 (N_17089,N_15619,N_15459);
or U17090 (N_17090,N_15005,N_15942);
or U17091 (N_17091,N_15889,N_15193);
nand U17092 (N_17092,N_15611,N_15608);
and U17093 (N_17093,N_15620,N_16084);
or U17094 (N_17094,N_15391,N_15670);
nand U17095 (N_17095,N_15941,N_15788);
xor U17096 (N_17096,N_16165,N_15942);
and U17097 (N_17097,N_15137,N_15894);
nor U17098 (N_17098,N_15786,N_15284);
nor U17099 (N_17099,N_15038,N_15477);
xnor U17100 (N_17100,N_16227,N_15171);
nand U17101 (N_17101,N_15868,N_16240);
nor U17102 (N_17102,N_16031,N_15439);
xor U17103 (N_17103,N_15277,N_16120);
nor U17104 (N_17104,N_15127,N_15685);
and U17105 (N_17105,N_15261,N_15417);
and U17106 (N_17106,N_15451,N_16028);
and U17107 (N_17107,N_15379,N_15015);
nand U17108 (N_17108,N_15780,N_15271);
nor U17109 (N_17109,N_15735,N_15097);
nand U17110 (N_17110,N_15883,N_15947);
nand U17111 (N_17111,N_15028,N_15658);
or U17112 (N_17112,N_16207,N_16166);
and U17113 (N_17113,N_15776,N_15320);
xnor U17114 (N_17114,N_15624,N_15440);
nand U17115 (N_17115,N_15003,N_15676);
and U17116 (N_17116,N_15075,N_15756);
xnor U17117 (N_17117,N_15913,N_15449);
nand U17118 (N_17118,N_15143,N_15321);
and U17119 (N_17119,N_15813,N_15097);
and U17120 (N_17120,N_16232,N_15163);
and U17121 (N_17121,N_16162,N_15993);
nor U17122 (N_17122,N_15766,N_15564);
xor U17123 (N_17123,N_15571,N_15223);
xnor U17124 (N_17124,N_15047,N_16186);
and U17125 (N_17125,N_15361,N_15123);
or U17126 (N_17126,N_16079,N_15513);
nand U17127 (N_17127,N_15141,N_16030);
and U17128 (N_17128,N_16146,N_15777);
nand U17129 (N_17129,N_15288,N_15446);
nor U17130 (N_17130,N_15218,N_15215);
nor U17131 (N_17131,N_15328,N_15819);
or U17132 (N_17132,N_15649,N_15606);
xor U17133 (N_17133,N_15691,N_16112);
nor U17134 (N_17134,N_15320,N_15146);
nor U17135 (N_17135,N_15108,N_15645);
and U17136 (N_17136,N_15405,N_15309);
or U17137 (N_17137,N_16056,N_15193);
or U17138 (N_17138,N_15830,N_15024);
xnor U17139 (N_17139,N_15021,N_15217);
or U17140 (N_17140,N_15661,N_15719);
or U17141 (N_17141,N_15333,N_15296);
nand U17142 (N_17142,N_15201,N_15877);
nor U17143 (N_17143,N_15383,N_16207);
nand U17144 (N_17144,N_16054,N_15658);
and U17145 (N_17145,N_16230,N_16055);
xor U17146 (N_17146,N_15550,N_16210);
and U17147 (N_17147,N_15188,N_15325);
xor U17148 (N_17148,N_15051,N_16033);
nand U17149 (N_17149,N_15778,N_16176);
nor U17150 (N_17150,N_15174,N_15530);
nand U17151 (N_17151,N_15080,N_15776);
nand U17152 (N_17152,N_16017,N_15742);
nand U17153 (N_17153,N_16231,N_15054);
xor U17154 (N_17154,N_15674,N_15471);
nor U17155 (N_17155,N_16217,N_16156);
nor U17156 (N_17156,N_15553,N_15652);
or U17157 (N_17157,N_16206,N_15278);
xor U17158 (N_17158,N_15170,N_15907);
nand U17159 (N_17159,N_15705,N_15586);
or U17160 (N_17160,N_15678,N_15191);
nand U17161 (N_17161,N_16213,N_15819);
xnor U17162 (N_17162,N_15658,N_16232);
nor U17163 (N_17163,N_15382,N_15569);
xor U17164 (N_17164,N_15132,N_16105);
nor U17165 (N_17165,N_16080,N_15594);
and U17166 (N_17166,N_15645,N_15727);
nand U17167 (N_17167,N_15007,N_15510);
and U17168 (N_17168,N_15508,N_15250);
nor U17169 (N_17169,N_15820,N_16099);
and U17170 (N_17170,N_15092,N_15927);
nor U17171 (N_17171,N_15100,N_15517);
nor U17172 (N_17172,N_15532,N_16225);
xnor U17173 (N_17173,N_15691,N_16082);
nand U17174 (N_17174,N_15196,N_15485);
or U17175 (N_17175,N_15572,N_15723);
nor U17176 (N_17176,N_15609,N_15308);
nor U17177 (N_17177,N_15896,N_15400);
and U17178 (N_17178,N_15976,N_15279);
xnor U17179 (N_17179,N_15508,N_15193);
nor U17180 (N_17180,N_16159,N_16166);
nor U17181 (N_17181,N_15862,N_15860);
nor U17182 (N_17182,N_15206,N_15191);
nor U17183 (N_17183,N_15682,N_15536);
and U17184 (N_17184,N_15432,N_16185);
and U17185 (N_17185,N_15394,N_15380);
xnor U17186 (N_17186,N_15834,N_15420);
nand U17187 (N_17187,N_15358,N_15254);
nor U17188 (N_17188,N_15267,N_15685);
nand U17189 (N_17189,N_16163,N_15212);
nand U17190 (N_17190,N_15992,N_15202);
and U17191 (N_17191,N_15584,N_15286);
xnor U17192 (N_17192,N_16151,N_16140);
xnor U17193 (N_17193,N_16099,N_16074);
or U17194 (N_17194,N_15496,N_16239);
xor U17195 (N_17195,N_15647,N_16028);
nand U17196 (N_17196,N_15262,N_15254);
nor U17197 (N_17197,N_15364,N_16178);
or U17198 (N_17198,N_15464,N_15125);
and U17199 (N_17199,N_15718,N_15654);
or U17200 (N_17200,N_15132,N_15668);
xnor U17201 (N_17201,N_15208,N_15858);
xnor U17202 (N_17202,N_16195,N_15909);
and U17203 (N_17203,N_15616,N_15260);
and U17204 (N_17204,N_15532,N_15175);
nor U17205 (N_17205,N_15174,N_15831);
and U17206 (N_17206,N_16100,N_15571);
and U17207 (N_17207,N_15132,N_15623);
or U17208 (N_17208,N_15137,N_15405);
nor U17209 (N_17209,N_15379,N_15611);
and U17210 (N_17210,N_16236,N_15032);
and U17211 (N_17211,N_16065,N_15138);
nor U17212 (N_17212,N_15041,N_15136);
xor U17213 (N_17213,N_15053,N_15925);
nor U17214 (N_17214,N_15497,N_15037);
nor U17215 (N_17215,N_15960,N_15912);
and U17216 (N_17216,N_15863,N_16075);
xnor U17217 (N_17217,N_16023,N_16240);
and U17218 (N_17218,N_15290,N_15814);
and U17219 (N_17219,N_15063,N_16127);
nand U17220 (N_17220,N_15616,N_15217);
nand U17221 (N_17221,N_15533,N_15113);
nand U17222 (N_17222,N_15892,N_15637);
xor U17223 (N_17223,N_15859,N_15530);
nand U17224 (N_17224,N_15785,N_15758);
xor U17225 (N_17225,N_15386,N_15331);
or U17226 (N_17226,N_16083,N_15990);
or U17227 (N_17227,N_15779,N_15628);
and U17228 (N_17228,N_16026,N_15223);
xor U17229 (N_17229,N_15986,N_15242);
nand U17230 (N_17230,N_15093,N_15837);
nand U17231 (N_17231,N_16030,N_15591);
and U17232 (N_17232,N_15593,N_15871);
or U17233 (N_17233,N_15441,N_15744);
xnor U17234 (N_17234,N_15730,N_15237);
xor U17235 (N_17235,N_15629,N_15695);
nand U17236 (N_17236,N_15590,N_15112);
and U17237 (N_17237,N_15714,N_15887);
and U17238 (N_17238,N_15362,N_15309);
xor U17239 (N_17239,N_15323,N_15427);
or U17240 (N_17240,N_15755,N_15536);
or U17241 (N_17241,N_16204,N_15102);
and U17242 (N_17242,N_16203,N_15159);
and U17243 (N_17243,N_16203,N_15364);
or U17244 (N_17244,N_15878,N_15953);
and U17245 (N_17245,N_16185,N_15158);
nand U17246 (N_17246,N_15109,N_15506);
nand U17247 (N_17247,N_15649,N_15961);
or U17248 (N_17248,N_15112,N_16091);
xnor U17249 (N_17249,N_15523,N_15387);
nand U17250 (N_17250,N_16064,N_15771);
nand U17251 (N_17251,N_15802,N_15864);
and U17252 (N_17252,N_15808,N_15765);
and U17253 (N_17253,N_16139,N_15561);
nand U17254 (N_17254,N_16116,N_15467);
and U17255 (N_17255,N_16021,N_15931);
or U17256 (N_17256,N_16225,N_15193);
and U17257 (N_17257,N_15752,N_15940);
or U17258 (N_17258,N_16242,N_15683);
nor U17259 (N_17259,N_15004,N_15778);
and U17260 (N_17260,N_15224,N_15753);
xor U17261 (N_17261,N_15825,N_15412);
nand U17262 (N_17262,N_15664,N_15769);
nor U17263 (N_17263,N_15959,N_15057);
nand U17264 (N_17264,N_15894,N_15316);
or U17265 (N_17265,N_15659,N_15516);
nor U17266 (N_17266,N_15534,N_15515);
nor U17267 (N_17267,N_15417,N_15668);
and U17268 (N_17268,N_16094,N_15864);
nor U17269 (N_17269,N_16029,N_15034);
or U17270 (N_17270,N_15377,N_16035);
nand U17271 (N_17271,N_15181,N_15082);
nand U17272 (N_17272,N_15918,N_15811);
nor U17273 (N_17273,N_15764,N_15351);
nor U17274 (N_17274,N_15613,N_15896);
and U17275 (N_17275,N_15842,N_15717);
nor U17276 (N_17276,N_15711,N_16002);
nand U17277 (N_17277,N_15916,N_16111);
nor U17278 (N_17278,N_15581,N_15980);
and U17279 (N_17279,N_15791,N_15969);
or U17280 (N_17280,N_15429,N_15333);
xor U17281 (N_17281,N_15565,N_15436);
and U17282 (N_17282,N_16138,N_15343);
nand U17283 (N_17283,N_15582,N_15871);
nand U17284 (N_17284,N_15303,N_15419);
nand U17285 (N_17285,N_15107,N_15354);
xor U17286 (N_17286,N_16189,N_16046);
nor U17287 (N_17287,N_15281,N_15751);
nand U17288 (N_17288,N_15585,N_15415);
nand U17289 (N_17289,N_15487,N_15099);
nand U17290 (N_17290,N_15857,N_15303);
nand U17291 (N_17291,N_15867,N_15253);
or U17292 (N_17292,N_15141,N_15790);
xor U17293 (N_17293,N_15933,N_15231);
or U17294 (N_17294,N_15273,N_15775);
nand U17295 (N_17295,N_15667,N_16190);
xnor U17296 (N_17296,N_15287,N_15247);
xor U17297 (N_17297,N_15941,N_15328);
nor U17298 (N_17298,N_15622,N_15895);
or U17299 (N_17299,N_16051,N_15876);
or U17300 (N_17300,N_15863,N_15299);
or U17301 (N_17301,N_15319,N_15581);
nand U17302 (N_17302,N_15014,N_15737);
xor U17303 (N_17303,N_15759,N_15967);
nor U17304 (N_17304,N_15467,N_15839);
nor U17305 (N_17305,N_15693,N_15350);
or U17306 (N_17306,N_16150,N_15099);
nand U17307 (N_17307,N_16185,N_15597);
or U17308 (N_17308,N_15105,N_15058);
xor U17309 (N_17309,N_16217,N_15862);
xor U17310 (N_17310,N_15657,N_15180);
and U17311 (N_17311,N_15830,N_16010);
nand U17312 (N_17312,N_15989,N_15619);
xnor U17313 (N_17313,N_16134,N_15712);
or U17314 (N_17314,N_16223,N_15414);
xor U17315 (N_17315,N_16210,N_15061);
nand U17316 (N_17316,N_15004,N_15182);
or U17317 (N_17317,N_15664,N_16232);
xor U17318 (N_17318,N_15513,N_15163);
nor U17319 (N_17319,N_15827,N_15200);
and U17320 (N_17320,N_16244,N_15557);
nand U17321 (N_17321,N_16177,N_15752);
or U17322 (N_17322,N_15794,N_15302);
nor U17323 (N_17323,N_15637,N_15488);
nand U17324 (N_17324,N_15381,N_15156);
and U17325 (N_17325,N_15033,N_15733);
or U17326 (N_17326,N_15128,N_15110);
nor U17327 (N_17327,N_15340,N_15413);
xnor U17328 (N_17328,N_15172,N_15543);
xor U17329 (N_17329,N_15712,N_15707);
nor U17330 (N_17330,N_15383,N_16155);
xor U17331 (N_17331,N_15529,N_15494);
or U17332 (N_17332,N_15780,N_16107);
nand U17333 (N_17333,N_15936,N_16228);
nand U17334 (N_17334,N_15168,N_15773);
nor U17335 (N_17335,N_15892,N_15662);
xnor U17336 (N_17336,N_16205,N_15197);
xnor U17337 (N_17337,N_15664,N_15286);
nand U17338 (N_17338,N_16056,N_15763);
nor U17339 (N_17339,N_15811,N_15283);
xor U17340 (N_17340,N_15843,N_15429);
or U17341 (N_17341,N_16222,N_15281);
or U17342 (N_17342,N_15110,N_15590);
or U17343 (N_17343,N_15759,N_15287);
and U17344 (N_17344,N_15589,N_16014);
or U17345 (N_17345,N_15844,N_16014);
xnor U17346 (N_17346,N_15051,N_15697);
nand U17347 (N_17347,N_15409,N_15006);
nand U17348 (N_17348,N_15612,N_16104);
xor U17349 (N_17349,N_15145,N_15303);
xnor U17350 (N_17350,N_16216,N_15017);
nand U17351 (N_17351,N_15495,N_15036);
and U17352 (N_17352,N_15241,N_15109);
xnor U17353 (N_17353,N_15210,N_15119);
xnor U17354 (N_17354,N_15412,N_16239);
or U17355 (N_17355,N_15198,N_15086);
nor U17356 (N_17356,N_15747,N_15311);
nand U17357 (N_17357,N_15713,N_15452);
nor U17358 (N_17358,N_15917,N_15344);
nand U17359 (N_17359,N_15172,N_15495);
or U17360 (N_17360,N_15846,N_15806);
nor U17361 (N_17361,N_15396,N_15347);
xnor U17362 (N_17362,N_16231,N_16021);
nor U17363 (N_17363,N_15754,N_16012);
xor U17364 (N_17364,N_15345,N_16142);
and U17365 (N_17365,N_15577,N_15611);
nand U17366 (N_17366,N_15535,N_16040);
and U17367 (N_17367,N_15225,N_15764);
and U17368 (N_17368,N_15037,N_16183);
xor U17369 (N_17369,N_15469,N_15686);
and U17370 (N_17370,N_16020,N_15789);
nor U17371 (N_17371,N_15199,N_15308);
and U17372 (N_17372,N_15798,N_15283);
xor U17373 (N_17373,N_15896,N_15661);
nor U17374 (N_17374,N_15819,N_15829);
nor U17375 (N_17375,N_15956,N_16016);
nand U17376 (N_17376,N_16000,N_15686);
or U17377 (N_17377,N_15302,N_15372);
nor U17378 (N_17378,N_15180,N_16246);
nand U17379 (N_17379,N_15467,N_15588);
and U17380 (N_17380,N_15951,N_16047);
nor U17381 (N_17381,N_16061,N_15818);
and U17382 (N_17382,N_15008,N_15505);
or U17383 (N_17383,N_16107,N_16192);
and U17384 (N_17384,N_15817,N_15069);
nor U17385 (N_17385,N_16047,N_15303);
nor U17386 (N_17386,N_15844,N_15565);
and U17387 (N_17387,N_15809,N_15048);
and U17388 (N_17388,N_15319,N_15492);
nor U17389 (N_17389,N_16042,N_15339);
xnor U17390 (N_17390,N_16178,N_15095);
xor U17391 (N_17391,N_15559,N_15568);
nand U17392 (N_17392,N_15949,N_15914);
nand U17393 (N_17393,N_15001,N_15698);
xor U17394 (N_17394,N_16010,N_16054);
or U17395 (N_17395,N_16240,N_15576);
nor U17396 (N_17396,N_15385,N_15951);
nand U17397 (N_17397,N_16026,N_15629);
or U17398 (N_17398,N_15957,N_15384);
or U17399 (N_17399,N_15868,N_15808);
and U17400 (N_17400,N_15685,N_15427);
nand U17401 (N_17401,N_15547,N_15667);
and U17402 (N_17402,N_15643,N_15338);
nand U17403 (N_17403,N_15547,N_16096);
nor U17404 (N_17404,N_15377,N_15945);
and U17405 (N_17405,N_15417,N_15414);
nand U17406 (N_17406,N_15111,N_15242);
nor U17407 (N_17407,N_16093,N_16157);
nand U17408 (N_17408,N_15082,N_15964);
nand U17409 (N_17409,N_15452,N_16165);
xnor U17410 (N_17410,N_15088,N_16146);
nand U17411 (N_17411,N_15821,N_15313);
and U17412 (N_17412,N_15438,N_15603);
nand U17413 (N_17413,N_15513,N_15639);
nand U17414 (N_17414,N_15988,N_15342);
xnor U17415 (N_17415,N_15212,N_15007);
nand U17416 (N_17416,N_16143,N_15800);
xor U17417 (N_17417,N_15014,N_16123);
nor U17418 (N_17418,N_16247,N_15163);
xnor U17419 (N_17419,N_15928,N_15002);
or U17420 (N_17420,N_15988,N_15222);
and U17421 (N_17421,N_15223,N_15544);
or U17422 (N_17422,N_16111,N_15702);
nor U17423 (N_17423,N_15939,N_15172);
and U17424 (N_17424,N_16120,N_15420);
nor U17425 (N_17425,N_15382,N_15639);
nand U17426 (N_17426,N_15022,N_15495);
and U17427 (N_17427,N_15152,N_15062);
xor U17428 (N_17428,N_16006,N_16112);
or U17429 (N_17429,N_15192,N_15722);
or U17430 (N_17430,N_15544,N_15887);
and U17431 (N_17431,N_15849,N_15349);
xnor U17432 (N_17432,N_15934,N_15345);
nand U17433 (N_17433,N_16220,N_15166);
or U17434 (N_17434,N_15306,N_15297);
and U17435 (N_17435,N_16242,N_15489);
xnor U17436 (N_17436,N_15412,N_15358);
nor U17437 (N_17437,N_15934,N_16041);
or U17438 (N_17438,N_15925,N_15001);
or U17439 (N_17439,N_16103,N_16084);
nor U17440 (N_17440,N_15837,N_15479);
xor U17441 (N_17441,N_15261,N_15501);
or U17442 (N_17442,N_15153,N_15762);
nor U17443 (N_17443,N_15591,N_15063);
nand U17444 (N_17444,N_15345,N_15031);
xor U17445 (N_17445,N_15899,N_15453);
nand U17446 (N_17446,N_15147,N_15268);
xnor U17447 (N_17447,N_16015,N_15796);
or U17448 (N_17448,N_15077,N_15102);
nor U17449 (N_17449,N_15438,N_15983);
nor U17450 (N_17450,N_15538,N_15740);
or U17451 (N_17451,N_15918,N_15935);
nor U17452 (N_17452,N_15588,N_15917);
or U17453 (N_17453,N_15673,N_15927);
and U17454 (N_17454,N_15962,N_15194);
or U17455 (N_17455,N_15183,N_15939);
xor U17456 (N_17456,N_15020,N_15207);
xnor U17457 (N_17457,N_16029,N_15925);
nor U17458 (N_17458,N_16141,N_16200);
nor U17459 (N_17459,N_16063,N_15816);
and U17460 (N_17460,N_15222,N_15331);
or U17461 (N_17461,N_15285,N_16214);
nand U17462 (N_17462,N_16203,N_15030);
nand U17463 (N_17463,N_15660,N_16038);
xor U17464 (N_17464,N_15214,N_15878);
nand U17465 (N_17465,N_15396,N_15942);
nand U17466 (N_17466,N_15438,N_15925);
or U17467 (N_17467,N_15716,N_16154);
nand U17468 (N_17468,N_15593,N_15203);
and U17469 (N_17469,N_15945,N_15336);
and U17470 (N_17470,N_15048,N_15005);
nor U17471 (N_17471,N_15582,N_15911);
nor U17472 (N_17472,N_15756,N_15132);
or U17473 (N_17473,N_15984,N_15265);
or U17474 (N_17474,N_15865,N_16123);
or U17475 (N_17475,N_15729,N_15040);
nand U17476 (N_17476,N_16202,N_16139);
xnor U17477 (N_17477,N_15612,N_15499);
nand U17478 (N_17478,N_15392,N_15116);
and U17479 (N_17479,N_15233,N_15311);
or U17480 (N_17480,N_16207,N_15835);
nand U17481 (N_17481,N_15176,N_15440);
nor U17482 (N_17482,N_15485,N_15128);
nand U17483 (N_17483,N_15292,N_15633);
nand U17484 (N_17484,N_15182,N_15370);
and U17485 (N_17485,N_16085,N_15989);
nand U17486 (N_17486,N_15013,N_15530);
and U17487 (N_17487,N_15184,N_15346);
nor U17488 (N_17488,N_15697,N_15307);
nand U17489 (N_17489,N_16180,N_15901);
nand U17490 (N_17490,N_16188,N_16224);
nand U17491 (N_17491,N_15111,N_16030);
nand U17492 (N_17492,N_15175,N_15177);
xor U17493 (N_17493,N_15617,N_15975);
xor U17494 (N_17494,N_15231,N_15719);
xnor U17495 (N_17495,N_15526,N_15497);
nor U17496 (N_17496,N_15088,N_15333);
nand U17497 (N_17497,N_15491,N_15512);
or U17498 (N_17498,N_15717,N_15087);
or U17499 (N_17499,N_15758,N_15537);
and U17500 (N_17500,N_16250,N_17453);
and U17501 (N_17501,N_16607,N_17040);
nor U17502 (N_17502,N_17039,N_16588);
and U17503 (N_17503,N_17410,N_16757);
nand U17504 (N_17504,N_16458,N_16787);
and U17505 (N_17505,N_16831,N_16288);
xor U17506 (N_17506,N_17428,N_17141);
and U17507 (N_17507,N_17245,N_17229);
and U17508 (N_17508,N_16571,N_16775);
and U17509 (N_17509,N_16911,N_17430);
nor U17510 (N_17510,N_17236,N_16611);
nand U17511 (N_17511,N_16315,N_17452);
nand U17512 (N_17512,N_16445,N_16296);
and U17513 (N_17513,N_16529,N_17016);
or U17514 (N_17514,N_16271,N_16992);
xnor U17515 (N_17515,N_17263,N_17486);
nor U17516 (N_17516,N_17457,N_17252);
nor U17517 (N_17517,N_16374,N_17179);
nand U17518 (N_17518,N_16847,N_17015);
nor U17519 (N_17519,N_17495,N_17339);
nor U17520 (N_17520,N_16953,N_17001);
nor U17521 (N_17521,N_16566,N_17412);
or U17522 (N_17522,N_16455,N_17093);
xor U17523 (N_17523,N_17357,N_16679);
xnor U17524 (N_17524,N_16998,N_16686);
xnor U17525 (N_17525,N_16474,N_17019);
nor U17526 (N_17526,N_17456,N_16584);
or U17527 (N_17527,N_16748,N_16415);
and U17528 (N_17528,N_16676,N_16930);
nor U17529 (N_17529,N_16887,N_16378);
nor U17530 (N_17530,N_16821,N_16361);
xnor U17531 (N_17531,N_16610,N_17075);
or U17532 (N_17532,N_16964,N_17369);
nand U17533 (N_17533,N_16903,N_16535);
nor U17534 (N_17534,N_17087,N_16791);
nand U17535 (N_17535,N_16266,N_17132);
and U17536 (N_17536,N_17111,N_17069);
nand U17537 (N_17537,N_17354,N_16582);
xor U17538 (N_17538,N_16262,N_17246);
xnor U17539 (N_17539,N_16294,N_17090);
or U17540 (N_17540,N_16491,N_17206);
xnor U17541 (N_17541,N_17215,N_16870);
nor U17542 (N_17542,N_17288,N_16554);
nor U17543 (N_17543,N_17313,N_16800);
xor U17544 (N_17544,N_16954,N_17492);
xor U17545 (N_17545,N_16927,N_17408);
nand U17546 (N_17546,N_17064,N_17284);
nand U17547 (N_17547,N_16916,N_16331);
or U17548 (N_17548,N_16984,N_16934);
nor U17549 (N_17549,N_16359,N_17325);
and U17550 (N_17550,N_16343,N_16258);
or U17551 (N_17551,N_16555,N_17375);
xor U17552 (N_17552,N_17405,N_16742);
nor U17553 (N_17553,N_16569,N_16747);
nand U17554 (N_17554,N_16260,N_16345);
or U17555 (N_17555,N_16739,N_16762);
nand U17556 (N_17556,N_16808,N_16325);
nand U17557 (N_17557,N_16809,N_16841);
or U17558 (N_17558,N_16446,N_16444);
nand U17559 (N_17559,N_16840,N_16436);
and U17560 (N_17560,N_16560,N_17218);
xor U17561 (N_17561,N_16494,N_16558);
and U17562 (N_17562,N_16805,N_17210);
nor U17563 (N_17563,N_17362,N_16790);
xor U17564 (N_17564,N_16810,N_16307);
nor U17565 (N_17565,N_17280,N_17458);
nand U17566 (N_17566,N_16779,N_16682);
xor U17567 (N_17567,N_17371,N_16854);
or U17568 (N_17568,N_17131,N_16699);
nor U17569 (N_17569,N_17176,N_16941);
or U17570 (N_17570,N_16741,N_16386);
and U17571 (N_17571,N_17349,N_16586);
xor U17572 (N_17572,N_16990,N_17009);
or U17573 (N_17573,N_16372,N_17464);
nand U17574 (N_17574,N_16332,N_16253);
or U17575 (N_17575,N_16723,N_17341);
and U17576 (N_17576,N_16279,N_17343);
or U17577 (N_17577,N_16310,N_16306);
and U17578 (N_17578,N_16363,N_16837);
nor U17579 (N_17579,N_16512,N_16721);
and U17580 (N_17580,N_17347,N_16724);
nand U17581 (N_17581,N_16380,N_16393);
xnor U17582 (N_17582,N_16399,N_17007);
or U17583 (N_17583,N_17474,N_17227);
nand U17584 (N_17584,N_16872,N_16576);
or U17585 (N_17585,N_16362,N_17329);
xnor U17586 (N_17586,N_17145,N_16634);
and U17587 (N_17587,N_17134,N_16842);
and U17588 (N_17588,N_17471,N_16908);
or U17589 (N_17589,N_16567,N_17373);
and U17590 (N_17590,N_16983,N_16920);
nand U17591 (N_17591,N_16475,N_16285);
nor U17592 (N_17592,N_17482,N_16918);
or U17593 (N_17593,N_16957,N_17282);
nand U17594 (N_17594,N_16794,N_17038);
nand U17595 (N_17595,N_16778,N_17006);
nor U17596 (N_17596,N_17254,N_17196);
and U17597 (N_17597,N_16795,N_16848);
xnor U17598 (N_17598,N_16284,N_17139);
or U17599 (N_17599,N_17382,N_16740);
xor U17600 (N_17600,N_17310,N_16855);
or U17601 (N_17601,N_17045,N_16340);
xor U17602 (N_17602,N_16546,N_16632);
nand U17603 (N_17603,N_16355,N_16326);
or U17604 (N_17604,N_16521,N_16898);
and U17605 (N_17605,N_17480,N_16614);
and U17606 (N_17606,N_16267,N_17345);
xor U17607 (N_17607,N_16956,N_16901);
nand U17608 (N_17608,N_16511,N_16286);
nor U17609 (N_17609,N_17125,N_17175);
xnor U17610 (N_17610,N_16532,N_17380);
nand U17611 (N_17611,N_17183,N_16961);
nor U17612 (N_17612,N_17372,N_17063);
xor U17613 (N_17613,N_16348,N_17494);
and U17614 (N_17614,N_16976,N_17318);
nor U17615 (N_17615,N_17002,N_17414);
xor U17616 (N_17616,N_16594,N_17022);
and U17617 (N_17617,N_16568,N_17352);
or U17618 (N_17618,N_16827,N_17127);
or U17619 (N_17619,N_16995,N_17048);
xor U17620 (N_17620,N_17117,N_16471);
and U17621 (N_17621,N_16688,N_16498);
nor U17622 (N_17622,N_16892,N_16745);
nor U17623 (N_17623,N_17182,N_16598);
nand U17624 (N_17624,N_16596,N_16356);
nand U17625 (N_17625,N_16252,N_17261);
or U17626 (N_17626,N_16483,N_16549);
xor U17627 (N_17627,N_17023,N_17376);
xnor U17628 (N_17628,N_16557,N_16410);
nand U17629 (N_17629,N_17350,N_16493);
nor U17630 (N_17630,N_16371,N_17332);
nand U17631 (N_17631,N_17481,N_17485);
xor U17632 (N_17632,N_16899,N_17126);
or U17633 (N_17633,N_16578,N_16756);
and U17634 (N_17634,N_17459,N_17420);
nor U17635 (N_17635,N_16650,N_17162);
nand U17636 (N_17636,N_17450,N_16979);
nor U17637 (N_17637,N_16781,N_17271);
xor U17638 (N_17638,N_17181,N_17461);
nand U17639 (N_17639,N_17011,N_17230);
or U17640 (N_17640,N_16300,N_16696);
xor U17641 (N_17641,N_16966,N_17028);
or U17642 (N_17642,N_16950,N_17171);
nor U17643 (N_17643,N_16274,N_17305);
or U17644 (N_17644,N_17205,N_16864);
and U17645 (N_17645,N_17164,N_16702);
and U17646 (N_17646,N_17036,N_16352);
or U17647 (N_17647,N_16403,N_17423);
and U17648 (N_17648,N_17312,N_17455);
xor U17649 (N_17649,N_17129,N_16360);
and U17650 (N_17650,N_16605,N_16706);
or U17651 (N_17651,N_17327,N_17399);
nor U17652 (N_17652,N_16564,N_16323);
nor U17653 (N_17653,N_16651,N_17026);
and U17654 (N_17654,N_17356,N_16713);
xnor U17655 (N_17655,N_16725,N_16656);
xor U17656 (N_17656,N_17014,N_16814);
or U17657 (N_17657,N_16720,N_16318);
and U17658 (N_17658,N_16648,N_16381);
or U17659 (N_17659,N_17066,N_17214);
nor U17660 (N_17660,N_17498,N_16430);
xnor U17661 (N_17661,N_17276,N_16574);
or U17662 (N_17662,N_17118,N_16945);
nor U17663 (N_17663,N_17300,N_17225);
and U17664 (N_17664,N_17315,N_17438);
xnor U17665 (N_17665,N_17445,N_16324);
nand U17666 (N_17666,N_17272,N_16602);
nand U17667 (N_17667,N_17470,N_16653);
and U17668 (N_17668,N_16871,N_16665);
or U17669 (N_17669,N_17081,N_16959);
or U17670 (N_17670,N_17419,N_16726);
and U17671 (N_17671,N_17085,N_16658);
and U17672 (N_17672,N_17432,N_16543);
xnor U17673 (N_17673,N_16777,N_16495);
nand U17674 (N_17674,N_17355,N_16452);
nand U17675 (N_17675,N_17324,N_16928);
and U17676 (N_17676,N_17243,N_17381);
nand U17677 (N_17677,N_16910,N_17274);
nor U17678 (N_17678,N_16350,N_16283);
nor U17679 (N_17679,N_17003,N_17483);
nand U17680 (N_17680,N_16680,N_17377);
nor U17681 (N_17681,N_17448,N_16876);
nor U17682 (N_17682,N_16733,N_17267);
and U17683 (N_17683,N_17247,N_16638);
or U17684 (N_17684,N_16986,N_17397);
and U17685 (N_17685,N_17005,N_16375);
nand U17686 (N_17686,N_16572,N_16963);
and U17687 (N_17687,N_16339,N_16946);
nor U17688 (N_17688,N_17437,N_16631);
or U17689 (N_17689,N_16552,N_17366);
nor U17690 (N_17690,N_17042,N_16465);
and U17691 (N_17691,N_16832,N_16636);
nor U17692 (N_17692,N_16402,N_17216);
xnor U17693 (N_17693,N_16320,N_16712);
nor U17694 (N_17694,N_17010,N_17211);
nor U17695 (N_17695,N_16974,N_16701);
nor U17696 (N_17696,N_16268,N_16993);
nor U17697 (N_17697,N_17108,N_16657);
nand U17698 (N_17698,N_16691,N_16478);
or U17699 (N_17699,N_16878,N_17058);
nand U17700 (N_17700,N_16488,N_16698);
and U17701 (N_17701,N_16782,N_16763);
or U17702 (N_17702,N_16642,N_17079);
nor U17703 (N_17703,N_16639,N_16731);
nor U17704 (N_17704,N_17113,N_17078);
and U17705 (N_17705,N_16786,N_16528);
and U17706 (N_17706,N_17049,N_16978);
or U17707 (N_17707,N_16666,N_17298);
or U17708 (N_17708,N_17497,N_16811);
and U17709 (N_17709,N_17037,N_17008);
and U17710 (N_17710,N_16663,N_16802);
or U17711 (N_17711,N_16856,N_17477);
nor U17712 (N_17712,N_17364,N_16687);
or U17713 (N_17713,N_16853,N_17188);
and U17714 (N_17714,N_16487,N_16513);
or U17715 (N_17715,N_16463,N_17240);
nand U17716 (N_17716,N_16818,N_16735);
and U17717 (N_17717,N_17451,N_16886);
nor U17718 (N_17718,N_17409,N_17148);
nor U17719 (N_17719,N_17223,N_16600);
nand U17720 (N_17720,N_17353,N_16670);
or U17721 (N_17721,N_16477,N_17441);
and U17722 (N_17722,N_16281,N_17433);
nand U17723 (N_17723,N_16681,N_16538);
or U17724 (N_17724,N_16462,N_16767);
and U17725 (N_17725,N_16617,N_17499);
or U17726 (N_17726,N_16647,N_16729);
nand U17727 (N_17727,N_17207,N_17199);
and U17728 (N_17728,N_17031,N_17241);
nand U17729 (N_17729,N_17157,N_17187);
nand U17730 (N_17730,N_17476,N_16585);
xor U17731 (N_17731,N_16287,N_16931);
nor U17732 (N_17732,N_16627,N_16385);
nand U17733 (N_17733,N_16317,N_17209);
nand U17734 (N_17734,N_16620,N_17059);
or U17735 (N_17735,N_17434,N_17344);
nand U17736 (N_17736,N_17238,N_17073);
and U17737 (N_17737,N_17116,N_17086);
or U17738 (N_17738,N_16664,N_16705);
nand U17739 (N_17739,N_17004,N_17147);
or U17740 (N_17740,N_16710,N_16815);
xor U17741 (N_17741,N_17138,N_16982);
nor U17742 (N_17742,N_16316,N_16387);
nor U17743 (N_17743,N_16812,N_16575);
or U17744 (N_17744,N_16604,N_17463);
and U17745 (N_17745,N_16865,N_16660);
xnor U17746 (N_17746,N_16932,N_16866);
and U17747 (N_17747,N_17197,N_17255);
nor U17748 (N_17748,N_16635,N_16960);
and U17749 (N_17749,N_17386,N_17025);
xnor U17750 (N_17750,N_16761,N_16760);
or U17751 (N_17751,N_17424,N_17060);
nor U17752 (N_17752,N_17133,N_16440);
or U17753 (N_17753,N_16637,N_16829);
nand U17754 (N_17754,N_16629,N_16625);
or U17755 (N_17755,N_16771,N_16434);
nand U17756 (N_17756,N_17057,N_17226);
xor U17757 (N_17757,N_17264,N_16376);
and U17758 (N_17758,N_16533,N_16755);
and U17759 (N_17759,N_17319,N_17235);
and U17760 (N_17760,N_16879,N_16674);
xor U17761 (N_17761,N_16358,N_16860);
or U17762 (N_17762,N_17365,N_16796);
xnor U17763 (N_17763,N_16780,N_16351);
xnor U17764 (N_17764,N_17102,N_17442);
or U17765 (N_17765,N_16801,N_17416);
or U17766 (N_17766,N_16861,N_16254);
and U17767 (N_17767,N_16923,N_16717);
or U17768 (N_17768,N_16844,N_16412);
nor U17769 (N_17769,N_17328,N_16426);
xor U17770 (N_17770,N_16792,N_16828);
nor U17771 (N_17771,N_16369,N_17484);
and U17772 (N_17772,N_17061,N_16883);
nor U17773 (N_17773,N_16621,N_17123);
or U17774 (N_17774,N_16438,N_16321);
or U17775 (N_17775,N_17121,N_17249);
or U17776 (N_17776,N_17444,N_16481);
nor U17777 (N_17777,N_17262,N_16514);
or U17778 (N_17778,N_16633,N_16357);
xor U17779 (N_17779,N_16389,N_17435);
xor U17780 (N_17780,N_16873,N_17251);
xnor U17781 (N_17781,N_17391,N_17311);
nand U17782 (N_17782,N_16644,N_16365);
or U17783 (N_17783,N_16496,N_17100);
nor U17784 (N_17784,N_17359,N_17077);
nor U17785 (N_17785,N_17177,N_16383);
or U17786 (N_17786,N_17259,N_17018);
nand U17787 (N_17787,N_17170,N_17286);
nand U17788 (N_17788,N_17469,N_17233);
or U17789 (N_17789,N_17265,N_16599);
nor U17790 (N_17790,N_17035,N_17335);
and U17791 (N_17791,N_17370,N_17208);
or U17792 (N_17792,N_17200,N_16969);
xnor U17793 (N_17793,N_17232,N_17260);
nand U17794 (N_17794,N_16601,N_17289);
and U17795 (N_17795,N_16457,N_17417);
and U17796 (N_17796,N_16830,N_17443);
nor U17797 (N_17797,N_17460,N_16673);
nand U17798 (N_17798,N_16367,N_17248);
and U17799 (N_17799,N_16895,N_16373);
nand U17800 (N_17800,N_17168,N_17389);
or U17801 (N_17801,N_16943,N_16508);
and U17802 (N_17802,N_17192,N_16404);
xor U17803 (N_17803,N_17411,N_16540);
and U17804 (N_17804,N_16292,N_17447);
and U17805 (N_17805,N_16833,N_16988);
nand U17806 (N_17806,N_17098,N_16622);
or U17807 (N_17807,N_17337,N_17115);
xor U17808 (N_17808,N_17186,N_17052);
xor U17809 (N_17809,N_16275,N_16551);
nand U17810 (N_17810,N_16518,N_16991);
xor U17811 (N_17811,N_17072,N_16784);
or U17812 (N_17812,N_16309,N_17128);
and U17813 (N_17813,N_17468,N_16759);
or U17814 (N_17814,N_16291,N_16849);
and U17815 (N_17815,N_17479,N_17393);
nand U17816 (N_17816,N_16424,N_16384);
nor U17817 (N_17817,N_17074,N_17488);
and U17818 (N_17818,N_17150,N_16751);
nand U17819 (N_17819,N_16606,N_16377);
xor U17820 (N_17820,N_17095,N_16265);
nand U17821 (N_17821,N_17269,N_16803);
or U17822 (N_17822,N_17043,N_16523);
xnor U17823 (N_17823,N_16732,N_16989);
and U17824 (N_17824,N_17462,N_17270);
and U17825 (N_17825,N_16938,N_16947);
nor U17826 (N_17826,N_16845,N_16573);
nand U17827 (N_17827,N_16823,N_17153);
or U17828 (N_17828,N_16531,N_16580);
or U17829 (N_17829,N_16290,N_16550);
and U17830 (N_17830,N_16539,N_16587);
nor U17831 (N_17831,N_16347,N_17051);
nand U17832 (N_17832,N_16689,N_16530);
xnor U17833 (N_17833,N_16464,N_16394);
nor U17834 (N_17834,N_16263,N_17496);
or U17835 (N_17835,N_16429,N_17279);
xor U17836 (N_17836,N_16589,N_16863);
or U17837 (N_17837,N_16485,N_16968);
xnor U17838 (N_17838,N_16972,N_16486);
nand U17839 (N_17839,N_17114,N_16277);
nor U17840 (N_17840,N_16505,N_16851);
and U17841 (N_17841,N_16738,N_16659);
or U17842 (N_17842,N_17068,N_17472);
or U17843 (N_17843,N_16921,N_17234);
nor U17844 (N_17844,N_17383,N_16652);
xor U17845 (N_17845,N_16750,N_16894);
nand U17846 (N_17846,N_17440,N_17449);
nor U17847 (N_17847,N_17071,N_17169);
xnor U17848 (N_17848,N_17309,N_16264);
or U17849 (N_17849,N_16545,N_16718);
nor U17850 (N_17850,N_16473,N_16330);
nor U17851 (N_17851,N_17160,N_16994);
nor U17852 (N_17852,N_17155,N_17487);
and U17853 (N_17853,N_16461,N_17213);
xor U17854 (N_17854,N_16447,N_16685);
or U17855 (N_17855,N_16337,N_16454);
xnor U17856 (N_17856,N_16562,N_17146);
nand U17857 (N_17857,N_16472,N_16527);
nand U17858 (N_17858,N_16534,N_17358);
xor U17859 (N_17859,N_17466,N_16619);
nand U17860 (N_17860,N_17094,N_16924);
and U17861 (N_17861,N_16907,N_16926);
and U17862 (N_17862,N_16734,N_16875);
or U17863 (N_17863,N_17439,N_16768);
xor U17864 (N_17864,N_16368,N_17221);
nand U17865 (N_17865,N_17159,N_16769);
and U17866 (N_17866,N_16765,N_17403);
or U17867 (N_17867,N_17422,N_16366);
nor U17868 (N_17868,N_17379,N_16379);
or U17869 (N_17869,N_16382,N_17275);
nor U17870 (N_17870,N_16344,N_17120);
xnor U17871 (N_17871,N_16719,N_17110);
or U17872 (N_17872,N_17491,N_16502);
nand U17873 (N_17873,N_16406,N_16824);
or U17874 (N_17874,N_17316,N_17388);
nor U17875 (N_17875,N_16933,N_16793);
xor U17876 (N_17876,N_16697,N_16459);
nor U17877 (N_17877,N_16515,N_17489);
and U17878 (N_17878,N_16418,N_16859);
nand U17879 (N_17879,N_16411,N_17180);
nand U17880 (N_17880,N_16925,N_16868);
and U17881 (N_17881,N_17107,N_16997);
nor U17882 (N_17882,N_16728,N_16655);
nand U17883 (N_17883,N_16590,N_17222);
or U17884 (N_17884,N_16788,N_16401);
and U17885 (N_17885,N_16407,N_16749);
nor U17886 (N_17886,N_16958,N_17163);
nand U17887 (N_17887,N_16419,N_16613);
xnor U17888 (N_17888,N_16730,N_16423);
nand U17889 (N_17889,N_16690,N_17030);
xor U17890 (N_17890,N_16583,N_16603);
or U17891 (N_17891,N_16985,N_17307);
xnor U17892 (N_17892,N_17446,N_17425);
and U17893 (N_17893,N_17166,N_16906);
or U17894 (N_17894,N_16479,N_16354);
nor U17895 (N_17895,N_16789,N_16295);
nor U17896 (N_17896,N_17290,N_16507);
or U17897 (N_17897,N_17143,N_16816);
and U17898 (N_17898,N_16737,N_17088);
or U17899 (N_17899,N_17224,N_16846);
nand U17900 (N_17900,N_17340,N_17415);
xor U17901 (N_17901,N_17253,N_16559);
and U17902 (N_17902,N_16396,N_16707);
nand U17903 (N_17903,N_16524,N_16333);
xnor U17904 (N_17904,N_16885,N_17101);
xnor U17905 (N_17905,N_17473,N_17135);
nor U17906 (N_17906,N_16677,N_16302);
or U17907 (N_17907,N_16301,N_16743);
nand U17908 (N_17908,N_17277,N_16962);
or U17909 (N_17909,N_17070,N_16807);
or U17910 (N_17910,N_17122,N_16987);
or U17911 (N_17911,N_16500,N_16497);
or U17912 (N_17912,N_16643,N_16970);
xnor U17913 (N_17913,N_17154,N_17326);
and U17914 (N_17914,N_17217,N_16826);
and U17915 (N_17915,N_16304,N_17161);
xor U17916 (N_17916,N_16476,N_16646);
nor U17917 (N_17917,N_16563,N_17055);
nor U17918 (N_17918,N_17395,N_17368);
nand U17919 (N_17919,N_16525,N_16273);
or U17920 (N_17920,N_16822,N_16715);
and U17921 (N_17921,N_16700,N_16744);
or U17922 (N_17922,N_17124,N_16276);
nand U17923 (N_17923,N_16595,N_17401);
and U17924 (N_17924,N_16764,N_16900);
or U17925 (N_17925,N_16397,N_16915);
xnor U17926 (N_17926,N_16427,N_17000);
nor U17927 (N_17927,N_16882,N_16722);
xor U17928 (N_17928,N_16547,N_16692);
or U17929 (N_17929,N_17297,N_16819);
xnor U17930 (N_17930,N_16467,N_17062);
and U17931 (N_17931,N_16649,N_17109);
xnor U17932 (N_17932,N_16694,N_17191);
nor U17933 (N_17933,N_16322,N_16683);
nand U17934 (N_17934,N_16869,N_16261);
nand U17935 (N_17935,N_16952,N_16449);
and U17936 (N_17936,N_16668,N_16570);
nor U17937 (N_17937,N_16392,N_17119);
nand U17938 (N_17938,N_17195,N_16289);
xnor U17939 (N_17939,N_16929,N_17091);
and U17940 (N_17940,N_16902,N_16951);
xor U17941 (N_17941,N_17454,N_17407);
xor U17942 (N_17942,N_16667,N_17156);
or U17943 (N_17943,N_16770,N_16612);
or U17944 (N_17944,N_16443,N_16398);
nor U17945 (N_17945,N_17065,N_17103);
nor U17946 (N_17946,N_16334,N_16618);
and U17947 (N_17947,N_16338,N_17152);
or U17948 (N_17948,N_17292,N_16400);
or U17949 (N_17949,N_16413,N_16797);
nand U17950 (N_17950,N_16433,N_16935);
nor U17951 (N_17951,N_16858,N_17304);
or U17952 (N_17952,N_16517,N_16949);
xor U17953 (N_17953,N_17220,N_17258);
nor U17954 (N_17954,N_17273,N_16272);
and U17955 (N_17955,N_17193,N_17418);
nor U17956 (N_17956,N_16884,N_16752);
or U17957 (N_17957,N_17080,N_17140);
xor U17958 (N_17958,N_17097,N_16942);
nand U17959 (N_17959,N_16624,N_16391);
nor U17960 (N_17960,N_17257,N_16628);
xor U17961 (N_17961,N_17020,N_17174);
nor U17962 (N_17962,N_16813,N_17167);
nand U17963 (N_17963,N_17212,N_16311);
and U17964 (N_17964,N_16695,N_17396);
nand U17965 (N_17965,N_16758,N_16675);
and U17966 (N_17966,N_16503,N_17266);
and U17967 (N_17967,N_16255,N_16460);
and U17968 (N_17968,N_16838,N_16936);
and U17969 (N_17969,N_16798,N_16684);
nand U17970 (N_17970,N_16280,N_16510);
nor U17971 (N_17971,N_17244,N_17321);
xnor U17972 (N_17972,N_16880,N_16727);
nand U17973 (N_17973,N_17320,N_16336);
nor U17974 (N_17974,N_16329,N_17178);
xor U17975 (N_17975,N_16482,N_16919);
xnor U17976 (N_17976,N_16672,N_16428);
and U17977 (N_17977,N_16640,N_17322);
nand U17978 (N_17978,N_16470,N_16616);
xnor U17979 (N_17979,N_16857,N_16509);
nand U17980 (N_17980,N_16328,N_16425);
nor U17981 (N_17981,N_16897,N_17190);
xor U17982 (N_17982,N_16492,N_16506);
nor U17983 (N_17983,N_16422,N_17041);
or U17984 (N_17984,N_17165,N_17427);
nand U17985 (N_17985,N_17392,N_16693);
xor U17986 (N_17986,N_16999,N_17294);
or U17987 (N_17987,N_16314,N_16349);
and U17988 (N_17988,N_16981,N_16917);
and U17989 (N_17989,N_17105,N_16421);
xnor U17990 (N_17990,N_16395,N_16416);
or U17991 (N_17991,N_17421,N_17490);
or U17992 (N_17992,N_16980,N_16913);
xor U17993 (N_17993,N_16904,N_16912);
or U17994 (N_17994,N_16626,N_17374);
nand U17995 (N_17995,N_16877,N_16453);
xnor U17996 (N_17996,N_17185,N_16537);
nor U17997 (N_17997,N_16327,N_16716);
or U17998 (N_17998,N_17184,N_17151);
nand U17999 (N_17999,N_16703,N_16390);
nor U18000 (N_18000,N_17099,N_17398);
or U18001 (N_18001,N_17172,N_17346);
xor U18002 (N_18002,N_17295,N_17402);
or U18003 (N_18003,N_17198,N_16937);
xnor U18004 (N_18004,N_16714,N_16776);
xnor U18005 (N_18005,N_16364,N_16592);
nor U18006 (N_18006,N_16519,N_16967);
xnor U18007 (N_18007,N_17283,N_17426);
or U18008 (N_18008,N_17342,N_16746);
xor U18009 (N_18009,N_16293,N_17334);
or U18010 (N_18010,N_17330,N_17201);
and U18011 (N_18011,N_17360,N_16939);
and U18012 (N_18012,N_16388,N_17351);
or U18013 (N_18013,N_17308,N_16893);
xor U18014 (N_18014,N_16298,N_16581);
nor U18015 (N_18015,N_16548,N_16420);
xor U18016 (N_18016,N_16480,N_16773);
nor U18017 (N_18017,N_17204,N_17256);
and U18018 (N_18018,N_17306,N_16278);
or U18019 (N_18019,N_16645,N_16704);
nor U18020 (N_18020,N_16820,N_16955);
xnor U18021 (N_18021,N_17384,N_16662);
or U18022 (N_18022,N_17385,N_16591);
xnor U18023 (N_18023,N_16414,N_16468);
nor U18024 (N_18024,N_16504,N_16909);
xor U18025 (N_18025,N_17149,N_16774);
or U18026 (N_18026,N_17189,N_17056);
nand U18027 (N_18027,N_16565,N_16839);
or U18028 (N_18028,N_17478,N_16442);
nor U18029 (N_18029,N_17436,N_16448);
or U18030 (N_18030,N_16862,N_17285);
nor U18031 (N_18031,N_17012,N_16437);
or U18032 (N_18032,N_16678,N_17219);
nand U18033 (N_18033,N_17046,N_17047);
nand U18034 (N_18034,N_16753,N_17013);
or U18035 (N_18035,N_17239,N_16541);
nand U18036 (N_18036,N_17034,N_17323);
nor U18037 (N_18037,N_16914,N_16708);
xnor U18038 (N_18038,N_17024,N_16405);
nand U18039 (N_18039,N_17076,N_16944);
nand U18040 (N_18040,N_17050,N_16711);
nand U18041 (N_18041,N_16466,N_17331);
xor U18042 (N_18042,N_16450,N_17429);
nor U18043 (N_18043,N_17202,N_17338);
xnor U18044 (N_18044,N_17021,N_16654);
or U18045 (N_18045,N_17296,N_16516);
and U18046 (N_18046,N_16905,N_17082);
or U18047 (N_18047,N_17336,N_16522);
and U18048 (N_18048,N_17106,N_16432);
xor U18049 (N_18049,N_16843,N_16825);
or U18050 (N_18050,N_17092,N_16269);
nor U18051 (N_18051,N_16305,N_16259);
nor U18052 (N_18052,N_17029,N_17173);
and U18053 (N_18053,N_17465,N_16874);
or U18054 (N_18054,N_17228,N_16597);
nand U18055 (N_18055,N_17137,N_16973);
nand U18056 (N_18056,N_16520,N_16661);
xnor U18057 (N_18057,N_17291,N_16456);
nor U18058 (N_18058,N_17302,N_17493);
or U18059 (N_18059,N_16888,N_17431);
nor U18060 (N_18060,N_16671,N_17278);
and U18061 (N_18061,N_16439,N_17083);
nand U18062 (N_18062,N_17237,N_17467);
and U18063 (N_18063,N_17281,N_17367);
nor U18064 (N_18064,N_17194,N_17017);
nand U18065 (N_18065,N_17130,N_17299);
nand U18066 (N_18066,N_17390,N_16451);
nor U18067 (N_18067,N_16353,N_16501);
and U18068 (N_18068,N_17142,N_16256);
xor U18069 (N_18069,N_16754,N_17104);
xor U18070 (N_18070,N_17033,N_17293);
and U18071 (N_18071,N_16896,N_16785);
nand U18072 (N_18072,N_17400,N_16889);
and U18073 (N_18073,N_16556,N_17314);
and U18074 (N_18074,N_16852,N_16409);
nand U18075 (N_18075,N_16608,N_16641);
and U18076 (N_18076,N_17363,N_16346);
nor U18077 (N_18077,N_17096,N_17394);
xor U18078 (N_18078,N_17054,N_16526);
nor U18079 (N_18079,N_16579,N_16577);
xnor U18080 (N_18080,N_17303,N_16490);
nand U18081 (N_18081,N_16303,N_17404);
xor U18082 (N_18082,N_17032,N_16850);
or U18083 (N_18083,N_16561,N_16544);
nor U18084 (N_18084,N_16881,N_16536);
or U18085 (N_18085,N_16891,N_16593);
xnor U18086 (N_18086,N_16996,N_16799);
nor U18087 (N_18087,N_17112,N_16971);
nand U18088 (N_18088,N_17144,N_16922);
xnor U18089 (N_18089,N_17067,N_16297);
xnor U18090 (N_18090,N_16806,N_17348);
nand U18091 (N_18091,N_17242,N_16313);
xor U18092 (N_18092,N_17158,N_16299);
xnor U18093 (N_18093,N_16335,N_16431);
nand U18094 (N_18094,N_16609,N_16615);
and U18095 (N_18095,N_17333,N_16417);
nor U18096 (N_18096,N_17413,N_17136);
xnor U18097 (N_18097,N_16835,N_16867);
nor U18098 (N_18098,N_16817,N_17027);
nor U18099 (N_18099,N_17387,N_16499);
and U18100 (N_18100,N_17378,N_16469);
nand U18101 (N_18101,N_16975,N_16977);
nor U18102 (N_18102,N_16630,N_16312);
and U18103 (N_18103,N_16257,N_16669);
nand U18104 (N_18104,N_16251,N_16836);
xnor U18105 (N_18105,N_17084,N_16308);
nor U18106 (N_18106,N_16489,N_17250);
xor U18107 (N_18107,N_17203,N_16370);
and U18108 (N_18108,N_16441,N_17268);
nor U18109 (N_18109,N_17053,N_17287);
nand U18110 (N_18110,N_16940,N_16965);
nor U18111 (N_18111,N_16623,N_16890);
and U18112 (N_18112,N_17044,N_16553);
nand U18113 (N_18113,N_16766,N_16948);
nand U18114 (N_18114,N_16783,N_16282);
nor U18115 (N_18115,N_16834,N_16542);
nor U18116 (N_18116,N_16484,N_17231);
nor U18117 (N_18117,N_16319,N_17406);
or U18118 (N_18118,N_16341,N_16408);
nand U18119 (N_18119,N_16709,N_17301);
nand U18120 (N_18120,N_16772,N_17089);
xnor U18121 (N_18121,N_17475,N_16804);
or U18122 (N_18122,N_16736,N_17317);
xor U18123 (N_18123,N_16435,N_16270);
nor U18124 (N_18124,N_17361,N_16342);
nor U18125 (N_18125,N_16519,N_17282);
and U18126 (N_18126,N_16425,N_17003);
nor U18127 (N_18127,N_16365,N_16612);
or U18128 (N_18128,N_17100,N_16385);
or U18129 (N_18129,N_17166,N_16630);
or U18130 (N_18130,N_17257,N_16442);
xor U18131 (N_18131,N_16970,N_16257);
and U18132 (N_18132,N_17014,N_16830);
nor U18133 (N_18133,N_17218,N_16431);
xnor U18134 (N_18134,N_17115,N_16442);
xor U18135 (N_18135,N_16288,N_17306);
and U18136 (N_18136,N_17031,N_17476);
or U18137 (N_18137,N_16464,N_16736);
and U18138 (N_18138,N_16297,N_17413);
nand U18139 (N_18139,N_16268,N_17405);
xor U18140 (N_18140,N_17260,N_16616);
and U18141 (N_18141,N_16382,N_17201);
nor U18142 (N_18142,N_16669,N_16892);
nand U18143 (N_18143,N_16857,N_17125);
nand U18144 (N_18144,N_17397,N_17112);
nand U18145 (N_18145,N_17054,N_16748);
nor U18146 (N_18146,N_16917,N_16681);
nand U18147 (N_18147,N_16730,N_16926);
nand U18148 (N_18148,N_16629,N_16672);
or U18149 (N_18149,N_17225,N_16289);
nand U18150 (N_18150,N_17067,N_16736);
and U18151 (N_18151,N_17130,N_17094);
nor U18152 (N_18152,N_16575,N_16348);
nor U18153 (N_18153,N_17279,N_16949);
nand U18154 (N_18154,N_16745,N_17446);
or U18155 (N_18155,N_17385,N_16959);
xnor U18156 (N_18156,N_16922,N_16522);
nor U18157 (N_18157,N_17100,N_17276);
and U18158 (N_18158,N_16766,N_16485);
xnor U18159 (N_18159,N_17276,N_17003);
nand U18160 (N_18160,N_16718,N_17474);
or U18161 (N_18161,N_16436,N_16532);
xor U18162 (N_18162,N_17290,N_16805);
nand U18163 (N_18163,N_16706,N_16554);
nand U18164 (N_18164,N_17303,N_16349);
or U18165 (N_18165,N_17202,N_16293);
xor U18166 (N_18166,N_17248,N_17360);
nand U18167 (N_18167,N_16945,N_16842);
or U18168 (N_18168,N_17095,N_17318);
or U18169 (N_18169,N_16771,N_17267);
nand U18170 (N_18170,N_17451,N_17362);
or U18171 (N_18171,N_16567,N_16783);
or U18172 (N_18172,N_17056,N_16567);
nor U18173 (N_18173,N_16816,N_16398);
xor U18174 (N_18174,N_17034,N_17393);
xnor U18175 (N_18175,N_17301,N_16436);
xor U18176 (N_18176,N_16490,N_17373);
and U18177 (N_18177,N_16338,N_16372);
or U18178 (N_18178,N_17318,N_16906);
xor U18179 (N_18179,N_17394,N_16544);
nor U18180 (N_18180,N_17484,N_17105);
nand U18181 (N_18181,N_17028,N_16863);
xor U18182 (N_18182,N_17445,N_16351);
and U18183 (N_18183,N_17115,N_17101);
nor U18184 (N_18184,N_17308,N_16850);
or U18185 (N_18185,N_17010,N_17290);
nand U18186 (N_18186,N_16363,N_16721);
and U18187 (N_18187,N_16441,N_17456);
and U18188 (N_18188,N_16304,N_16770);
nor U18189 (N_18189,N_16794,N_16874);
nor U18190 (N_18190,N_16803,N_16605);
or U18191 (N_18191,N_16790,N_17112);
and U18192 (N_18192,N_17097,N_16472);
nor U18193 (N_18193,N_17233,N_16797);
or U18194 (N_18194,N_16665,N_17265);
and U18195 (N_18195,N_16929,N_16925);
nand U18196 (N_18196,N_17082,N_17037);
and U18197 (N_18197,N_16284,N_16965);
and U18198 (N_18198,N_16400,N_16706);
nor U18199 (N_18199,N_16796,N_17371);
nand U18200 (N_18200,N_17088,N_17129);
nor U18201 (N_18201,N_16747,N_16920);
and U18202 (N_18202,N_17174,N_17085);
or U18203 (N_18203,N_17219,N_16932);
xnor U18204 (N_18204,N_17346,N_17385);
and U18205 (N_18205,N_16707,N_16449);
xor U18206 (N_18206,N_16404,N_17117);
nand U18207 (N_18207,N_16783,N_16646);
and U18208 (N_18208,N_16362,N_16305);
or U18209 (N_18209,N_16676,N_17178);
nand U18210 (N_18210,N_16939,N_17211);
and U18211 (N_18211,N_16991,N_16257);
xnor U18212 (N_18212,N_17336,N_16342);
xnor U18213 (N_18213,N_16906,N_16576);
xnor U18214 (N_18214,N_17460,N_16367);
and U18215 (N_18215,N_17300,N_16429);
or U18216 (N_18216,N_16258,N_17365);
and U18217 (N_18217,N_17452,N_16368);
nor U18218 (N_18218,N_16754,N_16305);
nor U18219 (N_18219,N_16489,N_16396);
and U18220 (N_18220,N_16896,N_16670);
nor U18221 (N_18221,N_16703,N_16968);
xor U18222 (N_18222,N_16987,N_16737);
and U18223 (N_18223,N_16547,N_17099);
xnor U18224 (N_18224,N_17148,N_16996);
xnor U18225 (N_18225,N_16343,N_17067);
and U18226 (N_18226,N_16813,N_17473);
nor U18227 (N_18227,N_17173,N_16751);
or U18228 (N_18228,N_16493,N_17222);
nor U18229 (N_18229,N_17484,N_16397);
or U18230 (N_18230,N_16844,N_16781);
nor U18231 (N_18231,N_17150,N_17398);
xnor U18232 (N_18232,N_17294,N_17013);
nand U18233 (N_18233,N_17075,N_16736);
and U18234 (N_18234,N_16762,N_16299);
nor U18235 (N_18235,N_16710,N_17339);
and U18236 (N_18236,N_17024,N_16346);
and U18237 (N_18237,N_16561,N_16522);
or U18238 (N_18238,N_16756,N_17257);
nand U18239 (N_18239,N_16829,N_16827);
nor U18240 (N_18240,N_16658,N_17057);
nor U18241 (N_18241,N_16637,N_17476);
nand U18242 (N_18242,N_16575,N_17097);
nor U18243 (N_18243,N_17063,N_17296);
xnor U18244 (N_18244,N_16417,N_16409);
nand U18245 (N_18245,N_16477,N_17219);
and U18246 (N_18246,N_16356,N_16739);
or U18247 (N_18247,N_16714,N_17254);
xnor U18248 (N_18248,N_17105,N_17358);
and U18249 (N_18249,N_16963,N_16768);
and U18250 (N_18250,N_17032,N_16557);
nor U18251 (N_18251,N_17156,N_16311);
xnor U18252 (N_18252,N_17264,N_16469);
or U18253 (N_18253,N_17284,N_16650);
nor U18254 (N_18254,N_16431,N_16424);
and U18255 (N_18255,N_16909,N_17443);
xor U18256 (N_18256,N_16901,N_16934);
and U18257 (N_18257,N_16254,N_17242);
nor U18258 (N_18258,N_16443,N_16969);
xnor U18259 (N_18259,N_16862,N_17493);
nor U18260 (N_18260,N_16576,N_17309);
nand U18261 (N_18261,N_17115,N_17005);
nor U18262 (N_18262,N_16276,N_16968);
or U18263 (N_18263,N_16411,N_16790);
or U18264 (N_18264,N_16393,N_17374);
nor U18265 (N_18265,N_16338,N_16588);
nand U18266 (N_18266,N_16338,N_17364);
xnor U18267 (N_18267,N_16808,N_17281);
nand U18268 (N_18268,N_16335,N_17432);
nor U18269 (N_18269,N_17307,N_16791);
nand U18270 (N_18270,N_16398,N_16418);
nor U18271 (N_18271,N_16702,N_16844);
nand U18272 (N_18272,N_17434,N_17241);
nor U18273 (N_18273,N_17172,N_17134);
nor U18274 (N_18274,N_17293,N_17481);
nor U18275 (N_18275,N_16580,N_16539);
nor U18276 (N_18276,N_16510,N_17355);
nand U18277 (N_18277,N_17450,N_16996);
and U18278 (N_18278,N_16353,N_17234);
nor U18279 (N_18279,N_17020,N_16899);
and U18280 (N_18280,N_17194,N_17356);
xnor U18281 (N_18281,N_16462,N_17463);
or U18282 (N_18282,N_17160,N_17194);
xor U18283 (N_18283,N_16353,N_16548);
xor U18284 (N_18284,N_17264,N_17253);
xnor U18285 (N_18285,N_17148,N_16951);
and U18286 (N_18286,N_16391,N_17154);
nor U18287 (N_18287,N_16555,N_16973);
and U18288 (N_18288,N_17426,N_16259);
xor U18289 (N_18289,N_17468,N_16884);
nor U18290 (N_18290,N_16602,N_16859);
nor U18291 (N_18291,N_16917,N_17073);
or U18292 (N_18292,N_16664,N_17421);
nand U18293 (N_18293,N_17352,N_16882);
or U18294 (N_18294,N_16790,N_16612);
nand U18295 (N_18295,N_17192,N_16773);
nor U18296 (N_18296,N_16527,N_16494);
xor U18297 (N_18297,N_16435,N_16749);
xnor U18298 (N_18298,N_16962,N_16683);
xor U18299 (N_18299,N_16933,N_16315);
nand U18300 (N_18300,N_16645,N_17086);
nand U18301 (N_18301,N_17299,N_16959);
or U18302 (N_18302,N_16838,N_17414);
or U18303 (N_18303,N_16322,N_17348);
nor U18304 (N_18304,N_16653,N_17413);
xnor U18305 (N_18305,N_17368,N_16878);
nor U18306 (N_18306,N_17444,N_16939);
or U18307 (N_18307,N_17390,N_16579);
and U18308 (N_18308,N_17429,N_16381);
nand U18309 (N_18309,N_16628,N_16481);
nand U18310 (N_18310,N_16547,N_17241);
nand U18311 (N_18311,N_16979,N_16500);
nor U18312 (N_18312,N_17370,N_16291);
nor U18313 (N_18313,N_17215,N_17112);
nand U18314 (N_18314,N_16983,N_16761);
and U18315 (N_18315,N_16342,N_16308);
nand U18316 (N_18316,N_16749,N_16891);
xor U18317 (N_18317,N_16272,N_16903);
or U18318 (N_18318,N_16651,N_17322);
and U18319 (N_18319,N_16301,N_17104);
nor U18320 (N_18320,N_17256,N_16532);
nor U18321 (N_18321,N_17449,N_16357);
xnor U18322 (N_18322,N_17122,N_16760);
or U18323 (N_18323,N_16471,N_17301);
or U18324 (N_18324,N_17248,N_17210);
or U18325 (N_18325,N_17446,N_16943);
xnor U18326 (N_18326,N_16258,N_16376);
and U18327 (N_18327,N_16997,N_17198);
nor U18328 (N_18328,N_16834,N_17062);
xor U18329 (N_18329,N_17169,N_16830);
and U18330 (N_18330,N_17144,N_16478);
or U18331 (N_18331,N_16953,N_17285);
xnor U18332 (N_18332,N_16567,N_16506);
nor U18333 (N_18333,N_17344,N_16767);
or U18334 (N_18334,N_16610,N_16606);
nand U18335 (N_18335,N_17227,N_16659);
and U18336 (N_18336,N_17220,N_17095);
or U18337 (N_18337,N_16753,N_16268);
and U18338 (N_18338,N_17460,N_16878);
and U18339 (N_18339,N_16322,N_16649);
nor U18340 (N_18340,N_16533,N_16821);
or U18341 (N_18341,N_17377,N_16574);
nand U18342 (N_18342,N_17301,N_16547);
and U18343 (N_18343,N_17446,N_17015);
and U18344 (N_18344,N_16334,N_16399);
and U18345 (N_18345,N_16833,N_16875);
xnor U18346 (N_18346,N_16644,N_16920);
nand U18347 (N_18347,N_17402,N_16336);
and U18348 (N_18348,N_16602,N_17067);
or U18349 (N_18349,N_16609,N_16291);
nor U18350 (N_18350,N_16473,N_16622);
nor U18351 (N_18351,N_16321,N_17335);
or U18352 (N_18352,N_16411,N_17242);
xnor U18353 (N_18353,N_16327,N_16341);
or U18354 (N_18354,N_17275,N_16828);
xnor U18355 (N_18355,N_16404,N_16312);
or U18356 (N_18356,N_17321,N_16638);
or U18357 (N_18357,N_17278,N_16695);
nor U18358 (N_18358,N_16731,N_17077);
nand U18359 (N_18359,N_16851,N_17046);
nor U18360 (N_18360,N_16575,N_16616);
xor U18361 (N_18361,N_17132,N_16502);
nand U18362 (N_18362,N_16951,N_16486);
and U18363 (N_18363,N_16842,N_17083);
or U18364 (N_18364,N_16748,N_16868);
xor U18365 (N_18365,N_16791,N_16877);
and U18366 (N_18366,N_16318,N_16639);
and U18367 (N_18367,N_16439,N_16256);
and U18368 (N_18368,N_17281,N_16859);
nand U18369 (N_18369,N_16909,N_17376);
nor U18370 (N_18370,N_16792,N_17287);
nand U18371 (N_18371,N_16841,N_16862);
nor U18372 (N_18372,N_17388,N_16626);
or U18373 (N_18373,N_17078,N_17020);
nor U18374 (N_18374,N_16830,N_16424);
and U18375 (N_18375,N_17477,N_17255);
or U18376 (N_18376,N_16558,N_16776);
xor U18377 (N_18377,N_17441,N_16955);
nand U18378 (N_18378,N_17091,N_16713);
nand U18379 (N_18379,N_17188,N_17091);
xor U18380 (N_18380,N_17419,N_16930);
nor U18381 (N_18381,N_16819,N_17280);
and U18382 (N_18382,N_16257,N_17027);
nand U18383 (N_18383,N_17321,N_17222);
nand U18384 (N_18384,N_17168,N_16820);
or U18385 (N_18385,N_17275,N_17240);
nand U18386 (N_18386,N_16257,N_16894);
and U18387 (N_18387,N_17127,N_16918);
xor U18388 (N_18388,N_17330,N_16463);
nor U18389 (N_18389,N_17463,N_16341);
and U18390 (N_18390,N_17315,N_16341);
and U18391 (N_18391,N_17249,N_17454);
and U18392 (N_18392,N_17002,N_17336);
or U18393 (N_18393,N_16282,N_16697);
xnor U18394 (N_18394,N_17076,N_17411);
nor U18395 (N_18395,N_16934,N_17473);
nand U18396 (N_18396,N_16827,N_16796);
or U18397 (N_18397,N_17359,N_17394);
nor U18398 (N_18398,N_16629,N_16478);
xor U18399 (N_18399,N_17381,N_17091);
or U18400 (N_18400,N_16865,N_16342);
xor U18401 (N_18401,N_16763,N_17091);
nor U18402 (N_18402,N_17432,N_17021);
and U18403 (N_18403,N_17231,N_16641);
and U18404 (N_18404,N_17189,N_16812);
nor U18405 (N_18405,N_17401,N_16603);
xor U18406 (N_18406,N_17256,N_17492);
nor U18407 (N_18407,N_16642,N_16538);
nand U18408 (N_18408,N_16970,N_17132);
nor U18409 (N_18409,N_17107,N_16276);
nor U18410 (N_18410,N_17189,N_16771);
xnor U18411 (N_18411,N_16323,N_16647);
xor U18412 (N_18412,N_17273,N_16254);
and U18413 (N_18413,N_17297,N_16324);
nor U18414 (N_18414,N_16679,N_16483);
nand U18415 (N_18415,N_17436,N_17040);
or U18416 (N_18416,N_16732,N_17086);
nand U18417 (N_18417,N_16467,N_16395);
nor U18418 (N_18418,N_16892,N_16829);
nand U18419 (N_18419,N_17376,N_17389);
and U18420 (N_18420,N_16653,N_16760);
and U18421 (N_18421,N_17129,N_17359);
xnor U18422 (N_18422,N_16842,N_16644);
nor U18423 (N_18423,N_16649,N_16315);
and U18424 (N_18424,N_17091,N_16954);
nor U18425 (N_18425,N_17191,N_16546);
xnor U18426 (N_18426,N_17364,N_17015);
nand U18427 (N_18427,N_17332,N_16859);
nor U18428 (N_18428,N_16476,N_17230);
nand U18429 (N_18429,N_17114,N_16665);
nor U18430 (N_18430,N_17234,N_16914);
xor U18431 (N_18431,N_16539,N_17120);
xor U18432 (N_18432,N_16738,N_16426);
xnor U18433 (N_18433,N_16509,N_17106);
or U18434 (N_18434,N_16418,N_17373);
nor U18435 (N_18435,N_17037,N_16736);
and U18436 (N_18436,N_17173,N_16912);
nand U18437 (N_18437,N_17420,N_17336);
nand U18438 (N_18438,N_16682,N_16432);
or U18439 (N_18439,N_16825,N_17324);
and U18440 (N_18440,N_16776,N_16818);
and U18441 (N_18441,N_17041,N_17017);
and U18442 (N_18442,N_16448,N_16534);
nand U18443 (N_18443,N_17376,N_17359);
nor U18444 (N_18444,N_16703,N_17085);
and U18445 (N_18445,N_16830,N_16414);
xnor U18446 (N_18446,N_17247,N_17087);
or U18447 (N_18447,N_16576,N_17073);
or U18448 (N_18448,N_16745,N_16845);
xor U18449 (N_18449,N_16513,N_16555);
nand U18450 (N_18450,N_16379,N_17279);
xnor U18451 (N_18451,N_16359,N_16468);
xor U18452 (N_18452,N_17134,N_17015);
nor U18453 (N_18453,N_16424,N_17011);
nand U18454 (N_18454,N_16299,N_17180);
or U18455 (N_18455,N_16919,N_16797);
nand U18456 (N_18456,N_17333,N_16624);
and U18457 (N_18457,N_16547,N_17262);
nand U18458 (N_18458,N_16564,N_16560);
and U18459 (N_18459,N_16485,N_16979);
and U18460 (N_18460,N_17461,N_17315);
nor U18461 (N_18461,N_17384,N_16950);
nand U18462 (N_18462,N_16959,N_17262);
nand U18463 (N_18463,N_16310,N_16505);
xnor U18464 (N_18464,N_16439,N_17390);
xnor U18465 (N_18465,N_16923,N_16311);
and U18466 (N_18466,N_17491,N_16897);
and U18467 (N_18467,N_16401,N_16502);
or U18468 (N_18468,N_16737,N_17130);
and U18469 (N_18469,N_16892,N_16415);
xor U18470 (N_18470,N_16738,N_16747);
nor U18471 (N_18471,N_17480,N_16626);
nor U18472 (N_18472,N_16458,N_17327);
xor U18473 (N_18473,N_16329,N_16728);
nand U18474 (N_18474,N_16785,N_16793);
or U18475 (N_18475,N_17161,N_16463);
nand U18476 (N_18476,N_17360,N_16500);
and U18477 (N_18477,N_16957,N_16502);
or U18478 (N_18478,N_17063,N_16506);
xor U18479 (N_18479,N_16966,N_16822);
nor U18480 (N_18480,N_16264,N_16950);
nor U18481 (N_18481,N_17272,N_17264);
and U18482 (N_18482,N_16966,N_17180);
or U18483 (N_18483,N_17312,N_16947);
nor U18484 (N_18484,N_16734,N_16630);
nand U18485 (N_18485,N_16991,N_16632);
nand U18486 (N_18486,N_16500,N_16751);
nor U18487 (N_18487,N_17054,N_16692);
nand U18488 (N_18488,N_16991,N_16370);
nor U18489 (N_18489,N_17147,N_17292);
nor U18490 (N_18490,N_17377,N_16978);
nor U18491 (N_18491,N_16395,N_16628);
and U18492 (N_18492,N_16470,N_16392);
nor U18493 (N_18493,N_16341,N_16725);
or U18494 (N_18494,N_16461,N_17028);
xor U18495 (N_18495,N_17024,N_17262);
and U18496 (N_18496,N_16475,N_17389);
nor U18497 (N_18497,N_16824,N_16837);
nand U18498 (N_18498,N_17155,N_17315);
xor U18499 (N_18499,N_16746,N_16897);
xor U18500 (N_18500,N_17004,N_16523);
xnor U18501 (N_18501,N_16738,N_16856);
nor U18502 (N_18502,N_16808,N_17129);
or U18503 (N_18503,N_17487,N_16839);
nor U18504 (N_18504,N_17433,N_17456);
nand U18505 (N_18505,N_17377,N_16554);
xnor U18506 (N_18506,N_16590,N_17246);
xor U18507 (N_18507,N_16756,N_17004);
nor U18508 (N_18508,N_16837,N_17114);
xnor U18509 (N_18509,N_16307,N_16530);
or U18510 (N_18510,N_17340,N_16396);
or U18511 (N_18511,N_17162,N_16845);
and U18512 (N_18512,N_17352,N_17227);
and U18513 (N_18513,N_16714,N_17219);
and U18514 (N_18514,N_17012,N_17425);
xnor U18515 (N_18515,N_16833,N_17374);
and U18516 (N_18516,N_16774,N_16420);
nand U18517 (N_18517,N_17255,N_16549);
or U18518 (N_18518,N_16989,N_16445);
xnor U18519 (N_18519,N_16557,N_16642);
or U18520 (N_18520,N_16808,N_16472);
nand U18521 (N_18521,N_16726,N_17300);
nand U18522 (N_18522,N_17200,N_17134);
or U18523 (N_18523,N_16934,N_17065);
or U18524 (N_18524,N_16883,N_17475);
nor U18525 (N_18525,N_16415,N_17096);
and U18526 (N_18526,N_16730,N_16750);
xor U18527 (N_18527,N_17138,N_16367);
nor U18528 (N_18528,N_16943,N_16944);
nor U18529 (N_18529,N_16339,N_17336);
nor U18530 (N_18530,N_17047,N_17364);
or U18531 (N_18531,N_17342,N_16810);
xor U18532 (N_18532,N_16644,N_17434);
and U18533 (N_18533,N_16596,N_17071);
nand U18534 (N_18534,N_17405,N_16454);
and U18535 (N_18535,N_16462,N_16460);
and U18536 (N_18536,N_16764,N_17488);
nor U18537 (N_18537,N_17357,N_17286);
or U18538 (N_18538,N_16760,N_16914);
nand U18539 (N_18539,N_16705,N_16577);
and U18540 (N_18540,N_16689,N_16561);
nand U18541 (N_18541,N_16298,N_17319);
and U18542 (N_18542,N_16255,N_17242);
xnor U18543 (N_18543,N_17475,N_17322);
xor U18544 (N_18544,N_16309,N_16549);
nand U18545 (N_18545,N_16731,N_16544);
nor U18546 (N_18546,N_16598,N_17169);
nor U18547 (N_18547,N_17285,N_16568);
and U18548 (N_18548,N_17275,N_16441);
xor U18549 (N_18549,N_16597,N_17112);
and U18550 (N_18550,N_16974,N_16923);
and U18551 (N_18551,N_16559,N_16871);
or U18552 (N_18552,N_16845,N_17266);
nor U18553 (N_18553,N_16826,N_16725);
or U18554 (N_18554,N_16824,N_16319);
nand U18555 (N_18555,N_16301,N_16730);
nor U18556 (N_18556,N_17278,N_16804);
xnor U18557 (N_18557,N_17416,N_16367);
or U18558 (N_18558,N_17277,N_17271);
and U18559 (N_18559,N_17427,N_16353);
or U18560 (N_18560,N_16513,N_17128);
xor U18561 (N_18561,N_17224,N_16586);
or U18562 (N_18562,N_17200,N_16556);
nor U18563 (N_18563,N_16641,N_16960);
nand U18564 (N_18564,N_17246,N_17307);
xnor U18565 (N_18565,N_16960,N_17195);
nand U18566 (N_18566,N_17370,N_16332);
nand U18567 (N_18567,N_17368,N_17162);
and U18568 (N_18568,N_16630,N_16890);
nand U18569 (N_18569,N_16662,N_17241);
or U18570 (N_18570,N_16259,N_16403);
or U18571 (N_18571,N_17329,N_16758);
and U18572 (N_18572,N_16869,N_17024);
or U18573 (N_18573,N_16670,N_17491);
or U18574 (N_18574,N_16918,N_16367);
and U18575 (N_18575,N_17180,N_16556);
nor U18576 (N_18576,N_17021,N_17213);
xnor U18577 (N_18577,N_17088,N_17045);
nand U18578 (N_18578,N_17186,N_17361);
nand U18579 (N_18579,N_16979,N_16703);
xnor U18580 (N_18580,N_16928,N_16429);
nor U18581 (N_18581,N_17285,N_16416);
nand U18582 (N_18582,N_17091,N_16799);
or U18583 (N_18583,N_16616,N_17352);
xor U18584 (N_18584,N_16980,N_17139);
nand U18585 (N_18585,N_17186,N_16279);
nand U18586 (N_18586,N_16507,N_16867);
and U18587 (N_18587,N_16428,N_16511);
and U18588 (N_18588,N_17305,N_16610);
and U18589 (N_18589,N_17102,N_16775);
xnor U18590 (N_18590,N_16287,N_16302);
and U18591 (N_18591,N_16536,N_16667);
or U18592 (N_18592,N_16731,N_16715);
xnor U18593 (N_18593,N_16992,N_16594);
nor U18594 (N_18594,N_16455,N_17155);
xor U18595 (N_18595,N_16337,N_17010);
nor U18596 (N_18596,N_17327,N_17469);
and U18597 (N_18597,N_16537,N_16932);
or U18598 (N_18598,N_16454,N_16767);
nand U18599 (N_18599,N_17443,N_17410);
nor U18600 (N_18600,N_16276,N_16662);
nor U18601 (N_18601,N_16694,N_16252);
and U18602 (N_18602,N_16283,N_16700);
nand U18603 (N_18603,N_17452,N_17121);
and U18604 (N_18604,N_16918,N_16942);
xor U18605 (N_18605,N_17185,N_16251);
nor U18606 (N_18606,N_16255,N_17207);
xor U18607 (N_18607,N_17016,N_16657);
nor U18608 (N_18608,N_16725,N_16485);
and U18609 (N_18609,N_16464,N_17166);
nor U18610 (N_18610,N_17093,N_16635);
nor U18611 (N_18611,N_17139,N_17037);
nand U18612 (N_18612,N_17346,N_16453);
xor U18613 (N_18613,N_16671,N_16832);
or U18614 (N_18614,N_16577,N_16943);
nor U18615 (N_18615,N_17178,N_16748);
xnor U18616 (N_18616,N_17449,N_17364);
and U18617 (N_18617,N_17416,N_17348);
xor U18618 (N_18618,N_17397,N_16514);
nand U18619 (N_18619,N_16674,N_16626);
and U18620 (N_18620,N_16287,N_17243);
nor U18621 (N_18621,N_17347,N_16385);
nor U18622 (N_18622,N_17318,N_17383);
nor U18623 (N_18623,N_16427,N_17267);
and U18624 (N_18624,N_16546,N_16459);
or U18625 (N_18625,N_16733,N_16757);
xor U18626 (N_18626,N_16987,N_16988);
or U18627 (N_18627,N_17366,N_16363);
xor U18628 (N_18628,N_17454,N_17292);
xor U18629 (N_18629,N_16421,N_16578);
xnor U18630 (N_18630,N_16762,N_16336);
or U18631 (N_18631,N_17321,N_16356);
nand U18632 (N_18632,N_17162,N_16326);
xnor U18633 (N_18633,N_16679,N_16550);
or U18634 (N_18634,N_17280,N_16549);
and U18635 (N_18635,N_17116,N_16569);
nand U18636 (N_18636,N_16928,N_17309);
nand U18637 (N_18637,N_16297,N_16620);
nor U18638 (N_18638,N_17210,N_17207);
nor U18639 (N_18639,N_16931,N_16541);
and U18640 (N_18640,N_16294,N_16852);
and U18641 (N_18641,N_16895,N_16390);
nor U18642 (N_18642,N_17410,N_17112);
and U18643 (N_18643,N_17077,N_16586);
or U18644 (N_18644,N_17223,N_16994);
nand U18645 (N_18645,N_16774,N_16372);
nor U18646 (N_18646,N_16603,N_16453);
or U18647 (N_18647,N_16832,N_17416);
nand U18648 (N_18648,N_17036,N_16330);
nand U18649 (N_18649,N_17263,N_17252);
nor U18650 (N_18650,N_16587,N_16652);
nor U18651 (N_18651,N_17232,N_17242);
xor U18652 (N_18652,N_16625,N_17292);
nor U18653 (N_18653,N_17254,N_17310);
xor U18654 (N_18654,N_16871,N_16562);
xor U18655 (N_18655,N_17020,N_17394);
xnor U18656 (N_18656,N_16933,N_16558);
and U18657 (N_18657,N_17257,N_17464);
and U18658 (N_18658,N_16552,N_16688);
and U18659 (N_18659,N_16551,N_16436);
xor U18660 (N_18660,N_16647,N_16264);
nand U18661 (N_18661,N_16938,N_17185);
nor U18662 (N_18662,N_17351,N_16868);
nor U18663 (N_18663,N_17170,N_17258);
nand U18664 (N_18664,N_17434,N_16392);
xnor U18665 (N_18665,N_17435,N_16711);
xor U18666 (N_18666,N_16673,N_17188);
xnor U18667 (N_18667,N_17404,N_16774);
nor U18668 (N_18668,N_16509,N_16831);
nor U18669 (N_18669,N_17337,N_17165);
and U18670 (N_18670,N_17221,N_16387);
xnor U18671 (N_18671,N_16657,N_17498);
or U18672 (N_18672,N_16748,N_17107);
xor U18673 (N_18673,N_16930,N_16873);
and U18674 (N_18674,N_17240,N_16418);
or U18675 (N_18675,N_16866,N_16808);
xnor U18676 (N_18676,N_16695,N_17077);
xor U18677 (N_18677,N_16567,N_16385);
nand U18678 (N_18678,N_17331,N_17155);
and U18679 (N_18679,N_16685,N_16462);
nor U18680 (N_18680,N_16372,N_16377);
and U18681 (N_18681,N_17095,N_17428);
nand U18682 (N_18682,N_16800,N_16541);
xor U18683 (N_18683,N_16410,N_16696);
xnor U18684 (N_18684,N_16947,N_17453);
or U18685 (N_18685,N_17335,N_17053);
xnor U18686 (N_18686,N_16699,N_17214);
nand U18687 (N_18687,N_16641,N_16793);
nand U18688 (N_18688,N_16476,N_17215);
nor U18689 (N_18689,N_16500,N_16814);
nor U18690 (N_18690,N_16856,N_16653);
nor U18691 (N_18691,N_16340,N_16798);
xnor U18692 (N_18692,N_16331,N_17435);
nor U18693 (N_18693,N_16334,N_16549);
and U18694 (N_18694,N_17114,N_17178);
and U18695 (N_18695,N_16764,N_17413);
xor U18696 (N_18696,N_17272,N_16764);
nor U18697 (N_18697,N_16436,N_16455);
xor U18698 (N_18698,N_16942,N_17302);
xor U18699 (N_18699,N_16739,N_16589);
nor U18700 (N_18700,N_16620,N_16734);
or U18701 (N_18701,N_16658,N_16406);
or U18702 (N_18702,N_16609,N_16640);
nor U18703 (N_18703,N_16592,N_17423);
or U18704 (N_18704,N_16482,N_16283);
nand U18705 (N_18705,N_16564,N_16660);
xnor U18706 (N_18706,N_16553,N_16637);
and U18707 (N_18707,N_16887,N_16885);
nand U18708 (N_18708,N_16911,N_16573);
nor U18709 (N_18709,N_17451,N_17159);
xnor U18710 (N_18710,N_16892,N_16476);
nand U18711 (N_18711,N_17325,N_16324);
and U18712 (N_18712,N_17212,N_17056);
xor U18713 (N_18713,N_16441,N_16571);
and U18714 (N_18714,N_16790,N_16536);
or U18715 (N_18715,N_16735,N_16473);
xor U18716 (N_18716,N_16917,N_17009);
or U18717 (N_18717,N_17147,N_16650);
and U18718 (N_18718,N_16698,N_16329);
and U18719 (N_18719,N_16934,N_17116);
xor U18720 (N_18720,N_17357,N_16579);
or U18721 (N_18721,N_17268,N_16931);
nor U18722 (N_18722,N_17217,N_17193);
and U18723 (N_18723,N_16411,N_17008);
and U18724 (N_18724,N_16499,N_17166);
and U18725 (N_18725,N_16509,N_16346);
xnor U18726 (N_18726,N_17181,N_16994);
nand U18727 (N_18727,N_16790,N_16794);
nand U18728 (N_18728,N_17456,N_17070);
xnor U18729 (N_18729,N_16602,N_17407);
nand U18730 (N_18730,N_17253,N_17293);
nor U18731 (N_18731,N_16541,N_16559);
nand U18732 (N_18732,N_17068,N_16342);
nand U18733 (N_18733,N_17253,N_16310);
nor U18734 (N_18734,N_17475,N_17016);
and U18735 (N_18735,N_17172,N_17049);
nand U18736 (N_18736,N_16515,N_16564);
xor U18737 (N_18737,N_16650,N_16437);
nor U18738 (N_18738,N_16564,N_16333);
nor U18739 (N_18739,N_16946,N_16909);
nor U18740 (N_18740,N_17229,N_16616);
nor U18741 (N_18741,N_17377,N_16530);
nor U18742 (N_18742,N_17395,N_16901);
nand U18743 (N_18743,N_16433,N_16269);
xnor U18744 (N_18744,N_16700,N_17048);
nor U18745 (N_18745,N_17185,N_17280);
xor U18746 (N_18746,N_17284,N_17055);
or U18747 (N_18747,N_17182,N_17153);
nor U18748 (N_18748,N_16906,N_16695);
nand U18749 (N_18749,N_16566,N_16805);
nor U18750 (N_18750,N_18371,N_18181);
xnor U18751 (N_18751,N_17850,N_17758);
nor U18752 (N_18752,N_18529,N_18676);
or U18753 (N_18753,N_17804,N_17774);
nor U18754 (N_18754,N_18111,N_18680);
nand U18755 (N_18755,N_18082,N_17766);
or U18756 (N_18756,N_17877,N_18241);
nor U18757 (N_18757,N_18234,N_17911);
and U18758 (N_18758,N_17579,N_18457);
xnor U18759 (N_18759,N_18744,N_18040);
and U18760 (N_18760,N_17888,N_18369);
nand U18761 (N_18761,N_17838,N_18413);
xnor U18762 (N_18762,N_17626,N_18123);
or U18763 (N_18763,N_18305,N_18162);
nor U18764 (N_18764,N_18533,N_18617);
nand U18765 (N_18765,N_18309,N_18386);
xor U18766 (N_18766,N_18404,N_18532);
xnor U18767 (N_18767,N_18577,N_18002);
nand U18768 (N_18768,N_18455,N_18745);
nand U18769 (N_18769,N_17999,N_17903);
and U18770 (N_18770,N_18128,N_18520);
and U18771 (N_18771,N_18535,N_18377);
nand U18772 (N_18772,N_18347,N_17519);
xor U18773 (N_18773,N_17778,N_18120);
nand U18774 (N_18774,N_17906,N_18094);
or U18775 (N_18775,N_17987,N_18236);
and U18776 (N_18776,N_17924,N_17973);
or U18777 (N_18777,N_17853,N_17709);
and U18778 (N_18778,N_17749,N_17539);
nor U18779 (N_18779,N_18585,N_17921);
nand U18780 (N_18780,N_17553,N_17633);
xor U18781 (N_18781,N_18013,N_18672);
or U18782 (N_18782,N_17568,N_17737);
xor U18783 (N_18783,N_18544,N_17677);
or U18784 (N_18784,N_18539,N_18280);
and U18785 (N_18785,N_18502,N_18050);
or U18786 (N_18786,N_18137,N_17615);
nand U18787 (N_18787,N_17963,N_17739);
nand U18788 (N_18788,N_17975,N_17538);
nand U18789 (N_18789,N_18285,N_17800);
xnor U18790 (N_18790,N_17544,N_17712);
xor U18791 (N_18791,N_18000,N_18126);
or U18792 (N_18792,N_18301,N_18109);
nor U18793 (N_18793,N_18553,N_17655);
nand U18794 (N_18794,N_18047,N_18452);
or U18795 (N_18795,N_17604,N_17708);
nand U18796 (N_18796,N_17979,N_17762);
nor U18797 (N_18797,N_18150,N_18392);
or U18798 (N_18798,N_18634,N_18567);
xor U18799 (N_18799,N_18068,N_18438);
nand U18800 (N_18800,N_17943,N_18558);
nand U18801 (N_18801,N_18546,N_18584);
or U18802 (N_18802,N_18025,N_18232);
or U18803 (N_18803,N_17754,N_18102);
nor U18804 (N_18804,N_18562,N_18433);
nand U18805 (N_18805,N_17535,N_18589);
and U18806 (N_18806,N_17831,N_18422);
xor U18807 (N_18807,N_18103,N_18063);
xnor U18808 (N_18808,N_18582,N_17680);
nor U18809 (N_18809,N_18435,N_18623);
and U18810 (N_18810,N_18415,N_18294);
xor U18811 (N_18811,N_17607,N_18208);
and U18812 (N_18812,N_18008,N_18210);
nand U18813 (N_18813,N_17893,N_18341);
and U18814 (N_18814,N_17522,N_18651);
nor U18815 (N_18815,N_18169,N_18700);
or U18816 (N_18816,N_18314,N_17767);
nand U18817 (N_18817,N_17736,N_17640);
nor U18818 (N_18818,N_18458,N_18159);
or U18819 (N_18819,N_17628,N_17833);
nand U18820 (N_18820,N_18317,N_17907);
nand U18821 (N_18821,N_18498,N_17944);
nand U18822 (N_18822,N_18657,N_18446);
nor U18823 (N_18823,N_18440,N_18054);
nor U18824 (N_18824,N_17554,N_17595);
nand U18825 (N_18825,N_17507,N_17878);
xor U18826 (N_18826,N_18555,N_17769);
and U18827 (N_18827,N_18110,N_18428);
or U18828 (N_18828,N_18659,N_17970);
and U18829 (N_18829,N_18340,N_17560);
and U18830 (N_18830,N_18607,N_18276);
nor U18831 (N_18831,N_18112,N_18543);
or U18832 (N_18832,N_18733,N_18015);
nand U18833 (N_18833,N_17997,N_18296);
or U18834 (N_18834,N_18702,N_17678);
or U18835 (N_18835,N_17891,N_17728);
and U18836 (N_18836,N_18175,N_17581);
xor U18837 (N_18837,N_18565,N_18603);
xor U18838 (N_18838,N_18564,N_17514);
nand U18839 (N_18839,N_18245,N_18287);
or U18840 (N_18840,N_18179,N_18005);
xor U18841 (N_18841,N_18174,N_17717);
or U18842 (N_18842,N_18714,N_17761);
and U18843 (N_18843,N_18077,N_18482);
nor U18844 (N_18844,N_17520,N_17613);
nor U18845 (N_18845,N_17741,N_18135);
and U18846 (N_18846,N_17948,N_17991);
nand U18847 (N_18847,N_18283,N_18673);
nand U18848 (N_18848,N_17793,N_18396);
or U18849 (N_18849,N_17646,N_18331);
and U18850 (N_18850,N_18719,N_17666);
nand U18851 (N_18851,N_18568,N_18662);
nand U18852 (N_18852,N_17618,N_18460);
or U18853 (N_18853,N_17842,N_18160);
xnor U18854 (N_18854,N_18715,N_18125);
nor U18855 (N_18855,N_18721,N_17720);
and U18856 (N_18856,N_17710,N_18749);
nor U18857 (N_18857,N_17608,N_18004);
or U18858 (N_18858,N_18027,N_18198);
or U18859 (N_18859,N_17593,N_17611);
nor U18860 (N_18860,N_18049,N_17691);
nor U18861 (N_18861,N_17781,N_17654);
xnor U18862 (N_18862,N_18207,N_18183);
xor U18863 (N_18863,N_17980,N_17798);
nor U18864 (N_18864,N_17589,N_17564);
nand U18865 (N_18865,N_18352,N_18081);
nor U18866 (N_18866,N_17860,N_17516);
nand U18867 (N_18867,N_18595,N_18664);
nor U18868 (N_18868,N_17662,N_17596);
and U18869 (N_18869,N_17733,N_18191);
xor U18870 (N_18870,N_17630,N_18221);
nand U18871 (N_18871,N_17658,N_17543);
nor U18872 (N_18872,N_18057,N_18261);
xnor U18873 (N_18873,N_17729,N_17967);
xor U18874 (N_18874,N_18140,N_18315);
or U18875 (N_18875,N_18594,N_18472);
xor U18876 (N_18876,N_18268,N_18747);
xnor U18877 (N_18877,N_18330,N_18693);
nor U18878 (N_18878,N_17650,N_17956);
nand U18879 (N_18879,N_18353,N_18566);
and U18880 (N_18880,N_18726,N_17609);
nand U18881 (N_18881,N_17964,N_18153);
or U18882 (N_18882,N_18441,N_18678);
or U18883 (N_18883,N_18333,N_18373);
and U18884 (N_18884,N_17847,N_17965);
xnor U18885 (N_18885,N_18053,N_17515);
and U18886 (N_18886,N_17526,N_17884);
and U18887 (N_18887,N_17835,N_18447);
and U18888 (N_18888,N_18591,N_18530);
and U18889 (N_18889,N_18439,N_18354);
xor U18890 (N_18890,N_18090,N_18394);
nand U18891 (N_18891,N_18319,N_18074);
xor U18892 (N_18892,N_17856,N_17585);
or U18893 (N_18893,N_17852,N_18148);
xnor U18894 (N_18894,N_18501,N_18638);
and U18895 (N_18895,N_17742,N_17692);
xnor U18896 (N_18896,N_18293,N_17636);
or U18897 (N_18897,N_17772,N_17527);
xor U18898 (N_18898,N_18092,N_18359);
or U18899 (N_18899,N_17916,N_17701);
nor U18900 (N_18900,N_18122,N_17575);
or U18901 (N_18901,N_17873,N_17722);
nand U18902 (N_18902,N_17969,N_18527);
nand U18903 (N_18903,N_18574,N_18610);
xor U18904 (N_18904,N_18172,N_18224);
or U18905 (N_18905,N_17718,N_18199);
or U18906 (N_18906,N_18557,N_18635);
nor U18907 (N_18907,N_17922,N_18030);
or U18908 (N_18908,N_18476,N_18096);
xnor U18909 (N_18909,N_18531,N_18541);
or U18910 (N_18910,N_18604,N_18216);
or U18911 (N_18911,N_18615,N_18576);
and U18912 (N_18912,N_17610,N_18338);
xor U18913 (N_18913,N_18098,N_18249);
and U18914 (N_18914,N_17686,N_18445);
and U18915 (N_18915,N_17962,N_18526);
nand U18916 (N_18916,N_18692,N_17752);
nand U18917 (N_18917,N_17525,N_17819);
or U18918 (N_18918,N_18034,N_17945);
and U18919 (N_18919,N_18259,N_18419);
or U18920 (N_18920,N_18266,N_17971);
and U18921 (N_18921,N_18704,N_18718);
nor U18922 (N_18922,N_17745,N_17669);
nand U18923 (N_18923,N_18402,N_18243);
xor U18924 (N_18924,N_18303,N_18361);
or U18925 (N_18925,N_17644,N_18357);
nor U18926 (N_18926,N_18376,N_18084);
nand U18927 (N_18927,N_18011,N_17990);
xnor U18928 (N_18928,N_17756,N_17574);
nor U18929 (N_18929,N_18345,N_18290);
nor U18930 (N_18930,N_18573,N_17801);
nand U18931 (N_18931,N_17513,N_17875);
nand U18932 (N_18932,N_18432,N_18674);
nand U18933 (N_18933,N_17989,N_17668);
or U18934 (N_18934,N_17941,N_18206);
nor U18935 (N_18935,N_18586,N_18026);
or U18936 (N_18936,N_18253,N_17889);
xnor U18937 (N_18937,N_17755,N_17620);
nor U18938 (N_18938,N_17510,N_17587);
and U18939 (N_18939,N_18188,N_17530);
or U18940 (N_18940,N_18348,N_18713);
or U18941 (N_18941,N_17748,N_18235);
xnor U18942 (N_18942,N_18547,N_18080);
nand U18943 (N_18943,N_18503,N_18258);
xor U18944 (N_18944,N_17857,N_18709);
xor U18945 (N_18945,N_17809,N_17919);
nor U18946 (N_18946,N_18580,N_18267);
xor U18947 (N_18947,N_17682,N_17994);
or U18948 (N_18948,N_18017,N_18456);
or U18949 (N_18949,N_18156,N_18654);
xor U18950 (N_18950,N_18029,N_17839);
or U18951 (N_18951,N_18540,N_17714);
and U18952 (N_18952,N_18480,N_18180);
xor U18953 (N_18953,N_17823,N_18740);
nor U18954 (N_18954,N_18563,N_18406);
xnor U18955 (N_18955,N_17663,N_17699);
xor U18956 (N_18956,N_18263,N_18114);
or U18957 (N_18957,N_17643,N_18738);
xor U18958 (N_18958,N_18523,N_18675);
or U18959 (N_18959,N_18323,N_18417);
or U18960 (N_18960,N_18147,N_18625);
or U18961 (N_18961,N_18048,N_18493);
and U18962 (N_18962,N_18157,N_18661);
and U18963 (N_18963,N_17672,N_17836);
xor U18964 (N_18964,N_17910,N_18132);
xnor U18965 (N_18965,N_18142,N_18233);
and U18966 (N_18966,N_18667,N_18411);
or U18967 (N_18967,N_18736,N_17719);
nand U18968 (N_18968,N_17625,N_18064);
and U18969 (N_18969,N_18105,N_17641);
nor U18970 (N_18970,N_18583,N_17946);
nor U18971 (N_18971,N_17558,N_17993);
nor U18972 (N_18972,N_18601,N_18737);
xor U18973 (N_18973,N_17547,N_17652);
xor U18974 (N_18974,N_18384,N_18600);
xor U18975 (N_18975,N_17784,N_18485);
xnor U18976 (N_18976,N_18450,N_17874);
xnor U18977 (N_18977,N_18743,N_18278);
or U18978 (N_18978,N_18219,N_17542);
nand U18979 (N_18979,N_18036,N_18133);
nand U18980 (N_18980,N_17932,N_18292);
and U18981 (N_18981,N_18382,N_17501);
nand U18982 (N_18982,N_17619,N_17811);
nor U18983 (N_18983,N_17697,N_17787);
or U18984 (N_18984,N_18538,N_17586);
and U18985 (N_18985,N_17828,N_18732);
and U18986 (N_18986,N_18307,N_17511);
or U18987 (N_18987,N_18100,N_18459);
and U18988 (N_18988,N_18149,N_18506);
xor U18989 (N_18989,N_18682,N_18729);
or U18990 (N_18990,N_18009,N_18071);
xor U18991 (N_18991,N_17707,N_18522);
and U18992 (N_18992,N_18627,N_18592);
xor U18993 (N_18993,N_18525,N_17978);
xor U18994 (N_18994,N_17660,N_17689);
nand U18995 (N_18995,N_18061,N_17930);
nor U18996 (N_18996,N_18468,N_18284);
and U18997 (N_18997,N_18368,N_18274);
xnor U18998 (N_18998,N_18426,N_17806);
nand U18999 (N_18999,N_18407,N_18537);
or U19000 (N_19000,N_18487,N_18521);
nor U19001 (N_19001,N_17812,N_18010);
or U19002 (N_19002,N_17934,N_17768);
and U19003 (N_19003,N_18681,N_18240);
nor U19004 (N_19004,N_17822,N_17982);
nor U19005 (N_19005,N_18237,N_17940);
or U19006 (N_19006,N_18614,N_18322);
nand U19007 (N_19007,N_18730,N_17909);
xor U19008 (N_19008,N_18524,N_18632);
nor U19009 (N_19009,N_17902,N_18701);
or U19010 (N_19010,N_17505,N_18182);
and U19011 (N_19011,N_17548,N_18746);
xor U19012 (N_19012,N_18028,N_17841);
nor U19013 (N_19013,N_18690,N_18629);
or U19014 (N_19014,N_17995,N_18511);
nand U19015 (N_19015,N_18488,N_18691);
or U19016 (N_19016,N_18257,N_18155);
or U19017 (N_19017,N_17675,N_18007);
nor U19018 (N_19018,N_17939,N_18479);
or U19019 (N_19019,N_17687,N_17676);
nand U19020 (N_19020,N_18337,N_18467);
or U19021 (N_19021,N_17876,N_18619);
and U19022 (N_19022,N_18260,N_17786);
or U19023 (N_19023,N_18003,N_17763);
xor U19024 (N_19024,N_17639,N_18121);
nand U19025 (N_19025,N_17753,N_18118);
nor U19026 (N_19026,N_18115,N_18051);
nand U19027 (N_19027,N_17740,N_18660);
xnor U19028 (N_19028,N_18019,N_18645);
nor U19029 (N_19029,N_18624,N_18088);
nand U19030 (N_19030,N_17817,N_18067);
xnor U19031 (N_19031,N_18325,N_18650);
or U19032 (N_19032,N_17540,N_18431);
or U19033 (N_19033,N_18470,N_18728);
or U19034 (N_19034,N_17868,N_18255);
nor U19035 (N_19035,N_17904,N_18443);
xnor U19036 (N_19036,N_18089,N_18575);
nand U19037 (N_19037,N_17532,N_17900);
or U19038 (N_19038,N_18289,N_18412);
xor U19039 (N_19039,N_17698,N_18041);
xnor U19040 (N_19040,N_18152,N_18213);
nand U19041 (N_19041,N_18324,N_17827);
xnor U19042 (N_19042,N_18087,N_18205);
xor U19043 (N_19043,N_18306,N_18463);
xnor U19044 (N_19044,N_18381,N_18262);
nand U19045 (N_19045,N_18666,N_17704);
xnor U19046 (N_19046,N_18039,N_17670);
and U19047 (N_19047,N_18668,N_18131);
nor U19048 (N_19048,N_18072,N_18058);
and U19049 (N_19049,N_17623,N_18549);
or U19050 (N_19050,N_17821,N_18542);
xor U19051 (N_19051,N_18490,N_17632);
nand U19052 (N_19052,N_17938,N_18193);
or U19053 (N_19053,N_18297,N_18197);
nand U19054 (N_19054,N_18722,N_17782);
xor U19055 (N_19055,N_17915,N_18395);
xor U19056 (N_19056,N_17914,N_18190);
nor U19057 (N_19057,N_17743,N_18326);
nor U19058 (N_19058,N_18454,N_18648);
and U19059 (N_19059,N_17832,N_17961);
nor U19060 (N_19060,N_17802,N_17614);
nand U19061 (N_19061,N_18229,N_18509);
nor U19062 (N_19062,N_17509,N_18708);
nand U19063 (N_19063,N_18579,N_18251);
nor U19064 (N_19064,N_18355,N_18069);
nand U19065 (N_19065,N_17984,N_18161);
or U19066 (N_19066,N_18697,N_18494);
or U19067 (N_19067,N_17949,N_18299);
nor U19068 (N_19068,N_17584,N_18343);
or U19069 (N_19069,N_18683,N_17805);
nor U19070 (N_19070,N_17985,N_17826);
nand U19071 (N_19071,N_17703,N_18598);
nand U19072 (N_19072,N_18066,N_17788);
or U19073 (N_19073,N_18688,N_17777);
nand U19074 (N_19074,N_17534,N_18185);
xor U19075 (N_19075,N_17917,N_17751);
and U19076 (N_19076,N_18165,N_18639);
nand U19077 (N_19077,N_18095,N_18130);
xnor U19078 (N_19078,N_17559,N_18416);
and U19079 (N_19079,N_18223,N_18390);
nand U19080 (N_19080,N_17523,N_17541);
and U19081 (N_19081,N_18741,N_18209);
or U19082 (N_19082,N_17923,N_17713);
xnor U19083 (N_19083,N_17517,N_17913);
nand U19084 (N_19084,N_17638,N_18196);
nand U19085 (N_19085,N_17550,N_18351);
nand U19086 (N_19086,N_18663,N_18497);
xor U19087 (N_19087,N_17594,N_18164);
or U19088 (N_19088,N_18134,N_17667);
xor U19089 (N_19089,N_18214,N_18158);
nor U19090 (N_19090,N_18246,N_18748);
nand U19091 (N_19091,N_17649,N_18486);
or U19092 (N_19092,N_18500,N_18363);
or U19093 (N_19093,N_18141,N_18146);
xnor U19094 (N_19094,N_17879,N_18033);
or U19095 (N_19095,N_17702,N_18403);
xnor U19096 (N_19096,N_17671,N_18554);
nand U19097 (N_19097,N_18641,N_17545);
nand U19098 (N_19098,N_17816,N_18366);
nor U19099 (N_19099,N_18630,N_18295);
or U19100 (N_19100,N_17750,N_17854);
nor U19101 (N_19101,N_17780,N_17790);
or U19102 (N_19102,N_17573,N_17651);
nor U19103 (N_19103,N_18018,N_18187);
nor U19104 (N_19104,N_17512,N_17706);
and U19105 (N_19105,N_17871,N_18186);
nand U19106 (N_19106,N_18194,N_18099);
nor U19107 (N_19107,N_18649,N_18587);
and U19108 (N_19108,N_18383,N_17583);
or U19109 (N_19109,N_17605,N_18313);
nand U19110 (N_19110,N_18101,N_18717);
nor U19111 (N_19111,N_18515,N_17795);
xor U19112 (N_19112,N_18024,N_17881);
and U19113 (N_19113,N_18212,N_17773);
or U19114 (N_19114,N_18372,N_17617);
and U19115 (N_19115,N_18388,N_17746);
nand U19116 (N_19116,N_18083,N_17657);
xor U19117 (N_19117,N_17684,N_18242);
nor U19118 (N_19118,N_18093,N_17601);
and U19119 (N_19119,N_18512,N_18465);
xnor U19120 (N_19120,N_18442,N_17616);
nand U19121 (N_19121,N_18510,N_18362);
nor U19122 (N_19122,N_17928,N_18477);
nand U19123 (N_19123,N_17679,N_18473);
nor U19124 (N_19124,N_18065,N_17950);
and U19125 (N_19125,N_17771,N_18217);
nor U19126 (N_19126,N_18086,N_18677);
and U19127 (N_19127,N_17834,N_17591);
nor U19128 (N_19128,N_17716,N_17775);
nor U19129 (N_19129,N_17927,N_18550);
nor U19130 (N_19130,N_17977,N_18508);
nor U19131 (N_19131,N_17642,N_17966);
or U19132 (N_19132,N_18076,N_18012);
nor U19133 (N_19133,N_17843,N_17936);
or U19134 (N_19134,N_18492,N_18184);
or U19135 (N_19135,N_17974,N_17606);
nor U19136 (N_19136,N_18312,N_17959);
nor U19137 (N_19137,N_17556,N_17688);
nor U19138 (N_19138,N_18646,N_18572);
xnor U19139 (N_19139,N_18356,N_17631);
xor U19140 (N_19140,N_18052,N_18723);
nor U19141 (N_19141,N_18517,N_18379);
nor U19142 (N_19142,N_18669,N_17863);
nor U19143 (N_19143,N_18484,N_18321);
or U19144 (N_19144,N_17957,N_18483);
xnor U19145 (N_19145,N_18265,N_18489);
nor U19146 (N_19146,N_17549,N_17905);
nand U19147 (N_19147,N_18588,N_17551);
xnor U19148 (N_19148,N_17955,N_17598);
and U19149 (N_19149,N_18350,N_17635);
xnor U19150 (N_19150,N_18329,N_17960);
xnor U19151 (N_19151,N_17685,N_18720);
xnor U19152 (N_19152,N_18006,N_18399);
xnor U19153 (N_19153,N_18023,N_17624);
nor U19154 (N_19154,N_18405,N_17599);
and U19155 (N_19155,N_17552,N_17791);
and U19156 (N_19156,N_18695,N_18075);
and U19157 (N_19157,N_18124,N_17637);
nand U19158 (N_19158,N_17858,N_18385);
xnor U19159 (N_19159,N_17731,N_18374);
or U19160 (N_19160,N_18593,N_17747);
nand U19161 (N_19161,N_17942,N_17757);
nor U19162 (N_19162,N_17518,N_17502);
or U19163 (N_19163,N_18079,N_17629);
nor U19164 (N_19164,N_18464,N_17500);
xnor U19165 (N_19165,N_18665,N_18408);
nand U19166 (N_19166,N_17715,N_18536);
nor U19167 (N_19167,N_17653,N_17765);
nor U19168 (N_19168,N_18252,N_18073);
or U19169 (N_19169,N_18401,N_18300);
xor U19170 (N_19170,N_17813,N_17845);
xnor U19171 (N_19171,N_17603,N_18308);
nand U19172 (N_19172,N_18062,N_18344);
xnor U19173 (N_19173,N_17890,N_17810);
or U19174 (N_19174,N_17645,N_17602);
or U19175 (N_19175,N_18696,N_18171);
xnor U19176 (N_19176,N_18277,N_18706);
and U19177 (N_19177,N_18104,N_17918);
and U19178 (N_19178,N_18398,N_18166);
or U19179 (N_19179,N_18612,N_17711);
nor U19180 (N_19180,N_18742,N_17700);
and U19181 (N_19181,N_17859,N_18670);
nor U19182 (N_19182,N_17565,N_17759);
nor U19183 (N_19183,N_18106,N_18545);
nand U19184 (N_19184,N_17531,N_17861);
nand U19185 (N_19185,N_18569,N_17869);
and U19186 (N_19186,N_18616,N_17794);
nor U19187 (N_19187,N_18671,N_17844);
and U19188 (N_19188,N_18712,N_18491);
nand U19189 (N_19189,N_18602,N_18304);
and U19190 (N_19190,N_17908,N_18302);
or U19191 (N_19191,N_17647,N_17533);
or U19192 (N_19192,N_18248,N_17572);
and U19193 (N_19193,N_18282,N_18453);
nand U19194 (N_19194,N_18250,N_18378);
nand U19195 (N_19195,N_18656,N_17735);
xnor U19196 (N_19196,N_17952,N_18551);
and U19197 (N_19197,N_18581,N_18621);
or U19198 (N_19198,N_17931,N_17954);
nand U19199 (N_19199,N_18727,N_17656);
xor U19200 (N_19200,N_18393,N_18225);
and U19201 (N_19201,N_18734,N_18699);
nand U19202 (N_19202,N_17665,N_18275);
nor U19203 (N_19203,N_18561,N_18475);
and U19204 (N_19204,N_18620,N_18514);
nor U19205 (N_19205,N_17933,N_17588);
nor U19206 (N_19206,N_18505,N_17725);
xnor U19207 (N_19207,N_18035,N_17892);
nor U19208 (N_19208,N_18410,N_18679);
xnor U19209 (N_19209,N_18154,N_18178);
xor U19210 (N_19210,N_18643,N_17726);
nor U19211 (N_19211,N_18332,N_18310);
nor U19212 (N_19212,N_18631,N_17988);
nor U19213 (N_19213,N_18270,N_17567);
nand U19214 (N_19214,N_18320,N_17947);
xor U19215 (N_19215,N_18045,N_17557);
nor U19216 (N_19216,N_17705,N_18144);
and U19217 (N_19217,N_18710,N_18238);
or U19218 (N_19218,N_18163,N_17571);
or U19219 (N_19219,N_18151,N_17661);
nor U19220 (N_19220,N_18247,N_18244);
or U19221 (N_19221,N_18055,N_18516);
nor U19222 (N_19222,N_17935,N_18342);
xnor U19223 (N_19223,N_18380,N_17951);
xor U19224 (N_19224,N_18552,N_17524);
nor U19225 (N_19225,N_18264,N_18097);
and U19226 (N_19226,N_18070,N_17724);
or U19227 (N_19227,N_18220,N_18414);
or U19228 (N_19228,N_18471,N_18195);
and U19229 (N_19229,N_18478,N_18496);
and U19230 (N_19230,N_18481,N_18420);
or U19231 (N_19231,N_17829,N_18031);
nand U19232 (N_19232,N_17760,N_18685);
xnor U19233 (N_19233,N_18316,N_17885);
or U19234 (N_19234,N_18429,N_18469);
nand U19235 (N_19235,N_17894,N_18436);
or U19236 (N_19236,N_18085,N_18548);
and U19237 (N_19237,N_18637,N_17506);
nand U19238 (N_19238,N_18400,N_18606);
and U19239 (N_19239,N_17880,N_18613);
nand U19240 (N_19240,N_18391,N_17764);
nand U19241 (N_19241,N_18640,N_18571);
xnor U19242 (N_19242,N_18626,N_18716);
and U19243 (N_19243,N_18168,N_17776);
or U19244 (N_19244,N_18117,N_18360);
xor U19245 (N_19245,N_18628,N_17566);
xnor U19246 (N_19246,N_18427,N_17681);
nor U19247 (N_19247,N_18618,N_17992);
or U19248 (N_19248,N_18387,N_18698);
nor U19249 (N_19249,N_18042,N_17851);
nor U19250 (N_19250,N_18037,N_18288);
or U19251 (N_19251,N_17503,N_18281);
xor U19252 (N_19252,N_18655,N_18254);
or U19253 (N_19253,N_18684,N_17899);
or U19254 (N_19254,N_18021,N_17848);
and U19255 (N_19255,N_18642,N_17830);
and U19256 (N_19256,N_18731,N_17958);
nor U19257 (N_19257,N_17744,N_18466);
nand U19258 (N_19258,N_17521,N_18652);
nor U19259 (N_19259,N_17528,N_17926);
or U19260 (N_19260,N_18364,N_17895);
nand U19261 (N_19261,N_17937,N_18725);
or U19262 (N_19262,N_18328,N_17862);
and U19263 (N_19263,N_18513,N_18059);
xnor U19264 (N_19264,N_18273,N_18611);
or U19265 (N_19265,N_17577,N_18534);
or U19266 (N_19266,N_18444,N_17693);
xor U19267 (N_19267,N_18409,N_17820);
and U19268 (N_19268,N_18686,N_17870);
xor U19269 (N_19269,N_18291,N_17855);
and U19270 (N_19270,N_18177,N_18001);
nand U19271 (N_19271,N_18375,N_18108);
nor U19272 (N_19272,N_18346,N_18056);
or U19273 (N_19273,N_17799,N_18334);
nor U19274 (N_19274,N_18425,N_18022);
and U19275 (N_19275,N_17897,N_17779);
xnor U19276 (N_19276,N_17696,N_17621);
xor U19277 (N_19277,N_18143,N_18694);
or U19278 (N_19278,N_18016,N_18707);
and U19279 (N_19279,N_17886,N_18578);
nand U19280 (N_19280,N_17986,N_17840);
nand U19281 (N_19281,N_18724,N_17582);
and U19282 (N_19282,N_18107,N_17953);
or U19283 (N_19283,N_18230,N_17818);
nor U19284 (N_19284,N_18367,N_17690);
and U19285 (N_19285,N_17674,N_18226);
nor U19286 (N_19286,N_18349,N_18129);
nor U19287 (N_19287,N_17546,N_17570);
xor U19288 (N_19288,N_18462,N_17770);
xnor U19289 (N_19289,N_17529,N_17864);
nor U19290 (N_19290,N_18271,N_17612);
and U19291 (N_19291,N_17673,N_18636);
xor U19292 (N_19292,N_18269,N_18437);
xnor U19293 (N_19293,N_17983,N_18227);
and U19294 (N_19294,N_17694,N_17837);
and U19295 (N_19295,N_17783,N_17732);
and U19296 (N_19296,N_17814,N_18078);
nor U19297 (N_19297,N_17508,N_17600);
nor U19298 (N_19298,N_18327,N_18590);
nand U19299 (N_19299,N_18318,N_18136);
nand U19300 (N_19300,N_18647,N_18622);
or U19301 (N_19301,N_18658,N_18139);
nand U19302 (N_19302,N_17622,N_18644);
xor U19303 (N_19303,N_18507,N_17883);
nor U19304 (N_19304,N_17627,N_18504);
and U19305 (N_19305,N_18609,N_17866);
and U19306 (N_19306,N_17563,N_18286);
nor U19307 (N_19307,N_17562,N_17882);
nand U19308 (N_19308,N_17659,N_18201);
nand U19309 (N_19309,N_18218,N_17561);
nor U19310 (N_19310,N_18597,N_18167);
or U19311 (N_19311,N_18599,N_17976);
xor U19312 (N_19312,N_17825,N_18204);
and U19313 (N_19313,N_17634,N_17865);
nor U19314 (N_19314,N_17597,N_18298);
nand U19315 (N_19315,N_18256,N_17846);
and U19316 (N_19316,N_17785,N_18605);
xnor U19317 (N_19317,N_17555,N_18397);
nand U19318 (N_19318,N_18339,N_18202);
and U19319 (N_19319,N_18272,N_18560);
xnor U19320 (N_19320,N_17727,N_17648);
or U19321 (N_19321,N_18044,N_17996);
or U19322 (N_19322,N_18633,N_18418);
nor U19323 (N_19323,N_18711,N_18739);
nand U19324 (N_19324,N_17590,N_18528);
nand U19325 (N_19325,N_18358,N_17807);
nor U19326 (N_19326,N_18365,N_18311);
nand U19327 (N_19327,N_18703,N_18145);
xnor U19328 (N_19328,N_18231,N_18389);
nor U19329 (N_19329,N_18173,N_18735);
or U19330 (N_19330,N_18138,N_18474);
or U19331 (N_19331,N_17808,N_17664);
and U19332 (N_19332,N_18518,N_17981);
nor U19333 (N_19333,N_18608,N_17504);
xor U19334 (N_19334,N_18043,N_18215);
nor U19335 (N_19335,N_18239,N_17925);
nand U19336 (N_19336,N_18434,N_17872);
nand U19337 (N_19337,N_18370,N_18421);
nand U19338 (N_19338,N_18192,N_17920);
xnor U19339 (N_19339,N_18200,N_17695);
nand U19340 (N_19340,N_18449,N_18559);
xnor U19341 (N_19341,N_18335,N_17968);
nor U19342 (N_19342,N_17569,N_18570);
or U19343 (N_19343,N_17815,N_18116);
and U19344 (N_19344,N_17578,N_17683);
nor U19345 (N_19345,N_17537,N_17896);
and U19346 (N_19346,N_17723,N_17738);
and U19347 (N_19347,N_18046,N_17592);
and U19348 (N_19348,N_18461,N_17576);
nor U19349 (N_19349,N_17887,N_17792);
nor U19350 (N_19350,N_18653,N_17898);
and U19351 (N_19351,N_18091,N_18424);
or U19352 (N_19352,N_18170,N_18689);
or U19353 (N_19353,N_18336,N_17580);
or U19354 (N_19354,N_17797,N_18430);
or U19355 (N_19355,N_18687,N_17867);
xnor U19356 (N_19356,N_18222,N_18451);
and U19357 (N_19357,N_18705,N_17789);
nand U19358 (N_19358,N_17734,N_17972);
xor U19359 (N_19359,N_17929,N_17803);
nor U19360 (N_19360,N_18038,N_18032);
or U19361 (N_19361,N_18495,N_17849);
and U19362 (N_19362,N_18014,N_18127);
or U19363 (N_19363,N_17730,N_18423);
nor U19364 (N_19364,N_18203,N_18211);
and U19365 (N_19365,N_18176,N_18448);
or U19366 (N_19366,N_17796,N_18519);
nand U19367 (N_19367,N_17721,N_18228);
xor U19368 (N_19368,N_18596,N_18020);
nand U19369 (N_19369,N_17536,N_18113);
or U19370 (N_19370,N_18499,N_17998);
or U19371 (N_19371,N_17901,N_18556);
xnor U19372 (N_19372,N_18279,N_18060);
or U19373 (N_19373,N_18119,N_17912);
nand U19374 (N_19374,N_17824,N_18189);
and U19375 (N_19375,N_18189,N_17537);
and U19376 (N_19376,N_18387,N_17793);
or U19377 (N_19377,N_18050,N_18398);
or U19378 (N_19378,N_18097,N_17864);
xor U19379 (N_19379,N_18293,N_18532);
nand U19380 (N_19380,N_18200,N_17886);
nand U19381 (N_19381,N_17675,N_18661);
or U19382 (N_19382,N_17739,N_17980);
nor U19383 (N_19383,N_18732,N_18406);
nor U19384 (N_19384,N_18005,N_17654);
or U19385 (N_19385,N_17999,N_17653);
xnor U19386 (N_19386,N_18165,N_18026);
nor U19387 (N_19387,N_17701,N_18605);
and U19388 (N_19388,N_17614,N_17724);
and U19389 (N_19389,N_18285,N_17801);
or U19390 (N_19390,N_18145,N_18542);
and U19391 (N_19391,N_17876,N_18467);
nand U19392 (N_19392,N_18508,N_18449);
or U19393 (N_19393,N_17503,N_18613);
xnor U19394 (N_19394,N_18467,N_18291);
or U19395 (N_19395,N_18448,N_18152);
nor U19396 (N_19396,N_18577,N_17605);
xnor U19397 (N_19397,N_17851,N_18703);
xnor U19398 (N_19398,N_18053,N_18605);
and U19399 (N_19399,N_18394,N_18461);
and U19400 (N_19400,N_18254,N_18743);
and U19401 (N_19401,N_18375,N_18512);
or U19402 (N_19402,N_18737,N_18203);
or U19403 (N_19403,N_18422,N_17880);
and U19404 (N_19404,N_18212,N_17590);
nor U19405 (N_19405,N_18675,N_18502);
and U19406 (N_19406,N_18525,N_18701);
nand U19407 (N_19407,N_18223,N_18269);
nand U19408 (N_19408,N_18179,N_17841);
xor U19409 (N_19409,N_18292,N_18136);
xnor U19410 (N_19410,N_18007,N_17866);
or U19411 (N_19411,N_18205,N_17772);
nor U19412 (N_19412,N_18088,N_17792);
and U19413 (N_19413,N_17624,N_18273);
and U19414 (N_19414,N_18514,N_17516);
nand U19415 (N_19415,N_18442,N_18007);
xor U19416 (N_19416,N_18133,N_18249);
and U19417 (N_19417,N_18600,N_18028);
and U19418 (N_19418,N_18329,N_18426);
nand U19419 (N_19419,N_18396,N_18162);
xnor U19420 (N_19420,N_18415,N_18489);
or U19421 (N_19421,N_18148,N_18094);
xor U19422 (N_19422,N_17814,N_18478);
or U19423 (N_19423,N_18462,N_17945);
or U19424 (N_19424,N_18088,N_17899);
or U19425 (N_19425,N_18098,N_18602);
or U19426 (N_19426,N_18193,N_18234);
nor U19427 (N_19427,N_18433,N_18496);
xnor U19428 (N_19428,N_17839,N_18695);
nor U19429 (N_19429,N_18020,N_18702);
or U19430 (N_19430,N_17941,N_18049);
xnor U19431 (N_19431,N_18231,N_17791);
nor U19432 (N_19432,N_17604,N_18142);
nor U19433 (N_19433,N_18281,N_18178);
or U19434 (N_19434,N_17691,N_18603);
nor U19435 (N_19435,N_17795,N_18176);
or U19436 (N_19436,N_18359,N_18685);
or U19437 (N_19437,N_18356,N_17739);
and U19438 (N_19438,N_17847,N_17956);
nor U19439 (N_19439,N_17818,N_17514);
nor U19440 (N_19440,N_18233,N_18631);
xor U19441 (N_19441,N_18613,N_18259);
xnor U19442 (N_19442,N_18479,N_18290);
xor U19443 (N_19443,N_18378,N_18230);
nor U19444 (N_19444,N_18588,N_18168);
or U19445 (N_19445,N_18200,N_18273);
nor U19446 (N_19446,N_18591,N_17540);
and U19447 (N_19447,N_18609,N_17632);
nand U19448 (N_19448,N_18193,N_18633);
or U19449 (N_19449,N_17577,N_18642);
nand U19450 (N_19450,N_17645,N_18501);
and U19451 (N_19451,N_18464,N_17616);
or U19452 (N_19452,N_17951,N_17854);
nand U19453 (N_19453,N_17914,N_17571);
nand U19454 (N_19454,N_17528,N_18177);
and U19455 (N_19455,N_18071,N_17770);
and U19456 (N_19456,N_18739,N_18040);
or U19457 (N_19457,N_18699,N_17663);
nand U19458 (N_19458,N_17579,N_17621);
or U19459 (N_19459,N_18270,N_18118);
nor U19460 (N_19460,N_18187,N_18722);
and U19461 (N_19461,N_18645,N_18414);
xnor U19462 (N_19462,N_17820,N_18652);
or U19463 (N_19463,N_18302,N_18158);
xor U19464 (N_19464,N_18662,N_18607);
nor U19465 (N_19465,N_17908,N_18174);
xor U19466 (N_19466,N_18553,N_17598);
nor U19467 (N_19467,N_18736,N_17765);
nand U19468 (N_19468,N_17899,N_17708);
and U19469 (N_19469,N_18359,N_18666);
nand U19470 (N_19470,N_17924,N_18202);
xor U19471 (N_19471,N_17783,N_17965);
and U19472 (N_19472,N_18657,N_17932);
nor U19473 (N_19473,N_18507,N_18304);
or U19474 (N_19474,N_17630,N_18723);
nor U19475 (N_19475,N_18174,N_17779);
nor U19476 (N_19476,N_17627,N_18306);
xnor U19477 (N_19477,N_17613,N_17957);
or U19478 (N_19478,N_17549,N_18484);
and U19479 (N_19479,N_18441,N_18394);
nand U19480 (N_19480,N_17860,N_18069);
or U19481 (N_19481,N_18708,N_18202);
nand U19482 (N_19482,N_17779,N_18699);
nor U19483 (N_19483,N_18722,N_18196);
and U19484 (N_19484,N_18411,N_18198);
xnor U19485 (N_19485,N_18065,N_17622);
and U19486 (N_19486,N_17549,N_17872);
nor U19487 (N_19487,N_17777,N_17766);
nor U19488 (N_19488,N_17714,N_17629);
and U19489 (N_19489,N_18051,N_17989);
xor U19490 (N_19490,N_18397,N_18712);
xor U19491 (N_19491,N_18688,N_18471);
and U19492 (N_19492,N_18264,N_18045);
nand U19493 (N_19493,N_17896,N_18424);
xor U19494 (N_19494,N_18034,N_18138);
xor U19495 (N_19495,N_18165,N_18305);
and U19496 (N_19496,N_17524,N_17861);
nor U19497 (N_19497,N_18391,N_18672);
or U19498 (N_19498,N_17999,N_17573);
xnor U19499 (N_19499,N_18738,N_18716);
and U19500 (N_19500,N_17500,N_18732);
xor U19501 (N_19501,N_18700,N_18376);
xor U19502 (N_19502,N_18613,N_18147);
nor U19503 (N_19503,N_18022,N_17933);
nor U19504 (N_19504,N_18038,N_18532);
xor U19505 (N_19505,N_18070,N_18225);
nor U19506 (N_19506,N_18107,N_18732);
nor U19507 (N_19507,N_18533,N_18183);
or U19508 (N_19508,N_18121,N_18101);
nor U19509 (N_19509,N_18612,N_17721);
and U19510 (N_19510,N_18549,N_17918);
nand U19511 (N_19511,N_18673,N_17507);
nand U19512 (N_19512,N_17841,N_17714);
or U19513 (N_19513,N_17509,N_18509);
nand U19514 (N_19514,N_18308,N_17511);
nand U19515 (N_19515,N_18481,N_18041);
or U19516 (N_19516,N_17772,N_18166);
xor U19517 (N_19517,N_17930,N_17808);
nand U19518 (N_19518,N_18068,N_17753);
and U19519 (N_19519,N_18216,N_18683);
or U19520 (N_19520,N_18287,N_18354);
xnor U19521 (N_19521,N_18192,N_18583);
xor U19522 (N_19522,N_18721,N_17972);
xnor U19523 (N_19523,N_18120,N_18004);
nand U19524 (N_19524,N_18111,N_17972);
xnor U19525 (N_19525,N_18601,N_17942);
nand U19526 (N_19526,N_17979,N_17892);
xor U19527 (N_19527,N_17933,N_18714);
and U19528 (N_19528,N_17960,N_17990);
nand U19529 (N_19529,N_17624,N_17928);
and U19530 (N_19530,N_17964,N_17801);
nor U19531 (N_19531,N_18070,N_17644);
or U19532 (N_19532,N_18405,N_18091);
and U19533 (N_19533,N_18182,N_17840);
nor U19534 (N_19534,N_18345,N_17649);
nand U19535 (N_19535,N_18730,N_17804);
and U19536 (N_19536,N_18250,N_18570);
or U19537 (N_19537,N_17632,N_17545);
nand U19538 (N_19538,N_17752,N_18223);
xor U19539 (N_19539,N_17676,N_18096);
nand U19540 (N_19540,N_18633,N_17774);
nor U19541 (N_19541,N_17866,N_18036);
nand U19542 (N_19542,N_18362,N_18652);
xnor U19543 (N_19543,N_18160,N_17742);
nor U19544 (N_19544,N_18546,N_18160);
nor U19545 (N_19545,N_17778,N_17576);
xnor U19546 (N_19546,N_18370,N_18155);
or U19547 (N_19547,N_18203,N_18420);
nand U19548 (N_19548,N_17536,N_18403);
xor U19549 (N_19549,N_17795,N_18186);
nand U19550 (N_19550,N_18745,N_18446);
xor U19551 (N_19551,N_17868,N_18431);
xnor U19552 (N_19552,N_17854,N_18503);
and U19553 (N_19553,N_18748,N_17571);
or U19554 (N_19554,N_18200,N_17858);
and U19555 (N_19555,N_18148,N_18219);
nand U19556 (N_19556,N_17729,N_18447);
nor U19557 (N_19557,N_18548,N_18021);
nor U19558 (N_19558,N_18108,N_17992);
and U19559 (N_19559,N_18692,N_17874);
nor U19560 (N_19560,N_17945,N_18124);
xor U19561 (N_19561,N_18404,N_17912);
nand U19562 (N_19562,N_18103,N_18143);
xnor U19563 (N_19563,N_18243,N_17874);
nor U19564 (N_19564,N_18133,N_17522);
nor U19565 (N_19565,N_18108,N_17549);
nor U19566 (N_19566,N_17509,N_18465);
xnor U19567 (N_19567,N_18376,N_17554);
nand U19568 (N_19568,N_17963,N_17992);
and U19569 (N_19569,N_18105,N_18576);
nand U19570 (N_19570,N_18574,N_18116);
and U19571 (N_19571,N_18109,N_17949);
nor U19572 (N_19572,N_17800,N_18161);
nand U19573 (N_19573,N_17867,N_17512);
or U19574 (N_19574,N_17528,N_17992);
and U19575 (N_19575,N_17723,N_18513);
nor U19576 (N_19576,N_18714,N_18022);
nand U19577 (N_19577,N_18293,N_17623);
xnor U19578 (N_19578,N_18051,N_18693);
nor U19579 (N_19579,N_17901,N_17772);
nor U19580 (N_19580,N_17870,N_18405);
or U19581 (N_19581,N_17998,N_17837);
nand U19582 (N_19582,N_17578,N_18149);
and U19583 (N_19583,N_18052,N_18640);
and U19584 (N_19584,N_17878,N_18388);
xor U19585 (N_19585,N_17647,N_17941);
nor U19586 (N_19586,N_17919,N_17631);
and U19587 (N_19587,N_18397,N_17681);
nor U19588 (N_19588,N_17855,N_18615);
nand U19589 (N_19589,N_18478,N_18011);
xor U19590 (N_19590,N_18132,N_17589);
nand U19591 (N_19591,N_18303,N_18108);
nand U19592 (N_19592,N_17764,N_18413);
nor U19593 (N_19593,N_17985,N_18692);
or U19594 (N_19594,N_18486,N_17580);
and U19595 (N_19595,N_18489,N_17855);
xor U19596 (N_19596,N_18597,N_18617);
nand U19597 (N_19597,N_17771,N_18492);
nand U19598 (N_19598,N_18657,N_18592);
nand U19599 (N_19599,N_18665,N_17774);
nor U19600 (N_19600,N_17860,N_18538);
xnor U19601 (N_19601,N_18428,N_18227);
and U19602 (N_19602,N_17831,N_17859);
nor U19603 (N_19603,N_18506,N_18056);
nor U19604 (N_19604,N_17904,N_17887);
nor U19605 (N_19605,N_18617,N_17868);
nand U19606 (N_19606,N_18346,N_17961);
nand U19607 (N_19607,N_18659,N_18565);
xnor U19608 (N_19608,N_17601,N_18424);
nand U19609 (N_19609,N_18749,N_18582);
nor U19610 (N_19610,N_18578,N_18205);
nor U19611 (N_19611,N_17657,N_17726);
xor U19612 (N_19612,N_18649,N_17689);
xnor U19613 (N_19613,N_17515,N_18714);
nand U19614 (N_19614,N_18712,N_17728);
nor U19615 (N_19615,N_17958,N_17711);
nand U19616 (N_19616,N_17711,N_18502);
xor U19617 (N_19617,N_18178,N_17941);
xor U19618 (N_19618,N_18225,N_18383);
xor U19619 (N_19619,N_18172,N_17863);
nor U19620 (N_19620,N_18228,N_18364);
xor U19621 (N_19621,N_17868,N_17819);
nor U19622 (N_19622,N_18536,N_17779);
or U19623 (N_19623,N_18651,N_17536);
nand U19624 (N_19624,N_17815,N_18360);
or U19625 (N_19625,N_18171,N_18251);
nand U19626 (N_19626,N_18204,N_17867);
and U19627 (N_19627,N_18205,N_18381);
nor U19628 (N_19628,N_18527,N_18677);
or U19629 (N_19629,N_17828,N_18410);
and U19630 (N_19630,N_17962,N_18636);
nor U19631 (N_19631,N_18167,N_17578);
nand U19632 (N_19632,N_17604,N_17633);
nor U19633 (N_19633,N_18484,N_17548);
nand U19634 (N_19634,N_18157,N_18495);
xnor U19635 (N_19635,N_18169,N_18198);
and U19636 (N_19636,N_18180,N_18211);
and U19637 (N_19637,N_17765,N_17528);
xor U19638 (N_19638,N_17585,N_17654);
nand U19639 (N_19639,N_17923,N_18738);
nand U19640 (N_19640,N_17827,N_17837);
and U19641 (N_19641,N_17661,N_17850);
nor U19642 (N_19642,N_18413,N_17623);
nand U19643 (N_19643,N_18071,N_17534);
xnor U19644 (N_19644,N_17767,N_18099);
or U19645 (N_19645,N_17570,N_18516);
nor U19646 (N_19646,N_17739,N_18507);
nand U19647 (N_19647,N_18391,N_17930);
and U19648 (N_19648,N_18660,N_18162);
xnor U19649 (N_19649,N_18004,N_17519);
nor U19650 (N_19650,N_18016,N_17560);
and U19651 (N_19651,N_17566,N_18568);
xor U19652 (N_19652,N_17844,N_17787);
xnor U19653 (N_19653,N_18205,N_18049);
and U19654 (N_19654,N_18287,N_18055);
nor U19655 (N_19655,N_17797,N_17625);
and U19656 (N_19656,N_18456,N_17570);
nor U19657 (N_19657,N_18422,N_18323);
nand U19658 (N_19658,N_18056,N_18261);
nand U19659 (N_19659,N_17558,N_18487);
or U19660 (N_19660,N_17741,N_18712);
nand U19661 (N_19661,N_17931,N_18118);
and U19662 (N_19662,N_18209,N_18544);
nor U19663 (N_19663,N_18077,N_18238);
nand U19664 (N_19664,N_17898,N_17944);
xor U19665 (N_19665,N_18472,N_17996);
or U19666 (N_19666,N_17887,N_18163);
nand U19667 (N_19667,N_17970,N_17931);
and U19668 (N_19668,N_18680,N_18212);
xor U19669 (N_19669,N_18307,N_18240);
xor U19670 (N_19670,N_17768,N_17613);
and U19671 (N_19671,N_18171,N_18277);
nor U19672 (N_19672,N_17578,N_17945);
and U19673 (N_19673,N_17992,N_17959);
nand U19674 (N_19674,N_18571,N_18279);
nand U19675 (N_19675,N_18066,N_18178);
xnor U19676 (N_19676,N_18471,N_18452);
and U19677 (N_19677,N_18563,N_18684);
nor U19678 (N_19678,N_18562,N_18401);
nor U19679 (N_19679,N_18037,N_18747);
or U19680 (N_19680,N_17599,N_18369);
or U19681 (N_19681,N_18053,N_17765);
nand U19682 (N_19682,N_18371,N_18713);
nand U19683 (N_19683,N_17999,N_17595);
nand U19684 (N_19684,N_18472,N_17805);
nor U19685 (N_19685,N_18087,N_18649);
and U19686 (N_19686,N_17786,N_17941);
nor U19687 (N_19687,N_18126,N_18165);
xor U19688 (N_19688,N_18170,N_17893);
nand U19689 (N_19689,N_18748,N_17519);
or U19690 (N_19690,N_17962,N_17807);
nor U19691 (N_19691,N_17833,N_17791);
and U19692 (N_19692,N_18509,N_18733);
and U19693 (N_19693,N_17579,N_18038);
nand U19694 (N_19694,N_18118,N_18307);
nor U19695 (N_19695,N_18707,N_17999);
and U19696 (N_19696,N_17969,N_18213);
nor U19697 (N_19697,N_17658,N_18316);
nand U19698 (N_19698,N_18451,N_18149);
xor U19699 (N_19699,N_17660,N_18151);
xor U19700 (N_19700,N_18389,N_18482);
xor U19701 (N_19701,N_18379,N_18252);
or U19702 (N_19702,N_17981,N_18600);
xnor U19703 (N_19703,N_17924,N_18179);
nor U19704 (N_19704,N_18513,N_18300);
and U19705 (N_19705,N_18559,N_18453);
nand U19706 (N_19706,N_18175,N_18283);
or U19707 (N_19707,N_18458,N_17925);
nor U19708 (N_19708,N_17889,N_18659);
nand U19709 (N_19709,N_18626,N_17653);
xnor U19710 (N_19710,N_18538,N_17911);
or U19711 (N_19711,N_17679,N_17993);
or U19712 (N_19712,N_18622,N_18689);
or U19713 (N_19713,N_17732,N_18061);
xnor U19714 (N_19714,N_17905,N_17604);
nand U19715 (N_19715,N_18415,N_17991);
and U19716 (N_19716,N_17676,N_18385);
nand U19717 (N_19717,N_17804,N_18386);
or U19718 (N_19718,N_18379,N_18372);
nor U19719 (N_19719,N_18164,N_17772);
xnor U19720 (N_19720,N_18081,N_18369);
nor U19721 (N_19721,N_18371,N_18384);
and U19722 (N_19722,N_18147,N_17672);
xor U19723 (N_19723,N_18726,N_17719);
and U19724 (N_19724,N_17630,N_17605);
or U19725 (N_19725,N_17891,N_18716);
nand U19726 (N_19726,N_18051,N_18035);
xor U19727 (N_19727,N_17642,N_17529);
or U19728 (N_19728,N_17887,N_18545);
or U19729 (N_19729,N_18364,N_17584);
nor U19730 (N_19730,N_17837,N_17901);
xor U19731 (N_19731,N_18006,N_17570);
nand U19732 (N_19732,N_18236,N_17981);
or U19733 (N_19733,N_17507,N_18416);
or U19734 (N_19734,N_17615,N_18002);
nor U19735 (N_19735,N_18655,N_18567);
nand U19736 (N_19736,N_17828,N_18003);
or U19737 (N_19737,N_18122,N_18501);
nor U19738 (N_19738,N_18179,N_17502);
nor U19739 (N_19739,N_17603,N_18084);
xor U19740 (N_19740,N_18503,N_18680);
or U19741 (N_19741,N_18591,N_18194);
nor U19742 (N_19742,N_17820,N_17750);
and U19743 (N_19743,N_18082,N_18185);
nand U19744 (N_19744,N_18022,N_18160);
or U19745 (N_19745,N_17946,N_17984);
nand U19746 (N_19746,N_18098,N_17677);
and U19747 (N_19747,N_17791,N_18447);
nor U19748 (N_19748,N_17594,N_18598);
or U19749 (N_19749,N_17779,N_17693);
nor U19750 (N_19750,N_18184,N_18552);
or U19751 (N_19751,N_18742,N_18713);
or U19752 (N_19752,N_17533,N_18210);
or U19753 (N_19753,N_17829,N_17515);
xor U19754 (N_19754,N_18130,N_17784);
nor U19755 (N_19755,N_18369,N_18558);
xnor U19756 (N_19756,N_18640,N_18548);
nor U19757 (N_19757,N_18069,N_18178);
nor U19758 (N_19758,N_18488,N_18295);
nor U19759 (N_19759,N_18293,N_17544);
xor U19760 (N_19760,N_18184,N_18298);
and U19761 (N_19761,N_17964,N_17584);
nand U19762 (N_19762,N_18352,N_17673);
nand U19763 (N_19763,N_18483,N_18056);
nand U19764 (N_19764,N_17735,N_18712);
nand U19765 (N_19765,N_17982,N_17688);
nor U19766 (N_19766,N_18714,N_17587);
xor U19767 (N_19767,N_17535,N_18627);
xnor U19768 (N_19768,N_18330,N_17922);
nor U19769 (N_19769,N_17862,N_18094);
nand U19770 (N_19770,N_18303,N_17991);
or U19771 (N_19771,N_17995,N_18718);
nor U19772 (N_19772,N_17578,N_17669);
xnor U19773 (N_19773,N_18665,N_18335);
nand U19774 (N_19774,N_18283,N_18675);
and U19775 (N_19775,N_17614,N_18730);
or U19776 (N_19776,N_18037,N_18607);
nand U19777 (N_19777,N_18723,N_18569);
nand U19778 (N_19778,N_18669,N_18024);
xnor U19779 (N_19779,N_17902,N_18663);
and U19780 (N_19780,N_17843,N_18080);
nand U19781 (N_19781,N_17530,N_18147);
or U19782 (N_19782,N_18119,N_18066);
or U19783 (N_19783,N_17854,N_18185);
and U19784 (N_19784,N_17560,N_17938);
nand U19785 (N_19785,N_18056,N_18196);
xor U19786 (N_19786,N_17678,N_17901);
or U19787 (N_19787,N_17654,N_18021);
or U19788 (N_19788,N_18091,N_17933);
nor U19789 (N_19789,N_18158,N_17881);
xnor U19790 (N_19790,N_18643,N_17657);
nand U19791 (N_19791,N_17971,N_17937);
or U19792 (N_19792,N_18039,N_17941);
nor U19793 (N_19793,N_18321,N_18074);
and U19794 (N_19794,N_18416,N_17879);
nand U19795 (N_19795,N_17890,N_18561);
nor U19796 (N_19796,N_18035,N_17830);
nor U19797 (N_19797,N_17867,N_17796);
or U19798 (N_19798,N_17663,N_17516);
xor U19799 (N_19799,N_18543,N_18378);
nor U19800 (N_19800,N_18512,N_18551);
nor U19801 (N_19801,N_17683,N_17511);
nand U19802 (N_19802,N_18171,N_17848);
or U19803 (N_19803,N_18133,N_18366);
nand U19804 (N_19804,N_17903,N_18698);
and U19805 (N_19805,N_17766,N_18279);
and U19806 (N_19806,N_17917,N_17695);
and U19807 (N_19807,N_18661,N_17816);
xnor U19808 (N_19808,N_18018,N_17949);
nand U19809 (N_19809,N_18604,N_18413);
nor U19810 (N_19810,N_18076,N_17867);
or U19811 (N_19811,N_18000,N_18400);
and U19812 (N_19812,N_18098,N_17731);
or U19813 (N_19813,N_18329,N_17563);
and U19814 (N_19814,N_17754,N_18142);
or U19815 (N_19815,N_17891,N_18497);
or U19816 (N_19816,N_17830,N_17533);
and U19817 (N_19817,N_18004,N_17535);
xnor U19818 (N_19818,N_18050,N_18727);
nand U19819 (N_19819,N_18414,N_17792);
nand U19820 (N_19820,N_17878,N_17684);
xor U19821 (N_19821,N_17696,N_17983);
nand U19822 (N_19822,N_18035,N_18079);
and U19823 (N_19823,N_18112,N_18066);
xor U19824 (N_19824,N_17595,N_18212);
and U19825 (N_19825,N_17949,N_17668);
and U19826 (N_19826,N_18576,N_17507);
or U19827 (N_19827,N_18133,N_18389);
and U19828 (N_19828,N_17684,N_17626);
and U19829 (N_19829,N_17886,N_17552);
nand U19830 (N_19830,N_18068,N_18230);
nand U19831 (N_19831,N_18357,N_18015);
nor U19832 (N_19832,N_18225,N_17800);
nor U19833 (N_19833,N_18207,N_18395);
or U19834 (N_19834,N_17905,N_17856);
and U19835 (N_19835,N_18346,N_17737);
nand U19836 (N_19836,N_18130,N_18050);
nor U19837 (N_19837,N_18229,N_17876);
xor U19838 (N_19838,N_18313,N_17924);
or U19839 (N_19839,N_18503,N_18494);
xnor U19840 (N_19840,N_18080,N_18546);
xnor U19841 (N_19841,N_18648,N_18616);
xor U19842 (N_19842,N_18683,N_17744);
or U19843 (N_19843,N_17548,N_18554);
and U19844 (N_19844,N_18034,N_18153);
or U19845 (N_19845,N_18429,N_18284);
or U19846 (N_19846,N_18013,N_17820);
nor U19847 (N_19847,N_18381,N_18674);
or U19848 (N_19848,N_18406,N_17530);
nor U19849 (N_19849,N_17822,N_17862);
nor U19850 (N_19850,N_17700,N_17849);
or U19851 (N_19851,N_18425,N_17917);
xnor U19852 (N_19852,N_18283,N_17969);
xnor U19853 (N_19853,N_17957,N_18476);
xnor U19854 (N_19854,N_18329,N_18685);
nor U19855 (N_19855,N_17615,N_18267);
xor U19856 (N_19856,N_17680,N_17879);
or U19857 (N_19857,N_17951,N_17621);
or U19858 (N_19858,N_17639,N_18581);
nand U19859 (N_19859,N_18739,N_18647);
and U19860 (N_19860,N_17811,N_18668);
xnor U19861 (N_19861,N_18028,N_17948);
and U19862 (N_19862,N_17655,N_17957);
xor U19863 (N_19863,N_18120,N_18746);
nand U19864 (N_19864,N_18730,N_18256);
or U19865 (N_19865,N_18471,N_18265);
or U19866 (N_19866,N_18360,N_18496);
nand U19867 (N_19867,N_18214,N_17730);
xor U19868 (N_19868,N_17793,N_18298);
nand U19869 (N_19869,N_18626,N_18456);
nand U19870 (N_19870,N_17897,N_18457);
and U19871 (N_19871,N_17657,N_18437);
or U19872 (N_19872,N_18700,N_17714);
nor U19873 (N_19873,N_18562,N_18051);
or U19874 (N_19874,N_17962,N_17508);
or U19875 (N_19875,N_18494,N_17626);
and U19876 (N_19876,N_17550,N_18636);
nor U19877 (N_19877,N_18103,N_18113);
xor U19878 (N_19878,N_17557,N_18446);
nor U19879 (N_19879,N_18602,N_18198);
nand U19880 (N_19880,N_18329,N_18252);
xor U19881 (N_19881,N_18377,N_18281);
or U19882 (N_19882,N_18067,N_17501);
nor U19883 (N_19883,N_18633,N_17828);
nor U19884 (N_19884,N_17889,N_18579);
and U19885 (N_19885,N_18000,N_17500);
nor U19886 (N_19886,N_18390,N_17891);
and U19887 (N_19887,N_17573,N_17966);
and U19888 (N_19888,N_18363,N_17509);
xnor U19889 (N_19889,N_17603,N_18062);
xor U19890 (N_19890,N_17645,N_18656);
nand U19891 (N_19891,N_17973,N_17710);
nand U19892 (N_19892,N_17954,N_18086);
nor U19893 (N_19893,N_18054,N_17950);
xnor U19894 (N_19894,N_18353,N_18738);
or U19895 (N_19895,N_17693,N_18328);
xnor U19896 (N_19896,N_17717,N_18541);
nand U19897 (N_19897,N_18254,N_17796);
xnor U19898 (N_19898,N_17846,N_17761);
nor U19899 (N_19899,N_18427,N_18695);
nand U19900 (N_19900,N_18413,N_17929);
xnor U19901 (N_19901,N_18003,N_17802);
xor U19902 (N_19902,N_18189,N_18180);
xnor U19903 (N_19903,N_18339,N_18192);
nor U19904 (N_19904,N_18682,N_18274);
or U19905 (N_19905,N_17811,N_18652);
nor U19906 (N_19906,N_17949,N_18061);
or U19907 (N_19907,N_18182,N_18533);
nand U19908 (N_19908,N_18671,N_17794);
nand U19909 (N_19909,N_18064,N_17964);
nand U19910 (N_19910,N_18584,N_18573);
or U19911 (N_19911,N_18641,N_17864);
and U19912 (N_19912,N_18591,N_18141);
and U19913 (N_19913,N_18489,N_18710);
and U19914 (N_19914,N_18044,N_17948);
nor U19915 (N_19915,N_18005,N_17822);
or U19916 (N_19916,N_18224,N_18047);
nor U19917 (N_19917,N_17989,N_17704);
nor U19918 (N_19918,N_17689,N_18371);
xnor U19919 (N_19919,N_17869,N_17798);
xnor U19920 (N_19920,N_17642,N_18621);
and U19921 (N_19921,N_17685,N_17895);
or U19922 (N_19922,N_18186,N_18683);
and U19923 (N_19923,N_18563,N_18028);
xor U19924 (N_19924,N_17687,N_18712);
xor U19925 (N_19925,N_18730,N_18624);
nor U19926 (N_19926,N_17533,N_18150);
nor U19927 (N_19927,N_18367,N_18460);
xnor U19928 (N_19928,N_18227,N_18181);
nor U19929 (N_19929,N_17704,N_18237);
nor U19930 (N_19930,N_18712,N_17851);
or U19931 (N_19931,N_18676,N_17897);
nor U19932 (N_19932,N_18635,N_18715);
and U19933 (N_19933,N_18444,N_18465);
nor U19934 (N_19934,N_18158,N_17629);
nand U19935 (N_19935,N_18275,N_17546);
and U19936 (N_19936,N_17613,N_17509);
xor U19937 (N_19937,N_17780,N_18416);
nor U19938 (N_19938,N_17879,N_17956);
and U19939 (N_19939,N_18670,N_18456);
nand U19940 (N_19940,N_18590,N_18506);
or U19941 (N_19941,N_17812,N_18396);
or U19942 (N_19942,N_17742,N_17586);
nand U19943 (N_19943,N_18687,N_17763);
xnor U19944 (N_19944,N_18373,N_18042);
xnor U19945 (N_19945,N_18118,N_18313);
or U19946 (N_19946,N_18258,N_18396);
and U19947 (N_19947,N_18690,N_18508);
nand U19948 (N_19948,N_18429,N_17925);
or U19949 (N_19949,N_18140,N_18740);
xor U19950 (N_19950,N_18028,N_18305);
and U19951 (N_19951,N_17824,N_18138);
nand U19952 (N_19952,N_18518,N_17872);
xnor U19953 (N_19953,N_18647,N_18473);
nor U19954 (N_19954,N_18360,N_18315);
nor U19955 (N_19955,N_17772,N_17976);
or U19956 (N_19956,N_18386,N_18582);
or U19957 (N_19957,N_17936,N_18181);
and U19958 (N_19958,N_17754,N_17840);
or U19959 (N_19959,N_17914,N_17520);
xnor U19960 (N_19960,N_17617,N_17659);
xnor U19961 (N_19961,N_18522,N_17762);
or U19962 (N_19962,N_17720,N_17830);
nor U19963 (N_19963,N_18739,N_18417);
nand U19964 (N_19964,N_17658,N_17537);
and U19965 (N_19965,N_17691,N_18641);
or U19966 (N_19966,N_17833,N_18435);
xor U19967 (N_19967,N_17639,N_18446);
or U19968 (N_19968,N_18561,N_18105);
nor U19969 (N_19969,N_17517,N_18749);
nand U19970 (N_19970,N_18666,N_18237);
and U19971 (N_19971,N_17700,N_18170);
or U19972 (N_19972,N_17865,N_18105);
and U19973 (N_19973,N_17966,N_18584);
nor U19974 (N_19974,N_17651,N_18523);
xor U19975 (N_19975,N_18610,N_17652);
xor U19976 (N_19976,N_18304,N_18495);
or U19977 (N_19977,N_18205,N_17803);
nand U19978 (N_19978,N_18432,N_17912);
nor U19979 (N_19979,N_17712,N_18038);
nand U19980 (N_19980,N_18461,N_18355);
nor U19981 (N_19981,N_17974,N_18622);
or U19982 (N_19982,N_17866,N_18739);
xor U19983 (N_19983,N_18072,N_18096);
nand U19984 (N_19984,N_18447,N_18371);
or U19985 (N_19985,N_18058,N_17505);
or U19986 (N_19986,N_17845,N_17880);
nor U19987 (N_19987,N_18355,N_18681);
and U19988 (N_19988,N_18638,N_18437);
and U19989 (N_19989,N_17694,N_17670);
xor U19990 (N_19990,N_18610,N_18088);
nand U19991 (N_19991,N_18723,N_17634);
xor U19992 (N_19992,N_18286,N_18324);
and U19993 (N_19993,N_17673,N_17745);
xor U19994 (N_19994,N_18725,N_18109);
xnor U19995 (N_19995,N_18126,N_18202);
xor U19996 (N_19996,N_18705,N_17614);
nor U19997 (N_19997,N_18330,N_17943);
and U19998 (N_19998,N_17965,N_18393);
xor U19999 (N_19999,N_18518,N_17752);
nor U20000 (N_20000,N_19797,N_19265);
and U20001 (N_20001,N_18776,N_19284);
or U20002 (N_20002,N_19206,N_19654);
nand U20003 (N_20003,N_19824,N_19735);
or U20004 (N_20004,N_19699,N_19293);
nor U20005 (N_20005,N_19328,N_19663);
or U20006 (N_20006,N_18933,N_18765);
xnor U20007 (N_20007,N_18863,N_19934);
nor U20008 (N_20008,N_19147,N_19862);
nand U20009 (N_20009,N_19003,N_19698);
nand U20010 (N_20010,N_19083,N_19789);
nor U20011 (N_20011,N_19307,N_19141);
nand U20012 (N_20012,N_19203,N_19425);
xnor U20013 (N_20013,N_19967,N_18986);
nand U20014 (N_20014,N_18750,N_19551);
or U20015 (N_20015,N_19977,N_19481);
or U20016 (N_20016,N_18910,N_18808);
xor U20017 (N_20017,N_18850,N_19343);
nand U20018 (N_20018,N_19847,N_19189);
or U20019 (N_20019,N_19867,N_19592);
and U20020 (N_20020,N_19113,N_19950);
and U20021 (N_20021,N_19619,N_18844);
nand U20022 (N_20022,N_19350,N_19010);
nand U20023 (N_20023,N_19721,N_19980);
or U20024 (N_20024,N_18780,N_19348);
or U20025 (N_20025,N_19471,N_19216);
or U20026 (N_20026,N_19391,N_19669);
nand U20027 (N_20027,N_19122,N_19812);
or U20028 (N_20028,N_18859,N_19543);
xnor U20029 (N_20029,N_19384,N_19016);
or U20030 (N_20030,N_19261,N_18928);
and U20031 (N_20031,N_18921,N_18895);
and U20032 (N_20032,N_18820,N_19837);
xnor U20033 (N_20033,N_19170,N_19869);
nor U20034 (N_20034,N_19478,N_19389);
xnor U20035 (N_20035,N_19930,N_19295);
and U20036 (N_20036,N_19532,N_19563);
and U20037 (N_20037,N_19683,N_18977);
or U20038 (N_20038,N_19406,N_19033);
xnor U20039 (N_20039,N_19136,N_19194);
xor U20040 (N_20040,N_19831,N_19883);
or U20041 (N_20041,N_19248,N_19052);
nor U20042 (N_20042,N_18826,N_19828);
and U20043 (N_20043,N_19430,N_19873);
xnor U20044 (N_20044,N_19360,N_19520);
nand U20045 (N_20045,N_19947,N_19125);
and U20046 (N_20046,N_19905,N_19413);
nand U20047 (N_20047,N_19457,N_19143);
and U20048 (N_20048,N_19848,N_19688);
and U20049 (N_20049,N_19130,N_19567);
and U20050 (N_20050,N_19103,N_19435);
nor U20051 (N_20051,N_18785,N_18969);
nand U20052 (N_20052,N_19943,N_19436);
and U20053 (N_20053,N_19954,N_19317);
or U20054 (N_20054,N_19054,N_19658);
and U20055 (N_20055,N_19507,N_19599);
nand U20056 (N_20056,N_19393,N_19465);
and U20057 (N_20057,N_19936,N_19111);
nor U20058 (N_20058,N_19585,N_19000);
or U20059 (N_20059,N_19020,N_19500);
and U20060 (N_20060,N_18796,N_19556);
xnor U20061 (N_20061,N_18817,N_19770);
xnor U20062 (N_20062,N_19530,N_19202);
xor U20063 (N_20063,N_19888,N_19925);
or U20064 (N_20064,N_19745,N_19615);
nand U20065 (N_20065,N_19055,N_19723);
or U20066 (N_20066,N_19605,N_19446);
xor U20067 (N_20067,N_19805,N_18752);
and U20068 (N_20068,N_19221,N_18990);
xor U20069 (N_20069,N_19233,N_18989);
xnor U20070 (N_20070,N_19749,N_18793);
xnor U20071 (N_20071,N_19537,N_19002);
nand U20072 (N_20072,N_18950,N_19262);
and U20073 (N_20073,N_19971,N_18922);
nor U20074 (N_20074,N_18811,N_19800);
nor U20075 (N_20075,N_19383,N_19292);
or U20076 (N_20076,N_19713,N_19795);
xor U20077 (N_20077,N_18880,N_19427);
xor U20078 (N_20078,N_19172,N_19548);
nor U20079 (N_20079,N_19414,N_19356);
nand U20080 (N_20080,N_19129,N_19839);
xor U20081 (N_20081,N_19112,N_18988);
or U20082 (N_20082,N_19833,N_19462);
nor U20083 (N_20083,N_18951,N_18919);
nor U20084 (N_20084,N_18941,N_19774);
nand U20085 (N_20085,N_18839,N_19149);
nand U20086 (N_20086,N_18886,N_19410);
nand U20087 (N_20087,N_19378,N_18974);
xor U20088 (N_20088,N_19140,N_19794);
nand U20089 (N_20089,N_18829,N_19322);
and U20090 (N_20090,N_19215,N_19526);
nand U20091 (N_20091,N_19246,N_18783);
nor U20092 (N_20092,N_18923,N_19309);
nor U20093 (N_20093,N_19429,N_18760);
nand U20094 (N_20094,N_19063,N_19305);
nand U20095 (N_20095,N_18966,N_19155);
nor U20096 (N_20096,N_19761,N_19211);
xor U20097 (N_20097,N_19252,N_19027);
nand U20098 (N_20098,N_19102,N_19842);
nand U20099 (N_20099,N_18991,N_19270);
and U20100 (N_20100,N_19240,N_19249);
or U20101 (N_20101,N_19219,N_19212);
xnor U20102 (N_20102,N_19546,N_18784);
xor U20103 (N_20103,N_18799,N_18984);
xor U20104 (N_20104,N_19926,N_19695);
xor U20105 (N_20105,N_18803,N_18963);
nand U20106 (N_20106,N_19659,N_19386);
nand U20107 (N_20107,N_19744,N_19999);
xnor U20108 (N_20108,N_19989,N_19367);
and U20109 (N_20109,N_19816,N_19299);
xnor U20110 (N_20110,N_19268,N_19983);
xnor U20111 (N_20111,N_18878,N_18836);
and U20112 (N_20112,N_19804,N_19998);
or U20113 (N_20113,N_19613,N_19696);
or U20114 (N_20114,N_18949,N_18864);
nand U20115 (N_20115,N_19354,N_19370);
and U20116 (N_20116,N_19453,N_19319);
or U20117 (N_20117,N_19612,N_19561);
nor U20118 (N_20118,N_19437,N_18889);
and U20119 (N_20119,N_19773,N_19618);
or U20120 (N_20120,N_19084,N_18893);
nor U20121 (N_20121,N_18801,N_19889);
xnor U20122 (N_20122,N_18792,N_19065);
xnor U20123 (N_20123,N_19985,N_18815);
nand U20124 (N_20124,N_18913,N_18993);
and U20125 (N_20125,N_19388,N_19637);
or U20126 (N_20126,N_19739,N_19362);
xnor U20127 (N_20127,N_19366,N_19036);
or U20128 (N_20128,N_19836,N_19979);
nand U20129 (N_20129,N_18885,N_19126);
nand U20130 (N_20130,N_19693,N_19668);
or U20131 (N_20131,N_18800,N_19379);
or U20132 (N_20132,N_19093,N_19604);
nor U20133 (N_20133,N_18944,N_19376);
nor U20134 (N_20134,N_19772,N_19336);
or U20135 (N_20135,N_19929,N_19256);
xnor U20136 (N_20136,N_18847,N_19893);
nor U20137 (N_20137,N_19857,N_19482);
and U20138 (N_20138,N_19213,N_19961);
or U20139 (N_20139,N_19234,N_19579);
or U20140 (N_20140,N_19959,N_19080);
xor U20141 (N_20141,N_19928,N_19062);
nor U20142 (N_20142,N_18809,N_19220);
xor U20143 (N_20143,N_19759,N_19920);
nor U20144 (N_20144,N_19371,N_19734);
xnor U20145 (N_20145,N_19667,N_19493);
and U20146 (N_20146,N_18825,N_19509);
or U20147 (N_20147,N_19756,N_19564);
and U20148 (N_20148,N_19499,N_19819);
nor U20149 (N_20149,N_19827,N_19621);
xnor U20150 (N_20150,N_19374,N_19455);
and U20151 (N_20151,N_19404,N_19135);
or U20152 (N_20152,N_18860,N_19022);
nor U20153 (N_20153,N_19301,N_18979);
and U20154 (N_20154,N_19898,N_19602);
or U20155 (N_20155,N_19673,N_19878);
nand U20156 (N_20156,N_19716,N_19958);
and U20157 (N_20157,N_18866,N_19214);
nand U20158 (N_20158,N_18753,N_18769);
nor U20159 (N_20159,N_19392,N_19736);
nor U20160 (N_20160,N_18952,N_18835);
nor U20161 (N_20161,N_19835,N_19448);
and U20162 (N_20162,N_19809,N_19165);
xnor U20163 (N_20163,N_18837,N_19762);
xor U20164 (N_20164,N_19200,N_19331);
nand U20165 (N_20165,N_18907,N_18787);
xnor U20166 (N_20166,N_19259,N_19900);
nand U20167 (N_20167,N_18828,N_19986);
xnor U20168 (N_20168,N_19045,N_19401);
or U20169 (N_20169,N_19689,N_19818);
nand U20170 (N_20170,N_19134,N_19487);
nand U20171 (N_20171,N_18940,N_19628);
or U20172 (N_20172,N_19533,N_18834);
or U20173 (N_20173,N_19450,N_19583);
nor U20174 (N_20174,N_18795,N_19005);
and U20175 (N_20175,N_18872,N_18773);
nand U20176 (N_20176,N_19163,N_19255);
nor U20177 (N_20177,N_18934,N_19086);
nand U20178 (N_20178,N_19609,N_19814);
nor U20179 (N_20179,N_18775,N_19335);
nand U20180 (N_20180,N_19186,N_18807);
or U20181 (N_20181,N_19639,N_19491);
or U20182 (N_20182,N_19232,N_18888);
nor U20183 (N_20183,N_18833,N_19917);
nand U20184 (N_20184,N_18911,N_19787);
or U20185 (N_20185,N_19880,N_19196);
nand U20186 (N_20186,N_19629,N_19960);
nor U20187 (N_20187,N_18915,N_19117);
xnor U20188 (N_20188,N_19865,N_19786);
or U20189 (N_20189,N_19159,N_19297);
nor U20190 (N_20190,N_19651,N_19251);
nand U20191 (N_20191,N_19238,N_18822);
and U20192 (N_20192,N_18912,N_19023);
and U20193 (N_20193,N_19421,N_19534);
and U20194 (N_20194,N_19486,N_19048);
nand U20195 (N_20195,N_18802,N_19638);
and U20196 (N_20196,N_19715,N_19451);
and U20197 (N_20197,N_19078,N_18967);
xor U20198 (N_20198,N_18790,N_19966);
nand U20199 (N_20199,N_19566,N_19190);
xnor U20200 (N_20200,N_19116,N_19510);
or U20201 (N_20201,N_18827,N_19664);
nand U20202 (N_20202,N_19737,N_19515);
and U20203 (N_20203,N_18840,N_19577);
nor U20204 (N_20204,N_19188,N_19718);
and U20205 (N_20205,N_19523,N_19044);
or U20206 (N_20206,N_19963,N_19817);
and U20207 (N_20207,N_18972,N_19908);
nor U20208 (N_20208,N_19105,N_19559);
nor U20209 (N_20209,N_19173,N_18946);
and U20210 (N_20210,N_18854,N_19702);
nor U20211 (N_20211,N_19802,N_19104);
nand U20212 (N_20212,N_19747,N_19792);
nor U20213 (N_20213,N_19394,N_19175);
or U20214 (N_20214,N_19552,N_19881);
or U20215 (N_20215,N_19131,N_19426);
nor U20216 (N_20216,N_19573,N_19813);
and U20217 (N_20217,N_19623,N_19607);
and U20218 (N_20218,N_18812,N_19239);
nor U20219 (N_20219,N_19514,N_19281);
nand U20220 (N_20220,N_19349,N_18848);
xor U20221 (N_20221,N_19082,N_18901);
nand U20222 (N_20222,N_19750,N_18973);
nor U20223 (N_20223,N_19488,N_19754);
xnor U20224 (N_20224,N_19850,N_19798);
and U20225 (N_20225,N_19570,N_19508);
xnor U20226 (N_20226,N_19919,N_19369);
xor U20227 (N_20227,N_19108,N_19397);
or U20228 (N_20228,N_19545,N_19539);
xor U20229 (N_20229,N_19464,N_19157);
nor U20230 (N_20230,N_19915,N_19832);
and U20231 (N_20231,N_19784,N_19625);
nor U20232 (N_20232,N_18905,N_19810);
or U20233 (N_20233,N_19118,N_19763);
or U20234 (N_20234,N_18824,N_19390);
nor U20235 (N_20235,N_19940,N_19517);
or U20236 (N_20236,N_19557,N_19286);
and U20237 (N_20237,N_19655,N_18892);
xor U20238 (N_20238,N_19923,N_19984);
nor U20239 (N_20239,N_19308,N_19886);
nor U20240 (N_20240,N_19475,N_19549);
xor U20241 (N_20241,N_19617,N_19632);
nor U20242 (N_20242,N_19304,N_19236);
nor U20243 (N_20243,N_18882,N_19871);
and U20244 (N_20244,N_19182,N_18939);
nand U20245 (N_20245,N_18903,N_19001);
and U20246 (N_20246,N_19645,N_19948);
xnor U20247 (N_20247,N_18948,N_19741);
and U20248 (N_20248,N_19909,N_19555);
xnor U20249 (N_20249,N_18992,N_19808);
and U20250 (N_20250,N_19161,N_18877);
xnor U20251 (N_20251,N_19185,N_18916);
and U20252 (N_20252,N_19064,N_19341);
nand U20253 (N_20253,N_19581,N_18960);
nand U20254 (N_20254,N_19851,N_18865);
or U20255 (N_20255,N_19043,N_19859);
xnor U20256 (N_20256,N_19142,N_19580);
or U20257 (N_20257,N_19438,N_19092);
xnor U20258 (N_20258,N_19137,N_19780);
xnor U20259 (N_20259,N_19941,N_19516);
nor U20260 (N_20260,N_19300,N_19004);
nand U20261 (N_20261,N_19433,N_18788);
nand U20262 (N_20262,N_18971,N_19152);
and U20263 (N_20263,N_19973,N_19075);
xor U20264 (N_20264,N_18902,N_18962);
or U20265 (N_20265,N_18798,N_19569);
and U20266 (N_20266,N_19965,N_18771);
or U20267 (N_20267,N_19160,N_19411);
nor U20268 (N_20268,N_19237,N_19423);
or U20269 (N_20269,N_19952,N_19697);
xnor U20270 (N_20270,N_19225,N_19751);
nor U20271 (N_20271,N_19024,N_19353);
nand U20272 (N_20272,N_19858,N_19642);
xnor U20273 (N_20273,N_19227,N_19049);
and U20274 (N_20274,N_19272,N_19562);
nor U20275 (N_20275,N_19907,N_19742);
and U20276 (N_20276,N_18861,N_18761);
xor U20277 (N_20277,N_18985,N_19266);
or U20278 (N_20278,N_19730,N_19606);
xnor U20279 (N_20279,N_19198,N_19710);
or U20280 (N_20280,N_19224,N_19492);
xnor U20281 (N_20281,N_18810,N_19096);
nand U20282 (N_20282,N_19626,N_19402);
and U20283 (N_20283,N_19806,N_19993);
or U20284 (N_20284,N_19167,N_19403);
nor U20285 (N_20285,N_19372,N_19290);
or U20286 (N_20286,N_19325,N_19724);
nor U20287 (N_20287,N_19456,N_19554);
xnor U20288 (N_20288,N_18898,N_19978);
nor U20289 (N_20289,N_19899,N_18929);
nand U20290 (N_20290,N_19826,N_19714);
or U20291 (N_20291,N_19076,N_19633);
and U20292 (N_20292,N_19743,N_19037);
or U20293 (N_20293,N_19729,N_19030);
nand U20294 (N_20294,N_19527,N_19995);
and U20295 (N_20295,N_19578,N_19686);
or U20296 (N_20296,N_19298,N_19375);
nand U20297 (N_20297,N_19138,N_19957);
and U20298 (N_20298,N_18978,N_19017);
nor U20299 (N_20299,N_19921,N_19692);
nand U20300 (N_20300,N_19834,N_19849);
nor U20301 (N_20301,N_19665,N_19241);
or U20302 (N_20302,N_19846,N_19187);
and U20303 (N_20303,N_19195,N_18982);
nand U20304 (N_20304,N_19422,N_19666);
or U20305 (N_20305,N_19904,N_19582);
nand U20306 (N_20306,N_19635,N_19156);
and U20307 (N_20307,N_18762,N_19649);
nand U20308 (N_20308,N_19407,N_19511);
and U20309 (N_20309,N_19882,N_18954);
or U20310 (N_20310,N_19418,N_19970);
nor U20311 (N_20311,N_19459,N_19019);
and U20312 (N_20312,N_19709,N_19193);
xnor U20313 (N_20313,N_19498,N_19988);
or U20314 (N_20314,N_19870,N_19652);
nand U20315 (N_20315,N_19646,N_19521);
nor U20316 (N_20316,N_19788,N_18959);
nor U20317 (N_20317,N_19106,N_19591);
xor U20318 (N_20318,N_19506,N_19822);
and U20319 (N_20319,N_19531,N_19364);
xnor U20320 (N_20320,N_19181,N_19755);
nor U20321 (N_20321,N_19553,N_19071);
and U20322 (N_20322,N_19326,N_19576);
xor U20323 (N_20323,N_18896,N_19672);
and U20324 (N_20324,N_19489,N_18937);
nand U20325 (N_20325,N_19535,N_19976);
xor U20326 (N_20326,N_19056,N_18876);
or U20327 (N_20327,N_19962,N_19110);
xor U20328 (N_20328,N_19708,N_18851);
nand U20329 (N_20329,N_19053,N_19616);
nand U20330 (N_20330,N_19614,N_19327);
or U20331 (N_20331,N_19903,N_19906);
nand U20332 (N_20332,N_19547,N_19895);
xor U20333 (N_20333,N_19031,N_19179);
and U20334 (N_20334,N_19280,N_19257);
nand U20335 (N_20335,N_19679,N_19365);
xnor U20336 (N_20336,N_19201,N_19294);
nor U20337 (N_20337,N_19235,N_19287);
nor U20338 (N_20338,N_19176,N_18887);
and U20339 (N_20339,N_18853,N_19911);
xor U20340 (N_20340,N_19409,N_18947);
nand U20341 (N_20341,N_18884,N_19853);
or U20342 (N_20342,N_19525,N_19914);
or U20343 (N_20343,N_19796,N_19345);
or U20344 (N_20344,N_19440,N_19408);
and U20345 (N_20345,N_19803,N_19811);
nor U20346 (N_20346,N_19154,N_19505);
or U20347 (N_20347,N_18754,N_18768);
and U20348 (N_20348,N_19332,N_19277);
xor U20349 (N_20349,N_19099,N_19497);
and U20350 (N_20350,N_18955,N_19191);
nor U20351 (N_20351,N_19843,N_19342);
and U20352 (N_20352,N_19166,N_19012);
or U20353 (N_20353,N_19197,N_19685);
or U20354 (N_20354,N_19671,N_19057);
xnor U20355 (N_20355,N_19283,N_19544);
xor U20356 (N_20356,N_19042,N_18816);
xor U20357 (N_20357,N_19779,N_19059);
xnor U20358 (N_20358,N_19495,N_18927);
nand U20359 (N_20359,N_19334,N_19677);
and U20360 (N_20360,N_19139,N_19969);
nor U20361 (N_20361,N_19434,N_19412);
xor U20362 (N_20362,N_19778,N_19598);
or U20363 (N_20363,N_19355,N_19385);
nand U20364 (N_20364,N_19400,N_18999);
nand U20365 (N_20365,N_19035,N_19089);
nand U20366 (N_20366,N_19069,N_19377);
or U20367 (N_20367,N_19706,N_18930);
xor U20368 (N_20368,N_19600,N_18821);
and U20369 (N_20369,N_19072,N_19018);
xnor U20370 (N_20370,N_19250,N_19046);
or U20371 (N_20371,N_19924,N_18909);
and U20372 (N_20372,N_19324,N_18994);
xor U20373 (N_20373,N_19479,N_19070);
xnor U20374 (N_20374,N_19177,N_19395);
or U20375 (N_20375,N_19522,N_18764);
nand U20376 (N_20376,N_19758,N_19469);
and U20377 (N_20377,N_18899,N_19114);
and U20378 (N_20378,N_19311,N_19123);
and U20379 (N_20379,N_18778,N_19560);
nand U20380 (N_20380,N_19991,N_18996);
xor U20381 (N_20381,N_18871,N_19678);
nand U20382 (N_20382,N_19145,N_19944);
and U20383 (N_20383,N_18814,N_19657);
or U20384 (N_20384,N_19029,N_19597);
nor U20385 (N_20385,N_19705,N_18856);
nor U20386 (N_20386,N_19443,N_19992);
and U20387 (N_20387,N_18805,N_18806);
or U20388 (N_20388,N_19861,N_18995);
nor U20389 (N_20389,N_19868,N_19068);
or U20390 (N_20390,N_19624,N_19968);
xor U20391 (N_20391,N_19051,N_18879);
xor U20392 (N_20392,N_19876,N_19329);
or U20393 (N_20393,N_19519,N_19931);
and U20394 (N_20394,N_18782,N_19278);
xnor U20395 (N_20395,N_19449,N_18897);
nor U20396 (N_20396,N_19444,N_19694);
nor U20397 (N_20397,N_19653,N_19513);
nor U20398 (N_20398,N_19279,N_19684);
xnor U20399 (N_20399,N_19222,N_19799);
and U20400 (N_20400,N_18770,N_18920);
or U20401 (N_20401,N_19447,N_18819);
and U20402 (N_20402,N_19040,N_18766);
nor U20403 (N_20403,N_19073,N_19034);
or U20404 (N_20404,N_19589,N_19975);
or U20405 (N_20405,N_19050,N_19707);
and U20406 (N_20406,N_19269,N_18794);
xnor U20407 (N_20407,N_19863,N_18874);
and U20408 (N_20408,N_19996,N_18759);
xor U20409 (N_20409,N_19276,N_19720);
nor U20410 (N_20410,N_19396,N_19011);
nand U20411 (N_20411,N_19782,N_19381);
or U20412 (N_20412,N_19872,N_18831);
or U20413 (N_20413,N_19601,N_18917);
nor U20414 (N_20414,N_18767,N_19387);
and U20415 (N_20415,N_18964,N_18818);
xnor U20416 (N_20416,N_19575,N_19061);
nor U20417 (N_20417,N_18965,N_19622);
nor U20418 (N_20418,N_19680,N_19949);
nand U20419 (N_20419,N_19725,N_19351);
xnor U20420 (N_20420,N_19641,N_19209);
nand U20421 (N_20421,N_18890,N_18774);
nor U20422 (N_20422,N_19727,N_19901);
nor U20423 (N_20423,N_19550,N_19226);
and U20424 (N_20424,N_18908,N_19006);
nor U20425 (N_20425,N_19128,N_18838);
and U20426 (N_20426,N_19074,N_19424);
or U20427 (N_20427,N_19910,N_19184);
and U20428 (N_20428,N_19603,N_19574);
nand U20429 (N_20429,N_18958,N_19503);
nor U20430 (N_20430,N_19518,N_19303);
or U20431 (N_20431,N_19229,N_19008);
nor U20432 (N_20432,N_18935,N_19169);
nand U20433 (N_20433,N_19494,N_19874);
or U20434 (N_20434,N_19087,N_19101);
xnor U20435 (N_20435,N_19662,N_19109);
nor U20436 (N_20436,N_19643,N_19468);
or U20437 (N_20437,N_19178,N_18813);
xor U20438 (N_20438,N_19890,N_18961);
nor U20439 (N_20439,N_19289,N_19100);
or U20440 (N_20440,N_18980,N_19793);
or U20441 (N_20441,N_19442,N_19254);
and U20442 (N_20442,N_19470,N_19891);
or U20443 (N_20443,N_19703,N_19913);
and U20444 (N_20444,N_18830,N_18924);
and U20445 (N_20445,N_19887,N_18956);
and U20446 (N_20446,N_19825,N_19361);
and U20447 (N_20447,N_19399,N_19768);
nor U20448 (N_20448,N_19912,N_19820);
and U20449 (N_20449,N_19733,N_19753);
xnor U20450 (N_20450,N_19452,N_19337);
nor U20451 (N_20451,N_19151,N_19719);
and U20452 (N_20452,N_19781,N_19852);
and U20453 (N_20453,N_19982,N_19608);
nand U20454 (N_20454,N_19752,N_19318);
xnor U20455 (N_20455,N_19260,N_19879);
and U20456 (N_20456,N_19015,N_19939);
nor U20457 (N_20457,N_19748,N_19997);
and U20458 (N_20458,N_19077,N_19210);
xor U20459 (N_20459,N_19807,N_19783);
nor U20460 (N_20460,N_19775,N_19765);
nand U20461 (N_20461,N_19458,N_19041);
xor U20462 (N_20462,N_19026,N_19524);
and U20463 (N_20463,N_18862,N_18900);
xnor U20464 (N_20464,N_19922,N_19081);
nor U20465 (N_20465,N_18843,N_19316);
nand U20466 (N_20466,N_19593,N_18906);
nor U20467 (N_20467,N_19660,N_19472);
or U20468 (N_20468,N_19158,N_18987);
xor U20469 (N_20469,N_18953,N_19476);
xnor U20470 (N_20470,N_18881,N_18931);
nor U20471 (N_20471,N_19338,N_18976);
or U20472 (N_20472,N_18868,N_19504);
and U20473 (N_20473,N_19009,N_19230);
or U20474 (N_20474,N_19636,N_19704);
nand U20475 (N_20475,N_19892,N_19528);
nor U20476 (N_20476,N_19382,N_19540);
and U20477 (N_20477,N_19032,N_19150);
and U20478 (N_20478,N_18823,N_19771);
nor U20479 (N_20479,N_19791,N_19007);
or U20480 (N_20480,N_19285,N_19946);
nor U20481 (N_20481,N_18781,N_19485);
nand U20482 (N_20482,N_19039,N_19572);
nand U20483 (N_20483,N_18870,N_19512);
and U20484 (N_20484,N_19315,N_18777);
or U20485 (N_20485,N_19320,N_19955);
or U20486 (N_20486,N_19314,N_19088);
and U20487 (N_20487,N_18757,N_19352);
nand U20488 (N_20488,N_19467,N_19640);
and U20489 (N_20489,N_19047,N_19496);
xnor U20490 (N_20490,N_19830,N_19483);
xor U20491 (N_20491,N_19712,N_19454);
xor U20492 (N_20492,N_18772,N_19769);
nand U20493 (N_20493,N_19359,N_19243);
nor U20494 (N_20494,N_19484,N_19885);
xor U20495 (N_20495,N_19542,N_19417);
or U20496 (N_20496,N_19231,N_19144);
or U20497 (N_20497,N_19956,N_19121);
nand U20498 (N_20498,N_18957,N_19306);
nor U20499 (N_20499,N_19648,N_18846);
nand U20500 (N_20500,N_19460,N_19363);
nor U20501 (N_20501,N_19821,N_19596);
nor U20502 (N_20502,N_19711,N_19757);
nand U20503 (N_20503,N_19823,N_18926);
nor U20504 (N_20504,N_18855,N_19529);
xor U20505 (N_20505,N_19380,N_19728);
and U20506 (N_20506,N_19066,N_19373);
xnor U20507 (N_20507,N_19933,N_19884);
nand U20508 (N_20508,N_18894,N_19937);
nand U20509 (N_20509,N_19875,N_19223);
and U20510 (N_20510,N_19098,N_19171);
xnor U20511 (N_20511,N_19148,N_19676);
nor U20512 (N_20512,N_18970,N_19358);
nor U20513 (N_20513,N_19945,N_19275);
xor U20514 (N_20514,N_19845,N_19133);
nor U20515 (N_20515,N_19687,N_19162);
nand U20516 (N_20516,N_19038,N_19815);
xnor U20517 (N_20517,N_19474,N_19731);
xor U20518 (N_20518,N_19981,N_19439);
nand U20519 (N_20519,N_19942,N_19333);
nor U20520 (N_20520,N_19856,N_19670);
and U20521 (N_20521,N_19726,N_19264);
xor U20522 (N_20522,N_19902,N_18981);
and U20523 (N_20523,N_19094,N_19538);
xor U20524 (N_20524,N_19310,N_18867);
xor U20525 (N_20525,N_19700,N_19079);
xor U20526 (N_20526,N_19296,N_19866);
nand U20527 (N_20527,N_19860,N_19199);
xor U20528 (N_20528,N_19247,N_19897);
xor U20529 (N_20529,N_19776,N_19766);
xor U20530 (N_20530,N_19953,N_19841);
nand U20531 (N_20531,N_19346,N_18983);
and U20532 (N_20532,N_19764,N_19935);
nand U20533 (N_20533,N_19661,N_19253);
nand U20534 (N_20534,N_18832,N_19312);
or U20535 (N_20535,N_18914,N_19650);
nor U20536 (N_20536,N_19441,N_19620);
xnor U20537 (N_20537,N_19674,N_19938);
nand U20538 (N_20538,N_19431,N_18869);
or U20539 (N_20539,N_18875,N_19398);
nor U20540 (N_20540,N_19801,N_19894);
or U20541 (N_20541,N_19445,N_19501);
nor U20542 (N_20542,N_19586,N_19119);
xor U20543 (N_20543,N_19245,N_19675);
xnor U20544 (N_20544,N_19419,N_18756);
nand U20545 (N_20545,N_18925,N_18858);
xnor U20546 (N_20546,N_18975,N_19558);
and U20547 (N_20547,N_18758,N_19477);
and U20548 (N_20548,N_19502,N_19288);
xor U20549 (N_20549,N_19990,N_19368);
nand U20550 (N_20550,N_19028,N_19584);
xnor U20551 (N_20551,N_19767,N_19595);
or U20552 (N_20552,N_19473,N_18968);
nand U20553 (N_20553,N_19014,N_19844);
nor U20554 (N_20554,N_19095,N_19571);
nand U20555 (N_20555,N_19656,N_18998);
xnor U20556 (N_20556,N_19717,N_19271);
xnor U20557 (N_20557,N_19263,N_19916);
nand U20558 (N_20558,N_19174,N_19242);
or U20559 (N_20559,N_19013,N_19060);
nand U20560 (N_20560,N_19205,N_19896);
nand U20561 (N_20561,N_19330,N_19644);
and U20562 (N_20562,N_19590,N_18797);
nand U20563 (N_20563,N_19097,N_19273);
and U20564 (N_20564,N_19339,N_19588);
and U20565 (N_20565,N_18779,N_19415);
nor U20566 (N_20566,N_18942,N_19701);
nor U20567 (N_20567,N_19740,N_19738);
xor U20568 (N_20568,N_18997,N_19428);
or U20569 (N_20569,N_19918,N_19480);
nor U20570 (N_20570,N_19168,N_19932);
xor U20571 (N_20571,N_18918,N_19994);
nand U20572 (N_20572,N_18849,N_19258);
nor U20573 (N_20573,N_19228,N_18804);
nand U20574 (N_20574,N_19274,N_19565);
and U20575 (N_20575,N_19972,N_19085);
nand U20576 (N_20576,N_19146,N_19777);
and U20577 (N_20577,N_19090,N_18842);
and U20578 (N_20578,N_19127,N_19405);
xnor U20579 (N_20579,N_19153,N_19855);
nand U20580 (N_20580,N_19927,N_19107);
nand U20581 (N_20581,N_19323,N_19067);
nor U20582 (N_20582,N_19951,N_19340);
or U20583 (N_20583,N_19877,N_18786);
and U20584 (N_20584,N_19987,N_19634);
or U20585 (N_20585,N_19690,N_19302);
nor U20586 (N_20586,N_19722,N_19760);
nand U20587 (N_20587,N_19785,N_19536);
and U20588 (N_20588,N_19461,N_19124);
or U20589 (N_20589,N_19091,N_19631);
and U20590 (N_20590,N_19291,N_19321);
nand U20591 (N_20591,N_19682,N_18883);
or U20592 (N_20592,N_19120,N_19192);
nor U20593 (N_20593,N_19974,N_19829);
nand U20594 (N_20594,N_18945,N_19164);
nand U20595 (N_20595,N_19541,N_19691);
and U20596 (N_20596,N_19204,N_18873);
and U20597 (N_20597,N_18891,N_19490);
and U20598 (N_20598,N_18943,N_18932);
nand U20599 (N_20599,N_19838,N_18763);
nor U20600 (N_20600,N_19347,N_19183);
nand U20601 (N_20601,N_19681,N_18936);
nor U20602 (N_20602,N_18841,N_18857);
nand U20603 (N_20603,N_19568,N_19357);
nor U20604 (N_20604,N_19611,N_18845);
nand U20605 (N_20605,N_18938,N_19466);
nand U20606 (N_20606,N_18791,N_19463);
and U20607 (N_20607,N_19267,N_19790);
and U20608 (N_20608,N_19218,N_19746);
and U20609 (N_20609,N_19420,N_19587);
and U20610 (N_20610,N_19610,N_19217);
nand U20611 (N_20611,N_19416,N_19180);
nor U20612 (N_20612,N_18852,N_19115);
nand U20613 (N_20613,N_18751,N_19630);
nand U20614 (N_20614,N_19647,N_19627);
or U20615 (N_20615,N_18904,N_19864);
or U20616 (N_20616,N_19282,N_19594);
nor U20617 (N_20617,N_18755,N_19432);
nor U20618 (N_20618,N_18789,N_19025);
xnor U20619 (N_20619,N_19840,N_19313);
nand U20620 (N_20620,N_19854,N_19244);
xor U20621 (N_20621,N_19344,N_19208);
nand U20622 (N_20622,N_19964,N_19732);
xnor U20623 (N_20623,N_19207,N_19058);
nand U20624 (N_20624,N_19021,N_19132);
xnor U20625 (N_20625,N_18995,N_19035);
and U20626 (N_20626,N_19227,N_19832);
xnor U20627 (N_20627,N_19274,N_19458);
or U20628 (N_20628,N_19044,N_19901);
xnor U20629 (N_20629,N_19337,N_19568);
xor U20630 (N_20630,N_19601,N_19133);
xnor U20631 (N_20631,N_19306,N_18782);
nand U20632 (N_20632,N_19407,N_19174);
nand U20633 (N_20633,N_18871,N_19451);
and U20634 (N_20634,N_19836,N_18899);
or U20635 (N_20635,N_19746,N_19253);
nand U20636 (N_20636,N_19497,N_18848);
xor U20637 (N_20637,N_19044,N_19557);
nor U20638 (N_20638,N_19320,N_19243);
nor U20639 (N_20639,N_18834,N_19900);
xor U20640 (N_20640,N_19917,N_18822);
and U20641 (N_20641,N_19772,N_19323);
or U20642 (N_20642,N_19474,N_19160);
or U20643 (N_20643,N_19548,N_19487);
nand U20644 (N_20644,N_19866,N_19689);
or U20645 (N_20645,N_19985,N_19659);
xor U20646 (N_20646,N_19904,N_19237);
nand U20647 (N_20647,N_19281,N_19831);
and U20648 (N_20648,N_19982,N_19000);
xor U20649 (N_20649,N_18855,N_19560);
nor U20650 (N_20650,N_19302,N_19530);
nor U20651 (N_20651,N_19565,N_19240);
or U20652 (N_20652,N_19245,N_19493);
or U20653 (N_20653,N_19777,N_19342);
or U20654 (N_20654,N_19409,N_18955);
and U20655 (N_20655,N_19275,N_19192);
nor U20656 (N_20656,N_19205,N_18794);
nor U20657 (N_20657,N_19203,N_19630);
nor U20658 (N_20658,N_19677,N_19011);
nor U20659 (N_20659,N_19265,N_19255);
and U20660 (N_20660,N_19761,N_19188);
xor U20661 (N_20661,N_19718,N_19934);
nand U20662 (N_20662,N_19923,N_19102);
nor U20663 (N_20663,N_19890,N_19948);
xor U20664 (N_20664,N_19236,N_19446);
and U20665 (N_20665,N_19580,N_18910);
and U20666 (N_20666,N_19603,N_19775);
xnor U20667 (N_20667,N_19104,N_18845);
and U20668 (N_20668,N_19588,N_19755);
or U20669 (N_20669,N_19537,N_19466);
nand U20670 (N_20670,N_18784,N_19247);
xnor U20671 (N_20671,N_18792,N_18970);
xor U20672 (N_20672,N_19264,N_19166);
nor U20673 (N_20673,N_19082,N_19838);
xnor U20674 (N_20674,N_19983,N_19648);
nand U20675 (N_20675,N_18794,N_18861);
or U20676 (N_20676,N_19266,N_18926);
nor U20677 (N_20677,N_19608,N_18994);
and U20678 (N_20678,N_18876,N_18936);
or U20679 (N_20679,N_18771,N_19130);
nor U20680 (N_20680,N_19619,N_18872);
and U20681 (N_20681,N_19309,N_19236);
and U20682 (N_20682,N_19722,N_19595);
and U20683 (N_20683,N_19825,N_18980);
nand U20684 (N_20684,N_19711,N_18990);
xnor U20685 (N_20685,N_19473,N_19322);
nor U20686 (N_20686,N_19775,N_19698);
and U20687 (N_20687,N_19709,N_19188);
or U20688 (N_20688,N_19389,N_19212);
nand U20689 (N_20689,N_19003,N_19174);
xnor U20690 (N_20690,N_19374,N_19367);
and U20691 (N_20691,N_18923,N_19706);
or U20692 (N_20692,N_19561,N_19270);
or U20693 (N_20693,N_18889,N_19208);
nand U20694 (N_20694,N_19406,N_19333);
or U20695 (N_20695,N_19518,N_19371);
nor U20696 (N_20696,N_19052,N_18865);
and U20697 (N_20697,N_19495,N_19293);
or U20698 (N_20698,N_19509,N_19882);
or U20699 (N_20699,N_19976,N_19624);
or U20700 (N_20700,N_19310,N_19934);
nor U20701 (N_20701,N_19978,N_19208);
nor U20702 (N_20702,N_18878,N_19845);
nor U20703 (N_20703,N_19642,N_18783);
xor U20704 (N_20704,N_19311,N_19883);
nor U20705 (N_20705,N_19050,N_18936);
and U20706 (N_20706,N_19555,N_18784);
or U20707 (N_20707,N_18897,N_19096);
or U20708 (N_20708,N_19009,N_19397);
nand U20709 (N_20709,N_19902,N_19224);
xor U20710 (N_20710,N_19486,N_19932);
or U20711 (N_20711,N_19878,N_19686);
nand U20712 (N_20712,N_19720,N_19067);
or U20713 (N_20713,N_19089,N_19716);
nand U20714 (N_20714,N_19911,N_19907);
and U20715 (N_20715,N_19250,N_19426);
or U20716 (N_20716,N_19125,N_19832);
nor U20717 (N_20717,N_19158,N_19260);
and U20718 (N_20718,N_18993,N_19660);
nor U20719 (N_20719,N_19600,N_19684);
or U20720 (N_20720,N_19606,N_19034);
and U20721 (N_20721,N_19935,N_19397);
and U20722 (N_20722,N_19679,N_19166);
nand U20723 (N_20723,N_19307,N_19965);
and U20724 (N_20724,N_19744,N_18839);
xor U20725 (N_20725,N_18791,N_19243);
and U20726 (N_20726,N_18994,N_19010);
and U20727 (N_20727,N_19868,N_19946);
or U20728 (N_20728,N_18966,N_19037);
nand U20729 (N_20729,N_18928,N_19651);
or U20730 (N_20730,N_19439,N_19885);
nand U20731 (N_20731,N_18988,N_19869);
or U20732 (N_20732,N_19726,N_19668);
nor U20733 (N_20733,N_19373,N_19219);
and U20734 (N_20734,N_19883,N_19030);
xnor U20735 (N_20735,N_19846,N_19981);
nor U20736 (N_20736,N_19137,N_19540);
nor U20737 (N_20737,N_18837,N_18898);
nand U20738 (N_20738,N_19807,N_19099);
nand U20739 (N_20739,N_19191,N_18901);
or U20740 (N_20740,N_19802,N_19984);
or U20741 (N_20741,N_19516,N_19857);
nand U20742 (N_20742,N_19587,N_18997);
nand U20743 (N_20743,N_18853,N_19155);
nand U20744 (N_20744,N_19929,N_19726);
nor U20745 (N_20745,N_18763,N_19909);
and U20746 (N_20746,N_19867,N_18820);
and U20747 (N_20747,N_19137,N_18887);
and U20748 (N_20748,N_18754,N_19559);
nand U20749 (N_20749,N_19563,N_18963);
nand U20750 (N_20750,N_19840,N_18947);
and U20751 (N_20751,N_19955,N_19276);
xor U20752 (N_20752,N_19957,N_18913);
and U20753 (N_20753,N_19696,N_19816);
nor U20754 (N_20754,N_19720,N_19097);
and U20755 (N_20755,N_19953,N_19884);
nand U20756 (N_20756,N_19859,N_19944);
and U20757 (N_20757,N_18978,N_19800);
and U20758 (N_20758,N_19712,N_19412);
nand U20759 (N_20759,N_19699,N_19810);
or U20760 (N_20760,N_19520,N_19870);
nor U20761 (N_20761,N_19300,N_19261);
xnor U20762 (N_20762,N_18935,N_19122);
and U20763 (N_20763,N_19330,N_19668);
or U20764 (N_20764,N_19086,N_19876);
nor U20765 (N_20765,N_19962,N_19246);
nand U20766 (N_20766,N_19586,N_19487);
nand U20767 (N_20767,N_19163,N_19882);
xor U20768 (N_20768,N_19993,N_18813);
nor U20769 (N_20769,N_19820,N_19929);
nor U20770 (N_20770,N_18848,N_18944);
or U20771 (N_20771,N_19039,N_19651);
xor U20772 (N_20772,N_19870,N_18884);
nor U20773 (N_20773,N_19811,N_18852);
or U20774 (N_20774,N_19508,N_19864);
and U20775 (N_20775,N_19554,N_19782);
and U20776 (N_20776,N_18930,N_19138);
nor U20777 (N_20777,N_19548,N_19903);
nor U20778 (N_20778,N_19968,N_18906);
nand U20779 (N_20779,N_19609,N_18762);
and U20780 (N_20780,N_19730,N_19513);
nor U20781 (N_20781,N_19636,N_19498);
nor U20782 (N_20782,N_19403,N_19165);
nor U20783 (N_20783,N_19392,N_19865);
nand U20784 (N_20784,N_19437,N_19898);
xor U20785 (N_20785,N_19089,N_19790);
and U20786 (N_20786,N_19407,N_19624);
nand U20787 (N_20787,N_19499,N_19376);
xor U20788 (N_20788,N_19164,N_19683);
or U20789 (N_20789,N_19953,N_19400);
and U20790 (N_20790,N_19892,N_19778);
xor U20791 (N_20791,N_18969,N_19091);
nor U20792 (N_20792,N_18865,N_19709);
nand U20793 (N_20793,N_19912,N_18927);
xnor U20794 (N_20794,N_19831,N_19338);
nand U20795 (N_20795,N_19816,N_18864);
and U20796 (N_20796,N_19965,N_19538);
nor U20797 (N_20797,N_19337,N_19684);
nor U20798 (N_20798,N_19647,N_19193);
nor U20799 (N_20799,N_19909,N_19031);
and U20800 (N_20800,N_19457,N_18774);
nor U20801 (N_20801,N_19259,N_19508);
nand U20802 (N_20802,N_19468,N_19909);
nor U20803 (N_20803,N_19624,N_19439);
and U20804 (N_20804,N_18810,N_19058);
or U20805 (N_20805,N_18836,N_18943);
nor U20806 (N_20806,N_19076,N_19026);
or U20807 (N_20807,N_19241,N_19008);
nor U20808 (N_20808,N_19344,N_19258);
xor U20809 (N_20809,N_18988,N_18894);
nand U20810 (N_20810,N_18770,N_19292);
nand U20811 (N_20811,N_19237,N_19698);
and U20812 (N_20812,N_19391,N_19888);
and U20813 (N_20813,N_18848,N_19426);
xor U20814 (N_20814,N_19271,N_19173);
nor U20815 (N_20815,N_19230,N_19840);
or U20816 (N_20816,N_19846,N_19228);
nand U20817 (N_20817,N_19304,N_19913);
nand U20818 (N_20818,N_19924,N_19897);
and U20819 (N_20819,N_19500,N_18764);
nand U20820 (N_20820,N_19520,N_19197);
or U20821 (N_20821,N_19620,N_19398);
or U20822 (N_20822,N_19581,N_19777);
or U20823 (N_20823,N_19701,N_19851);
nor U20824 (N_20824,N_19135,N_19659);
or U20825 (N_20825,N_19887,N_19536);
nor U20826 (N_20826,N_19867,N_18885);
nor U20827 (N_20827,N_19343,N_19577);
nand U20828 (N_20828,N_19413,N_19719);
or U20829 (N_20829,N_19999,N_19294);
nand U20830 (N_20830,N_19229,N_19226);
nor U20831 (N_20831,N_19442,N_19950);
nor U20832 (N_20832,N_19744,N_19839);
nand U20833 (N_20833,N_19269,N_19950);
and U20834 (N_20834,N_18947,N_18839);
nand U20835 (N_20835,N_18949,N_19759);
and U20836 (N_20836,N_18958,N_18778);
and U20837 (N_20837,N_19895,N_19099);
or U20838 (N_20838,N_19087,N_18931);
or U20839 (N_20839,N_19415,N_19057);
nor U20840 (N_20840,N_19129,N_18792);
and U20841 (N_20841,N_18963,N_19836);
nand U20842 (N_20842,N_19475,N_19538);
nand U20843 (N_20843,N_18947,N_19374);
xnor U20844 (N_20844,N_19730,N_19992);
xnor U20845 (N_20845,N_19527,N_18912);
and U20846 (N_20846,N_18927,N_19526);
nand U20847 (N_20847,N_19364,N_19147);
nand U20848 (N_20848,N_19030,N_19667);
nand U20849 (N_20849,N_19845,N_18885);
or U20850 (N_20850,N_19439,N_19293);
nor U20851 (N_20851,N_18799,N_19409);
and U20852 (N_20852,N_19176,N_18863);
nand U20853 (N_20853,N_19734,N_18908);
and U20854 (N_20854,N_19457,N_19776);
and U20855 (N_20855,N_19546,N_19938);
nand U20856 (N_20856,N_19922,N_18862);
and U20857 (N_20857,N_19491,N_19411);
nor U20858 (N_20858,N_19527,N_19804);
or U20859 (N_20859,N_19970,N_19136);
or U20860 (N_20860,N_19597,N_19797);
and U20861 (N_20861,N_19515,N_19166);
xnor U20862 (N_20862,N_19725,N_19115);
and U20863 (N_20863,N_19606,N_19288);
nor U20864 (N_20864,N_19126,N_18798);
xnor U20865 (N_20865,N_19148,N_19577);
nor U20866 (N_20866,N_18985,N_18769);
nor U20867 (N_20867,N_19684,N_19699);
nor U20868 (N_20868,N_19023,N_19215);
and U20869 (N_20869,N_19307,N_19420);
or U20870 (N_20870,N_18858,N_19566);
nand U20871 (N_20871,N_19383,N_19087);
and U20872 (N_20872,N_19840,N_18876);
nand U20873 (N_20873,N_19092,N_19713);
xor U20874 (N_20874,N_19201,N_18963);
or U20875 (N_20875,N_18841,N_18904);
or U20876 (N_20876,N_19260,N_19399);
nor U20877 (N_20877,N_19291,N_18781);
nand U20878 (N_20878,N_19349,N_19633);
xnor U20879 (N_20879,N_19242,N_19003);
and U20880 (N_20880,N_19852,N_19515);
xnor U20881 (N_20881,N_18827,N_19594);
xor U20882 (N_20882,N_19825,N_19454);
or U20883 (N_20883,N_18972,N_19570);
or U20884 (N_20884,N_19269,N_19487);
or U20885 (N_20885,N_19606,N_18975);
or U20886 (N_20886,N_19182,N_19327);
or U20887 (N_20887,N_19982,N_18810);
and U20888 (N_20888,N_19306,N_18779);
nand U20889 (N_20889,N_18964,N_18895);
or U20890 (N_20890,N_19297,N_19700);
and U20891 (N_20891,N_19471,N_19314);
or U20892 (N_20892,N_19595,N_19128);
nand U20893 (N_20893,N_18941,N_19314);
and U20894 (N_20894,N_19263,N_19130);
nor U20895 (N_20895,N_19900,N_18866);
or U20896 (N_20896,N_18885,N_19822);
nand U20897 (N_20897,N_19221,N_19520);
nor U20898 (N_20898,N_19839,N_18859);
nand U20899 (N_20899,N_19276,N_19374);
and U20900 (N_20900,N_19884,N_19593);
nor U20901 (N_20901,N_19289,N_19960);
nor U20902 (N_20902,N_19648,N_19600);
and U20903 (N_20903,N_19432,N_19924);
xor U20904 (N_20904,N_19292,N_18875);
or U20905 (N_20905,N_18958,N_19665);
and U20906 (N_20906,N_19543,N_19681);
xnor U20907 (N_20907,N_19958,N_19202);
nor U20908 (N_20908,N_19877,N_19719);
nand U20909 (N_20909,N_19040,N_19166);
xnor U20910 (N_20910,N_18847,N_19784);
xor U20911 (N_20911,N_19173,N_19494);
and U20912 (N_20912,N_19599,N_19561);
nand U20913 (N_20913,N_19199,N_19638);
and U20914 (N_20914,N_18801,N_19176);
or U20915 (N_20915,N_18961,N_18906);
nand U20916 (N_20916,N_18766,N_18870);
or U20917 (N_20917,N_19440,N_19813);
nor U20918 (N_20918,N_19868,N_19094);
nor U20919 (N_20919,N_19896,N_19658);
xor U20920 (N_20920,N_19272,N_19055);
and U20921 (N_20921,N_19980,N_19713);
and U20922 (N_20922,N_19303,N_19919);
xnor U20923 (N_20923,N_19112,N_19093);
and U20924 (N_20924,N_19491,N_19546);
nor U20925 (N_20925,N_19333,N_19773);
xnor U20926 (N_20926,N_18960,N_19584);
or U20927 (N_20927,N_19305,N_19473);
nand U20928 (N_20928,N_19939,N_19993);
and U20929 (N_20929,N_19499,N_19323);
and U20930 (N_20930,N_18917,N_19871);
nor U20931 (N_20931,N_18833,N_19372);
or U20932 (N_20932,N_19160,N_19593);
and U20933 (N_20933,N_19691,N_18827);
nor U20934 (N_20934,N_19314,N_19896);
or U20935 (N_20935,N_19481,N_19134);
or U20936 (N_20936,N_19489,N_19607);
nand U20937 (N_20937,N_19433,N_19280);
and U20938 (N_20938,N_19082,N_19458);
or U20939 (N_20939,N_19686,N_19690);
xnor U20940 (N_20940,N_19211,N_19693);
or U20941 (N_20941,N_18848,N_19085);
nand U20942 (N_20942,N_19293,N_19237);
xor U20943 (N_20943,N_19484,N_18903);
and U20944 (N_20944,N_19425,N_19454);
or U20945 (N_20945,N_19755,N_19809);
xnor U20946 (N_20946,N_19553,N_19791);
nor U20947 (N_20947,N_18944,N_19128);
or U20948 (N_20948,N_19986,N_19995);
or U20949 (N_20949,N_19171,N_19488);
or U20950 (N_20950,N_19992,N_19426);
and U20951 (N_20951,N_19507,N_19908);
nand U20952 (N_20952,N_19352,N_19169);
xnor U20953 (N_20953,N_18780,N_19905);
xnor U20954 (N_20954,N_19646,N_19075);
xnor U20955 (N_20955,N_18976,N_19842);
xnor U20956 (N_20956,N_19028,N_19298);
or U20957 (N_20957,N_19993,N_19944);
xor U20958 (N_20958,N_18869,N_18823);
and U20959 (N_20959,N_19001,N_19192);
nand U20960 (N_20960,N_19121,N_19653);
nor U20961 (N_20961,N_19088,N_19356);
nand U20962 (N_20962,N_19406,N_19667);
or U20963 (N_20963,N_19149,N_19512);
or U20964 (N_20964,N_19313,N_19088);
and U20965 (N_20965,N_19787,N_19158);
and U20966 (N_20966,N_19645,N_19614);
or U20967 (N_20967,N_19031,N_19422);
nor U20968 (N_20968,N_19725,N_19975);
and U20969 (N_20969,N_19957,N_19014);
xor U20970 (N_20970,N_19886,N_19577);
or U20971 (N_20971,N_19044,N_18805);
and U20972 (N_20972,N_19598,N_19071);
xor U20973 (N_20973,N_19832,N_19628);
nand U20974 (N_20974,N_19027,N_19566);
nand U20975 (N_20975,N_18958,N_19675);
xnor U20976 (N_20976,N_19825,N_19112);
and U20977 (N_20977,N_19969,N_19461);
nand U20978 (N_20978,N_18895,N_19833);
or U20979 (N_20979,N_19623,N_19559);
or U20980 (N_20980,N_19095,N_19272);
and U20981 (N_20981,N_18793,N_18994);
nand U20982 (N_20982,N_18767,N_19273);
or U20983 (N_20983,N_19185,N_19288);
nor U20984 (N_20984,N_19013,N_19204);
nand U20985 (N_20985,N_19433,N_19906);
or U20986 (N_20986,N_19218,N_19848);
and U20987 (N_20987,N_19126,N_18754);
or U20988 (N_20988,N_18903,N_19380);
nand U20989 (N_20989,N_18954,N_19580);
or U20990 (N_20990,N_18768,N_18921);
nand U20991 (N_20991,N_19758,N_19682);
nor U20992 (N_20992,N_19343,N_19536);
or U20993 (N_20993,N_19071,N_19804);
nor U20994 (N_20994,N_19478,N_18831);
nand U20995 (N_20995,N_18766,N_19484);
and U20996 (N_20996,N_19937,N_19738);
or U20997 (N_20997,N_18881,N_19855);
nand U20998 (N_20998,N_19349,N_19545);
xnor U20999 (N_20999,N_19172,N_19332);
or U21000 (N_21000,N_18802,N_18978);
and U21001 (N_21001,N_19376,N_19519);
xor U21002 (N_21002,N_18823,N_19261);
xor U21003 (N_21003,N_19778,N_18885);
nand U21004 (N_21004,N_18810,N_19739);
nand U21005 (N_21005,N_18962,N_19730);
or U21006 (N_21006,N_19271,N_19703);
nor U21007 (N_21007,N_19941,N_19438);
and U21008 (N_21008,N_19235,N_19711);
xnor U21009 (N_21009,N_18980,N_19282);
xor U21010 (N_21010,N_19418,N_19180);
nand U21011 (N_21011,N_19962,N_18948);
or U21012 (N_21012,N_19278,N_18862);
and U21013 (N_21013,N_18812,N_19955);
and U21014 (N_21014,N_19749,N_19618);
nand U21015 (N_21015,N_19768,N_19479);
xor U21016 (N_21016,N_18798,N_19405);
or U21017 (N_21017,N_19407,N_19926);
and U21018 (N_21018,N_19224,N_18826);
nor U21019 (N_21019,N_19312,N_19172);
nor U21020 (N_21020,N_19181,N_19148);
xor U21021 (N_21021,N_19879,N_19998);
or U21022 (N_21022,N_19895,N_19644);
or U21023 (N_21023,N_18977,N_19013);
and U21024 (N_21024,N_19136,N_19500);
xor U21025 (N_21025,N_19837,N_19618);
nand U21026 (N_21026,N_19583,N_19355);
xnor U21027 (N_21027,N_19273,N_19060);
xnor U21028 (N_21028,N_19282,N_19325);
nor U21029 (N_21029,N_19600,N_19415);
and U21030 (N_21030,N_19882,N_19450);
nor U21031 (N_21031,N_18814,N_18817);
and U21032 (N_21032,N_19572,N_19501);
nand U21033 (N_21033,N_19982,N_18797);
nand U21034 (N_21034,N_19538,N_18967);
xor U21035 (N_21035,N_19337,N_18808);
nand U21036 (N_21036,N_18835,N_19686);
nor U21037 (N_21037,N_19077,N_19037);
or U21038 (N_21038,N_18842,N_19031);
xor U21039 (N_21039,N_18953,N_19466);
xnor U21040 (N_21040,N_19554,N_19200);
nor U21041 (N_21041,N_19220,N_19614);
or U21042 (N_21042,N_19008,N_19574);
nand U21043 (N_21043,N_19507,N_19102);
xor U21044 (N_21044,N_18977,N_19686);
xor U21045 (N_21045,N_19811,N_19821);
xnor U21046 (N_21046,N_19485,N_19865);
and U21047 (N_21047,N_19309,N_19034);
and U21048 (N_21048,N_19492,N_18794);
or U21049 (N_21049,N_19041,N_19698);
xnor U21050 (N_21050,N_19001,N_19422);
and U21051 (N_21051,N_19349,N_19606);
or U21052 (N_21052,N_19339,N_19184);
xnor U21053 (N_21053,N_19674,N_18956);
nand U21054 (N_21054,N_19016,N_19509);
xnor U21055 (N_21055,N_18862,N_19820);
and U21056 (N_21056,N_18968,N_19597);
nand U21057 (N_21057,N_19170,N_19970);
xnor U21058 (N_21058,N_18879,N_19812);
or U21059 (N_21059,N_19342,N_19097);
or U21060 (N_21060,N_19032,N_19919);
nor U21061 (N_21061,N_19708,N_19660);
and U21062 (N_21062,N_19944,N_18750);
or U21063 (N_21063,N_19140,N_19549);
and U21064 (N_21064,N_19900,N_19075);
xor U21065 (N_21065,N_19270,N_19235);
xnor U21066 (N_21066,N_19429,N_19667);
xnor U21067 (N_21067,N_19556,N_19640);
xnor U21068 (N_21068,N_19369,N_19942);
nor U21069 (N_21069,N_18811,N_18904);
xnor U21070 (N_21070,N_19526,N_19888);
xnor U21071 (N_21071,N_19197,N_19935);
and U21072 (N_21072,N_18765,N_19973);
or U21073 (N_21073,N_19162,N_19808);
nand U21074 (N_21074,N_19798,N_19527);
xor U21075 (N_21075,N_18926,N_19109);
or U21076 (N_21076,N_18815,N_19885);
nor U21077 (N_21077,N_19424,N_19436);
nor U21078 (N_21078,N_19187,N_19792);
or U21079 (N_21079,N_19217,N_18752);
nand U21080 (N_21080,N_19480,N_19009);
xor U21081 (N_21081,N_18803,N_19969);
nand U21082 (N_21082,N_19765,N_19668);
nand U21083 (N_21083,N_19490,N_18850);
nor U21084 (N_21084,N_19777,N_19055);
nor U21085 (N_21085,N_19214,N_19077);
nor U21086 (N_21086,N_19892,N_19805);
nand U21087 (N_21087,N_18890,N_19694);
nand U21088 (N_21088,N_19383,N_19576);
and U21089 (N_21089,N_19757,N_19014);
nand U21090 (N_21090,N_19711,N_19458);
or U21091 (N_21091,N_19457,N_19439);
nand U21092 (N_21092,N_19706,N_18852);
or U21093 (N_21093,N_19252,N_19824);
xnor U21094 (N_21094,N_19287,N_19298);
or U21095 (N_21095,N_19726,N_19742);
or U21096 (N_21096,N_19671,N_19979);
nor U21097 (N_21097,N_19545,N_18839);
xor U21098 (N_21098,N_19008,N_18927);
and U21099 (N_21099,N_19688,N_19185);
nand U21100 (N_21100,N_19183,N_19736);
xnor U21101 (N_21101,N_19095,N_19711);
nand U21102 (N_21102,N_19533,N_19555);
or U21103 (N_21103,N_19258,N_19716);
nand U21104 (N_21104,N_19188,N_19333);
or U21105 (N_21105,N_19672,N_19764);
nor U21106 (N_21106,N_19772,N_19960);
or U21107 (N_21107,N_19883,N_19949);
and U21108 (N_21108,N_19802,N_19209);
nand U21109 (N_21109,N_19324,N_19180);
xnor U21110 (N_21110,N_19595,N_18958);
or U21111 (N_21111,N_19171,N_19234);
nand U21112 (N_21112,N_19176,N_19912);
and U21113 (N_21113,N_19876,N_19373);
or U21114 (N_21114,N_19142,N_19549);
or U21115 (N_21115,N_19818,N_18984);
nor U21116 (N_21116,N_19446,N_19603);
or U21117 (N_21117,N_19685,N_18951);
and U21118 (N_21118,N_19773,N_18915);
xor U21119 (N_21119,N_19142,N_18890);
nand U21120 (N_21120,N_19220,N_19435);
nand U21121 (N_21121,N_19925,N_19643);
nor U21122 (N_21122,N_18959,N_19429);
xor U21123 (N_21123,N_19544,N_19008);
nor U21124 (N_21124,N_18996,N_19637);
and U21125 (N_21125,N_19544,N_18929);
and U21126 (N_21126,N_19498,N_19875);
nand U21127 (N_21127,N_19187,N_19834);
xor U21128 (N_21128,N_19485,N_19848);
xnor U21129 (N_21129,N_19262,N_19092);
or U21130 (N_21130,N_19954,N_18959);
nor U21131 (N_21131,N_19076,N_19773);
or U21132 (N_21132,N_19474,N_19751);
and U21133 (N_21133,N_19457,N_19236);
or U21134 (N_21134,N_19039,N_19256);
xor U21135 (N_21135,N_19460,N_19002);
nand U21136 (N_21136,N_19545,N_19705);
and U21137 (N_21137,N_19004,N_19383);
xor U21138 (N_21138,N_19804,N_18867);
nand U21139 (N_21139,N_19736,N_19125);
nor U21140 (N_21140,N_19411,N_19533);
nand U21141 (N_21141,N_18937,N_19639);
xnor U21142 (N_21142,N_19007,N_19163);
xor U21143 (N_21143,N_19850,N_19653);
nor U21144 (N_21144,N_19589,N_18886);
xnor U21145 (N_21145,N_19512,N_19974);
or U21146 (N_21146,N_19517,N_19879);
nand U21147 (N_21147,N_19662,N_18989);
or U21148 (N_21148,N_19022,N_18851);
nand U21149 (N_21149,N_19530,N_19985);
nand U21150 (N_21150,N_19527,N_19128);
and U21151 (N_21151,N_19463,N_19723);
or U21152 (N_21152,N_19704,N_19523);
nand U21153 (N_21153,N_19387,N_19189);
or U21154 (N_21154,N_19017,N_19606);
nand U21155 (N_21155,N_19406,N_19707);
nor U21156 (N_21156,N_18772,N_19698);
nor U21157 (N_21157,N_19375,N_19661);
nor U21158 (N_21158,N_19612,N_19779);
and U21159 (N_21159,N_19813,N_18824);
nand U21160 (N_21160,N_19525,N_19488);
and U21161 (N_21161,N_19232,N_19646);
xor U21162 (N_21162,N_19877,N_19620);
nand U21163 (N_21163,N_19721,N_19892);
nand U21164 (N_21164,N_19063,N_19910);
xnor U21165 (N_21165,N_18913,N_19084);
xnor U21166 (N_21166,N_18948,N_19827);
xnor U21167 (N_21167,N_18851,N_19928);
or U21168 (N_21168,N_19799,N_19317);
nor U21169 (N_21169,N_19615,N_19430);
xnor U21170 (N_21170,N_18909,N_19125);
xnor U21171 (N_21171,N_19471,N_19201);
or U21172 (N_21172,N_19948,N_19611);
and U21173 (N_21173,N_19757,N_19675);
or U21174 (N_21174,N_19163,N_19490);
nor U21175 (N_21175,N_19802,N_19054);
nor U21176 (N_21176,N_19594,N_19566);
and U21177 (N_21177,N_18961,N_19875);
xor U21178 (N_21178,N_19478,N_19807);
or U21179 (N_21179,N_19006,N_19246);
or U21180 (N_21180,N_18764,N_19838);
nand U21181 (N_21181,N_19132,N_18795);
and U21182 (N_21182,N_19740,N_19759);
xor U21183 (N_21183,N_18879,N_19155);
xnor U21184 (N_21184,N_18807,N_18819);
nand U21185 (N_21185,N_19165,N_18935);
nor U21186 (N_21186,N_19093,N_19403);
nor U21187 (N_21187,N_19220,N_19584);
xor U21188 (N_21188,N_19803,N_18928);
xor U21189 (N_21189,N_19741,N_19674);
xnor U21190 (N_21190,N_19380,N_18946);
nor U21191 (N_21191,N_19444,N_18998);
xnor U21192 (N_21192,N_18781,N_19352);
and U21193 (N_21193,N_19627,N_18965);
or U21194 (N_21194,N_18801,N_19006);
nor U21195 (N_21195,N_19902,N_19065);
nor U21196 (N_21196,N_18774,N_19554);
nand U21197 (N_21197,N_19439,N_19764);
and U21198 (N_21198,N_19943,N_19156);
and U21199 (N_21199,N_18760,N_18828);
nor U21200 (N_21200,N_19233,N_19493);
nand U21201 (N_21201,N_19897,N_18951);
nand U21202 (N_21202,N_19852,N_19355);
nand U21203 (N_21203,N_19420,N_18871);
xnor U21204 (N_21204,N_19998,N_19880);
nor U21205 (N_21205,N_19705,N_19782);
and U21206 (N_21206,N_19030,N_19972);
or U21207 (N_21207,N_19008,N_19887);
xnor U21208 (N_21208,N_19993,N_19900);
nand U21209 (N_21209,N_19706,N_19697);
and U21210 (N_21210,N_19410,N_18966);
xor U21211 (N_21211,N_19854,N_19669);
or U21212 (N_21212,N_19067,N_18865);
and U21213 (N_21213,N_19017,N_19784);
and U21214 (N_21214,N_19415,N_19984);
or U21215 (N_21215,N_19362,N_19125);
nor U21216 (N_21216,N_19782,N_19891);
and U21217 (N_21217,N_19983,N_19763);
xor U21218 (N_21218,N_19902,N_19814);
and U21219 (N_21219,N_18780,N_18771);
xor U21220 (N_21220,N_19433,N_19625);
and U21221 (N_21221,N_19841,N_19472);
xor U21222 (N_21222,N_19901,N_19872);
or U21223 (N_21223,N_19473,N_19818);
and U21224 (N_21224,N_19671,N_19247);
and U21225 (N_21225,N_19136,N_18962);
and U21226 (N_21226,N_19102,N_18937);
or U21227 (N_21227,N_19221,N_18929);
and U21228 (N_21228,N_19868,N_19546);
and U21229 (N_21229,N_19185,N_19740);
and U21230 (N_21230,N_18903,N_19259);
or U21231 (N_21231,N_19568,N_19839);
or U21232 (N_21232,N_19992,N_19088);
and U21233 (N_21233,N_18961,N_19074);
nor U21234 (N_21234,N_19197,N_19998);
or U21235 (N_21235,N_19017,N_19393);
xor U21236 (N_21236,N_19054,N_18977);
xnor U21237 (N_21237,N_19628,N_19192);
or U21238 (N_21238,N_19499,N_18916);
nand U21239 (N_21239,N_19220,N_19546);
xor U21240 (N_21240,N_19924,N_19581);
or U21241 (N_21241,N_19488,N_19730);
or U21242 (N_21242,N_19251,N_18915);
or U21243 (N_21243,N_19882,N_19402);
or U21244 (N_21244,N_18761,N_19436);
nor U21245 (N_21245,N_19760,N_19277);
or U21246 (N_21246,N_18937,N_18903);
xnor U21247 (N_21247,N_18868,N_18906);
or U21248 (N_21248,N_19203,N_19695);
nor U21249 (N_21249,N_19932,N_19651);
and U21250 (N_21250,N_21092,N_20537);
nand U21251 (N_21251,N_20355,N_21008);
or U21252 (N_21252,N_21203,N_21167);
xnor U21253 (N_21253,N_20288,N_20322);
nor U21254 (N_21254,N_20492,N_20824);
or U21255 (N_21255,N_20217,N_20014);
xnor U21256 (N_21256,N_20941,N_21122);
nor U21257 (N_21257,N_21088,N_21082);
xor U21258 (N_21258,N_20967,N_20857);
nor U21259 (N_21259,N_20135,N_20045);
nand U21260 (N_21260,N_20575,N_21141);
or U21261 (N_21261,N_20481,N_20635);
nor U21262 (N_21262,N_20034,N_20546);
nor U21263 (N_21263,N_20345,N_20885);
nand U21264 (N_21264,N_20634,N_20675);
xor U21265 (N_21265,N_20037,N_21155);
nand U21266 (N_21266,N_21146,N_20376);
nor U21267 (N_21267,N_21103,N_20658);
or U21268 (N_21268,N_20505,N_20980);
xor U21269 (N_21269,N_20465,N_20101);
nand U21270 (N_21270,N_21044,N_21175);
and U21271 (N_21271,N_20300,N_20805);
nor U21272 (N_21272,N_20527,N_21192);
or U21273 (N_21273,N_20147,N_20951);
xor U21274 (N_21274,N_20704,N_20396);
nand U21275 (N_21275,N_21202,N_20640);
nor U21276 (N_21276,N_20990,N_20063);
or U21277 (N_21277,N_20336,N_20818);
nor U21278 (N_21278,N_20298,N_20861);
nand U21279 (N_21279,N_20406,N_20287);
nor U21280 (N_21280,N_20269,N_20359);
nand U21281 (N_21281,N_20272,N_20447);
or U21282 (N_21282,N_20853,N_20562);
and U21283 (N_21283,N_20715,N_21235);
nor U21284 (N_21284,N_20612,N_21228);
nand U21285 (N_21285,N_20840,N_20219);
xor U21286 (N_21286,N_20190,N_20632);
nor U21287 (N_21287,N_20954,N_21150);
and U21288 (N_21288,N_20314,N_20566);
or U21289 (N_21289,N_20491,N_20810);
xor U21290 (N_21290,N_20551,N_20468);
nor U21291 (N_21291,N_20787,N_20904);
or U21292 (N_21292,N_20381,N_20471);
nor U21293 (N_21293,N_21210,N_20567);
nand U21294 (N_21294,N_20455,N_21191);
or U21295 (N_21295,N_20297,N_20850);
nor U21296 (N_21296,N_20835,N_20080);
xor U21297 (N_21297,N_20870,N_20246);
and U21298 (N_21298,N_20942,N_20498);
or U21299 (N_21299,N_20457,N_20800);
or U21300 (N_21300,N_21112,N_20846);
nand U21301 (N_21301,N_20115,N_20531);
nand U21302 (N_21302,N_21027,N_20369);
xnor U21303 (N_21303,N_20563,N_20930);
nor U21304 (N_21304,N_20175,N_21095);
and U21305 (N_21305,N_20596,N_20018);
xnor U21306 (N_21306,N_20698,N_20616);
or U21307 (N_21307,N_20024,N_20153);
nand U21308 (N_21308,N_21186,N_20451);
nand U21309 (N_21309,N_20561,N_20858);
nand U21310 (N_21310,N_20865,N_20433);
xor U21311 (N_21311,N_21035,N_20149);
or U21312 (N_21312,N_20871,N_20874);
and U21313 (N_21313,N_20162,N_20366);
xor U21314 (N_21314,N_20020,N_21166);
nor U21315 (N_21315,N_20694,N_20050);
xor U21316 (N_21316,N_20347,N_20273);
or U21317 (N_21317,N_20814,N_21230);
nand U21318 (N_21318,N_20332,N_20876);
and U21319 (N_21319,N_20720,N_20072);
and U21320 (N_21320,N_20279,N_20485);
or U21321 (N_21321,N_20318,N_20048);
nand U21322 (N_21322,N_20660,N_20134);
or U21323 (N_21323,N_21090,N_20242);
or U21324 (N_21324,N_21098,N_21173);
and U21325 (N_21325,N_21179,N_20388);
or U21326 (N_21326,N_20986,N_20483);
nand U21327 (N_21327,N_20431,N_20801);
nor U21328 (N_21328,N_20644,N_20588);
nor U21329 (N_21329,N_20856,N_20822);
xnor U21330 (N_21330,N_20906,N_20121);
or U21331 (N_21331,N_21214,N_21057);
or U21332 (N_21332,N_20619,N_20569);
nand U21333 (N_21333,N_20157,N_21028);
or U21334 (N_21334,N_20864,N_20985);
and U21335 (N_21335,N_20005,N_20570);
or U21336 (N_21336,N_20795,N_20540);
or U21337 (N_21337,N_20979,N_20205);
or U21338 (N_21338,N_20262,N_20617);
or U21339 (N_21339,N_21133,N_21209);
xor U21340 (N_21340,N_20953,N_20069);
or U21341 (N_21341,N_20912,N_20486);
or U21342 (N_21342,N_21212,N_20118);
or U21343 (N_21343,N_20823,N_20257);
and U21344 (N_21344,N_20449,N_20519);
nor U21345 (N_21345,N_20712,N_20978);
and U21346 (N_21346,N_20664,N_21229);
nand U21347 (N_21347,N_21128,N_20316);
nand U21348 (N_21348,N_20681,N_20143);
nor U21349 (N_21349,N_20295,N_20933);
nand U21350 (N_21350,N_20815,N_20197);
or U21351 (N_21351,N_20525,N_20998);
and U21352 (N_21352,N_21196,N_20282);
and U21353 (N_21353,N_21104,N_20999);
nor U21354 (N_21354,N_21094,N_21237);
nor U21355 (N_21355,N_20132,N_21165);
nor U21356 (N_21356,N_20091,N_21107);
nor U21357 (N_21357,N_20384,N_20429);
xnor U21358 (N_21358,N_20290,N_20541);
xor U21359 (N_21359,N_20252,N_20643);
xnor U21360 (N_21360,N_20574,N_20896);
or U21361 (N_21361,N_20777,N_20004);
or U21362 (N_21362,N_21052,N_20754);
or U21363 (N_21363,N_20827,N_20875);
xnor U21364 (N_21364,N_20208,N_20592);
and U21365 (N_21365,N_20439,N_20375);
nand U21366 (N_21366,N_20065,N_20277);
nand U21367 (N_21367,N_20225,N_20117);
xnor U21368 (N_21368,N_20104,N_21216);
nor U21369 (N_21369,N_21074,N_20301);
xor U21370 (N_21370,N_21248,N_20428);
nor U21371 (N_21371,N_20201,N_20070);
nor U21372 (N_21372,N_20144,N_20848);
nand U21373 (N_21373,N_20244,N_20475);
nand U21374 (N_21374,N_20834,N_20544);
or U21375 (N_21375,N_20283,N_21077);
and U21376 (N_21376,N_20995,N_21071);
nand U21377 (N_21377,N_20905,N_20446);
xnor U21378 (N_21378,N_20114,N_20372);
nor U21379 (N_21379,N_20745,N_20515);
nand U21380 (N_21380,N_20419,N_20031);
xnor U21381 (N_21381,N_20207,N_20554);
or U21382 (N_21382,N_20956,N_21013);
xnor U21383 (N_21383,N_20749,N_20676);
nor U21384 (N_21384,N_20994,N_21168);
and U21385 (N_21385,N_20582,N_20703);
xor U21386 (N_21386,N_20487,N_20189);
and U21387 (N_21387,N_20509,N_20180);
or U21388 (N_21388,N_20412,N_20129);
nand U21389 (N_21389,N_20761,N_20378);
xnor U21390 (N_21390,N_20006,N_20211);
or U21391 (N_21391,N_20338,N_20728);
nand U21392 (N_21392,N_20459,N_21055);
nor U21393 (N_21393,N_20265,N_21149);
nand U21394 (N_21394,N_20983,N_21063);
nor U21395 (N_21395,N_20329,N_20280);
nand U21396 (N_21396,N_20167,N_20666);
xor U21397 (N_21397,N_20379,N_20845);
or U21398 (N_21398,N_20928,N_20752);
and U21399 (N_21399,N_21117,N_20552);
and U21400 (N_21400,N_20656,N_20838);
xnor U21401 (N_21401,N_21051,N_20142);
nor U21402 (N_21402,N_20511,N_20131);
nor U21403 (N_21403,N_20274,N_21182);
nand U21404 (N_21404,N_21037,N_20714);
or U21405 (N_21405,N_20791,N_20187);
or U21406 (N_21406,N_20738,N_20241);
xor U21407 (N_21407,N_21121,N_20312);
or U21408 (N_21408,N_20514,N_20520);
xnor U21409 (N_21409,N_20737,N_20231);
nand U21410 (N_21410,N_20935,N_20969);
xor U21411 (N_21411,N_21111,N_20929);
xnor U21412 (N_21412,N_21067,N_20108);
nor U21413 (N_21413,N_20276,N_20442);
or U21414 (N_21414,N_20002,N_20568);
xor U21415 (N_21415,N_20011,N_20164);
xnor U21416 (N_21416,N_20328,N_21050);
and U21417 (N_21417,N_20176,N_20109);
or U21418 (N_21418,N_20747,N_20615);
and U21419 (N_21419,N_20123,N_20478);
nor U21420 (N_21420,N_20077,N_21208);
nor U21421 (N_21421,N_20860,N_20598);
nand U21422 (N_21422,N_20216,N_20326);
nor U21423 (N_21423,N_20548,N_20363);
nand U21424 (N_21424,N_20543,N_20767);
nor U21425 (N_21425,N_20590,N_20042);
nor U21426 (N_21426,N_20170,N_20398);
and U21427 (N_21427,N_21038,N_20008);
nor U21428 (N_21428,N_20784,N_20706);
nor U21429 (N_21429,N_20901,N_20560);
and U21430 (N_21430,N_20696,N_20251);
and U21431 (N_21431,N_20766,N_20623);
xnor U21432 (N_21432,N_21145,N_20719);
nand U21433 (N_21433,N_21240,N_20833);
xor U21434 (N_21434,N_20539,N_20627);
xor U21435 (N_21435,N_21096,N_21194);
xor U21436 (N_21436,N_20309,N_20830);
or U21437 (N_21437,N_21118,N_20053);
xor U21438 (N_21438,N_20807,N_20195);
nor U21439 (N_21439,N_20218,N_20305);
xor U21440 (N_21440,N_20270,N_20184);
or U21441 (N_21441,N_20756,N_20610);
nand U21442 (N_21442,N_20090,N_20213);
nor U21443 (N_21443,N_21217,N_20772);
xnor U21444 (N_21444,N_20545,N_20693);
nand U21445 (N_21445,N_20403,N_20235);
nor U21446 (N_21446,N_21031,N_20669);
nand U21447 (N_21447,N_20711,N_20155);
xnor U21448 (N_21448,N_20094,N_20368);
nand U21449 (N_21449,N_20458,N_20636);
xnor U21450 (N_21450,N_20339,N_20557);
and U21451 (N_21451,N_21059,N_20591);
nor U21452 (N_21452,N_21198,N_21181);
nor U21453 (N_21453,N_20771,N_20237);
xnor U21454 (N_21454,N_21241,N_20193);
xor U21455 (N_21455,N_21159,N_20400);
or U21456 (N_21456,N_20097,N_20992);
and U21457 (N_21457,N_20817,N_21042);
nand U21458 (N_21458,N_20432,N_20880);
xnor U21459 (N_21459,N_20401,N_20707);
and U21460 (N_21460,N_20816,N_20702);
xor U21461 (N_21461,N_20963,N_20899);
nor U21462 (N_21462,N_20385,N_20095);
or U21463 (N_21463,N_21218,N_20120);
and U21464 (N_21464,N_20556,N_20604);
or U21465 (N_21465,N_20832,N_21246);
or U21466 (N_21466,N_20421,N_20405);
nand U21467 (N_21467,N_21172,N_21232);
or U21468 (N_21468,N_20415,N_20606);
xor U21469 (N_21469,N_20950,N_20946);
nor U21470 (N_21470,N_20370,N_20934);
nor U21471 (N_21471,N_20182,N_21124);
nor U21472 (N_21472,N_20099,N_20585);
xor U21473 (N_21473,N_20284,N_20357);
nand U21474 (N_21474,N_21003,N_21040);
and U21475 (N_21475,N_20324,N_20970);
and U21476 (N_21476,N_20673,N_20759);
xnor U21477 (N_21477,N_20278,N_20526);
nor U21478 (N_21478,N_20017,N_20159);
and U21479 (N_21479,N_21199,N_21076);
nor U21480 (N_21480,N_20734,N_20528);
and U21481 (N_21481,N_20461,N_20670);
nand U21482 (N_21482,N_20051,N_20226);
xnor U21483 (N_21483,N_20087,N_21221);
or U21484 (N_21484,N_20410,N_20342);
or U21485 (N_21485,N_20908,N_21041);
and U21486 (N_21486,N_20549,N_20625);
or U21487 (N_21487,N_20862,N_20106);
and U21488 (N_21488,N_20281,N_21151);
xnor U21489 (N_21489,N_20721,N_20140);
or U21490 (N_21490,N_21207,N_20151);
nor U21491 (N_21491,N_20828,N_21070);
nor U21492 (N_21492,N_20056,N_20613);
nor U21493 (N_21493,N_20717,N_21000);
nand U21494 (N_21494,N_20049,N_20925);
xor U21495 (N_21495,N_20055,N_20086);
nor U21496 (N_21496,N_21195,N_20183);
nand U21497 (N_21497,N_21085,N_20092);
or U21498 (N_21498,N_20174,N_20402);
nor U21499 (N_21499,N_20234,N_20843);
and U21500 (N_21500,N_20320,N_20444);
nand U21501 (N_21501,N_20576,N_20809);
nor U21502 (N_21502,N_21080,N_21201);
or U21503 (N_21503,N_21187,N_20033);
nand U21504 (N_21504,N_20416,N_20013);
nor U21505 (N_21505,N_21177,N_21053);
nor U21506 (N_21506,N_20536,N_20466);
xnor U21507 (N_21507,N_20082,N_20774);
or U21508 (N_21508,N_21029,N_21125);
xnor U21509 (N_21509,N_21136,N_20701);
nor U21510 (N_21510,N_20629,N_20911);
or U21511 (N_21511,N_20327,N_20671);
or U21512 (N_21512,N_20012,N_20224);
nor U21513 (N_21513,N_20916,N_20130);
nand U21514 (N_21514,N_21189,N_20286);
and U21515 (N_21515,N_20230,N_20510);
and U21516 (N_21516,N_20829,N_20081);
nand U21517 (N_21517,N_21073,N_20009);
or U21518 (N_21518,N_20258,N_20364);
xor U21519 (N_21519,N_21058,N_20587);
and U21520 (N_21520,N_20323,N_20424);
and U21521 (N_21521,N_20622,N_20878);
nor U21522 (N_21522,N_21176,N_20028);
or U21523 (N_21523,N_20073,N_20726);
nand U21524 (N_21524,N_20245,N_20395);
nand U21525 (N_21525,N_21046,N_20695);
and U21526 (N_21526,N_20173,N_20330);
xor U21527 (N_21527,N_20602,N_20547);
nand U21528 (N_21528,N_20380,N_20373);
nand U21529 (N_21529,N_20869,N_20775);
or U21530 (N_21530,N_20762,N_20920);
or U21531 (N_21531,N_20315,N_20909);
nor U21532 (N_21532,N_20200,N_20168);
xor U21533 (N_21533,N_20501,N_20010);
or U21534 (N_21534,N_20516,N_21062);
and U21535 (N_21535,N_21142,N_21012);
and U21536 (N_21536,N_21022,N_20477);
and U21537 (N_21537,N_21227,N_20365);
nor U21538 (N_21538,N_20573,N_20199);
nor U21539 (N_21539,N_20264,N_20456);
or U21540 (N_21540,N_21033,N_20819);
or U21541 (N_21541,N_20007,N_20163);
nand U21542 (N_21542,N_21161,N_20639);
and U21543 (N_21543,N_21120,N_20799);
nand U21544 (N_21544,N_20993,N_20303);
nor U21545 (N_21545,N_21068,N_20507);
nand U21546 (N_21546,N_20866,N_21231);
nor U21547 (N_21547,N_20931,N_20887);
or U21548 (N_21548,N_21220,N_20076);
xnor U21549 (N_21549,N_20302,N_20663);
or U21550 (N_21550,N_20572,N_20260);
and U21551 (N_21551,N_20145,N_20959);
and U21552 (N_21552,N_21106,N_21023);
nor U21553 (N_21553,N_20882,N_20792);
or U21554 (N_21554,N_21020,N_20736);
xnor U21555 (N_21555,N_21060,N_20786);
or U21556 (N_21556,N_20524,N_20188);
nor U21557 (N_21557,N_20594,N_21153);
xor U21558 (N_21558,N_20488,N_21169);
and U21559 (N_21559,N_21157,N_20987);
xor U21560 (N_21560,N_21147,N_20674);
nand U21561 (N_21561,N_21086,N_20098);
xor U21562 (N_21562,N_21030,N_20154);
nand U21563 (N_21563,N_20680,N_20232);
or U21564 (N_21564,N_20735,N_20036);
nor U21565 (N_21565,N_21109,N_20710);
xor U21566 (N_21566,N_20291,N_20340);
or U21567 (N_21567,N_20452,N_20445);
or U21568 (N_21568,N_20881,N_20351);
nand U21569 (N_21569,N_20437,N_20965);
and U21570 (N_21570,N_20689,N_20944);
nand U21571 (N_21571,N_20961,N_20440);
and U21572 (N_21572,N_20932,N_20185);
nor U21573 (N_21573,N_20222,N_20947);
xnor U21574 (N_21574,N_20898,N_20382);
or U21575 (N_21575,N_21015,N_20855);
nor U21576 (N_21576,N_20684,N_20849);
xor U21577 (N_21577,N_20678,N_20377);
nor U21578 (N_21578,N_20236,N_20955);
nand U21579 (N_21579,N_20506,N_20753);
xnor U21580 (N_21580,N_20133,N_20839);
nand U21581 (N_21581,N_21171,N_20872);
nor U21582 (N_21582,N_20780,N_20397);
nand U21583 (N_21583,N_20266,N_20782);
nor U21584 (N_21584,N_20317,N_20078);
nand U21585 (N_21585,N_20744,N_20025);
nand U21586 (N_21586,N_20641,N_20583);
nor U21587 (N_21587,N_20088,N_20128);
nor U21588 (N_21588,N_21001,N_20127);
nor U21589 (N_21589,N_20884,N_20742);
xnor U21590 (N_21590,N_20859,N_21226);
or U21591 (N_21591,N_20648,N_20289);
nand U21592 (N_21592,N_21011,N_20346);
xnor U21593 (N_21593,N_20550,N_20480);
nand U21594 (N_21594,N_20124,N_20067);
or U21595 (N_21595,N_20022,N_20812);
nand U21596 (N_21596,N_21064,N_20495);
nand U21597 (N_21597,N_20075,N_20976);
or U21598 (N_21598,N_20467,N_20060);
nor U21599 (N_21599,N_20386,N_21009);
nand U21600 (N_21600,N_20599,N_20581);
xnor U21601 (N_21601,N_21211,N_21139);
xor U21602 (N_21602,N_20443,N_20249);
nor U21603 (N_21603,N_21079,N_20331);
nor U21604 (N_21604,N_20621,N_20141);
xnor U21605 (N_21605,N_20668,N_20785);
and U21606 (N_21606,N_20997,N_20253);
nor U21607 (N_21607,N_20358,N_21091);
nor U21608 (N_21608,N_20387,N_20781);
or U21609 (N_21609,N_21245,N_20179);
nor U21610 (N_21610,N_20408,N_20657);
or U21611 (N_21611,N_20394,N_20892);
nand U21612 (N_21612,N_21239,N_20152);
nand U21613 (N_21613,N_20064,N_20068);
and U21614 (N_21614,N_20299,N_20221);
nor U21615 (N_21615,N_20794,N_20600);
or U21616 (N_21616,N_20915,N_21010);
nand U21617 (N_21617,N_21123,N_20229);
nand U21618 (N_21618,N_20250,N_20161);
nand U21619 (N_21619,N_21116,N_20441);
nor U21620 (N_21620,N_20977,N_20027);
xnor U21621 (N_21621,N_21002,N_21108);
xor U21622 (N_21622,N_20019,N_20578);
and U21623 (N_21623,N_20972,N_20293);
and U21624 (N_21624,N_20895,N_20769);
and U21625 (N_21625,N_20608,N_20725);
nor U21626 (N_21626,N_20212,N_20665);
nor U21627 (N_21627,N_20939,N_20662);
nor U21628 (N_21628,N_20879,N_21223);
nor U21629 (N_21629,N_20584,N_20733);
and U21630 (N_21630,N_20058,N_21129);
nand U21631 (N_21631,N_20268,N_20620);
nor U21632 (N_21632,N_20609,N_20350);
nor U21633 (N_21633,N_20389,N_20374);
nand U21634 (N_21634,N_20001,N_20982);
and U21635 (N_21635,N_20746,N_20523);
and U21636 (N_21636,N_20427,N_20923);
xnor U21637 (N_21637,N_20015,N_20448);
xnor U21638 (N_21638,N_20043,N_20741);
nor U21639 (N_21639,N_20903,N_21007);
xnor U21640 (N_21640,N_20649,N_20227);
nor U21641 (N_21641,N_20209,N_20697);
xnor U21642 (N_21642,N_20659,N_20198);
or U21643 (N_21643,N_20851,N_20938);
nand U21644 (N_21644,N_20897,N_20631);
nor U21645 (N_21645,N_20138,N_20748);
nand U21646 (N_21646,N_20789,N_20793);
or U21647 (N_21647,N_20473,N_21102);
nand U21648 (N_21648,N_20362,N_20059);
nand U21649 (N_21649,N_20926,N_21036);
nor U21650 (N_21650,N_20732,N_20204);
and U21651 (N_21651,N_20661,N_20044);
or U21652 (N_21652,N_20958,N_20166);
and U21653 (N_21653,N_20093,N_20113);
xor U21654 (N_21654,N_20731,N_20513);
xor U21655 (N_21655,N_21144,N_20066);
xnor U21656 (N_21656,N_20893,N_20722);
xor U21657 (N_21657,N_20420,N_20047);
or U21658 (N_21658,N_20413,N_21093);
or U21659 (N_21659,N_21222,N_20924);
or U21660 (N_21660,N_21078,N_21016);
nor U21661 (N_21661,N_21045,N_21005);
nand U21662 (N_21662,N_20655,N_20831);
xor U21663 (N_21663,N_21215,N_20259);
nor U21664 (N_21664,N_20319,N_20984);
and U21665 (N_21665,N_20256,N_20751);
xnor U21666 (N_21666,N_21190,N_20646);
xnor U21667 (N_21667,N_21204,N_20802);
nand U21668 (N_21668,N_20089,N_20263);
xor U21669 (N_21669,N_20156,N_20718);
xnor U21670 (N_21670,N_20438,N_20571);
nand U21671 (N_21671,N_20535,N_20790);
nand U21672 (N_21672,N_21024,N_20335);
xnor U21673 (N_21673,N_20215,N_20148);
nor U21674 (N_21674,N_20463,N_21018);
nor U21675 (N_21675,N_20797,N_20922);
xor U21676 (N_21676,N_20907,N_20914);
and U21677 (N_21677,N_20529,N_20146);
or U21678 (N_21678,N_21138,N_20096);
and U21679 (N_21679,N_20618,N_20434);
nor U21680 (N_21680,N_21006,N_21162);
or U21681 (N_21681,N_20645,N_20533);
nand U21682 (N_21682,N_20962,N_20624);
and U21683 (N_21683,N_20032,N_20111);
or U21684 (N_21684,N_21249,N_20071);
or U21685 (N_21685,N_21099,N_20796);
nor U21686 (N_21686,N_20223,N_21114);
nor U21687 (N_21687,N_20079,N_20417);
nor U21688 (N_21688,N_20808,N_20023);
nand U21689 (N_21689,N_20530,N_21026);
nor U21690 (N_21690,N_20764,N_20074);
nor U21691 (N_21691,N_20354,N_20353);
xnor U21692 (N_21692,N_20178,N_20936);
and U21693 (N_21693,N_21174,N_20690);
xor U21694 (N_21694,N_20344,N_20798);
nor U21695 (N_21695,N_20886,N_20597);
and U21696 (N_21696,N_20254,N_20974);
and U21697 (N_21697,N_20565,N_20683);
nor U21698 (N_21698,N_21081,N_20407);
and U21699 (N_21699,N_20029,N_21043);
or U21700 (N_21700,N_20988,N_21100);
or U21701 (N_21701,N_20595,N_21193);
and U21702 (N_21702,N_20682,N_20700);
xnor U21703 (N_21703,N_20743,N_20479);
and U21704 (N_21704,N_20913,N_20943);
xnor U21705 (N_21705,N_21137,N_21048);
xnor U21706 (N_21706,N_20558,N_20383);
nor U21707 (N_21707,N_20484,N_20638);
and U21708 (N_21708,N_20041,N_20160);
and U21709 (N_21709,N_20247,N_20952);
xor U21710 (N_21710,N_20460,N_20083);
and U21711 (N_21711,N_20057,N_20292);
or U21712 (N_21712,N_20390,N_20371);
xnor U21713 (N_21713,N_20806,N_21017);
and U21714 (N_21714,N_20169,N_21243);
and U21715 (N_21715,N_20888,N_21127);
nand U21716 (N_21716,N_21143,N_20103);
and U21717 (N_21717,N_20430,N_20973);
and U21718 (N_21718,N_20240,N_21115);
nand U21719 (N_21719,N_20220,N_20085);
nand U21720 (N_21720,N_21019,N_20716);
and U21721 (N_21721,N_20532,N_20811);
or U21722 (N_21722,N_20654,N_20628);
nand U21723 (N_21723,N_20891,N_20489);
or U21724 (N_21724,N_20713,N_20820);
nor U21725 (N_21725,N_20825,N_20770);
and U21726 (N_21726,N_20306,N_20534);
or U21727 (N_21727,N_21188,N_20779);
xor U21728 (N_21728,N_20740,N_20294);
nor U21729 (N_21729,N_21097,N_20186);
nor U21730 (N_21730,N_20119,N_20577);
or U21731 (N_21731,N_21247,N_20494);
nor U21732 (N_21732,N_20553,N_20642);
or U21733 (N_21733,N_20894,N_20776);
nor U21734 (N_21734,N_21130,N_21213);
nor U21735 (N_21735,N_21032,N_20607);
or U21736 (N_21736,N_21160,N_20172);
and U21737 (N_21737,N_20687,N_20110);
xor U21738 (N_21738,N_20196,N_20307);
nand U21739 (N_21739,N_21061,N_20727);
nand U21740 (N_21740,N_20136,N_20462);
nand U21741 (N_21741,N_20971,N_20472);
nor U21742 (N_21742,N_20308,N_20685);
or U21743 (N_21743,N_20758,N_20739);
xor U21744 (N_21744,N_20100,N_20046);
nand U21745 (N_21745,N_20267,N_20757);
and U21746 (N_21746,N_20768,N_20423);
or U21747 (N_21747,N_20837,N_20393);
xnor U21748 (N_21748,N_21154,N_21132);
or U21749 (N_21749,N_20334,N_20729);
or U21750 (N_21750,N_20902,N_20210);
nand U21751 (N_21751,N_20989,N_21164);
and U21752 (N_21752,N_20248,N_20867);
or U21753 (N_21753,N_21244,N_20579);
nand U21754 (N_21754,N_21200,N_21126);
nand U21755 (N_21755,N_20116,N_20233);
nand U21756 (N_21756,N_20699,N_20868);
xnor U21757 (N_21757,N_20788,N_20504);
nor U21758 (N_21758,N_20436,N_20411);
xor U21759 (N_21759,N_20966,N_20203);
nor U21760 (N_21760,N_20626,N_21119);
nor U21761 (N_21761,N_20945,N_20325);
xnor U21762 (N_21762,N_20021,N_20271);
and U21763 (N_21763,N_20181,N_20202);
nor U21764 (N_21764,N_21205,N_20844);
or U21765 (N_21765,N_20691,N_20672);
xor U21766 (N_21766,N_21083,N_20016);
nor U21767 (N_21767,N_20311,N_20877);
nor U21768 (N_21768,N_21025,N_20927);
nor U21769 (N_21769,N_21054,N_20321);
or U21770 (N_21770,N_20137,N_20239);
nor U21771 (N_21771,N_21047,N_20500);
xnor U21772 (N_21772,N_20705,N_20062);
or U21773 (N_21773,N_21021,N_21158);
nor U21774 (N_21774,N_20341,N_20647);
xor U21775 (N_21775,N_20508,N_21197);
and U21776 (N_21776,N_20503,N_20158);
or U21777 (N_21777,N_20490,N_20105);
xnor U21778 (N_21778,N_20755,N_20343);
or U21779 (N_21779,N_20593,N_20349);
and U21780 (N_21780,N_20863,N_21039);
xnor U21781 (N_21781,N_20453,N_20026);
nand U21782 (N_21782,N_21004,N_20910);
nand U21783 (N_21783,N_20564,N_20688);
nor U21784 (N_21784,N_21069,N_20773);
and U21785 (N_21785,N_20653,N_20852);
nand U21786 (N_21786,N_20667,N_20333);
xnor U21787 (N_21787,N_21087,N_20949);
nor U21788 (N_21788,N_20633,N_20679);
nand U21789 (N_21789,N_20192,N_20964);
xnor U21790 (N_21790,N_20650,N_21233);
nor U21791 (N_21791,N_21105,N_20917);
xnor U21792 (N_21792,N_20813,N_21152);
and U21793 (N_21793,N_20206,N_21178);
or U21794 (N_21794,N_20228,N_20054);
or U21795 (N_21795,N_20361,N_20521);
or U21796 (N_21796,N_21140,N_20783);
and U21797 (N_21797,N_20102,N_20765);
xor U21798 (N_21798,N_20723,N_20611);
nor U21799 (N_21799,N_20692,N_20310);
and U21800 (N_21800,N_20651,N_20414);
or U21801 (N_21801,N_20589,N_20040);
nor U21802 (N_21802,N_20356,N_21185);
nor U21803 (N_21803,N_21183,N_20854);
or U21804 (N_21804,N_20803,N_21101);
nor U21805 (N_21805,N_20177,N_21131);
nor U21806 (N_21806,N_20555,N_20518);
and U21807 (N_21807,N_20760,N_21219);
or U21808 (N_21808,N_20150,N_20313);
nor U21809 (N_21809,N_20841,N_20873);
and U21810 (N_21810,N_21148,N_20360);
nand U21811 (N_21811,N_21242,N_20512);
and U21812 (N_21812,N_20352,N_20968);
and U21813 (N_21813,N_20296,N_20522);
or U21814 (N_21814,N_20470,N_21072);
nor U21815 (N_21815,N_20348,N_21034);
xor U21816 (N_21816,N_20285,N_21113);
and U21817 (N_21817,N_20399,N_21224);
xor U21818 (N_21818,N_20493,N_20605);
or U21819 (N_21819,N_20847,N_20122);
nor U21820 (N_21820,N_20243,N_20940);
nor U21821 (N_21821,N_20708,N_20425);
nor U21822 (N_21822,N_21134,N_20981);
nand U21823 (N_21823,N_20948,N_20061);
nor U21824 (N_21824,N_20586,N_20337);
nand U21825 (N_21825,N_20601,N_20038);
nor U21826 (N_21826,N_20422,N_20804);
and U21827 (N_21827,N_20409,N_21056);
and U21828 (N_21828,N_20107,N_20391);
or U21829 (N_21829,N_20730,N_21049);
xor U21830 (N_21830,N_20637,N_20125);
and U21831 (N_21831,N_20039,N_20750);
nand U21832 (N_21832,N_20469,N_20538);
nor U21833 (N_21833,N_20921,N_20559);
nor U21834 (N_21834,N_20474,N_20517);
nor U21835 (N_21835,N_21156,N_20975);
nand U21836 (N_21836,N_20763,N_20194);
nand U21837 (N_21837,N_21014,N_20255);
and U21838 (N_21838,N_21236,N_20883);
and U21839 (N_21839,N_20084,N_20000);
or U21840 (N_21840,N_20686,N_20542);
and U21841 (N_21841,N_20464,N_20214);
or U21842 (N_21842,N_20709,N_20821);
and U21843 (N_21843,N_20724,N_20991);
xnor U21844 (N_21844,N_20030,N_20937);
and U21845 (N_21845,N_20418,N_20996);
and U21846 (N_21846,N_21180,N_21065);
and U21847 (N_21847,N_20112,N_20842);
xnor U21848 (N_21848,N_20890,N_20392);
nand U21849 (N_21849,N_20482,N_21184);
or U21850 (N_21850,N_20426,N_21163);
nand U21851 (N_21851,N_20603,N_20450);
nor U21852 (N_21852,N_20502,N_20171);
nor U21853 (N_21853,N_20035,N_20496);
nor U21854 (N_21854,N_21238,N_20052);
and U21855 (N_21855,N_20003,N_21234);
nand U21856 (N_21856,N_20191,N_20126);
nor U21857 (N_21857,N_20499,N_20304);
xor U21858 (N_21858,N_20275,N_20630);
and U21859 (N_21859,N_21110,N_21135);
or U21860 (N_21860,N_20261,N_20614);
xor U21861 (N_21861,N_20652,N_21206);
and U21862 (N_21862,N_20826,N_21225);
xor U21863 (N_21863,N_20367,N_21066);
nor U21864 (N_21864,N_20960,N_20139);
xnor U21865 (N_21865,N_20918,N_20580);
or U21866 (N_21866,N_20836,N_20919);
or U21867 (N_21867,N_20435,N_20957);
xor U21868 (N_21868,N_20238,N_20778);
or U21869 (N_21869,N_20497,N_21170);
nand U21870 (N_21870,N_20404,N_21084);
and U21871 (N_21871,N_20454,N_21075);
nor U21872 (N_21872,N_20165,N_21089);
xor U21873 (N_21873,N_20900,N_20476);
xor U21874 (N_21874,N_20677,N_20889);
and U21875 (N_21875,N_20408,N_20858);
nor U21876 (N_21876,N_20151,N_21004);
nand U21877 (N_21877,N_20095,N_20059);
nor U21878 (N_21878,N_20451,N_21229);
nor U21879 (N_21879,N_20393,N_20249);
and U21880 (N_21880,N_20577,N_20706);
nor U21881 (N_21881,N_21206,N_20066);
nor U21882 (N_21882,N_20964,N_20817);
xnor U21883 (N_21883,N_20170,N_21056);
or U21884 (N_21884,N_20191,N_20979);
nand U21885 (N_21885,N_20965,N_20458);
or U21886 (N_21886,N_20481,N_20351);
or U21887 (N_21887,N_20565,N_20159);
xnor U21888 (N_21888,N_20522,N_20492);
or U21889 (N_21889,N_20849,N_20547);
nand U21890 (N_21890,N_20456,N_20379);
or U21891 (N_21891,N_20310,N_20606);
or U21892 (N_21892,N_20350,N_20625);
xor U21893 (N_21893,N_20530,N_20031);
and U21894 (N_21894,N_20471,N_21007);
and U21895 (N_21895,N_20676,N_20922);
and U21896 (N_21896,N_20431,N_20764);
nand U21897 (N_21897,N_20583,N_21072);
nand U21898 (N_21898,N_20444,N_21177);
or U21899 (N_21899,N_20094,N_20828);
nor U21900 (N_21900,N_20935,N_20181);
nand U21901 (N_21901,N_20752,N_20824);
or U21902 (N_21902,N_20820,N_20693);
xor U21903 (N_21903,N_20253,N_21180);
xnor U21904 (N_21904,N_20186,N_20579);
or U21905 (N_21905,N_20788,N_20799);
nor U21906 (N_21906,N_20027,N_20116);
nor U21907 (N_21907,N_21212,N_20226);
nand U21908 (N_21908,N_20141,N_20026);
xnor U21909 (N_21909,N_20001,N_20421);
nor U21910 (N_21910,N_20284,N_20405);
or U21911 (N_21911,N_20678,N_21158);
xor U21912 (N_21912,N_20163,N_20178);
xor U21913 (N_21913,N_20467,N_20537);
nor U21914 (N_21914,N_21213,N_20545);
xnor U21915 (N_21915,N_20898,N_20591);
xor U21916 (N_21916,N_20490,N_20052);
nor U21917 (N_21917,N_20915,N_21215);
nor U21918 (N_21918,N_20969,N_20146);
or U21919 (N_21919,N_20470,N_20576);
nand U21920 (N_21920,N_20529,N_21171);
nand U21921 (N_21921,N_21019,N_21118);
or U21922 (N_21922,N_20626,N_20787);
nor U21923 (N_21923,N_20165,N_20957);
xor U21924 (N_21924,N_21069,N_20198);
nor U21925 (N_21925,N_20803,N_20542);
nand U21926 (N_21926,N_20176,N_20926);
xnor U21927 (N_21927,N_20952,N_20617);
nor U21928 (N_21928,N_20087,N_20308);
nand U21929 (N_21929,N_21214,N_21186);
nand U21930 (N_21930,N_20994,N_20061);
nand U21931 (N_21931,N_21087,N_20996);
xnor U21932 (N_21932,N_20929,N_21028);
nand U21933 (N_21933,N_20693,N_20256);
nand U21934 (N_21934,N_20348,N_20816);
xnor U21935 (N_21935,N_20920,N_20463);
xnor U21936 (N_21936,N_20091,N_20901);
nor U21937 (N_21937,N_20098,N_20962);
nand U21938 (N_21938,N_20150,N_21034);
nand U21939 (N_21939,N_21003,N_20223);
xnor U21940 (N_21940,N_21152,N_20555);
nor U21941 (N_21941,N_20044,N_20988);
or U21942 (N_21942,N_20481,N_21218);
nor U21943 (N_21943,N_20676,N_20945);
nor U21944 (N_21944,N_20473,N_20878);
or U21945 (N_21945,N_20679,N_20536);
xnor U21946 (N_21946,N_20619,N_21169);
xnor U21947 (N_21947,N_20185,N_20626);
or U21948 (N_21948,N_20459,N_20497);
nor U21949 (N_21949,N_20071,N_20016);
nand U21950 (N_21950,N_20817,N_20505);
xnor U21951 (N_21951,N_20143,N_20025);
nand U21952 (N_21952,N_20731,N_21166);
nand U21953 (N_21953,N_20172,N_20416);
or U21954 (N_21954,N_20890,N_20190);
or U21955 (N_21955,N_21187,N_20479);
and U21956 (N_21956,N_20455,N_20160);
nand U21957 (N_21957,N_21190,N_21013);
xnor U21958 (N_21958,N_20587,N_20866);
xnor U21959 (N_21959,N_20539,N_21031);
and U21960 (N_21960,N_21167,N_21080);
nand U21961 (N_21961,N_21066,N_20409);
and U21962 (N_21962,N_20359,N_20784);
nand U21963 (N_21963,N_20195,N_21012);
nand U21964 (N_21964,N_21056,N_20319);
and U21965 (N_21965,N_20038,N_20359);
xor U21966 (N_21966,N_20232,N_20361);
and U21967 (N_21967,N_20825,N_21188);
and U21968 (N_21968,N_20658,N_20286);
or U21969 (N_21969,N_20082,N_20799);
or U21970 (N_21970,N_20991,N_20511);
or U21971 (N_21971,N_20680,N_21247);
and U21972 (N_21972,N_20754,N_21228);
nor U21973 (N_21973,N_20591,N_21010);
nor U21974 (N_21974,N_20722,N_20317);
nand U21975 (N_21975,N_20338,N_21240);
xnor U21976 (N_21976,N_20147,N_20710);
and U21977 (N_21977,N_20609,N_20369);
or U21978 (N_21978,N_20440,N_21233);
xnor U21979 (N_21979,N_20075,N_20093);
or U21980 (N_21980,N_20088,N_20913);
nand U21981 (N_21981,N_20306,N_20104);
xnor U21982 (N_21982,N_20410,N_20421);
nand U21983 (N_21983,N_20083,N_21141);
nor U21984 (N_21984,N_20717,N_20590);
nor U21985 (N_21985,N_21206,N_20920);
or U21986 (N_21986,N_20471,N_21195);
and U21987 (N_21987,N_20799,N_21122);
nand U21988 (N_21988,N_20205,N_21004);
xnor U21989 (N_21989,N_20711,N_20081);
and U21990 (N_21990,N_20666,N_20496);
and U21991 (N_21991,N_20064,N_20238);
and U21992 (N_21992,N_21195,N_20957);
nor U21993 (N_21993,N_20636,N_20345);
nor U21994 (N_21994,N_21099,N_20591);
xnor U21995 (N_21995,N_20265,N_20724);
or U21996 (N_21996,N_20721,N_20163);
nand U21997 (N_21997,N_20417,N_20294);
or U21998 (N_21998,N_20775,N_20456);
nor U21999 (N_21999,N_20388,N_20065);
nand U22000 (N_22000,N_21070,N_21115);
and U22001 (N_22001,N_21236,N_20572);
nor U22002 (N_22002,N_20881,N_20414);
and U22003 (N_22003,N_20636,N_20763);
or U22004 (N_22004,N_20086,N_20992);
or U22005 (N_22005,N_20260,N_20722);
nand U22006 (N_22006,N_20608,N_20194);
nor U22007 (N_22007,N_20846,N_20847);
xor U22008 (N_22008,N_21099,N_20252);
nor U22009 (N_22009,N_20453,N_21200);
or U22010 (N_22010,N_20661,N_20539);
or U22011 (N_22011,N_20672,N_21021);
xor U22012 (N_22012,N_20279,N_20651);
and U22013 (N_22013,N_20425,N_20749);
nor U22014 (N_22014,N_21136,N_20219);
and U22015 (N_22015,N_20077,N_20473);
or U22016 (N_22016,N_20362,N_20297);
xor U22017 (N_22017,N_20005,N_20998);
nor U22018 (N_22018,N_20715,N_21131);
and U22019 (N_22019,N_20918,N_20274);
xor U22020 (N_22020,N_20364,N_20113);
or U22021 (N_22021,N_20239,N_20602);
and U22022 (N_22022,N_20572,N_20518);
nor U22023 (N_22023,N_21112,N_20204);
xnor U22024 (N_22024,N_20475,N_21105);
and U22025 (N_22025,N_20100,N_20761);
xor U22026 (N_22026,N_20332,N_20474);
nor U22027 (N_22027,N_20473,N_20033);
and U22028 (N_22028,N_20464,N_21145);
or U22029 (N_22029,N_20887,N_20664);
nor U22030 (N_22030,N_20983,N_20005);
xor U22031 (N_22031,N_20430,N_20822);
and U22032 (N_22032,N_20460,N_21203);
nor U22033 (N_22033,N_20566,N_21158);
xnor U22034 (N_22034,N_20077,N_20263);
and U22035 (N_22035,N_20425,N_20440);
nor U22036 (N_22036,N_20816,N_20427);
xnor U22037 (N_22037,N_20862,N_21141);
xor U22038 (N_22038,N_20649,N_20231);
and U22039 (N_22039,N_20300,N_20966);
nand U22040 (N_22040,N_20426,N_20632);
nor U22041 (N_22041,N_20301,N_20432);
or U22042 (N_22042,N_21139,N_20367);
and U22043 (N_22043,N_20244,N_21133);
nor U22044 (N_22044,N_20594,N_21091);
or U22045 (N_22045,N_20992,N_20539);
xor U22046 (N_22046,N_20614,N_21161);
or U22047 (N_22047,N_21033,N_20307);
and U22048 (N_22048,N_20963,N_20261);
xnor U22049 (N_22049,N_20370,N_20251);
nand U22050 (N_22050,N_20213,N_20019);
or U22051 (N_22051,N_20252,N_20587);
nand U22052 (N_22052,N_21023,N_20766);
and U22053 (N_22053,N_20433,N_20754);
and U22054 (N_22054,N_20334,N_20032);
or U22055 (N_22055,N_20136,N_20279);
xnor U22056 (N_22056,N_20456,N_21199);
or U22057 (N_22057,N_20278,N_20119);
xor U22058 (N_22058,N_20717,N_21161);
nor U22059 (N_22059,N_20796,N_20175);
and U22060 (N_22060,N_20597,N_20209);
nor U22061 (N_22061,N_20037,N_20564);
nor U22062 (N_22062,N_21178,N_21190);
nor U22063 (N_22063,N_21067,N_20771);
nand U22064 (N_22064,N_20177,N_20445);
nor U22065 (N_22065,N_20046,N_21209);
xor U22066 (N_22066,N_21041,N_20048);
and U22067 (N_22067,N_20847,N_20383);
or U22068 (N_22068,N_20853,N_21242);
nor U22069 (N_22069,N_20679,N_20333);
xor U22070 (N_22070,N_20534,N_20318);
nand U22071 (N_22071,N_21078,N_21001);
and U22072 (N_22072,N_20272,N_20664);
xnor U22073 (N_22073,N_20678,N_20091);
or U22074 (N_22074,N_20095,N_20197);
and U22075 (N_22075,N_21119,N_21096);
nand U22076 (N_22076,N_21018,N_20328);
nand U22077 (N_22077,N_20486,N_20505);
nand U22078 (N_22078,N_20617,N_20535);
nor U22079 (N_22079,N_20723,N_20907);
xor U22080 (N_22080,N_20810,N_20392);
nand U22081 (N_22081,N_20834,N_20916);
nor U22082 (N_22082,N_20523,N_20875);
nand U22083 (N_22083,N_20040,N_21220);
or U22084 (N_22084,N_20054,N_20800);
xor U22085 (N_22085,N_20586,N_21138);
or U22086 (N_22086,N_20783,N_21168);
xor U22087 (N_22087,N_20012,N_20962);
xnor U22088 (N_22088,N_20811,N_21206);
nor U22089 (N_22089,N_20960,N_21121);
or U22090 (N_22090,N_20581,N_20268);
nor U22091 (N_22091,N_20523,N_20847);
nor U22092 (N_22092,N_20429,N_20870);
and U22093 (N_22093,N_20750,N_20022);
xor U22094 (N_22094,N_20859,N_20074);
and U22095 (N_22095,N_20375,N_20214);
nor U22096 (N_22096,N_20092,N_21196);
and U22097 (N_22097,N_20294,N_20626);
nor U22098 (N_22098,N_21058,N_20771);
nor U22099 (N_22099,N_20594,N_21092);
nand U22100 (N_22100,N_20095,N_20552);
and U22101 (N_22101,N_20546,N_21163);
xnor U22102 (N_22102,N_20818,N_20254);
xor U22103 (N_22103,N_20164,N_20381);
nor U22104 (N_22104,N_20243,N_20864);
or U22105 (N_22105,N_20275,N_20525);
xnor U22106 (N_22106,N_21242,N_21064);
and U22107 (N_22107,N_20001,N_20257);
nand U22108 (N_22108,N_20679,N_21246);
nor U22109 (N_22109,N_20894,N_20269);
nand U22110 (N_22110,N_20943,N_21124);
xnor U22111 (N_22111,N_20809,N_20885);
xnor U22112 (N_22112,N_20654,N_20806);
nor U22113 (N_22113,N_20266,N_20034);
nand U22114 (N_22114,N_20592,N_20326);
nor U22115 (N_22115,N_20504,N_20667);
and U22116 (N_22116,N_21225,N_20308);
xor U22117 (N_22117,N_21163,N_21088);
or U22118 (N_22118,N_20758,N_20186);
and U22119 (N_22119,N_20236,N_20078);
nor U22120 (N_22120,N_20720,N_20549);
or U22121 (N_22121,N_20013,N_21067);
nor U22122 (N_22122,N_20006,N_21167);
or U22123 (N_22123,N_20794,N_20795);
or U22124 (N_22124,N_20968,N_21213);
xnor U22125 (N_22125,N_20558,N_20633);
or U22126 (N_22126,N_20589,N_20334);
or U22127 (N_22127,N_20637,N_20274);
or U22128 (N_22128,N_20177,N_20755);
and U22129 (N_22129,N_20848,N_21244);
nor U22130 (N_22130,N_20782,N_20362);
and U22131 (N_22131,N_20455,N_20205);
or U22132 (N_22132,N_20718,N_20769);
nor U22133 (N_22133,N_21097,N_20425);
xnor U22134 (N_22134,N_20472,N_20282);
nor U22135 (N_22135,N_21024,N_20331);
nor U22136 (N_22136,N_21013,N_20646);
or U22137 (N_22137,N_20061,N_20487);
or U22138 (N_22138,N_20375,N_20722);
and U22139 (N_22139,N_20768,N_20755);
or U22140 (N_22140,N_20117,N_20754);
xnor U22141 (N_22141,N_21130,N_20731);
or U22142 (N_22142,N_20193,N_20569);
nor U22143 (N_22143,N_20866,N_20454);
nand U22144 (N_22144,N_20025,N_20011);
xnor U22145 (N_22145,N_20480,N_20405);
nand U22146 (N_22146,N_21061,N_20577);
nand U22147 (N_22147,N_20039,N_20836);
xor U22148 (N_22148,N_21078,N_21239);
xnor U22149 (N_22149,N_20952,N_20637);
and U22150 (N_22150,N_20619,N_20249);
nand U22151 (N_22151,N_20111,N_20209);
xor U22152 (N_22152,N_21128,N_20457);
xnor U22153 (N_22153,N_20357,N_20939);
xnor U22154 (N_22154,N_20485,N_20642);
and U22155 (N_22155,N_20061,N_20919);
or U22156 (N_22156,N_20949,N_21046);
xnor U22157 (N_22157,N_20546,N_20701);
nor U22158 (N_22158,N_21135,N_20306);
and U22159 (N_22159,N_20511,N_21011);
nor U22160 (N_22160,N_21040,N_20411);
and U22161 (N_22161,N_20250,N_20700);
and U22162 (N_22162,N_20336,N_21235);
and U22163 (N_22163,N_20310,N_20268);
and U22164 (N_22164,N_20920,N_20032);
or U22165 (N_22165,N_20933,N_20534);
nor U22166 (N_22166,N_20215,N_20912);
nand U22167 (N_22167,N_20298,N_21210);
nand U22168 (N_22168,N_20771,N_20386);
nor U22169 (N_22169,N_21163,N_20729);
xor U22170 (N_22170,N_20828,N_20542);
xnor U22171 (N_22171,N_20216,N_20412);
and U22172 (N_22172,N_20409,N_20713);
nand U22173 (N_22173,N_21231,N_20383);
and U22174 (N_22174,N_21050,N_20980);
nor U22175 (N_22175,N_20675,N_20425);
or U22176 (N_22176,N_21172,N_20892);
nor U22177 (N_22177,N_20511,N_20575);
xor U22178 (N_22178,N_20430,N_21117);
and U22179 (N_22179,N_20022,N_20540);
or U22180 (N_22180,N_20394,N_20321);
nand U22181 (N_22181,N_21075,N_20841);
nor U22182 (N_22182,N_20645,N_20787);
and U22183 (N_22183,N_21084,N_20804);
or U22184 (N_22184,N_21189,N_20666);
xnor U22185 (N_22185,N_20508,N_20978);
or U22186 (N_22186,N_20739,N_20668);
nor U22187 (N_22187,N_21235,N_20209);
nor U22188 (N_22188,N_20170,N_20006);
xnor U22189 (N_22189,N_20828,N_20847);
or U22190 (N_22190,N_20329,N_20121);
nand U22191 (N_22191,N_20571,N_20358);
or U22192 (N_22192,N_21222,N_20076);
nor U22193 (N_22193,N_20917,N_20991);
nand U22194 (N_22194,N_20888,N_20060);
xnor U22195 (N_22195,N_21229,N_21220);
nand U22196 (N_22196,N_20480,N_20610);
and U22197 (N_22197,N_20406,N_20949);
nand U22198 (N_22198,N_20000,N_20144);
nor U22199 (N_22199,N_21072,N_20999);
nor U22200 (N_22200,N_20777,N_20591);
nand U22201 (N_22201,N_20551,N_21015);
and U22202 (N_22202,N_20410,N_20626);
nor U22203 (N_22203,N_20574,N_20580);
xor U22204 (N_22204,N_20703,N_20540);
and U22205 (N_22205,N_20042,N_20993);
xnor U22206 (N_22206,N_20170,N_20468);
xnor U22207 (N_22207,N_21203,N_21227);
and U22208 (N_22208,N_20444,N_20569);
and U22209 (N_22209,N_20029,N_20524);
nand U22210 (N_22210,N_20972,N_20175);
or U22211 (N_22211,N_20301,N_20679);
nand U22212 (N_22212,N_20434,N_20596);
and U22213 (N_22213,N_20026,N_20165);
and U22214 (N_22214,N_20677,N_21239);
nor U22215 (N_22215,N_20101,N_20287);
xnor U22216 (N_22216,N_20196,N_20935);
xnor U22217 (N_22217,N_20371,N_20591);
xnor U22218 (N_22218,N_20960,N_20356);
nor U22219 (N_22219,N_20281,N_20696);
xor U22220 (N_22220,N_20169,N_20019);
nand U22221 (N_22221,N_20823,N_20163);
and U22222 (N_22222,N_20827,N_20882);
and U22223 (N_22223,N_20853,N_20742);
and U22224 (N_22224,N_20144,N_20562);
nor U22225 (N_22225,N_20304,N_20323);
and U22226 (N_22226,N_20272,N_20163);
nand U22227 (N_22227,N_21048,N_20688);
nor U22228 (N_22228,N_20897,N_20650);
xnor U22229 (N_22229,N_20692,N_21063);
or U22230 (N_22230,N_20210,N_20087);
and U22231 (N_22231,N_20939,N_20097);
xor U22232 (N_22232,N_20480,N_20250);
or U22233 (N_22233,N_20921,N_20507);
and U22234 (N_22234,N_20042,N_20217);
or U22235 (N_22235,N_20280,N_21110);
and U22236 (N_22236,N_20589,N_20408);
nand U22237 (N_22237,N_20661,N_20425);
and U22238 (N_22238,N_20202,N_20045);
nand U22239 (N_22239,N_20255,N_20587);
nand U22240 (N_22240,N_20188,N_21219);
xor U22241 (N_22241,N_20428,N_20905);
nor U22242 (N_22242,N_20196,N_20191);
xnor U22243 (N_22243,N_20673,N_20799);
xor U22244 (N_22244,N_20362,N_20171);
nor U22245 (N_22245,N_20928,N_20343);
and U22246 (N_22246,N_20047,N_20331);
and U22247 (N_22247,N_20315,N_20075);
and U22248 (N_22248,N_20454,N_20125);
and U22249 (N_22249,N_20225,N_20238);
nand U22250 (N_22250,N_20918,N_20894);
nand U22251 (N_22251,N_20004,N_20813);
or U22252 (N_22252,N_20420,N_20009);
nor U22253 (N_22253,N_20436,N_20022);
and U22254 (N_22254,N_21132,N_20648);
nor U22255 (N_22255,N_20881,N_20475);
or U22256 (N_22256,N_20372,N_20416);
xor U22257 (N_22257,N_20459,N_20613);
xor U22258 (N_22258,N_20165,N_20791);
nor U22259 (N_22259,N_20033,N_20255);
nor U22260 (N_22260,N_20013,N_21206);
nor U22261 (N_22261,N_21070,N_20486);
and U22262 (N_22262,N_20623,N_21000);
xnor U22263 (N_22263,N_20917,N_20113);
nand U22264 (N_22264,N_20711,N_21082);
nand U22265 (N_22265,N_21209,N_20938);
or U22266 (N_22266,N_20110,N_20631);
and U22267 (N_22267,N_20936,N_20836);
nor U22268 (N_22268,N_20548,N_20554);
or U22269 (N_22269,N_20612,N_20850);
nand U22270 (N_22270,N_20059,N_20696);
or U22271 (N_22271,N_20356,N_21034);
xor U22272 (N_22272,N_20607,N_21192);
and U22273 (N_22273,N_20054,N_20441);
nor U22274 (N_22274,N_20713,N_20612);
xor U22275 (N_22275,N_21090,N_21147);
nand U22276 (N_22276,N_20077,N_20321);
and U22277 (N_22277,N_20256,N_20841);
nor U22278 (N_22278,N_20675,N_20277);
and U22279 (N_22279,N_21124,N_21014);
or U22280 (N_22280,N_20610,N_20839);
nor U22281 (N_22281,N_20486,N_20883);
and U22282 (N_22282,N_20579,N_20260);
nor U22283 (N_22283,N_20061,N_21041);
or U22284 (N_22284,N_20040,N_20102);
xnor U22285 (N_22285,N_20664,N_20982);
and U22286 (N_22286,N_21110,N_20950);
or U22287 (N_22287,N_20308,N_20688);
nor U22288 (N_22288,N_21174,N_21109);
nand U22289 (N_22289,N_20956,N_20354);
nand U22290 (N_22290,N_20878,N_20407);
and U22291 (N_22291,N_20925,N_20867);
xor U22292 (N_22292,N_21241,N_20759);
xor U22293 (N_22293,N_20532,N_20587);
or U22294 (N_22294,N_20062,N_20628);
and U22295 (N_22295,N_20973,N_20672);
nand U22296 (N_22296,N_20924,N_20591);
and U22297 (N_22297,N_20761,N_20522);
xnor U22298 (N_22298,N_20541,N_20132);
nand U22299 (N_22299,N_20052,N_20025);
xnor U22300 (N_22300,N_21247,N_20577);
nand U22301 (N_22301,N_20969,N_21067);
and U22302 (N_22302,N_20294,N_20460);
xnor U22303 (N_22303,N_20926,N_20929);
xnor U22304 (N_22304,N_20666,N_20341);
or U22305 (N_22305,N_20782,N_20950);
and U22306 (N_22306,N_21166,N_20541);
or U22307 (N_22307,N_20438,N_20989);
xnor U22308 (N_22308,N_20309,N_21066);
and U22309 (N_22309,N_20136,N_20094);
xor U22310 (N_22310,N_20747,N_20995);
or U22311 (N_22311,N_20106,N_21149);
nand U22312 (N_22312,N_20645,N_20731);
nor U22313 (N_22313,N_20877,N_20750);
nand U22314 (N_22314,N_20393,N_20903);
and U22315 (N_22315,N_20060,N_20387);
xnor U22316 (N_22316,N_20084,N_20840);
nand U22317 (N_22317,N_20225,N_20698);
and U22318 (N_22318,N_20796,N_21082);
xnor U22319 (N_22319,N_21141,N_20248);
xnor U22320 (N_22320,N_21070,N_20201);
or U22321 (N_22321,N_20856,N_20046);
xor U22322 (N_22322,N_20972,N_20843);
nor U22323 (N_22323,N_20121,N_20320);
nor U22324 (N_22324,N_20249,N_20194);
and U22325 (N_22325,N_21201,N_20897);
nand U22326 (N_22326,N_20575,N_20361);
or U22327 (N_22327,N_21158,N_20070);
or U22328 (N_22328,N_20674,N_20436);
or U22329 (N_22329,N_20816,N_21044);
xor U22330 (N_22330,N_20715,N_21150);
nand U22331 (N_22331,N_21167,N_20259);
nand U22332 (N_22332,N_21162,N_20664);
nor U22333 (N_22333,N_20448,N_20974);
nor U22334 (N_22334,N_20363,N_20562);
and U22335 (N_22335,N_20620,N_20015);
or U22336 (N_22336,N_20536,N_20333);
nor U22337 (N_22337,N_20783,N_20768);
nor U22338 (N_22338,N_20880,N_20526);
nor U22339 (N_22339,N_20602,N_21248);
nand U22340 (N_22340,N_20456,N_20207);
nand U22341 (N_22341,N_21179,N_20644);
or U22342 (N_22342,N_21144,N_20684);
nor U22343 (N_22343,N_20481,N_21231);
nand U22344 (N_22344,N_20344,N_20601);
xor U22345 (N_22345,N_20454,N_20489);
nand U22346 (N_22346,N_20705,N_20580);
or U22347 (N_22347,N_20438,N_20483);
nand U22348 (N_22348,N_20104,N_20038);
or U22349 (N_22349,N_20084,N_21124);
and U22350 (N_22350,N_20765,N_20559);
nor U22351 (N_22351,N_20365,N_20800);
nand U22352 (N_22352,N_21086,N_20211);
or U22353 (N_22353,N_20645,N_20540);
xor U22354 (N_22354,N_20603,N_20106);
or U22355 (N_22355,N_21056,N_20021);
and U22356 (N_22356,N_20859,N_20992);
nor U22357 (N_22357,N_20424,N_20786);
xnor U22358 (N_22358,N_20165,N_20824);
and U22359 (N_22359,N_20452,N_21099);
or U22360 (N_22360,N_20066,N_20271);
nor U22361 (N_22361,N_20954,N_20173);
nand U22362 (N_22362,N_20930,N_20147);
nor U22363 (N_22363,N_20031,N_20983);
and U22364 (N_22364,N_20540,N_20036);
nor U22365 (N_22365,N_21234,N_20572);
nor U22366 (N_22366,N_21053,N_20047);
nand U22367 (N_22367,N_21228,N_20013);
nand U22368 (N_22368,N_20748,N_20978);
nor U22369 (N_22369,N_20649,N_21220);
xor U22370 (N_22370,N_20410,N_20379);
nor U22371 (N_22371,N_20231,N_20085);
nor U22372 (N_22372,N_20716,N_21182);
and U22373 (N_22373,N_21026,N_20361);
and U22374 (N_22374,N_20420,N_20045);
nand U22375 (N_22375,N_21059,N_21021);
xnor U22376 (N_22376,N_20350,N_20461);
nand U22377 (N_22377,N_20988,N_20950);
xor U22378 (N_22378,N_21049,N_21228);
and U22379 (N_22379,N_20039,N_20889);
and U22380 (N_22380,N_21140,N_20852);
or U22381 (N_22381,N_20298,N_20083);
and U22382 (N_22382,N_20646,N_20420);
nor U22383 (N_22383,N_20000,N_20551);
xor U22384 (N_22384,N_20833,N_20182);
and U22385 (N_22385,N_21225,N_20579);
or U22386 (N_22386,N_20692,N_20724);
nand U22387 (N_22387,N_21057,N_20277);
nor U22388 (N_22388,N_20810,N_21239);
xor U22389 (N_22389,N_20409,N_20056);
and U22390 (N_22390,N_20736,N_20835);
and U22391 (N_22391,N_20550,N_20921);
and U22392 (N_22392,N_20733,N_20580);
nor U22393 (N_22393,N_20091,N_21030);
or U22394 (N_22394,N_20509,N_20338);
or U22395 (N_22395,N_20917,N_20653);
nor U22396 (N_22396,N_20556,N_20854);
nor U22397 (N_22397,N_20906,N_21225);
xor U22398 (N_22398,N_20834,N_20518);
nand U22399 (N_22399,N_20149,N_20811);
nor U22400 (N_22400,N_21054,N_20615);
nand U22401 (N_22401,N_21005,N_20368);
nand U22402 (N_22402,N_21138,N_20486);
nor U22403 (N_22403,N_20847,N_20825);
nor U22404 (N_22404,N_20708,N_20650);
xor U22405 (N_22405,N_20898,N_20096);
or U22406 (N_22406,N_20946,N_20250);
nand U22407 (N_22407,N_20981,N_20776);
nand U22408 (N_22408,N_20884,N_20016);
or U22409 (N_22409,N_20521,N_20782);
or U22410 (N_22410,N_20061,N_21073);
xor U22411 (N_22411,N_20283,N_20285);
and U22412 (N_22412,N_21200,N_20948);
and U22413 (N_22413,N_21053,N_20881);
nor U22414 (N_22414,N_20541,N_20237);
or U22415 (N_22415,N_20777,N_20594);
nand U22416 (N_22416,N_20144,N_20807);
nand U22417 (N_22417,N_21109,N_20867);
nand U22418 (N_22418,N_21168,N_20759);
or U22419 (N_22419,N_20253,N_20832);
or U22420 (N_22420,N_21058,N_20564);
nor U22421 (N_22421,N_20697,N_21135);
nand U22422 (N_22422,N_21019,N_21024);
or U22423 (N_22423,N_20465,N_20751);
xor U22424 (N_22424,N_20283,N_21046);
nand U22425 (N_22425,N_20797,N_20477);
nand U22426 (N_22426,N_20556,N_20182);
nor U22427 (N_22427,N_21240,N_20101);
xor U22428 (N_22428,N_20572,N_21040);
or U22429 (N_22429,N_20240,N_20999);
nand U22430 (N_22430,N_21171,N_21218);
xor U22431 (N_22431,N_20246,N_20825);
and U22432 (N_22432,N_20602,N_20898);
and U22433 (N_22433,N_20001,N_20451);
nor U22434 (N_22434,N_21211,N_21203);
and U22435 (N_22435,N_20773,N_20373);
or U22436 (N_22436,N_20677,N_20810);
nand U22437 (N_22437,N_20666,N_21111);
and U22438 (N_22438,N_20441,N_20433);
and U22439 (N_22439,N_20506,N_20515);
or U22440 (N_22440,N_20892,N_20559);
nor U22441 (N_22441,N_20668,N_20321);
and U22442 (N_22442,N_20033,N_20264);
xnor U22443 (N_22443,N_21245,N_21106);
or U22444 (N_22444,N_20003,N_20454);
or U22445 (N_22445,N_20983,N_20931);
and U22446 (N_22446,N_21232,N_20448);
nand U22447 (N_22447,N_20338,N_20899);
and U22448 (N_22448,N_20458,N_21244);
xnor U22449 (N_22449,N_20391,N_20586);
or U22450 (N_22450,N_20585,N_21059);
or U22451 (N_22451,N_20411,N_20458);
or U22452 (N_22452,N_21052,N_20707);
and U22453 (N_22453,N_20885,N_20985);
nand U22454 (N_22454,N_20281,N_20348);
and U22455 (N_22455,N_21237,N_21109);
or U22456 (N_22456,N_20953,N_20355);
nand U22457 (N_22457,N_20098,N_20095);
and U22458 (N_22458,N_20550,N_20993);
nand U22459 (N_22459,N_20288,N_20517);
and U22460 (N_22460,N_20279,N_20647);
nand U22461 (N_22461,N_20594,N_20154);
nor U22462 (N_22462,N_20689,N_20945);
nand U22463 (N_22463,N_21150,N_21213);
or U22464 (N_22464,N_20228,N_21133);
or U22465 (N_22465,N_20954,N_20857);
nor U22466 (N_22466,N_21133,N_21061);
and U22467 (N_22467,N_20528,N_20448);
xnor U22468 (N_22468,N_20187,N_20624);
nand U22469 (N_22469,N_21032,N_20812);
nor U22470 (N_22470,N_21172,N_21235);
nand U22471 (N_22471,N_20510,N_20004);
nand U22472 (N_22472,N_20856,N_21116);
xor U22473 (N_22473,N_20705,N_20312);
nor U22474 (N_22474,N_21038,N_20624);
xor U22475 (N_22475,N_20848,N_20448);
or U22476 (N_22476,N_20527,N_20044);
or U22477 (N_22477,N_20873,N_20443);
or U22478 (N_22478,N_20020,N_20624);
and U22479 (N_22479,N_20570,N_20120);
and U22480 (N_22480,N_20975,N_20625);
nand U22481 (N_22481,N_20901,N_20610);
or U22482 (N_22482,N_20073,N_21106);
nor U22483 (N_22483,N_20099,N_20678);
and U22484 (N_22484,N_20914,N_20692);
and U22485 (N_22485,N_20695,N_20583);
nor U22486 (N_22486,N_20153,N_20336);
nand U22487 (N_22487,N_20459,N_20578);
nand U22488 (N_22488,N_20365,N_20086);
nor U22489 (N_22489,N_20583,N_20957);
nand U22490 (N_22490,N_20186,N_20200);
xnor U22491 (N_22491,N_21178,N_20505);
xnor U22492 (N_22492,N_20652,N_20425);
or U22493 (N_22493,N_20056,N_21114);
xnor U22494 (N_22494,N_20741,N_20009);
and U22495 (N_22495,N_20475,N_20106);
or U22496 (N_22496,N_20129,N_21119);
nor U22497 (N_22497,N_20821,N_20136);
nand U22498 (N_22498,N_20727,N_20552);
or U22499 (N_22499,N_20302,N_20963);
and U22500 (N_22500,N_21812,N_21870);
and U22501 (N_22501,N_21409,N_21810);
xnor U22502 (N_22502,N_21802,N_21835);
nand U22503 (N_22503,N_21291,N_21990);
or U22504 (N_22504,N_21253,N_22337);
and U22505 (N_22505,N_21633,N_21745);
nor U22506 (N_22506,N_21662,N_22125);
nand U22507 (N_22507,N_21906,N_22017);
and U22508 (N_22508,N_22084,N_21814);
nor U22509 (N_22509,N_21735,N_21374);
or U22510 (N_22510,N_22474,N_21577);
xnor U22511 (N_22511,N_21665,N_21534);
or U22512 (N_22512,N_22422,N_21561);
nor U22513 (N_22513,N_21329,N_21889);
xnor U22514 (N_22514,N_22215,N_21498);
nor U22515 (N_22515,N_22134,N_21296);
nor U22516 (N_22516,N_22245,N_21258);
nor U22517 (N_22517,N_22317,N_21923);
xor U22518 (N_22518,N_21618,N_21920);
nand U22519 (N_22519,N_22008,N_21953);
and U22520 (N_22520,N_21940,N_21685);
or U22521 (N_22521,N_21673,N_21469);
nand U22522 (N_22522,N_22114,N_21670);
xnor U22523 (N_22523,N_21638,N_22123);
nor U22524 (N_22524,N_22265,N_21384);
nor U22525 (N_22525,N_21493,N_21679);
nand U22526 (N_22526,N_22316,N_21407);
xor U22527 (N_22527,N_22395,N_21734);
nor U22528 (N_22528,N_22392,N_21857);
xnor U22529 (N_22529,N_22381,N_22147);
or U22530 (N_22530,N_21448,N_21731);
nand U22531 (N_22531,N_21402,N_22361);
xor U22532 (N_22532,N_22441,N_22448);
or U22533 (N_22533,N_21737,N_21915);
or U22534 (N_22534,N_21369,N_21982);
nand U22535 (N_22535,N_22351,N_21925);
nand U22536 (N_22536,N_22176,N_22193);
nand U22537 (N_22537,N_21688,N_21471);
nor U22538 (N_22538,N_22075,N_22177);
nand U22539 (N_22539,N_21437,N_21256);
nor U22540 (N_22540,N_22210,N_21758);
and U22541 (N_22541,N_21749,N_22168);
and U22542 (N_22542,N_21455,N_21529);
nor U22543 (N_22543,N_22179,N_21309);
xnor U22544 (N_22544,N_22314,N_22077);
and U22545 (N_22545,N_21317,N_21397);
or U22546 (N_22546,N_22399,N_22110);
and U22547 (N_22547,N_21949,N_22431);
nand U22548 (N_22548,N_22266,N_21672);
nor U22549 (N_22549,N_21339,N_22243);
nor U22550 (N_22550,N_22459,N_21261);
xor U22551 (N_22551,N_21525,N_22439);
nor U22552 (N_22552,N_22409,N_21739);
nand U22553 (N_22553,N_21605,N_21974);
or U22554 (N_22554,N_21817,N_22447);
xor U22555 (N_22555,N_22228,N_21929);
nor U22556 (N_22556,N_21349,N_22246);
and U22557 (N_22557,N_22032,N_22241);
nor U22558 (N_22558,N_21487,N_21364);
xnor U22559 (N_22559,N_22031,N_21599);
nor U22560 (N_22560,N_21410,N_21896);
nor U22561 (N_22561,N_22423,N_21403);
or U22562 (N_22562,N_21547,N_21546);
and U22563 (N_22563,N_21632,N_21959);
nor U22564 (N_22564,N_21716,N_21341);
nor U22565 (N_22565,N_22052,N_21474);
and U22566 (N_22566,N_21483,N_22343);
xor U22567 (N_22567,N_22277,N_21993);
and U22568 (N_22568,N_21729,N_21967);
nor U22569 (N_22569,N_21895,N_22222);
and U22570 (N_22570,N_21962,N_21771);
xnor U22571 (N_22571,N_21821,N_22238);
or U22572 (N_22572,N_22479,N_21634);
xor U22573 (N_22573,N_22461,N_22309);
nor U22574 (N_22574,N_22234,N_21502);
nand U22575 (N_22575,N_21572,N_21690);
and U22576 (N_22576,N_21352,N_22132);
and U22577 (N_22577,N_22372,N_21921);
xor U22578 (N_22578,N_21666,N_22319);
nor U22579 (N_22579,N_22019,N_21645);
nand U22580 (N_22580,N_22371,N_21726);
and U22581 (N_22581,N_21418,N_22034);
or U22582 (N_22582,N_21894,N_21926);
xnor U22583 (N_22583,N_22041,N_21357);
nor U22584 (N_22584,N_22208,N_21548);
nand U22585 (N_22585,N_22364,N_22021);
xnor U22586 (N_22586,N_22185,N_21543);
nor U22587 (N_22587,N_21527,N_22435);
or U22588 (N_22588,N_22023,N_22213);
and U22589 (N_22589,N_21890,N_22487);
nand U22590 (N_22590,N_22236,N_21678);
nor U22591 (N_22591,N_22252,N_22494);
xnor U22592 (N_22592,N_22336,N_22360);
nand U22593 (N_22593,N_22492,N_22264);
xnor U22594 (N_22594,N_21664,N_22088);
or U22595 (N_22595,N_22211,N_21520);
and U22596 (N_22596,N_21887,N_21311);
or U22597 (N_22597,N_22156,N_22359);
xor U22598 (N_22598,N_21683,N_21554);
nand U22599 (N_22599,N_22338,N_21540);
and U22600 (N_22600,N_21533,N_21293);
or U22601 (N_22601,N_21934,N_21280);
or U22602 (N_22602,N_21303,N_22477);
or U22603 (N_22603,N_22167,N_21558);
and U22604 (N_22604,N_22128,N_21278);
or U22605 (N_22605,N_22036,N_21837);
xnor U22606 (N_22606,N_21438,N_22289);
nand U22607 (N_22607,N_21732,N_22254);
nor U22608 (N_22608,N_21935,N_21715);
or U22609 (N_22609,N_21500,N_21452);
nand U22610 (N_22610,N_21700,N_22257);
nand U22611 (N_22611,N_22443,N_22226);
xor U22612 (N_22612,N_22383,N_21963);
xnor U22613 (N_22613,N_21893,N_22356);
nand U22614 (N_22614,N_22182,N_21697);
xor U22615 (N_22615,N_21326,N_21375);
or U22616 (N_22616,N_22432,N_22282);
nor U22617 (N_22617,N_22051,N_21754);
or U22618 (N_22618,N_21299,N_22109);
nor U22619 (N_22619,N_21612,N_21508);
and U22620 (N_22620,N_22293,N_21456);
nand U22621 (N_22621,N_21382,N_21691);
or U22622 (N_22622,N_21760,N_21839);
or U22623 (N_22623,N_22380,N_21408);
or U22624 (N_22624,N_22410,N_22046);
and U22625 (N_22625,N_21616,N_21955);
or U22626 (N_22626,N_22229,N_22368);
nor U22627 (N_22627,N_21902,N_22239);
or U22628 (N_22628,N_22199,N_21914);
or U22629 (N_22629,N_21578,N_21968);
nor U22630 (N_22630,N_21701,N_21260);
or U22631 (N_22631,N_22348,N_21722);
nor U22632 (N_22632,N_21328,N_22442);
or U22633 (N_22633,N_21304,N_22152);
and U22634 (N_22634,N_21900,N_21947);
or U22635 (N_22635,N_21601,N_21782);
xnor U22636 (N_22636,N_21689,N_22205);
and U22637 (N_22637,N_21386,N_22398);
xnor U22638 (N_22638,N_22404,N_21800);
nor U22639 (N_22639,N_21453,N_22022);
nor U22640 (N_22640,N_21724,N_22452);
and U22641 (N_22641,N_22318,N_21593);
and U22642 (N_22642,N_21987,N_22158);
and U22643 (N_22643,N_21985,N_21830);
nand U22644 (N_22644,N_21342,N_22366);
nand U22645 (N_22645,N_21322,N_21343);
and U22646 (N_22646,N_22406,N_22064);
and U22647 (N_22647,N_21553,N_21769);
nor U22648 (N_22648,N_22073,N_21770);
or U22649 (N_22649,N_21806,N_22043);
and U22650 (N_22650,N_22030,N_21294);
or U22651 (N_22651,N_21706,N_21551);
nand U22652 (N_22652,N_21852,N_22137);
xnor U22653 (N_22653,N_21766,N_21415);
nor U22654 (N_22654,N_21517,N_22172);
nor U22655 (N_22655,N_21399,N_22071);
and U22656 (N_22656,N_21753,N_21658);
and U22657 (N_22657,N_21711,N_21834);
and U22658 (N_22658,N_22148,N_21305);
or U22659 (N_22659,N_21798,N_21521);
nand U22660 (N_22660,N_21287,N_22163);
or U22661 (N_22661,N_21995,N_21492);
nand U22662 (N_22662,N_21905,N_21536);
and U22663 (N_22663,N_21478,N_22292);
and U22664 (N_22664,N_21392,N_21752);
nand U22665 (N_22665,N_21602,N_22278);
nor U22666 (N_22666,N_22445,N_21587);
nor U22667 (N_22667,N_21930,N_21466);
and U22668 (N_22668,N_21768,N_21477);
xor U22669 (N_22669,N_22072,N_22397);
nor U22670 (N_22670,N_22263,N_22499);
nand U22671 (N_22671,N_22207,N_21432);
nor U22672 (N_22672,N_21489,N_22391);
and U22673 (N_22673,N_21820,N_21333);
nor U22674 (N_22674,N_22027,N_21838);
or U22675 (N_22675,N_21285,N_21986);
nand U22676 (N_22676,N_21796,N_22183);
or U22677 (N_22677,N_22294,N_22290);
and U22678 (N_22678,N_22054,N_21370);
and U22679 (N_22679,N_21791,N_22061);
and U22680 (N_22680,N_22029,N_21494);
xor U22681 (N_22681,N_22175,N_21473);
xnor U22682 (N_22682,N_21832,N_22298);
or U22683 (N_22683,N_22483,N_22272);
nor U22684 (N_22684,N_21289,N_21956);
nand U22685 (N_22685,N_21516,N_21822);
nor U22686 (N_22686,N_21348,N_21526);
nand U22687 (N_22687,N_22198,N_22260);
nor U22688 (N_22688,N_21610,N_22416);
and U22689 (N_22689,N_21876,N_22214);
xor U22690 (N_22690,N_21366,N_22322);
and U22691 (N_22691,N_21899,N_22446);
nor U22692 (N_22692,N_22345,N_21863);
or U22693 (N_22693,N_21625,N_22157);
or U22694 (N_22694,N_21695,N_22330);
xnor U22695 (N_22695,N_22310,N_22066);
or U22696 (N_22696,N_22341,N_21396);
or U22697 (N_22697,N_21686,N_22120);
nand U22698 (N_22698,N_22186,N_22151);
and U22699 (N_22699,N_21831,N_22413);
nand U22700 (N_22700,N_22115,N_21552);
nor U22701 (N_22701,N_21480,N_21594);
and U22702 (N_22702,N_21428,N_21564);
nor U22703 (N_22703,N_21450,N_21510);
nand U22704 (N_22704,N_22408,N_22411);
and U22705 (N_22705,N_21479,N_22387);
or U22706 (N_22706,N_22324,N_22333);
nand U22707 (N_22707,N_22457,N_22015);
nand U22708 (N_22708,N_21816,N_21845);
nand U22709 (N_22709,N_21266,N_21394);
xor U22710 (N_22710,N_22108,N_21677);
nand U22711 (N_22711,N_21515,N_21585);
nand U22712 (N_22712,N_21747,N_22011);
nor U22713 (N_22713,N_21661,N_21624);
and U22714 (N_22714,N_21530,N_21542);
nand U22715 (N_22715,N_21354,N_21524);
nor U22716 (N_22716,N_22419,N_21776);
xor U22717 (N_22717,N_22393,N_21998);
xnor U22718 (N_22718,N_22468,N_21576);
or U22719 (N_22719,N_21292,N_21254);
nor U22720 (N_22720,N_21641,N_22386);
xor U22721 (N_22721,N_21829,N_22057);
nor U22722 (N_22722,N_21644,N_21416);
xnor U22723 (N_22723,N_22217,N_21522);
and U22724 (N_22724,N_22065,N_21999);
nand U22725 (N_22725,N_22189,N_21808);
or U22726 (N_22726,N_22178,N_22480);
and U22727 (N_22727,N_22143,N_22276);
nor U22728 (N_22728,N_22074,N_21581);
xnor U22729 (N_22729,N_21579,N_21325);
and U22730 (N_22730,N_21847,N_22112);
nor U22731 (N_22731,N_21908,N_22369);
or U22732 (N_22732,N_22003,N_21560);
and U22733 (N_22733,N_21273,N_21582);
xnor U22734 (N_22734,N_21262,N_21475);
xnor U22735 (N_22735,N_22047,N_21388);
and U22736 (N_22736,N_21545,N_21751);
or U22737 (N_22737,N_21848,N_21775);
nor U22738 (N_22738,N_22083,N_21781);
nand U22739 (N_22739,N_21295,N_22303);
and U22740 (N_22740,N_21763,N_21746);
xnor U22741 (N_22741,N_21575,N_22300);
nand U22742 (N_22742,N_22042,N_21608);
and U22743 (N_22743,N_21767,N_21503);
and U22744 (N_22744,N_22235,N_21843);
or U22745 (N_22745,N_21809,N_22327);
and U22746 (N_22746,N_22164,N_22230);
and U22747 (N_22747,N_22321,N_21795);
nand U22748 (N_22748,N_21713,N_21321);
or U22749 (N_22749,N_21338,N_22104);
or U22750 (N_22750,N_21482,N_21360);
or U22751 (N_22751,N_21302,N_22069);
xnor U22752 (N_22752,N_21652,N_21785);
or U22753 (N_22753,N_22224,N_22142);
nand U22754 (N_22754,N_22297,N_21933);
nor U22755 (N_22755,N_22204,N_21372);
or U22756 (N_22756,N_21756,N_22286);
nor U22757 (N_22757,N_21460,N_21660);
xor U22758 (N_22758,N_21977,N_22390);
nand U22759 (N_22759,N_21653,N_22091);
and U22760 (N_22760,N_22497,N_22203);
xor U22761 (N_22761,N_21353,N_22382);
and U22762 (N_22762,N_21362,N_22059);
xnor U22763 (N_22763,N_22180,N_22472);
nor U22764 (N_22764,N_21301,N_22133);
or U22765 (N_22765,N_22420,N_21481);
xor U22766 (N_22766,N_22296,N_21907);
nand U22767 (N_22767,N_22216,N_21306);
or U22768 (N_22768,N_21316,N_21345);
and U22769 (N_22769,N_21710,N_21764);
nor U22770 (N_22770,N_21513,N_21454);
nor U22771 (N_22771,N_22259,N_21903);
nand U22772 (N_22772,N_22449,N_21844);
and U22773 (N_22773,N_22450,N_21854);
or U22774 (N_22774,N_21412,N_22020);
nor U22775 (N_22775,N_21314,N_21356);
or U22776 (N_22776,N_21346,N_21656);
nand U22777 (N_22777,N_21331,N_21406);
nor U22778 (N_22778,N_21787,N_21320);
and U22779 (N_22779,N_21901,N_21580);
nand U22780 (N_22780,N_22190,N_22090);
nor U22781 (N_22781,N_22375,N_22040);
and U22782 (N_22782,N_22130,N_22106);
nand U22783 (N_22783,N_22462,N_21988);
xnor U22784 (N_22784,N_22365,N_21523);
nand U22785 (N_22785,N_21367,N_21468);
and U22786 (N_22786,N_21390,N_22103);
xnor U22787 (N_22787,N_21417,N_22427);
xnor U22788 (N_22788,N_22227,N_21420);
and U22789 (N_22789,N_22295,N_21978);
nand U22790 (N_22790,N_21877,N_21431);
xor U22791 (N_22791,N_22223,N_21850);
nand U22792 (N_22792,N_22454,N_21441);
nand U22793 (N_22793,N_21404,N_21668);
or U22794 (N_22794,N_22135,N_22247);
nor U22795 (N_22795,N_21574,N_22326);
and U22796 (N_22796,N_21627,N_22006);
nor U22797 (N_22797,N_22484,N_22490);
nand U22798 (N_22798,N_22433,N_21436);
nand U22799 (N_22799,N_21922,N_21840);
and U22800 (N_22800,N_21675,N_22153);
xor U22801 (N_22801,N_21337,N_21405);
and U22802 (N_22802,N_21755,N_21620);
xnor U22803 (N_22803,N_21797,N_21430);
or U22804 (N_22804,N_21784,N_21259);
nor U22805 (N_22805,N_21556,N_21937);
and U22806 (N_22806,N_21853,N_22038);
and U22807 (N_22807,N_22225,N_21954);
or U22808 (N_22808,N_21957,N_21344);
or U22809 (N_22809,N_22187,N_21598);
or U22810 (N_22810,N_21472,N_21702);
xnor U22811 (N_22811,N_22181,N_21932);
nor U22812 (N_22812,N_22424,N_21590);
xor U22813 (N_22813,N_21931,N_21461);
nor U22814 (N_22814,N_21698,N_21445);
nand U22815 (N_22815,N_22160,N_22473);
and U22816 (N_22816,N_22232,N_21970);
or U22817 (N_22817,N_22437,N_21973);
xor U22818 (N_22818,N_21310,N_21757);
xnor U22819 (N_22819,N_21861,N_21569);
and U22820 (N_22820,N_21421,N_21786);
nand U22821 (N_22821,N_21308,N_21792);
nor U22822 (N_22822,N_21819,N_21506);
and U22823 (N_22823,N_22460,N_21823);
or U22824 (N_22824,N_22358,N_22078);
nand U22825 (N_22825,N_21825,N_21692);
nand U22826 (N_22826,N_21950,N_21457);
and U22827 (N_22827,N_21267,N_21635);
and U22828 (N_22828,N_22354,N_21484);
nand U22829 (N_22829,N_22414,N_21811);
nand U22830 (N_22830,N_21693,N_21413);
xnor U22831 (N_22831,N_22488,N_21570);
xor U22832 (N_22832,N_21671,N_22304);
and U22833 (N_22833,N_21426,N_21712);
nor U22834 (N_22834,N_22161,N_21268);
and U22835 (N_22835,N_21676,N_22093);
nand U22836 (N_22836,N_21912,N_21774);
or U22837 (N_22837,N_21788,N_22016);
xor U22838 (N_22838,N_22403,N_22220);
xnor U22839 (N_22839,N_21714,N_21687);
nand U22840 (N_22840,N_22146,N_22346);
and U22841 (N_22841,N_22384,N_21257);
and U22842 (N_22842,N_21433,N_21879);
xor U22843 (N_22843,N_21836,N_21589);
or U22844 (N_22844,N_21497,N_21741);
or U22845 (N_22845,N_22325,N_22010);
nor U22846 (N_22846,N_22258,N_21762);
and U22847 (N_22847,N_22089,N_21277);
nand U22848 (N_22848,N_22094,N_21748);
or U22849 (N_22849,N_21365,N_22287);
xnor U22850 (N_22850,N_22116,N_21884);
nor U22851 (N_22851,N_21470,N_21462);
nand U22852 (N_22852,N_22056,N_21860);
or U22853 (N_22853,N_21419,N_22050);
xor U22854 (N_22854,N_21319,N_22126);
or U22855 (N_22855,N_21980,N_22063);
nor U22856 (N_22856,N_21779,N_22444);
or U22857 (N_22857,N_21379,N_22139);
xor U22858 (N_22858,N_21491,N_22253);
xor U22859 (N_22859,N_22305,N_22035);
xnor U22860 (N_22860,N_21898,N_21703);
and U22861 (N_22861,N_22212,N_21380);
nor U22862 (N_22862,N_21655,N_22458);
nor U22863 (N_22863,N_22113,N_22470);
nand U22864 (N_22864,N_22350,N_22430);
xnor U22865 (N_22865,N_22005,N_21359);
nand U22866 (N_22866,N_21272,N_21640);
and U22867 (N_22867,N_22053,N_22194);
or U22868 (N_22868,N_22012,N_21916);
nand U22869 (N_22869,N_21946,N_21401);
nand U22870 (N_22870,N_22367,N_22170);
nand U22871 (N_22871,N_21965,N_21709);
or U22872 (N_22872,N_21532,N_21743);
nor U22873 (N_22873,N_22291,N_21892);
nand U22874 (N_22874,N_21674,N_22357);
xnor U22875 (N_22875,N_21571,N_21911);
or U22876 (N_22876,N_22024,N_21793);
nand U22877 (N_22877,N_21750,N_22136);
nor U22878 (N_22878,N_21778,N_22100);
nor U22879 (N_22879,N_21442,N_21623);
and U22880 (N_22880,N_21443,N_22482);
nand U22881 (N_22881,N_21867,N_22376);
xor U22882 (N_22882,N_21376,N_22082);
and U22883 (N_22883,N_22481,N_21592);
xor U22884 (N_22884,N_21476,N_21684);
nor U22885 (N_22885,N_22493,N_21424);
or U22886 (N_22886,N_21727,N_21288);
or U22887 (N_22887,N_22173,N_22284);
and U22888 (N_22888,N_21393,N_21423);
nand U22889 (N_22889,N_22440,N_21621);
or U22890 (N_22890,N_22080,N_21567);
xnor U22891 (N_22891,N_22248,N_21917);
nor U22892 (N_22892,N_22119,N_21596);
nor U22893 (N_22893,N_21391,N_22149);
or U22894 (N_22894,N_21449,N_21340);
nor U22895 (N_22895,N_22251,N_22313);
nor U22896 (N_22896,N_21518,N_22412);
nand U22897 (N_22897,N_22340,N_22067);
or U22898 (N_22898,N_21613,N_22344);
and U22899 (N_22899,N_21351,N_21603);
nor U22900 (N_22900,N_22013,N_21972);
xor U22901 (N_22901,N_21948,N_22465);
nand U22902 (N_22902,N_21439,N_21313);
or U22903 (N_22903,N_21960,N_22328);
xnor U22904 (N_22904,N_21429,N_22107);
and U22905 (N_22905,N_22092,N_22044);
nand U22906 (N_22906,N_22274,N_21389);
or U22907 (N_22907,N_21446,N_21467);
and U22908 (N_22908,N_22200,N_21614);
and U22909 (N_22909,N_21385,N_22261);
nor U22910 (N_22910,N_22415,N_21654);
or U22911 (N_22911,N_21519,N_21856);
nand U22912 (N_22912,N_22456,N_21334);
xnor U22913 (N_22913,N_21447,N_22355);
or U22914 (N_22914,N_22288,N_22018);
xor U22915 (N_22915,N_22396,N_22209);
xor U22916 (N_22916,N_22374,N_22273);
and U22917 (N_22917,N_22425,N_22202);
or U22918 (N_22918,N_22055,N_21794);
nor U22919 (N_22919,N_21958,N_22122);
nand U22920 (N_22920,N_21490,N_22159);
and U22921 (N_22921,N_22102,N_21680);
or U22922 (N_22922,N_22280,N_22138);
xor U22923 (N_22923,N_21913,N_21381);
nor U22924 (N_22924,N_21263,N_22192);
nor U22925 (N_22925,N_22485,N_22062);
xor U22926 (N_22926,N_21704,N_22049);
or U22927 (N_22927,N_21643,N_22184);
or U22928 (N_22928,N_22169,N_21528);
xor U22929 (N_22929,N_21550,N_21881);
or U22930 (N_22930,N_22155,N_21855);
or U22931 (N_22931,N_22307,N_21777);
and U22932 (N_22932,N_22007,N_21891);
xnor U22933 (N_22933,N_21780,N_21717);
nor U22934 (N_22934,N_21251,N_21992);
xor U22935 (N_22935,N_22096,N_21886);
and U22936 (N_22936,N_21647,N_21505);
nand U22937 (N_22937,N_22377,N_21549);
or U22938 (N_22938,N_22463,N_21807);
nand U22939 (N_22939,N_21979,N_21307);
or U22940 (N_22940,N_22141,N_22476);
xor U22941 (N_22941,N_21789,N_21875);
nand U22942 (N_22942,N_22095,N_21300);
nor U22943 (N_22943,N_21265,N_22400);
xnor U22944 (N_22944,N_22174,N_22453);
and U22945 (N_22945,N_21846,N_22455);
nand U22946 (N_22946,N_21873,N_21813);
nand U22947 (N_22947,N_22352,N_22331);
nor U22948 (N_22948,N_21398,N_22118);
nor U22949 (N_22949,N_22312,N_22166);
nor U22950 (N_22950,N_22275,N_21562);
nand U22951 (N_22951,N_21804,N_22131);
nand U22952 (N_22952,N_22342,N_21286);
or U22953 (N_22953,N_22353,N_21595);
and U22954 (N_22954,N_21639,N_22339);
nor U22955 (N_22955,N_22299,N_21565);
xor U22956 (N_22956,N_21928,N_22249);
and U22957 (N_22957,N_22025,N_21942);
nor U22958 (N_22958,N_21994,N_21951);
or U22959 (N_22959,N_21918,N_21361);
and U22960 (N_22960,N_21862,N_21363);
xor U22961 (N_22961,N_21606,N_21327);
or U22962 (N_22962,N_21961,N_21864);
nand U22963 (N_22963,N_21971,N_21842);
or U22964 (N_22964,N_21607,N_21910);
and U22965 (N_22965,N_21269,N_21435);
or U22966 (N_22966,N_22434,N_21725);
nand U22967 (N_22967,N_22121,N_22467);
nor U22968 (N_22968,N_21719,N_22233);
nand U22969 (N_22969,N_22009,N_22039);
and U22970 (N_22970,N_21504,N_22436);
nor U22971 (N_22971,N_21927,N_22329);
or U22972 (N_22972,N_21966,N_22283);
nand U22973 (N_22973,N_22242,N_21650);
nor U22974 (N_22974,N_21738,N_21588);
nor U22975 (N_22975,N_21969,N_21514);
or U22976 (N_22976,N_21919,N_21411);
nor U22977 (N_22977,N_21874,N_21537);
or U22978 (N_22978,N_21833,N_21274);
or U22979 (N_22979,N_21939,N_21667);
nand U22980 (N_22980,N_21284,N_22349);
and U22981 (N_22981,N_21591,N_21499);
nor U22982 (N_22982,N_21451,N_22262);
nand U22983 (N_22983,N_21945,N_22058);
or U22984 (N_22984,N_21648,N_22335);
xor U22985 (N_22985,N_21859,N_21255);
or U22986 (N_22986,N_21271,N_21646);
nand U22987 (N_22987,N_21312,N_21531);
and U22988 (N_22988,N_22099,N_21600);
or U22989 (N_22989,N_22070,N_22429);
or U22990 (N_22990,N_21721,N_21444);
nand U22991 (N_22991,N_21728,N_21723);
nand U22992 (N_22992,N_22347,N_21742);
or U22993 (N_22993,N_21669,N_22466);
xor U22994 (N_22994,N_21459,N_21651);
xnor U22995 (N_22995,N_21350,N_22281);
nand U22996 (N_22996,N_21872,N_22255);
nand U22997 (N_22997,N_21264,N_21373);
nor U22998 (N_22998,N_21496,N_21324);
and U22999 (N_22999,N_22219,N_21828);
or U23000 (N_23000,N_21279,N_22495);
nand U23001 (N_23001,N_22129,N_21984);
xor U23002 (N_23002,N_21659,N_22270);
and U23003 (N_23003,N_21878,N_21851);
nand U23004 (N_23004,N_21583,N_21622);
and U23005 (N_23005,N_21841,N_21883);
xnor U23006 (N_23006,N_21276,N_22068);
xnor U23007 (N_23007,N_21976,N_22407);
xor U23008 (N_23008,N_22195,N_21885);
xnor U23009 (N_23009,N_21315,N_22271);
nand U23010 (N_23010,N_21283,N_22196);
xor U23011 (N_23011,N_21952,N_21705);
nand U23012 (N_23012,N_22323,N_22206);
and U23013 (N_23013,N_22124,N_22469);
nor U23014 (N_23014,N_21290,N_21297);
or U23015 (N_23015,N_22489,N_21538);
and U23016 (N_23016,N_22218,N_22165);
xor U23017 (N_23017,N_22221,N_22417);
or U23018 (N_23018,N_21630,N_21458);
or U23019 (N_23019,N_22250,N_22379);
nor U23020 (N_23020,N_21378,N_21387);
and U23021 (N_23021,N_21615,N_22478);
nor U23022 (N_23022,N_21604,N_21996);
nand U23023 (N_23023,N_21395,N_22154);
or U23024 (N_23024,N_22048,N_21488);
nand U23025 (N_23025,N_21869,N_21535);
nand U23026 (N_23026,N_22000,N_21941);
nor U23027 (N_23027,N_22111,N_21733);
or U23028 (N_23028,N_21282,N_22098);
or U23029 (N_23029,N_21332,N_22301);
or U23030 (N_23030,N_22498,N_21657);
or U23031 (N_23031,N_22311,N_21335);
nor U23032 (N_23032,N_21636,N_21541);
or U23033 (N_23033,N_22244,N_21740);
or U23034 (N_23034,N_22389,N_21252);
nand U23035 (N_23035,N_22471,N_21539);
nand U23036 (N_23036,N_22127,N_21681);
xnor U23037 (N_23037,N_21501,N_21981);
xor U23038 (N_23038,N_21440,N_22486);
xor U23039 (N_23039,N_21368,N_21663);
nor U23040 (N_23040,N_22426,N_21544);
or U23041 (N_23041,N_21761,N_21465);
nand U23042 (N_23042,N_21975,N_21512);
and U23043 (N_23043,N_21619,N_21559);
and U23044 (N_23044,N_21938,N_22334);
nor U23045 (N_23045,N_22370,N_21347);
nor U23046 (N_23046,N_21699,N_21944);
nand U23047 (N_23047,N_21772,N_22105);
xnor U23048 (N_23048,N_22451,N_22081);
xnor U23049 (N_23049,N_22240,N_21924);
and U23050 (N_23050,N_21318,N_21507);
nand U23051 (N_23051,N_22117,N_21696);
or U23052 (N_23052,N_21485,N_21557);
or U23053 (N_23053,N_22418,N_22385);
nor U23054 (N_23054,N_21708,N_21826);
or U23055 (N_23055,N_21355,N_21815);
and U23056 (N_23056,N_22302,N_21765);
or U23057 (N_23057,N_21991,N_21377);
xor U23058 (N_23058,N_22496,N_21801);
nor U23059 (N_23059,N_22267,N_21434);
nand U23060 (N_23060,N_21936,N_22076);
nand U23061 (N_23061,N_21275,N_21631);
or U23062 (N_23062,N_21868,N_21642);
and U23063 (N_23063,N_22464,N_21904);
and U23064 (N_23064,N_22162,N_22308);
or U23065 (N_23065,N_22197,N_21464);
and U23066 (N_23066,N_22421,N_22004);
nor U23067 (N_23067,N_21358,N_21568);
nand U23068 (N_23068,N_21888,N_22037);
nand U23069 (N_23069,N_21744,N_21849);
nor U23070 (N_23070,N_22279,N_22101);
and U23071 (N_23071,N_21336,N_21720);
or U23072 (N_23072,N_21573,N_21718);
nand U23073 (N_23073,N_21427,N_22401);
or U23074 (N_23074,N_22145,N_21383);
nor U23075 (N_23075,N_21943,N_22256);
nor U23076 (N_23076,N_21989,N_21824);
nand U23077 (N_23077,N_21511,N_22191);
xor U23078 (N_23078,N_22140,N_21250);
xnor U23079 (N_23079,N_21799,N_21773);
nor U23080 (N_23080,N_21425,N_22438);
nand U23081 (N_23081,N_21997,N_21858);
xnor U23082 (N_23082,N_22026,N_22014);
nand U23083 (N_23083,N_22363,N_21694);
xor U23084 (N_23084,N_22001,N_21880);
or U23085 (N_23085,N_22378,N_21298);
or U23086 (N_23086,N_21818,N_22428);
or U23087 (N_23087,N_21486,N_21597);
or U23088 (N_23088,N_22201,N_21783);
and U23089 (N_23089,N_22079,N_21371);
or U23090 (N_23090,N_22405,N_21495);
or U23091 (N_23091,N_22028,N_22306);
and U23092 (N_23092,N_21637,N_21805);
nand U23093 (N_23093,N_22402,N_22237);
xor U23094 (N_23094,N_22144,N_21509);
and U23095 (N_23095,N_21827,N_21865);
xor U23096 (N_23096,N_22002,N_21281);
xnor U23097 (N_23097,N_21629,N_21323);
nor U23098 (N_23098,N_22171,N_21414);
nand U23099 (N_23099,N_21617,N_22097);
or U23100 (N_23100,N_21682,N_22268);
nor U23101 (N_23101,N_21897,N_21555);
nor U23102 (N_23102,N_21563,N_21803);
and U23103 (N_23103,N_21790,N_22060);
and U23104 (N_23104,N_21909,N_21626);
nor U23105 (N_23105,N_21882,N_22231);
or U23106 (N_23106,N_22150,N_22033);
nand U23107 (N_23107,N_21611,N_22320);
nor U23108 (N_23108,N_22394,N_21584);
nor U23109 (N_23109,N_21628,N_22188);
or U23110 (N_23110,N_21964,N_21609);
nand U23111 (N_23111,N_21330,N_22087);
or U23112 (N_23112,N_21983,N_21649);
xnor U23113 (N_23113,N_21736,N_22475);
xnor U23114 (N_23114,N_22388,N_21707);
nand U23115 (N_23115,N_21730,N_22086);
nand U23116 (N_23116,N_21270,N_22045);
or U23117 (N_23117,N_21566,N_21866);
nand U23118 (N_23118,N_21759,N_22373);
and U23119 (N_23119,N_22285,N_21586);
or U23120 (N_23120,N_22332,N_22491);
nor U23121 (N_23121,N_21871,N_21422);
or U23122 (N_23122,N_22315,N_22269);
and U23123 (N_23123,N_21463,N_22362);
nor U23124 (N_23124,N_22085,N_21400);
or U23125 (N_23125,N_21824,N_21747);
and U23126 (N_23126,N_21719,N_21254);
nor U23127 (N_23127,N_21270,N_22348);
and U23128 (N_23128,N_21473,N_22195);
nor U23129 (N_23129,N_21832,N_21875);
nor U23130 (N_23130,N_22475,N_22210);
xor U23131 (N_23131,N_22269,N_22048);
xnor U23132 (N_23132,N_22207,N_21880);
and U23133 (N_23133,N_21800,N_21918);
xor U23134 (N_23134,N_21729,N_21721);
and U23135 (N_23135,N_21534,N_21778);
nor U23136 (N_23136,N_21834,N_21365);
nand U23137 (N_23137,N_22483,N_22107);
or U23138 (N_23138,N_22398,N_22289);
nand U23139 (N_23139,N_22000,N_21669);
xnor U23140 (N_23140,N_22445,N_21451);
and U23141 (N_23141,N_21919,N_21328);
nand U23142 (N_23142,N_21551,N_22465);
nand U23143 (N_23143,N_21781,N_22425);
nand U23144 (N_23144,N_21775,N_21689);
and U23145 (N_23145,N_21875,N_21692);
or U23146 (N_23146,N_22307,N_22192);
nand U23147 (N_23147,N_21953,N_22369);
nor U23148 (N_23148,N_22441,N_21535);
and U23149 (N_23149,N_21326,N_21916);
nand U23150 (N_23150,N_21720,N_22351);
nor U23151 (N_23151,N_22458,N_21922);
xor U23152 (N_23152,N_21943,N_22492);
nor U23153 (N_23153,N_21453,N_22480);
nor U23154 (N_23154,N_22076,N_21986);
or U23155 (N_23155,N_22054,N_21316);
nand U23156 (N_23156,N_21539,N_21965);
nor U23157 (N_23157,N_21544,N_21441);
and U23158 (N_23158,N_21564,N_21326);
nand U23159 (N_23159,N_21444,N_22045);
nand U23160 (N_23160,N_21277,N_22307);
nand U23161 (N_23161,N_21713,N_21868);
and U23162 (N_23162,N_21995,N_21250);
nor U23163 (N_23163,N_22402,N_21962);
or U23164 (N_23164,N_22055,N_22046);
and U23165 (N_23165,N_21958,N_21293);
nand U23166 (N_23166,N_21984,N_22069);
xnor U23167 (N_23167,N_21889,N_21958);
and U23168 (N_23168,N_22228,N_21914);
nand U23169 (N_23169,N_21788,N_22315);
nand U23170 (N_23170,N_22423,N_22175);
nor U23171 (N_23171,N_21930,N_21341);
nand U23172 (N_23172,N_21387,N_21793);
nor U23173 (N_23173,N_22463,N_21985);
and U23174 (N_23174,N_21292,N_21559);
or U23175 (N_23175,N_22252,N_21419);
or U23176 (N_23176,N_22446,N_22249);
or U23177 (N_23177,N_21740,N_22474);
nor U23178 (N_23178,N_22375,N_21425);
or U23179 (N_23179,N_22015,N_22321);
and U23180 (N_23180,N_22445,N_22392);
nor U23181 (N_23181,N_21665,N_22443);
nand U23182 (N_23182,N_21431,N_22294);
nand U23183 (N_23183,N_21384,N_22418);
nand U23184 (N_23184,N_22250,N_22374);
nor U23185 (N_23185,N_22457,N_22263);
or U23186 (N_23186,N_21485,N_22184);
nor U23187 (N_23187,N_21372,N_21415);
and U23188 (N_23188,N_21549,N_21598);
xor U23189 (N_23189,N_21550,N_22092);
nor U23190 (N_23190,N_22296,N_21408);
xor U23191 (N_23191,N_21264,N_22444);
nor U23192 (N_23192,N_21513,N_21539);
or U23193 (N_23193,N_21351,N_21889);
or U23194 (N_23194,N_21451,N_22085);
nand U23195 (N_23195,N_21343,N_21547);
or U23196 (N_23196,N_21829,N_21465);
xnor U23197 (N_23197,N_21839,N_22144);
nand U23198 (N_23198,N_21484,N_22174);
and U23199 (N_23199,N_22421,N_21850);
nor U23200 (N_23200,N_21292,N_21902);
and U23201 (N_23201,N_22154,N_21725);
or U23202 (N_23202,N_22179,N_22283);
xor U23203 (N_23203,N_21257,N_21884);
nor U23204 (N_23204,N_21656,N_21497);
nor U23205 (N_23205,N_21405,N_21486);
xnor U23206 (N_23206,N_21944,N_22446);
and U23207 (N_23207,N_21661,N_22104);
and U23208 (N_23208,N_22128,N_22067);
or U23209 (N_23209,N_21987,N_21291);
nand U23210 (N_23210,N_21808,N_22129);
or U23211 (N_23211,N_22233,N_22071);
xnor U23212 (N_23212,N_21725,N_21580);
or U23213 (N_23213,N_22221,N_22274);
nand U23214 (N_23214,N_21273,N_22488);
xnor U23215 (N_23215,N_21399,N_22115);
and U23216 (N_23216,N_21690,N_21861);
and U23217 (N_23217,N_21398,N_22008);
xnor U23218 (N_23218,N_21252,N_22162);
and U23219 (N_23219,N_21303,N_21674);
xor U23220 (N_23220,N_22208,N_21841);
or U23221 (N_23221,N_21296,N_21436);
nand U23222 (N_23222,N_21655,N_21375);
nor U23223 (N_23223,N_21745,N_21899);
nor U23224 (N_23224,N_22345,N_21446);
and U23225 (N_23225,N_22091,N_22096);
nand U23226 (N_23226,N_21683,N_22126);
and U23227 (N_23227,N_21777,N_21784);
or U23228 (N_23228,N_22331,N_22060);
nand U23229 (N_23229,N_21686,N_21481);
xnor U23230 (N_23230,N_21913,N_21969);
or U23231 (N_23231,N_22396,N_22439);
or U23232 (N_23232,N_22299,N_22440);
nand U23233 (N_23233,N_21298,N_21421);
and U23234 (N_23234,N_21853,N_22408);
and U23235 (N_23235,N_21718,N_21551);
nand U23236 (N_23236,N_22138,N_22063);
nand U23237 (N_23237,N_21691,N_21815);
xor U23238 (N_23238,N_21425,N_22447);
nand U23239 (N_23239,N_22437,N_22227);
nor U23240 (N_23240,N_21787,N_21466);
xnor U23241 (N_23241,N_21846,N_21962);
nor U23242 (N_23242,N_21328,N_21583);
and U23243 (N_23243,N_21717,N_22150);
nand U23244 (N_23244,N_21450,N_21803);
or U23245 (N_23245,N_22388,N_22184);
nand U23246 (N_23246,N_21575,N_21944);
or U23247 (N_23247,N_21781,N_21274);
or U23248 (N_23248,N_22028,N_21317);
nand U23249 (N_23249,N_21775,N_21722);
nor U23250 (N_23250,N_22460,N_21907);
and U23251 (N_23251,N_21384,N_22476);
or U23252 (N_23252,N_21944,N_21410);
xnor U23253 (N_23253,N_22145,N_21475);
and U23254 (N_23254,N_21866,N_21843);
and U23255 (N_23255,N_21785,N_22192);
or U23256 (N_23256,N_21782,N_21586);
nor U23257 (N_23257,N_22410,N_22314);
xnor U23258 (N_23258,N_21654,N_21768);
or U23259 (N_23259,N_22008,N_22068);
or U23260 (N_23260,N_21855,N_22010);
nand U23261 (N_23261,N_22127,N_21698);
nor U23262 (N_23262,N_21754,N_22201);
or U23263 (N_23263,N_21281,N_21836);
and U23264 (N_23264,N_21877,N_22191);
nor U23265 (N_23265,N_22420,N_21713);
nand U23266 (N_23266,N_22459,N_21568);
nor U23267 (N_23267,N_22495,N_22411);
and U23268 (N_23268,N_22331,N_22376);
nor U23269 (N_23269,N_22317,N_21598);
nand U23270 (N_23270,N_21325,N_22336);
or U23271 (N_23271,N_22155,N_22350);
or U23272 (N_23272,N_21331,N_22447);
nor U23273 (N_23273,N_21424,N_21477);
and U23274 (N_23274,N_22010,N_22239);
xnor U23275 (N_23275,N_21713,N_22306);
nor U23276 (N_23276,N_21455,N_21874);
or U23277 (N_23277,N_22117,N_21354);
xnor U23278 (N_23278,N_21714,N_22073);
and U23279 (N_23279,N_21893,N_21958);
and U23280 (N_23280,N_21715,N_21439);
nor U23281 (N_23281,N_22318,N_21699);
nor U23282 (N_23282,N_21421,N_21620);
or U23283 (N_23283,N_21939,N_21878);
xor U23284 (N_23284,N_21775,N_21917);
and U23285 (N_23285,N_21880,N_22328);
nand U23286 (N_23286,N_21364,N_22358);
nand U23287 (N_23287,N_22440,N_21792);
xor U23288 (N_23288,N_21648,N_22323);
or U23289 (N_23289,N_22355,N_21472);
xor U23290 (N_23290,N_21417,N_21627);
xnor U23291 (N_23291,N_22433,N_21362);
or U23292 (N_23292,N_22427,N_21992);
nor U23293 (N_23293,N_21835,N_21410);
nor U23294 (N_23294,N_22050,N_22364);
xor U23295 (N_23295,N_21623,N_21856);
xor U23296 (N_23296,N_21419,N_22106);
nor U23297 (N_23297,N_22195,N_22356);
and U23298 (N_23298,N_21861,N_22374);
nor U23299 (N_23299,N_22300,N_22029);
and U23300 (N_23300,N_21293,N_21288);
nor U23301 (N_23301,N_21864,N_21627);
or U23302 (N_23302,N_22335,N_22117);
nand U23303 (N_23303,N_22250,N_22350);
and U23304 (N_23304,N_22278,N_22405);
xnor U23305 (N_23305,N_22257,N_22142);
nand U23306 (N_23306,N_22297,N_22258);
nor U23307 (N_23307,N_22464,N_21525);
or U23308 (N_23308,N_22327,N_21337);
or U23309 (N_23309,N_21789,N_22319);
nand U23310 (N_23310,N_22016,N_22087);
and U23311 (N_23311,N_21843,N_21436);
and U23312 (N_23312,N_21557,N_21353);
or U23313 (N_23313,N_21909,N_22486);
or U23314 (N_23314,N_21444,N_22053);
or U23315 (N_23315,N_21724,N_21800);
nor U23316 (N_23316,N_21263,N_21639);
nand U23317 (N_23317,N_21864,N_21263);
or U23318 (N_23318,N_22311,N_21656);
nand U23319 (N_23319,N_21602,N_22354);
xor U23320 (N_23320,N_21545,N_22012);
or U23321 (N_23321,N_21278,N_21313);
or U23322 (N_23322,N_21592,N_21471);
or U23323 (N_23323,N_22303,N_21526);
xor U23324 (N_23324,N_21752,N_22393);
and U23325 (N_23325,N_21656,N_22421);
or U23326 (N_23326,N_21890,N_22472);
and U23327 (N_23327,N_22155,N_21909);
nor U23328 (N_23328,N_22349,N_21317);
xor U23329 (N_23329,N_22353,N_21591);
nand U23330 (N_23330,N_21863,N_21915);
and U23331 (N_23331,N_21468,N_22254);
nor U23332 (N_23332,N_22146,N_21323);
and U23333 (N_23333,N_22246,N_21637);
or U23334 (N_23334,N_21879,N_22374);
and U23335 (N_23335,N_21349,N_22228);
and U23336 (N_23336,N_21622,N_22042);
xor U23337 (N_23337,N_22265,N_21918);
nor U23338 (N_23338,N_22199,N_21316);
and U23339 (N_23339,N_22212,N_21734);
nor U23340 (N_23340,N_21478,N_22378);
and U23341 (N_23341,N_21383,N_22223);
xor U23342 (N_23342,N_21472,N_21609);
nand U23343 (N_23343,N_22121,N_21349);
and U23344 (N_23344,N_22494,N_22014);
or U23345 (N_23345,N_21671,N_22273);
and U23346 (N_23346,N_22017,N_22494);
nand U23347 (N_23347,N_21301,N_22299);
or U23348 (N_23348,N_21876,N_21502);
and U23349 (N_23349,N_21932,N_21930);
and U23350 (N_23350,N_22060,N_22396);
xor U23351 (N_23351,N_21466,N_21634);
nand U23352 (N_23352,N_21489,N_21427);
or U23353 (N_23353,N_21977,N_22459);
xor U23354 (N_23354,N_21455,N_22169);
xnor U23355 (N_23355,N_21620,N_22068);
xnor U23356 (N_23356,N_21684,N_22286);
or U23357 (N_23357,N_21269,N_22114);
xor U23358 (N_23358,N_21855,N_21444);
xor U23359 (N_23359,N_21844,N_22326);
nand U23360 (N_23360,N_21831,N_21463);
or U23361 (N_23361,N_21859,N_22475);
or U23362 (N_23362,N_21883,N_21674);
nor U23363 (N_23363,N_22045,N_22046);
xor U23364 (N_23364,N_22299,N_21534);
or U23365 (N_23365,N_22327,N_22338);
nand U23366 (N_23366,N_21377,N_21422);
and U23367 (N_23367,N_22037,N_21458);
or U23368 (N_23368,N_21418,N_22213);
and U23369 (N_23369,N_21974,N_21996);
nand U23370 (N_23370,N_22426,N_21331);
and U23371 (N_23371,N_22324,N_21819);
and U23372 (N_23372,N_22103,N_21862);
nor U23373 (N_23373,N_22096,N_21588);
or U23374 (N_23374,N_21377,N_21621);
or U23375 (N_23375,N_22208,N_21682);
xnor U23376 (N_23376,N_22351,N_22451);
nor U23377 (N_23377,N_21865,N_21637);
nand U23378 (N_23378,N_21824,N_21306);
or U23379 (N_23379,N_21735,N_22216);
nand U23380 (N_23380,N_22450,N_22401);
or U23381 (N_23381,N_22329,N_21607);
nor U23382 (N_23382,N_22066,N_21725);
or U23383 (N_23383,N_21519,N_21459);
nand U23384 (N_23384,N_22400,N_21973);
and U23385 (N_23385,N_21641,N_21284);
xnor U23386 (N_23386,N_21909,N_21775);
xnor U23387 (N_23387,N_21409,N_21504);
or U23388 (N_23388,N_21769,N_21559);
and U23389 (N_23389,N_22000,N_22410);
and U23390 (N_23390,N_21738,N_21686);
or U23391 (N_23391,N_21606,N_21450);
or U23392 (N_23392,N_22443,N_21383);
nor U23393 (N_23393,N_22037,N_22352);
xnor U23394 (N_23394,N_22354,N_21937);
or U23395 (N_23395,N_22376,N_22274);
nand U23396 (N_23396,N_22227,N_21640);
nor U23397 (N_23397,N_22117,N_22327);
xor U23398 (N_23398,N_21694,N_21516);
nand U23399 (N_23399,N_21859,N_21727);
xor U23400 (N_23400,N_21669,N_21812);
and U23401 (N_23401,N_22161,N_21281);
or U23402 (N_23402,N_22384,N_22163);
xor U23403 (N_23403,N_22062,N_21813);
and U23404 (N_23404,N_22032,N_22266);
nand U23405 (N_23405,N_22074,N_21314);
nor U23406 (N_23406,N_21310,N_21452);
and U23407 (N_23407,N_22044,N_22178);
xor U23408 (N_23408,N_21785,N_21695);
xnor U23409 (N_23409,N_22432,N_22395);
and U23410 (N_23410,N_21895,N_22108);
nor U23411 (N_23411,N_22179,N_22409);
nor U23412 (N_23412,N_21542,N_22009);
and U23413 (N_23413,N_22318,N_21912);
xnor U23414 (N_23414,N_21329,N_21546);
or U23415 (N_23415,N_22062,N_22379);
or U23416 (N_23416,N_22484,N_22160);
nand U23417 (N_23417,N_21953,N_22401);
and U23418 (N_23418,N_21495,N_21787);
xnor U23419 (N_23419,N_21919,N_21469);
nand U23420 (N_23420,N_22113,N_21974);
xor U23421 (N_23421,N_21619,N_21355);
nor U23422 (N_23422,N_21896,N_21739);
nand U23423 (N_23423,N_22077,N_21320);
nand U23424 (N_23424,N_22113,N_22198);
and U23425 (N_23425,N_21289,N_21450);
or U23426 (N_23426,N_22187,N_22093);
nand U23427 (N_23427,N_22480,N_21455);
and U23428 (N_23428,N_22332,N_21685);
and U23429 (N_23429,N_21390,N_21690);
xnor U23430 (N_23430,N_21757,N_21688);
or U23431 (N_23431,N_22002,N_22129);
and U23432 (N_23432,N_22298,N_21869);
and U23433 (N_23433,N_21382,N_21732);
and U23434 (N_23434,N_21859,N_22369);
and U23435 (N_23435,N_22139,N_22428);
xnor U23436 (N_23436,N_21312,N_21650);
and U23437 (N_23437,N_21933,N_21702);
nand U23438 (N_23438,N_21814,N_22173);
and U23439 (N_23439,N_21722,N_21771);
or U23440 (N_23440,N_22321,N_21616);
or U23441 (N_23441,N_22239,N_22068);
and U23442 (N_23442,N_22459,N_21958);
nand U23443 (N_23443,N_21476,N_21380);
nand U23444 (N_23444,N_22029,N_21709);
and U23445 (N_23445,N_21471,N_21988);
and U23446 (N_23446,N_21379,N_22047);
and U23447 (N_23447,N_22356,N_22455);
nand U23448 (N_23448,N_22269,N_21633);
and U23449 (N_23449,N_22028,N_22018);
and U23450 (N_23450,N_21423,N_21451);
xor U23451 (N_23451,N_22467,N_21892);
xor U23452 (N_23452,N_22198,N_22030);
xor U23453 (N_23453,N_22049,N_21496);
xor U23454 (N_23454,N_21968,N_21961);
or U23455 (N_23455,N_21737,N_21352);
or U23456 (N_23456,N_21826,N_21347);
and U23457 (N_23457,N_22078,N_21450);
nand U23458 (N_23458,N_22392,N_21507);
nand U23459 (N_23459,N_22104,N_22464);
nor U23460 (N_23460,N_21289,N_21744);
or U23461 (N_23461,N_21442,N_21854);
and U23462 (N_23462,N_21947,N_22077);
nand U23463 (N_23463,N_21560,N_21841);
nor U23464 (N_23464,N_21884,N_22457);
xor U23465 (N_23465,N_21733,N_21253);
and U23466 (N_23466,N_21321,N_22169);
nand U23467 (N_23467,N_22436,N_21962);
xnor U23468 (N_23468,N_21470,N_21515);
or U23469 (N_23469,N_21646,N_22352);
nor U23470 (N_23470,N_21853,N_22452);
nor U23471 (N_23471,N_22084,N_22058);
xor U23472 (N_23472,N_22178,N_22495);
nor U23473 (N_23473,N_22215,N_22050);
or U23474 (N_23474,N_22201,N_21514);
or U23475 (N_23475,N_21730,N_21628);
nor U23476 (N_23476,N_21648,N_21902);
nor U23477 (N_23477,N_21291,N_21281);
nor U23478 (N_23478,N_21436,N_21575);
nor U23479 (N_23479,N_21643,N_21534);
xnor U23480 (N_23480,N_22332,N_21911);
nor U23481 (N_23481,N_21453,N_22069);
xnor U23482 (N_23482,N_21411,N_21341);
or U23483 (N_23483,N_21843,N_22001);
or U23484 (N_23484,N_22480,N_22289);
and U23485 (N_23485,N_21555,N_21652);
and U23486 (N_23486,N_21541,N_21674);
nor U23487 (N_23487,N_22052,N_21802);
or U23488 (N_23488,N_21618,N_21706);
or U23489 (N_23489,N_21929,N_21522);
and U23490 (N_23490,N_21791,N_21463);
xnor U23491 (N_23491,N_22241,N_21679);
nand U23492 (N_23492,N_21948,N_21671);
xnor U23493 (N_23493,N_21640,N_21687);
xnor U23494 (N_23494,N_22377,N_21561);
or U23495 (N_23495,N_22028,N_22020);
nor U23496 (N_23496,N_22065,N_21602);
nand U23497 (N_23497,N_21570,N_22195);
or U23498 (N_23498,N_21352,N_21320);
nor U23499 (N_23499,N_21631,N_21407);
nor U23500 (N_23500,N_21765,N_22327);
or U23501 (N_23501,N_22015,N_21693);
nor U23502 (N_23502,N_21586,N_21734);
nand U23503 (N_23503,N_21767,N_21313);
nand U23504 (N_23504,N_22475,N_22285);
nor U23505 (N_23505,N_22312,N_22145);
nor U23506 (N_23506,N_22181,N_21735);
or U23507 (N_23507,N_22431,N_22136);
nand U23508 (N_23508,N_21752,N_22352);
or U23509 (N_23509,N_21673,N_22405);
nand U23510 (N_23510,N_22362,N_21880);
nand U23511 (N_23511,N_22077,N_22422);
nor U23512 (N_23512,N_22115,N_21930);
nor U23513 (N_23513,N_21872,N_22340);
and U23514 (N_23514,N_21380,N_22088);
xnor U23515 (N_23515,N_21605,N_22066);
nand U23516 (N_23516,N_22426,N_21675);
nor U23517 (N_23517,N_22325,N_21340);
or U23518 (N_23518,N_21687,N_21897);
or U23519 (N_23519,N_22420,N_21562);
xnor U23520 (N_23520,N_21452,N_21755);
or U23521 (N_23521,N_21318,N_22152);
nor U23522 (N_23522,N_22393,N_21706);
and U23523 (N_23523,N_21944,N_21625);
and U23524 (N_23524,N_22291,N_22457);
xor U23525 (N_23525,N_21667,N_21826);
or U23526 (N_23526,N_21859,N_22146);
and U23527 (N_23527,N_21614,N_21542);
nand U23528 (N_23528,N_21840,N_22357);
nand U23529 (N_23529,N_21915,N_21978);
and U23530 (N_23530,N_21678,N_21784);
and U23531 (N_23531,N_21743,N_21555);
or U23532 (N_23532,N_22313,N_21542);
and U23533 (N_23533,N_21761,N_21373);
xor U23534 (N_23534,N_22216,N_21806);
or U23535 (N_23535,N_21882,N_21357);
xnor U23536 (N_23536,N_22272,N_22250);
xnor U23537 (N_23537,N_21262,N_22271);
and U23538 (N_23538,N_22107,N_21621);
nor U23539 (N_23539,N_22419,N_22237);
xnor U23540 (N_23540,N_22168,N_22068);
nor U23541 (N_23541,N_21746,N_21594);
xor U23542 (N_23542,N_21737,N_21251);
nor U23543 (N_23543,N_21619,N_21878);
xnor U23544 (N_23544,N_21782,N_21645);
nand U23545 (N_23545,N_22224,N_21466);
and U23546 (N_23546,N_21545,N_22109);
and U23547 (N_23547,N_22047,N_21835);
nor U23548 (N_23548,N_22393,N_21438);
nor U23549 (N_23549,N_21516,N_21508);
nand U23550 (N_23550,N_21959,N_21563);
xnor U23551 (N_23551,N_21604,N_21627);
nand U23552 (N_23552,N_22440,N_21844);
or U23553 (N_23553,N_21646,N_21302);
and U23554 (N_23554,N_21517,N_21456);
nor U23555 (N_23555,N_21457,N_22135);
and U23556 (N_23556,N_22259,N_21495);
and U23557 (N_23557,N_21629,N_21918);
nor U23558 (N_23558,N_21865,N_22288);
nor U23559 (N_23559,N_21683,N_22162);
xor U23560 (N_23560,N_22081,N_21884);
or U23561 (N_23561,N_22359,N_22322);
and U23562 (N_23562,N_21526,N_22382);
nor U23563 (N_23563,N_21774,N_22194);
xnor U23564 (N_23564,N_22313,N_21369);
xor U23565 (N_23565,N_22169,N_22455);
nand U23566 (N_23566,N_21536,N_21361);
and U23567 (N_23567,N_21384,N_22348);
nand U23568 (N_23568,N_22065,N_21703);
and U23569 (N_23569,N_21813,N_21414);
nor U23570 (N_23570,N_21835,N_22239);
xor U23571 (N_23571,N_21835,N_22164);
xnor U23572 (N_23572,N_21933,N_21695);
xnor U23573 (N_23573,N_21889,N_21278);
xnor U23574 (N_23574,N_21574,N_22061);
xnor U23575 (N_23575,N_22281,N_21397);
xnor U23576 (N_23576,N_21272,N_21641);
and U23577 (N_23577,N_22491,N_22334);
and U23578 (N_23578,N_21456,N_22258);
nor U23579 (N_23579,N_21801,N_22050);
nor U23580 (N_23580,N_22250,N_21642);
nor U23581 (N_23581,N_22098,N_22336);
nor U23582 (N_23582,N_21711,N_21423);
nor U23583 (N_23583,N_22244,N_21360);
nand U23584 (N_23584,N_22244,N_22194);
nand U23585 (N_23585,N_22029,N_22450);
and U23586 (N_23586,N_21411,N_22277);
xor U23587 (N_23587,N_22271,N_21535);
nor U23588 (N_23588,N_21690,N_21737);
nand U23589 (N_23589,N_21254,N_22056);
nand U23590 (N_23590,N_21483,N_21869);
and U23591 (N_23591,N_21837,N_22471);
nand U23592 (N_23592,N_21259,N_22265);
xnor U23593 (N_23593,N_22442,N_21816);
nand U23594 (N_23594,N_22361,N_22331);
nand U23595 (N_23595,N_22313,N_22323);
nand U23596 (N_23596,N_21673,N_22369);
xor U23597 (N_23597,N_21928,N_22212);
or U23598 (N_23598,N_21923,N_21478);
nor U23599 (N_23599,N_21739,N_21620);
or U23600 (N_23600,N_21452,N_22344);
xnor U23601 (N_23601,N_22078,N_21647);
nor U23602 (N_23602,N_21919,N_21951);
xnor U23603 (N_23603,N_21265,N_22044);
nor U23604 (N_23604,N_21334,N_21895);
and U23605 (N_23605,N_22237,N_21253);
nand U23606 (N_23606,N_21800,N_22352);
or U23607 (N_23607,N_21871,N_22476);
nor U23608 (N_23608,N_21672,N_21745);
xor U23609 (N_23609,N_21436,N_22296);
nand U23610 (N_23610,N_21295,N_22385);
xnor U23611 (N_23611,N_22111,N_21454);
nor U23612 (N_23612,N_21829,N_21686);
xor U23613 (N_23613,N_22466,N_22106);
nor U23614 (N_23614,N_21493,N_21522);
xor U23615 (N_23615,N_21576,N_22237);
nor U23616 (N_23616,N_22102,N_21841);
xnor U23617 (N_23617,N_22457,N_21602);
or U23618 (N_23618,N_22393,N_21434);
and U23619 (N_23619,N_22405,N_22113);
or U23620 (N_23620,N_21557,N_22379);
xor U23621 (N_23621,N_22227,N_21750);
and U23622 (N_23622,N_22337,N_21326);
nand U23623 (N_23623,N_21932,N_21290);
nor U23624 (N_23624,N_21780,N_21549);
xor U23625 (N_23625,N_22144,N_21840);
nor U23626 (N_23626,N_21622,N_21884);
xnor U23627 (N_23627,N_21542,N_21485);
xnor U23628 (N_23628,N_22148,N_21295);
nor U23629 (N_23629,N_21634,N_21885);
or U23630 (N_23630,N_21546,N_21777);
and U23631 (N_23631,N_21790,N_21439);
nor U23632 (N_23632,N_21687,N_21359);
and U23633 (N_23633,N_21284,N_21872);
and U23634 (N_23634,N_22335,N_22173);
and U23635 (N_23635,N_21713,N_21495);
or U23636 (N_23636,N_21627,N_21438);
xnor U23637 (N_23637,N_22324,N_21336);
xor U23638 (N_23638,N_21629,N_21633);
nor U23639 (N_23639,N_21368,N_22391);
nand U23640 (N_23640,N_21824,N_22065);
nor U23641 (N_23641,N_22304,N_22313);
and U23642 (N_23642,N_21590,N_22316);
xnor U23643 (N_23643,N_21764,N_21586);
and U23644 (N_23644,N_21344,N_21876);
xor U23645 (N_23645,N_21528,N_22194);
and U23646 (N_23646,N_22481,N_22010);
nor U23647 (N_23647,N_22015,N_22263);
and U23648 (N_23648,N_21562,N_21549);
xor U23649 (N_23649,N_22313,N_22148);
and U23650 (N_23650,N_21940,N_22126);
nand U23651 (N_23651,N_21426,N_22305);
xnor U23652 (N_23652,N_21495,N_21802);
and U23653 (N_23653,N_21932,N_22322);
and U23654 (N_23654,N_21925,N_21606);
or U23655 (N_23655,N_22136,N_21615);
nand U23656 (N_23656,N_22037,N_22183);
xnor U23657 (N_23657,N_21354,N_21982);
and U23658 (N_23658,N_21687,N_21813);
xor U23659 (N_23659,N_21396,N_21416);
nand U23660 (N_23660,N_21653,N_22274);
nand U23661 (N_23661,N_21551,N_22076);
xor U23662 (N_23662,N_21901,N_21977);
and U23663 (N_23663,N_21846,N_22368);
or U23664 (N_23664,N_21773,N_21557);
nor U23665 (N_23665,N_21449,N_21507);
nor U23666 (N_23666,N_22145,N_22349);
or U23667 (N_23667,N_21912,N_22267);
nor U23668 (N_23668,N_21490,N_21307);
xnor U23669 (N_23669,N_22318,N_21881);
and U23670 (N_23670,N_22107,N_21304);
or U23671 (N_23671,N_22045,N_21339);
xnor U23672 (N_23672,N_22332,N_22360);
nand U23673 (N_23673,N_22242,N_21786);
and U23674 (N_23674,N_22407,N_22202);
nor U23675 (N_23675,N_21563,N_22389);
and U23676 (N_23676,N_21789,N_21588);
nor U23677 (N_23677,N_22257,N_22276);
or U23678 (N_23678,N_21338,N_22209);
or U23679 (N_23679,N_21711,N_21483);
nand U23680 (N_23680,N_21535,N_21842);
xor U23681 (N_23681,N_21373,N_21539);
or U23682 (N_23682,N_21667,N_21557);
or U23683 (N_23683,N_22439,N_21406);
nand U23684 (N_23684,N_22121,N_21846);
nand U23685 (N_23685,N_21820,N_22043);
nor U23686 (N_23686,N_21390,N_21855);
nor U23687 (N_23687,N_21898,N_22234);
nand U23688 (N_23688,N_21293,N_21422);
xor U23689 (N_23689,N_22367,N_21833);
and U23690 (N_23690,N_21696,N_21410);
and U23691 (N_23691,N_21580,N_21484);
nor U23692 (N_23692,N_22029,N_21264);
nor U23693 (N_23693,N_21674,N_21774);
and U23694 (N_23694,N_22091,N_21862);
or U23695 (N_23695,N_21980,N_21410);
nand U23696 (N_23696,N_21658,N_21667);
or U23697 (N_23697,N_21730,N_22311);
and U23698 (N_23698,N_21686,N_21789);
and U23699 (N_23699,N_21839,N_21920);
and U23700 (N_23700,N_22294,N_22412);
or U23701 (N_23701,N_21706,N_22412);
or U23702 (N_23702,N_21366,N_21954);
nand U23703 (N_23703,N_22285,N_22087);
nor U23704 (N_23704,N_22225,N_21757);
and U23705 (N_23705,N_22435,N_21906);
or U23706 (N_23706,N_21330,N_21807);
nand U23707 (N_23707,N_22110,N_21791);
or U23708 (N_23708,N_21955,N_22007);
nand U23709 (N_23709,N_22128,N_21252);
nand U23710 (N_23710,N_22141,N_21403);
nand U23711 (N_23711,N_22193,N_21964);
nor U23712 (N_23712,N_22439,N_22182);
nor U23713 (N_23713,N_21379,N_21278);
nor U23714 (N_23714,N_21435,N_21443);
nand U23715 (N_23715,N_22428,N_22496);
nor U23716 (N_23716,N_22290,N_22247);
or U23717 (N_23717,N_21668,N_22036);
nand U23718 (N_23718,N_22382,N_21355);
or U23719 (N_23719,N_21453,N_21816);
xnor U23720 (N_23720,N_22254,N_22079);
or U23721 (N_23721,N_22049,N_22092);
nor U23722 (N_23722,N_22013,N_21307);
and U23723 (N_23723,N_22129,N_21560);
nor U23724 (N_23724,N_22261,N_22437);
and U23725 (N_23725,N_21953,N_21509);
nor U23726 (N_23726,N_22166,N_21692);
xnor U23727 (N_23727,N_21737,N_22154);
or U23728 (N_23728,N_22215,N_22156);
nand U23729 (N_23729,N_22415,N_21321);
xnor U23730 (N_23730,N_22246,N_22373);
nor U23731 (N_23731,N_22019,N_22230);
or U23732 (N_23732,N_21785,N_21882);
or U23733 (N_23733,N_21749,N_21947);
nand U23734 (N_23734,N_21624,N_22181);
and U23735 (N_23735,N_21616,N_21478);
xor U23736 (N_23736,N_22438,N_21834);
or U23737 (N_23737,N_22344,N_21750);
and U23738 (N_23738,N_21333,N_21282);
nor U23739 (N_23739,N_21590,N_21785);
nand U23740 (N_23740,N_21768,N_22004);
xnor U23741 (N_23741,N_22497,N_22285);
or U23742 (N_23742,N_22499,N_22275);
xor U23743 (N_23743,N_22048,N_22256);
nand U23744 (N_23744,N_21836,N_22152);
nand U23745 (N_23745,N_21782,N_21848);
and U23746 (N_23746,N_21473,N_22118);
nor U23747 (N_23747,N_21782,N_21778);
nor U23748 (N_23748,N_21373,N_21816);
xor U23749 (N_23749,N_21416,N_22350);
nand U23750 (N_23750,N_22841,N_22875);
nand U23751 (N_23751,N_22811,N_23459);
xor U23752 (N_23752,N_22592,N_23419);
nand U23753 (N_23753,N_23441,N_23457);
nor U23754 (N_23754,N_22827,N_22505);
and U23755 (N_23755,N_23378,N_23034);
nor U23756 (N_23756,N_22544,N_23136);
or U23757 (N_23757,N_22671,N_23511);
nand U23758 (N_23758,N_23232,N_22750);
and U23759 (N_23759,N_22680,N_23663);
nor U23760 (N_23760,N_22936,N_23729);
nand U23761 (N_23761,N_22663,N_22596);
and U23762 (N_23762,N_22534,N_22729);
and U23763 (N_23763,N_22763,N_22990);
nand U23764 (N_23764,N_23572,N_23116);
xnor U23765 (N_23765,N_23520,N_23696);
nor U23766 (N_23766,N_22714,N_23235);
nor U23767 (N_23767,N_23125,N_22994);
xnor U23768 (N_23768,N_23166,N_23635);
or U23769 (N_23769,N_23623,N_23415);
nor U23770 (N_23770,N_22880,N_23484);
nand U23771 (N_23771,N_23610,N_22611);
and U23772 (N_23772,N_23108,N_22650);
or U23773 (N_23773,N_22560,N_23720);
or U23774 (N_23774,N_23042,N_23372);
and U23775 (N_23775,N_22806,N_23045);
nand U23776 (N_23776,N_22546,N_23399);
nor U23777 (N_23777,N_23532,N_23576);
nor U23778 (N_23778,N_22745,N_22710);
xnor U23779 (N_23779,N_22629,N_23214);
xor U23780 (N_23780,N_23287,N_22620);
nand U23781 (N_23781,N_22588,N_23543);
and U23782 (N_23782,N_22801,N_22830);
and U23783 (N_23783,N_23551,N_23335);
xor U23784 (N_23784,N_23434,N_22631);
nor U23785 (N_23785,N_22539,N_22789);
and U23786 (N_23786,N_22838,N_23657);
nand U23787 (N_23787,N_22869,N_23546);
and U23788 (N_23788,N_23703,N_23028);
xnor U23789 (N_23789,N_23365,N_23246);
or U23790 (N_23790,N_22832,N_22787);
or U23791 (N_23791,N_22943,N_23070);
nor U23792 (N_23792,N_23278,N_23143);
xnor U23793 (N_23793,N_22567,N_23435);
and U23794 (N_23794,N_23529,N_22939);
nand U23795 (N_23795,N_22898,N_23407);
nor U23796 (N_23796,N_23651,N_22824);
nand U23797 (N_23797,N_23142,N_22595);
nand U23798 (N_23798,N_23380,N_23425);
and U23799 (N_23799,N_22513,N_23749);
nand U23800 (N_23800,N_22713,N_22857);
and U23801 (N_23801,N_22615,N_23538);
nand U23802 (N_23802,N_23063,N_23173);
nor U23803 (N_23803,N_22905,N_22897);
nor U23804 (N_23804,N_22780,N_22711);
and U23805 (N_23805,N_22719,N_23440);
nor U23806 (N_23806,N_23376,N_23452);
and U23807 (N_23807,N_23171,N_23517);
and U23808 (N_23808,N_22549,N_23619);
xnor U23809 (N_23809,N_23496,N_23408);
nand U23810 (N_23810,N_23698,N_23224);
nor U23811 (N_23811,N_23454,N_22540);
nor U23812 (N_23812,N_23715,N_22632);
nand U23813 (N_23813,N_22609,N_23015);
or U23814 (N_23814,N_22538,N_22687);
and U23815 (N_23815,N_22746,N_23343);
xor U23816 (N_23816,N_23398,N_23726);
and U23817 (N_23817,N_23205,N_22533);
xnor U23818 (N_23818,N_22951,N_23662);
and U23819 (N_23819,N_22508,N_23445);
or U23820 (N_23820,N_23183,N_23602);
and U23821 (N_23821,N_23683,N_23067);
xor U23822 (N_23822,N_23233,N_23119);
nor U23823 (N_23823,N_23225,N_23585);
and U23824 (N_23824,N_23601,N_23073);
or U23825 (N_23825,N_23467,N_23327);
nand U23826 (N_23826,N_23148,N_22522);
nand U23827 (N_23827,N_22656,N_23540);
or U23828 (N_23828,N_23331,N_23675);
or U23829 (N_23829,N_23220,N_22678);
xor U23830 (N_23830,N_23075,N_23172);
and U23831 (N_23831,N_22602,N_23025);
or U23832 (N_23832,N_23210,N_23262);
and U23833 (N_23833,N_22863,N_23204);
nand U23834 (N_23834,N_22575,N_22755);
or U23835 (N_23835,N_23126,N_22563);
xnor U23836 (N_23836,N_22800,N_22870);
or U23837 (N_23837,N_23266,N_23253);
nor U23838 (N_23838,N_22784,N_23490);
xor U23839 (N_23839,N_23003,N_23134);
xor U23840 (N_23840,N_23570,N_22695);
or U23841 (N_23841,N_23443,N_23433);
xor U23842 (N_23842,N_23049,N_23040);
nor U23843 (N_23843,N_23492,N_23303);
xnor U23844 (N_23844,N_22941,N_22574);
xor U23845 (N_23845,N_22966,N_23221);
nor U23846 (N_23846,N_22531,N_22665);
nand U23847 (N_23847,N_22682,N_23724);
or U23848 (N_23848,N_22614,N_23087);
nor U23849 (N_23849,N_23285,N_22970);
nor U23850 (N_23850,N_22584,N_23109);
and U23851 (N_23851,N_23313,N_23052);
nor U23852 (N_23852,N_23397,N_23153);
or U23853 (N_23853,N_22786,N_23130);
xnor U23854 (N_23854,N_22555,N_22778);
nand U23855 (N_23855,N_22667,N_22621);
xor U23856 (N_23856,N_23339,N_23530);
and U23857 (N_23857,N_23627,N_22652);
or U23858 (N_23858,N_23731,N_22934);
or U23859 (N_23859,N_22581,N_22747);
nand U23860 (N_23860,N_22954,N_23298);
or U23861 (N_23861,N_22762,N_22967);
or U23862 (N_23862,N_22925,N_22895);
or U23863 (N_23863,N_23323,N_23456);
nor U23864 (N_23864,N_22541,N_22702);
xnor U23865 (N_23865,N_22879,N_23636);
nor U23866 (N_23866,N_23550,N_22878);
nand U23867 (N_23867,N_23249,N_23737);
or U23868 (N_23868,N_23702,N_23088);
nand U23869 (N_23869,N_22674,N_22888);
or U23870 (N_23870,N_23306,N_23678);
or U23871 (N_23871,N_22782,N_23212);
nand U23872 (N_23872,N_22660,N_22706);
xnor U23873 (N_23873,N_23414,N_23213);
and U23874 (N_23874,N_23436,N_23138);
xnor U23875 (N_23875,N_23643,N_23605);
xnor U23876 (N_23876,N_22518,N_23163);
nor U23877 (N_23877,N_23290,N_23730);
xnor U23878 (N_23878,N_23017,N_23613);
and U23879 (N_23879,N_22666,N_22769);
xnor U23880 (N_23880,N_23647,N_23681);
nor U23881 (N_23881,N_22507,N_23571);
xor U23882 (N_23882,N_23207,N_23367);
nand U23883 (N_23883,N_23498,N_23389);
nor U23884 (N_23884,N_22950,N_23732);
nand U23885 (N_23885,N_22669,N_22753);
xor U23886 (N_23886,N_23476,N_23057);
or U23887 (N_23887,N_22552,N_23451);
xnor U23888 (N_23888,N_23641,N_23309);
nor U23889 (N_23889,N_22573,N_23320);
and U23890 (N_23890,N_22593,N_22924);
and U23891 (N_23891,N_23533,N_23453);
and U23892 (N_23892,N_23267,N_22808);
nor U23893 (N_23893,N_23628,N_22709);
xnor U23894 (N_23894,N_22532,N_23649);
nor U23895 (N_23895,N_22772,N_23591);
and U23896 (N_23896,N_22884,N_23107);
and U23897 (N_23897,N_22585,N_22633);
xnor U23898 (N_23898,N_23547,N_22908);
xor U23899 (N_23899,N_22591,N_23429);
xor U23900 (N_23900,N_22501,N_23666);
nand U23901 (N_23901,N_23008,N_22873);
or U23902 (N_23902,N_22969,N_23727);
nand U23903 (N_23903,N_22771,N_23607);
nor U23904 (N_23904,N_23553,N_22960);
nor U23905 (N_23905,N_23507,N_22985);
nor U23906 (N_23906,N_22959,N_23653);
xor U23907 (N_23907,N_23240,N_23076);
and U23908 (N_23908,N_22701,N_23346);
or U23909 (N_23909,N_22984,N_23528);
nand U23910 (N_23910,N_23735,N_23481);
xor U23911 (N_23911,N_23264,N_22752);
and U23912 (N_23912,N_23086,N_23395);
nor U23913 (N_23913,N_22610,N_22881);
nor U23914 (N_23914,N_22860,N_22697);
xor U23915 (N_23915,N_22707,N_23127);
or U23916 (N_23916,N_23223,N_23072);
nor U23917 (N_23917,N_23560,N_22933);
nand U23918 (N_23918,N_22728,N_23349);
or U23919 (N_23919,N_23182,N_23275);
xor U23920 (N_23920,N_22599,N_22818);
xnor U23921 (N_23921,N_22802,N_22642);
and U23922 (N_23922,N_23710,N_23631);
nand U23923 (N_23923,N_22644,N_23286);
and U23924 (N_23924,N_23679,N_22686);
or U23925 (N_23925,N_23305,N_23404);
or U23926 (N_23926,N_23633,N_23449);
and U23927 (N_23927,N_22562,N_23312);
or U23928 (N_23928,N_22963,N_23699);
or U23929 (N_23929,N_23310,N_22910);
xor U23930 (N_23930,N_22866,N_22504);
and U23931 (N_23931,N_22502,N_23314);
nor U23932 (N_23932,N_22834,N_22547);
nor U23933 (N_23933,N_22740,N_23200);
nor U23934 (N_23934,N_23373,N_23186);
nand U23935 (N_23935,N_22766,N_22576);
or U23936 (N_23936,N_23640,N_23377);
or U23937 (N_23937,N_22848,N_23743);
nand U23938 (N_23938,N_22964,N_22862);
nand U23939 (N_23939,N_23512,N_23552);
or U23940 (N_23940,N_23615,N_23439);
nand U23941 (N_23941,N_22657,N_23013);
and U23942 (N_23942,N_22989,N_23472);
or U23943 (N_23943,N_23341,N_22675);
or U23944 (N_23944,N_22828,N_23606);
xor U23945 (N_23945,N_23642,N_23104);
and U23946 (N_23946,N_23078,N_23600);
xnor U23947 (N_23947,N_22927,N_22916);
nor U23948 (N_23948,N_23079,N_22991);
and U23949 (N_23949,N_22942,N_23632);
nand U23950 (N_23950,N_22708,N_23069);
and U23951 (N_23951,N_23096,N_23742);
and U23952 (N_23952,N_23021,N_23676);
nor U23953 (N_23953,N_23508,N_22521);
and U23954 (N_23954,N_23250,N_23243);
nor U23955 (N_23955,N_23318,N_23744);
xor U23956 (N_23956,N_22906,N_23444);
nor U23957 (N_23957,N_22703,N_23721);
xnor U23958 (N_23958,N_22823,N_23705);
nand U23959 (N_23959,N_23603,N_23736);
nor U23960 (N_23960,N_23061,N_22949);
xor U23961 (N_23961,N_23673,N_22980);
nor U23962 (N_23962,N_22922,N_22699);
and U23963 (N_23963,N_22516,N_23248);
or U23964 (N_23964,N_22907,N_22993);
or U23965 (N_23965,N_23252,N_23035);
nand U23966 (N_23966,N_23189,N_23195);
nand U23967 (N_23967,N_23409,N_23217);
xnor U23968 (N_23968,N_23599,N_22545);
or U23969 (N_23969,N_23621,N_23241);
and U23970 (N_23970,N_22972,N_23670);
xnor U23971 (N_23971,N_23717,N_23468);
and U23972 (N_23972,N_22958,N_23251);
nand U23973 (N_23973,N_22770,N_23258);
nand U23974 (N_23974,N_23020,N_23450);
xor U23975 (N_23975,N_23350,N_23272);
nand U23976 (N_23976,N_22572,N_23392);
or U23977 (N_23977,N_23105,N_23165);
nor U23978 (N_23978,N_23351,N_22810);
nor U23979 (N_23979,N_22654,N_23374);
and U23980 (N_23980,N_22978,N_23030);
nor U23981 (N_23981,N_22515,N_23145);
nor U23982 (N_23982,N_23010,N_23301);
xnor U23983 (N_23983,N_22788,N_22730);
or U23984 (N_23984,N_23483,N_23411);
xnor U23985 (N_23985,N_23348,N_22512);
nand U23986 (N_23986,N_22874,N_22809);
nor U23987 (N_23987,N_22684,N_23626);
or U23988 (N_23988,N_22836,N_22727);
xor U23989 (N_23989,N_22510,N_23499);
nand U23990 (N_23990,N_23300,N_23537);
xnor U23991 (N_23991,N_23405,N_22524);
xor U23992 (N_23992,N_22992,N_23677);
xnor U23993 (N_23993,N_22847,N_23523);
and U23994 (N_23994,N_23048,N_22506);
xnor U23995 (N_23995,N_23463,N_23497);
or U23996 (N_23996,N_23384,N_22833);
nand U23997 (N_23997,N_23009,N_23674);
nor U23998 (N_23998,N_23355,N_23427);
xor U23999 (N_23999,N_22672,N_23222);
or U24000 (N_24000,N_23328,N_22913);
or U24001 (N_24001,N_22998,N_23158);
xor U24002 (N_24002,N_23667,N_22726);
and U24003 (N_24003,N_23442,N_22931);
nand U24004 (N_24004,N_23489,N_22759);
or U24005 (N_24005,N_22887,N_23334);
nand U24006 (N_24006,N_22635,N_23315);
nand U24007 (N_24007,N_23304,N_23245);
nor U24008 (N_24008,N_23693,N_23029);
nor U24009 (N_24009,N_23039,N_22914);
nor U24010 (N_24010,N_23132,N_23032);
and U24011 (N_24011,N_23283,N_23518);
and U24012 (N_24012,N_23092,N_22689);
nand U24013 (N_24013,N_22628,N_22817);
and U24014 (N_24014,N_22872,N_22751);
or U24015 (N_24015,N_23470,N_23332);
and U24016 (N_24016,N_23006,N_22804);
or U24017 (N_24017,N_23082,N_22733);
and U24018 (N_24018,N_23123,N_22662);
nand U24019 (N_24019,N_22867,N_23708);
nand U24020 (N_24020,N_23236,N_22673);
nand U24021 (N_24021,N_22921,N_23639);
or U24022 (N_24022,N_23084,N_22854);
nor U24023 (N_24023,N_23360,N_22937);
nand U24024 (N_24024,N_23162,N_22626);
and U24025 (N_24025,N_23541,N_22917);
or U24026 (N_24026,N_23579,N_23595);
nor U24027 (N_24027,N_22586,N_22556);
or U24028 (N_24028,N_23176,N_23050);
nand U24029 (N_24029,N_23027,N_23475);
or U24030 (N_24030,N_23375,N_23358);
nor U24031 (N_24031,N_23549,N_23118);
nor U24032 (N_24032,N_22821,N_22903);
or U24033 (N_24033,N_23161,N_23525);
nand U24034 (N_24034,N_22700,N_23329);
nand U24035 (N_24035,N_22739,N_23352);
xor U24036 (N_24036,N_22928,N_23519);
nand U24037 (N_24037,N_23685,N_23011);
nor U24038 (N_24038,N_22825,N_23159);
nand U24039 (N_24039,N_22600,N_22839);
or U24040 (N_24040,N_23294,N_23692);
xnor U24041 (N_24041,N_23170,N_23277);
nand U24042 (N_24042,N_23326,N_23357);
xnor U24043 (N_24043,N_22736,N_23437);
and U24044 (N_24044,N_23137,N_23056);
or U24045 (N_24045,N_22935,N_23098);
xor U24046 (N_24046,N_23055,N_22957);
nand U24047 (N_24047,N_23568,N_23612);
nand U24048 (N_24048,N_22911,N_23263);
or U24049 (N_24049,N_22630,N_22637);
xnor U24050 (N_24050,N_22734,N_22568);
nand U24051 (N_24051,N_23164,N_22803);
and U24052 (N_24052,N_22999,N_23094);
xnor U24053 (N_24053,N_23645,N_23388);
xnor U24054 (N_24054,N_22845,N_23062);
and U24055 (N_24055,N_23071,N_23700);
xor U24056 (N_24056,N_23191,N_23578);
or U24057 (N_24057,N_23120,N_22775);
or U24058 (N_24058,N_22659,N_22822);
nand U24059 (N_24059,N_22981,N_23493);
nor U24060 (N_24060,N_23690,N_23292);
and U24061 (N_24061,N_22738,N_23167);
nand U24062 (N_24062,N_22798,N_23714);
or U24063 (N_24063,N_22525,N_22519);
and U24064 (N_24064,N_23064,N_23382);
nand U24065 (N_24065,N_22988,N_22855);
or U24066 (N_24066,N_23261,N_22676);
nand U24067 (N_24067,N_23113,N_22975);
and U24068 (N_24068,N_22816,N_23187);
nor U24069 (N_24069,N_22997,N_23354);
nor U24070 (N_24070,N_23366,N_23115);
nand U24071 (N_24071,N_23002,N_22718);
and U24072 (N_24072,N_23394,N_23316);
nor U24073 (N_24073,N_22956,N_23573);
xor U24074 (N_24074,N_23097,N_23622);
nand U24075 (N_24075,N_22773,N_23733);
nor U24076 (N_24076,N_23671,N_23184);
nor U24077 (N_24077,N_23402,N_22899);
nand U24078 (N_24078,N_23648,N_22590);
nand U24079 (N_24079,N_22594,N_23296);
and U24080 (N_24080,N_23426,N_23307);
or U24081 (N_24081,N_23041,N_23000);
nor U24082 (N_24082,N_22996,N_22612);
xor U24083 (N_24083,N_23144,N_23117);
xnor U24084 (N_24084,N_23480,N_22724);
and U24085 (N_24085,N_22831,N_23629);
or U24086 (N_24086,N_22826,N_23654);
nor U24087 (N_24087,N_22514,N_22643);
and U24088 (N_24088,N_23746,N_22776);
and U24089 (N_24089,N_22756,N_23129);
nand U24090 (N_24090,N_22876,N_22731);
nand U24091 (N_24091,N_22843,N_23403);
xor U24092 (N_24092,N_22894,N_23077);
nand U24093 (N_24093,N_23128,N_22646);
or U24094 (N_24094,N_23110,N_22690);
nand U24095 (N_24095,N_23256,N_22570);
nor U24096 (N_24096,N_23141,N_22840);
and U24097 (N_24097,N_22923,N_23385);
nor U24098 (N_24098,N_22692,N_23276);
or U24099 (N_24099,N_23046,N_22946);
nand U24100 (N_24100,N_23637,N_22932);
and U24101 (N_24101,N_22500,N_23151);
nor U24102 (N_24102,N_23099,N_23422);
nor U24103 (N_24103,N_23215,N_22799);
nand U24104 (N_24104,N_23381,N_22623);
nand U24105 (N_24105,N_23695,N_23282);
or U24106 (N_24106,N_23669,N_22744);
nor U24107 (N_24107,N_23417,N_23157);
or U24108 (N_24108,N_22953,N_22685);
nor U24109 (N_24109,N_23455,N_23058);
nand U24110 (N_24110,N_22622,N_23739);
nand U24111 (N_24111,N_22566,N_23515);
nand U24112 (N_24112,N_23524,N_22597);
nor U24113 (N_24113,N_22636,N_23093);
and U24114 (N_24114,N_23004,N_23682);
xor U24115 (N_24115,N_23139,N_23562);
and U24116 (N_24116,N_22886,N_23201);
or U24117 (N_24117,N_23535,N_23299);
and U24118 (N_24118,N_22902,N_22649);
nor U24119 (N_24119,N_22987,N_23644);
and U24120 (N_24120,N_23133,N_23347);
nand U24121 (N_24121,N_23228,N_22580);
or U24122 (N_24122,N_23598,N_23270);
nor U24123 (N_24123,N_23580,N_23706);
nor U24124 (N_24124,N_23206,N_22704);
nor U24125 (N_24125,N_23680,N_22774);
and U24126 (N_24126,N_23593,N_22578);
and U24127 (N_24127,N_23741,N_22829);
xor U24128 (N_24128,N_22767,N_22837);
or U24129 (N_24129,N_22794,N_22948);
xor U24130 (N_24130,N_22758,N_23477);
nand U24131 (N_24131,N_23154,N_22995);
and U24132 (N_24132,N_23396,N_22901);
nor U24133 (N_24133,N_22792,N_22553);
or U24134 (N_24134,N_23242,N_22651);
xnor U24135 (N_24135,N_22864,N_23043);
nand U24136 (N_24136,N_22737,N_23059);
nor U24137 (N_24137,N_23361,N_23464);
and U24138 (N_24138,N_23620,N_23689);
or U24139 (N_24139,N_23630,N_23566);
nor U24140 (N_24140,N_22940,N_23302);
or U24141 (N_24141,N_23646,N_23211);
or U24142 (N_24142,N_23462,N_23234);
nor U24143 (N_24143,N_23694,N_22764);
nor U24144 (N_24144,N_22721,N_23103);
nor U24145 (N_24145,N_23660,N_23418);
xor U24146 (N_24146,N_23718,N_22893);
or U24147 (N_24147,N_22819,N_22781);
xnor U24148 (N_24148,N_23121,N_22768);
nand U24149 (N_24149,N_23012,N_23446);
and U24150 (N_24150,N_23268,N_23036);
or U24151 (N_24151,N_23659,N_22749);
nand U24152 (N_24152,N_23448,N_23582);
nor U24153 (N_24153,N_23711,N_23255);
nor U24154 (N_24154,N_22616,N_23725);
xnor U24155 (N_24155,N_23311,N_23413);
nor U24156 (N_24156,N_23391,N_22688);
xnor U24157 (N_24157,N_23218,N_22741);
xor U24158 (N_24158,N_22529,N_23563);
nor U24159 (N_24159,N_23295,N_23140);
xnor U24160 (N_24160,N_23716,N_23734);
and U24161 (N_24161,N_23555,N_23344);
or U24162 (N_24162,N_22761,N_22909);
xnor U24163 (N_24163,N_22640,N_23474);
nor U24164 (N_24164,N_23155,N_22900);
nand U24165 (N_24165,N_23308,N_23018);
and U24166 (N_24166,N_23065,N_23393);
nor U24167 (N_24167,N_22890,N_22743);
and U24168 (N_24168,N_22589,N_23432);
and U24169 (N_24169,N_23420,N_23370);
xnor U24170 (N_24170,N_23168,N_23428);
nor U24171 (N_24171,N_22868,N_22815);
or U24172 (N_24172,N_22582,N_22624);
nor U24173 (N_24173,N_23514,N_22952);
xor U24174 (N_24174,N_23565,N_23527);
nor U24175 (N_24175,N_23597,N_22796);
nor U24176 (N_24176,N_22835,N_23424);
and U24177 (N_24177,N_22677,N_23400);
or U24178 (N_24178,N_23704,N_23430);
xnor U24179 (N_24179,N_22944,N_22564);
xnor U24180 (N_24180,N_23485,N_22859);
xnor U24181 (N_24181,N_23333,N_22526);
and U24182 (N_24182,N_22965,N_22604);
nand U24183 (N_24183,N_23135,N_22955);
or U24184 (N_24184,N_23356,N_23661);
xor U24185 (N_24185,N_22785,N_22891);
and U24186 (N_24186,N_23713,N_23177);
xnor U24187 (N_24187,N_23719,N_23471);
nand U24188 (N_24188,N_23487,N_23581);
nand U24189 (N_24189,N_23247,N_23491);
nor U24190 (N_24190,N_23421,N_22974);
nand U24191 (N_24191,N_22765,N_22717);
nor U24192 (N_24192,N_23353,N_22691);
xor U24193 (N_24193,N_23583,N_23510);
or U24194 (N_24194,N_23274,N_22904);
and U24195 (N_24195,N_22561,N_22805);
and U24196 (N_24196,N_22783,N_23687);
nand U24197 (N_24197,N_23509,N_22723);
and U24198 (N_24198,N_23656,N_23410);
or U24199 (N_24199,N_23198,N_23122);
nand U24200 (N_24200,N_22748,N_22754);
xor U24201 (N_24201,N_23588,N_22814);
nand U24202 (N_24202,N_22977,N_22947);
or U24203 (N_24203,N_23482,N_23548);
and U24204 (N_24204,N_22537,N_23178);
xnor U24205 (N_24205,N_23539,N_22606);
nor U24206 (N_24206,N_23095,N_23513);
xor U24207 (N_24207,N_22971,N_23216);
nor U24208 (N_24208,N_22962,N_22760);
xnor U24209 (N_24209,N_22797,N_22926);
and U24210 (N_24210,N_23209,N_23617);
and U24211 (N_24211,N_23616,N_22858);
or U24212 (N_24212,N_22511,N_23458);
nand U24213 (N_24213,N_22655,N_23574);
or U24214 (N_24214,N_23265,N_23239);
and U24215 (N_24215,N_23208,N_22715);
nor U24216 (N_24216,N_23586,N_23567);
or U24217 (N_24217,N_23723,N_23544);
or U24218 (N_24218,N_23460,N_22607);
or U24219 (N_24219,N_22634,N_23363);
nand U24220 (N_24220,N_23230,N_23074);
nor U24221 (N_24221,N_22844,N_22536);
nand U24222 (N_24222,N_22535,N_23494);
nand U24223 (N_24223,N_22871,N_23297);
nand U24224 (N_24224,N_22938,N_23709);
or U24225 (N_24225,N_23534,N_23317);
or U24226 (N_24226,N_23081,N_23701);
or U24227 (N_24227,N_22961,N_23169);
nor U24228 (N_24228,N_23387,N_23390);
nor U24229 (N_24229,N_22613,N_23738);
nand U24230 (N_24230,N_22681,N_23345);
xnor U24231 (N_24231,N_23279,N_22527);
or U24232 (N_24232,N_22577,N_23495);
nor U24233 (N_24233,N_22982,N_22850);
nor U24234 (N_24234,N_23054,N_22852);
and U24235 (N_24235,N_23665,N_23066);
nor U24236 (N_24236,N_23728,N_23625);
nand U24237 (N_24237,N_23146,N_22919);
or U24238 (N_24238,N_23545,N_23342);
xor U24239 (N_24239,N_22885,N_23199);
and U24240 (N_24240,N_22777,N_23577);
and U24241 (N_24241,N_23338,N_22598);
xnor U24242 (N_24242,N_23614,N_23007);
xnor U24243 (N_24243,N_23180,N_23505);
xnor U24244 (N_24244,N_23371,N_22779);
nor U24245 (N_24245,N_22571,N_23044);
or U24246 (N_24246,N_23336,N_23016);
nand U24247 (N_24247,N_23416,N_22587);
or U24248 (N_24248,N_23037,N_22661);
nand U24249 (N_24249,N_23479,N_22503);
xor U24250 (N_24250,N_23634,N_23269);
and U24251 (N_24251,N_23090,N_23522);
nor U24252 (N_24252,N_22583,N_23196);
nor U24253 (N_24253,N_22523,N_23500);
and U24254 (N_24254,N_23112,N_23280);
nand U24255 (N_24255,N_22856,N_23594);
and U24256 (N_24256,N_22968,N_23100);
nor U24257 (N_24257,N_22653,N_23503);
nor U24258 (N_24258,N_23672,N_23324);
xor U24259 (N_24259,N_23083,N_23589);
nor U24260 (N_24260,N_23284,N_23194);
nor U24261 (N_24261,N_23556,N_23273);
nor U24262 (N_24262,N_23053,N_22664);
nand U24263 (N_24263,N_23260,N_23051);
nor U24264 (N_24264,N_22853,N_23229);
nor U24265 (N_24265,N_22557,N_23111);
xor U24266 (N_24266,N_23526,N_23575);
and U24267 (N_24267,N_22812,N_23748);
and U24268 (N_24268,N_23592,N_23147);
and U24269 (N_24269,N_23038,N_23536);
or U24270 (N_24270,N_22735,N_22559);
nand U24271 (N_24271,N_23684,N_22716);
xnor U24272 (N_24272,N_22882,N_23596);
xor U24273 (N_24273,N_23340,N_23219);
or U24274 (N_24274,N_22929,N_23152);
and U24275 (N_24275,N_22793,N_23190);
and U24276 (N_24276,N_23559,N_23506);
nand U24277 (N_24277,N_22645,N_23237);
xor U24278 (N_24278,N_22722,N_23712);
and U24279 (N_24279,N_23026,N_22791);
nor U24280 (N_24280,N_23608,N_23558);
nor U24281 (N_24281,N_22725,N_23447);
nor U24282 (N_24282,N_22569,N_23359);
and U24283 (N_24283,N_23697,N_23181);
nand U24284 (N_24284,N_22912,N_23293);
and U24285 (N_24285,N_23174,N_22542);
xor U24286 (N_24286,N_22605,N_23022);
or U24287 (N_24287,N_23244,N_23412);
xnor U24288 (N_24288,N_23587,N_23150);
nand U24289 (N_24289,N_22861,N_23542);
or U24290 (N_24290,N_22720,N_22896);
and U24291 (N_24291,N_22693,N_23722);
and U24292 (N_24292,N_23379,N_23257);
nor U24293 (N_24293,N_23114,N_23466);
xnor U24294 (N_24294,N_22889,N_23488);
nor U24295 (N_24295,N_23238,N_23254);
and U24296 (N_24296,N_23707,N_23655);
xor U24297 (N_24297,N_22530,N_22920);
nand U24298 (N_24298,N_22976,N_22842);
or U24299 (N_24299,N_23478,N_23185);
nor U24300 (N_24300,N_23033,N_23197);
xor U24301 (N_24301,N_22548,N_23438);
nor U24302 (N_24302,N_22668,N_23618);
and U24303 (N_24303,N_23383,N_23465);
nand U24304 (N_24304,N_22618,N_22930);
nand U24305 (N_24305,N_22790,N_23291);
nand U24306 (N_24306,N_23686,N_23330);
and U24307 (N_24307,N_23271,N_22979);
or U24308 (N_24308,N_22603,N_22647);
nand U24309 (N_24309,N_22619,N_23624);
and U24310 (N_24310,N_22846,N_23203);
and U24311 (N_24311,N_23486,N_22757);
nand U24312 (N_24312,N_22617,N_23024);
and U24313 (N_24313,N_22742,N_23089);
or U24314 (N_24314,N_22986,N_23564);
nand U24315 (N_24315,N_23001,N_23369);
xnor U24316 (N_24316,N_23386,N_22509);
nand U24317 (N_24317,N_23611,N_23469);
xor U24318 (N_24318,N_23584,N_22945);
or U24319 (N_24319,N_23068,N_22973);
nand U24320 (N_24320,N_23557,N_22892);
xor U24321 (N_24321,N_23288,N_23202);
or U24322 (N_24322,N_22732,N_23688);
nor U24323 (N_24323,N_22639,N_22918);
or U24324 (N_24324,N_22520,N_23019);
xor U24325 (N_24325,N_22608,N_22877);
nand U24326 (N_24326,N_23160,N_23226);
xnor U24327 (N_24327,N_22641,N_22670);
nand U24328 (N_24328,N_22983,N_22543);
xor U24329 (N_24329,N_22558,N_23259);
xnor U24330 (N_24330,N_22683,N_23060);
nand U24331 (N_24331,N_23691,N_22601);
nand U24332 (N_24332,N_23747,N_23231);
nand U24333 (N_24333,N_23325,N_23740);
nor U24334 (N_24334,N_23504,N_23102);
or U24335 (N_24335,N_23604,N_23080);
nand U24336 (N_24336,N_23175,N_23501);
nor U24337 (N_24337,N_23101,N_23192);
and U24338 (N_24338,N_22849,N_23227);
nor U24339 (N_24339,N_23569,N_23091);
nor U24340 (N_24340,N_23023,N_23554);
nor U24341 (N_24341,N_23609,N_22627);
nand U24342 (N_24342,N_22528,N_23156);
xor U24343 (N_24343,N_23638,N_22820);
or U24344 (N_24344,N_22865,N_22658);
xnor U24345 (N_24345,N_23473,N_22851);
nor U24346 (N_24346,N_23668,N_23031);
or U24347 (N_24347,N_23321,N_22517);
xor U24348 (N_24348,N_23319,N_23431);
nand U24349 (N_24349,N_23362,N_23106);
or U24350 (N_24350,N_23461,N_22883);
and U24351 (N_24351,N_23516,N_23561);
and U24352 (N_24352,N_23149,N_22807);
nor U24353 (N_24353,N_23193,N_22694);
or U24354 (N_24354,N_23521,N_22579);
nor U24355 (N_24355,N_23368,N_23364);
or U24356 (N_24356,N_22813,N_23047);
xnor U24357 (N_24357,N_22625,N_22638);
or U24358 (N_24358,N_23179,N_22565);
xnor U24359 (N_24359,N_22696,N_22712);
and U24360 (N_24360,N_23590,N_22550);
and U24361 (N_24361,N_23531,N_23745);
nor U24362 (N_24362,N_23337,N_22915);
xnor U24363 (N_24363,N_23014,N_22679);
nand U24364 (N_24364,N_22648,N_23085);
and U24365 (N_24365,N_22795,N_23401);
or U24366 (N_24366,N_23658,N_22705);
xnor U24367 (N_24367,N_23005,N_23423);
nor U24368 (N_24368,N_23124,N_23322);
nor U24369 (N_24369,N_23502,N_23281);
xnor U24370 (N_24370,N_23188,N_22554);
nor U24371 (N_24371,N_23131,N_23650);
and U24372 (N_24372,N_23664,N_23406);
nor U24373 (N_24373,N_23289,N_22698);
nand U24374 (N_24374,N_22551,N_23652);
or U24375 (N_24375,N_22831,N_22646);
nand U24376 (N_24376,N_23454,N_22915);
and U24377 (N_24377,N_22843,N_23481);
nor U24378 (N_24378,N_23421,N_23187);
and U24379 (N_24379,N_23556,N_23345);
and U24380 (N_24380,N_23156,N_23454);
xor U24381 (N_24381,N_22924,N_22835);
nor U24382 (N_24382,N_22886,N_23587);
or U24383 (N_24383,N_23364,N_23203);
or U24384 (N_24384,N_23686,N_23675);
xor U24385 (N_24385,N_22503,N_22869);
xnor U24386 (N_24386,N_22541,N_23190);
nor U24387 (N_24387,N_23188,N_23492);
nor U24388 (N_24388,N_23140,N_23437);
or U24389 (N_24389,N_23727,N_23472);
and U24390 (N_24390,N_22630,N_22807);
xnor U24391 (N_24391,N_23293,N_23360);
nor U24392 (N_24392,N_22921,N_22683);
or U24393 (N_24393,N_23549,N_22820);
nor U24394 (N_24394,N_22503,N_23561);
xor U24395 (N_24395,N_23614,N_23553);
xor U24396 (N_24396,N_23592,N_23713);
nand U24397 (N_24397,N_23128,N_23553);
nor U24398 (N_24398,N_23135,N_23372);
and U24399 (N_24399,N_22755,N_23203);
xor U24400 (N_24400,N_23142,N_22714);
nand U24401 (N_24401,N_23227,N_22857);
and U24402 (N_24402,N_22526,N_23007);
xnor U24403 (N_24403,N_22827,N_23666);
or U24404 (N_24404,N_23712,N_22912);
or U24405 (N_24405,N_23306,N_23298);
nand U24406 (N_24406,N_22756,N_22898);
or U24407 (N_24407,N_22693,N_22781);
nand U24408 (N_24408,N_23153,N_22689);
xor U24409 (N_24409,N_23395,N_23678);
nand U24410 (N_24410,N_23081,N_22855);
nor U24411 (N_24411,N_23301,N_23699);
nand U24412 (N_24412,N_23562,N_23323);
nand U24413 (N_24413,N_22962,N_23627);
nand U24414 (N_24414,N_23082,N_22561);
and U24415 (N_24415,N_22928,N_23410);
and U24416 (N_24416,N_22619,N_22759);
and U24417 (N_24417,N_23355,N_23613);
nand U24418 (N_24418,N_23365,N_23512);
nor U24419 (N_24419,N_22578,N_23396);
or U24420 (N_24420,N_23144,N_23522);
or U24421 (N_24421,N_23012,N_23258);
and U24422 (N_24422,N_23571,N_23434);
nand U24423 (N_24423,N_22982,N_23049);
xor U24424 (N_24424,N_23401,N_23011);
nand U24425 (N_24425,N_23709,N_23026);
xor U24426 (N_24426,N_22894,N_23340);
and U24427 (N_24427,N_22747,N_23507);
xor U24428 (N_24428,N_23481,N_22714);
nor U24429 (N_24429,N_22761,N_23304);
xor U24430 (N_24430,N_22611,N_22554);
nand U24431 (N_24431,N_22584,N_22845);
or U24432 (N_24432,N_23103,N_23267);
xor U24433 (N_24433,N_23676,N_23087);
nand U24434 (N_24434,N_22961,N_22760);
nand U24435 (N_24435,N_22645,N_23197);
xor U24436 (N_24436,N_22987,N_23518);
or U24437 (N_24437,N_23667,N_23392);
and U24438 (N_24438,N_23068,N_23100);
and U24439 (N_24439,N_22762,N_23037);
or U24440 (N_24440,N_23679,N_22564);
or U24441 (N_24441,N_22834,N_23033);
and U24442 (N_24442,N_23130,N_22517);
nand U24443 (N_24443,N_23346,N_23625);
nor U24444 (N_24444,N_23692,N_22994);
nand U24445 (N_24445,N_22704,N_23301);
xor U24446 (N_24446,N_23510,N_23143);
and U24447 (N_24447,N_23521,N_23441);
xor U24448 (N_24448,N_23559,N_22939);
or U24449 (N_24449,N_22996,N_23620);
and U24450 (N_24450,N_22900,N_23443);
nor U24451 (N_24451,N_23737,N_23337);
nor U24452 (N_24452,N_23006,N_22560);
and U24453 (N_24453,N_22947,N_22554);
nand U24454 (N_24454,N_23152,N_23621);
nor U24455 (N_24455,N_23556,N_22727);
nand U24456 (N_24456,N_22506,N_22808);
nor U24457 (N_24457,N_23561,N_23052);
nor U24458 (N_24458,N_22610,N_23007);
nor U24459 (N_24459,N_23606,N_23114);
nor U24460 (N_24460,N_23735,N_23360);
nand U24461 (N_24461,N_23380,N_22793);
xnor U24462 (N_24462,N_23606,N_23318);
and U24463 (N_24463,N_22513,N_23517);
nand U24464 (N_24464,N_23334,N_23547);
and U24465 (N_24465,N_23470,N_22978);
or U24466 (N_24466,N_23442,N_22928);
nor U24467 (N_24467,N_23652,N_23603);
nor U24468 (N_24468,N_23613,N_22601);
nand U24469 (N_24469,N_23449,N_23265);
xnor U24470 (N_24470,N_22917,N_23439);
or U24471 (N_24471,N_23190,N_23742);
and U24472 (N_24472,N_23093,N_23583);
or U24473 (N_24473,N_23643,N_23360);
nand U24474 (N_24474,N_22796,N_22595);
nand U24475 (N_24475,N_23332,N_23651);
and U24476 (N_24476,N_22980,N_23294);
nand U24477 (N_24477,N_22636,N_22896);
nand U24478 (N_24478,N_22641,N_23288);
or U24479 (N_24479,N_22957,N_23572);
nand U24480 (N_24480,N_22972,N_23435);
and U24481 (N_24481,N_22697,N_23610);
nor U24482 (N_24482,N_23123,N_22661);
and U24483 (N_24483,N_23268,N_22683);
xnor U24484 (N_24484,N_22963,N_23682);
nor U24485 (N_24485,N_23182,N_23123);
nor U24486 (N_24486,N_23399,N_23537);
and U24487 (N_24487,N_23269,N_23298);
and U24488 (N_24488,N_22682,N_22735);
and U24489 (N_24489,N_23689,N_22614);
xor U24490 (N_24490,N_22712,N_23608);
xor U24491 (N_24491,N_22860,N_22636);
xnor U24492 (N_24492,N_22608,N_22545);
xnor U24493 (N_24493,N_23479,N_22553);
nor U24494 (N_24494,N_23073,N_23050);
nand U24495 (N_24495,N_23107,N_22842);
nor U24496 (N_24496,N_22904,N_23567);
nor U24497 (N_24497,N_23160,N_22972);
xnor U24498 (N_24498,N_22960,N_23699);
nor U24499 (N_24499,N_23479,N_22671);
nand U24500 (N_24500,N_22802,N_23069);
nor U24501 (N_24501,N_22900,N_23337);
xor U24502 (N_24502,N_22609,N_23652);
nand U24503 (N_24503,N_23263,N_23471);
nor U24504 (N_24504,N_22895,N_23108);
or U24505 (N_24505,N_23597,N_23254);
nor U24506 (N_24506,N_23274,N_22827);
nand U24507 (N_24507,N_22924,N_23568);
nor U24508 (N_24508,N_23263,N_23747);
xnor U24509 (N_24509,N_23436,N_23555);
and U24510 (N_24510,N_22811,N_23272);
xor U24511 (N_24511,N_22528,N_23512);
xnor U24512 (N_24512,N_22864,N_23381);
and U24513 (N_24513,N_23402,N_23514);
and U24514 (N_24514,N_23740,N_23608);
nand U24515 (N_24515,N_22825,N_23515);
nand U24516 (N_24516,N_22838,N_23186);
xnor U24517 (N_24517,N_23556,N_23424);
or U24518 (N_24518,N_23220,N_23072);
or U24519 (N_24519,N_22831,N_22535);
and U24520 (N_24520,N_22591,N_23637);
or U24521 (N_24521,N_23077,N_23516);
xor U24522 (N_24522,N_23339,N_22813);
or U24523 (N_24523,N_23423,N_23599);
xnor U24524 (N_24524,N_23644,N_22716);
xor U24525 (N_24525,N_23117,N_23329);
or U24526 (N_24526,N_23006,N_23036);
nand U24527 (N_24527,N_22741,N_23658);
and U24528 (N_24528,N_23555,N_23247);
and U24529 (N_24529,N_23246,N_23596);
or U24530 (N_24530,N_23052,N_22862);
nor U24531 (N_24531,N_23606,N_22540);
nand U24532 (N_24532,N_23117,N_22953);
xnor U24533 (N_24533,N_22570,N_22957);
nand U24534 (N_24534,N_23015,N_23641);
and U24535 (N_24535,N_23184,N_23230);
or U24536 (N_24536,N_22566,N_22559);
nand U24537 (N_24537,N_23518,N_23284);
nand U24538 (N_24538,N_22553,N_22514);
or U24539 (N_24539,N_22536,N_23538);
nand U24540 (N_24540,N_23402,N_23433);
nor U24541 (N_24541,N_22695,N_22860);
xor U24542 (N_24542,N_23467,N_23182);
nand U24543 (N_24543,N_22644,N_23411);
nor U24544 (N_24544,N_22725,N_22552);
and U24545 (N_24545,N_23675,N_22796);
nor U24546 (N_24546,N_22888,N_23002);
xor U24547 (N_24547,N_23263,N_23317);
nor U24548 (N_24548,N_23383,N_22603);
or U24549 (N_24549,N_22962,N_23045);
nand U24550 (N_24550,N_22855,N_22863);
nand U24551 (N_24551,N_22944,N_23746);
nand U24552 (N_24552,N_23684,N_23407);
nor U24553 (N_24553,N_23219,N_23739);
xnor U24554 (N_24554,N_23437,N_22563);
or U24555 (N_24555,N_22972,N_23521);
nand U24556 (N_24556,N_23728,N_23321);
nand U24557 (N_24557,N_23477,N_23618);
xor U24558 (N_24558,N_22878,N_23081);
nor U24559 (N_24559,N_23690,N_23159);
xor U24560 (N_24560,N_22814,N_22748);
and U24561 (N_24561,N_23045,N_23048);
and U24562 (N_24562,N_22733,N_23496);
or U24563 (N_24563,N_23345,N_22519);
nand U24564 (N_24564,N_23321,N_22515);
nor U24565 (N_24565,N_23204,N_23407);
and U24566 (N_24566,N_22856,N_22729);
nand U24567 (N_24567,N_22683,N_23412);
xor U24568 (N_24568,N_22931,N_23372);
nor U24569 (N_24569,N_22595,N_23612);
nand U24570 (N_24570,N_23278,N_22852);
nor U24571 (N_24571,N_22705,N_22532);
xor U24572 (N_24572,N_23506,N_23194);
nand U24573 (N_24573,N_23671,N_22568);
and U24574 (N_24574,N_23687,N_23354);
nor U24575 (N_24575,N_22824,N_23616);
or U24576 (N_24576,N_22920,N_23174);
xnor U24577 (N_24577,N_23087,N_23520);
nand U24578 (N_24578,N_22746,N_23683);
nor U24579 (N_24579,N_23206,N_23009);
nand U24580 (N_24580,N_23044,N_23736);
or U24581 (N_24581,N_23373,N_22918);
nand U24582 (N_24582,N_23271,N_23250);
nand U24583 (N_24583,N_23504,N_22768);
or U24584 (N_24584,N_22660,N_23035);
nand U24585 (N_24585,N_23284,N_22807);
and U24586 (N_24586,N_23072,N_22839);
nor U24587 (N_24587,N_23724,N_22603);
nor U24588 (N_24588,N_23551,N_23373);
xnor U24589 (N_24589,N_23051,N_22664);
nor U24590 (N_24590,N_22949,N_22883);
xor U24591 (N_24591,N_23447,N_23057);
and U24592 (N_24592,N_22794,N_23721);
and U24593 (N_24593,N_23510,N_23431);
xnor U24594 (N_24594,N_22987,N_23256);
nand U24595 (N_24595,N_23007,N_22584);
nor U24596 (N_24596,N_23523,N_23420);
or U24597 (N_24597,N_23361,N_22810);
or U24598 (N_24598,N_23360,N_23748);
nor U24599 (N_24599,N_22825,N_22830);
and U24600 (N_24600,N_22665,N_23050);
or U24601 (N_24601,N_23535,N_23048);
nand U24602 (N_24602,N_23287,N_23279);
or U24603 (N_24603,N_23170,N_22543);
xnor U24604 (N_24604,N_23566,N_23062);
nand U24605 (N_24605,N_22833,N_22777);
and U24606 (N_24606,N_23734,N_22812);
nand U24607 (N_24607,N_23713,N_23022);
nor U24608 (N_24608,N_23183,N_22741);
nor U24609 (N_24609,N_23509,N_22602);
xor U24610 (N_24610,N_22953,N_22579);
nor U24611 (N_24611,N_23010,N_23236);
xnor U24612 (N_24612,N_23644,N_22842);
xor U24613 (N_24613,N_22922,N_22547);
and U24614 (N_24614,N_22555,N_23234);
nor U24615 (N_24615,N_22740,N_22677);
nand U24616 (N_24616,N_23217,N_22569);
and U24617 (N_24617,N_23621,N_22703);
xnor U24618 (N_24618,N_22609,N_22659);
nand U24619 (N_24619,N_23559,N_22755);
or U24620 (N_24620,N_23305,N_22702);
nor U24621 (N_24621,N_23620,N_22547);
xor U24622 (N_24622,N_23021,N_23370);
or U24623 (N_24623,N_23488,N_23237);
or U24624 (N_24624,N_23491,N_23225);
xor U24625 (N_24625,N_22881,N_22647);
or U24626 (N_24626,N_22787,N_23321);
nand U24627 (N_24627,N_23595,N_22683);
and U24628 (N_24628,N_23448,N_22517);
nor U24629 (N_24629,N_22929,N_22606);
xnor U24630 (N_24630,N_23065,N_22511);
xnor U24631 (N_24631,N_23367,N_23275);
and U24632 (N_24632,N_23204,N_23168);
or U24633 (N_24633,N_23073,N_23076);
nor U24634 (N_24634,N_23248,N_23714);
and U24635 (N_24635,N_22569,N_22561);
nor U24636 (N_24636,N_22859,N_23104);
nor U24637 (N_24637,N_23383,N_23501);
or U24638 (N_24638,N_22934,N_23287);
nand U24639 (N_24639,N_22572,N_22801);
nor U24640 (N_24640,N_22575,N_22708);
and U24641 (N_24641,N_23217,N_23456);
nor U24642 (N_24642,N_22777,N_23018);
or U24643 (N_24643,N_23556,N_22728);
and U24644 (N_24644,N_22730,N_22535);
nand U24645 (N_24645,N_22765,N_23389);
nand U24646 (N_24646,N_23647,N_23152);
or U24647 (N_24647,N_22537,N_22896);
nor U24648 (N_24648,N_23304,N_23587);
nor U24649 (N_24649,N_22681,N_22882);
and U24650 (N_24650,N_23637,N_22823);
and U24651 (N_24651,N_23645,N_22802);
and U24652 (N_24652,N_23277,N_22748);
and U24653 (N_24653,N_23481,N_23036);
nor U24654 (N_24654,N_23290,N_23334);
nor U24655 (N_24655,N_22865,N_22945);
xnor U24656 (N_24656,N_23716,N_23102);
and U24657 (N_24657,N_22712,N_23639);
nor U24658 (N_24658,N_22567,N_22673);
nor U24659 (N_24659,N_22701,N_22785);
xor U24660 (N_24660,N_23162,N_23672);
xor U24661 (N_24661,N_23061,N_22886);
xnor U24662 (N_24662,N_22677,N_23465);
or U24663 (N_24663,N_22756,N_22579);
or U24664 (N_24664,N_23481,N_23352);
and U24665 (N_24665,N_23484,N_23170);
and U24666 (N_24666,N_22557,N_23007);
nor U24667 (N_24667,N_23031,N_22625);
xnor U24668 (N_24668,N_23384,N_23577);
xor U24669 (N_24669,N_23158,N_22892);
or U24670 (N_24670,N_23425,N_22635);
xnor U24671 (N_24671,N_23553,N_23414);
or U24672 (N_24672,N_23150,N_23575);
nor U24673 (N_24673,N_23676,N_23234);
and U24674 (N_24674,N_22751,N_23507);
nor U24675 (N_24675,N_23538,N_22921);
xor U24676 (N_24676,N_23383,N_23419);
nand U24677 (N_24677,N_22681,N_23606);
nor U24678 (N_24678,N_23404,N_23335);
and U24679 (N_24679,N_23586,N_23476);
or U24680 (N_24680,N_22562,N_23364);
nand U24681 (N_24681,N_22675,N_22560);
nor U24682 (N_24682,N_23646,N_22514);
nand U24683 (N_24683,N_22750,N_22808);
and U24684 (N_24684,N_22873,N_22912);
xnor U24685 (N_24685,N_22744,N_22560);
or U24686 (N_24686,N_23161,N_23160);
xnor U24687 (N_24687,N_22992,N_23694);
xnor U24688 (N_24688,N_23328,N_23127);
or U24689 (N_24689,N_23507,N_23669);
and U24690 (N_24690,N_22799,N_23399);
xor U24691 (N_24691,N_23102,N_22810);
xor U24692 (N_24692,N_22948,N_22539);
nor U24693 (N_24693,N_23322,N_23508);
nor U24694 (N_24694,N_23359,N_23044);
nor U24695 (N_24695,N_23638,N_23040);
and U24696 (N_24696,N_23288,N_23532);
nor U24697 (N_24697,N_22891,N_23678);
or U24698 (N_24698,N_23266,N_22999);
xnor U24699 (N_24699,N_23390,N_23607);
or U24700 (N_24700,N_23043,N_23392);
nand U24701 (N_24701,N_22881,N_23516);
nor U24702 (N_24702,N_22875,N_23357);
and U24703 (N_24703,N_23144,N_23445);
nor U24704 (N_24704,N_22542,N_23419);
or U24705 (N_24705,N_23268,N_23378);
nand U24706 (N_24706,N_23051,N_22873);
nand U24707 (N_24707,N_22901,N_22927);
nor U24708 (N_24708,N_23375,N_22926);
and U24709 (N_24709,N_22578,N_22805);
nor U24710 (N_24710,N_23049,N_23526);
xnor U24711 (N_24711,N_23409,N_23634);
xnor U24712 (N_24712,N_23204,N_23249);
nand U24713 (N_24713,N_23470,N_22833);
or U24714 (N_24714,N_22763,N_22748);
and U24715 (N_24715,N_23428,N_23660);
and U24716 (N_24716,N_23369,N_23476);
xnor U24717 (N_24717,N_22655,N_23149);
nor U24718 (N_24718,N_23050,N_22722);
nand U24719 (N_24719,N_22523,N_22611);
and U24720 (N_24720,N_23039,N_23359);
and U24721 (N_24721,N_23345,N_22546);
and U24722 (N_24722,N_22562,N_22622);
nand U24723 (N_24723,N_23399,N_22840);
nor U24724 (N_24724,N_23111,N_23550);
xnor U24725 (N_24725,N_23747,N_22643);
and U24726 (N_24726,N_22701,N_23696);
and U24727 (N_24727,N_22713,N_22663);
xor U24728 (N_24728,N_22575,N_22519);
nand U24729 (N_24729,N_23424,N_23561);
and U24730 (N_24730,N_23557,N_22640);
or U24731 (N_24731,N_23188,N_22639);
nor U24732 (N_24732,N_23335,N_23531);
nand U24733 (N_24733,N_23369,N_23258);
xnor U24734 (N_24734,N_23663,N_23326);
or U24735 (N_24735,N_23465,N_23420);
xor U24736 (N_24736,N_23509,N_22539);
or U24737 (N_24737,N_23064,N_23265);
and U24738 (N_24738,N_22646,N_22720);
xor U24739 (N_24739,N_23718,N_22783);
and U24740 (N_24740,N_23653,N_23734);
or U24741 (N_24741,N_22921,N_23313);
nor U24742 (N_24742,N_23664,N_23317);
xnor U24743 (N_24743,N_23263,N_23479);
and U24744 (N_24744,N_22699,N_23739);
xnor U24745 (N_24745,N_23493,N_23746);
nor U24746 (N_24746,N_22967,N_23689);
nor U24747 (N_24747,N_22936,N_22959);
and U24748 (N_24748,N_22708,N_23236);
nor U24749 (N_24749,N_23402,N_22878);
and U24750 (N_24750,N_23146,N_23719);
nand U24751 (N_24751,N_23223,N_22854);
xnor U24752 (N_24752,N_22776,N_23055);
nand U24753 (N_24753,N_23651,N_22702);
nand U24754 (N_24754,N_23159,N_23387);
nand U24755 (N_24755,N_23347,N_23155);
nor U24756 (N_24756,N_23437,N_22576);
or U24757 (N_24757,N_23749,N_23465);
and U24758 (N_24758,N_23717,N_23518);
xor U24759 (N_24759,N_22944,N_22604);
nor U24760 (N_24760,N_23705,N_23656);
or U24761 (N_24761,N_23125,N_22619);
xnor U24762 (N_24762,N_23187,N_22506);
or U24763 (N_24763,N_22878,N_22999);
xor U24764 (N_24764,N_22980,N_23387);
xor U24765 (N_24765,N_23380,N_23318);
xnor U24766 (N_24766,N_23262,N_22548);
or U24767 (N_24767,N_23267,N_23155);
and U24768 (N_24768,N_22845,N_23118);
and U24769 (N_24769,N_22782,N_23680);
or U24770 (N_24770,N_23481,N_23252);
and U24771 (N_24771,N_23337,N_23713);
or U24772 (N_24772,N_22636,N_22763);
and U24773 (N_24773,N_22889,N_23331);
nand U24774 (N_24774,N_23127,N_22568);
nand U24775 (N_24775,N_23003,N_23519);
xor U24776 (N_24776,N_23157,N_22835);
and U24777 (N_24777,N_22714,N_23377);
xor U24778 (N_24778,N_23210,N_22913);
nor U24779 (N_24779,N_23417,N_23229);
xor U24780 (N_24780,N_23207,N_23371);
xnor U24781 (N_24781,N_22874,N_23248);
xor U24782 (N_24782,N_23057,N_23496);
nand U24783 (N_24783,N_23169,N_22834);
or U24784 (N_24784,N_22866,N_23473);
or U24785 (N_24785,N_23392,N_22998);
xor U24786 (N_24786,N_22970,N_23115);
nand U24787 (N_24787,N_22989,N_23419);
nor U24788 (N_24788,N_22837,N_23179);
or U24789 (N_24789,N_23349,N_23497);
xor U24790 (N_24790,N_22950,N_23418);
nor U24791 (N_24791,N_23211,N_23673);
nand U24792 (N_24792,N_23316,N_22813);
or U24793 (N_24793,N_22855,N_23544);
or U24794 (N_24794,N_23203,N_23675);
and U24795 (N_24795,N_22736,N_22716);
nand U24796 (N_24796,N_22764,N_23126);
xnor U24797 (N_24797,N_22826,N_22614);
and U24798 (N_24798,N_22696,N_23507);
and U24799 (N_24799,N_23075,N_22859);
xor U24800 (N_24800,N_23073,N_23052);
nor U24801 (N_24801,N_22678,N_23522);
nand U24802 (N_24802,N_23600,N_23230);
and U24803 (N_24803,N_23720,N_23332);
nand U24804 (N_24804,N_22847,N_23476);
nor U24805 (N_24805,N_23107,N_23638);
or U24806 (N_24806,N_23464,N_23482);
nand U24807 (N_24807,N_22679,N_22883);
or U24808 (N_24808,N_22823,N_22727);
nor U24809 (N_24809,N_22767,N_22507);
nand U24810 (N_24810,N_23530,N_23119);
nor U24811 (N_24811,N_23291,N_23676);
nand U24812 (N_24812,N_22981,N_22810);
nand U24813 (N_24813,N_22609,N_23580);
and U24814 (N_24814,N_23414,N_23442);
xnor U24815 (N_24815,N_23626,N_23601);
nor U24816 (N_24816,N_23550,N_23269);
xnor U24817 (N_24817,N_22652,N_22900);
nand U24818 (N_24818,N_23688,N_23227);
and U24819 (N_24819,N_23171,N_22763);
nor U24820 (N_24820,N_23564,N_22890);
and U24821 (N_24821,N_22619,N_23042);
or U24822 (N_24822,N_23191,N_22683);
and U24823 (N_24823,N_23668,N_23073);
xor U24824 (N_24824,N_23535,N_22633);
and U24825 (N_24825,N_22732,N_22730);
or U24826 (N_24826,N_22598,N_23156);
or U24827 (N_24827,N_23253,N_23474);
nand U24828 (N_24828,N_22508,N_23640);
and U24829 (N_24829,N_22715,N_23022);
xnor U24830 (N_24830,N_23272,N_22931);
or U24831 (N_24831,N_22870,N_22700);
nand U24832 (N_24832,N_22732,N_23212);
nand U24833 (N_24833,N_23639,N_23019);
and U24834 (N_24834,N_23675,N_23481);
nor U24835 (N_24835,N_23192,N_22909);
or U24836 (N_24836,N_23567,N_22841);
nor U24837 (N_24837,N_22906,N_23339);
nor U24838 (N_24838,N_23164,N_23100);
nor U24839 (N_24839,N_22585,N_22535);
nand U24840 (N_24840,N_23084,N_23062);
xnor U24841 (N_24841,N_23150,N_22953);
nand U24842 (N_24842,N_23278,N_23329);
nand U24843 (N_24843,N_22866,N_22848);
or U24844 (N_24844,N_22926,N_23124);
or U24845 (N_24845,N_23075,N_23326);
and U24846 (N_24846,N_23576,N_23638);
nand U24847 (N_24847,N_23252,N_22742);
xnor U24848 (N_24848,N_22781,N_22858);
and U24849 (N_24849,N_22798,N_23670);
or U24850 (N_24850,N_23479,N_23052);
nand U24851 (N_24851,N_22551,N_23748);
nand U24852 (N_24852,N_23029,N_22754);
xor U24853 (N_24853,N_23018,N_23126);
or U24854 (N_24854,N_23249,N_22664);
xnor U24855 (N_24855,N_22696,N_23129);
and U24856 (N_24856,N_23564,N_22648);
nand U24857 (N_24857,N_23021,N_23443);
or U24858 (N_24858,N_23120,N_23006);
nand U24859 (N_24859,N_23317,N_23164);
nand U24860 (N_24860,N_22586,N_23326);
nand U24861 (N_24861,N_23149,N_22842);
nand U24862 (N_24862,N_22553,N_23015);
nand U24863 (N_24863,N_22759,N_23736);
xor U24864 (N_24864,N_22752,N_23033);
or U24865 (N_24865,N_23430,N_23359);
nand U24866 (N_24866,N_23599,N_23019);
nor U24867 (N_24867,N_23333,N_23075);
nand U24868 (N_24868,N_22787,N_22645);
xnor U24869 (N_24869,N_23130,N_23630);
nor U24870 (N_24870,N_22780,N_22969);
xor U24871 (N_24871,N_22810,N_23557);
nand U24872 (N_24872,N_23704,N_22707);
nand U24873 (N_24873,N_23599,N_23354);
and U24874 (N_24874,N_22783,N_23147);
and U24875 (N_24875,N_23319,N_22818);
xor U24876 (N_24876,N_22509,N_23471);
nand U24877 (N_24877,N_22517,N_22533);
nand U24878 (N_24878,N_22641,N_23549);
nor U24879 (N_24879,N_23270,N_23675);
and U24880 (N_24880,N_23266,N_23013);
or U24881 (N_24881,N_23390,N_23080);
or U24882 (N_24882,N_23008,N_22685);
nand U24883 (N_24883,N_22913,N_23302);
xnor U24884 (N_24884,N_23704,N_22531);
nand U24885 (N_24885,N_23445,N_22979);
or U24886 (N_24886,N_23386,N_22831);
nor U24887 (N_24887,N_23705,N_22998);
and U24888 (N_24888,N_23563,N_23564);
nand U24889 (N_24889,N_23401,N_23734);
or U24890 (N_24890,N_22523,N_23221);
or U24891 (N_24891,N_22602,N_23608);
nor U24892 (N_24892,N_22838,N_22967);
or U24893 (N_24893,N_23606,N_23636);
nand U24894 (N_24894,N_23296,N_22894);
nor U24895 (N_24895,N_23361,N_23340);
xnor U24896 (N_24896,N_22808,N_23442);
and U24897 (N_24897,N_23149,N_23055);
nand U24898 (N_24898,N_23515,N_23109);
or U24899 (N_24899,N_23639,N_22536);
nor U24900 (N_24900,N_22736,N_23506);
or U24901 (N_24901,N_22516,N_23424);
nand U24902 (N_24902,N_22916,N_23112);
nand U24903 (N_24903,N_23164,N_23177);
xor U24904 (N_24904,N_22915,N_23053);
nand U24905 (N_24905,N_23746,N_22517);
nand U24906 (N_24906,N_22704,N_22892);
nand U24907 (N_24907,N_22804,N_23616);
or U24908 (N_24908,N_23690,N_22723);
nor U24909 (N_24909,N_23107,N_23329);
or U24910 (N_24910,N_23266,N_22649);
nand U24911 (N_24911,N_22777,N_22897);
nand U24912 (N_24912,N_23193,N_23720);
and U24913 (N_24913,N_23088,N_23584);
or U24914 (N_24914,N_23028,N_22679);
nand U24915 (N_24915,N_22939,N_23444);
or U24916 (N_24916,N_23557,N_23240);
nand U24917 (N_24917,N_23183,N_23051);
or U24918 (N_24918,N_23685,N_22917);
nand U24919 (N_24919,N_22808,N_22855);
or U24920 (N_24920,N_22709,N_22518);
xnor U24921 (N_24921,N_23288,N_22907);
or U24922 (N_24922,N_22776,N_22922);
and U24923 (N_24923,N_22646,N_23685);
nand U24924 (N_24924,N_23037,N_22961);
nor U24925 (N_24925,N_22804,N_22815);
nor U24926 (N_24926,N_22801,N_23578);
nor U24927 (N_24927,N_22935,N_23588);
xor U24928 (N_24928,N_23627,N_23246);
nor U24929 (N_24929,N_22936,N_22502);
nand U24930 (N_24930,N_23419,N_22740);
and U24931 (N_24931,N_23209,N_23696);
or U24932 (N_24932,N_23228,N_23490);
or U24933 (N_24933,N_22725,N_22925);
nand U24934 (N_24934,N_22656,N_23272);
xnor U24935 (N_24935,N_23661,N_23322);
nor U24936 (N_24936,N_23078,N_23583);
xnor U24937 (N_24937,N_23664,N_23090);
xor U24938 (N_24938,N_22569,N_23693);
nor U24939 (N_24939,N_23465,N_23585);
or U24940 (N_24940,N_23562,N_22696);
and U24941 (N_24941,N_22651,N_22708);
or U24942 (N_24942,N_22778,N_23729);
xnor U24943 (N_24943,N_23741,N_22578);
nand U24944 (N_24944,N_23321,N_23284);
and U24945 (N_24945,N_22812,N_22942);
and U24946 (N_24946,N_22805,N_23043);
nand U24947 (N_24947,N_23045,N_23318);
nand U24948 (N_24948,N_22614,N_23099);
and U24949 (N_24949,N_23477,N_23374);
and U24950 (N_24950,N_23361,N_22664);
xnor U24951 (N_24951,N_23503,N_23725);
xnor U24952 (N_24952,N_23543,N_22575);
and U24953 (N_24953,N_23537,N_23277);
nand U24954 (N_24954,N_22831,N_23512);
or U24955 (N_24955,N_23235,N_22521);
xor U24956 (N_24956,N_23008,N_23036);
or U24957 (N_24957,N_22934,N_22832);
or U24958 (N_24958,N_22793,N_22605);
xor U24959 (N_24959,N_22688,N_22964);
nor U24960 (N_24960,N_22975,N_22896);
and U24961 (N_24961,N_23302,N_22659);
or U24962 (N_24962,N_23034,N_23636);
nand U24963 (N_24963,N_23281,N_22659);
xor U24964 (N_24964,N_23333,N_23350);
nand U24965 (N_24965,N_23439,N_23142);
nand U24966 (N_24966,N_23372,N_23204);
nand U24967 (N_24967,N_22998,N_23255);
xnor U24968 (N_24968,N_22574,N_23235);
nor U24969 (N_24969,N_23072,N_22926);
nor U24970 (N_24970,N_23004,N_22911);
and U24971 (N_24971,N_23029,N_22746);
and U24972 (N_24972,N_23567,N_23390);
nor U24973 (N_24973,N_23604,N_22577);
nor U24974 (N_24974,N_22525,N_22546);
or U24975 (N_24975,N_23005,N_22608);
xor U24976 (N_24976,N_23007,N_23707);
and U24977 (N_24977,N_23425,N_23517);
xnor U24978 (N_24978,N_22729,N_23657);
nand U24979 (N_24979,N_22904,N_23426);
and U24980 (N_24980,N_23037,N_23360);
xnor U24981 (N_24981,N_23403,N_23594);
xor U24982 (N_24982,N_23347,N_22783);
xor U24983 (N_24983,N_23671,N_22504);
nand U24984 (N_24984,N_23524,N_22553);
nor U24985 (N_24985,N_22746,N_22691);
or U24986 (N_24986,N_23747,N_23062);
xnor U24987 (N_24987,N_23614,N_23210);
and U24988 (N_24988,N_23279,N_23594);
nand U24989 (N_24989,N_23634,N_23637);
nand U24990 (N_24990,N_22742,N_23633);
nor U24991 (N_24991,N_22596,N_23705);
or U24992 (N_24992,N_23477,N_23111);
and U24993 (N_24993,N_22682,N_22923);
or U24994 (N_24994,N_23205,N_22567);
xnor U24995 (N_24995,N_23721,N_23524);
nor U24996 (N_24996,N_22586,N_22718);
and U24997 (N_24997,N_23338,N_23518);
and U24998 (N_24998,N_22809,N_23213);
and U24999 (N_24999,N_22705,N_22766);
and UO_0 (O_0,N_24798,N_24079);
xor UO_1 (O_1,N_23888,N_23852);
nand UO_2 (O_2,N_23963,N_24607);
and UO_3 (O_3,N_24669,N_23896);
nand UO_4 (O_4,N_24427,N_24791);
and UO_5 (O_5,N_24944,N_23926);
and UO_6 (O_6,N_24176,N_23804);
nor UO_7 (O_7,N_24747,N_24536);
nor UO_8 (O_8,N_24312,N_24450);
xnor UO_9 (O_9,N_24443,N_24012);
nand UO_10 (O_10,N_24453,N_24821);
and UO_11 (O_11,N_23948,N_24761);
and UO_12 (O_12,N_24721,N_24744);
nor UO_13 (O_13,N_24003,N_24413);
xor UO_14 (O_14,N_24974,N_24947);
xnor UO_15 (O_15,N_24618,N_23970);
and UO_16 (O_16,N_24781,N_24058);
and UO_17 (O_17,N_24817,N_24473);
nand UO_18 (O_18,N_23788,N_24051);
or UO_19 (O_19,N_24589,N_24709);
and UO_20 (O_20,N_24516,N_24188);
and UO_21 (O_21,N_24389,N_24895);
xor UO_22 (O_22,N_24004,N_24294);
and UO_23 (O_23,N_24788,N_24616);
xor UO_24 (O_24,N_24093,N_24907);
and UO_25 (O_25,N_24057,N_24769);
nor UO_26 (O_26,N_24503,N_24643);
and UO_27 (O_27,N_23791,N_24157);
xnor UO_28 (O_28,N_24298,N_24726);
and UO_29 (O_29,N_23934,N_24491);
nor UO_30 (O_30,N_24667,N_24455);
nor UO_31 (O_31,N_23812,N_24860);
and UO_32 (O_32,N_24594,N_24403);
or UO_33 (O_33,N_23995,N_24556);
and UO_34 (O_34,N_24644,N_24734);
nor UO_35 (O_35,N_23760,N_24840);
nand UO_36 (O_36,N_23997,N_24988);
and UO_37 (O_37,N_24710,N_24574);
xor UO_38 (O_38,N_24697,N_24303);
xor UO_39 (O_39,N_24893,N_24692);
and UO_40 (O_40,N_24320,N_24513);
and UO_41 (O_41,N_24489,N_23763);
or UO_42 (O_42,N_23814,N_24115);
and UO_43 (O_43,N_23778,N_24684);
nor UO_44 (O_44,N_24028,N_24000);
nor UO_45 (O_45,N_24421,N_24471);
nand UO_46 (O_46,N_24061,N_24066);
xnor UO_47 (O_47,N_24071,N_24475);
and UO_48 (O_48,N_24660,N_24689);
nand UO_49 (O_49,N_24903,N_24610);
or UO_50 (O_50,N_24016,N_23750);
nor UO_51 (O_51,N_24719,N_24756);
nand UO_52 (O_52,N_24933,N_24444);
or UO_53 (O_53,N_23858,N_24996);
or UO_54 (O_54,N_24477,N_23921);
nand UO_55 (O_55,N_24210,N_24577);
nand UO_56 (O_56,N_24573,N_24940);
nand UO_57 (O_57,N_23947,N_24950);
xor UO_58 (O_58,N_24131,N_24278);
nand UO_59 (O_59,N_23932,N_24199);
and UO_60 (O_60,N_24155,N_24168);
and UO_61 (O_61,N_23933,N_24982);
nand UO_62 (O_62,N_24038,N_24366);
nor UO_63 (O_63,N_24322,N_24362);
xor UO_64 (O_64,N_24775,N_24390);
nor UO_65 (O_65,N_24258,N_24263);
xnor UO_66 (O_66,N_24106,N_24136);
and UO_67 (O_67,N_24883,N_24158);
nand UO_68 (O_68,N_24122,N_24957);
or UO_69 (O_69,N_23936,N_24013);
and UO_70 (O_70,N_24955,N_23761);
or UO_71 (O_71,N_24546,N_24031);
or UO_72 (O_72,N_24463,N_24614);
and UO_73 (O_73,N_24025,N_24161);
xor UO_74 (O_74,N_23923,N_24792);
or UO_75 (O_75,N_24102,N_24454);
or UO_76 (O_76,N_24901,N_24581);
or UO_77 (O_77,N_23833,N_24623);
and UO_78 (O_78,N_23983,N_24178);
nand UO_79 (O_79,N_24027,N_23918);
nor UO_80 (O_80,N_24645,N_24172);
nor UO_81 (O_81,N_24074,N_24009);
nor UO_82 (O_82,N_24571,N_24805);
and UO_83 (O_83,N_24282,N_24945);
xor UO_84 (O_84,N_24241,N_24419);
xor UO_85 (O_85,N_24668,N_24807);
nand UO_86 (O_86,N_24356,N_24948);
and UO_87 (O_87,N_24409,N_24396);
and UO_88 (O_88,N_24240,N_24078);
nand UO_89 (O_89,N_23958,N_24209);
or UO_90 (O_90,N_23842,N_24711);
nor UO_91 (O_91,N_23895,N_23922);
xnor UO_92 (O_92,N_24002,N_24724);
nand UO_93 (O_93,N_24869,N_23952);
or UO_94 (O_94,N_23879,N_24208);
nor UO_95 (O_95,N_24867,N_24741);
and UO_96 (O_96,N_23767,N_24637);
and UO_97 (O_97,N_24297,N_23951);
xnor UO_98 (O_98,N_23903,N_23859);
nand UO_99 (O_99,N_24142,N_24946);
and UO_100 (O_100,N_24559,N_24024);
nand UO_101 (O_101,N_24108,N_23935);
nor UO_102 (O_102,N_23999,N_23953);
nand UO_103 (O_103,N_24773,N_24963);
nand UO_104 (O_104,N_24851,N_24561);
xor UO_105 (O_105,N_24519,N_24202);
xor UO_106 (O_106,N_23904,N_24796);
or UO_107 (O_107,N_24984,N_24152);
or UO_108 (O_108,N_24033,N_24921);
nor UO_109 (O_109,N_24395,N_24431);
or UO_110 (O_110,N_24306,N_24401);
nand UO_111 (O_111,N_24994,N_24225);
or UO_112 (O_112,N_24289,N_24254);
nand UO_113 (O_113,N_24968,N_24865);
nor UO_114 (O_114,N_24315,N_24731);
or UO_115 (O_115,N_24498,N_24888);
and UO_116 (O_116,N_24582,N_23775);
and UO_117 (O_117,N_24077,N_24457);
xor UO_118 (O_118,N_23940,N_24970);
or UO_119 (O_119,N_23831,N_24146);
nand UO_120 (O_120,N_23809,N_24462);
and UO_121 (O_121,N_24327,N_23773);
nand UO_122 (O_122,N_23962,N_24750);
or UO_123 (O_123,N_23803,N_24759);
or UO_124 (O_124,N_24999,N_24599);
and UO_125 (O_125,N_24232,N_24934);
nor UO_126 (O_126,N_24564,N_23768);
nor UO_127 (O_127,N_24174,N_23915);
and UO_128 (O_128,N_23880,N_24405);
xnor UO_129 (O_129,N_24195,N_24615);
nand UO_130 (O_130,N_24980,N_24590);
nand UO_131 (O_131,N_24149,N_24839);
nor UO_132 (O_132,N_24262,N_24110);
xnor UO_133 (O_133,N_23781,N_24835);
nor UO_134 (O_134,N_24735,N_24780);
nor UO_135 (O_135,N_24191,N_24635);
xor UO_136 (O_136,N_23798,N_24517);
and UO_137 (O_137,N_24100,N_23978);
or UO_138 (O_138,N_24993,N_23843);
xor UO_139 (O_139,N_24598,N_24636);
nor UO_140 (O_140,N_24797,N_24085);
nor UO_141 (O_141,N_24237,N_24430);
nor UO_142 (O_142,N_23982,N_24766);
xor UO_143 (O_143,N_24399,N_24221);
xnor UO_144 (O_144,N_24483,N_24808);
and UO_145 (O_145,N_24397,N_24165);
nor UO_146 (O_146,N_24460,N_24114);
nor UO_147 (O_147,N_24558,N_24246);
nand UO_148 (O_148,N_24526,N_24260);
or UO_149 (O_149,N_24505,N_23954);
nand UO_150 (O_150,N_24323,N_24586);
nand UO_151 (O_151,N_24981,N_24998);
xnor UO_152 (O_152,N_24416,N_23916);
or UO_153 (O_153,N_24676,N_23938);
or UO_154 (O_154,N_24374,N_23985);
or UO_155 (O_155,N_24657,N_24036);
nand UO_156 (O_156,N_24398,N_24153);
xor UO_157 (O_157,N_24605,N_23930);
nor UO_158 (O_158,N_24973,N_24552);
and UO_159 (O_159,N_24743,N_24482);
xor UO_160 (O_160,N_23974,N_24467);
xor UO_161 (O_161,N_24445,N_24509);
or UO_162 (O_162,N_24834,N_23980);
xor UO_163 (O_163,N_24705,N_24602);
or UO_164 (O_164,N_24717,N_24820);
or UO_165 (O_165,N_24704,N_23969);
and UO_166 (O_166,N_24273,N_24583);
and UO_167 (O_167,N_24341,N_23866);
nand UO_168 (O_168,N_24097,N_24287);
xnor UO_169 (O_169,N_24402,N_24037);
and UO_170 (O_170,N_24997,N_24017);
nor UO_171 (O_171,N_24307,N_24723);
and UO_172 (O_172,N_24065,N_24976);
nor UO_173 (O_173,N_24005,N_24107);
or UO_174 (O_174,N_23805,N_23876);
nand UO_175 (O_175,N_24548,N_24699);
nor UO_176 (O_176,N_24587,N_24141);
nand UO_177 (O_177,N_24674,N_24203);
nor UO_178 (O_178,N_24958,N_24338);
and UO_179 (O_179,N_24010,N_24420);
or UO_180 (O_180,N_24658,N_24528);
xor UO_181 (O_181,N_23841,N_24681);
xor UO_182 (O_182,N_24259,N_24139);
and UO_183 (O_183,N_24218,N_24889);
or UO_184 (O_184,N_23813,N_24291);
or UO_185 (O_185,N_24803,N_24795);
and UO_186 (O_186,N_23769,N_24529);
or UO_187 (O_187,N_24686,N_24228);
xor UO_188 (O_188,N_24328,N_23881);
nor UO_189 (O_189,N_24733,N_24638);
nor UO_190 (O_190,N_24170,N_24771);
or UO_191 (O_191,N_24147,N_24148);
nor UO_192 (O_192,N_24653,N_24140);
nor UO_193 (O_193,N_24922,N_24030);
or UO_194 (O_194,N_24633,N_23782);
nor UO_195 (O_195,N_23984,N_24479);
or UO_196 (O_196,N_24370,N_24631);
or UO_197 (O_197,N_24707,N_24732);
xnor UO_198 (O_198,N_23801,N_24861);
or UO_199 (O_199,N_24916,N_24729);
nor UO_200 (O_200,N_23939,N_23973);
and UO_201 (O_201,N_24779,N_24261);
and UO_202 (O_202,N_23942,N_23826);
or UO_203 (O_203,N_24299,N_24290);
nand UO_204 (O_204,N_24601,N_24035);
nor UO_205 (O_205,N_24608,N_24632);
xnor UO_206 (O_206,N_24964,N_24716);
nor UO_207 (O_207,N_24989,N_24512);
and UO_208 (O_208,N_24971,N_23802);
or UO_209 (O_209,N_24145,N_24569);
xnor UO_210 (O_210,N_24377,N_24991);
nor UO_211 (O_211,N_24647,N_24314);
xnor UO_212 (O_212,N_24350,N_24639);
or UO_213 (O_213,N_24422,N_23869);
and UO_214 (O_214,N_24696,N_23840);
nor UO_215 (O_215,N_24864,N_24234);
nor UO_216 (O_216,N_23764,N_24619);
nor UO_217 (O_217,N_24335,N_24047);
or UO_218 (O_218,N_23960,N_23865);
or UO_219 (O_219,N_24006,N_24281);
nand UO_220 (O_220,N_24083,N_23822);
and UO_221 (O_221,N_24393,N_24748);
nand UO_222 (O_222,N_23887,N_24504);
or UO_223 (O_223,N_24326,N_24810);
xor UO_224 (O_224,N_24470,N_23882);
and UO_225 (O_225,N_24032,N_23765);
or UO_226 (O_226,N_24109,N_24339);
xor UO_227 (O_227,N_24242,N_24793);
or UO_228 (O_228,N_24486,N_24845);
nand UO_229 (O_229,N_24132,N_24880);
and UO_230 (O_230,N_24391,N_24055);
nor UO_231 (O_231,N_24522,N_24833);
xor UO_232 (O_232,N_24159,N_24224);
nand UO_233 (O_233,N_24346,N_23968);
or UO_234 (O_234,N_24956,N_24103);
and UO_235 (O_235,N_24368,N_24112);
xnor UO_236 (O_236,N_24878,N_23821);
xnor UO_237 (O_237,N_24879,N_24364);
and UO_238 (O_238,N_24042,N_24160);
xnor UO_239 (O_239,N_24662,N_24424);
xor UO_240 (O_240,N_23956,N_24768);
nand UO_241 (O_241,N_24348,N_24321);
nor UO_242 (O_242,N_24011,N_24975);
nand UO_243 (O_243,N_23818,N_24099);
or UO_244 (O_244,N_24056,N_24856);
and UO_245 (O_245,N_24309,N_24270);
xor UO_246 (O_246,N_24836,N_23762);
xor UO_247 (O_247,N_23806,N_24511);
and UO_248 (O_248,N_24620,N_24238);
nand UO_249 (O_249,N_23850,N_24597);
xnor UO_250 (O_250,N_24182,N_24437);
and UO_251 (O_251,N_24824,N_24113);
and UO_252 (O_252,N_23911,N_23860);
xnor UO_253 (O_253,N_24245,N_24920);
or UO_254 (O_254,N_24310,N_24596);
and UO_255 (O_255,N_24641,N_24855);
nand UO_256 (O_256,N_23975,N_24818);
or UO_257 (O_257,N_24650,N_24926);
nand UO_258 (O_258,N_24340,N_24537);
or UO_259 (O_259,N_24806,N_23941);
xor UO_260 (O_260,N_24720,N_23910);
nor UO_261 (O_261,N_23885,N_23898);
nand UO_262 (O_262,N_24654,N_24352);
nand UO_263 (O_263,N_24205,N_23851);
and UO_264 (O_264,N_24737,N_24677);
nand UO_265 (O_265,N_24854,N_24767);
nand UO_266 (O_266,N_24969,N_24624);
nand UO_267 (O_267,N_24930,N_24995);
nor UO_268 (O_268,N_24815,N_24685);
nor UO_269 (O_269,N_24630,N_24318);
nor UO_270 (O_270,N_23823,N_23971);
nor UO_271 (O_271,N_24698,N_24887);
nor UO_272 (O_272,N_24871,N_24502);
nor UO_273 (O_273,N_23884,N_23830);
nor UO_274 (O_274,N_24541,N_23785);
or UO_275 (O_275,N_24844,N_24611);
nand UO_276 (O_276,N_24184,N_24466);
nor UO_277 (O_277,N_24876,N_24757);
nand UO_278 (O_278,N_24841,N_24754);
xnor UO_279 (O_279,N_23987,N_24900);
xnor UO_280 (O_280,N_24215,N_24219);
xnor UO_281 (O_281,N_23966,N_24019);
and UO_282 (O_282,N_24177,N_24800);
and UO_283 (O_283,N_24799,N_24150);
or UO_284 (O_284,N_24156,N_24388);
nand UO_285 (O_285,N_24591,N_24333);
nor UO_286 (O_286,N_24648,N_24764);
or UO_287 (O_287,N_24008,N_24084);
nand UO_288 (O_288,N_24041,N_23981);
nand UO_289 (O_289,N_24830,N_24429);
xnor UO_290 (O_290,N_23990,N_24274);
xor UO_291 (O_291,N_24763,N_24915);
and UO_292 (O_292,N_24337,N_24386);
nand UO_293 (O_293,N_24555,N_24300);
or UO_294 (O_294,N_23752,N_24557);
or UO_295 (O_295,N_23796,N_23862);
and UO_296 (O_296,N_23874,N_24465);
or UO_297 (O_297,N_24311,N_24007);
and UO_298 (O_298,N_24656,N_24565);
xor UO_299 (O_299,N_24360,N_23836);
nor UO_300 (O_300,N_23756,N_24069);
nor UO_301 (O_301,N_24544,N_24135);
or UO_302 (O_302,N_24411,N_24862);
nand UO_303 (O_303,N_23899,N_24595);
nand UO_304 (O_304,N_24250,N_24527);
xnor UO_305 (O_305,N_23955,N_24436);
and UO_306 (O_306,N_24123,N_24313);
xor UO_307 (O_307,N_24938,N_24089);
nor UO_308 (O_308,N_24521,N_24910);
nor UO_309 (O_309,N_24917,N_24914);
xor UO_310 (O_310,N_23811,N_24380);
or UO_311 (O_311,N_24562,N_24464);
and UO_312 (O_312,N_24593,N_24972);
xor UO_313 (O_313,N_23846,N_24050);
xnor UO_314 (O_314,N_24943,N_24813);
xnor UO_315 (O_315,N_24325,N_24739);
nand UO_316 (O_316,N_24253,N_24449);
nor UO_317 (O_317,N_24899,N_24022);
nand UO_318 (O_318,N_24354,N_23871);
nor UO_319 (O_319,N_24746,N_24954);
xnor UO_320 (O_320,N_24180,N_23996);
and UO_321 (O_321,N_24098,N_24912);
and UO_322 (O_322,N_24230,N_24279);
xor UO_323 (O_323,N_24469,N_24925);
nand UO_324 (O_324,N_24343,N_24052);
xor UO_325 (O_325,N_24220,N_24540);
and UO_326 (O_326,N_24823,N_24183);
nand UO_327 (O_327,N_24592,N_24217);
nor UO_328 (O_328,N_24134,N_24962);
and UO_329 (O_329,N_23766,N_24932);
nor UO_330 (O_330,N_24295,N_23931);
nand UO_331 (O_331,N_24096,N_24138);
xor UO_332 (O_332,N_24837,N_24931);
nor UO_333 (O_333,N_24683,N_24927);
nand UO_334 (O_334,N_23817,N_24829);
nand UO_335 (O_335,N_24266,N_24197);
or UO_336 (O_336,N_23861,N_24550);
and UO_337 (O_337,N_23891,N_23794);
nor UO_338 (O_338,N_24870,N_24929);
nand UO_339 (O_339,N_24407,N_24578);
nor UO_340 (O_340,N_24367,N_23815);
xnor UO_341 (O_341,N_23901,N_23946);
nand UO_342 (O_342,N_24935,N_24257);
and UO_343 (O_343,N_24133,N_24301);
or UO_344 (O_344,N_24353,N_24501);
and UO_345 (O_345,N_23993,N_24198);
or UO_346 (O_346,N_24143,N_24678);
and UO_347 (O_347,N_24695,N_24227);
xor UO_348 (O_348,N_24488,N_24394);
and UO_349 (O_349,N_24977,N_23890);
nor UO_350 (O_350,N_23949,N_24939);
nand UO_351 (O_351,N_24722,N_24440);
xor UO_352 (O_352,N_24979,N_24244);
and UO_353 (O_353,N_23967,N_24873);
xor UO_354 (O_354,N_24378,N_24179);
nand UO_355 (O_355,N_24777,N_24786);
or UO_356 (O_356,N_24832,N_24673);
or UO_357 (O_357,N_24474,N_24866);
nor UO_358 (O_358,N_24770,N_24015);
xor UO_359 (O_359,N_24566,N_24116);
nor UO_360 (O_360,N_24524,N_24271);
xnor UO_361 (O_361,N_24908,N_24852);
and UO_362 (O_362,N_24809,N_24130);
and UO_363 (O_363,N_24949,N_24120);
nand UO_364 (O_364,N_24772,N_24308);
xnor UO_365 (O_365,N_24252,N_24428);
or UO_366 (O_366,N_23827,N_23800);
or UO_367 (O_367,N_24026,N_24822);
xnor UO_368 (O_368,N_24542,N_24048);
or UO_369 (O_369,N_24942,N_24649);
nand UO_370 (O_370,N_24406,N_24890);
xnor UO_371 (O_371,N_24062,N_24622);
or UO_372 (O_372,N_24236,N_23902);
nor UO_373 (O_373,N_23770,N_23906);
and UO_374 (O_374,N_24603,N_24909);
nor UO_375 (O_375,N_23959,N_23897);
nor UO_376 (O_376,N_24213,N_23784);
xor UO_377 (O_377,N_23816,N_24500);
or UO_378 (O_378,N_23937,N_24408);
or UO_379 (O_379,N_23912,N_24790);
xnor UO_380 (O_380,N_24941,N_24627);
xor UO_381 (O_381,N_23920,N_23789);
or UO_382 (O_382,N_23844,N_24877);
xor UO_383 (O_383,N_24251,N_24691);
or UO_384 (O_384,N_24714,N_24264);
and UO_385 (O_385,N_24186,N_24441);
xor UO_386 (O_386,N_24609,N_23799);
nor UO_387 (O_387,N_24296,N_24898);
xor UO_388 (O_388,N_23790,N_24802);
or UO_389 (O_389,N_23807,N_24478);
nor UO_390 (O_390,N_23964,N_24572);
and UO_391 (O_391,N_24514,N_24842);
and UO_392 (O_392,N_24304,N_23927);
or UO_393 (O_393,N_24382,N_24285);
xnor UO_394 (O_394,N_24438,N_24670);
nor UO_395 (O_395,N_24742,N_24359);
xor UO_396 (O_396,N_24214,N_24095);
nand UO_397 (O_397,N_24532,N_23925);
and UO_398 (O_398,N_24919,N_24092);
nand UO_399 (O_399,N_24936,N_23839);
nor UO_400 (O_400,N_24570,N_24881);
nand UO_401 (O_401,N_24439,N_24425);
or UO_402 (O_402,N_24499,N_24211);
nor UO_403 (O_403,N_24828,N_24575);
nand UO_404 (O_404,N_24495,N_23873);
or UO_405 (O_405,N_24280,N_24715);
and UO_406 (O_406,N_24316,N_24204);
nor UO_407 (O_407,N_24520,N_23758);
nor UO_408 (O_408,N_24167,N_24730);
xor UO_409 (O_409,N_24187,N_23992);
xor UO_410 (O_410,N_24690,N_24530);
xnor UO_411 (O_411,N_24154,N_24345);
and UO_412 (O_412,N_24459,N_24072);
nor UO_413 (O_413,N_24554,N_24535);
nand UO_414 (O_414,N_24302,N_24090);
and UO_415 (O_415,N_24358,N_24196);
nand UO_416 (O_416,N_23832,N_23998);
nand UO_417 (O_417,N_24200,N_24646);
nor UO_418 (O_418,N_24442,N_24319);
and UO_419 (O_419,N_24882,N_23777);
nor UO_420 (O_420,N_24848,N_24361);
and UO_421 (O_421,N_24913,N_24105);
xnor UO_422 (O_422,N_24787,N_24468);
or UO_423 (O_423,N_24905,N_24175);
nand UO_424 (O_424,N_24543,N_24412);
nand UO_425 (O_425,N_24563,N_24021);
xor UO_426 (O_426,N_23924,N_23919);
xor UO_427 (O_427,N_24446,N_24703);
nand UO_428 (O_428,N_24672,N_23838);
xor UO_429 (O_429,N_24659,N_24904);
nor UO_430 (O_430,N_23976,N_24604);
xor UO_431 (O_431,N_24081,N_24189);
or UO_432 (O_432,N_24222,N_24018);
nor UO_433 (O_433,N_24827,N_24265);
xor UO_434 (O_434,N_24118,N_24451);
or UO_435 (O_435,N_24060,N_24125);
nand UO_436 (O_436,N_24275,N_24447);
nand UO_437 (O_437,N_24054,N_24288);
xnor UO_438 (O_438,N_24235,N_24902);
xor UO_439 (O_439,N_24738,N_23870);
and UO_440 (O_440,N_23853,N_24070);
and UO_441 (O_441,N_24712,N_24371);
or UO_442 (O_442,N_24986,N_24753);
xnor UO_443 (O_443,N_24363,N_24694);
and UO_444 (O_444,N_24838,N_23849);
xor UO_445 (O_445,N_24978,N_24063);
and UO_446 (O_446,N_23786,N_24101);
xnor UO_447 (O_447,N_24082,N_23759);
xor UO_448 (O_448,N_24560,N_24494);
xor UO_449 (O_449,N_24992,N_24020);
nor UO_450 (O_450,N_23751,N_24506);
or UO_451 (O_451,N_24128,N_24508);
or UO_452 (O_452,N_23783,N_24664);
and UO_453 (O_453,N_24347,N_24379);
xnor UO_454 (O_454,N_24736,N_24727);
nor UO_455 (O_455,N_24706,N_24249);
nand UO_456 (O_456,N_24785,N_24765);
xor UO_457 (O_457,N_24682,N_24029);
nor UO_458 (O_458,N_24523,N_24661);
and UO_459 (O_459,N_24617,N_23894);
xor UO_460 (O_460,N_23872,N_24372);
xnor UO_461 (O_461,N_23771,N_23988);
xnor UO_462 (O_462,N_24385,N_24344);
nor UO_463 (O_463,N_24718,N_24671);
xor UO_464 (O_464,N_24216,N_24376);
xnor UO_465 (O_465,N_24126,N_23864);
xnor UO_466 (O_466,N_24192,N_24434);
and UO_467 (O_467,N_24846,N_24663);
and UO_468 (O_468,N_24740,N_24655);
and UO_469 (O_469,N_24534,N_24080);
or UO_470 (O_470,N_24190,N_24952);
and UO_471 (O_471,N_24276,N_24497);
or UO_472 (O_472,N_24875,N_24336);
xnor UO_473 (O_473,N_24417,N_24960);
nor UO_474 (O_474,N_24819,N_23845);
xor UO_475 (O_475,N_24194,N_24169);
or UO_476 (O_476,N_24868,N_24816);
nor UO_477 (O_477,N_23779,N_24928);
xnor UO_478 (O_478,N_24044,N_24001);
nand UO_479 (O_479,N_23854,N_23857);
xor UO_480 (O_480,N_24783,N_24243);
or UO_481 (O_481,N_23917,N_24277);
or UO_482 (O_482,N_24119,N_24383);
or UO_483 (O_483,N_24104,N_24384);
and UO_484 (O_484,N_23905,N_23979);
or UO_485 (O_485,N_24452,N_23950);
nor UO_486 (O_486,N_24373,N_23886);
or UO_487 (O_487,N_23757,N_24349);
xor UO_488 (O_488,N_24375,N_24127);
and UO_489 (O_489,N_24634,N_24778);
and UO_490 (O_490,N_24111,N_24164);
and UO_491 (O_491,N_24525,N_24687);
xor UO_492 (O_492,N_23893,N_24226);
xor UO_493 (O_493,N_24351,N_24043);
nor UO_494 (O_494,N_23994,N_24531);
nor UO_495 (O_495,N_24567,N_24539);
or UO_496 (O_496,N_24863,N_24162);
and UO_497 (O_497,N_23977,N_23848);
or UO_498 (O_498,N_24269,N_24496);
nand UO_499 (O_499,N_24688,N_24814);
nor UO_500 (O_500,N_24458,N_23908);
nand UO_501 (O_501,N_23957,N_24064);
nor UO_502 (O_502,N_23913,N_24959);
nand UO_503 (O_503,N_24752,N_24621);
and UO_504 (O_504,N_24897,N_24924);
and UO_505 (O_505,N_24576,N_24894);
nor UO_506 (O_506,N_24987,N_23868);
nand UO_507 (O_507,N_23835,N_24223);
and UO_508 (O_508,N_24293,N_24751);
or UO_509 (O_509,N_23755,N_23909);
nand UO_510 (O_510,N_24518,N_23834);
or UO_511 (O_511,N_23847,N_24515);
nand UO_512 (O_512,N_24357,N_23961);
nor UO_513 (O_513,N_24794,N_24255);
nor UO_514 (O_514,N_24843,N_24549);
nand UO_515 (O_515,N_23819,N_23797);
and UO_516 (O_516,N_24825,N_24625);
and UO_517 (O_517,N_24283,N_24423);
and UO_518 (O_518,N_23772,N_24324);
xor UO_519 (O_519,N_24911,N_24680);
nor UO_520 (O_520,N_24966,N_24045);
nor UO_521 (O_521,N_23776,N_24053);
xnor UO_522 (O_522,N_23829,N_24049);
nand UO_523 (O_523,N_24233,N_24039);
nor UO_524 (O_524,N_24585,N_23855);
or UO_525 (O_525,N_24642,N_24268);
xnor UO_526 (O_526,N_24404,N_24811);
and UO_527 (O_527,N_24481,N_24923);
and UO_528 (O_528,N_23892,N_24068);
xnor UO_529 (O_529,N_24612,N_24801);
and UO_530 (O_530,N_24628,N_24144);
xnor UO_531 (O_531,N_24201,N_23863);
and UO_532 (O_532,N_24713,N_24762);
or UO_533 (O_533,N_24046,N_23900);
nor UO_534 (O_534,N_24831,N_23972);
and UO_535 (O_535,N_23991,N_24884);
xor UO_536 (O_536,N_24588,N_24284);
and UO_537 (O_537,N_24472,N_23824);
or UO_538 (O_538,N_24967,N_24342);
nor UO_539 (O_539,N_24749,N_24129);
and UO_540 (O_540,N_24426,N_24094);
nand UO_541 (O_541,N_23792,N_24305);
or UO_542 (O_542,N_24675,N_24490);
nor UO_543 (O_543,N_23914,N_23780);
xor UO_544 (O_544,N_24332,N_24414);
nand UO_545 (O_545,N_24418,N_24784);
nor UO_546 (O_546,N_23856,N_24181);
xor UO_547 (O_547,N_24448,N_24387);
nor UO_548 (O_548,N_24073,N_24510);
xnor UO_549 (O_549,N_24415,N_24076);
or UO_550 (O_550,N_24613,N_24480);
nand UO_551 (O_551,N_24492,N_24651);
and UO_552 (O_552,N_24185,N_24745);
and UO_553 (O_553,N_24606,N_24693);
xnor UO_554 (O_554,N_24476,N_24137);
nand UO_555 (O_555,N_24331,N_24826);
nand UO_556 (O_556,N_24568,N_24317);
or UO_557 (O_557,N_24918,N_24906);
or UO_558 (O_558,N_24075,N_24166);
xnor UO_559 (O_559,N_23989,N_23965);
or UO_560 (O_560,N_24121,N_23877);
or UO_561 (O_561,N_24087,N_23867);
and UO_562 (O_562,N_24758,N_24891);
or UO_563 (O_563,N_23986,N_24990);
nor UO_564 (O_564,N_24626,N_24961);
or UO_565 (O_565,N_24725,N_24040);
and UO_566 (O_566,N_24533,N_24484);
and UO_567 (O_567,N_24239,N_24124);
xnor UO_568 (O_568,N_24088,N_24435);
nand UO_569 (O_569,N_24173,N_24776);
nor UO_570 (O_570,N_23810,N_24171);
and UO_571 (O_571,N_23787,N_24885);
nand UO_572 (O_572,N_24163,N_24728);
xnor UO_573 (O_573,N_24059,N_24292);
xnor UO_574 (O_574,N_23774,N_24701);
nor UO_575 (O_575,N_24272,N_24507);
and UO_576 (O_576,N_24229,N_24086);
nor UO_577 (O_577,N_24896,N_24789);
and UO_578 (O_578,N_24551,N_24151);
or UO_579 (O_579,N_23828,N_23875);
nand UO_580 (O_580,N_24334,N_23929);
or UO_581 (O_581,N_24708,N_24652);
nor UO_582 (O_582,N_24247,N_24206);
xor UO_583 (O_583,N_24755,N_24760);
xnor UO_584 (O_584,N_24392,N_24937);
nand UO_585 (O_585,N_23878,N_24212);
nor UO_586 (O_586,N_24953,N_23825);
nand UO_587 (O_587,N_24547,N_24872);
nor UO_588 (O_588,N_23945,N_24433);
nand UO_589 (O_589,N_24983,N_23793);
and UO_590 (O_590,N_23944,N_23837);
or UO_591 (O_591,N_23820,N_24355);
and UO_592 (O_592,N_24410,N_24640);
and UO_593 (O_593,N_24329,N_24485);
nand UO_594 (O_594,N_24487,N_23889);
or UO_595 (O_595,N_23883,N_24965);
and UO_596 (O_596,N_24286,N_23754);
and UO_597 (O_597,N_24014,N_24267);
and UO_598 (O_598,N_24985,N_24886);
nor UO_599 (O_599,N_24849,N_24369);
and UO_600 (O_600,N_24330,N_24207);
nand UO_601 (O_601,N_24117,N_24665);
nand UO_602 (O_602,N_24702,N_24853);
nor UO_603 (O_603,N_24091,N_23943);
and UO_604 (O_604,N_23907,N_24847);
nor UO_605 (O_605,N_24600,N_24679);
or UO_606 (O_606,N_24951,N_24629);
and UO_607 (O_607,N_24256,N_24774);
xor UO_608 (O_608,N_24700,N_23808);
or UO_609 (O_609,N_23795,N_24545);
xnor UO_610 (O_610,N_24858,N_24857);
nand UO_611 (O_611,N_24365,N_24493);
xnor UO_612 (O_612,N_24584,N_23928);
nor UO_613 (O_613,N_23753,N_24023);
nand UO_614 (O_614,N_24553,N_24892);
and UO_615 (O_615,N_24381,N_24400);
nand UO_616 (O_616,N_24193,N_24538);
or UO_617 (O_617,N_24034,N_24850);
xnor UO_618 (O_618,N_24859,N_24804);
nor UO_619 (O_619,N_24067,N_24432);
nand UO_620 (O_620,N_24580,N_24782);
or UO_621 (O_621,N_24579,N_24461);
nand UO_622 (O_622,N_24456,N_24874);
and UO_623 (O_623,N_24812,N_24231);
xor UO_624 (O_624,N_24248,N_24666);
or UO_625 (O_625,N_24486,N_24973);
nand UO_626 (O_626,N_23811,N_24996);
and UO_627 (O_627,N_24063,N_24053);
and UO_628 (O_628,N_24959,N_23867);
or UO_629 (O_629,N_24723,N_24151);
xor UO_630 (O_630,N_24201,N_24220);
xnor UO_631 (O_631,N_24753,N_24101);
or UO_632 (O_632,N_23999,N_24594);
or UO_633 (O_633,N_24677,N_24199);
or UO_634 (O_634,N_24522,N_24886);
nor UO_635 (O_635,N_24604,N_24459);
xor UO_636 (O_636,N_24036,N_24334);
nand UO_637 (O_637,N_24330,N_23781);
nand UO_638 (O_638,N_24302,N_24646);
xnor UO_639 (O_639,N_24854,N_24362);
nor UO_640 (O_640,N_24426,N_24111);
nand UO_641 (O_641,N_24908,N_23878);
or UO_642 (O_642,N_24697,N_24848);
xnor UO_643 (O_643,N_24665,N_23785);
or UO_644 (O_644,N_24085,N_24597);
nor UO_645 (O_645,N_23762,N_24426);
and UO_646 (O_646,N_24332,N_24198);
nand UO_647 (O_647,N_24846,N_24237);
xnor UO_648 (O_648,N_23863,N_24104);
xor UO_649 (O_649,N_24054,N_23922);
xor UO_650 (O_650,N_24141,N_23940);
nand UO_651 (O_651,N_23799,N_24269);
xnor UO_652 (O_652,N_24640,N_24453);
or UO_653 (O_653,N_24423,N_24170);
nand UO_654 (O_654,N_24254,N_24738);
nand UO_655 (O_655,N_24011,N_24724);
or UO_656 (O_656,N_24373,N_23763);
xor UO_657 (O_657,N_24841,N_24077);
and UO_658 (O_658,N_23791,N_24120);
nand UO_659 (O_659,N_24209,N_24302);
and UO_660 (O_660,N_24264,N_24818);
xor UO_661 (O_661,N_23810,N_23814);
and UO_662 (O_662,N_24695,N_24873);
nand UO_663 (O_663,N_24742,N_24415);
or UO_664 (O_664,N_24070,N_24922);
or UO_665 (O_665,N_24986,N_23826);
and UO_666 (O_666,N_24759,N_24914);
nand UO_667 (O_667,N_24028,N_24470);
or UO_668 (O_668,N_24496,N_23791);
and UO_669 (O_669,N_24467,N_24205);
nor UO_670 (O_670,N_24887,N_24083);
or UO_671 (O_671,N_24433,N_23750);
and UO_672 (O_672,N_24221,N_24368);
nor UO_673 (O_673,N_24980,N_24876);
nor UO_674 (O_674,N_24465,N_24655);
xor UO_675 (O_675,N_24885,N_24703);
xnor UO_676 (O_676,N_24541,N_24311);
or UO_677 (O_677,N_24315,N_24721);
and UO_678 (O_678,N_24291,N_24045);
and UO_679 (O_679,N_24167,N_24288);
and UO_680 (O_680,N_23892,N_23905);
and UO_681 (O_681,N_24055,N_24957);
xor UO_682 (O_682,N_24977,N_24414);
or UO_683 (O_683,N_24107,N_24283);
nor UO_684 (O_684,N_24180,N_23814);
and UO_685 (O_685,N_24154,N_24036);
and UO_686 (O_686,N_24530,N_24115);
xnor UO_687 (O_687,N_23752,N_24885);
xnor UO_688 (O_688,N_23809,N_24266);
or UO_689 (O_689,N_24138,N_24836);
xnor UO_690 (O_690,N_24063,N_24259);
nor UO_691 (O_691,N_24369,N_24473);
nor UO_692 (O_692,N_23872,N_23862);
nor UO_693 (O_693,N_24806,N_24927);
nor UO_694 (O_694,N_24766,N_24230);
nor UO_695 (O_695,N_24830,N_24618);
nor UO_696 (O_696,N_23783,N_24864);
or UO_697 (O_697,N_24100,N_23861);
xor UO_698 (O_698,N_24689,N_23816);
or UO_699 (O_699,N_23842,N_24297);
nor UO_700 (O_700,N_24872,N_24362);
xor UO_701 (O_701,N_24041,N_24603);
or UO_702 (O_702,N_23851,N_24116);
or UO_703 (O_703,N_24616,N_23993);
or UO_704 (O_704,N_24630,N_24485);
nand UO_705 (O_705,N_24737,N_24117);
xor UO_706 (O_706,N_23987,N_23846);
or UO_707 (O_707,N_24263,N_24165);
nand UO_708 (O_708,N_23826,N_24521);
nand UO_709 (O_709,N_24129,N_23770);
or UO_710 (O_710,N_24616,N_24348);
or UO_711 (O_711,N_23905,N_24363);
or UO_712 (O_712,N_24198,N_24834);
xnor UO_713 (O_713,N_23960,N_23754);
nand UO_714 (O_714,N_24404,N_24350);
nand UO_715 (O_715,N_24782,N_24469);
and UO_716 (O_716,N_24617,N_23783);
nor UO_717 (O_717,N_23936,N_24482);
xor UO_718 (O_718,N_24777,N_24312);
xnor UO_719 (O_719,N_24293,N_24260);
xnor UO_720 (O_720,N_24142,N_24467);
and UO_721 (O_721,N_24368,N_24202);
or UO_722 (O_722,N_24763,N_24266);
and UO_723 (O_723,N_24562,N_24004);
nand UO_724 (O_724,N_24820,N_23900);
nor UO_725 (O_725,N_24244,N_24534);
xnor UO_726 (O_726,N_24706,N_24993);
nor UO_727 (O_727,N_24309,N_23782);
or UO_728 (O_728,N_24959,N_24690);
xnor UO_729 (O_729,N_24618,N_24982);
or UO_730 (O_730,N_24550,N_24964);
and UO_731 (O_731,N_24517,N_24002);
nand UO_732 (O_732,N_24256,N_23856);
nand UO_733 (O_733,N_24246,N_24916);
nor UO_734 (O_734,N_23946,N_23909);
and UO_735 (O_735,N_24596,N_24482);
and UO_736 (O_736,N_24007,N_24216);
xnor UO_737 (O_737,N_24187,N_24432);
and UO_738 (O_738,N_24502,N_24192);
nor UO_739 (O_739,N_24702,N_24097);
and UO_740 (O_740,N_24389,N_24377);
and UO_741 (O_741,N_24678,N_24472);
and UO_742 (O_742,N_24731,N_24735);
and UO_743 (O_743,N_24346,N_24311);
nor UO_744 (O_744,N_24642,N_24680);
or UO_745 (O_745,N_24067,N_24586);
nand UO_746 (O_746,N_24663,N_24251);
and UO_747 (O_747,N_23870,N_24839);
and UO_748 (O_748,N_24067,N_23974);
nor UO_749 (O_749,N_24362,N_23996);
nor UO_750 (O_750,N_24904,N_24066);
and UO_751 (O_751,N_23912,N_24090);
or UO_752 (O_752,N_24250,N_24456);
and UO_753 (O_753,N_23938,N_24657);
and UO_754 (O_754,N_24333,N_24773);
nand UO_755 (O_755,N_24410,N_24304);
nor UO_756 (O_756,N_23769,N_23882);
or UO_757 (O_757,N_24385,N_24247);
or UO_758 (O_758,N_24948,N_23769);
xnor UO_759 (O_759,N_24495,N_24422);
nor UO_760 (O_760,N_23902,N_24483);
nor UO_761 (O_761,N_24839,N_23934);
and UO_762 (O_762,N_24094,N_24559);
nor UO_763 (O_763,N_24911,N_24073);
or UO_764 (O_764,N_24671,N_24171);
xor UO_765 (O_765,N_24062,N_24849);
or UO_766 (O_766,N_24549,N_23868);
xnor UO_767 (O_767,N_23879,N_23769);
xnor UO_768 (O_768,N_23805,N_24239);
or UO_769 (O_769,N_24029,N_24932);
or UO_770 (O_770,N_23869,N_23850);
or UO_771 (O_771,N_23925,N_24810);
and UO_772 (O_772,N_24538,N_24990);
and UO_773 (O_773,N_24799,N_24665);
xnor UO_774 (O_774,N_23937,N_24052);
and UO_775 (O_775,N_23882,N_24866);
or UO_776 (O_776,N_24519,N_23923);
or UO_777 (O_777,N_24775,N_24444);
xor UO_778 (O_778,N_24881,N_24967);
nor UO_779 (O_779,N_23916,N_24354);
xnor UO_780 (O_780,N_24212,N_23825);
xnor UO_781 (O_781,N_24204,N_23802);
xnor UO_782 (O_782,N_24857,N_24118);
nor UO_783 (O_783,N_23943,N_24683);
nand UO_784 (O_784,N_24954,N_24609);
xnor UO_785 (O_785,N_24885,N_24926);
or UO_786 (O_786,N_24866,N_23780);
or UO_787 (O_787,N_24010,N_24532);
nand UO_788 (O_788,N_24977,N_24445);
and UO_789 (O_789,N_23987,N_23974);
xor UO_790 (O_790,N_24078,N_23892);
nand UO_791 (O_791,N_24220,N_24983);
and UO_792 (O_792,N_24996,N_24189);
nand UO_793 (O_793,N_24832,N_24397);
nor UO_794 (O_794,N_24628,N_24068);
and UO_795 (O_795,N_24010,N_24620);
nand UO_796 (O_796,N_24818,N_24166);
or UO_797 (O_797,N_24753,N_24203);
or UO_798 (O_798,N_24858,N_24556);
nor UO_799 (O_799,N_24418,N_24265);
or UO_800 (O_800,N_23980,N_24327);
nand UO_801 (O_801,N_24098,N_24904);
or UO_802 (O_802,N_23791,N_24882);
or UO_803 (O_803,N_24113,N_24880);
and UO_804 (O_804,N_23839,N_24084);
or UO_805 (O_805,N_24482,N_24071);
xor UO_806 (O_806,N_23824,N_24031);
nand UO_807 (O_807,N_24893,N_24251);
and UO_808 (O_808,N_23836,N_23909);
xnor UO_809 (O_809,N_24890,N_24830);
and UO_810 (O_810,N_24671,N_23910);
xnor UO_811 (O_811,N_23950,N_23929);
nand UO_812 (O_812,N_23945,N_24495);
or UO_813 (O_813,N_24830,N_24245);
nor UO_814 (O_814,N_24619,N_23888);
nor UO_815 (O_815,N_24588,N_24501);
and UO_816 (O_816,N_24530,N_24851);
or UO_817 (O_817,N_24580,N_24522);
or UO_818 (O_818,N_24347,N_24967);
or UO_819 (O_819,N_24569,N_24177);
nand UO_820 (O_820,N_24244,N_23837);
nand UO_821 (O_821,N_24444,N_24024);
or UO_822 (O_822,N_24572,N_24026);
nor UO_823 (O_823,N_24800,N_23844);
or UO_824 (O_824,N_24249,N_24340);
or UO_825 (O_825,N_24841,N_23887);
xor UO_826 (O_826,N_23986,N_24066);
and UO_827 (O_827,N_23797,N_24732);
and UO_828 (O_828,N_23938,N_23782);
or UO_829 (O_829,N_24258,N_24443);
xor UO_830 (O_830,N_24111,N_24219);
and UO_831 (O_831,N_24188,N_24154);
and UO_832 (O_832,N_24164,N_24125);
and UO_833 (O_833,N_23955,N_23855);
or UO_834 (O_834,N_24687,N_24994);
nand UO_835 (O_835,N_24475,N_23908);
nand UO_836 (O_836,N_23941,N_24530);
nand UO_837 (O_837,N_23870,N_24737);
nor UO_838 (O_838,N_23944,N_24725);
or UO_839 (O_839,N_24067,N_23832);
or UO_840 (O_840,N_24365,N_24350);
or UO_841 (O_841,N_23953,N_23885);
or UO_842 (O_842,N_24363,N_24960);
xor UO_843 (O_843,N_24838,N_23794);
xor UO_844 (O_844,N_24847,N_24759);
nor UO_845 (O_845,N_24442,N_23963);
xor UO_846 (O_846,N_24528,N_24891);
or UO_847 (O_847,N_24711,N_23958);
nand UO_848 (O_848,N_24002,N_24567);
nor UO_849 (O_849,N_24583,N_24310);
nand UO_850 (O_850,N_24796,N_24473);
nand UO_851 (O_851,N_24412,N_24845);
xnor UO_852 (O_852,N_24628,N_23952);
or UO_853 (O_853,N_24464,N_24051);
or UO_854 (O_854,N_24791,N_23807);
and UO_855 (O_855,N_24536,N_24149);
xnor UO_856 (O_856,N_24397,N_24491);
nand UO_857 (O_857,N_23969,N_24136);
and UO_858 (O_858,N_23752,N_24251);
nor UO_859 (O_859,N_24030,N_23923);
nor UO_860 (O_860,N_23759,N_23815);
and UO_861 (O_861,N_23930,N_23752);
nand UO_862 (O_862,N_24110,N_23812);
nand UO_863 (O_863,N_24572,N_24977);
xnor UO_864 (O_864,N_24995,N_24740);
nand UO_865 (O_865,N_24606,N_24703);
nor UO_866 (O_866,N_24566,N_24230);
and UO_867 (O_867,N_24551,N_24373);
and UO_868 (O_868,N_24353,N_24701);
or UO_869 (O_869,N_24253,N_23907);
or UO_870 (O_870,N_24469,N_24071);
nand UO_871 (O_871,N_24164,N_24460);
nand UO_872 (O_872,N_24000,N_24074);
nand UO_873 (O_873,N_24779,N_24831);
xor UO_874 (O_874,N_24220,N_23782);
nor UO_875 (O_875,N_24476,N_24567);
nand UO_876 (O_876,N_24346,N_24675);
or UO_877 (O_877,N_24966,N_24694);
nand UO_878 (O_878,N_23870,N_24592);
nand UO_879 (O_879,N_24291,N_24139);
xnor UO_880 (O_880,N_23801,N_24189);
nand UO_881 (O_881,N_24988,N_24827);
nand UO_882 (O_882,N_24575,N_24060);
nor UO_883 (O_883,N_24862,N_23982);
nand UO_884 (O_884,N_24453,N_24602);
or UO_885 (O_885,N_24958,N_24536);
xnor UO_886 (O_886,N_24552,N_24101);
xnor UO_887 (O_887,N_23770,N_24678);
xor UO_888 (O_888,N_24518,N_24970);
nor UO_889 (O_889,N_23948,N_24678);
or UO_890 (O_890,N_24971,N_24203);
nor UO_891 (O_891,N_24344,N_23962);
nand UO_892 (O_892,N_24079,N_24048);
and UO_893 (O_893,N_24698,N_23913);
nor UO_894 (O_894,N_23909,N_24576);
or UO_895 (O_895,N_24011,N_24477);
xnor UO_896 (O_896,N_23864,N_24723);
or UO_897 (O_897,N_24101,N_24732);
or UO_898 (O_898,N_24847,N_24267);
nor UO_899 (O_899,N_24732,N_23773);
nand UO_900 (O_900,N_23758,N_24351);
and UO_901 (O_901,N_23927,N_23921);
nand UO_902 (O_902,N_24274,N_24977);
or UO_903 (O_903,N_24329,N_24407);
nand UO_904 (O_904,N_24429,N_24824);
and UO_905 (O_905,N_24083,N_23924);
nand UO_906 (O_906,N_23958,N_24857);
and UO_907 (O_907,N_24278,N_24656);
xor UO_908 (O_908,N_24016,N_24285);
xor UO_909 (O_909,N_24653,N_24803);
and UO_910 (O_910,N_24250,N_23986);
nor UO_911 (O_911,N_24304,N_24198);
nor UO_912 (O_912,N_24524,N_24996);
xnor UO_913 (O_913,N_23898,N_24487);
nor UO_914 (O_914,N_24116,N_23904);
xnor UO_915 (O_915,N_23961,N_23969);
xnor UO_916 (O_916,N_24311,N_23963);
nand UO_917 (O_917,N_24101,N_23769);
and UO_918 (O_918,N_24239,N_24418);
nand UO_919 (O_919,N_24938,N_24245);
or UO_920 (O_920,N_24010,N_23767);
and UO_921 (O_921,N_24159,N_24505);
nor UO_922 (O_922,N_23864,N_24097);
xor UO_923 (O_923,N_24637,N_23978);
or UO_924 (O_924,N_23865,N_23776);
nor UO_925 (O_925,N_24729,N_23866);
or UO_926 (O_926,N_24240,N_24330);
or UO_927 (O_927,N_24780,N_24517);
and UO_928 (O_928,N_24624,N_23796);
nor UO_929 (O_929,N_24230,N_24358);
nor UO_930 (O_930,N_24894,N_23996);
and UO_931 (O_931,N_24695,N_24200);
or UO_932 (O_932,N_24189,N_24641);
nand UO_933 (O_933,N_24420,N_24948);
xnor UO_934 (O_934,N_24708,N_24367);
xnor UO_935 (O_935,N_23951,N_24029);
xor UO_936 (O_936,N_24042,N_24989);
or UO_937 (O_937,N_24956,N_24473);
and UO_938 (O_938,N_24218,N_24852);
or UO_939 (O_939,N_24152,N_24852);
and UO_940 (O_940,N_24066,N_24696);
nor UO_941 (O_941,N_24438,N_23946);
nor UO_942 (O_942,N_24704,N_24268);
or UO_943 (O_943,N_24343,N_23771);
nor UO_944 (O_944,N_24633,N_24495);
nor UO_945 (O_945,N_24886,N_24057);
and UO_946 (O_946,N_24070,N_24378);
or UO_947 (O_947,N_24867,N_24312);
nor UO_948 (O_948,N_24170,N_24188);
and UO_949 (O_949,N_24078,N_24195);
or UO_950 (O_950,N_24955,N_24760);
xnor UO_951 (O_951,N_24709,N_24447);
nor UO_952 (O_952,N_24217,N_24370);
nor UO_953 (O_953,N_23763,N_24260);
xor UO_954 (O_954,N_24187,N_24922);
nand UO_955 (O_955,N_24354,N_24608);
or UO_956 (O_956,N_23782,N_24160);
nor UO_957 (O_957,N_24524,N_24330);
nand UO_958 (O_958,N_24924,N_24186);
nor UO_959 (O_959,N_24835,N_23957);
and UO_960 (O_960,N_24082,N_23897);
and UO_961 (O_961,N_24449,N_23911);
xnor UO_962 (O_962,N_24610,N_24790);
nor UO_963 (O_963,N_24239,N_24957);
nor UO_964 (O_964,N_24390,N_24651);
or UO_965 (O_965,N_23769,N_24677);
or UO_966 (O_966,N_24906,N_24640);
nor UO_967 (O_967,N_24846,N_24295);
or UO_968 (O_968,N_24772,N_23783);
nor UO_969 (O_969,N_24809,N_24149);
nor UO_970 (O_970,N_24426,N_24411);
and UO_971 (O_971,N_24057,N_24175);
or UO_972 (O_972,N_24905,N_24568);
and UO_973 (O_973,N_23862,N_23963);
xnor UO_974 (O_974,N_23938,N_24462);
nand UO_975 (O_975,N_23970,N_23793);
nor UO_976 (O_976,N_24542,N_24656);
nand UO_977 (O_977,N_24509,N_24346);
or UO_978 (O_978,N_23869,N_24074);
or UO_979 (O_979,N_24930,N_24733);
nor UO_980 (O_980,N_24954,N_24864);
nor UO_981 (O_981,N_24666,N_24980);
xnor UO_982 (O_982,N_24694,N_24108);
nor UO_983 (O_983,N_24648,N_24007);
nand UO_984 (O_984,N_24199,N_23808);
nor UO_985 (O_985,N_24752,N_23969);
nor UO_986 (O_986,N_24291,N_23948);
nand UO_987 (O_987,N_24362,N_24196);
nand UO_988 (O_988,N_24448,N_24597);
and UO_989 (O_989,N_24284,N_24235);
nor UO_990 (O_990,N_24846,N_23839);
nand UO_991 (O_991,N_24513,N_23828);
or UO_992 (O_992,N_24399,N_24120);
or UO_993 (O_993,N_24962,N_24323);
or UO_994 (O_994,N_24023,N_24695);
nand UO_995 (O_995,N_24952,N_24335);
xnor UO_996 (O_996,N_24304,N_24210);
xor UO_997 (O_997,N_23891,N_24258);
nand UO_998 (O_998,N_24850,N_24397);
and UO_999 (O_999,N_24614,N_24692);
xor UO_1000 (O_1000,N_24656,N_24001);
and UO_1001 (O_1001,N_24937,N_24940);
or UO_1002 (O_1002,N_24534,N_24940);
xor UO_1003 (O_1003,N_24720,N_24199);
and UO_1004 (O_1004,N_24179,N_23758);
nand UO_1005 (O_1005,N_24738,N_24674);
and UO_1006 (O_1006,N_24674,N_24158);
nor UO_1007 (O_1007,N_24546,N_24807);
xnor UO_1008 (O_1008,N_23837,N_23866);
or UO_1009 (O_1009,N_24539,N_24481);
or UO_1010 (O_1010,N_24420,N_24951);
nand UO_1011 (O_1011,N_24678,N_23780);
and UO_1012 (O_1012,N_24562,N_23823);
nor UO_1013 (O_1013,N_24683,N_24084);
xor UO_1014 (O_1014,N_24164,N_24527);
or UO_1015 (O_1015,N_24574,N_23829);
nand UO_1016 (O_1016,N_24090,N_23886);
xor UO_1017 (O_1017,N_23984,N_24535);
nand UO_1018 (O_1018,N_24878,N_24656);
xor UO_1019 (O_1019,N_24537,N_24199);
nor UO_1020 (O_1020,N_24737,N_24291);
or UO_1021 (O_1021,N_24087,N_23873);
xor UO_1022 (O_1022,N_24923,N_24841);
and UO_1023 (O_1023,N_23760,N_24138);
nand UO_1024 (O_1024,N_24131,N_24100);
xor UO_1025 (O_1025,N_24369,N_23881);
and UO_1026 (O_1026,N_24016,N_24592);
and UO_1027 (O_1027,N_24316,N_24509);
and UO_1028 (O_1028,N_24561,N_24933);
and UO_1029 (O_1029,N_24733,N_24271);
or UO_1030 (O_1030,N_24430,N_24858);
and UO_1031 (O_1031,N_24598,N_24388);
nor UO_1032 (O_1032,N_23985,N_24708);
nand UO_1033 (O_1033,N_23776,N_24213);
nor UO_1034 (O_1034,N_24140,N_24357);
or UO_1035 (O_1035,N_23780,N_24584);
and UO_1036 (O_1036,N_24139,N_24069);
or UO_1037 (O_1037,N_24527,N_23766);
nand UO_1038 (O_1038,N_24123,N_24442);
or UO_1039 (O_1039,N_24855,N_24212);
xor UO_1040 (O_1040,N_24171,N_24922);
nand UO_1041 (O_1041,N_24684,N_24682);
nor UO_1042 (O_1042,N_24334,N_24802);
and UO_1043 (O_1043,N_23904,N_24718);
and UO_1044 (O_1044,N_23922,N_24567);
and UO_1045 (O_1045,N_24081,N_24198);
nor UO_1046 (O_1046,N_24751,N_24727);
or UO_1047 (O_1047,N_24079,N_24939);
nor UO_1048 (O_1048,N_24491,N_24852);
xnor UO_1049 (O_1049,N_23763,N_24076);
or UO_1050 (O_1050,N_24519,N_24630);
or UO_1051 (O_1051,N_24546,N_23856);
nand UO_1052 (O_1052,N_24063,N_23921);
and UO_1053 (O_1053,N_24047,N_23924);
xor UO_1054 (O_1054,N_24558,N_24615);
xnor UO_1055 (O_1055,N_24946,N_24572);
xor UO_1056 (O_1056,N_24314,N_24320);
nor UO_1057 (O_1057,N_24677,N_23989);
nand UO_1058 (O_1058,N_24050,N_24761);
nor UO_1059 (O_1059,N_24281,N_24484);
and UO_1060 (O_1060,N_24064,N_24632);
xor UO_1061 (O_1061,N_23768,N_24936);
nor UO_1062 (O_1062,N_24750,N_23893);
nor UO_1063 (O_1063,N_24683,N_24923);
nand UO_1064 (O_1064,N_23999,N_24567);
nor UO_1065 (O_1065,N_24367,N_24721);
nor UO_1066 (O_1066,N_24478,N_23989);
nor UO_1067 (O_1067,N_24200,N_24920);
or UO_1068 (O_1068,N_24963,N_23967);
nand UO_1069 (O_1069,N_23960,N_24566);
nor UO_1070 (O_1070,N_23791,N_24696);
xnor UO_1071 (O_1071,N_24531,N_24161);
or UO_1072 (O_1072,N_24076,N_24160);
and UO_1073 (O_1073,N_24936,N_24938);
nand UO_1074 (O_1074,N_24026,N_24880);
or UO_1075 (O_1075,N_23831,N_24063);
xor UO_1076 (O_1076,N_24579,N_24804);
nor UO_1077 (O_1077,N_24326,N_24532);
nand UO_1078 (O_1078,N_24129,N_24966);
nor UO_1079 (O_1079,N_24058,N_24264);
or UO_1080 (O_1080,N_24016,N_24169);
nand UO_1081 (O_1081,N_24768,N_24669);
xnor UO_1082 (O_1082,N_24079,N_24056);
xor UO_1083 (O_1083,N_24466,N_23788);
nor UO_1084 (O_1084,N_24575,N_24902);
xor UO_1085 (O_1085,N_24957,N_23901);
and UO_1086 (O_1086,N_24097,N_24183);
nor UO_1087 (O_1087,N_24226,N_24560);
and UO_1088 (O_1088,N_24415,N_24491);
or UO_1089 (O_1089,N_24296,N_23955);
and UO_1090 (O_1090,N_24542,N_24072);
and UO_1091 (O_1091,N_23759,N_24869);
nand UO_1092 (O_1092,N_24658,N_24717);
xnor UO_1093 (O_1093,N_24868,N_24258);
nand UO_1094 (O_1094,N_24030,N_24575);
xnor UO_1095 (O_1095,N_24861,N_24531);
nand UO_1096 (O_1096,N_23893,N_23948);
nor UO_1097 (O_1097,N_24474,N_24206);
or UO_1098 (O_1098,N_24759,N_23795);
nand UO_1099 (O_1099,N_23833,N_24053);
nand UO_1100 (O_1100,N_23862,N_24494);
nor UO_1101 (O_1101,N_24898,N_24313);
or UO_1102 (O_1102,N_23806,N_24793);
or UO_1103 (O_1103,N_24882,N_23815);
and UO_1104 (O_1104,N_24923,N_23803);
and UO_1105 (O_1105,N_24832,N_24393);
xnor UO_1106 (O_1106,N_24959,N_24442);
nor UO_1107 (O_1107,N_24947,N_24178);
nor UO_1108 (O_1108,N_24815,N_24058);
nand UO_1109 (O_1109,N_23999,N_24417);
nor UO_1110 (O_1110,N_24241,N_24194);
nor UO_1111 (O_1111,N_24840,N_23969);
or UO_1112 (O_1112,N_23853,N_23981);
xor UO_1113 (O_1113,N_24941,N_24524);
and UO_1114 (O_1114,N_24766,N_24608);
nand UO_1115 (O_1115,N_24985,N_24752);
xor UO_1116 (O_1116,N_24285,N_23853);
or UO_1117 (O_1117,N_24975,N_24653);
and UO_1118 (O_1118,N_24093,N_24394);
and UO_1119 (O_1119,N_24621,N_23780);
nor UO_1120 (O_1120,N_24069,N_24550);
or UO_1121 (O_1121,N_23855,N_24111);
or UO_1122 (O_1122,N_24054,N_24784);
or UO_1123 (O_1123,N_24758,N_24505);
nor UO_1124 (O_1124,N_24441,N_24730);
nor UO_1125 (O_1125,N_23827,N_24653);
and UO_1126 (O_1126,N_23896,N_23775);
nand UO_1127 (O_1127,N_24692,N_24569);
and UO_1128 (O_1128,N_24711,N_24798);
xor UO_1129 (O_1129,N_24374,N_24491);
xor UO_1130 (O_1130,N_24461,N_23822);
and UO_1131 (O_1131,N_24785,N_24015);
nand UO_1132 (O_1132,N_23969,N_24503);
xnor UO_1133 (O_1133,N_23816,N_23953);
and UO_1134 (O_1134,N_24213,N_23946);
xor UO_1135 (O_1135,N_24505,N_24176);
and UO_1136 (O_1136,N_24366,N_23869);
nor UO_1137 (O_1137,N_24609,N_24993);
and UO_1138 (O_1138,N_23859,N_24024);
and UO_1139 (O_1139,N_24650,N_24585);
nor UO_1140 (O_1140,N_24861,N_24512);
nand UO_1141 (O_1141,N_24324,N_24889);
nand UO_1142 (O_1142,N_24138,N_24427);
xnor UO_1143 (O_1143,N_24682,N_23864);
or UO_1144 (O_1144,N_24578,N_24354);
nor UO_1145 (O_1145,N_24946,N_24419);
or UO_1146 (O_1146,N_24533,N_24273);
xor UO_1147 (O_1147,N_23800,N_24898);
nor UO_1148 (O_1148,N_24073,N_24326);
and UO_1149 (O_1149,N_24703,N_23911);
nand UO_1150 (O_1150,N_24011,N_24840);
nand UO_1151 (O_1151,N_23771,N_24695);
nor UO_1152 (O_1152,N_23887,N_24864);
and UO_1153 (O_1153,N_24788,N_23991);
and UO_1154 (O_1154,N_24631,N_24821);
and UO_1155 (O_1155,N_23971,N_23786);
or UO_1156 (O_1156,N_24725,N_24705);
xnor UO_1157 (O_1157,N_23819,N_24356);
and UO_1158 (O_1158,N_24328,N_23936);
xor UO_1159 (O_1159,N_24686,N_24313);
nand UO_1160 (O_1160,N_24543,N_24941);
and UO_1161 (O_1161,N_24969,N_24203);
nor UO_1162 (O_1162,N_24276,N_24308);
nand UO_1163 (O_1163,N_24876,N_24769);
nor UO_1164 (O_1164,N_24213,N_24925);
and UO_1165 (O_1165,N_24429,N_24129);
or UO_1166 (O_1166,N_24048,N_24095);
nor UO_1167 (O_1167,N_23864,N_24734);
and UO_1168 (O_1168,N_24557,N_24239);
and UO_1169 (O_1169,N_24513,N_23924);
or UO_1170 (O_1170,N_24913,N_24853);
and UO_1171 (O_1171,N_24578,N_23891);
nor UO_1172 (O_1172,N_24478,N_24491);
or UO_1173 (O_1173,N_23753,N_24511);
nor UO_1174 (O_1174,N_24313,N_24671);
or UO_1175 (O_1175,N_23816,N_24425);
xnor UO_1176 (O_1176,N_24900,N_23862);
xor UO_1177 (O_1177,N_24970,N_24011);
nand UO_1178 (O_1178,N_24535,N_24082);
or UO_1179 (O_1179,N_24444,N_24795);
nor UO_1180 (O_1180,N_23943,N_24777);
and UO_1181 (O_1181,N_23784,N_24184);
and UO_1182 (O_1182,N_24142,N_24351);
and UO_1183 (O_1183,N_24815,N_24297);
and UO_1184 (O_1184,N_24421,N_23763);
nor UO_1185 (O_1185,N_24848,N_23867);
or UO_1186 (O_1186,N_24698,N_24001);
nor UO_1187 (O_1187,N_24738,N_24287);
or UO_1188 (O_1188,N_24828,N_24751);
and UO_1189 (O_1189,N_24679,N_24104);
nor UO_1190 (O_1190,N_24939,N_24390);
nand UO_1191 (O_1191,N_24943,N_24181);
nand UO_1192 (O_1192,N_24111,N_24265);
and UO_1193 (O_1193,N_24398,N_24209);
xor UO_1194 (O_1194,N_23868,N_24033);
nor UO_1195 (O_1195,N_24185,N_24026);
or UO_1196 (O_1196,N_24521,N_24400);
xor UO_1197 (O_1197,N_23884,N_24133);
xor UO_1198 (O_1198,N_24905,N_24355);
nand UO_1199 (O_1199,N_24706,N_24523);
or UO_1200 (O_1200,N_24505,N_24247);
nand UO_1201 (O_1201,N_24424,N_24446);
nor UO_1202 (O_1202,N_23962,N_23782);
and UO_1203 (O_1203,N_23778,N_23849);
nand UO_1204 (O_1204,N_23786,N_24362);
nor UO_1205 (O_1205,N_24822,N_23922);
xor UO_1206 (O_1206,N_23753,N_24433);
xnor UO_1207 (O_1207,N_24998,N_24230);
and UO_1208 (O_1208,N_24038,N_24865);
xor UO_1209 (O_1209,N_24218,N_23833);
xor UO_1210 (O_1210,N_24106,N_24772);
nor UO_1211 (O_1211,N_24152,N_24781);
or UO_1212 (O_1212,N_24842,N_24447);
and UO_1213 (O_1213,N_24938,N_24990);
or UO_1214 (O_1214,N_23884,N_24871);
or UO_1215 (O_1215,N_23935,N_24554);
and UO_1216 (O_1216,N_23769,N_24256);
nor UO_1217 (O_1217,N_24149,N_23972);
nor UO_1218 (O_1218,N_24050,N_23781);
xnor UO_1219 (O_1219,N_24178,N_24549);
xor UO_1220 (O_1220,N_24026,N_24051);
nor UO_1221 (O_1221,N_24289,N_24213);
xnor UO_1222 (O_1222,N_24571,N_24999);
xnor UO_1223 (O_1223,N_23830,N_23849);
nand UO_1224 (O_1224,N_24642,N_24358);
nand UO_1225 (O_1225,N_24118,N_24726);
nand UO_1226 (O_1226,N_23791,N_24359);
nand UO_1227 (O_1227,N_24833,N_24280);
and UO_1228 (O_1228,N_24268,N_24255);
or UO_1229 (O_1229,N_23925,N_24574);
or UO_1230 (O_1230,N_23925,N_24493);
and UO_1231 (O_1231,N_24879,N_24621);
xnor UO_1232 (O_1232,N_24999,N_23781);
nand UO_1233 (O_1233,N_23797,N_24390);
and UO_1234 (O_1234,N_24200,N_23831);
xnor UO_1235 (O_1235,N_24901,N_24894);
nor UO_1236 (O_1236,N_24907,N_24845);
xor UO_1237 (O_1237,N_24115,N_24366);
xor UO_1238 (O_1238,N_24727,N_24281);
nor UO_1239 (O_1239,N_23804,N_24531);
and UO_1240 (O_1240,N_23830,N_24667);
and UO_1241 (O_1241,N_24231,N_23835);
nor UO_1242 (O_1242,N_24660,N_23926);
and UO_1243 (O_1243,N_23994,N_23867);
nor UO_1244 (O_1244,N_24110,N_23834);
xor UO_1245 (O_1245,N_24054,N_24540);
nand UO_1246 (O_1246,N_24549,N_24719);
xnor UO_1247 (O_1247,N_24817,N_24192);
and UO_1248 (O_1248,N_24107,N_23836);
or UO_1249 (O_1249,N_23948,N_24479);
nor UO_1250 (O_1250,N_24304,N_24034);
nand UO_1251 (O_1251,N_23776,N_24628);
nand UO_1252 (O_1252,N_24316,N_24908);
xor UO_1253 (O_1253,N_24405,N_24643);
and UO_1254 (O_1254,N_24115,N_23847);
and UO_1255 (O_1255,N_24266,N_24546);
xor UO_1256 (O_1256,N_24224,N_24698);
nor UO_1257 (O_1257,N_24047,N_24344);
xnor UO_1258 (O_1258,N_23812,N_23884);
nor UO_1259 (O_1259,N_24235,N_24815);
nor UO_1260 (O_1260,N_24146,N_24141);
xnor UO_1261 (O_1261,N_24528,N_24727);
or UO_1262 (O_1262,N_24288,N_24033);
xor UO_1263 (O_1263,N_24446,N_24311);
xnor UO_1264 (O_1264,N_23799,N_23911);
nand UO_1265 (O_1265,N_23866,N_24925);
nor UO_1266 (O_1266,N_23881,N_24842);
xnor UO_1267 (O_1267,N_24668,N_24592);
or UO_1268 (O_1268,N_24397,N_23883);
and UO_1269 (O_1269,N_24011,N_24951);
nand UO_1270 (O_1270,N_24150,N_24215);
nor UO_1271 (O_1271,N_24689,N_24666);
xnor UO_1272 (O_1272,N_24543,N_23809);
nand UO_1273 (O_1273,N_24253,N_24315);
nand UO_1274 (O_1274,N_24279,N_24051);
nor UO_1275 (O_1275,N_24630,N_23806);
nand UO_1276 (O_1276,N_24792,N_24162);
or UO_1277 (O_1277,N_24826,N_24188);
nor UO_1278 (O_1278,N_24703,N_24702);
nand UO_1279 (O_1279,N_24139,N_24470);
and UO_1280 (O_1280,N_23895,N_24777);
and UO_1281 (O_1281,N_24699,N_23988);
nand UO_1282 (O_1282,N_24008,N_24600);
xor UO_1283 (O_1283,N_24643,N_24947);
xor UO_1284 (O_1284,N_23892,N_24312);
xor UO_1285 (O_1285,N_24877,N_24627);
nor UO_1286 (O_1286,N_24882,N_24908);
nor UO_1287 (O_1287,N_24192,N_24783);
xnor UO_1288 (O_1288,N_23814,N_24458);
nor UO_1289 (O_1289,N_24565,N_24753);
nand UO_1290 (O_1290,N_24464,N_24888);
and UO_1291 (O_1291,N_24128,N_24254);
and UO_1292 (O_1292,N_24745,N_24165);
xor UO_1293 (O_1293,N_24981,N_24743);
xor UO_1294 (O_1294,N_23880,N_24676);
and UO_1295 (O_1295,N_24869,N_24410);
xor UO_1296 (O_1296,N_24289,N_23752);
nand UO_1297 (O_1297,N_23783,N_23955);
xor UO_1298 (O_1298,N_24167,N_24329);
nand UO_1299 (O_1299,N_24170,N_23801);
or UO_1300 (O_1300,N_24291,N_24644);
and UO_1301 (O_1301,N_23804,N_24494);
and UO_1302 (O_1302,N_24042,N_24235);
nand UO_1303 (O_1303,N_24327,N_24783);
and UO_1304 (O_1304,N_24388,N_24188);
and UO_1305 (O_1305,N_24227,N_24895);
nand UO_1306 (O_1306,N_23776,N_24554);
xor UO_1307 (O_1307,N_23750,N_23812);
and UO_1308 (O_1308,N_24300,N_24568);
and UO_1309 (O_1309,N_24967,N_24858);
or UO_1310 (O_1310,N_24018,N_24232);
or UO_1311 (O_1311,N_23996,N_24118);
or UO_1312 (O_1312,N_24980,N_24041);
or UO_1313 (O_1313,N_24794,N_24090);
nor UO_1314 (O_1314,N_24404,N_24471);
nor UO_1315 (O_1315,N_24938,N_23923);
nor UO_1316 (O_1316,N_23914,N_24148);
or UO_1317 (O_1317,N_24616,N_23787);
xor UO_1318 (O_1318,N_23876,N_23793);
nor UO_1319 (O_1319,N_24131,N_24515);
nor UO_1320 (O_1320,N_24291,N_24433);
nor UO_1321 (O_1321,N_24146,N_24776);
and UO_1322 (O_1322,N_24158,N_24825);
nand UO_1323 (O_1323,N_23801,N_24791);
and UO_1324 (O_1324,N_24775,N_23974);
or UO_1325 (O_1325,N_24777,N_24724);
and UO_1326 (O_1326,N_24515,N_24928);
and UO_1327 (O_1327,N_24645,N_24817);
nor UO_1328 (O_1328,N_24525,N_24417);
nand UO_1329 (O_1329,N_24443,N_24669);
and UO_1330 (O_1330,N_23764,N_23957);
nand UO_1331 (O_1331,N_24315,N_24768);
nor UO_1332 (O_1332,N_24845,N_23772);
nand UO_1333 (O_1333,N_24962,N_24723);
nor UO_1334 (O_1334,N_24363,N_24989);
nor UO_1335 (O_1335,N_24488,N_24346);
xor UO_1336 (O_1336,N_23775,N_23995);
or UO_1337 (O_1337,N_24786,N_24939);
or UO_1338 (O_1338,N_24294,N_24835);
or UO_1339 (O_1339,N_23858,N_23814);
and UO_1340 (O_1340,N_24151,N_24477);
nor UO_1341 (O_1341,N_24419,N_24766);
nand UO_1342 (O_1342,N_24475,N_24782);
nor UO_1343 (O_1343,N_23810,N_24944);
or UO_1344 (O_1344,N_24945,N_24379);
nand UO_1345 (O_1345,N_23810,N_24446);
or UO_1346 (O_1346,N_24617,N_24093);
nor UO_1347 (O_1347,N_24629,N_24862);
and UO_1348 (O_1348,N_24563,N_24119);
and UO_1349 (O_1349,N_24136,N_24190);
nand UO_1350 (O_1350,N_23844,N_23752);
nor UO_1351 (O_1351,N_24510,N_24723);
xor UO_1352 (O_1352,N_24100,N_24237);
nor UO_1353 (O_1353,N_24225,N_24012);
or UO_1354 (O_1354,N_24743,N_23791);
and UO_1355 (O_1355,N_24917,N_23829);
xnor UO_1356 (O_1356,N_24073,N_24085);
or UO_1357 (O_1357,N_24376,N_24482);
and UO_1358 (O_1358,N_24932,N_23764);
and UO_1359 (O_1359,N_24065,N_24043);
xor UO_1360 (O_1360,N_24207,N_24697);
and UO_1361 (O_1361,N_24623,N_24794);
or UO_1362 (O_1362,N_24349,N_24115);
nand UO_1363 (O_1363,N_24515,N_24624);
and UO_1364 (O_1364,N_23798,N_24375);
nand UO_1365 (O_1365,N_24340,N_24107);
or UO_1366 (O_1366,N_23787,N_24726);
nand UO_1367 (O_1367,N_24153,N_24171);
or UO_1368 (O_1368,N_24803,N_24819);
nand UO_1369 (O_1369,N_24158,N_24840);
or UO_1370 (O_1370,N_24948,N_24668);
or UO_1371 (O_1371,N_24982,N_24549);
or UO_1372 (O_1372,N_24212,N_23982);
nand UO_1373 (O_1373,N_24641,N_24466);
nor UO_1374 (O_1374,N_24974,N_24805);
nor UO_1375 (O_1375,N_23947,N_24845);
or UO_1376 (O_1376,N_24515,N_24334);
and UO_1377 (O_1377,N_24872,N_23750);
or UO_1378 (O_1378,N_24390,N_24731);
nor UO_1379 (O_1379,N_24282,N_24898);
and UO_1380 (O_1380,N_24863,N_23932);
or UO_1381 (O_1381,N_24770,N_24548);
and UO_1382 (O_1382,N_24386,N_24492);
xor UO_1383 (O_1383,N_24951,N_23927);
or UO_1384 (O_1384,N_24463,N_23821);
and UO_1385 (O_1385,N_24499,N_24532);
nor UO_1386 (O_1386,N_23762,N_24140);
and UO_1387 (O_1387,N_24294,N_24680);
nand UO_1388 (O_1388,N_24347,N_24674);
and UO_1389 (O_1389,N_24848,N_24491);
nand UO_1390 (O_1390,N_24342,N_24098);
xor UO_1391 (O_1391,N_24024,N_23806);
nor UO_1392 (O_1392,N_24231,N_24036);
xor UO_1393 (O_1393,N_24010,N_23870);
or UO_1394 (O_1394,N_24746,N_24886);
xor UO_1395 (O_1395,N_24908,N_24562);
nand UO_1396 (O_1396,N_24786,N_24468);
or UO_1397 (O_1397,N_24376,N_24398);
or UO_1398 (O_1398,N_23968,N_24442);
nor UO_1399 (O_1399,N_24104,N_23918);
nand UO_1400 (O_1400,N_23824,N_24642);
nand UO_1401 (O_1401,N_24915,N_23994);
and UO_1402 (O_1402,N_24538,N_24861);
nor UO_1403 (O_1403,N_24397,N_24583);
and UO_1404 (O_1404,N_24219,N_24474);
or UO_1405 (O_1405,N_24383,N_24466);
xor UO_1406 (O_1406,N_24147,N_24750);
and UO_1407 (O_1407,N_24310,N_24505);
and UO_1408 (O_1408,N_24815,N_24502);
nor UO_1409 (O_1409,N_24674,N_24202);
and UO_1410 (O_1410,N_23783,N_24721);
nand UO_1411 (O_1411,N_23907,N_24296);
or UO_1412 (O_1412,N_24830,N_24885);
or UO_1413 (O_1413,N_24603,N_24068);
nor UO_1414 (O_1414,N_24983,N_24404);
xor UO_1415 (O_1415,N_23862,N_23861);
nand UO_1416 (O_1416,N_24675,N_24320);
or UO_1417 (O_1417,N_24164,N_24571);
xnor UO_1418 (O_1418,N_24266,N_24570);
xor UO_1419 (O_1419,N_24249,N_24161);
xor UO_1420 (O_1420,N_24815,N_23785);
and UO_1421 (O_1421,N_24354,N_24270);
or UO_1422 (O_1422,N_24663,N_24637);
xnor UO_1423 (O_1423,N_24367,N_23972);
and UO_1424 (O_1424,N_24680,N_24613);
nor UO_1425 (O_1425,N_23798,N_24791);
nand UO_1426 (O_1426,N_24727,N_24289);
and UO_1427 (O_1427,N_24024,N_24292);
or UO_1428 (O_1428,N_24442,N_24742);
or UO_1429 (O_1429,N_23921,N_24180);
nor UO_1430 (O_1430,N_24208,N_24924);
nor UO_1431 (O_1431,N_24386,N_24950);
xnor UO_1432 (O_1432,N_24321,N_24937);
and UO_1433 (O_1433,N_24724,N_24137);
nand UO_1434 (O_1434,N_23974,N_24321);
xor UO_1435 (O_1435,N_23870,N_23920);
or UO_1436 (O_1436,N_24482,N_24145);
and UO_1437 (O_1437,N_24435,N_23934);
or UO_1438 (O_1438,N_24500,N_24762);
and UO_1439 (O_1439,N_23760,N_24419);
and UO_1440 (O_1440,N_24591,N_23977);
and UO_1441 (O_1441,N_24292,N_23988);
nand UO_1442 (O_1442,N_24615,N_24546);
nand UO_1443 (O_1443,N_24261,N_24248);
nand UO_1444 (O_1444,N_24488,N_23854);
nor UO_1445 (O_1445,N_23828,N_23999);
or UO_1446 (O_1446,N_24269,N_24660);
or UO_1447 (O_1447,N_24424,N_24012);
nand UO_1448 (O_1448,N_23998,N_24093);
xnor UO_1449 (O_1449,N_24281,N_23883);
nand UO_1450 (O_1450,N_24697,N_24316);
nand UO_1451 (O_1451,N_24877,N_24801);
or UO_1452 (O_1452,N_23975,N_23753);
xnor UO_1453 (O_1453,N_24659,N_24653);
and UO_1454 (O_1454,N_23846,N_24917);
or UO_1455 (O_1455,N_24454,N_23926);
nand UO_1456 (O_1456,N_24148,N_24489);
nand UO_1457 (O_1457,N_24565,N_24163);
or UO_1458 (O_1458,N_24359,N_24973);
or UO_1459 (O_1459,N_24139,N_24087);
and UO_1460 (O_1460,N_24127,N_24534);
xnor UO_1461 (O_1461,N_24775,N_24660);
and UO_1462 (O_1462,N_23802,N_24538);
nor UO_1463 (O_1463,N_23924,N_23943);
nor UO_1464 (O_1464,N_24122,N_24133);
or UO_1465 (O_1465,N_24777,N_24300);
or UO_1466 (O_1466,N_24461,N_23783);
nor UO_1467 (O_1467,N_24749,N_24982);
or UO_1468 (O_1468,N_23893,N_24715);
or UO_1469 (O_1469,N_24284,N_23987);
and UO_1470 (O_1470,N_24525,N_24219);
or UO_1471 (O_1471,N_24518,N_24533);
and UO_1472 (O_1472,N_24909,N_24895);
nor UO_1473 (O_1473,N_24379,N_24417);
and UO_1474 (O_1474,N_24864,N_24313);
nand UO_1475 (O_1475,N_23830,N_23779);
nor UO_1476 (O_1476,N_24900,N_24410);
nor UO_1477 (O_1477,N_24896,N_24598);
or UO_1478 (O_1478,N_24476,N_24223);
or UO_1479 (O_1479,N_24847,N_24029);
nor UO_1480 (O_1480,N_24661,N_23813);
and UO_1481 (O_1481,N_23813,N_23818);
xnor UO_1482 (O_1482,N_24798,N_24113);
and UO_1483 (O_1483,N_23931,N_24588);
or UO_1484 (O_1484,N_24955,N_24376);
and UO_1485 (O_1485,N_24290,N_24255);
xnor UO_1486 (O_1486,N_24120,N_24488);
xor UO_1487 (O_1487,N_24743,N_24372);
nand UO_1488 (O_1488,N_23914,N_24960);
nor UO_1489 (O_1489,N_24542,N_24644);
or UO_1490 (O_1490,N_24223,N_24725);
and UO_1491 (O_1491,N_23764,N_23904);
or UO_1492 (O_1492,N_24827,N_24459);
nand UO_1493 (O_1493,N_23905,N_24707);
xor UO_1494 (O_1494,N_24525,N_24725);
or UO_1495 (O_1495,N_24883,N_24323);
and UO_1496 (O_1496,N_24151,N_24989);
and UO_1497 (O_1497,N_23878,N_24552);
nor UO_1498 (O_1498,N_24613,N_23882);
xor UO_1499 (O_1499,N_24707,N_24884);
xnor UO_1500 (O_1500,N_24069,N_24908);
and UO_1501 (O_1501,N_24596,N_24232);
nand UO_1502 (O_1502,N_24632,N_23775);
nor UO_1503 (O_1503,N_24994,N_24989);
xnor UO_1504 (O_1504,N_24506,N_24405);
and UO_1505 (O_1505,N_24496,N_24932);
nor UO_1506 (O_1506,N_24230,N_23987);
nand UO_1507 (O_1507,N_24423,N_23884);
nor UO_1508 (O_1508,N_24572,N_24179);
and UO_1509 (O_1509,N_23902,N_24313);
and UO_1510 (O_1510,N_24132,N_24160);
xnor UO_1511 (O_1511,N_24355,N_24419);
xnor UO_1512 (O_1512,N_23986,N_24355);
or UO_1513 (O_1513,N_24270,N_23971);
nor UO_1514 (O_1514,N_23881,N_24896);
and UO_1515 (O_1515,N_24030,N_24853);
nand UO_1516 (O_1516,N_24561,N_23899);
and UO_1517 (O_1517,N_24817,N_24430);
xnor UO_1518 (O_1518,N_24798,N_24489);
or UO_1519 (O_1519,N_24461,N_24026);
nor UO_1520 (O_1520,N_24185,N_23783);
xor UO_1521 (O_1521,N_23964,N_24335);
xnor UO_1522 (O_1522,N_23796,N_24649);
or UO_1523 (O_1523,N_24842,N_24080);
nor UO_1524 (O_1524,N_23880,N_23852);
xor UO_1525 (O_1525,N_24493,N_24303);
nand UO_1526 (O_1526,N_24234,N_24943);
nand UO_1527 (O_1527,N_24749,N_24493);
xnor UO_1528 (O_1528,N_24072,N_24223);
or UO_1529 (O_1529,N_23767,N_24474);
and UO_1530 (O_1530,N_24199,N_24160);
or UO_1531 (O_1531,N_24785,N_23844);
or UO_1532 (O_1532,N_24562,N_24461);
and UO_1533 (O_1533,N_24668,N_24879);
nand UO_1534 (O_1534,N_24433,N_23943);
or UO_1535 (O_1535,N_24998,N_24707);
nand UO_1536 (O_1536,N_24168,N_24754);
xor UO_1537 (O_1537,N_24432,N_24153);
or UO_1538 (O_1538,N_24322,N_23971);
nor UO_1539 (O_1539,N_23946,N_24176);
nand UO_1540 (O_1540,N_24332,N_24989);
xnor UO_1541 (O_1541,N_24047,N_24760);
nand UO_1542 (O_1542,N_24332,N_24852);
nor UO_1543 (O_1543,N_24087,N_23836);
xnor UO_1544 (O_1544,N_24944,N_24007);
nor UO_1545 (O_1545,N_24859,N_24770);
xor UO_1546 (O_1546,N_24488,N_24594);
or UO_1547 (O_1547,N_24584,N_23883);
and UO_1548 (O_1548,N_24318,N_23773);
xnor UO_1549 (O_1549,N_24908,N_24991);
xor UO_1550 (O_1550,N_24853,N_24706);
xor UO_1551 (O_1551,N_24328,N_24998);
nor UO_1552 (O_1552,N_24410,N_24921);
nor UO_1553 (O_1553,N_24878,N_24802);
xor UO_1554 (O_1554,N_24858,N_24102);
nand UO_1555 (O_1555,N_24700,N_24699);
or UO_1556 (O_1556,N_24988,N_24129);
xnor UO_1557 (O_1557,N_24858,N_24986);
nor UO_1558 (O_1558,N_23986,N_23908);
or UO_1559 (O_1559,N_23876,N_24768);
xor UO_1560 (O_1560,N_23845,N_23905);
or UO_1561 (O_1561,N_24198,N_23928);
and UO_1562 (O_1562,N_24155,N_24278);
or UO_1563 (O_1563,N_24855,N_24410);
xnor UO_1564 (O_1564,N_24785,N_24546);
and UO_1565 (O_1565,N_24567,N_23947);
and UO_1566 (O_1566,N_24594,N_24962);
nand UO_1567 (O_1567,N_24833,N_24583);
nor UO_1568 (O_1568,N_23825,N_24784);
and UO_1569 (O_1569,N_24729,N_24905);
nand UO_1570 (O_1570,N_24864,N_24943);
and UO_1571 (O_1571,N_24962,N_24105);
xor UO_1572 (O_1572,N_24324,N_24931);
nor UO_1573 (O_1573,N_23998,N_24291);
nand UO_1574 (O_1574,N_23870,N_24061);
and UO_1575 (O_1575,N_24147,N_24152);
or UO_1576 (O_1576,N_24958,N_24647);
nor UO_1577 (O_1577,N_24134,N_24416);
nor UO_1578 (O_1578,N_24970,N_24720);
nand UO_1579 (O_1579,N_24972,N_24949);
xnor UO_1580 (O_1580,N_24110,N_24200);
nor UO_1581 (O_1581,N_24758,N_24788);
nand UO_1582 (O_1582,N_24511,N_23791);
nand UO_1583 (O_1583,N_24917,N_24501);
nand UO_1584 (O_1584,N_24479,N_23985);
and UO_1585 (O_1585,N_24305,N_24072);
nand UO_1586 (O_1586,N_24417,N_24729);
nor UO_1587 (O_1587,N_23967,N_23900);
or UO_1588 (O_1588,N_24975,N_24644);
nor UO_1589 (O_1589,N_24865,N_23843);
or UO_1590 (O_1590,N_23979,N_24829);
or UO_1591 (O_1591,N_24803,N_24378);
nor UO_1592 (O_1592,N_24003,N_24684);
and UO_1593 (O_1593,N_24399,N_23958);
nand UO_1594 (O_1594,N_24607,N_24904);
xnor UO_1595 (O_1595,N_23958,N_24102);
nor UO_1596 (O_1596,N_23904,N_24975);
xnor UO_1597 (O_1597,N_24481,N_24430);
and UO_1598 (O_1598,N_24538,N_24617);
nor UO_1599 (O_1599,N_24758,N_24103);
or UO_1600 (O_1600,N_24955,N_24893);
nor UO_1601 (O_1601,N_23902,N_24955);
nor UO_1602 (O_1602,N_23861,N_24308);
nor UO_1603 (O_1603,N_24079,N_24868);
nor UO_1604 (O_1604,N_23994,N_24791);
xor UO_1605 (O_1605,N_23899,N_24881);
and UO_1606 (O_1606,N_24691,N_23959);
nor UO_1607 (O_1607,N_24729,N_24508);
xor UO_1608 (O_1608,N_23842,N_24289);
and UO_1609 (O_1609,N_24426,N_23786);
xnor UO_1610 (O_1610,N_24684,N_24552);
xnor UO_1611 (O_1611,N_23823,N_24308);
xor UO_1612 (O_1612,N_24837,N_24332);
xnor UO_1613 (O_1613,N_24527,N_24939);
or UO_1614 (O_1614,N_23774,N_24649);
nor UO_1615 (O_1615,N_24837,N_24746);
nand UO_1616 (O_1616,N_24829,N_23934);
or UO_1617 (O_1617,N_24773,N_23791);
xor UO_1618 (O_1618,N_24904,N_23873);
or UO_1619 (O_1619,N_24811,N_24937);
nor UO_1620 (O_1620,N_24656,N_24703);
and UO_1621 (O_1621,N_23820,N_24760);
nor UO_1622 (O_1622,N_23863,N_23752);
nand UO_1623 (O_1623,N_24125,N_24763);
and UO_1624 (O_1624,N_24284,N_24086);
or UO_1625 (O_1625,N_24966,N_24533);
xnor UO_1626 (O_1626,N_23763,N_24533);
or UO_1627 (O_1627,N_24302,N_24575);
or UO_1628 (O_1628,N_24857,N_24707);
nor UO_1629 (O_1629,N_24078,N_23815);
nand UO_1630 (O_1630,N_24091,N_24947);
and UO_1631 (O_1631,N_24865,N_23758);
xnor UO_1632 (O_1632,N_24559,N_24656);
or UO_1633 (O_1633,N_23909,N_24572);
or UO_1634 (O_1634,N_23767,N_24028);
xor UO_1635 (O_1635,N_24662,N_23852);
xnor UO_1636 (O_1636,N_24654,N_24336);
and UO_1637 (O_1637,N_23964,N_24826);
nand UO_1638 (O_1638,N_24505,N_24826);
xnor UO_1639 (O_1639,N_24233,N_24280);
xnor UO_1640 (O_1640,N_23974,N_24486);
xnor UO_1641 (O_1641,N_24416,N_24890);
or UO_1642 (O_1642,N_23967,N_23805);
or UO_1643 (O_1643,N_23993,N_23798);
nand UO_1644 (O_1644,N_24386,N_24373);
nand UO_1645 (O_1645,N_24553,N_24520);
xnor UO_1646 (O_1646,N_24812,N_24143);
and UO_1647 (O_1647,N_24682,N_24477);
xnor UO_1648 (O_1648,N_24419,N_23821);
nand UO_1649 (O_1649,N_24522,N_24136);
xor UO_1650 (O_1650,N_24399,N_24795);
nand UO_1651 (O_1651,N_24815,N_24521);
nor UO_1652 (O_1652,N_24832,N_24340);
or UO_1653 (O_1653,N_23819,N_24161);
and UO_1654 (O_1654,N_24902,N_24805);
and UO_1655 (O_1655,N_24468,N_24329);
or UO_1656 (O_1656,N_24286,N_24926);
nand UO_1657 (O_1657,N_24758,N_24267);
xnor UO_1658 (O_1658,N_24748,N_24495);
nor UO_1659 (O_1659,N_24770,N_24289);
and UO_1660 (O_1660,N_24507,N_24813);
xnor UO_1661 (O_1661,N_23813,N_24019);
xnor UO_1662 (O_1662,N_23878,N_23923);
xor UO_1663 (O_1663,N_23775,N_23922);
and UO_1664 (O_1664,N_24857,N_24820);
and UO_1665 (O_1665,N_23919,N_24118);
or UO_1666 (O_1666,N_24261,N_24090);
or UO_1667 (O_1667,N_24049,N_24486);
or UO_1668 (O_1668,N_24873,N_24211);
nand UO_1669 (O_1669,N_24875,N_23800);
nand UO_1670 (O_1670,N_24002,N_24342);
nand UO_1671 (O_1671,N_24040,N_24655);
nand UO_1672 (O_1672,N_23865,N_24165);
nor UO_1673 (O_1673,N_23851,N_24582);
and UO_1674 (O_1674,N_24357,N_24852);
xor UO_1675 (O_1675,N_24680,N_24531);
nand UO_1676 (O_1676,N_24955,N_24153);
xor UO_1677 (O_1677,N_24940,N_24355);
xnor UO_1678 (O_1678,N_24566,N_23801);
xnor UO_1679 (O_1679,N_24603,N_24074);
xnor UO_1680 (O_1680,N_24805,N_24578);
xnor UO_1681 (O_1681,N_24057,N_24212);
xnor UO_1682 (O_1682,N_24727,N_24655);
nor UO_1683 (O_1683,N_24671,N_24627);
xor UO_1684 (O_1684,N_24007,N_23876);
and UO_1685 (O_1685,N_24214,N_24145);
nand UO_1686 (O_1686,N_24448,N_24233);
or UO_1687 (O_1687,N_24268,N_24146);
nor UO_1688 (O_1688,N_24949,N_23767);
or UO_1689 (O_1689,N_23838,N_23756);
nor UO_1690 (O_1690,N_24824,N_24132);
nand UO_1691 (O_1691,N_23953,N_24881);
and UO_1692 (O_1692,N_24695,N_24560);
and UO_1693 (O_1693,N_23881,N_24204);
and UO_1694 (O_1694,N_24273,N_24013);
or UO_1695 (O_1695,N_24171,N_24250);
nand UO_1696 (O_1696,N_24608,N_23792);
nand UO_1697 (O_1697,N_24643,N_24356);
and UO_1698 (O_1698,N_24737,N_24320);
or UO_1699 (O_1699,N_24789,N_24242);
xnor UO_1700 (O_1700,N_23813,N_24719);
xnor UO_1701 (O_1701,N_23949,N_24121);
nand UO_1702 (O_1702,N_24779,N_23802);
nor UO_1703 (O_1703,N_24034,N_24711);
nand UO_1704 (O_1704,N_23997,N_23965);
or UO_1705 (O_1705,N_24033,N_24492);
or UO_1706 (O_1706,N_24442,N_24318);
nand UO_1707 (O_1707,N_24268,N_24303);
or UO_1708 (O_1708,N_24139,N_24080);
xnor UO_1709 (O_1709,N_24073,N_24601);
nor UO_1710 (O_1710,N_24295,N_24650);
and UO_1711 (O_1711,N_23783,N_24044);
and UO_1712 (O_1712,N_24625,N_24275);
and UO_1713 (O_1713,N_24730,N_24270);
nand UO_1714 (O_1714,N_24046,N_24733);
nand UO_1715 (O_1715,N_23830,N_24930);
nor UO_1716 (O_1716,N_24132,N_24907);
xnor UO_1717 (O_1717,N_24366,N_23780);
xor UO_1718 (O_1718,N_24821,N_24372);
or UO_1719 (O_1719,N_24206,N_24096);
nand UO_1720 (O_1720,N_23797,N_24840);
and UO_1721 (O_1721,N_24839,N_23927);
xnor UO_1722 (O_1722,N_24579,N_24538);
and UO_1723 (O_1723,N_24254,N_24353);
and UO_1724 (O_1724,N_24214,N_24552);
nor UO_1725 (O_1725,N_24612,N_24459);
xnor UO_1726 (O_1726,N_24948,N_23891);
or UO_1727 (O_1727,N_24653,N_24182);
and UO_1728 (O_1728,N_23941,N_24820);
or UO_1729 (O_1729,N_24383,N_24633);
nand UO_1730 (O_1730,N_23841,N_24869);
xnor UO_1731 (O_1731,N_24780,N_24384);
xor UO_1732 (O_1732,N_24690,N_24488);
xnor UO_1733 (O_1733,N_24452,N_24147);
and UO_1734 (O_1734,N_24929,N_24186);
or UO_1735 (O_1735,N_24994,N_23824);
or UO_1736 (O_1736,N_24069,N_23928);
nand UO_1737 (O_1737,N_23963,N_24532);
xor UO_1738 (O_1738,N_24088,N_23798);
or UO_1739 (O_1739,N_24466,N_24816);
or UO_1740 (O_1740,N_24491,N_23890);
nor UO_1741 (O_1741,N_24171,N_24389);
nor UO_1742 (O_1742,N_24858,N_24365);
xor UO_1743 (O_1743,N_24085,N_24171);
nand UO_1744 (O_1744,N_24958,N_24087);
and UO_1745 (O_1745,N_23970,N_24803);
xnor UO_1746 (O_1746,N_24755,N_24373);
nor UO_1747 (O_1747,N_24487,N_23977);
or UO_1748 (O_1748,N_24877,N_24189);
nand UO_1749 (O_1749,N_24903,N_23756);
or UO_1750 (O_1750,N_23781,N_24178);
xnor UO_1751 (O_1751,N_24862,N_24437);
or UO_1752 (O_1752,N_24057,N_24996);
and UO_1753 (O_1753,N_24879,N_23833);
or UO_1754 (O_1754,N_23866,N_24274);
nor UO_1755 (O_1755,N_24950,N_24580);
or UO_1756 (O_1756,N_24337,N_24653);
xor UO_1757 (O_1757,N_24212,N_24323);
nand UO_1758 (O_1758,N_24378,N_24506);
or UO_1759 (O_1759,N_23803,N_24079);
or UO_1760 (O_1760,N_23986,N_24539);
nand UO_1761 (O_1761,N_24349,N_24223);
xor UO_1762 (O_1762,N_24124,N_24190);
nand UO_1763 (O_1763,N_24198,N_24817);
or UO_1764 (O_1764,N_24134,N_24020);
nor UO_1765 (O_1765,N_24847,N_24441);
xor UO_1766 (O_1766,N_24947,N_24949);
xnor UO_1767 (O_1767,N_24651,N_24310);
nor UO_1768 (O_1768,N_24373,N_24459);
xnor UO_1769 (O_1769,N_24931,N_24843);
and UO_1770 (O_1770,N_24663,N_24340);
nor UO_1771 (O_1771,N_24019,N_24202);
or UO_1772 (O_1772,N_24942,N_24651);
nand UO_1773 (O_1773,N_24204,N_23947);
and UO_1774 (O_1774,N_23972,N_24820);
xnor UO_1775 (O_1775,N_24708,N_23944);
nor UO_1776 (O_1776,N_23991,N_24323);
xor UO_1777 (O_1777,N_23975,N_24758);
nor UO_1778 (O_1778,N_24341,N_23895);
or UO_1779 (O_1779,N_24943,N_23966);
xor UO_1780 (O_1780,N_24202,N_24595);
xnor UO_1781 (O_1781,N_24349,N_24393);
and UO_1782 (O_1782,N_24827,N_23976);
nand UO_1783 (O_1783,N_24188,N_23823);
or UO_1784 (O_1784,N_24753,N_24671);
xor UO_1785 (O_1785,N_24620,N_24499);
and UO_1786 (O_1786,N_24690,N_23947);
or UO_1787 (O_1787,N_24154,N_24569);
nor UO_1788 (O_1788,N_24674,N_24008);
and UO_1789 (O_1789,N_24223,N_24754);
and UO_1790 (O_1790,N_24198,N_23942);
xor UO_1791 (O_1791,N_23766,N_24250);
or UO_1792 (O_1792,N_24206,N_24953);
or UO_1793 (O_1793,N_24463,N_23832);
nand UO_1794 (O_1794,N_23894,N_24080);
nand UO_1795 (O_1795,N_24964,N_24114);
or UO_1796 (O_1796,N_24678,N_24544);
or UO_1797 (O_1797,N_24086,N_24085);
or UO_1798 (O_1798,N_24686,N_24871);
or UO_1799 (O_1799,N_23934,N_24279);
and UO_1800 (O_1800,N_24539,N_24131);
and UO_1801 (O_1801,N_23944,N_24306);
nor UO_1802 (O_1802,N_24672,N_24941);
nand UO_1803 (O_1803,N_23888,N_23930);
xor UO_1804 (O_1804,N_24163,N_24556);
xor UO_1805 (O_1805,N_24947,N_24113);
xor UO_1806 (O_1806,N_24397,N_24674);
or UO_1807 (O_1807,N_24459,N_23855);
nor UO_1808 (O_1808,N_24070,N_24871);
nor UO_1809 (O_1809,N_24940,N_24144);
nor UO_1810 (O_1810,N_24728,N_24551);
nand UO_1811 (O_1811,N_24577,N_24864);
nand UO_1812 (O_1812,N_24258,N_24865);
nand UO_1813 (O_1813,N_23880,N_23864);
and UO_1814 (O_1814,N_24057,N_24575);
or UO_1815 (O_1815,N_24273,N_23939);
and UO_1816 (O_1816,N_24029,N_24285);
nand UO_1817 (O_1817,N_24352,N_24636);
nor UO_1818 (O_1818,N_24244,N_23792);
or UO_1819 (O_1819,N_24594,N_24660);
nor UO_1820 (O_1820,N_24157,N_24985);
and UO_1821 (O_1821,N_24524,N_24848);
nor UO_1822 (O_1822,N_24435,N_24795);
xor UO_1823 (O_1823,N_24055,N_24965);
nor UO_1824 (O_1824,N_24668,N_24466);
nand UO_1825 (O_1825,N_24761,N_24347);
xor UO_1826 (O_1826,N_24860,N_24004);
and UO_1827 (O_1827,N_24058,N_24744);
nand UO_1828 (O_1828,N_24965,N_24345);
nand UO_1829 (O_1829,N_24361,N_24830);
nor UO_1830 (O_1830,N_24089,N_24294);
nand UO_1831 (O_1831,N_23838,N_24173);
or UO_1832 (O_1832,N_23951,N_24651);
or UO_1833 (O_1833,N_23945,N_24934);
or UO_1834 (O_1834,N_24955,N_24852);
nor UO_1835 (O_1835,N_24259,N_23888);
nor UO_1836 (O_1836,N_24078,N_24311);
nand UO_1837 (O_1837,N_24268,N_24881);
and UO_1838 (O_1838,N_24388,N_24241);
xnor UO_1839 (O_1839,N_24294,N_24266);
xor UO_1840 (O_1840,N_24841,N_24040);
nor UO_1841 (O_1841,N_23982,N_24709);
and UO_1842 (O_1842,N_23759,N_24323);
nand UO_1843 (O_1843,N_24869,N_24221);
and UO_1844 (O_1844,N_24135,N_24717);
xnor UO_1845 (O_1845,N_24233,N_24391);
nor UO_1846 (O_1846,N_23914,N_24333);
or UO_1847 (O_1847,N_24417,N_24329);
xor UO_1848 (O_1848,N_24768,N_24591);
or UO_1849 (O_1849,N_24197,N_24322);
or UO_1850 (O_1850,N_24175,N_24195);
or UO_1851 (O_1851,N_24242,N_23976);
or UO_1852 (O_1852,N_24315,N_24143);
or UO_1853 (O_1853,N_24406,N_24994);
nor UO_1854 (O_1854,N_24419,N_24040);
nor UO_1855 (O_1855,N_24174,N_24004);
nor UO_1856 (O_1856,N_24035,N_23812);
nand UO_1857 (O_1857,N_24616,N_23802);
nand UO_1858 (O_1858,N_23834,N_24595);
xnor UO_1859 (O_1859,N_24503,N_24851);
nor UO_1860 (O_1860,N_23799,N_24542);
nor UO_1861 (O_1861,N_24957,N_24093);
nor UO_1862 (O_1862,N_23782,N_24219);
and UO_1863 (O_1863,N_24580,N_24430);
nand UO_1864 (O_1864,N_24855,N_24792);
or UO_1865 (O_1865,N_24673,N_24378);
or UO_1866 (O_1866,N_24700,N_24510);
nor UO_1867 (O_1867,N_24770,N_24199);
or UO_1868 (O_1868,N_24085,N_24128);
and UO_1869 (O_1869,N_23954,N_24770);
or UO_1870 (O_1870,N_24455,N_24530);
xor UO_1871 (O_1871,N_24780,N_23879);
nand UO_1872 (O_1872,N_24095,N_23767);
nor UO_1873 (O_1873,N_24769,N_23959);
xor UO_1874 (O_1874,N_24719,N_24230);
nor UO_1875 (O_1875,N_23805,N_23826);
and UO_1876 (O_1876,N_23871,N_24064);
and UO_1877 (O_1877,N_23841,N_24694);
or UO_1878 (O_1878,N_24746,N_24573);
or UO_1879 (O_1879,N_24202,N_24083);
and UO_1880 (O_1880,N_24300,N_23919);
and UO_1881 (O_1881,N_24189,N_24220);
xor UO_1882 (O_1882,N_24253,N_24818);
and UO_1883 (O_1883,N_23811,N_24369);
and UO_1884 (O_1884,N_23868,N_24774);
or UO_1885 (O_1885,N_24514,N_24791);
or UO_1886 (O_1886,N_24124,N_24338);
nand UO_1887 (O_1887,N_24584,N_24530);
nor UO_1888 (O_1888,N_24162,N_24237);
nand UO_1889 (O_1889,N_24889,N_24077);
or UO_1890 (O_1890,N_23868,N_24031);
xor UO_1891 (O_1891,N_24592,N_24730);
nor UO_1892 (O_1892,N_24526,N_24116);
or UO_1893 (O_1893,N_24665,N_24154);
nor UO_1894 (O_1894,N_24061,N_24362);
nand UO_1895 (O_1895,N_23790,N_24448);
nor UO_1896 (O_1896,N_24486,N_24793);
nor UO_1897 (O_1897,N_23898,N_24070);
and UO_1898 (O_1898,N_24958,N_24374);
or UO_1899 (O_1899,N_23946,N_24679);
nor UO_1900 (O_1900,N_24763,N_23905);
nand UO_1901 (O_1901,N_24792,N_24214);
nand UO_1902 (O_1902,N_23945,N_24219);
and UO_1903 (O_1903,N_24690,N_24135);
and UO_1904 (O_1904,N_23776,N_24069);
nand UO_1905 (O_1905,N_24317,N_24766);
or UO_1906 (O_1906,N_24235,N_24636);
nand UO_1907 (O_1907,N_24971,N_24848);
nor UO_1908 (O_1908,N_24245,N_24931);
nand UO_1909 (O_1909,N_24627,N_24359);
nand UO_1910 (O_1910,N_24115,N_24113);
xor UO_1911 (O_1911,N_24047,N_24844);
nand UO_1912 (O_1912,N_23886,N_24156);
or UO_1913 (O_1913,N_24229,N_24973);
and UO_1914 (O_1914,N_24254,N_24808);
or UO_1915 (O_1915,N_24364,N_24888);
or UO_1916 (O_1916,N_24405,N_24757);
xnor UO_1917 (O_1917,N_24461,N_24556);
or UO_1918 (O_1918,N_24276,N_23847);
nand UO_1919 (O_1919,N_24045,N_23764);
xor UO_1920 (O_1920,N_24393,N_24055);
xor UO_1921 (O_1921,N_24262,N_24854);
nor UO_1922 (O_1922,N_24958,N_23868);
or UO_1923 (O_1923,N_24339,N_24646);
nand UO_1924 (O_1924,N_23804,N_24435);
and UO_1925 (O_1925,N_24471,N_24982);
nand UO_1926 (O_1926,N_24107,N_24611);
xor UO_1927 (O_1927,N_24122,N_24479);
xor UO_1928 (O_1928,N_24118,N_24616);
or UO_1929 (O_1929,N_24954,N_24060);
nor UO_1930 (O_1930,N_24216,N_24819);
nor UO_1931 (O_1931,N_24864,N_23832);
nor UO_1932 (O_1932,N_24789,N_23928);
nor UO_1933 (O_1933,N_24484,N_24859);
xor UO_1934 (O_1934,N_24298,N_24457);
xnor UO_1935 (O_1935,N_24522,N_24998);
and UO_1936 (O_1936,N_24554,N_24618);
xnor UO_1937 (O_1937,N_24541,N_24125);
nand UO_1938 (O_1938,N_24257,N_24195);
nor UO_1939 (O_1939,N_24109,N_24131);
or UO_1940 (O_1940,N_24604,N_24752);
nor UO_1941 (O_1941,N_24450,N_23891);
nor UO_1942 (O_1942,N_24559,N_24234);
or UO_1943 (O_1943,N_24562,N_24475);
or UO_1944 (O_1944,N_24430,N_24240);
nor UO_1945 (O_1945,N_24586,N_24307);
xnor UO_1946 (O_1946,N_24809,N_24096);
and UO_1947 (O_1947,N_24873,N_24182);
nor UO_1948 (O_1948,N_24009,N_24934);
nor UO_1949 (O_1949,N_23842,N_24095);
and UO_1950 (O_1950,N_24886,N_24983);
and UO_1951 (O_1951,N_24756,N_24300);
and UO_1952 (O_1952,N_24150,N_23857);
nor UO_1953 (O_1953,N_24569,N_24397);
and UO_1954 (O_1954,N_24073,N_24760);
nor UO_1955 (O_1955,N_24017,N_24239);
nand UO_1956 (O_1956,N_24456,N_23809);
xnor UO_1957 (O_1957,N_24911,N_23860);
or UO_1958 (O_1958,N_24502,N_24230);
and UO_1959 (O_1959,N_24908,N_24159);
xnor UO_1960 (O_1960,N_23905,N_24101);
nand UO_1961 (O_1961,N_23873,N_24942);
and UO_1962 (O_1962,N_24250,N_24622);
and UO_1963 (O_1963,N_23897,N_24309);
nand UO_1964 (O_1964,N_23864,N_23877);
xnor UO_1965 (O_1965,N_24004,N_24368);
nor UO_1966 (O_1966,N_24796,N_24041);
nor UO_1967 (O_1967,N_23816,N_24907);
nor UO_1968 (O_1968,N_24733,N_23774);
nand UO_1969 (O_1969,N_24004,N_24000);
nand UO_1970 (O_1970,N_24991,N_24119);
and UO_1971 (O_1971,N_24679,N_24715);
nor UO_1972 (O_1972,N_24582,N_24706);
and UO_1973 (O_1973,N_24202,N_24366);
and UO_1974 (O_1974,N_23764,N_24538);
xor UO_1975 (O_1975,N_24843,N_24989);
xnor UO_1976 (O_1976,N_23866,N_24087);
or UO_1977 (O_1977,N_24443,N_24440);
nor UO_1978 (O_1978,N_23814,N_24935);
or UO_1979 (O_1979,N_23812,N_24265);
nand UO_1980 (O_1980,N_23779,N_24779);
or UO_1981 (O_1981,N_23979,N_24350);
nor UO_1982 (O_1982,N_24504,N_24885);
and UO_1983 (O_1983,N_23803,N_24147);
nand UO_1984 (O_1984,N_24857,N_24625);
or UO_1985 (O_1985,N_24041,N_24532);
and UO_1986 (O_1986,N_24172,N_24710);
nor UO_1987 (O_1987,N_24311,N_24613);
nand UO_1988 (O_1988,N_24588,N_24645);
and UO_1989 (O_1989,N_24343,N_24168);
nand UO_1990 (O_1990,N_24598,N_24858);
xnor UO_1991 (O_1991,N_24060,N_24676);
or UO_1992 (O_1992,N_24951,N_24525);
nor UO_1993 (O_1993,N_24619,N_24466);
and UO_1994 (O_1994,N_23898,N_24670);
and UO_1995 (O_1995,N_24511,N_23832);
nand UO_1996 (O_1996,N_24225,N_24175);
and UO_1997 (O_1997,N_24679,N_24375);
nor UO_1998 (O_1998,N_24949,N_24590);
nor UO_1999 (O_1999,N_24870,N_24729);
and UO_2000 (O_2000,N_24936,N_24970);
xnor UO_2001 (O_2001,N_24060,N_23904);
xnor UO_2002 (O_2002,N_23796,N_24384);
nor UO_2003 (O_2003,N_24993,N_24696);
nor UO_2004 (O_2004,N_23949,N_24425);
nor UO_2005 (O_2005,N_23753,N_24349);
or UO_2006 (O_2006,N_24193,N_24493);
and UO_2007 (O_2007,N_24862,N_24817);
nor UO_2008 (O_2008,N_24300,N_24962);
xor UO_2009 (O_2009,N_24656,N_24419);
nor UO_2010 (O_2010,N_24998,N_24909);
nor UO_2011 (O_2011,N_24242,N_24130);
and UO_2012 (O_2012,N_24327,N_24630);
nor UO_2013 (O_2013,N_24724,N_24504);
and UO_2014 (O_2014,N_24547,N_24902);
nor UO_2015 (O_2015,N_24447,N_24137);
xor UO_2016 (O_2016,N_24680,N_24653);
and UO_2017 (O_2017,N_24484,N_23961);
xor UO_2018 (O_2018,N_24425,N_24238);
nor UO_2019 (O_2019,N_24121,N_24987);
nand UO_2020 (O_2020,N_23981,N_24813);
nand UO_2021 (O_2021,N_24963,N_24503);
or UO_2022 (O_2022,N_24508,N_24081);
and UO_2023 (O_2023,N_24236,N_23932);
and UO_2024 (O_2024,N_24583,N_24848);
nor UO_2025 (O_2025,N_24204,N_23825);
and UO_2026 (O_2026,N_24749,N_23979);
nand UO_2027 (O_2027,N_24090,N_24941);
xnor UO_2028 (O_2028,N_24284,N_24340);
nand UO_2029 (O_2029,N_24381,N_23783);
xor UO_2030 (O_2030,N_24997,N_24877);
and UO_2031 (O_2031,N_24059,N_24737);
or UO_2032 (O_2032,N_23921,N_24325);
or UO_2033 (O_2033,N_24669,N_24197);
nand UO_2034 (O_2034,N_24137,N_24380);
nor UO_2035 (O_2035,N_24786,N_24759);
or UO_2036 (O_2036,N_24634,N_23841);
xnor UO_2037 (O_2037,N_24545,N_24004);
xor UO_2038 (O_2038,N_24178,N_23772);
xor UO_2039 (O_2039,N_24704,N_24478);
nor UO_2040 (O_2040,N_24958,N_24401);
or UO_2041 (O_2041,N_23869,N_24447);
nor UO_2042 (O_2042,N_24329,N_24959);
and UO_2043 (O_2043,N_24577,N_24951);
and UO_2044 (O_2044,N_24317,N_24783);
or UO_2045 (O_2045,N_24117,N_24031);
nor UO_2046 (O_2046,N_24074,N_24863);
nand UO_2047 (O_2047,N_24292,N_24819);
nor UO_2048 (O_2048,N_24156,N_24987);
and UO_2049 (O_2049,N_23933,N_23752);
and UO_2050 (O_2050,N_24206,N_24726);
nand UO_2051 (O_2051,N_24164,N_24497);
nand UO_2052 (O_2052,N_23887,N_23842);
nand UO_2053 (O_2053,N_24477,N_24520);
nor UO_2054 (O_2054,N_24761,N_23999);
and UO_2055 (O_2055,N_24145,N_24017);
or UO_2056 (O_2056,N_24556,N_24941);
and UO_2057 (O_2057,N_24143,N_24020);
xor UO_2058 (O_2058,N_24815,N_24878);
and UO_2059 (O_2059,N_24277,N_24064);
nand UO_2060 (O_2060,N_24130,N_24388);
nand UO_2061 (O_2061,N_24146,N_23941);
and UO_2062 (O_2062,N_23782,N_23927);
and UO_2063 (O_2063,N_24041,N_24607);
xor UO_2064 (O_2064,N_24822,N_24749);
and UO_2065 (O_2065,N_23963,N_24079);
nand UO_2066 (O_2066,N_23915,N_24694);
or UO_2067 (O_2067,N_24544,N_24796);
nand UO_2068 (O_2068,N_24778,N_24686);
and UO_2069 (O_2069,N_24927,N_24075);
xor UO_2070 (O_2070,N_24474,N_23816);
nand UO_2071 (O_2071,N_23804,N_24059);
nor UO_2072 (O_2072,N_24264,N_24382);
or UO_2073 (O_2073,N_24628,N_24345);
nand UO_2074 (O_2074,N_24414,N_24549);
xor UO_2075 (O_2075,N_24531,N_23807);
and UO_2076 (O_2076,N_24556,N_24651);
xor UO_2077 (O_2077,N_24207,N_24627);
or UO_2078 (O_2078,N_24973,N_24439);
nand UO_2079 (O_2079,N_24640,N_24018);
nor UO_2080 (O_2080,N_24009,N_24683);
nand UO_2081 (O_2081,N_24624,N_23799);
xor UO_2082 (O_2082,N_23826,N_24443);
nand UO_2083 (O_2083,N_24449,N_23762);
nor UO_2084 (O_2084,N_24283,N_24091);
or UO_2085 (O_2085,N_23948,N_24962);
and UO_2086 (O_2086,N_24975,N_24719);
xor UO_2087 (O_2087,N_24352,N_24374);
and UO_2088 (O_2088,N_23952,N_24396);
nor UO_2089 (O_2089,N_24266,N_24615);
nor UO_2090 (O_2090,N_24665,N_24673);
nand UO_2091 (O_2091,N_24693,N_23843);
nor UO_2092 (O_2092,N_24836,N_24500);
nor UO_2093 (O_2093,N_24245,N_24042);
and UO_2094 (O_2094,N_23878,N_23959);
xnor UO_2095 (O_2095,N_23929,N_24743);
xor UO_2096 (O_2096,N_24286,N_24417);
nor UO_2097 (O_2097,N_23979,N_24127);
nand UO_2098 (O_2098,N_23876,N_24306);
nor UO_2099 (O_2099,N_24643,N_24772);
xor UO_2100 (O_2100,N_23926,N_23775);
or UO_2101 (O_2101,N_24077,N_23827);
xnor UO_2102 (O_2102,N_24036,N_24543);
xor UO_2103 (O_2103,N_24980,N_24141);
xnor UO_2104 (O_2104,N_24466,N_24345);
nand UO_2105 (O_2105,N_24465,N_24256);
and UO_2106 (O_2106,N_23944,N_24020);
nand UO_2107 (O_2107,N_24043,N_24074);
and UO_2108 (O_2108,N_24910,N_24233);
nand UO_2109 (O_2109,N_24331,N_24373);
or UO_2110 (O_2110,N_24865,N_24275);
or UO_2111 (O_2111,N_24661,N_23844);
and UO_2112 (O_2112,N_23761,N_24535);
xor UO_2113 (O_2113,N_23881,N_24602);
or UO_2114 (O_2114,N_24696,N_23800);
or UO_2115 (O_2115,N_24959,N_24023);
or UO_2116 (O_2116,N_23833,N_24785);
or UO_2117 (O_2117,N_23769,N_24250);
or UO_2118 (O_2118,N_23972,N_24079);
xnor UO_2119 (O_2119,N_24403,N_23948);
nor UO_2120 (O_2120,N_24039,N_24034);
and UO_2121 (O_2121,N_23968,N_24672);
and UO_2122 (O_2122,N_24725,N_24007);
or UO_2123 (O_2123,N_24530,N_24951);
xor UO_2124 (O_2124,N_23925,N_24010);
nor UO_2125 (O_2125,N_24365,N_24506);
xor UO_2126 (O_2126,N_24232,N_24043);
nand UO_2127 (O_2127,N_24219,N_23984);
nor UO_2128 (O_2128,N_24360,N_24832);
or UO_2129 (O_2129,N_24414,N_24267);
and UO_2130 (O_2130,N_23846,N_24915);
nor UO_2131 (O_2131,N_24723,N_24806);
and UO_2132 (O_2132,N_23882,N_23873);
nand UO_2133 (O_2133,N_23968,N_24332);
nor UO_2134 (O_2134,N_24822,N_24996);
xor UO_2135 (O_2135,N_24912,N_24154);
xnor UO_2136 (O_2136,N_23825,N_24752);
xor UO_2137 (O_2137,N_24694,N_23830);
xor UO_2138 (O_2138,N_23781,N_24642);
and UO_2139 (O_2139,N_24118,N_24310);
or UO_2140 (O_2140,N_24943,N_24463);
and UO_2141 (O_2141,N_24272,N_24981);
nand UO_2142 (O_2142,N_23915,N_24458);
or UO_2143 (O_2143,N_24783,N_24429);
nor UO_2144 (O_2144,N_24955,N_24815);
or UO_2145 (O_2145,N_24678,N_24515);
or UO_2146 (O_2146,N_23844,N_24038);
or UO_2147 (O_2147,N_24695,N_24119);
nand UO_2148 (O_2148,N_24374,N_24713);
or UO_2149 (O_2149,N_24478,N_24573);
nand UO_2150 (O_2150,N_24647,N_24735);
and UO_2151 (O_2151,N_24434,N_24796);
nand UO_2152 (O_2152,N_23834,N_24170);
and UO_2153 (O_2153,N_24286,N_24521);
xnor UO_2154 (O_2154,N_24427,N_23874);
nand UO_2155 (O_2155,N_24460,N_24850);
or UO_2156 (O_2156,N_24473,N_24498);
nand UO_2157 (O_2157,N_24328,N_24279);
nor UO_2158 (O_2158,N_23811,N_24365);
nand UO_2159 (O_2159,N_24692,N_24655);
or UO_2160 (O_2160,N_24963,N_24554);
or UO_2161 (O_2161,N_23910,N_24605);
nand UO_2162 (O_2162,N_24223,N_24300);
or UO_2163 (O_2163,N_24986,N_24337);
or UO_2164 (O_2164,N_24903,N_23807);
and UO_2165 (O_2165,N_24835,N_23844);
or UO_2166 (O_2166,N_23907,N_24897);
nand UO_2167 (O_2167,N_24932,N_24199);
nor UO_2168 (O_2168,N_23939,N_24562);
xor UO_2169 (O_2169,N_23998,N_24255);
nor UO_2170 (O_2170,N_24239,N_23851);
nor UO_2171 (O_2171,N_24567,N_24310);
nand UO_2172 (O_2172,N_24884,N_24481);
nand UO_2173 (O_2173,N_24224,N_23916);
xor UO_2174 (O_2174,N_24189,N_24295);
xor UO_2175 (O_2175,N_24733,N_24868);
and UO_2176 (O_2176,N_24251,N_24123);
nor UO_2177 (O_2177,N_23878,N_24886);
and UO_2178 (O_2178,N_24249,N_24685);
or UO_2179 (O_2179,N_24642,N_24439);
nor UO_2180 (O_2180,N_24457,N_24095);
or UO_2181 (O_2181,N_24103,N_23843);
nand UO_2182 (O_2182,N_24382,N_24372);
xnor UO_2183 (O_2183,N_24378,N_24278);
and UO_2184 (O_2184,N_24141,N_24156);
nor UO_2185 (O_2185,N_23852,N_24434);
xnor UO_2186 (O_2186,N_24573,N_24101);
xor UO_2187 (O_2187,N_24472,N_24062);
nand UO_2188 (O_2188,N_24426,N_24763);
nand UO_2189 (O_2189,N_24382,N_24923);
or UO_2190 (O_2190,N_24316,N_24758);
or UO_2191 (O_2191,N_24278,N_24672);
xor UO_2192 (O_2192,N_24976,N_24234);
xnor UO_2193 (O_2193,N_23890,N_24547);
xnor UO_2194 (O_2194,N_24327,N_23776);
xnor UO_2195 (O_2195,N_24156,N_24656);
and UO_2196 (O_2196,N_24786,N_24330);
nand UO_2197 (O_2197,N_24608,N_23929);
and UO_2198 (O_2198,N_24091,N_24489);
xor UO_2199 (O_2199,N_23846,N_24925);
or UO_2200 (O_2200,N_24977,N_24616);
and UO_2201 (O_2201,N_23798,N_24171);
nand UO_2202 (O_2202,N_24670,N_24439);
nor UO_2203 (O_2203,N_24617,N_24053);
or UO_2204 (O_2204,N_24908,N_24567);
xor UO_2205 (O_2205,N_24989,N_24015);
or UO_2206 (O_2206,N_24383,N_24995);
nor UO_2207 (O_2207,N_24958,N_24730);
nor UO_2208 (O_2208,N_24862,N_23975);
xnor UO_2209 (O_2209,N_24808,N_24275);
and UO_2210 (O_2210,N_24522,N_24881);
and UO_2211 (O_2211,N_23877,N_24872);
nor UO_2212 (O_2212,N_24009,N_24575);
nor UO_2213 (O_2213,N_24751,N_24670);
or UO_2214 (O_2214,N_24966,N_24796);
nand UO_2215 (O_2215,N_24101,N_24160);
xnor UO_2216 (O_2216,N_23971,N_23917);
and UO_2217 (O_2217,N_23828,N_24141);
and UO_2218 (O_2218,N_24905,N_24527);
nor UO_2219 (O_2219,N_24463,N_24393);
nor UO_2220 (O_2220,N_24372,N_24178);
xor UO_2221 (O_2221,N_24969,N_24415);
nand UO_2222 (O_2222,N_24193,N_23768);
or UO_2223 (O_2223,N_23963,N_24183);
xor UO_2224 (O_2224,N_24630,N_24321);
xnor UO_2225 (O_2225,N_24825,N_24237);
or UO_2226 (O_2226,N_24644,N_24164);
and UO_2227 (O_2227,N_24007,N_24411);
and UO_2228 (O_2228,N_24479,N_23914);
and UO_2229 (O_2229,N_24342,N_24318);
xnor UO_2230 (O_2230,N_24651,N_24040);
and UO_2231 (O_2231,N_24239,N_24582);
and UO_2232 (O_2232,N_24172,N_24181);
or UO_2233 (O_2233,N_24273,N_24935);
nor UO_2234 (O_2234,N_24882,N_24098);
nor UO_2235 (O_2235,N_24577,N_24894);
nand UO_2236 (O_2236,N_24350,N_24904);
xor UO_2237 (O_2237,N_24514,N_23876);
nand UO_2238 (O_2238,N_23931,N_24330);
nand UO_2239 (O_2239,N_24263,N_23788);
or UO_2240 (O_2240,N_24380,N_24598);
nand UO_2241 (O_2241,N_24155,N_24957);
xnor UO_2242 (O_2242,N_24210,N_24088);
nor UO_2243 (O_2243,N_24597,N_24079);
xor UO_2244 (O_2244,N_24227,N_24629);
nor UO_2245 (O_2245,N_24913,N_24063);
or UO_2246 (O_2246,N_24306,N_24828);
nand UO_2247 (O_2247,N_23872,N_24306);
nor UO_2248 (O_2248,N_24615,N_24732);
nor UO_2249 (O_2249,N_24565,N_24728);
nor UO_2250 (O_2250,N_24634,N_24387);
and UO_2251 (O_2251,N_23972,N_24255);
nor UO_2252 (O_2252,N_24185,N_24188);
nor UO_2253 (O_2253,N_24146,N_24841);
nor UO_2254 (O_2254,N_24364,N_24188);
and UO_2255 (O_2255,N_24321,N_24208);
or UO_2256 (O_2256,N_23774,N_24762);
and UO_2257 (O_2257,N_24182,N_24619);
or UO_2258 (O_2258,N_24273,N_24899);
and UO_2259 (O_2259,N_24679,N_24924);
and UO_2260 (O_2260,N_24150,N_24465);
nand UO_2261 (O_2261,N_24132,N_23939);
nand UO_2262 (O_2262,N_24487,N_24127);
or UO_2263 (O_2263,N_24850,N_24560);
nor UO_2264 (O_2264,N_24753,N_24402);
nor UO_2265 (O_2265,N_24079,N_24504);
or UO_2266 (O_2266,N_24260,N_24448);
and UO_2267 (O_2267,N_24400,N_24436);
or UO_2268 (O_2268,N_24833,N_24127);
nor UO_2269 (O_2269,N_23910,N_23793);
nand UO_2270 (O_2270,N_24402,N_24638);
and UO_2271 (O_2271,N_24927,N_24213);
nor UO_2272 (O_2272,N_23993,N_24375);
nor UO_2273 (O_2273,N_24861,N_23905);
and UO_2274 (O_2274,N_24680,N_24013);
nand UO_2275 (O_2275,N_24908,N_24524);
nand UO_2276 (O_2276,N_24851,N_23996);
or UO_2277 (O_2277,N_24517,N_24018);
xor UO_2278 (O_2278,N_24540,N_24934);
nand UO_2279 (O_2279,N_24673,N_24235);
nor UO_2280 (O_2280,N_24041,N_24398);
xnor UO_2281 (O_2281,N_24451,N_23818);
or UO_2282 (O_2282,N_24798,N_24907);
xnor UO_2283 (O_2283,N_23767,N_24054);
xor UO_2284 (O_2284,N_24862,N_23813);
nor UO_2285 (O_2285,N_24029,N_24830);
or UO_2286 (O_2286,N_24436,N_24763);
nand UO_2287 (O_2287,N_24977,N_24814);
or UO_2288 (O_2288,N_24855,N_23799);
or UO_2289 (O_2289,N_23934,N_24408);
or UO_2290 (O_2290,N_24870,N_23837);
xnor UO_2291 (O_2291,N_24586,N_24898);
nand UO_2292 (O_2292,N_24448,N_24966);
xor UO_2293 (O_2293,N_24553,N_24826);
and UO_2294 (O_2294,N_24516,N_24620);
xnor UO_2295 (O_2295,N_24445,N_24297);
xor UO_2296 (O_2296,N_24005,N_23766);
xor UO_2297 (O_2297,N_24566,N_23970);
xor UO_2298 (O_2298,N_24225,N_23843);
xnor UO_2299 (O_2299,N_23998,N_24614);
or UO_2300 (O_2300,N_24399,N_23881);
and UO_2301 (O_2301,N_23938,N_24287);
nor UO_2302 (O_2302,N_23909,N_23969);
and UO_2303 (O_2303,N_24616,N_23861);
and UO_2304 (O_2304,N_24423,N_24744);
xor UO_2305 (O_2305,N_24954,N_24504);
nand UO_2306 (O_2306,N_24242,N_24985);
xnor UO_2307 (O_2307,N_24453,N_24107);
nor UO_2308 (O_2308,N_24430,N_23883);
nor UO_2309 (O_2309,N_24596,N_24165);
xor UO_2310 (O_2310,N_24255,N_24432);
nor UO_2311 (O_2311,N_23943,N_24219);
xnor UO_2312 (O_2312,N_24350,N_24308);
and UO_2313 (O_2313,N_24739,N_24061);
or UO_2314 (O_2314,N_24917,N_24509);
nand UO_2315 (O_2315,N_24414,N_24845);
and UO_2316 (O_2316,N_23949,N_23846);
and UO_2317 (O_2317,N_23985,N_24765);
and UO_2318 (O_2318,N_24690,N_24293);
or UO_2319 (O_2319,N_24908,N_24510);
nand UO_2320 (O_2320,N_24076,N_24659);
or UO_2321 (O_2321,N_23752,N_24658);
xnor UO_2322 (O_2322,N_24656,N_24213);
nand UO_2323 (O_2323,N_24481,N_24862);
and UO_2324 (O_2324,N_24977,N_24664);
nor UO_2325 (O_2325,N_24876,N_23755);
nand UO_2326 (O_2326,N_23816,N_24145);
nand UO_2327 (O_2327,N_24523,N_24745);
nor UO_2328 (O_2328,N_24457,N_24562);
nor UO_2329 (O_2329,N_24060,N_24785);
and UO_2330 (O_2330,N_24668,N_24917);
xnor UO_2331 (O_2331,N_24960,N_24837);
xnor UO_2332 (O_2332,N_24520,N_24700);
nand UO_2333 (O_2333,N_24065,N_24412);
nor UO_2334 (O_2334,N_24646,N_24981);
xor UO_2335 (O_2335,N_24124,N_23930);
xor UO_2336 (O_2336,N_24120,N_24172);
nand UO_2337 (O_2337,N_24335,N_24009);
xor UO_2338 (O_2338,N_24303,N_24785);
and UO_2339 (O_2339,N_23978,N_24468);
or UO_2340 (O_2340,N_24921,N_24920);
and UO_2341 (O_2341,N_23872,N_24825);
nand UO_2342 (O_2342,N_24976,N_24660);
or UO_2343 (O_2343,N_24653,N_24290);
or UO_2344 (O_2344,N_24769,N_24269);
and UO_2345 (O_2345,N_24889,N_24041);
and UO_2346 (O_2346,N_24420,N_23859);
xor UO_2347 (O_2347,N_24747,N_24907);
xnor UO_2348 (O_2348,N_24051,N_24816);
nand UO_2349 (O_2349,N_23977,N_23812);
nand UO_2350 (O_2350,N_24631,N_23796);
xor UO_2351 (O_2351,N_24684,N_24328);
and UO_2352 (O_2352,N_24922,N_24659);
nor UO_2353 (O_2353,N_23991,N_24593);
and UO_2354 (O_2354,N_24154,N_24099);
and UO_2355 (O_2355,N_24432,N_24481);
nor UO_2356 (O_2356,N_23841,N_24163);
and UO_2357 (O_2357,N_24342,N_24860);
nand UO_2358 (O_2358,N_24406,N_24819);
nor UO_2359 (O_2359,N_24044,N_24574);
nand UO_2360 (O_2360,N_24216,N_24753);
or UO_2361 (O_2361,N_23799,N_24458);
xnor UO_2362 (O_2362,N_24552,N_24691);
nand UO_2363 (O_2363,N_24022,N_24116);
nand UO_2364 (O_2364,N_23995,N_23950);
nand UO_2365 (O_2365,N_24430,N_24458);
nand UO_2366 (O_2366,N_23809,N_24001);
or UO_2367 (O_2367,N_23781,N_24525);
xnor UO_2368 (O_2368,N_24576,N_24959);
or UO_2369 (O_2369,N_24512,N_24622);
nand UO_2370 (O_2370,N_24488,N_24597);
xor UO_2371 (O_2371,N_24905,N_24249);
or UO_2372 (O_2372,N_24498,N_24677);
nor UO_2373 (O_2373,N_24918,N_24142);
nand UO_2374 (O_2374,N_23769,N_24808);
xor UO_2375 (O_2375,N_24844,N_24283);
nor UO_2376 (O_2376,N_23816,N_24577);
or UO_2377 (O_2377,N_24108,N_23880);
or UO_2378 (O_2378,N_24341,N_24383);
nand UO_2379 (O_2379,N_24972,N_23824);
nand UO_2380 (O_2380,N_24392,N_24372);
nor UO_2381 (O_2381,N_24461,N_23852);
nand UO_2382 (O_2382,N_23853,N_24132);
and UO_2383 (O_2383,N_23880,N_23757);
and UO_2384 (O_2384,N_24735,N_24247);
nand UO_2385 (O_2385,N_24917,N_24393);
and UO_2386 (O_2386,N_24544,N_24675);
xnor UO_2387 (O_2387,N_24887,N_24785);
or UO_2388 (O_2388,N_24189,N_24917);
and UO_2389 (O_2389,N_24703,N_24516);
xnor UO_2390 (O_2390,N_24211,N_24957);
or UO_2391 (O_2391,N_23798,N_24732);
nand UO_2392 (O_2392,N_24666,N_24621);
nand UO_2393 (O_2393,N_24041,N_24382);
xor UO_2394 (O_2394,N_24195,N_24932);
nor UO_2395 (O_2395,N_24482,N_24190);
or UO_2396 (O_2396,N_23854,N_24861);
and UO_2397 (O_2397,N_24006,N_24853);
nand UO_2398 (O_2398,N_24895,N_24817);
xor UO_2399 (O_2399,N_24142,N_24197);
or UO_2400 (O_2400,N_24078,N_24224);
nor UO_2401 (O_2401,N_24240,N_24757);
xor UO_2402 (O_2402,N_24949,N_23799);
nor UO_2403 (O_2403,N_24791,N_23986);
and UO_2404 (O_2404,N_24417,N_24240);
nand UO_2405 (O_2405,N_24641,N_24725);
or UO_2406 (O_2406,N_24638,N_24883);
nor UO_2407 (O_2407,N_24736,N_23835);
or UO_2408 (O_2408,N_24335,N_24583);
and UO_2409 (O_2409,N_24300,N_24263);
nand UO_2410 (O_2410,N_24859,N_24469);
and UO_2411 (O_2411,N_24871,N_24143);
and UO_2412 (O_2412,N_24692,N_24364);
nand UO_2413 (O_2413,N_24190,N_23801);
or UO_2414 (O_2414,N_24192,N_24847);
or UO_2415 (O_2415,N_24609,N_24751);
nand UO_2416 (O_2416,N_24111,N_24445);
xnor UO_2417 (O_2417,N_24808,N_24369);
or UO_2418 (O_2418,N_24473,N_24385);
and UO_2419 (O_2419,N_24186,N_24549);
and UO_2420 (O_2420,N_24830,N_24430);
or UO_2421 (O_2421,N_24867,N_24296);
xnor UO_2422 (O_2422,N_24842,N_24553);
nand UO_2423 (O_2423,N_24152,N_24295);
nor UO_2424 (O_2424,N_24016,N_24959);
and UO_2425 (O_2425,N_24901,N_24921);
and UO_2426 (O_2426,N_24292,N_23781);
nand UO_2427 (O_2427,N_23897,N_24965);
nand UO_2428 (O_2428,N_23880,N_24592);
or UO_2429 (O_2429,N_24083,N_24734);
nand UO_2430 (O_2430,N_24059,N_24198);
nand UO_2431 (O_2431,N_24382,N_24098);
nand UO_2432 (O_2432,N_24708,N_23997);
nor UO_2433 (O_2433,N_24118,N_24787);
nand UO_2434 (O_2434,N_24937,N_23790);
and UO_2435 (O_2435,N_24847,N_23947);
nand UO_2436 (O_2436,N_24819,N_24098);
and UO_2437 (O_2437,N_24342,N_24325);
xnor UO_2438 (O_2438,N_24556,N_23851);
and UO_2439 (O_2439,N_24079,N_24670);
xor UO_2440 (O_2440,N_24236,N_24747);
or UO_2441 (O_2441,N_24266,N_23802);
xnor UO_2442 (O_2442,N_24840,N_23913);
nor UO_2443 (O_2443,N_24726,N_24002);
and UO_2444 (O_2444,N_24785,N_24547);
nand UO_2445 (O_2445,N_23849,N_24018);
nand UO_2446 (O_2446,N_24036,N_24402);
nand UO_2447 (O_2447,N_24133,N_24250);
xor UO_2448 (O_2448,N_24660,N_24173);
xnor UO_2449 (O_2449,N_24363,N_24341);
nor UO_2450 (O_2450,N_24666,N_24239);
nor UO_2451 (O_2451,N_24052,N_24803);
nor UO_2452 (O_2452,N_24220,N_24965);
nor UO_2453 (O_2453,N_24292,N_24073);
and UO_2454 (O_2454,N_24600,N_24555);
nand UO_2455 (O_2455,N_23984,N_24585);
and UO_2456 (O_2456,N_24133,N_24051);
nand UO_2457 (O_2457,N_24046,N_24304);
nand UO_2458 (O_2458,N_23828,N_24976);
xnor UO_2459 (O_2459,N_24002,N_24872);
or UO_2460 (O_2460,N_23917,N_24301);
and UO_2461 (O_2461,N_23930,N_24183);
xnor UO_2462 (O_2462,N_24146,N_24449);
and UO_2463 (O_2463,N_24074,N_23885);
nand UO_2464 (O_2464,N_23974,N_24969);
xor UO_2465 (O_2465,N_24822,N_24742);
and UO_2466 (O_2466,N_24850,N_24112);
xnor UO_2467 (O_2467,N_24823,N_24674);
and UO_2468 (O_2468,N_24595,N_24338);
and UO_2469 (O_2469,N_24816,N_23978);
xnor UO_2470 (O_2470,N_24414,N_24535);
xor UO_2471 (O_2471,N_24670,N_24719);
and UO_2472 (O_2472,N_24016,N_24166);
nand UO_2473 (O_2473,N_23817,N_24280);
nor UO_2474 (O_2474,N_24050,N_24729);
xnor UO_2475 (O_2475,N_24159,N_24340);
and UO_2476 (O_2476,N_24596,N_24814);
xnor UO_2477 (O_2477,N_24200,N_24103);
nor UO_2478 (O_2478,N_24550,N_23865);
and UO_2479 (O_2479,N_24687,N_24368);
and UO_2480 (O_2480,N_24888,N_24969);
nand UO_2481 (O_2481,N_24822,N_24962);
and UO_2482 (O_2482,N_24684,N_24597);
nand UO_2483 (O_2483,N_23902,N_24047);
nand UO_2484 (O_2484,N_23798,N_24633);
nor UO_2485 (O_2485,N_24864,N_24578);
xor UO_2486 (O_2486,N_24617,N_24194);
or UO_2487 (O_2487,N_24245,N_23772);
nor UO_2488 (O_2488,N_24650,N_24079);
nor UO_2489 (O_2489,N_24671,N_24460);
and UO_2490 (O_2490,N_24890,N_24036);
nor UO_2491 (O_2491,N_24603,N_24852);
xor UO_2492 (O_2492,N_24411,N_24377);
xor UO_2493 (O_2493,N_23956,N_24200);
nor UO_2494 (O_2494,N_24104,N_24199);
or UO_2495 (O_2495,N_24161,N_24248);
and UO_2496 (O_2496,N_24779,N_24640);
or UO_2497 (O_2497,N_24592,N_24700);
and UO_2498 (O_2498,N_23871,N_23844);
xor UO_2499 (O_2499,N_24882,N_24772);
or UO_2500 (O_2500,N_23891,N_24710);
xnor UO_2501 (O_2501,N_23780,N_24903);
and UO_2502 (O_2502,N_24208,N_23814);
or UO_2503 (O_2503,N_23809,N_24089);
or UO_2504 (O_2504,N_24127,N_24801);
nand UO_2505 (O_2505,N_24894,N_24798);
or UO_2506 (O_2506,N_24408,N_23939);
nand UO_2507 (O_2507,N_24627,N_24072);
or UO_2508 (O_2508,N_24878,N_24021);
xnor UO_2509 (O_2509,N_24637,N_24845);
and UO_2510 (O_2510,N_23854,N_24128);
xor UO_2511 (O_2511,N_24074,N_24233);
and UO_2512 (O_2512,N_24908,N_24255);
xnor UO_2513 (O_2513,N_24194,N_24709);
nand UO_2514 (O_2514,N_24776,N_24799);
nor UO_2515 (O_2515,N_24324,N_24496);
nor UO_2516 (O_2516,N_24804,N_24254);
and UO_2517 (O_2517,N_24542,N_23760);
nand UO_2518 (O_2518,N_23842,N_24333);
nand UO_2519 (O_2519,N_24547,N_23983);
xor UO_2520 (O_2520,N_24764,N_24784);
nand UO_2521 (O_2521,N_24676,N_24741);
or UO_2522 (O_2522,N_24984,N_23804);
nand UO_2523 (O_2523,N_24234,N_24846);
xor UO_2524 (O_2524,N_24475,N_24848);
nand UO_2525 (O_2525,N_23810,N_24891);
nand UO_2526 (O_2526,N_24619,N_23873);
and UO_2527 (O_2527,N_24419,N_23966);
and UO_2528 (O_2528,N_23838,N_24284);
nor UO_2529 (O_2529,N_24550,N_23856);
nand UO_2530 (O_2530,N_24109,N_24864);
nor UO_2531 (O_2531,N_24618,N_24445);
nor UO_2532 (O_2532,N_24067,N_23826);
or UO_2533 (O_2533,N_24554,N_24894);
or UO_2534 (O_2534,N_24313,N_23810);
nand UO_2535 (O_2535,N_24304,N_24940);
nand UO_2536 (O_2536,N_24670,N_23966);
and UO_2537 (O_2537,N_23945,N_24814);
and UO_2538 (O_2538,N_24542,N_23949);
and UO_2539 (O_2539,N_24817,N_24525);
nand UO_2540 (O_2540,N_23776,N_23852);
nand UO_2541 (O_2541,N_24008,N_24957);
nand UO_2542 (O_2542,N_24148,N_24213);
nor UO_2543 (O_2543,N_24948,N_24526);
xor UO_2544 (O_2544,N_24539,N_24233);
xor UO_2545 (O_2545,N_24611,N_24582);
nor UO_2546 (O_2546,N_24509,N_24344);
xnor UO_2547 (O_2547,N_23923,N_24158);
and UO_2548 (O_2548,N_24452,N_24826);
nand UO_2549 (O_2549,N_23890,N_24526);
nor UO_2550 (O_2550,N_24991,N_24497);
nor UO_2551 (O_2551,N_24054,N_24683);
nand UO_2552 (O_2552,N_24760,N_24968);
xor UO_2553 (O_2553,N_24632,N_24920);
nor UO_2554 (O_2554,N_24864,N_24902);
nor UO_2555 (O_2555,N_24470,N_24332);
nand UO_2556 (O_2556,N_24334,N_24314);
xnor UO_2557 (O_2557,N_24054,N_24021);
and UO_2558 (O_2558,N_24171,N_24149);
or UO_2559 (O_2559,N_23767,N_24321);
nand UO_2560 (O_2560,N_23876,N_24343);
xnor UO_2561 (O_2561,N_24879,N_24493);
xor UO_2562 (O_2562,N_24279,N_24865);
nor UO_2563 (O_2563,N_24613,N_24111);
and UO_2564 (O_2564,N_24510,N_24670);
nand UO_2565 (O_2565,N_24030,N_23788);
or UO_2566 (O_2566,N_24011,N_24204);
xor UO_2567 (O_2567,N_24452,N_24664);
xnor UO_2568 (O_2568,N_24656,N_23973);
or UO_2569 (O_2569,N_24406,N_23769);
and UO_2570 (O_2570,N_24278,N_24382);
nand UO_2571 (O_2571,N_24804,N_24854);
and UO_2572 (O_2572,N_24306,N_24737);
and UO_2573 (O_2573,N_24749,N_24425);
and UO_2574 (O_2574,N_24250,N_24505);
or UO_2575 (O_2575,N_24652,N_24220);
nor UO_2576 (O_2576,N_24317,N_24933);
nor UO_2577 (O_2577,N_24498,N_24534);
nor UO_2578 (O_2578,N_23798,N_24069);
or UO_2579 (O_2579,N_24615,N_23846);
nor UO_2580 (O_2580,N_24060,N_24398);
xnor UO_2581 (O_2581,N_24161,N_24778);
or UO_2582 (O_2582,N_24659,N_24455);
nor UO_2583 (O_2583,N_24225,N_24481);
and UO_2584 (O_2584,N_24898,N_24255);
and UO_2585 (O_2585,N_24357,N_24681);
nand UO_2586 (O_2586,N_24980,N_24677);
or UO_2587 (O_2587,N_23908,N_24763);
xor UO_2588 (O_2588,N_23908,N_23849);
xor UO_2589 (O_2589,N_24722,N_23847);
nor UO_2590 (O_2590,N_24942,N_24199);
nand UO_2591 (O_2591,N_24366,N_24268);
and UO_2592 (O_2592,N_23853,N_24214);
nor UO_2593 (O_2593,N_24009,N_24827);
and UO_2594 (O_2594,N_24970,N_23884);
xor UO_2595 (O_2595,N_24726,N_24455);
xor UO_2596 (O_2596,N_24733,N_24038);
and UO_2597 (O_2597,N_24238,N_24758);
or UO_2598 (O_2598,N_24917,N_23950);
or UO_2599 (O_2599,N_24186,N_24750);
xnor UO_2600 (O_2600,N_24719,N_24178);
xor UO_2601 (O_2601,N_24500,N_24383);
xor UO_2602 (O_2602,N_24225,N_24355);
nor UO_2603 (O_2603,N_24821,N_23872);
or UO_2604 (O_2604,N_24928,N_24516);
and UO_2605 (O_2605,N_24805,N_24590);
xor UO_2606 (O_2606,N_24337,N_24602);
and UO_2607 (O_2607,N_23988,N_24686);
and UO_2608 (O_2608,N_24877,N_24247);
nand UO_2609 (O_2609,N_24149,N_24002);
xnor UO_2610 (O_2610,N_24741,N_24265);
xor UO_2611 (O_2611,N_24261,N_23971);
or UO_2612 (O_2612,N_23946,N_23995);
or UO_2613 (O_2613,N_23952,N_24506);
and UO_2614 (O_2614,N_24300,N_24888);
xor UO_2615 (O_2615,N_24358,N_24428);
or UO_2616 (O_2616,N_24910,N_24816);
nor UO_2617 (O_2617,N_24645,N_24035);
nor UO_2618 (O_2618,N_24616,N_24524);
and UO_2619 (O_2619,N_24518,N_24866);
nand UO_2620 (O_2620,N_23827,N_24735);
nand UO_2621 (O_2621,N_24472,N_24602);
and UO_2622 (O_2622,N_24272,N_23858);
and UO_2623 (O_2623,N_24037,N_24448);
or UO_2624 (O_2624,N_24840,N_24426);
or UO_2625 (O_2625,N_24952,N_24490);
xor UO_2626 (O_2626,N_24561,N_24161);
or UO_2627 (O_2627,N_24519,N_24616);
and UO_2628 (O_2628,N_24214,N_23872);
xnor UO_2629 (O_2629,N_24589,N_24775);
and UO_2630 (O_2630,N_23784,N_24309);
nor UO_2631 (O_2631,N_24374,N_24253);
nor UO_2632 (O_2632,N_24806,N_23976);
and UO_2633 (O_2633,N_24324,N_24030);
nor UO_2634 (O_2634,N_24502,N_24781);
nand UO_2635 (O_2635,N_24121,N_24608);
nand UO_2636 (O_2636,N_24156,N_24812);
nor UO_2637 (O_2637,N_23957,N_24732);
nand UO_2638 (O_2638,N_24996,N_23931);
nor UO_2639 (O_2639,N_24340,N_24978);
xor UO_2640 (O_2640,N_24054,N_23927);
nor UO_2641 (O_2641,N_24864,N_24169);
xnor UO_2642 (O_2642,N_24372,N_23782);
and UO_2643 (O_2643,N_23839,N_23895);
xor UO_2644 (O_2644,N_24977,N_24622);
nor UO_2645 (O_2645,N_24639,N_24369);
xor UO_2646 (O_2646,N_24791,N_24626);
nand UO_2647 (O_2647,N_24548,N_24268);
and UO_2648 (O_2648,N_24806,N_24629);
or UO_2649 (O_2649,N_24202,N_24854);
nand UO_2650 (O_2650,N_24223,N_24729);
and UO_2651 (O_2651,N_24879,N_23975);
nand UO_2652 (O_2652,N_24954,N_24780);
and UO_2653 (O_2653,N_24541,N_23950);
xor UO_2654 (O_2654,N_24080,N_23928);
xnor UO_2655 (O_2655,N_24843,N_24905);
xnor UO_2656 (O_2656,N_23943,N_24955);
or UO_2657 (O_2657,N_24641,N_24024);
xnor UO_2658 (O_2658,N_23906,N_24961);
xor UO_2659 (O_2659,N_24875,N_24244);
nor UO_2660 (O_2660,N_23880,N_24375);
or UO_2661 (O_2661,N_23819,N_24756);
xor UO_2662 (O_2662,N_24340,N_23867);
xor UO_2663 (O_2663,N_24883,N_24650);
xor UO_2664 (O_2664,N_24914,N_24157);
and UO_2665 (O_2665,N_24968,N_24244);
and UO_2666 (O_2666,N_24357,N_23870);
or UO_2667 (O_2667,N_23781,N_24258);
nand UO_2668 (O_2668,N_23783,N_24489);
or UO_2669 (O_2669,N_24730,N_24208);
and UO_2670 (O_2670,N_24412,N_24242);
and UO_2671 (O_2671,N_23804,N_24524);
xor UO_2672 (O_2672,N_24889,N_24882);
and UO_2673 (O_2673,N_24864,N_23773);
xnor UO_2674 (O_2674,N_24419,N_24627);
or UO_2675 (O_2675,N_24611,N_24001);
xor UO_2676 (O_2676,N_24079,N_24213);
and UO_2677 (O_2677,N_24450,N_23765);
xor UO_2678 (O_2678,N_24566,N_24064);
and UO_2679 (O_2679,N_23873,N_24017);
xnor UO_2680 (O_2680,N_23815,N_24016);
or UO_2681 (O_2681,N_24602,N_24878);
nor UO_2682 (O_2682,N_24137,N_24561);
nand UO_2683 (O_2683,N_23958,N_24086);
xor UO_2684 (O_2684,N_24142,N_24666);
or UO_2685 (O_2685,N_23751,N_24050);
xnor UO_2686 (O_2686,N_23982,N_24719);
nand UO_2687 (O_2687,N_24090,N_23869);
or UO_2688 (O_2688,N_24119,N_23839);
or UO_2689 (O_2689,N_24698,N_23955);
nand UO_2690 (O_2690,N_24051,N_24711);
or UO_2691 (O_2691,N_24188,N_24824);
and UO_2692 (O_2692,N_24548,N_23767);
and UO_2693 (O_2693,N_24120,N_24483);
or UO_2694 (O_2694,N_24834,N_23876);
xor UO_2695 (O_2695,N_24921,N_24754);
nor UO_2696 (O_2696,N_24798,N_24423);
nor UO_2697 (O_2697,N_24794,N_24996);
nand UO_2698 (O_2698,N_23764,N_23984);
xnor UO_2699 (O_2699,N_24106,N_24360);
nand UO_2700 (O_2700,N_24482,N_24318);
xor UO_2701 (O_2701,N_24727,N_24988);
nor UO_2702 (O_2702,N_24540,N_23884);
xor UO_2703 (O_2703,N_24989,N_23841);
nand UO_2704 (O_2704,N_24814,N_23955);
and UO_2705 (O_2705,N_24213,N_24388);
nand UO_2706 (O_2706,N_24682,N_24412);
xor UO_2707 (O_2707,N_24020,N_24922);
xor UO_2708 (O_2708,N_24596,N_24499);
nand UO_2709 (O_2709,N_24474,N_23905);
and UO_2710 (O_2710,N_24850,N_24356);
nand UO_2711 (O_2711,N_24052,N_24685);
and UO_2712 (O_2712,N_24728,N_23840);
xnor UO_2713 (O_2713,N_24604,N_24501);
nand UO_2714 (O_2714,N_24146,N_24952);
or UO_2715 (O_2715,N_24239,N_24317);
and UO_2716 (O_2716,N_24777,N_24240);
xnor UO_2717 (O_2717,N_24844,N_24822);
or UO_2718 (O_2718,N_24451,N_24709);
and UO_2719 (O_2719,N_23830,N_24789);
nor UO_2720 (O_2720,N_24270,N_24077);
and UO_2721 (O_2721,N_24248,N_24728);
nand UO_2722 (O_2722,N_23895,N_24134);
xnor UO_2723 (O_2723,N_24672,N_23948);
nand UO_2724 (O_2724,N_24521,N_24539);
nor UO_2725 (O_2725,N_24780,N_24520);
or UO_2726 (O_2726,N_24542,N_24054);
and UO_2727 (O_2727,N_24885,N_24288);
or UO_2728 (O_2728,N_24879,N_23870);
and UO_2729 (O_2729,N_24417,N_24802);
and UO_2730 (O_2730,N_24713,N_24206);
nor UO_2731 (O_2731,N_24729,N_24391);
xnor UO_2732 (O_2732,N_24518,N_23990);
nand UO_2733 (O_2733,N_24103,N_24806);
nand UO_2734 (O_2734,N_24991,N_24433);
nor UO_2735 (O_2735,N_23920,N_24492);
nor UO_2736 (O_2736,N_24632,N_24349);
nand UO_2737 (O_2737,N_24257,N_24922);
and UO_2738 (O_2738,N_23809,N_23753);
nor UO_2739 (O_2739,N_23920,N_23849);
nand UO_2740 (O_2740,N_24772,N_24675);
and UO_2741 (O_2741,N_24196,N_23763);
xnor UO_2742 (O_2742,N_24356,N_24940);
or UO_2743 (O_2743,N_24599,N_24029);
nor UO_2744 (O_2744,N_24013,N_24187);
xor UO_2745 (O_2745,N_23967,N_24519);
and UO_2746 (O_2746,N_23907,N_24403);
or UO_2747 (O_2747,N_24913,N_24960);
and UO_2748 (O_2748,N_24564,N_24678);
nor UO_2749 (O_2749,N_23876,N_24115);
and UO_2750 (O_2750,N_24646,N_24050);
and UO_2751 (O_2751,N_23976,N_23950);
nor UO_2752 (O_2752,N_24346,N_24251);
xor UO_2753 (O_2753,N_23882,N_24762);
and UO_2754 (O_2754,N_24350,N_24527);
xnor UO_2755 (O_2755,N_24421,N_24266);
nand UO_2756 (O_2756,N_24702,N_24530);
xnor UO_2757 (O_2757,N_23909,N_23849);
xnor UO_2758 (O_2758,N_24017,N_24765);
and UO_2759 (O_2759,N_24435,N_24854);
nor UO_2760 (O_2760,N_24584,N_24218);
and UO_2761 (O_2761,N_23943,N_24312);
nor UO_2762 (O_2762,N_24755,N_23769);
nand UO_2763 (O_2763,N_24241,N_24452);
or UO_2764 (O_2764,N_24613,N_24974);
or UO_2765 (O_2765,N_24566,N_24217);
and UO_2766 (O_2766,N_24053,N_23895);
nor UO_2767 (O_2767,N_24687,N_24850);
nand UO_2768 (O_2768,N_24293,N_23825);
and UO_2769 (O_2769,N_24937,N_23799);
nor UO_2770 (O_2770,N_24977,N_24730);
nand UO_2771 (O_2771,N_24157,N_24048);
and UO_2772 (O_2772,N_24611,N_24778);
and UO_2773 (O_2773,N_23870,N_24413);
or UO_2774 (O_2774,N_24866,N_23967);
or UO_2775 (O_2775,N_24057,N_24254);
or UO_2776 (O_2776,N_24721,N_24894);
or UO_2777 (O_2777,N_24693,N_23962);
and UO_2778 (O_2778,N_24835,N_24308);
xor UO_2779 (O_2779,N_23857,N_24626);
nand UO_2780 (O_2780,N_24707,N_24734);
or UO_2781 (O_2781,N_24492,N_24298);
xor UO_2782 (O_2782,N_24102,N_23984);
and UO_2783 (O_2783,N_24119,N_24903);
or UO_2784 (O_2784,N_23886,N_23819);
xnor UO_2785 (O_2785,N_24681,N_24044);
xnor UO_2786 (O_2786,N_24433,N_24626);
nand UO_2787 (O_2787,N_24735,N_24178);
and UO_2788 (O_2788,N_24010,N_24036);
nand UO_2789 (O_2789,N_24753,N_24987);
nor UO_2790 (O_2790,N_24734,N_24256);
and UO_2791 (O_2791,N_24789,N_24129);
nand UO_2792 (O_2792,N_24123,N_23810);
xnor UO_2793 (O_2793,N_24346,N_23856);
xnor UO_2794 (O_2794,N_24840,N_23888);
nor UO_2795 (O_2795,N_24813,N_24956);
xnor UO_2796 (O_2796,N_24217,N_24201);
xor UO_2797 (O_2797,N_24300,N_24716);
or UO_2798 (O_2798,N_23778,N_24260);
nand UO_2799 (O_2799,N_24979,N_23920);
and UO_2800 (O_2800,N_24236,N_24091);
nor UO_2801 (O_2801,N_24433,N_24467);
xor UO_2802 (O_2802,N_24618,N_24790);
nand UO_2803 (O_2803,N_24399,N_24031);
nor UO_2804 (O_2804,N_23878,N_24829);
and UO_2805 (O_2805,N_24050,N_24436);
nand UO_2806 (O_2806,N_24287,N_24936);
nand UO_2807 (O_2807,N_24232,N_24587);
or UO_2808 (O_2808,N_24082,N_24215);
or UO_2809 (O_2809,N_24373,N_24731);
and UO_2810 (O_2810,N_24268,N_23837);
xor UO_2811 (O_2811,N_24539,N_24228);
xor UO_2812 (O_2812,N_24332,N_24569);
nor UO_2813 (O_2813,N_23922,N_24475);
nor UO_2814 (O_2814,N_24038,N_24041);
xor UO_2815 (O_2815,N_23887,N_24462);
nand UO_2816 (O_2816,N_24592,N_24659);
xnor UO_2817 (O_2817,N_24664,N_24602);
xnor UO_2818 (O_2818,N_24119,N_24190);
nor UO_2819 (O_2819,N_24091,N_23954);
and UO_2820 (O_2820,N_24866,N_23914);
and UO_2821 (O_2821,N_24445,N_24146);
xnor UO_2822 (O_2822,N_24348,N_24299);
xor UO_2823 (O_2823,N_23998,N_24770);
or UO_2824 (O_2824,N_24723,N_24741);
and UO_2825 (O_2825,N_24165,N_24339);
xnor UO_2826 (O_2826,N_24430,N_24789);
and UO_2827 (O_2827,N_24336,N_23941);
or UO_2828 (O_2828,N_24893,N_24176);
nor UO_2829 (O_2829,N_24001,N_24221);
nand UO_2830 (O_2830,N_23865,N_24011);
nor UO_2831 (O_2831,N_23995,N_24599);
nor UO_2832 (O_2832,N_24615,N_24351);
or UO_2833 (O_2833,N_24097,N_24050);
nor UO_2834 (O_2834,N_23803,N_24123);
nor UO_2835 (O_2835,N_24629,N_24359);
or UO_2836 (O_2836,N_24679,N_24308);
nand UO_2837 (O_2837,N_24052,N_24776);
nand UO_2838 (O_2838,N_24204,N_23828);
xor UO_2839 (O_2839,N_24664,N_23827);
nand UO_2840 (O_2840,N_24389,N_24842);
xor UO_2841 (O_2841,N_23891,N_24815);
xnor UO_2842 (O_2842,N_23773,N_24117);
and UO_2843 (O_2843,N_24050,N_24831);
nand UO_2844 (O_2844,N_23856,N_24111);
nand UO_2845 (O_2845,N_24517,N_24020);
and UO_2846 (O_2846,N_24905,N_24354);
and UO_2847 (O_2847,N_24804,N_24076);
nand UO_2848 (O_2848,N_24864,N_24508);
and UO_2849 (O_2849,N_24893,N_23945);
xnor UO_2850 (O_2850,N_24357,N_24723);
nand UO_2851 (O_2851,N_24853,N_24829);
nor UO_2852 (O_2852,N_23936,N_24473);
nor UO_2853 (O_2853,N_24877,N_24102);
and UO_2854 (O_2854,N_23819,N_24589);
and UO_2855 (O_2855,N_24079,N_24047);
xnor UO_2856 (O_2856,N_24324,N_24247);
nand UO_2857 (O_2857,N_24126,N_24423);
and UO_2858 (O_2858,N_24674,N_24562);
nor UO_2859 (O_2859,N_24548,N_23809);
xor UO_2860 (O_2860,N_24087,N_24969);
or UO_2861 (O_2861,N_23829,N_24880);
xnor UO_2862 (O_2862,N_23956,N_24252);
nand UO_2863 (O_2863,N_24723,N_24117);
xnor UO_2864 (O_2864,N_24978,N_24645);
xor UO_2865 (O_2865,N_24674,N_24773);
or UO_2866 (O_2866,N_24460,N_23998);
and UO_2867 (O_2867,N_24658,N_23766);
xnor UO_2868 (O_2868,N_24822,N_24964);
xor UO_2869 (O_2869,N_24247,N_24605);
xnor UO_2870 (O_2870,N_24419,N_23974);
nor UO_2871 (O_2871,N_24791,N_24121);
xnor UO_2872 (O_2872,N_24953,N_23898);
or UO_2873 (O_2873,N_23893,N_24617);
xnor UO_2874 (O_2874,N_24025,N_23919);
and UO_2875 (O_2875,N_24055,N_24755);
and UO_2876 (O_2876,N_24876,N_24682);
and UO_2877 (O_2877,N_24362,N_24142);
or UO_2878 (O_2878,N_24635,N_24828);
and UO_2879 (O_2879,N_24081,N_24276);
nand UO_2880 (O_2880,N_24597,N_23774);
nor UO_2881 (O_2881,N_24480,N_23781);
or UO_2882 (O_2882,N_24186,N_24704);
and UO_2883 (O_2883,N_24779,N_24521);
nand UO_2884 (O_2884,N_24450,N_23881);
or UO_2885 (O_2885,N_24177,N_24784);
xnor UO_2886 (O_2886,N_23865,N_24512);
nor UO_2887 (O_2887,N_23868,N_24573);
and UO_2888 (O_2888,N_24579,N_24486);
or UO_2889 (O_2889,N_24929,N_23793);
and UO_2890 (O_2890,N_24690,N_23966);
nand UO_2891 (O_2891,N_23752,N_23880);
nor UO_2892 (O_2892,N_24351,N_24642);
nand UO_2893 (O_2893,N_23957,N_24438);
nand UO_2894 (O_2894,N_24738,N_24335);
xor UO_2895 (O_2895,N_24634,N_24542);
or UO_2896 (O_2896,N_24413,N_24494);
nand UO_2897 (O_2897,N_24905,N_24316);
nand UO_2898 (O_2898,N_24053,N_24951);
xnor UO_2899 (O_2899,N_24113,N_24508);
and UO_2900 (O_2900,N_24883,N_24221);
or UO_2901 (O_2901,N_23752,N_24734);
and UO_2902 (O_2902,N_24609,N_24852);
nand UO_2903 (O_2903,N_23993,N_24363);
nand UO_2904 (O_2904,N_24007,N_24140);
and UO_2905 (O_2905,N_24350,N_24380);
and UO_2906 (O_2906,N_23938,N_23984);
and UO_2907 (O_2907,N_23770,N_24245);
nor UO_2908 (O_2908,N_24313,N_24984);
xnor UO_2909 (O_2909,N_24333,N_23806);
nand UO_2910 (O_2910,N_24873,N_24263);
or UO_2911 (O_2911,N_24189,N_24212);
nand UO_2912 (O_2912,N_24692,N_24214);
or UO_2913 (O_2913,N_24439,N_24127);
nand UO_2914 (O_2914,N_24737,N_24671);
xnor UO_2915 (O_2915,N_24196,N_24881);
and UO_2916 (O_2916,N_23876,N_24786);
xnor UO_2917 (O_2917,N_23966,N_24242);
or UO_2918 (O_2918,N_24342,N_24138);
nand UO_2919 (O_2919,N_24317,N_24956);
nand UO_2920 (O_2920,N_24239,N_23915);
or UO_2921 (O_2921,N_24781,N_24327);
nand UO_2922 (O_2922,N_24818,N_24142);
and UO_2923 (O_2923,N_24902,N_23995);
or UO_2924 (O_2924,N_23935,N_24722);
and UO_2925 (O_2925,N_23845,N_24414);
xnor UO_2926 (O_2926,N_24462,N_24975);
or UO_2927 (O_2927,N_24308,N_24134);
xor UO_2928 (O_2928,N_24748,N_24053);
or UO_2929 (O_2929,N_24870,N_24326);
nor UO_2930 (O_2930,N_24177,N_23892);
or UO_2931 (O_2931,N_23860,N_23890);
xor UO_2932 (O_2932,N_24552,N_24040);
and UO_2933 (O_2933,N_23902,N_24960);
or UO_2934 (O_2934,N_24219,N_24696);
nand UO_2935 (O_2935,N_24506,N_24523);
nor UO_2936 (O_2936,N_23825,N_23876);
xor UO_2937 (O_2937,N_24471,N_24723);
or UO_2938 (O_2938,N_24759,N_23928);
nand UO_2939 (O_2939,N_23956,N_23808);
and UO_2940 (O_2940,N_24454,N_24516);
nor UO_2941 (O_2941,N_24334,N_24155);
and UO_2942 (O_2942,N_23865,N_23916);
nand UO_2943 (O_2943,N_24370,N_24110);
nor UO_2944 (O_2944,N_24817,N_24124);
nor UO_2945 (O_2945,N_23949,N_23955);
nor UO_2946 (O_2946,N_24390,N_24626);
or UO_2947 (O_2947,N_24459,N_24776);
or UO_2948 (O_2948,N_24716,N_24425);
xor UO_2949 (O_2949,N_24509,N_23796);
or UO_2950 (O_2950,N_24973,N_24361);
or UO_2951 (O_2951,N_24091,N_24057);
xnor UO_2952 (O_2952,N_23908,N_23835);
nor UO_2953 (O_2953,N_24401,N_24878);
or UO_2954 (O_2954,N_24231,N_24840);
and UO_2955 (O_2955,N_24482,N_24263);
xnor UO_2956 (O_2956,N_24381,N_24736);
nor UO_2957 (O_2957,N_24317,N_24420);
and UO_2958 (O_2958,N_24234,N_24909);
and UO_2959 (O_2959,N_24386,N_24388);
or UO_2960 (O_2960,N_23755,N_23942);
or UO_2961 (O_2961,N_24944,N_24201);
nand UO_2962 (O_2962,N_24748,N_24003);
nand UO_2963 (O_2963,N_24603,N_24583);
xnor UO_2964 (O_2964,N_24467,N_23877);
nor UO_2965 (O_2965,N_23935,N_24659);
and UO_2966 (O_2966,N_24776,N_24311);
and UO_2967 (O_2967,N_24002,N_23913);
nand UO_2968 (O_2968,N_24323,N_24944);
nand UO_2969 (O_2969,N_24163,N_24943);
or UO_2970 (O_2970,N_24891,N_24622);
nand UO_2971 (O_2971,N_24755,N_24123);
and UO_2972 (O_2972,N_24972,N_24170);
or UO_2973 (O_2973,N_24635,N_24921);
xor UO_2974 (O_2974,N_24960,N_24867);
or UO_2975 (O_2975,N_24017,N_24503);
or UO_2976 (O_2976,N_24365,N_24782);
nand UO_2977 (O_2977,N_24775,N_24000);
nand UO_2978 (O_2978,N_23938,N_24323);
xor UO_2979 (O_2979,N_24939,N_24655);
xor UO_2980 (O_2980,N_23987,N_24288);
nor UO_2981 (O_2981,N_24896,N_24059);
xnor UO_2982 (O_2982,N_24083,N_24442);
nor UO_2983 (O_2983,N_24884,N_24526);
or UO_2984 (O_2984,N_24395,N_24409);
nor UO_2985 (O_2985,N_24968,N_24928);
or UO_2986 (O_2986,N_24986,N_24586);
or UO_2987 (O_2987,N_24041,N_24801);
nand UO_2988 (O_2988,N_24154,N_24322);
nand UO_2989 (O_2989,N_24167,N_24412);
and UO_2990 (O_2990,N_24203,N_23763);
and UO_2991 (O_2991,N_23939,N_24771);
and UO_2992 (O_2992,N_24393,N_23755);
or UO_2993 (O_2993,N_24296,N_24810);
or UO_2994 (O_2994,N_24664,N_24976);
nand UO_2995 (O_2995,N_24151,N_24956);
nor UO_2996 (O_2996,N_24530,N_24212);
nor UO_2997 (O_2997,N_24669,N_23969);
and UO_2998 (O_2998,N_24878,N_24613);
nand UO_2999 (O_2999,N_24356,N_24202);
endmodule