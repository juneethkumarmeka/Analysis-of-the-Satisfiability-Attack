module basic_1500_15000_2000_50_levels_10xor_6(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999;
nand U0 (N_0,In_774,In_210);
nand U1 (N_1,In_536,In_1088);
or U2 (N_2,In_1083,In_162);
and U3 (N_3,In_245,In_34);
xor U4 (N_4,In_105,In_575);
and U5 (N_5,In_967,In_1321);
xnor U6 (N_6,In_308,In_765);
and U7 (N_7,In_716,In_840);
nor U8 (N_8,In_60,In_289);
and U9 (N_9,In_1468,In_251);
and U10 (N_10,In_750,In_305);
nand U11 (N_11,In_612,In_992);
or U12 (N_12,In_880,In_703);
or U13 (N_13,In_257,In_1408);
nor U14 (N_14,In_1036,In_410);
or U15 (N_15,In_464,In_1396);
xnor U16 (N_16,In_1051,In_911);
xor U17 (N_17,In_600,In_1472);
and U18 (N_18,In_955,In_174);
or U19 (N_19,In_1336,In_824);
nor U20 (N_20,In_810,In_467);
and U21 (N_21,In_1459,In_482);
nand U22 (N_22,In_195,In_639);
or U23 (N_23,In_1290,In_404);
or U24 (N_24,In_486,In_31);
or U25 (N_25,In_673,In_391);
nand U26 (N_26,In_1369,In_772);
nand U27 (N_27,In_1042,In_879);
nand U28 (N_28,In_690,In_336);
nor U29 (N_29,In_958,In_281);
nand U30 (N_30,In_1143,In_1301);
and U31 (N_31,In_269,In_114);
nand U32 (N_32,In_295,In_469);
nand U33 (N_33,In_509,In_539);
nand U34 (N_34,In_571,In_1102);
xor U35 (N_35,In_1226,In_889);
nor U36 (N_36,In_679,In_1018);
and U37 (N_37,In_781,In_1441);
or U38 (N_38,In_1454,In_1490);
nand U39 (N_39,In_522,In_1469);
nand U40 (N_40,In_273,In_276);
and U41 (N_41,In_1116,In_595);
xor U42 (N_42,In_495,In_277);
or U43 (N_43,In_1305,In_1465);
xor U44 (N_44,In_294,In_483);
and U45 (N_45,In_392,In_325);
and U46 (N_46,In_922,In_1047);
nor U47 (N_47,In_1000,In_159);
nor U48 (N_48,In_903,In_650);
and U49 (N_49,In_88,In_1232);
nand U50 (N_50,In_364,In_437);
and U51 (N_51,In_1110,In_1195);
xor U52 (N_52,In_86,In_50);
and U53 (N_53,In_1428,In_492);
xor U54 (N_54,In_490,In_535);
nand U55 (N_55,In_488,In_828);
nand U56 (N_56,In_1164,In_1225);
or U57 (N_57,In_1265,In_1084);
nor U58 (N_58,In_523,In_1275);
xor U59 (N_59,In_1357,In_601);
nand U60 (N_60,In_823,In_939);
or U61 (N_61,In_1078,In_735);
nand U62 (N_62,In_183,In_951);
and U63 (N_63,In_950,In_450);
and U64 (N_64,In_1280,In_1160);
nor U65 (N_65,In_82,In_384);
nand U66 (N_66,In_1029,In_1244);
nor U67 (N_67,In_339,In_813);
nand U68 (N_68,In_701,In_783);
or U69 (N_69,In_15,In_444);
nor U70 (N_70,In_969,In_368);
xor U71 (N_71,In_332,In_386);
or U72 (N_72,In_1401,In_1363);
or U73 (N_73,In_1495,In_713);
or U74 (N_74,In_1438,In_1481);
xor U75 (N_75,In_373,In_1306);
and U76 (N_76,In_811,In_763);
nand U77 (N_77,In_1403,In_1256);
or U78 (N_78,In_362,In_876);
nand U79 (N_79,In_1138,In_1249);
and U80 (N_80,In_1020,In_704);
xnor U81 (N_81,In_948,In_1048);
or U82 (N_82,In_632,In_507);
nor U83 (N_83,In_1261,In_1482);
or U84 (N_84,In_663,In_1080);
nand U85 (N_85,In_1434,In_1033);
nand U86 (N_86,In_1317,In_1005);
or U87 (N_87,In_985,In_644);
xnor U88 (N_88,In_931,In_1485);
nand U89 (N_89,In_789,In_942);
or U90 (N_90,In_478,In_573);
nand U91 (N_91,In_285,In_1330);
nor U92 (N_92,In_725,In_794);
nand U93 (N_93,In_1057,In_293);
nor U94 (N_94,In_473,In_1156);
and U95 (N_95,In_1134,In_831);
xnor U96 (N_96,In_1219,In_1298);
and U97 (N_97,In_715,In_1151);
nor U98 (N_98,In_1340,In_1450);
nand U99 (N_99,In_381,In_407);
nand U100 (N_100,In_846,In_1121);
or U101 (N_101,In_420,In_652);
nand U102 (N_102,In_1262,In_378);
xnor U103 (N_103,In_1356,In_871);
xor U104 (N_104,In_1483,In_149);
xor U105 (N_105,In_57,In_1139);
or U106 (N_106,In_957,In_1133);
nand U107 (N_107,In_306,In_1115);
and U108 (N_108,In_1329,In_560);
or U109 (N_109,In_795,In_981);
xnor U110 (N_110,In_1235,In_1202);
xnor U111 (N_111,In_247,In_436);
and U112 (N_112,In_206,In_460);
nand U113 (N_113,In_1346,In_884);
xor U114 (N_114,In_702,In_812);
nor U115 (N_115,In_610,In_791);
or U116 (N_116,In_45,In_959);
xor U117 (N_117,In_401,In_1189);
nand U118 (N_118,In_904,In_833);
and U119 (N_119,In_1370,In_146);
nand U120 (N_120,In_1193,In_683);
or U121 (N_121,In_116,In_254);
nor U122 (N_122,In_790,In_572);
or U123 (N_123,In_870,In_80);
xor U124 (N_124,In_74,In_688);
or U125 (N_125,In_1291,In_141);
xor U126 (N_126,In_852,In_1263);
xor U127 (N_127,In_416,In_164);
or U128 (N_128,In_785,In_1386);
nor U129 (N_129,In_775,In_1268);
nand U130 (N_130,In_1090,In_1471);
nor U131 (N_131,In_236,In_102);
xor U132 (N_132,In_842,In_1400);
nand U133 (N_133,In_869,In_394);
and U134 (N_134,In_899,In_1347);
nor U135 (N_135,In_590,In_624);
xnor U136 (N_136,In_61,In_36);
nand U137 (N_137,In_798,In_500);
nor U138 (N_138,In_1251,In_565);
xor U139 (N_139,In_875,In_463);
or U140 (N_140,In_352,In_597);
and U141 (N_141,In_96,In_1382);
xor U142 (N_142,In_960,In_253);
xnor U143 (N_143,In_768,In_710);
nor U144 (N_144,In_1368,In_658);
nor U145 (N_145,In_479,In_95);
or U146 (N_146,In_949,In_1191);
xor U147 (N_147,In_426,In_711);
nor U148 (N_148,In_1049,In_203);
and U149 (N_149,In_278,In_941);
or U150 (N_150,In_1281,In_766);
nor U151 (N_151,In_973,In_1058);
nor U152 (N_152,In_1052,In_481);
nor U153 (N_153,In_909,In_1350);
xor U154 (N_154,In_705,In_890);
and U155 (N_155,In_48,In_707);
nand U156 (N_156,In_1435,In_1034);
and U157 (N_157,In_1070,In_970);
and U158 (N_158,In_54,In_648);
or U159 (N_159,In_1152,In_1276);
and U160 (N_160,In_168,In_1026);
and U161 (N_161,In_1066,In_487);
nand U162 (N_162,In_125,In_1008);
or U163 (N_163,In_261,In_804);
nor U164 (N_164,In_531,In_365);
nand U165 (N_165,In_435,In_173);
and U166 (N_166,In_1171,In_583);
xor U167 (N_167,In_671,In_591);
nor U168 (N_168,In_1079,In_1176);
nand U169 (N_169,In_7,In_406);
xnor U170 (N_170,In_1319,In_927);
and U171 (N_171,In_1073,In_240);
nor U172 (N_172,In_1241,In_402);
or U173 (N_173,In_20,In_627);
and U174 (N_174,In_1300,In_302);
or U175 (N_175,In_1109,In_71);
and U176 (N_176,In_1028,In_620);
nand U177 (N_177,In_917,In_1129);
nand U178 (N_178,In_1192,In_27);
nand U179 (N_179,In_337,In_579);
xor U180 (N_180,In_342,In_1492);
and U181 (N_181,In_1213,In_28);
xor U182 (N_182,In_631,In_1443);
xor U183 (N_183,In_980,In_241);
nor U184 (N_184,In_25,In_313);
xor U185 (N_185,In_264,In_1447);
nor U186 (N_186,In_510,In_1326);
xor U187 (N_187,In_457,In_986);
nor U188 (N_188,In_190,In_219);
nand U189 (N_189,In_11,In_1339);
and U190 (N_190,In_611,In_1407);
or U191 (N_191,In_314,In_316);
and U192 (N_192,In_643,In_1215);
nand U193 (N_193,In_641,In_636);
or U194 (N_194,In_218,In_1162);
xor U195 (N_195,In_1092,In_1168);
xor U196 (N_196,In_63,In_237);
and U197 (N_197,In_516,In_1214);
nand U198 (N_198,In_514,In_329);
xnor U199 (N_199,In_428,In_979);
xor U200 (N_200,In_576,In_1126);
nand U201 (N_201,In_398,In_258);
xor U202 (N_202,In_12,In_370);
nand U203 (N_203,In_820,In_533);
nand U204 (N_204,In_292,In_1453);
or U205 (N_205,In_217,In_230);
or U206 (N_206,In_966,In_1253);
nand U207 (N_207,In_945,In_1075);
and U208 (N_208,In_477,In_89);
xor U209 (N_209,In_1422,In_385);
xnor U210 (N_210,In_214,In_1136);
or U211 (N_211,In_607,In_838);
xnor U212 (N_212,In_300,In_1044);
and U213 (N_213,In_562,In_987);
or U214 (N_214,In_229,In_1433);
nand U215 (N_215,In_431,In_1361);
or U216 (N_216,In_578,In_603);
nor U217 (N_217,In_1313,In_1155);
nand U218 (N_218,In_642,In_260);
xor U219 (N_219,In_100,In_929);
and U220 (N_220,In_204,In_147);
xor U221 (N_221,In_892,In_1395);
nor U222 (N_222,In_1444,In_807);
xnor U223 (N_223,In_226,In_782);
nor U224 (N_224,In_433,In_693);
and U225 (N_225,In_1440,In_324);
xor U226 (N_226,In_1476,In_956);
nor U227 (N_227,In_676,In_496);
and U228 (N_228,In_517,In_1479);
and U229 (N_229,In_1056,In_994);
nand U230 (N_230,In_1285,In_803);
xor U231 (N_231,In_424,In_1413);
xnor U232 (N_232,In_24,In_863);
xor U233 (N_233,In_1394,In_443);
nand U234 (N_234,In_1446,In_609);
or U235 (N_235,In_1093,In_201);
nor U236 (N_236,In_749,In_882);
nor U237 (N_237,In_886,In_826);
and U238 (N_238,In_996,In_462);
xnor U239 (N_239,In_1274,In_982);
or U240 (N_240,In_1224,In_1296);
and U241 (N_241,In_593,In_282);
nand U242 (N_242,In_371,In_1098);
or U243 (N_243,In_35,In_170);
nor U244 (N_244,In_885,In_744);
nand U245 (N_245,In_596,In_221);
xnor U246 (N_246,In_532,In_568);
xor U247 (N_247,In_301,In_736);
and U248 (N_248,In_832,In_1242);
xor U249 (N_249,In_117,In_746);
or U250 (N_250,In_1266,In_1200);
xnor U251 (N_251,In_127,In_296);
nand U252 (N_252,In_505,In_1430);
and U253 (N_253,In_816,In_363);
nand U254 (N_254,In_1431,In_1295);
nor U255 (N_255,In_1166,In_235);
nor U256 (N_256,In_421,In_780);
xnor U257 (N_257,In_1384,In_920);
or U258 (N_258,In_1062,In_315);
nor U259 (N_259,In_318,In_312);
or U260 (N_260,In_861,In_1488);
nor U261 (N_261,In_757,In_604);
or U262 (N_262,In_938,In_65);
or U263 (N_263,In_1040,In_64);
nor U264 (N_264,In_847,In_860);
nand U265 (N_265,In_1167,In_694);
or U266 (N_266,In_1030,In_718);
or U267 (N_267,In_135,In_1470);
xor U268 (N_268,In_119,In_1123);
or U269 (N_269,In_1137,In_1383);
or U270 (N_270,In_359,In_354);
nor U271 (N_271,In_1074,In_23);
and U272 (N_272,In_42,In_274);
and U273 (N_273,In_376,In_76);
xor U274 (N_274,In_1072,In_1016);
nor U275 (N_275,In_825,In_223);
and U276 (N_276,In_341,In_255);
xor U277 (N_277,In_103,In_738);
nor U278 (N_278,In_19,In_954);
and U279 (N_279,In_1458,In_307);
nor U280 (N_280,In_144,In_788);
or U281 (N_281,In_549,In_724);
nor U282 (N_282,In_1053,In_429);
nand U283 (N_283,In_582,In_910);
xnor U284 (N_284,In_618,In_1333);
nor U285 (N_285,In_70,In_55);
and U286 (N_286,In_239,In_665);
nand U287 (N_287,In_1315,In_1304);
or U288 (N_288,In_913,In_585);
xnor U289 (N_289,In_111,In_1148);
xor U290 (N_290,In_918,In_1231);
nand U291 (N_291,In_1345,In_901);
and U292 (N_292,In_646,In_1038);
nand U293 (N_293,In_349,In_1452);
nand U294 (N_294,In_133,In_1427);
xor U295 (N_295,In_708,In_819);
or U296 (N_296,In_1130,In_850);
or U297 (N_297,In_543,In_343);
or U298 (N_298,In_1282,In_730);
xor U299 (N_299,In_234,In_353);
or U300 (N_300,In_1119,In_972);
or U301 (N_301,N_86,N_10);
and U302 (N_302,N_253,N_32);
and U303 (N_303,N_99,In_1194);
xnor U304 (N_304,In_280,In_962);
and U305 (N_305,In_108,N_73);
or U306 (N_306,N_96,In_1484);
nand U307 (N_307,N_57,In_1222);
or U308 (N_308,In_171,In_559);
or U309 (N_309,In_858,In_1218);
nor U310 (N_310,N_179,In_182);
nand U311 (N_311,In_242,In_1269);
nand U312 (N_312,In_761,In_1445);
nor U313 (N_313,N_24,In_461);
nand U314 (N_314,In_143,In_961);
or U315 (N_315,In_1323,N_31);
or U316 (N_316,In_1348,In_541);
and U317 (N_317,In_1294,N_201);
xor U318 (N_318,N_299,In_843);
nand U319 (N_319,In_1489,N_164);
nor U320 (N_320,In_706,In_120);
xnor U321 (N_321,N_55,In_654);
nor U322 (N_322,In_672,In_580);
nor U323 (N_323,In_66,N_59);
and U324 (N_324,N_0,In_995);
xnor U325 (N_325,In_914,In_835);
or U326 (N_326,In_212,N_7);
xnor U327 (N_327,N_44,In_335);
nand U328 (N_328,In_645,In_1397);
and U329 (N_329,In_1111,In_1095);
xnor U330 (N_330,In_1014,In_1010);
nor U331 (N_331,N_292,In_659);
and U332 (N_332,In_130,N_200);
or U333 (N_333,In_1420,In_474);
and U334 (N_334,N_88,In_1406);
xor U335 (N_335,In_664,In_334);
nand U336 (N_336,In_213,In_1353);
nand U337 (N_337,N_134,In_569);
xor U338 (N_338,In_608,In_1071);
nor U339 (N_339,N_276,In_403);
or U340 (N_340,In_647,In_767);
and U341 (N_341,N_245,In_37);
nand U342 (N_342,N_26,N_30);
nand U343 (N_343,In_1055,In_161);
or U344 (N_344,In_1343,N_252);
or U345 (N_345,In_309,In_106);
and U346 (N_346,In_1037,In_399);
or U347 (N_347,In_586,In_1318);
and U348 (N_348,In_881,In_267);
and U349 (N_349,N_85,In_243);
nor U350 (N_350,In_442,In_38);
nor U351 (N_351,In_198,In_1206);
nand U352 (N_352,In_943,In_1067);
xor U353 (N_353,N_266,In_321);
and U354 (N_354,In_734,N_289);
xor U355 (N_355,In_1497,In_682);
xnor U356 (N_356,N_177,In_1354);
or U357 (N_357,In_287,In_1365);
and U358 (N_358,In_771,N_20);
and U359 (N_359,N_291,N_283);
nand U360 (N_360,In_1196,N_9);
xnor U361 (N_361,In_1436,In_923);
nor U362 (N_362,In_501,In_379);
and U363 (N_363,In_452,In_263);
nor U364 (N_364,N_156,In_1157);
and U365 (N_365,N_255,In_908);
nand U366 (N_366,N_191,N_72);
or U367 (N_367,N_175,In_1077);
nand U368 (N_368,In_244,In_1417);
nor U369 (N_369,In_47,N_285);
or U370 (N_370,In_1355,In_21);
and U371 (N_371,In_755,In_515);
and U372 (N_372,In_1118,N_165);
or U373 (N_373,N_81,N_21);
xnor U374 (N_374,N_115,In_839);
nor U375 (N_375,In_1104,In_689);
nand U376 (N_376,In_1106,In_638);
nand U377 (N_377,In_1103,In_1292);
and U378 (N_378,In_169,In_445);
nor U379 (N_379,In_419,In_1019);
xnor U380 (N_380,N_92,In_976);
nand U381 (N_381,N_145,In_367);
nor U382 (N_382,In_1149,In_1412);
nor U383 (N_383,In_94,N_71);
nand U384 (N_384,N_279,N_89);
nand U385 (N_385,In_1204,In_151);
xor U386 (N_386,In_126,In_829);
or U387 (N_387,N_280,In_1388);
nand U388 (N_388,In_1087,In_1257);
or U389 (N_389,N_269,In_1374);
and U390 (N_390,In_556,N_181);
and U391 (N_391,In_1082,N_220);
or U392 (N_392,N_163,N_77);
and U393 (N_393,In_1174,In_1423);
nand U394 (N_394,In_1493,In_545);
nand U395 (N_395,In_1324,N_239);
xnor U396 (N_396,In_792,In_546);
nor U397 (N_397,In_1342,In_1494);
and U398 (N_398,In_484,In_1227);
xnor U399 (N_399,In_350,In_977);
nand U400 (N_400,In_844,In_347);
nand U401 (N_401,In_1277,In_92);
or U402 (N_402,In_947,In_1418);
xnor U403 (N_403,N_37,N_112);
or U404 (N_404,In_1158,N_4);
nor U405 (N_405,In_395,In_1212);
nor U406 (N_406,In_1007,N_287);
nor U407 (N_407,In_594,N_80);
or U408 (N_408,In_0,In_1352);
and U409 (N_409,In_856,In_605);
and U410 (N_410,In_374,In_1411);
nand U411 (N_411,In_513,In_696);
xor U412 (N_412,N_79,N_90);
xor U413 (N_413,In_1169,In_1175);
nand U414 (N_414,In_1108,In_1183);
or U415 (N_415,In_808,In_476);
or U416 (N_416,N_13,In_454);
and U417 (N_417,In_731,In_1096);
xor U418 (N_418,In_383,In_921);
or U419 (N_419,N_51,N_159);
and U420 (N_420,N_65,In_93);
nor U421 (N_421,N_62,In_382);
xor U422 (N_422,In_121,In_1011);
and U423 (N_423,In_1284,In_250);
or U424 (N_424,In_155,In_369);
nor U425 (N_425,In_1349,N_46);
nor U426 (N_426,N_206,In_1310);
or U427 (N_427,N_277,In_551);
nand U428 (N_428,In_916,N_243);
xnor U429 (N_429,In_104,In_1211);
or U430 (N_430,In_669,In_552);
and U431 (N_431,In_1230,N_2);
and U432 (N_432,N_34,In_475);
and U433 (N_433,N_202,N_39);
xor U434 (N_434,In_160,In_98);
nand U435 (N_435,In_388,In_786);
nor U436 (N_436,In_153,In_319);
nand U437 (N_437,N_122,In_157);
nor U438 (N_438,N_263,In_1069);
nor U439 (N_439,N_161,N_211);
and U440 (N_440,In_998,In_150);
xor U441 (N_441,N_108,In_864);
and U442 (N_442,N_149,N_148);
nand U443 (N_443,N_60,In_323);
xnor U444 (N_444,In_599,N_53);
or U445 (N_445,In_113,In_112);
and U446 (N_446,In_259,N_273);
xor U447 (N_447,In_32,In_1101);
nor U448 (N_448,In_723,In_529);
nor U449 (N_449,In_1405,In_859);
nor U450 (N_450,N_33,In_547);
nand U451 (N_451,In_284,N_249);
xnor U452 (N_452,In_619,N_267);
and U453 (N_453,In_651,N_133);
nor U454 (N_454,N_111,In_1208);
or U455 (N_455,In_1061,N_128);
nor U456 (N_456,In_97,In_926);
and U457 (N_457,In_1320,In_233);
nand U458 (N_458,In_1,N_70);
and U459 (N_459,In_1337,In_439);
xnor U460 (N_460,In_1364,In_412);
and U461 (N_461,N_187,In_299);
nor U462 (N_462,In_1247,In_784);
nor U463 (N_463,In_1351,In_657);
or U464 (N_464,In_1089,N_69);
nand U465 (N_465,In_1135,In_666);
xor U466 (N_466,In_1238,In_1376);
nor U467 (N_467,In_733,In_1437);
xor U468 (N_468,In_200,N_188);
or U469 (N_469,N_208,In_326);
nand U470 (N_470,In_246,In_1163);
nor U471 (N_471,In_91,N_215);
nand U472 (N_472,In_1178,N_8);
nor U473 (N_473,In_118,In_304);
nor U474 (N_474,In_851,N_125);
and U475 (N_475,N_48,In_1059);
xor U476 (N_476,In_361,N_235);
and U477 (N_477,N_218,In_577);
and U478 (N_478,In_272,In_145);
nand U479 (N_479,In_1462,In_49);
or U480 (N_480,In_194,In_331);
or U481 (N_481,In_53,In_732);
nand U482 (N_482,In_1477,In_540);
xor U483 (N_483,In_1460,In_1409);
or U484 (N_484,In_1228,In_465);
nor U485 (N_485,N_56,N_262);
nand U486 (N_486,N_16,In_874);
and U487 (N_487,N_143,N_93);
nor U488 (N_488,In_360,In_697);
xnor U489 (N_489,In_466,In_357);
nor U490 (N_490,In_896,In_472);
nor U491 (N_491,N_294,In_1022);
or U492 (N_492,In_558,N_141);
nand U493 (N_493,In_900,In_887);
nor U494 (N_494,In_830,In_743);
or U495 (N_495,In_177,In_667);
or U496 (N_496,In_275,N_84);
xnor U497 (N_497,In_494,In_628);
nand U498 (N_498,N_258,N_256);
nand U499 (N_499,N_36,In_470);
xnor U500 (N_500,In_1377,In_208);
nand U501 (N_501,In_993,In_39);
nor U502 (N_502,In_22,N_50);
nand U503 (N_503,In_418,In_1076);
or U504 (N_504,In_566,In_185);
xnor U505 (N_505,In_8,N_66);
xnor U506 (N_506,In_563,In_504);
or U507 (N_507,In_1498,In_1378);
nand U508 (N_508,N_98,N_157);
or U509 (N_509,In_207,In_1267);
and U510 (N_510,In_897,In_834);
or U511 (N_511,In_1201,In_1021);
and U512 (N_512,In_1127,N_212);
nand U513 (N_513,In_303,In_317);
and U514 (N_514,In_988,N_282);
and U515 (N_515,In_1054,N_268);
and U516 (N_516,In_393,In_935);
or U517 (N_517,In_493,In_1017);
nor U518 (N_518,In_936,N_295);
and U519 (N_519,In_451,N_248);
nand U520 (N_520,In_1147,In_564);
or U521 (N_521,In_1186,In_574);
and U522 (N_522,In_1264,In_1327);
or U523 (N_523,In_762,In_542);
nand U524 (N_524,N_203,In_753);
xor U525 (N_525,N_124,In_649);
nand U526 (N_526,In_184,In_101);
nand U527 (N_527,N_25,In_1117);
nand U528 (N_528,In_1181,N_42);
and U529 (N_529,In_148,In_888);
nor U530 (N_530,N_63,N_233);
nand U531 (N_531,In_425,In_983);
nand U532 (N_532,In_1198,In_290);
nor U533 (N_533,In_46,In_167);
nand U534 (N_534,N_217,In_924);
nor U535 (N_535,In_188,In_422);
or U536 (N_536,In_415,In_2);
nor U537 (N_537,In_1322,In_742);
nor U538 (N_538,In_202,In_625);
xnor U539 (N_539,In_554,In_1451);
nor U540 (N_540,In_737,In_1332);
nand U541 (N_541,N_118,In_1172);
and U542 (N_542,N_91,N_286);
nand U543 (N_543,N_12,In_634);
xnor U544 (N_544,In_99,In_1288);
nor U545 (N_545,N_107,In_1113);
or U546 (N_546,In_770,N_147);
nor U547 (N_547,In_441,In_686);
xor U548 (N_548,In_1091,In_1448);
or U549 (N_549,N_284,In_796);
and U550 (N_550,In_1125,N_126);
nand U551 (N_551,In_131,In_538);
nor U552 (N_552,In_152,In_1421);
and U553 (N_553,N_189,In_739);
nand U554 (N_554,In_1128,In_526);
nor U555 (N_555,N_209,In_351);
nand U556 (N_556,In_1278,In_512);
and U557 (N_557,In_1414,In_934);
or U558 (N_558,In_209,N_173);
nand U559 (N_559,In_142,In_1245);
nand U560 (N_560,N_241,N_250);
or U561 (N_561,N_182,In_912);
or U562 (N_562,N_199,In_1404);
nand U563 (N_563,N_45,In_1486);
xnor U564 (N_564,In_915,In_1252);
nand U565 (N_565,In_256,In_266);
or U566 (N_566,In_802,In_175);
xnor U567 (N_567,In_1105,N_227);
xnor U568 (N_568,In_878,In_1272);
or U569 (N_569,In_511,In_506);
nand U570 (N_570,In_974,N_52);
nand U571 (N_571,In_837,In_660);
and U572 (N_572,In_137,In_44);
and U573 (N_573,In_197,In_1311);
nand U574 (N_574,In_1132,In_989);
nand U575 (N_575,N_130,In_1273);
xnor U576 (N_576,In_907,In_1372);
nand U577 (N_577,In_930,In_1146);
nand U578 (N_578,In_894,In_67);
xor U579 (N_579,In_355,In_854);
nor U580 (N_580,N_74,In_1496);
nand U581 (N_581,In_158,In_172);
and U582 (N_582,In_1025,In_968);
nand U583 (N_583,N_137,In_1112);
nor U584 (N_584,In_115,N_222);
nor U585 (N_585,In_971,In_700);
nor U586 (N_586,In_1424,In_1254);
nor U587 (N_587,N_261,In_1250);
xnor U588 (N_588,In_822,N_281);
xor U589 (N_589,N_297,In_944);
xor U590 (N_590,N_192,In_51);
nor U591 (N_591,In_758,N_109);
nand U592 (N_592,In_1279,In_138);
nor U593 (N_593,In_937,In_128);
and U594 (N_594,In_166,N_228);
or U595 (N_595,In_189,In_773);
nor U596 (N_596,N_61,N_101);
xor U597 (N_597,In_748,In_390);
or U598 (N_598,In_1154,In_1107);
nor U599 (N_599,In_637,In_196);
nand U600 (N_600,In_1473,N_207);
and U601 (N_601,In_584,In_163);
or U602 (N_602,N_594,N_254);
nand U603 (N_603,N_22,N_364);
nor U604 (N_604,N_1,In_1380);
or U605 (N_605,In_283,N_553);
nand U606 (N_606,N_437,N_470);
nand U607 (N_607,In_187,N_471);
xnor U608 (N_608,N_311,N_324);
and U609 (N_609,In_699,In_1475);
xnor U610 (N_610,In_1381,N_154);
nand U611 (N_611,N_353,In_1203);
or U612 (N_612,N_598,In_616);
or U613 (N_613,In_893,N_338);
and U614 (N_614,In_1187,In_87);
or U615 (N_615,N_365,In_633);
or U616 (N_616,In_434,N_373);
and U617 (N_617,In_40,N_534);
or U618 (N_618,In_1302,In_62);
xnor U619 (N_619,N_350,In_1419);
xor U620 (N_620,N_378,N_240);
nor U621 (N_621,In_787,N_585);
or U622 (N_622,N_396,N_376);
or U623 (N_623,In_225,In_653);
nand U624 (N_624,N_275,N_117);
and U625 (N_625,In_1032,In_866);
and U626 (N_626,In_891,In_340);
nand U627 (N_627,N_583,In_1499);
nand U628 (N_628,In_1463,In_1124);
nand U629 (N_629,N_447,In_447);
xnor U630 (N_630,In_1165,In_1131);
nor U631 (N_631,N_290,In_1012);
and U632 (N_632,In_978,In_408);
or U633 (N_633,N_131,N_526);
xor U634 (N_634,N_388,In_1006);
nor U635 (N_635,N_488,N_19);
or U636 (N_636,In_1309,N_18);
nor U637 (N_637,N_216,N_544);
xnor U638 (N_638,In_1210,In_1297);
nand U639 (N_639,In_1050,In_192);
nand U640 (N_640,N_404,N_567);
and U641 (N_641,N_418,In_1328);
and U642 (N_642,N_225,N_95);
nand U643 (N_643,N_473,In_1046);
nand U644 (N_644,In_75,N_416);
xnor U645 (N_645,N_476,N_270);
and U646 (N_646,In_925,N_41);
and U647 (N_647,N_409,In_489);
and U648 (N_648,N_231,N_423);
nor U649 (N_649,N_491,In_867);
nor U650 (N_650,N_555,N_441);
nor U651 (N_651,In_220,N_412);
or U652 (N_652,In_1389,N_482);
xor U653 (N_653,In_503,In_59);
or U654 (N_654,In_1338,In_1255);
nand U655 (N_655,In_81,N_509);
or U656 (N_656,In_1344,N_574);
nor U657 (N_657,In_1170,N_139);
or U658 (N_658,N_307,N_410);
xor U659 (N_659,In_405,N_543);
nor U660 (N_660,N_563,In_1043);
or U661 (N_661,In_107,In_83);
and U662 (N_662,N_466,In_853);
nor U663 (N_663,In_779,N_27);
xnor U664 (N_664,N_510,In_898);
nand U665 (N_665,N_438,N_226);
nand U666 (N_666,N_310,N_460);
nand U667 (N_667,In_1426,N_369);
nor U668 (N_668,N_427,In_238);
and U669 (N_669,In_933,N_195);
or U670 (N_670,In_677,In_799);
nor U671 (N_671,N_426,N_352);
and U672 (N_672,In_684,N_76);
or U673 (N_673,In_855,In_181);
or U674 (N_674,In_1335,N_152);
xnor U675 (N_675,N_448,N_104);
and U676 (N_676,N_459,N_102);
nand U677 (N_677,In_1161,In_905);
or U678 (N_678,In_1229,In_519);
nand U679 (N_679,In_17,N_545);
nor U680 (N_680,In_10,N_340);
nand U681 (N_681,In_698,N_486);
nor U682 (N_682,In_1270,N_524);
xnor U683 (N_683,In_491,In_1027);
nor U684 (N_684,In_179,N_481);
and U685 (N_685,In_997,N_158);
xnor U686 (N_686,In_1120,N_257);
nor U687 (N_687,N_576,N_452);
nor U688 (N_688,In_5,N_308);
xor U689 (N_689,In_685,N_106);
xor U690 (N_690,N_453,N_484);
nand U691 (N_691,In_1003,N_508);
and U692 (N_692,In_3,In_1243);
xnor U693 (N_693,In_1039,In_26);
nor U694 (N_694,N_430,N_329);
and U695 (N_695,In_1140,N_123);
xor U696 (N_696,In_79,In_311);
or U697 (N_697,In_1220,N_361);
xor U698 (N_698,In_695,N_530);
or U699 (N_699,In_1190,In_836);
and U700 (N_700,N_569,In_640);
nand U701 (N_701,N_325,N_330);
xnor U702 (N_702,N_238,In_722);
or U703 (N_703,In_109,In_186);
nor U704 (N_704,N_549,In_1480);
and U705 (N_705,N_120,N_537);
nor U706 (N_706,In_530,N_337);
nor U707 (N_707,In_1177,N_5);
xor U708 (N_708,N_516,In_320);
and U709 (N_709,N_171,In_806);
nor U710 (N_710,In_1429,In_747);
nor U711 (N_711,N_597,N_523);
xnor U712 (N_712,N_205,N_110);
xnor U713 (N_713,N_464,N_587);
or U714 (N_714,N_445,N_363);
or U715 (N_715,N_334,In_1416);
and U716 (N_716,N_301,In_1236);
or U717 (N_717,N_496,In_760);
xor U718 (N_718,N_505,In_30);
or U719 (N_719,N_132,N_540);
nor U720 (N_720,N_54,In_1086);
nor U721 (N_721,N_43,In_1197);
xor U722 (N_722,N_506,N_390);
and U723 (N_723,In_1442,In_199);
and U724 (N_724,In_29,In_176);
nand U725 (N_725,In_124,In_122);
xnor U726 (N_726,N_136,N_467);
nor U727 (N_727,In_726,N_454);
or U728 (N_728,In_1015,N_527);
xor U729 (N_729,N_113,In_1325);
xnor U730 (N_730,N_213,N_579);
or U731 (N_731,In_1188,N_370);
nor U732 (N_732,N_229,In_110);
nand U733 (N_733,In_821,N_146);
nor U734 (N_734,In_224,In_553);
xor U735 (N_735,In_814,In_377);
nor U736 (N_736,N_483,N_15);
nand U737 (N_737,In_90,N_393);
nand U738 (N_738,N_23,In_946);
nand U739 (N_739,N_347,In_1002);
nand U740 (N_740,N_381,In_759);
or U741 (N_741,In_1004,In_227);
or U742 (N_742,In_629,N_6);
nand U743 (N_743,N_194,In_740);
nand U744 (N_744,In_588,N_372);
and U745 (N_745,In_271,In_1293);
and U746 (N_746,N_64,N_475);
or U747 (N_747,N_414,N_489);
xnor U748 (N_748,In_1246,In_841);
and U749 (N_749,In_123,In_1314);
and U750 (N_750,In_745,In_1001);
nor U751 (N_751,N_477,N_186);
or U752 (N_752,N_546,N_395);
or U753 (N_753,N_78,In_544);
nor U754 (N_754,N_572,N_357);
and U755 (N_755,N_321,N_244);
or U756 (N_756,In_338,In_587);
nand U757 (N_757,In_1063,N_419);
and U758 (N_758,In_1457,In_999);
nand U759 (N_759,In_635,N_315);
xnor U760 (N_760,In_1385,N_319);
xor U761 (N_761,N_592,In_1312);
or U762 (N_762,In_719,N_443);
or U763 (N_763,In_680,N_582);
xor U764 (N_764,In_499,N_490);
or U765 (N_765,In_518,In_570);
xnor U766 (N_766,In_1392,In_1179);
nor U767 (N_767,N_359,N_382);
xor U768 (N_768,N_331,In_868);
or U769 (N_769,N_58,N_339);
and U770 (N_770,In_883,N_306);
nand U771 (N_771,N_599,N_446);
and U772 (N_772,N_584,N_429);
or U773 (N_773,In_1122,In_1287);
xnor U774 (N_774,In_615,In_18);
nor U775 (N_775,In_621,N_312);
and U776 (N_776,In_33,N_500);
or U777 (N_777,In_1182,N_442);
or U778 (N_778,In_1060,N_428);
or U779 (N_779,In_670,N_193);
or U780 (N_780,N_144,In_623);
or U781 (N_781,In_528,N_518);
or U782 (N_782,In_691,In_14);
and U783 (N_783,N_531,N_94);
or U784 (N_784,In_1387,In_1237);
xor U785 (N_785,N_561,N_392);
xnor U786 (N_786,N_439,In_16);
nand U787 (N_787,In_668,In_1456);
nand U788 (N_788,N_578,In_502);
or U789 (N_789,In_895,In_752);
or U790 (N_790,In_661,N_380);
nor U791 (N_791,In_56,In_1097);
xor U792 (N_792,N_502,In_1391);
or U793 (N_793,N_138,In_727);
nand U794 (N_794,In_1415,In_262);
xor U795 (N_795,N_511,N_444);
and U796 (N_796,N_541,In_456);
or U797 (N_797,In_1398,N_407);
nor U798 (N_798,In_1045,N_185);
xnor U799 (N_799,In_1410,N_265);
or U800 (N_800,N_224,In_298);
and U801 (N_801,In_438,N_458);
or U802 (N_802,In_1491,In_656);
nand U803 (N_803,In_1159,N_271);
or U804 (N_804,N_28,N_397);
nand U805 (N_805,In_380,In_675);
or U806 (N_806,In_932,N_420);
or U807 (N_807,N_575,In_555);
xnor U808 (N_808,In_602,N_302);
and U809 (N_809,In_1331,In_581);
and U810 (N_810,In_769,N_377);
nand U811 (N_811,N_119,In_1455);
nand U812 (N_812,N_316,N_303);
xnor U813 (N_813,In_205,N_166);
and U814 (N_814,In_1013,In_873);
xor U815 (N_815,N_180,In_327);
nor U816 (N_816,N_183,In_1358);
xnor U817 (N_817,N_210,N_29);
nor U818 (N_818,In_845,N_538);
and U819 (N_819,In_140,In_288);
nand U820 (N_820,In_606,In_1239);
or U821 (N_821,In_906,In_1375);
nand U822 (N_822,N_551,N_432);
xnor U823 (N_823,N_230,In_1467);
or U824 (N_824,In_440,N_422);
nand U825 (N_825,In_6,In_964);
or U826 (N_826,In_387,In_1307);
xnor U827 (N_827,N_162,In_965);
xnor U828 (N_828,N_293,N_313);
nand U829 (N_829,N_348,In_567);
nand U830 (N_830,In_72,In_191);
nand U831 (N_831,In_228,N_326);
nor U832 (N_832,N_142,In_614);
and U833 (N_833,N_463,N_362);
and U834 (N_834,In_728,N_167);
or U835 (N_835,In_1031,N_371);
or U836 (N_836,In_1432,N_503);
nor U837 (N_837,In_741,N_513);
nor U838 (N_838,In_754,In_1289);
xnor U839 (N_839,In_1185,In_252);
xnor U840 (N_840,N_379,N_323);
xor U841 (N_841,N_344,N_114);
and U842 (N_842,N_398,In_333);
nor U843 (N_843,In_471,In_345);
and U844 (N_844,In_550,N_385);
and U845 (N_845,N_160,In_279);
nand U846 (N_846,In_344,In_681);
and U847 (N_847,N_155,N_237);
xor U848 (N_848,N_554,In_692);
nor U849 (N_849,N_296,In_1035);
nor U850 (N_850,In_330,N_596);
and U851 (N_851,N_368,In_537);
and U852 (N_852,N_406,In_1217);
nand U853 (N_853,In_1362,N_288);
xnor U854 (N_854,In_712,N_487);
xnor U855 (N_855,N_556,In_414);
or U856 (N_856,In_849,N_176);
nand U857 (N_857,In_430,N_197);
nor U858 (N_858,In_534,In_297);
xnor U859 (N_859,N_366,In_400);
xor U860 (N_860,In_346,In_1360);
and U861 (N_861,In_1393,N_214);
nor U862 (N_862,In_793,N_100);
xor U863 (N_863,In_9,N_577);
or U864 (N_864,In_1023,In_1399);
or U865 (N_865,In_751,N_455);
and U866 (N_866,N_251,In_358);
nand U867 (N_867,In_180,N_515);
nand U868 (N_868,N_184,N_355);
and U869 (N_869,N_558,In_975);
or U870 (N_870,N_542,N_153);
nor U871 (N_871,In_1234,N_127);
xor U872 (N_872,In_524,N_593);
nor U873 (N_873,In_827,N_559);
xnor U874 (N_874,In_348,N_595);
or U875 (N_875,N_298,N_571);
nor U876 (N_876,N_151,N_450);
or U877 (N_877,In_508,In_136);
or U878 (N_878,N_403,In_497);
and U879 (N_879,In_721,In_366);
nor U880 (N_880,N_67,N_400);
nor U881 (N_881,In_375,N_386);
and U882 (N_882,In_1366,In_1390);
xor U883 (N_883,N_387,In_1439);
or U884 (N_884,In_232,In_678);
xnor U885 (N_885,In_78,In_372);
or U886 (N_886,N_436,In_1173);
nand U887 (N_887,In_817,N_40);
xnor U888 (N_888,N_478,In_1207);
and U889 (N_889,N_568,In_777);
or U890 (N_890,N_402,N_457);
and U891 (N_891,N_512,N_140);
nor U892 (N_892,N_358,In_216);
nor U893 (N_893,N_168,N_528);
and U894 (N_894,N_384,N_465);
and U895 (N_895,N_383,N_178);
and U896 (N_896,In_984,N_532);
nor U897 (N_897,N_305,In_248);
xnor U898 (N_898,N_341,N_264);
nor U899 (N_899,In_409,N_566);
or U900 (N_900,N_767,N_761);
and U901 (N_901,In_778,N_731);
nand U902 (N_902,N_557,In_709);
xnor U903 (N_903,N_878,N_709);
nor U904 (N_904,N_718,In_776);
nand U905 (N_905,N_415,In_872);
nand U906 (N_906,In_630,N_812);
xor U907 (N_907,In_598,N_848);
nor U908 (N_908,N_884,N_610);
nand U909 (N_909,N_843,N_717);
and U910 (N_910,In_1379,N_898);
nor U911 (N_911,N_501,In_1478);
xnor U912 (N_912,N_701,N_169);
or U913 (N_913,In_13,N_866);
xor U914 (N_914,N_654,N_776);
nor U915 (N_915,N_771,N_839);
and U916 (N_916,N_735,N_838);
nand U917 (N_917,In_592,N_399);
xor U918 (N_918,In_520,In_1240);
nand U919 (N_919,N_346,In_626);
nand U920 (N_920,N_790,N_723);
nor U921 (N_921,N_719,N_885);
nand U922 (N_922,N_689,N_774);
nand U923 (N_923,N_590,N_886);
and U924 (N_924,N_525,N_562);
nor U925 (N_925,N_435,N_603);
and U926 (N_926,N_691,In_43);
nor U927 (N_927,N_608,N_850);
and U928 (N_928,N_768,N_698);
xor U929 (N_929,N_799,In_270);
xor U930 (N_930,N_636,N_869);
nand U931 (N_931,N_68,N_623);
nand U932 (N_932,N_780,N_684);
and U933 (N_933,N_859,N_97);
or U934 (N_934,N_232,In_714);
or U935 (N_935,N_641,N_860);
and U936 (N_936,N_656,N_389);
nor U937 (N_937,In_1373,N_711);
xor U938 (N_938,In_548,In_1041);
xnor U939 (N_939,N_785,N_891);
xnor U940 (N_940,N_796,N_521);
nor U941 (N_941,N_815,N_659);
nand U942 (N_942,N_849,In_1153);
or U943 (N_943,In_617,N_833);
or U944 (N_944,N_504,N_729);
nor U945 (N_945,N_652,N_784);
and U946 (N_946,In_1367,In_1425);
and U947 (N_947,In_1081,N_679);
or U948 (N_948,N_685,N_710);
and U949 (N_949,N_888,N_880);
nor U950 (N_950,In_52,N_825);
or U951 (N_951,N_198,In_818);
xor U952 (N_952,N_394,N_824);
xor U953 (N_953,In_165,N_635);
nand U954 (N_954,N_514,In_427);
or U955 (N_955,N_272,N_712);
xnor U956 (N_956,N_855,N_650);
or U957 (N_957,N_811,N_822);
nor U958 (N_958,N_736,N_818);
nor U959 (N_959,N_494,N_876);
and U960 (N_960,In_1184,N_788);
nor U961 (N_961,N_817,N_890);
and U962 (N_962,N_857,N_791);
xnor U963 (N_963,N_831,In_1308);
xnor U964 (N_964,N_360,N_686);
nand U965 (N_965,N_533,N_662);
and U966 (N_966,N_621,N_259);
xor U967 (N_967,N_536,N_170);
or U968 (N_968,N_658,N_696);
and U969 (N_969,N_674,N_535);
and U970 (N_970,In_417,N_417);
nor U971 (N_971,N_680,In_389);
nor U972 (N_972,N_520,N_672);
nand U973 (N_973,N_87,N_121);
xor U974 (N_974,N_793,N_675);
and U975 (N_975,N_327,N_612);
nand U976 (N_976,In_877,N_589);
xnor U977 (N_977,N_451,N_236);
nand U978 (N_978,N_498,N_580);
xor U979 (N_979,N_690,N_865);
or U980 (N_980,N_485,N_687);
xor U981 (N_981,N_547,N_345);
nor U982 (N_982,In_919,N_573);
nand U983 (N_983,N_832,N_628);
and U984 (N_984,N_278,In_557);
or U985 (N_985,In_1341,In_249);
and U986 (N_986,In_156,N_657);
nor U987 (N_987,N_17,N_522);
or U988 (N_988,In_1259,N_75);
or U989 (N_989,N_300,N_304);
or U990 (N_990,N_560,N_671);
and U991 (N_991,In_1150,N_668);
xnor U992 (N_992,N_797,N_367);
nand U993 (N_993,N_751,N_204);
nor U994 (N_994,N_755,N_425);
or U995 (N_995,N_829,N_651);
or U996 (N_996,N_116,N_550);
xor U997 (N_997,N_480,N_856);
nor U998 (N_998,N_601,N_769);
nand U999 (N_999,N_744,N_309);
or U1000 (N_1000,N_682,N_499);
nand U1001 (N_1001,N_845,In_720);
nand U1002 (N_1002,N_827,N_782);
xnor U1003 (N_1003,In_459,In_1094);
xor U1004 (N_1004,N_764,N_507);
and U1005 (N_1005,N_646,N_552);
nor U1006 (N_1006,In_801,In_1099);
xnor U1007 (N_1007,N_591,N_725);
or U1008 (N_1008,N_424,N_882);
and U1009 (N_1009,N_242,N_617);
and U1010 (N_1010,N_874,In_498);
or U1011 (N_1011,N_720,N_851);
or U1012 (N_1012,N_697,N_661);
nand U1013 (N_1013,N_821,N_816);
and U1014 (N_1014,N_677,N_411);
nor U1015 (N_1015,N_634,N_343);
or U1016 (N_1016,N_683,N_694);
or U1017 (N_1017,N_605,N_631);
xor U1018 (N_1018,N_517,In_413);
or U1019 (N_1019,N_642,N_622);
nand U1020 (N_1020,N_495,N_802);
nor U1021 (N_1021,N_190,N_391);
and U1022 (N_1022,N_630,In_561);
nor U1023 (N_1023,N_196,N_633);
nand U1024 (N_1024,N_748,N_778);
nor U1025 (N_1025,N_640,In_521);
or U1026 (N_1026,In_1221,N_11);
and U1027 (N_1027,N_529,N_732);
nand U1028 (N_1028,In_1144,N_150);
nand U1029 (N_1029,N_648,N_421);
and U1030 (N_1030,N_862,N_320);
nand U1031 (N_1031,N_440,In_1466);
nand U1032 (N_1032,In_729,In_815);
nand U1033 (N_1033,N_638,N_607);
xnor U1034 (N_1034,In_1487,N_759);
or U1035 (N_1035,In_1271,In_1205);
nand U1036 (N_1036,In_139,N_336);
nor U1037 (N_1037,N_830,N_472);
or U1038 (N_1038,N_749,In_613);
nor U1039 (N_1039,In_1286,In_1248);
or U1040 (N_1040,N_223,N_738);
nand U1041 (N_1041,N_706,In_448);
nor U1042 (N_1042,N_609,In_1359);
nand U1043 (N_1043,N_864,In_1145);
nand U1044 (N_1044,N_669,N_693);
xor U1045 (N_1045,In_1449,N_655);
or U1046 (N_1046,N_374,In_68);
and U1047 (N_1047,In_589,N_333);
or U1048 (N_1048,N_632,N_743);
or U1049 (N_1049,In_990,N_332);
nand U1050 (N_1050,In_85,In_1371);
and U1051 (N_1051,N_750,N_846);
nand U1052 (N_1052,In_662,In_952);
xnor U1053 (N_1053,In_928,N_762);
nand U1054 (N_1054,In_41,In_73);
nor U1055 (N_1055,N_813,N_234);
or U1056 (N_1056,N_820,In_655);
xnor U1057 (N_1057,In_862,N_647);
nor U1058 (N_1058,In_423,N_375);
xnor U1059 (N_1059,N_493,N_730);
nand U1060 (N_1060,N_760,N_405);
or U1061 (N_1061,N_809,N_318);
xor U1062 (N_1062,N_840,In_453);
nand U1063 (N_1063,In_940,N_800);
and U1064 (N_1064,N_614,N_806);
xnor U1065 (N_1065,In_4,N_335);
xnor U1066 (N_1066,In_132,N_604);
nand U1067 (N_1067,N_863,N_896);
nor U1068 (N_1068,N_756,In_1316);
nor U1069 (N_1069,N_624,N_787);
or U1070 (N_1070,N_172,N_754);
xnor U1071 (N_1071,In_1085,In_622);
or U1072 (N_1072,N_274,In_991);
or U1073 (N_1073,N_870,N_322);
and U1074 (N_1074,In_809,N_667);
xor U1075 (N_1075,N_354,In_687);
or U1076 (N_1076,N_716,N_826);
xor U1077 (N_1077,N_847,N_783);
nand U1078 (N_1078,N_798,In_1299);
xor U1079 (N_1079,N_739,N_781);
xnor U1080 (N_1080,N_431,In_154);
xor U1081 (N_1081,N_342,N_721);
nand U1082 (N_1082,N_328,N_792);
and U1083 (N_1083,In_455,N_707);
xnor U1084 (N_1084,N_873,N_861);
nand U1085 (N_1085,N_14,N_852);
and U1086 (N_1086,In_222,N_700);
xor U1087 (N_1087,N_666,N_618);
nor U1088 (N_1088,In_1223,N_834);
nand U1089 (N_1089,In_1100,N_616);
and U1090 (N_1090,In_1464,N_889);
and U1091 (N_1091,N_408,N_469);
and U1092 (N_1092,N_492,N_479);
xor U1093 (N_1093,N_47,In_865);
or U1094 (N_1094,In_1402,In_446);
and U1095 (N_1095,N_49,N_606);
nor U1096 (N_1096,N_715,In_902);
and U1097 (N_1097,In_1283,In_215);
and U1098 (N_1098,In_797,N_837);
or U1099 (N_1099,N_629,In_134);
and U1100 (N_1100,N_804,N_814);
nand U1101 (N_1101,In_1334,N_673);
or U1102 (N_1102,In_356,N_726);
and U1103 (N_1103,N_219,N_681);
nor U1104 (N_1104,N_625,In_58);
and U1105 (N_1105,In_77,N_789);
xor U1106 (N_1106,N_83,N_548);
xnor U1107 (N_1107,In_1064,In_268);
nor U1108 (N_1108,N_611,N_351);
nand U1109 (N_1109,N_828,In_69);
or U1110 (N_1110,N_619,N_246);
nor U1111 (N_1111,N_626,N_461);
nor U1112 (N_1112,N_895,N_260);
or U1113 (N_1113,N_705,N_714);
nor U1114 (N_1114,N_713,N_875);
nor U1115 (N_1115,N_615,N_670);
or U1116 (N_1116,N_703,In_397);
and U1117 (N_1117,N_737,In_193);
nor U1118 (N_1118,N_899,In_231);
xnor U1119 (N_1119,N_844,In_764);
or U1120 (N_1120,N_356,N_742);
or U1121 (N_1121,N_757,N_678);
xnor U1122 (N_1122,In_1009,N_349);
nand U1123 (N_1123,N_639,N_897);
nor U1124 (N_1124,In_84,N_872);
xnor U1125 (N_1125,N_835,In_963);
nand U1126 (N_1126,N_724,N_777);
xnor U1127 (N_1127,N_688,In_1209);
and U1128 (N_1128,N_564,N_613);
and U1129 (N_1129,In_717,In_432);
xor U1130 (N_1130,N_766,In_178);
nand U1131 (N_1131,N_881,In_1303);
xnor U1132 (N_1132,In_800,N_775);
xor U1133 (N_1133,N_519,In_1260);
xor U1134 (N_1134,In_1199,N_858);
xnor U1135 (N_1135,N_702,N_35);
and U1136 (N_1136,N_600,N_727);
or U1137 (N_1137,In_322,N_734);
nand U1138 (N_1138,N_795,N_803);
nor U1139 (N_1139,In_1141,N_38);
nor U1140 (N_1140,N_665,N_314);
nand U1141 (N_1141,N_765,N_722);
or U1142 (N_1142,N_644,N_823);
and U1143 (N_1143,N_449,N_753);
and U1144 (N_1144,In_458,N_413);
nor U1145 (N_1145,N_434,N_794);
xnor U1146 (N_1146,N_401,In_129);
and U1147 (N_1147,N_570,In_468);
xor U1148 (N_1148,N_433,In_265);
and U1149 (N_1149,N_801,N_317);
nand U1150 (N_1150,N_773,N_468);
nand U1151 (N_1151,In_805,N_221);
and U1152 (N_1152,In_1114,N_877);
and U1153 (N_1153,N_745,In_396);
nand U1154 (N_1154,N_649,N_620);
nor U1155 (N_1155,In_1233,N_645);
xor U1156 (N_1156,N_497,N_708);
or U1157 (N_1157,In_1216,N_462);
and U1158 (N_1158,N_660,N_695);
and U1159 (N_1159,N_893,N_627);
nor U1160 (N_1160,In_674,N_836);
xnor U1161 (N_1161,N_894,N_779);
and U1162 (N_1162,N_103,In_211);
xnor U1163 (N_1163,N_752,In_449);
or U1164 (N_1164,N_786,N_841);
or U1165 (N_1165,In_480,In_1142);
nor U1166 (N_1166,N_805,In_1258);
nand U1167 (N_1167,N_747,N_174);
nand U1168 (N_1168,N_853,N_704);
and U1169 (N_1169,N_653,N_868);
or U1170 (N_1170,N_588,N_664);
nand U1171 (N_1171,N_842,In_485);
nor U1172 (N_1172,N_637,N_699);
xor U1173 (N_1173,N_740,In_1461);
xnor U1174 (N_1174,N_135,In_286);
nand U1175 (N_1175,In_848,In_411);
or U1176 (N_1176,N_474,N_807);
and U1177 (N_1177,N_770,N_247);
or U1178 (N_1178,In_291,In_953);
xnor U1179 (N_1179,N_871,N_565);
or U1180 (N_1180,In_328,N_883);
nand U1181 (N_1181,N_741,In_1180);
nand U1182 (N_1182,N_581,In_527);
or U1183 (N_1183,N_758,N_456);
and U1184 (N_1184,N_82,In_1068);
or U1185 (N_1185,N_819,N_728);
xor U1186 (N_1186,In_1065,N_643);
nor U1187 (N_1187,N_539,N_854);
and U1188 (N_1188,N_887,N_763);
xnor U1189 (N_1189,N_892,N_129);
nand U1190 (N_1190,N_772,N_586);
xor U1191 (N_1191,In_525,In_1024);
and U1192 (N_1192,N_663,N_733);
xnor U1193 (N_1193,N_808,N_867);
and U1194 (N_1194,In_1474,N_105);
nand U1195 (N_1195,N_692,N_3);
xor U1196 (N_1196,N_879,In_310);
xnor U1197 (N_1197,In_756,N_746);
and U1198 (N_1198,N_810,N_602);
and U1199 (N_1199,In_857,N_676);
nor U1200 (N_1200,N_1030,N_1106);
nor U1201 (N_1201,N_1125,N_1036);
xnor U1202 (N_1202,N_1105,N_1063);
and U1203 (N_1203,N_1012,N_1195);
and U1204 (N_1204,N_1042,N_1190);
nand U1205 (N_1205,N_955,N_998);
or U1206 (N_1206,N_1034,N_1184);
nor U1207 (N_1207,N_991,N_1076);
nand U1208 (N_1208,N_1019,N_1109);
nor U1209 (N_1209,N_1081,N_1112);
or U1210 (N_1210,N_1182,N_1183);
nor U1211 (N_1211,N_1122,N_951);
or U1212 (N_1212,N_942,N_1000);
and U1213 (N_1213,N_1194,N_956);
xor U1214 (N_1214,N_1044,N_1160);
nor U1215 (N_1215,N_968,N_1010);
xor U1216 (N_1216,N_1186,N_1046);
xor U1217 (N_1217,N_961,N_1196);
xnor U1218 (N_1218,N_1007,N_1021);
nand U1219 (N_1219,N_1116,N_1004);
nor U1220 (N_1220,N_949,N_1079);
xor U1221 (N_1221,N_1199,N_1126);
and U1222 (N_1222,N_1101,N_1165);
xor U1223 (N_1223,N_935,N_1005);
nor U1224 (N_1224,N_1049,N_1098);
or U1225 (N_1225,N_916,N_1048);
xor U1226 (N_1226,N_1020,N_946);
xnor U1227 (N_1227,N_1108,N_1028);
nor U1228 (N_1228,N_1060,N_939);
nand U1229 (N_1229,N_1135,N_1100);
and U1230 (N_1230,N_1128,N_959);
and U1231 (N_1231,N_958,N_1158);
nor U1232 (N_1232,N_982,N_1003);
and U1233 (N_1233,N_1023,N_990);
or U1234 (N_1234,N_1163,N_967);
and U1235 (N_1235,N_1144,N_1154);
xnor U1236 (N_1236,N_999,N_1185);
or U1237 (N_1237,N_1155,N_997);
and U1238 (N_1238,N_953,N_1059);
and U1239 (N_1239,N_1124,N_902);
or U1240 (N_1240,N_952,N_1051);
nand U1241 (N_1241,N_1031,N_1169);
nor U1242 (N_1242,N_930,N_1131);
nor U1243 (N_1243,N_954,N_986);
xor U1244 (N_1244,N_1107,N_1039);
nor U1245 (N_1245,N_912,N_1167);
xor U1246 (N_1246,N_1172,N_1159);
or U1247 (N_1247,N_1179,N_1175);
and U1248 (N_1248,N_941,N_1157);
or U1249 (N_1249,N_1080,N_1070);
xnor U1250 (N_1250,N_964,N_1002);
and U1251 (N_1251,N_985,N_957);
nand U1252 (N_1252,N_1087,N_1166);
nand U1253 (N_1253,N_1022,N_915);
or U1254 (N_1254,N_1127,N_1174);
nor U1255 (N_1255,N_1095,N_1145);
nor U1256 (N_1256,N_1191,N_1103);
or U1257 (N_1257,N_987,N_1027);
xnor U1258 (N_1258,N_1180,N_975);
nand U1259 (N_1259,N_1143,N_1008);
xor U1260 (N_1260,N_1173,N_932);
xnor U1261 (N_1261,N_1198,N_1137);
xor U1262 (N_1262,N_979,N_1114);
xor U1263 (N_1263,N_937,N_1168);
nor U1264 (N_1264,N_1018,N_929);
nand U1265 (N_1265,N_1140,N_1024);
and U1266 (N_1266,N_1142,N_931);
or U1267 (N_1267,N_1016,N_1147);
nor U1268 (N_1268,N_1001,N_947);
nand U1269 (N_1269,N_1110,N_1193);
nand U1270 (N_1270,N_973,N_984);
nand U1271 (N_1271,N_1075,N_948);
and U1272 (N_1272,N_1141,N_904);
or U1273 (N_1273,N_983,N_1134);
xor U1274 (N_1274,N_1009,N_1015);
and U1275 (N_1275,N_903,N_906);
nor U1276 (N_1276,N_992,N_1130);
nor U1277 (N_1277,N_1156,N_1078);
and U1278 (N_1278,N_1071,N_1099);
or U1279 (N_1279,N_1104,N_1006);
xor U1280 (N_1280,N_1111,N_1136);
nand U1281 (N_1281,N_1052,N_1097);
and U1282 (N_1282,N_1177,N_981);
or U1283 (N_1283,N_962,N_1187);
xnor U1284 (N_1284,N_1088,N_1056);
nand U1285 (N_1285,N_921,N_993);
xor U1286 (N_1286,N_922,N_1153);
or U1287 (N_1287,N_944,N_1055);
xor U1288 (N_1288,N_1032,N_1038);
xor U1289 (N_1289,N_1045,N_908);
nand U1290 (N_1290,N_1133,N_918);
or U1291 (N_1291,N_1058,N_960);
or U1292 (N_1292,N_1050,N_1014);
xor U1293 (N_1293,N_1066,N_1162);
or U1294 (N_1294,N_1054,N_927);
or U1295 (N_1295,N_928,N_1151);
and U1296 (N_1296,N_920,N_965);
or U1297 (N_1297,N_1091,N_969);
nor U1298 (N_1298,N_934,N_1035);
or U1299 (N_1299,N_940,N_910);
nor U1300 (N_1300,N_923,N_971);
xnor U1301 (N_1301,N_1171,N_1119);
or U1302 (N_1302,N_1096,N_1040);
and U1303 (N_1303,N_1065,N_1084);
nor U1304 (N_1304,N_1094,N_1026);
nor U1305 (N_1305,N_1069,N_1149);
nand U1306 (N_1306,N_1089,N_989);
or U1307 (N_1307,N_1073,N_1170);
xor U1308 (N_1308,N_1017,N_1057);
nor U1309 (N_1309,N_963,N_911);
xnor U1310 (N_1310,N_917,N_1102);
or U1311 (N_1311,N_1132,N_978);
nor U1312 (N_1312,N_1164,N_996);
nand U1313 (N_1313,N_1189,N_972);
nor U1314 (N_1314,N_943,N_1090);
and U1315 (N_1315,N_988,N_1139);
or U1316 (N_1316,N_1061,N_1152);
xor U1317 (N_1317,N_1037,N_1138);
nor U1318 (N_1318,N_1118,N_1025);
nand U1319 (N_1319,N_1148,N_977);
or U1320 (N_1320,N_1146,N_938);
nand U1321 (N_1321,N_970,N_950);
and U1322 (N_1322,N_900,N_1161);
xnor U1323 (N_1323,N_1178,N_1083);
or U1324 (N_1324,N_1011,N_1033);
xnor U1325 (N_1325,N_1197,N_980);
or U1326 (N_1326,N_1117,N_1192);
or U1327 (N_1327,N_1082,N_933);
and U1328 (N_1328,N_1043,N_1067);
nand U1329 (N_1329,N_1123,N_1086);
nand U1330 (N_1330,N_1029,N_1068);
nand U1331 (N_1331,N_1062,N_1064);
xnor U1332 (N_1332,N_1121,N_1113);
nor U1333 (N_1333,N_1129,N_1047);
and U1334 (N_1334,N_966,N_1176);
xnor U1335 (N_1335,N_1093,N_974);
xor U1336 (N_1336,N_1077,N_925);
nor U1337 (N_1337,N_907,N_1053);
or U1338 (N_1338,N_926,N_905);
nor U1339 (N_1339,N_1115,N_1085);
xor U1340 (N_1340,N_936,N_1074);
xor U1341 (N_1341,N_1092,N_1188);
xnor U1342 (N_1342,N_913,N_914);
or U1343 (N_1343,N_1041,N_919);
xor U1344 (N_1344,N_909,N_1072);
nor U1345 (N_1345,N_901,N_994);
and U1346 (N_1346,N_1181,N_1120);
xnor U1347 (N_1347,N_976,N_1150);
nor U1348 (N_1348,N_1013,N_945);
nor U1349 (N_1349,N_995,N_924);
and U1350 (N_1350,N_943,N_973);
nand U1351 (N_1351,N_1197,N_1150);
xor U1352 (N_1352,N_977,N_1000);
xnor U1353 (N_1353,N_1135,N_965);
nor U1354 (N_1354,N_951,N_1100);
or U1355 (N_1355,N_1157,N_1169);
or U1356 (N_1356,N_992,N_1159);
nor U1357 (N_1357,N_1053,N_1120);
nand U1358 (N_1358,N_1072,N_939);
nor U1359 (N_1359,N_1149,N_1027);
nor U1360 (N_1360,N_1197,N_1058);
nor U1361 (N_1361,N_1078,N_1013);
nand U1362 (N_1362,N_1065,N_932);
xnor U1363 (N_1363,N_1129,N_933);
and U1364 (N_1364,N_1073,N_1079);
or U1365 (N_1365,N_1090,N_992);
or U1366 (N_1366,N_904,N_942);
or U1367 (N_1367,N_1089,N_1031);
or U1368 (N_1368,N_1012,N_1181);
xnor U1369 (N_1369,N_940,N_986);
nor U1370 (N_1370,N_986,N_1115);
xnor U1371 (N_1371,N_1027,N_1157);
and U1372 (N_1372,N_986,N_1065);
nor U1373 (N_1373,N_1197,N_983);
nor U1374 (N_1374,N_1185,N_1142);
nand U1375 (N_1375,N_1038,N_1107);
nand U1376 (N_1376,N_914,N_1004);
nor U1377 (N_1377,N_1095,N_1093);
or U1378 (N_1378,N_1128,N_1057);
or U1379 (N_1379,N_1129,N_981);
xnor U1380 (N_1380,N_1181,N_1103);
nand U1381 (N_1381,N_1186,N_1179);
and U1382 (N_1382,N_982,N_1063);
and U1383 (N_1383,N_1099,N_1130);
nor U1384 (N_1384,N_1014,N_953);
or U1385 (N_1385,N_1129,N_1087);
xor U1386 (N_1386,N_1065,N_1122);
and U1387 (N_1387,N_1007,N_1054);
nor U1388 (N_1388,N_1135,N_1080);
nor U1389 (N_1389,N_1162,N_1169);
nor U1390 (N_1390,N_1026,N_1193);
nand U1391 (N_1391,N_969,N_966);
nand U1392 (N_1392,N_1109,N_1186);
nor U1393 (N_1393,N_1051,N_1178);
and U1394 (N_1394,N_926,N_1166);
or U1395 (N_1395,N_959,N_943);
and U1396 (N_1396,N_1112,N_1141);
xor U1397 (N_1397,N_935,N_901);
xor U1398 (N_1398,N_948,N_1187);
or U1399 (N_1399,N_1136,N_1140);
nand U1400 (N_1400,N_992,N_1118);
xnor U1401 (N_1401,N_960,N_1127);
xnor U1402 (N_1402,N_1072,N_1000);
nor U1403 (N_1403,N_1154,N_1004);
nor U1404 (N_1404,N_1032,N_1116);
nand U1405 (N_1405,N_996,N_1128);
and U1406 (N_1406,N_1124,N_1010);
nor U1407 (N_1407,N_1142,N_1163);
xnor U1408 (N_1408,N_1150,N_1092);
nand U1409 (N_1409,N_955,N_906);
nand U1410 (N_1410,N_941,N_991);
or U1411 (N_1411,N_1197,N_1063);
nand U1412 (N_1412,N_1172,N_1083);
and U1413 (N_1413,N_932,N_1056);
or U1414 (N_1414,N_1163,N_955);
or U1415 (N_1415,N_920,N_1032);
and U1416 (N_1416,N_1144,N_1115);
nor U1417 (N_1417,N_987,N_1113);
nand U1418 (N_1418,N_1071,N_1035);
and U1419 (N_1419,N_986,N_1191);
and U1420 (N_1420,N_992,N_1036);
and U1421 (N_1421,N_1188,N_1161);
or U1422 (N_1422,N_906,N_915);
nor U1423 (N_1423,N_1078,N_1007);
nand U1424 (N_1424,N_925,N_1170);
nor U1425 (N_1425,N_1193,N_1143);
and U1426 (N_1426,N_1134,N_1024);
nand U1427 (N_1427,N_1063,N_1186);
nand U1428 (N_1428,N_1046,N_1076);
xnor U1429 (N_1429,N_1070,N_971);
nand U1430 (N_1430,N_1153,N_986);
nand U1431 (N_1431,N_954,N_939);
nor U1432 (N_1432,N_944,N_991);
and U1433 (N_1433,N_984,N_924);
xor U1434 (N_1434,N_930,N_1010);
xor U1435 (N_1435,N_1136,N_1068);
xnor U1436 (N_1436,N_1059,N_982);
and U1437 (N_1437,N_923,N_1198);
nor U1438 (N_1438,N_1074,N_904);
nor U1439 (N_1439,N_959,N_1098);
and U1440 (N_1440,N_1099,N_984);
xor U1441 (N_1441,N_1061,N_1160);
nor U1442 (N_1442,N_990,N_1155);
and U1443 (N_1443,N_1145,N_1155);
and U1444 (N_1444,N_1101,N_1086);
or U1445 (N_1445,N_938,N_1019);
xor U1446 (N_1446,N_1022,N_1010);
nand U1447 (N_1447,N_1046,N_920);
or U1448 (N_1448,N_959,N_1094);
nor U1449 (N_1449,N_1138,N_1164);
nand U1450 (N_1450,N_1145,N_970);
or U1451 (N_1451,N_938,N_1000);
nor U1452 (N_1452,N_1002,N_1184);
nor U1453 (N_1453,N_1092,N_1156);
nor U1454 (N_1454,N_1051,N_934);
xnor U1455 (N_1455,N_1165,N_1075);
xor U1456 (N_1456,N_1172,N_1154);
nor U1457 (N_1457,N_1056,N_921);
or U1458 (N_1458,N_1195,N_1161);
or U1459 (N_1459,N_1131,N_1088);
nor U1460 (N_1460,N_1089,N_1166);
and U1461 (N_1461,N_983,N_1030);
nand U1462 (N_1462,N_996,N_1127);
or U1463 (N_1463,N_972,N_1157);
xnor U1464 (N_1464,N_959,N_966);
nor U1465 (N_1465,N_934,N_986);
nor U1466 (N_1466,N_1010,N_1043);
nand U1467 (N_1467,N_1138,N_917);
nor U1468 (N_1468,N_1106,N_982);
or U1469 (N_1469,N_1100,N_1011);
nand U1470 (N_1470,N_945,N_1014);
nor U1471 (N_1471,N_1004,N_1131);
and U1472 (N_1472,N_1021,N_901);
nor U1473 (N_1473,N_937,N_1094);
and U1474 (N_1474,N_990,N_1138);
nor U1475 (N_1475,N_960,N_996);
xor U1476 (N_1476,N_919,N_1076);
or U1477 (N_1477,N_1024,N_1169);
nor U1478 (N_1478,N_1076,N_944);
and U1479 (N_1479,N_1148,N_1107);
nand U1480 (N_1480,N_1072,N_1110);
or U1481 (N_1481,N_999,N_1128);
xor U1482 (N_1482,N_1190,N_940);
and U1483 (N_1483,N_963,N_925);
or U1484 (N_1484,N_1002,N_942);
xor U1485 (N_1485,N_1180,N_1184);
or U1486 (N_1486,N_1153,N_1183);
and U1487 (N_1487,N_1103,N_979);
nor U1488 (N_1488,N_1126,N_1043);
or U1489 (N_1489,N_959,N_910);
or U1490 (N_1490,N_1197,N_1140);
nand U1491 (N_1491,N_1157,N_929);
nand U1492 (N_1492,N_1042,N_1079);
nor U1493 (N_1493,N_901,N_1090);
and U1494 (N_1494,N_985,N_969);
or U1495 (N_1495,N_1054,N_1186);
nand U1496 (N_1496,N_1193,N_1156);
nor U1497 (N_1497,N_1120,N_1132);
or U1498 (N_1498,N_913,N_1085);
or U1499 (N_1499,N_1094,N_1174);
and U1500 (N_1500,N_1315,N_1319);
and U1501 (N_1501,N_1239,N_1408);
xor U1502 (N_1502,N_1230,N_1255);
and U1503 (N_1503,N_1286,N_1298);
nand U1504 (N_1504,N_1451,N_1450);
and U1505 (N_1505,N_1378,N_1256);
nand U1506 (N_1506,N_1453,N_1471);
nor U1507 (N_1507,N_1497,N_1200);
and U1508 (N_1508,N_1322,N_1262);
xnor U1509 (N_1509,N_1488,N_1339);
xnor U1510 (N_1510,N_1351,N_1251);
nor U1511 (N_1511,N_1456,N_1430);
or U1512 (N_1512,N_1482,N_1336);
xor U1513 (N_1513,N_1473,N_1463);
and U1514 (N_1514,N_1287,N_1429);
or U1515 (N_1515,N_1310,N_1417);
or U1516 (N_1516,N_1387,N_1419);
nor U1517 (N_1517,N_1377,N_1445);
or U1518 (N_1518,N_1284,N_1457);
and U1519 (N_1519,N_1276,N_1323);
nand U1520 (N_1520,N_1369,N_1206);
xor U1521 (N_1521,N_1259,N_1309);
or U1522 (N_1522,N_1333,N_1345);
or U1523 (N_1523,N_1263,N_1289);
nor U1524 (N_1524,N_1320,N_1335);
and U1525 (N_1525,N_1352,N_1253);
and U1526 (N_1526,N_1212,N_1228);
nor U1527 (N_1527,N_1402,N_1381);
nor U1528 (N_1528,N_1407,N_1208);
nand U1529 (N_1529,N_1346,N_1413);
and U1530 (N_1530,N_1411,N_1410);
or U1531 (N_1531,N_1350,N_1404);
xor U1532 (N_1532,N_1278,N_1330);
nor U1533 (N_1533,N_1421,N_1397);
or U1534 (N_1534,N_1476,N_1422);
xor U1535 (N_1535,N_1481,N_1388);
and U1536 (N_1536,N_1393,N_1271);
nand U1537 (N_1537,N_1232,N_1210);
nor U1538 (N_1538,N_1275,N_1426);
xor U1539 (N_1539,N_1223,N_1297);
or U1540 (N_1540,N_1358,N_1440);
or U1541 (N_1541,N_1483,N_1291);
or U1542 (N_1542,N_1341,N_1443);
nand U1543 (N_1543,N_1209,N_1279);
and U1544 (N_1544,N_1204,N_1398);
nor U1545 (N_1545,N_1329,N_1317);
xor U1546 (N_1546,N_1401,N_1405);
nand U1547 (N_1547,N_1406,N_1460);
and U1548 (N_1548,N_1360,N_1418);
xor U1549 (N_1549,N_1490,N_1416);
nor U1550 (N_1550,N_1318,N_1334);
xnor U1551 (N_1551,N_1288,N_1226);
or U1552 (N_1552,N_1436,N_1229);
nand U1553 (N_1553,N_1498,N_1285);
xnor U1554 (N_1554,N_1234,N_1280);
xnor U1555 (N_1555,N_1296,N_1383);
nand U1556 (N_1556,N_1475,N_1477);
and U1557 (N_1557,N_1273,N_1268);
nand U1558 (N_1558,N_1241,N_1431);
or U1559 (N_1559,N_1356,N_1294);
and U1560 (N_1560,N_1363,N_1269);
and U1561 (N_1561,N_1361,N_1220);
and U1562 (N_1562,N_1292,N_1302);
or U1563 (N_1563,N_1313,N_1207);
nor U1564 (N_1564,N_1264,N_1290);
xnor U1565 (N_1565,N_1427,N_1458);
or U1566 (N_1566,N_1392,N_1247);
nor U1567 (N_1567,N_1424,N_1432);
or U1568 (N_1568,N_1267,N_1308);
nor U1569 (N_1569,N_1362,N_1250);
or U1570 (N_1570,N_1214,N_1277);
nor U1571 (N_1571,N_1217,N_1487);
xor U1572 (N_1572,N_1303,N_1466);
and U1573 (N_1573,N_1367,N_1373);
and U1574 (N_1574,N_1328,N_1400);
and U1575 (N_1575,N_1492,N_1257);
xor U1576 (N_1576,N_1371,N_1359);
nor U1577 (N_1577,N_1365,N_1441);
xnor U1578 (N_1578,N_1237,N_1394);
xnor U1579 (N_1579,N_1258,N_1435);
or U1580 (N_1580,N_1412,N_1254);
xor U1581 (N_1581,N_1243,N_1382);
nand U1582 (N_1582,N_1357,N_1312);
nor U1583 (N_1583,N_1470,N_1205);
and U1584 (N_1584,N_1233,N_1274);
and U1585 (N_1585,N_1238,N_1353);
or U1586 (N_1586,N_1438,N_1465);
or U1587 (N_1587,N_1225,N_1235);
nor U1588 (N_1588,N_1467,N_1366);
nand U1589 (N_1589,N_1478,N_1252);
nand U1590 (N_1590,N_1433,N_1464);
xnor U1591 (N_1591,N_1236,N_1215);
xor U1592 (N_1592,N_1386,N_1491);
nand U1593 (N_1593,N_1316,N_1244);
nand U1594 (N_1594,N_1472,N_1375);
nor U1595 (N_1595,N_1265,N_1203);
and U1596 (N_1596,N_1389,N_1272);
xor U1597 (N_1597,N_1231,N_1266);
nand U1598 (N_1598,N_1454,N_1403);
nand U1599 (N_1599,N_1240,N_1349);
nand U1600 (N_1600,N_1282,N_1423);
xnor U1601 (N_1601,N_1299,N_1372);
nor U1602 (N_1602,N_1213,N_1489);
and U1603 (N_1603,N_1376,N_1260);
or U1604 (N_1604,N_1459,N_1305);
and U1605 (N_1605,N_1224,N_1364);
xnor U1606 (N_1606,N_1304,N_1496);
nand U1607 (N_1607,N_1379,N_1347);
nor U1608 (N_1608,N_1409,N_1380);
xor U1609 (N_1609,N_1300,N_1449);
or U1610 (N_1610,N_1338,N_1370);
nor U1611 (N_1611,N_1211,N_1307);
nor U1612 (N_1612,N_1479,N_1219);
nor U1613 (N_1613,N_1425,N_1499);
and U1614 (N_1614,N_1484,N_1332);
xor U1615 (N_1615,N_1248,N_1348);
nor U1616 (N_1616,N_1202,N_1395);
nor U1617 (N_1617,N_1428,N_1444);
nor U1618 (N_1618,N_1246,N_1494);
nor U1619 (N_1619,N_1415,N_1455);
xnor U1620 (N_1620,N_1437,N_1218);
xnor U1621 (N_1621,N_1399,N_1469);
nor U1622 (N_1622,N_1355,N_1324);
nor U1623 (N_1623,N_1495,N_1222);
xor U1624 (N_1624,N_1325,N_1314);
nor U1625 (N_1625,N_1396,N_1448);
or U1626 (N_1626,N_1327,N_1452);
or U1627 (N_1627,N_1340,N_1242);
nand U1628 (N_1628,N_1485,N_1227);
nor U1629 (N_1629,N_1344,N_1439);
nor U1630 (N_1630,N_1447,N_1391);
or U1631 (N_1631,N_1337,N_1221);
and U1632 (N_1632,N_1368,N_1249);
nand U1633 (N_1633,N_1321,N_1343);
or U1634 (N_1634,N_1311,N_1281);
nand U1635 (N_1635,N_1293,N_1216);
nand U1636 (N_1636,N_1480,N_1326);
xor U1637 (N_1637,N_1374,N_1434);
nor U1638 (N_1638,N_1354,N_1442);
xnor U1639 (N_1639,N_1462,N_1493);
or U1640 (N_1640,N_1384,N_1261);
and U1641 (N_1641,N_1461,N_1342);
nand U1642 (N_1642,N_1385,N_1468);
nand U1643 (N_1643,N_1474,N_1420);
xnor U1644 (N_1644,N_1331,N_1414);
or U1645 (N_1645,N_1283,N_1486);
nor U1646 (N_1646,N_1270,N_1390);
or U1647 (N_1647,N_1306,N_1446);
xnor U1648 (N_1648,N_1301,N_1295);
nand U1649 (N_1649,N_1201,N_1245);
xnor U1650 (N_1650,N_1362,N_1423);
nand U1651 (N_1651,N_1263,N_1243);
or U1652 (N_1652,N_1404,N_1383);
nor U1653 (N_1653,N_1256,N_1274);
and U1654 (N_1654,N_1475,N_1210);
nor U1655 (N_1655,N_1288,N_1441);
nand U1656 (N_1656,N_1409,N_1439);
or U1657 (N_1657,N_1225,N_1214);
nand U1658 (N_1658,N_1211,N_1312);
nand U1659 (N_1659,N_1286,N_1391);
nor U1660 (N_1660,N_1465,N_1422);
nor U1661 (N_1661,N_1235,N_1461);
and U1662 (N_1662,N_1296,N_1235);
or U1663 (N_1663,N_1258,N_1394);
or U1664 (N_1664,N_1355,N_1228);
nand U1665 (N_1665,N_1479,N_1399);
xnor U1666 (N_1666,N_1484,N_1372);
xor U1667 (N_1667,N_1488,N_1290);
nor U1668 (N_1668,N_1206,N_1489);
nor U1669 (N_1669,N_1329,N_1477);
nor U1670 (N_1670,N_1462,N_1445);
xor U1671 (N_1671,N_1458,N_1449);
nor U1672 (N_1672,N_1494,N_1271);
nor U1673 (N_1673,N_1324,N_1315);
xor U1674 (N_1674,N_1351,N_1303);
xnor U1675 (N_1675,N_1294,N_1291);
or U1676 (N_1676,N_1361,N_1354);
nand U1677 (N_1677,N_1395,N_1282);
and U1678 (N_1678,N_1219,N_1260);
xor U1679 (N_1679,N_1390,N_1305);
or U1680 (N_1680,N_1442,N_1313);
and U1681 (N_1681,N_1266,N_1225);
or U1682 (N_1682,N_1261,N_1371);
and U1683 (N_1683,N_1427,N_1294);
xnor U1684 (N_1684,N_1223,N_1268);
xnor U1685 (N_1685,N_1340,N_1410);
and U1686 (N_1686,N_1383,N_1387);
xor U1687 (N_1687,N_1315,N_1367);
and U1688 (N_1688,N_1303,N_1290);
and U1689 (N_1689,N_1227,N_1219);
xor U1690 (N_1690,N_1349,N_1419);
and U1691 (N_1691,N_1211,N_1412);
nand U1692 (N_1692,N_1465,N_1336);
or U1693 (N_1693,N_1398,N_1229);
nor U1694 (N_1694,N_1221,N_1398);
nor U1695 (N_1695,N_1279,N_1273);
and U1696 (N_1696,N_1353,N_1365);
xnor U1697 (N_1697,N_1263,N_1425);
nand U1698 (N_1698,N_1339,N_1428);
or U1699 (N_1699,N_1332,N_1248);
xnor U1700 (N_1700,N_1217,N_1288);
xor U1701 (N_1701,N_1363,N_1486);
xnor U1702 (N_1702,N_1302,N_1380);
and U1703 (N_1703,N_1369,N_1373);
xnor U1704 (N_1704,N_1431,N_1398);
xor U1705 (N_1705,N_1411,N_1268);
nor U1706 (N_1706,N_1324,N_1446);
and U1707 (N_1707,N_1347,N_1309);
xnor U1708 (N_1708,N_1305,N_1461);
or U1709 (N_1709,N_1238,N_1445);
xnor U1710 (N_1710,N_1272,N_1372);
and U1711 (N_1711,N_1441,N_1317);
nand U1712 (N_1712,N_1441,N_1222);
nor U1713 (N_1713,N_1219,N_1221);
and U1714 (N_1714,N_1208,N_1289);
or U1715 (N_1715,N_1417,N_1318);
nand U1716 (N_1716,N_1248,N_1457);
or U1717 (N_1717,N_1284,N_1352);
or U1718 (N_1718,N_1265,N_1348);
xnor U1719 (N_1719,N_1311,N_1294);
and U1720 (N_1720,N_1330,N_1409);
xor U1721 (N_1721,N_1320,N_1365);
nor U1722 (N_1722,N_1388,N_1301);
and U1723 (N_1723,N_1296,N_1472);
and U1724 (N_1724,N_1374,N_1283);
nor U1725 (N_1725,N_1333,N_1314);
xor U1726 (N_1726,N_1210,N_1258);
xnor U1727 (N_1727,N_1283,N_1334);
nor U1728 (N_1728,N_1214,N_1405);
nor U1729 (N_1729,N_1436,N_1200);
or U1730 (N_1730,N_1407,N_1405);
xor U1731 (N_1731,N_1212,N_1375);
or U1732 (N_1732,N_1260,N_1484);
nand U1733 (N_1733,N_1370,N_1350);
nor U1734 (N_1734,N_1357,N_1360);
xnor U1735 (N_1735,N_1365,N_1471);
nand U1736 (N_1736,N_1381,N_1430);
xnor U1737 (N_1737,N_1444,N_1272);
nor U1738 (N_1738,N_1207,N_1274);
or U1739 (N_1739,N_1394,N_1225);
nand U1740 (N_1740,N_1445,N_1316);
or U1741 (N_1741,N_1292,N_1357);
and U1742 (N_1742,N_1235,N_1272);
nor U1743 (N_1743,N_1367,N_1394);
and U1744 (N_1744,N_1492,N_1471);
xnor U1745 (N_1745,N_1387,N_1322);
or U1746 (N_1746,N_1295,N_1352);
nor U1747 (N_1747,N_1463,N_1415);
nor U1748 (N_1748,N_1469,N_1233);
nand U1749 (N_1749,N_1389,N_1348);
nand U1750 (N_1750,N_1317,N_1380);
nor U1751 (N_1751,N_1365,N_1269);
nor U1752 (N_1752,N_1365,N_1356);
xor U1753 (N_1753,N_1281,N_1257);
and U1754 (N_1754,N_1202,N_1212);
xor U1755 (N_1755,N_1383,N_1423);
nor U1756 (N_1756,N_1399,N_1319);
and U1757 (N_1757,N_1378,N_1224);
nor U1758 (N_1758,N_1271,N_1286);
nor U1759 (N_1759,N_1418,N_1348);
and U1760 (N_1760,N_1315,N_1343);
or U1761 (N_1761,N_1295,N_1333);
and U1762 (N_1762,N_1496,N_1344);
or U1763 (N_1763,N_1255,N_1211);
nand U1764 (N_1764,N_1490,N_1425);
nor U1765 (N_1765,N_1360,N_1297);
or U1766 (N_1766,N_1405,N_1264);
or U1767 (N_1767,N_1472,N_1384);
nand U1768 (N_1768,N_1314,N_1305);
xnor U1769 (N_1769,N_1445,N_1260);
nor U1770 (N_1770,N_1464,N_1319);
nand U1771 (N_1771,N_1485,N_1412);
nor U1772 (N_1772,N_1390,N_1219);
and U1773 (N_1773,N_1270,N_1401);
nor U1774 (N_1774,N_1218,N_1458);
xor U1775 (N_1775,N_1400,N_1233);
nor U1776 (N_1776,N_1233,N_1402);
xnor U1777 (N_1777,N_1265,N_1473);
nand U1778 (N_1778,N_1359,N_1416);
or U1779 (N_1779,N_1396,N_1384);
or U1780 (N_1780,N_1282,N_1387);
nor U1781 (N_1781,N_1361,N_1267);
xor U1782 (N_1782,N_1303,N_1214);
xor U1783 (N_1783,N_1309,N_1427);
xor U1784 (N_1784,N_1409,N_1456);
or U1785 (N_1785,N_1453,N_1475);
nor U1786 (N_1786,N_1331,N_1356);
and U1787 (N_1787,N_1388,N_1241);
xor U1788 (N_1788,N_1397,N_1302);
xnor U1789 (N_1789,N_1315,N_1229);
and U1790 (N_1790,N_1202,N_1482);
and U1791 (N_1791,N_1396,N_1391);
nand U1792 (N_1792,N_1341,N_1474);
nand U1793 (N_1793,N_1449,N_1291);
or U1794 (N_1794,N_1339,N_1374);
or U1795 (N_1795,N_1321,N_1496);
xnor U1796 (N_1796,N_1325,N_1336);
xnor U1797 (N_1797,N_1452,N_1265);
and U1798 (N_1798,N_1392,N_1497);
xor U1799 (N_1799,N_1481,N_1497);
xor U1800 (N_1800,N_1609,N_1633);
nand U1801 (N_1801,N_1763,N_1637);
nor U1802 (N_1802,N_1699,N_1624);
and U1803 (N_1803,N_1590,N_1658);
nor U1804 (N_1804,N_1631,N_1589);
nor U1805 (N_1805,N_1749,N_1772);
and U1806 (N_1806,N_1758,N_1720);
nand U1807 (N_1807,N_1782,N_1615);
xor U1808 (N_1808,N_1536,N_1646);
xnor U1809 (N_1809,N_1706,N_1565);
and U1810 (N_1810,N_1604,N_1632);
nand U1811 (N_1811,N_1744,N_1503);
nor U1812 (N_1812,N_1783,N_1550);
nor U1813 (N_1813,N_1725,N_1579);
or U1814 (N_1814,N_1515,N_1520);
or U1815 (N_1815,N_1771,N_1788);
nand U1816 (N_1816,N_1601,N_1618);
or U1817 (N_1817,N_1792,N_1648);
and U1818 (N_1818,N_1678,N_1671);
nand U1819 (N_1819,N_1751,N_1689);
nand U1820 (N_1820,N_1681,N_1574);
nor U1821 (N_1821,N_1755,N_1791);
xnor U1822 (N_1822,N_1661,N_1641);
nor U1823 (N_1823,N_1533,N_1760);
nand U1824 (N_1824,N_1716,N_1532);
nand U1825 (N_1825,N_1786,N_1713);
nand U1826 (N_1826,N_1572,N_1683);
and U1827 (N_1827,N_1636,N_1587);
and U1828 (N_1828,N_1710,N_1531);
xor U1829 (N_1829,N_1701,N_1798);
or U1830 (N_1830,N_1659,N_1595);
xnor U1831 (N_1831,N_1656,N_1748);
xnor U1832 (N_1832,N_1702,N_1573);
nor U1833 (N_1833,N_1688,N_1784);
nand U1834 (N_1834,N_1500,N_1645);
and U1835 (N_1835,N_1665,N_1516);
nand U1836 (N_1836,N_1700,N_1558);
nor U1837 (N_1837,N_1630,N_1793);
xnor U1838 (N_1838,N_1727,N_1651);
xnor U1839 (N_1839,N_1660,N_1704);
nand U1840 (N_1840,N_1785,N_1757);
nor U1841 (N_1841,N_1605,N_1745);
xor U1842 (N_1842,N_1512,N_1570);
xor U1843 (N_1843,N_1717,N_1740);
and U1844 (N_1844,N_1542,N_1730);
nor U1845 (N_1845,N_1790,N_1649);
xnor U1846 (N_1846,N_1567,N_1770);
xor U1847 (N_1847,N_1626,N_1766);
nand U1848 (N_1848,N_1606,N_1509);
or U1849 (N_1849,N_1682,N_1508);
xor U1850 (N_1850,N_1707,N_1692);
or U1851 (N_1851,N_1623,N_1639);
xor U1852 (N_1852,N_1582,N_1691);
xor U1853 (N_1853,N_1724,N_1553);
xnor U1854 (N_1854,N_1764,N_1657);
nand U1855 (N_1855,N_1663,N_1610);
xnor U1856 (N_1856,N_1695,N_1625);
nand U1857 (N_1857,N_1685,N_1735);
xor U1858 (N_1858,N_1799,N_1577);
and U1859 (N_1859,N_1709,N_1591);
and U1860 (N_1860,N_1539,N_1737);
or U1861 (N_1861,N_1547,N_1712);
nand U1862 (N_1862,N_1540,N_1629);
nor U1863 (N_1863,N_1680,N_1753);
and U1864 (N_1864,N_1543,N_1673);
nor U1865 (N_1865,N_1557,N_1675);
xor U1866 (N_1866,N_1527,N_1703);
nor U1867 (N_1867,N_1722,N_1654);
and U1868 (N_1868,N_1777,N_1664);
or U1869 (N_1869,N_1655,N_1779);
nand U1870 (N_1870,N_1562,N_1556);
nand U1871 (N_1871,N_1555,N_1768);
and U1872 (N_1872,N_1732,N_1674);
nand U1873 (N_1873,N_1686,N_1599);
nand U1874 (N_1874,N_1693,N_1612);
nor U1875 (N_1875,N_1723,N_1514);
and U1876 (N_1876,N_1787,N_1511);
xnor U1877 (N_1877,N_1552,N_1564);
xor U1878 (N_1878,N_1726,N_1690);
or U1879 (N_1879,N_1521,N_1635);
xnor U1880 (N_1880,N_1642,N_1721);
or U1881 (N_1881,N_1506,N_1667);
and U1882 (N_1882,N_1714,N_1580);
nand U1883 (N_1883,N_1762,N_1780);
nand U1884 (N_1884,N_1687,N_1597);
nor U1885 (N_1885,N_1734,N_1526);
or U1886 (N_1886,N_1694,N_1608);
xnor U1887 (N_1887,N_1541,N_1617);
xor U1888 (N_1888,N_1769,N_1776);
nand U1889 (N_1889,N_1593,N_1781);
nand U1890 (N_1890,N_1736,N_1621);
and U1891 (N_1891,N_1743,N_1505);
nor U1892 (N_1892,N_1662,N_1530);
nor U1893 (N_1893,N_1602,N_1554);
xnor U1894 (N_1894,N_1747,N_1560);
and U1895 (N_1895,N_1775,N_1529);
xor U1896 (N_1896,N_1698,N_1568);
and U1897 (N_1897,N_1611,N_1718);
xnor U1898 (N_1898,N_1729,N_1644);
and U1899 (N_1899,N_1739,N_1652);
and U1900 (N_1900,N_1634,N_1679);
or U1901 (N_1901,N_1517,N_1684);
nand U1902 (N_1902,N_1669,N_1650);
xnor U1903 (N_1903,N_1607,N_1584);
xnor U1904 (N_1904,N_1696,N_1738);
nand U1905 (N_1905,N_1549,N_1594);
or U1906 (N_1906,N_1619,N_1653);
xnor U1907 (N_1907,N_1666,N_1774);
or U1908 (N_1908,N_1742,N_1566);
xnor U1909 (N_1909,N_1647,N_1754);
nand U1910 (N_1910,N_1537,N_1583);
nor U1911 (N_1911,N_1796,N_1705);
nor U1912 (N_1912,N_1643,N_1773);
or U1913 (N_1913,N_1524,N_1640);
and U1914 (N_1914,N_1789,N_1596);
nand U1915 (N_1915,N_1510,N_1563);
or U1916 (N_1916,N_1676,N_1546);
or U1917 (N_1917,N_1588,N_1585);
xor U1918 (N_1918,N_1741,N_1561);
nand U1919 (N_1919,N_1711,N_1519);
nor U1920 (N_1920,N_1613,N_1797);
nor U1921 (N_1921,N_1750,N_1767);
xor U1922 (N_1922,N_1668,N_1616);
nor U1923 (N_1923,N_1528,N_1534);
nor U1924 (N_1924,N_1501,N_1627);
nand U1925 (N_1925,N_1746,N_1614);
nand U1926 (N_1926,N_1507,N_1545);
xor U1927 (N_1927,N_1733,N_1715);
xnor U1928 (N_1928,N_1544,N_1759);
or U1929 (N_1929,N_1677,N_1628);
and U1930 (N_1930,N_1622,N_1581);
or U1931 (N_1931,N_1752,N_1765);
or U1932 (N_1932,N_1523,N_1620);
xnor U1933 (N_1933,N_1559,N_1522);
and U1934 (N_1934,N_1504,N_1794);
xor U1935 (N_1935,N_1535,N_1525);
xor U1936 (N_1936,N_1670,N_1598);
nand U1937 (N_1937,N_1571,N_1502);
nor U1938 (N_1938,N_1586,N_1600);
xnor U1939 (N_1939,N_1548,N_1578);
or U1940 (N_1940,N_1697,N_1672);
xnor U1941 (N_1941,N_1551,N_1592);
xnor U1942 (N_1942,N_1603,N_1731);
nand U1943 (N_1943,N_1569,N_1575);
nand U1944 (N_1944,N_1795,N_1576);
and U1945 (N_1945,N_1538,N_1778);
xor U1946 (N_1946,N_1756,N_1708);
nor U1947 (N_1947,N_1719,N_1638);
nor U1948 (N_1948,N_1513,N_1728);
nor U1949 (N_1949,N_1761,N_1518);
or U1950 (N_1950,N_1588,N_1500);
nand U1951 (N_1951,N_1602,N_1622);
nand U1952 (N_1952,N_1754,N_1675);
nand U1953 (N_1953,N_1762,N_1618);
and U1954 (N_1954,N_1646,N_1645);
or U1955 (N_1955,N_1755,N_1564);
xnor U1956 (N_1956,N_1750,N_1633);
and U1957 (N_1957,N_1659,N_1775);
nor U1958 (N_1958,N_1696,N_1598);
or U1959 (N_1959,N_1503,N_1576);
or U1960 (N_1960,N_1558,N_1782);
or U1961 (N_1961,N_1572,N_1676);
nor U1962 (N_1962,N_1571,N_1548);
or U1963 (N_1963,N_1555,N_1529);
xor U1964 (N_1964,N_1618,N_1777);
nand U1965 (N_1965,N_1688,N_1568);
nor U1966 (N_1966,N_1515,N_1502);
or U1967 (N_1967,N_1676,N_1607);
nand U1968 (N_1968,N_1551,N_1720);
or U1969 (N_1969,N_1515,N_1556);
or U1970 (N_1970,N_1768,N_1697);
nand U1971 (N_1971,N_1595,N_1711);
xnor U1972 (N_1972,N_1633,N_1791);
and U1973 (N_1973,N_1686,N_1549);
nand U1974 (N_1974,N_1504,N_1734);
and U1975 (N_1975,N_1697,N_1792);
and U1976 (N_1976,N_1772,N_1783);
nand U1977 (N_1977,N_1566,N_1547);
xnor U1978 (N_1978,N_1777,N_1588);
or U1979 (N_1979,N_1689,N_1667);
xor U1980 (N_1980,N_1567,N_1778);
nand U1981 (N_1981,N_1665,N_1648);
or U1982 (N_1982,N_1639,N_1650);
xor U1983 (N_1983,N_1526,N_1588);
xnor U1984 (N_1984,N_1714,N_1754);
or U1985 (N_1985,N_1564,N_1765);
xnor U1986 (N_1986,N_1739,N_1601);
xor U1987 (N_1987,N_1570,N_1684);
nor U1988 (N_1988,N_1638,N_1531);
nor U1989 (N_1989,N_1524,N_1617);
nand U1990 (N_1990,N_1543,N_1512);
nor U1991 (N_1991,N_1566,N_1683);
and U1992 (N_1992,N_1774,N_1518);
nor U1993 (N_1993,N_1722,N_1703);
xnor U1994 (N_1994,N_1762,N_1570);
or U1995 (N_1995,N_1600,N_1523);
xor U1996 (N_1996,N_1503,N_1644);
nand U1997 (N_1997,N_1611,N_1721);
nand U1998 (N_1998,N_1742,N_1682);
nor U1999 (N_1999,N_1602,N_1728);
or U2000 (N_2000,N_1779,N_1631);
or U2001 (N_2001,N_1658,N_1672);
nor U2002 (N_2002,N_1500,N_1542);
xnor U2003 (N_2003,N_1567,N_1501);
nand U2004 (N_2004,N_1767,N_1688);
nand U2005 (N_2005,N_1793,N_1779);
nor U2006 (N_2006,N_1604,N_1784);
nor U2007 (N_2007,N_1623,N_1532);
or U2008 (N_2008,N_1562,N_1698);
nand U2009 (N_2009,N_1764,N_1580);
nor U2010 (N_2010,N_1636,N_1578);
and U2011 (N_2011,N_1796,N_1751);
xor U2012 (N_2012,N_1664,N_1665);
nor U2013 (N_2013,N_1742,N_1650);
and U2014 (N_2014,N_1596,N_1692);
nor U2015 (N_2015,N_1781,N_1706);
nor U2016 (N_2016,N_1544,N_1722);
xor U2017 (N_2017,N_1501,N_1580);
xnor U2018 (N_2018,N_1691,N_1571);
nor U2019 (N_2019,N_1622,N_1528);
xnor U2020 (N_2020,N_1518,N_1753);
xor U2021 (N_2021,N_1556,N_1596);
and U2022 (N_2022,N_1788,N_1577);
or U2023 (N_2023,N_1538,N_1526);
or U2024 (N_2024,N_1633,N_1714);
and U2025 (N_2025,N_1587,N_1649);
nand U2026 (N_2026,N_1710,N_1589);
or U2027 (N_2027,N_1507,N_1725);
nor U2028 (N_2028,N_1547,N_1543);
nor U2029 (N_2029,N_1530,N_1663);
xnor U2030 (N_2030,N_1799,N_1775);
xor U2031 (N_2031,N_1743,N_1671);
nor U2032 (N_2032,N_1704,N_1636);
nand U2033 (N_2033,N_1763,N_1685);
and U2034 (N_2034,N_1581,N_1656);
and U2035 (N_2035,N_1726,N_1728);
nor U2036 (N_2036,N_1654,N_1513);
xor U2037 (N_2037,N_1673,N_1684);
or U2038 (N_2038,N_1639,N_1798);
or U2039 (N_2039,N_1721,N_1724);
nor U2040 (N_2040,N_1504,N_1793);
xor U2041 (N_2041,N_1616,N_1664);
and U2042 (N_2042,N_1582,N_1579);
xor U2043 (N_2043,N_1599,N_1506);
xor U2044 (N_2044,N_1762,N_1538);
and U2045 (N_2045,N_1673,N_1525);
nand U2046 (N_2046,N_1668,N_1650);
or U2047 (N_2047,N_1642,N_1750);
nand U2048 (N_2048,N_1585,N_1647);
or U2049 (N_2049,N_1617,N_1575);
nor U2050 (N_2050,N_1730,N_1587);
or U2051 (N_2051,N_1691,N_1710);
nand U2052 (N_2052,N_1501,N_1584);
or U2053 (N_2053,N_1535,N_1519);
nand U2054 (N_2054,N_1559,N_1642);
or U2055 (N_2055,N_1528,N_1728);
or U2056 (N_2056,N_1620,N_1648);
nand U2057 (N_2057,N_1606,N_1575);
nand U2058 (N_2058,N_1556,N_1663);
and U2059 (N_2059,N_1717,N_1662);
nor U2060 (N_2060,N_1762,N_1643);
and U2061 (N_2061,N_1533,N_1742);
nor U2062 (N_2062,N_1576,N_1799);
or U2063 (N_2063,N_1662,N_1668);
nand U2064 (N_2064,N_1573,N_1563);
xor U2065 (N_2065,N_1549,N_1692);
and U2066 (N_2066,N_1694,N_1733);
nand U2067 (N_2067,N_1530,N_1532);
nand U2068 (N_2068,N_1539,N_1529);
nor U2069 (N_2069,N_1649,N_1750);
xnor U2070 (N_2070,N_1630,N_1570);
and U2071 (N_2071,N_1598,N_1776);
nor U2072 (N_2072,N_1523,N_1646);
nand U2073 (N_2073,N_1565,N_1663);
nand U2074 (N_2074,N_1614,N_1734);
or U2075 (N_2075,N_1724,N_1620);
or U2076 (N_2076,N_1524,N_1656);
nor U2077 (N_2077,N_1758,N_1799);
nor U2078 (N_2078,N_1506,N_1581);
nor U2079 (N_2079,N_1620,N_1785);
nor U2080 (N_2080,N_1798,N_1510);
and U2081 (N_2081,N_1683,N_1553);
nor U2082 (N_2082,N_1638,N_1591);
or U2083 (N_2083,N_1598,N_1608);
xnor U2084 (N_2084,N_1596,N_1612);
nor U2085 (N_2085,N_1505,N_1639);
or U2086 (N_2086,N_1789,N_1551);
or U2087 (N_2087,N_1619,N_1668);
and U2088 (N_2088,N_1606,N_1570);
xor U2089 (N_2089,N_1699,N_1701);
or U2090 (N_2090,N_1717,N_1770);
and U2091 (N_2091,N_1504,N_1646);
nand U2092 (N_2092,N_1563,N_1585);
xnor U2093 (N_2093,N_1554,N_1576);
and U2094 (N_2094,N_1688,N_1570);
or U2095 (N_2095,N_1729,N_1531);
or U2096 (N_2096,N_1792,N_1667);
and U2097 (N_2097,N_1520,N_1567);
and U2098 (N_2098,N_1505,N_1667);
nand U2099 (N_2099,N_1565,N_1765);
nand U2100 (N_2100,N_1955,N_2005);
and U2101 (N_2101,N_2001,N_2074);
or U2102 (N_2102,N_2020,N_1837);
or U2103 (N_2103,N_2063,N_2078);
nand U2104 (N_2104,N_1801,N_2077);
or U2105 (N_2105,N_1853,N_1977);
nor U2106 (N_2106,N_1831,N_1859);
and U2107 (N_2107,N_2013,N_2099);
or U2108 (N_2108,N_1940,N_1805);
xnor U2109 (N_2109,N_2095,N_1843);
and U2110 (N_2110,N_1972,N_1881);
or U2111 (N_2111,N_1849,N_1941);
nand U2112 (N_2112,N_2058,N_1932);
and U2113 (N_2113,N_1855,N_1850);
nand U2114 (N_2114,N_1839,N_1872);
or U2115 (N_2115,N_2067,N_2047);
nand U2116 (N_2116,N_1998,N_1844);
nor U2117 (N_2117,N_1988,N_2002);
and U2118 (N_2118,N_1928,N_1866);
and U2119 (N_2119,N_1820,N_1981);
and U2120 (N_2120,N_1807,N_1826);
nand U2121 (N_2121,N_2019,N_1957);
and U2122 (N_2122,N_2083,N_1838);
nor U2123 (N_2123,N_1871,N_1834);
xnor U2124 (N_2124,N_2043,N_2096);
nor U2125 (N_2125,N_1821,N_2040);
or U2126 (N_2126,N_1817,N_1861);
nand U2127 (N_2127,N_1912,N_2000);
xnor U2128 (N_2128,N_2012,N_1914);
or U2129 (N_2129,N_1814,N_1869);
nor U2130 (N_2130,N_2036,N_1951);
nand U2131 (N_2131,N_1999,N_1898);
xnor U2132 (N_2132,N_1846,N_1904);
xor U2133 (N_2133,N_1994,N_2051);
and U2134 (N_2134,N_1931,N_1933);
and U2135 (N_2135,N_2084,N_1927);
nand U2136 (N_2136,N_1873,N_2009);
nor U2137 (N_2137,N_1929,N_1895);
nor U2138 (N_2138,N_2094,N_2022);
nor U2139 (N_2139,N_1910,N_2089);
nand U2140 (N_2140,N_2090,N_2097);
and U2141 (N_2141,N_1970,N_1891);
and U2142 (N_2142,N_2070,N_1811);
xor U2143 (N_2143,N_1857,N_2024);
nand U2144 (N_2144,N_2007,N_1824);
nor U2145 (N_2145,N_1819,N_1980);
or U2146 (N_2146,N_2080,N_1863);
or U2147 (N_2147,N_2011,N_1847);
or U2148 (N_2148,N_1806,N_1969);
nand U2149 (N_2149,N_2098,N_1973);
nand U2150 (N_2150,N_2082,N_1887);
nor U2151 (N_2151,N_1936,N_1832);
and U2152 (N_2152,N_2032,N_2057);
nor U2153 (N_2153,N_1854,N_2065);
xor U2154 (N_2154,N_1939,N_1968);
nand U2155 (N_2155,N_1874,N_1845);
or U2156 (N_2156,N_2062,N_2091);
and U2157 (N_2157,N_1935,N_1996);
nor U2158 (N_2158,N_2041,N_1848);
and U2159 (N_2159,N_1860,N_2087);
and U2160 (N_2160,N_1841,N_1946);
and U2161 (N_2161,N_2044,N_1802);
or U2162 (N_2162,N_1913,N_2055);
xnor U2163 (N_2163,N_1890,N_1959);
nand U2164 (N_2164,N_1963,N_1903);
nand U2165 (N_2165,N_1956,N_1856);
nand U2166 (N_2166,N_2086,N_2072);
nor U2167 (N_2167,N_1897,N_1810);
nor U2168 (N_2168,N_1813,N_1923);
nand U2169 (N_2169,N_2033,N_1938);
or U2170 (N_2170,N_2008,N_1985);
xnor U2171 (N_2171,N_2054,N_2034);
or U2172 (N_2172,N_1883,N_1888);
and U2173 (N_2173,N_2004,N_2010);
or U2174 (N_2174,N_2035,N_1829);
or U2175 (N_2175,N_1907,N_1880);
nand U2176 (N_2176,N_1930,N_1879);
xor U2177 (N_2177,N_1840,N_2059);
nand U2178 (N_2178,N_1948,N_2030);
nor U2179 (N_2179,N_1962,N_1809);
or U2180 (N_2180,N_2068,N_1989);
nor U2181 (N_2181,N_1919,N_2092);
and U2182 (N_2182,N_1833,N_1953);
or U2183 (N_2183,N_1920,N_1918);
nand U2184 (N_2184,N_1876,N_1896);
nor U2185 (N_2185,N_2079,N_2073);
xnor U2186 (N_2186,N_2017,N_2014);
nand U2187 (N_2187,N_2060,N_1967);
nand U2188 (N_2188,N_2046,N_1925);
nor U2189 (N_2189,N_1842,N_1945);
nand U2190 (N_2190,N_1952,N_1892);
or U2191 (N_2191,N_1954,N_2064);
and U2192 (N_2192,N_2026,N_1862);
xnor U2193 (N_2193,N_2069,N_1991);
and U2194 (N_2194,N_2045,N_2038);
nand U2195 (N_2195,N_1978,N_1905);
nand U2196 (N_2196,N_1965,N_2021);
and U2197 (N_2197,N_1894,N_1966);
or U2198 (N_2198,N_2088,N_1867);
nand U2199 (N_2199,N_1902,N_1958);
and U2200 (N_2200,N_1922,N_1858);
xnor U2201 (N_2201,N_2056,N_1868);
and U2202 (N_2202,N_1818,N_1815);
nand U2203 (N_2203,N_1816,N_1964);
xnor U2204 (N_2204,N_1979,N_1911);
and U2205 (N_2205,N_2075,N_2027);
and U2206 (N_2206,N_1915,N_1906);
and U2207 (N_2207,N_2076,N_2071);
xor U2208 (N_2208,N_1835,N_1943);
nor U2209 (N_2209,N_1983,N_2015);
or U2210 (N_2210,N_1825,N_1934);
xnor U2211 (N_2211,N_1900,N_1974);
xnor U2212 (N_2212,N_1917,N_1921);
and U2213 (N_2213,N_1916,N_1947);
xnor U2214 (N_2214,N_2050,N_1942);
xnor U2215 (N_2215,N_1830,N_2039);
nor U2216 (N_2216,N_1975,N_2006);
xnor U2217 (N_2217,N_2025,N_1870);
nor U2218 (N_2218,N_2052,N_2049);
and U2219 (N_2219,N_1995,N_1808);
nand U2220 (N_2220,N_1949,N_2029);
nand U2221 (N_2221,N_1950,N_1909);
and U2222 (N_2222,N_1877,N_1990);
and U2223 (N_2223,N_1926,N_1800);
and U2224 (N_2224,N_1827,N_2061);
and U2225 (N_2225,N_2066,N_2053);
nand U2226 (N_2226,N_2031,N_1893);
or U2227 (N_2227,N_1886,N_2003);
xnor U2228 (N_2228,N_1889,N_1982);
nand U2229 (N_2229,N_1993,N_1937);
or U2230 (N_2230,N_1823,N_2023);
xor U2231 (N_2231,N_1822,N_1864);
nor U2232 (N_2232,N_1901,N_2081);
or U2233 (N_2233,N_1961,N_1992);
xnor U2234 (N_2234,N_1984,N_1851);
nor U2235 (N_2235,N_1836,N_1803);
nor U2236 (N_2236,N_1924,N_1987);
xor U2237 (N_2237,N_2037,N_2028);
nor U2238 (N_2238,N_1884,N_1882);
nand U2239 (N_2239,N_2085,N_2016);
nand U2240 (N_2240,N_1971,N_1885);
or U2241 (N_2241,N_1944,N_1997);
xor U2242 (N_2242,N_2042,N_1878);
nor U2243 (N_2243,N_1812,N_2048);
nor U2244 (N_2244,N_2018,N_1852);
xnor U2245 (N_2245,N_2093,N_1804);
or U2246 (N_2246,N_1899,N_1986);
nand U2247 (N_2247,N_1875,N_1960);
nor U2248 (N_2248,N_1976,N_1828);
and U2249 (N_2249,N_1865,N_1908);
nand U2250 (N_2250,N_1868,N_1988);
nor U2251 (N_2251,N_1869,N_1812);
xnor U2252 (N_2252,N_1866,N_1957);
nor U2253 (N_2253,N_2040,N_1841);
nor U2254 (N_2254,N_1969,N_1923);
nand U2255 (N_2255,N_2052,N_2062);
or U2256 (N_2256,N_1971,N_1967);
nor U2257 (N_2257,N_1872,N_2070);
nor U2258 (N_2258,N_1916,N_1836);
nor U2259 (N_2259,N_1856,N_1948);
nand U2260 (N_2260,N_1988,N_1985);
or U2261 (N_2261,N_2071,N_1855);
nand U2262 (N_2262,N_2099,N_1819);
nand U2263 (N_2263,N_1921,N_1972);
or U2264 (N_2264,N_1811,N_1900);
xor U2265 (N_2265,N_1997,N_2067);
xnor U2266 (N_2266,N_1893,N_1911);
and U2267 (N_2267,N_1832,N_1938);
nand U2268 (N_2268,N_1822,N_2010);
and U2269 (N_2269,N_1805,N_1911);
nand U2270 (N_2270,N_2084,N_1885);
or U2271 (N_2271,N_1954,N_1951);
nor U2272 (N_2272,N_1983,N_2051);
xnor U2273 (N_2273,N_1835,N_1888);
nor U2274 (N_2274,N_1808,N_2098);
or U2275 (N_2275,N_2040,N_2018);
nor U2276 (N_2276,N_2079,N_2016);
xor U2277 (N_2277,N_2097,N_1899);
and U2278 (N_2278,N_2041,N_1894);
nor U2279 (N_2279,N_1961,N_1878);
nor U2280 (N_2280,N_1905,N_1879);
xor U2281 (N_2281,N_1921,N_1800);
and U2282 (N_2282,N_1911,N_2041);
nor U2283 (N_2283,N_2015,N_1924);
nor U2284 (N_2284,N_1919,N_1942);
nand U2285 (N_2285,N_1864,N_1868);
xnor U2286 (N_2286,N_2042,N_2003);
nor U2287 (N_2287,N_1893,N_1833);
nand U2288 (N_2288,N_1817,N_1971);
and U2289 (N_2289,N_1867,N_1895);
or U2290 (N_2290,N_1833,N_1841);
nor U2291 (N_2291,N_2028,N_1852);
xnor U2292 (N_2292,N_2065,N_1944);
and U2293 (N_2293,N_2080,N_1967);
nor U2294 (N_2294,N_1881,N_2061);
or U2295 (N_2295,N_2035,N_1952);
nand U2296 (N_2296,N_1947,N_1997);
nand U2297 (N_2297,N_1896,N_2040);
and U2298 (N_2298,N_1968,N_1985);
or U2299 (N_2299,N_2098,N_2005);
and U2300 (N_2300,N_1871,N_1899);
nor U2301 (N_2301,N_1907,N_1961);
xnor U2302 (N_2302,N_1850,N_2098);
nand U2303 (N_2303,N_2094,N_1917);
nand U2304 (N_2304,N_1852,N_1891);
xnor U2305 (N_2305,N_2070,N_1936);
nor U2306 (N_2306,N_2037,N_1932);
and U2307 (N_2307,N_1962,N_1845);
or U2308 (N_2308,N_1969,N_1996);
xor U2309 (N_2309,N_2052,N_1821);
nor U2310 (N_2310,N_1835,N_1865);
nand U2311 (N_2311,N_1898,N_1932);
xnor U2312 (N_2312,N_1832,N_2034);
and U2313 (N_2313,N_2099,N_2098);
nand U2314 (N_2314,N_2020,N_2076);
or U2315 (N_2315,N_2004,N_1836);
xnor U2316 (N_2316,N_1966,N_2034);
or U2317 (N_2317,N_1884,N_1969);
xor U2318 (N_2318,N_1959,N_1990);
nand U2319 (N_2319,N_1932,N_1807);
nor U2320 (N_2320,N_1860,N_1812);
or U2321 (N_2321,N_2022,N_1857);
xor U2322 (N_2322,N_1934,N_2077);
or U2323 (N_2323,N_2076,N_1937);
nor U2324 (N_2324,N_1945,N_1876);
xor U2325 (N_2325,N_2072,N_1971);
and U2326 (N_2326,N_2039,N_2062);
xor U2327 (N_2327,N_2087,N_1800);
and U2328 (N_2328,N_2083,N_1923);
nor U2329 (N_2329,N_2061,N_1851);
xnor U2330 (N_2330,N_2007,N_1870);
nor U2331 (N_2331,N_1848,N_1819);
nand U2332 (N_2332,N_2051,N_2071);
or U2333 (N_2333,N_2073,N_1940);
and U2334 (N_2334,N_1932,N_1964);
or U2335 (N_2335,N_2052,N_1961);
xnor U2336 (N_2336,N_2017,N_2050);
xor U2337 (N_2337,N_1934,N_1986);
and U2338 (N_2338,N_1884,N_1837);
or U2339 (N_2339,N_1840,N_1950);
nand U2340 (N_2340,N_1967,N_2022);
nand U2341 (N_2341,N_1859,N_2067);
and U2342 (N_2342,N_1982,N_2057);
nand U2343 (N_2343,N_2029,N_2036);
xnor U2344 (N_2344,N_2034,N_1882);
nand U2345 (N_2345,N_1950,N_1831);
nor U2346 (N_2346,N_2001,N_1808);
nor U2347 (N_2347,N_1877,N_2066);
or U2348 (N_2348,N_1834,N_2087);
nor U2349 (N_2349,N_1861,N_2098);
nor U2350 (N_2350,N_1896,N_2084);
nand U2351 (N_2351,N_1834,N_2073);
nand U2352 (N_2352,N_1872,N_1966);
or U2353 (N_2353,N_1973,N_2053);
nand U2354 (N_2354,N_1853,N_1831);
nand U2355 (N_2355,N_2083,N_1900);
xnor U2356 (N_2356,N_1933,N_2028);
or U2357 (N_2357,N_1858,N_2086);
and U2358 (N_2358,N_1861,N_1949);
nor U2359 (N_2359,N_2029,N_1848);
nand U2360 (N_2360,N_2060,N_1880);
nor U2361 (N_2361,N_1905,N_2064);
nor U2362 (N_2362,N_1802,N_1884);
nor U2363 (N_2363,N_1962,N_1874);
or U2364 (N_2364,N_1841,N_1819);
xnor U2365 (N_2365,N_1895,N_2020);
and U2366 (N_2366,N_1927,N_1868);
or U2367 (N_2367,N_2044,N_2094);
xor U2368 (N_2368,N_1822,N_2006);
nand U2369 (N_2369,N_2048,N_2030);
xnor U2370 (N_2370,N_1945,N_1954);
xnor U2371 (N_2371,N_1878,N_2047);
or U2372 (N_2372,N_1905,N_1962);
and U2373 (N_2373,N_1846,N_1808);
nor U2374 (N_2374,N_1892,N_1909);
nor U2375 (N_2375,N_1859,N_1989);
nand U2376 (N_2376,N_1970,N_1816);
or U2377 (N_2377,N_2088,N_2066);
and U2378 (N_2378,N_1878,N_1837);
nand U2379 (N_2379,N_2028,N_2088);
nor U2380 (N_2380,N_2023,N_1945);
or U2381 (N_2381,N_1839,N_1821);
nand U2382 (N_2382,N_2043,N_1860);
nand U2383 (N_2383,N_1955,N_2065);
xnor U2384 (N_2384,N_1815,N_2025);
xnor U2385 (N_2385,N_1882,N_2058);
nor U2386 (N_2386,N_1801,N_1828);
and U2387 (N_2387,N_2002,N_1820);
xnor U2388 (N_2388,N_2003,N_1816);
nand U2389 (N_2389,N_1982,N_1845);
or U2390 (N_2390,N_1883,N_1860);
or U2391 (N_2391,N_1965,N_1827);
and U2392 (N_2392,N_2092,N_2088);
xor U2393 (N_2393,N_1942,N_1890);
xnor U2394 (N_2394,N_1957,N_2051);
nor U2395 (N_2395,N_1949,N_1955);
nand U2396 (N_2396,N_1866,N_1925);
nand U2397 (N_2397,N_1844,N_2070);
nand U2398 (N_2398,N_2040,N_2031);
or U2399 (N_2399,N_1907,N_1964);
or U2400 (N_2400,N_2356,N_2145);
xnor U2401 (N_2401,N_2141,N_2261);
xnor U2402 (N_2402,N_2366,N_2334);
or U2403 (N_2403,N_2367,N_2355);
or U2404 (N_2404,N_2387,N_2287);
and U2405 (N_2405,N_2299,N_2307);
nand U2406 (N_2406,N_2330,N_2123);
or U2407 (N_2407,N_2276,N_2227);
nand U2408 (N_2408,N_2375,N_2247);
and U2409 (N_2409,N_2280,N_2328);
nand U2410 (N_2410,N_2369,N_2309);
or U2411 (N_2411,N_2115,N_2197);
or U2412 (N_2412,N_2170,N_2274);
or U2413 (N_2413,N_2198,N_2399);
or U2414 (N_2414,N_2228,N_2207);
nor U2415 (N_2415,N_2325,N_2353);
xor U2416 (N_2416,N_2386,N_2181);
or U2417 (N_2417,N_2351,N_2234);
xor U2418 (N_2418,N_2314,N_2229);
or U2419 (N_2419,N_2251,N_2200);
xor U2420 (N_2420,N_2180,N_2245);
or U2421 (N_2421,N_2297,N_2294);
nand U2422 (N_2422,N_2352,N_2102);
nor U2423 (N_2423,N_2390,N_2360);
and U2424 (N_2424,N_2184,N_2389);
xnor U2425 (N_2425,N_2370,N_2343);
nand U2426 (N_2426,N_2254,N_2174);
or U2427 (N_2427,N_2196,N_2110);
xnor U2428 (N_2428,N_2209,N_2371);
or U2429 (N_2429,N_2290,N_2154);
nand U2430 (N_2430,N_2277,N_2347);
xor U2431 (N_2431,N_2398,N_2288);
nand U2432 (N_2432,N_2226,N_2373);
nor U2433 (N_2433,N_2357,N_2124);
xor U2434 (N_2434,N_2150,N_2364);
or U2435 (N_2435,N_2383,N_2268);
and U2436 (N_2436,N_2361,N_2362);
xnor U2437 (N_2437,N_2354,N_2233);
nor U2438 (N_2438,N_2368,N_2295);
or U2439 (N_2439,N_2324,N_2376);
xnor U2440 (N_2440,N_2118,N_2281);
or U2441 (N_2441,N_2379,N_2250);
and U2442 (N_2442,N_2318,N_2240);
nor U2443 (N_2443,N_2338,N_2131);
nand U2444 (N_2444,N_2293,N_2291);
xnor U2445 (N_2445,N_2262,N_2103);
nor U2446 (N_2446,N_2193,N_2242);
nor U2447 (N_2447,N_2119,N_2265);
and U2448 (N_2448,N_2204,N_2199);
nor U2449 (N_2449,N_2125,N_2305);
xnor U2450 (N_2450,N_2231,N_2208);
and U2451 (N_2451,N_2216,N_2140);
nand U2452 (N_2452,N_2335,N_2313);
nand U2453 (N_2453,N_2302,N_2202);
nand U2454 (N_2454,N_2310,N_2165);
or U2455 (N_2455,N_2134,N_2378);
xor U2456 (N_2456,N_2253,N_2126);
nand U2457 (N_2457,N_2363,N_2256);
and U2458 (N_2458,N_2358,N_2116);
or U2459 (N_2459,N_2215,N_2139);
xnor U2460 (N_2460,N_2339,N_2206);
nand U2461 (N_2461,N_2286,N_2275);
nor U2462 (N_2462,N_2346,N_2201);
or U2463 (N_2463,N_2266,N_2223);
and U2464 (N_2464,N_2260,N_2169);
and U2465 (N_2465,N_2298,N_2185);
nor U2466 (N_2466,N_2127,N_2248);
or U2467 (N_2467,N_2108,N_2385);
nand U2468 (N_2468,N_2271,N_2306);
xnor U2469 (N_2469,N_2136,N_2349);
nand U2470 (N_2470,N_2388,N_2257);
or U2471 (N_2471,N_2188,N_2173);
xnor U2472 (N_2472,N_2301,N_2331);
xnor U2473 (N_2473,N_2192,N_2155);
xnor U2474 (N_2474,N_2267,N_2397);
and U2475 (N_2475,N_2393,N_2359);
nand U2476 (N_2476,N_2146,N_2241);
or U2477 (N_2477,N_2292,N_2382);
or U2478 (N_2478,N_2117,N_2308);
or U2479 (N_2479,N_2232,N_2342);
nand U2480 (N_2480,N_2168,N_2249);
nand U2481 (N_2481,N_2121,N_2273);
or U2482 (N_2482,N_2321,N_2323);
and U2483 (N_2483,N_2160,N_2135);
or U2484 (N_2484,N_2176,N_2164);
nor U2485 (N_2485,N_2300,N_2182);
and U2486 (N_2486,N_2104,N_2345);
and U2487 (N_2487,N_2317,N_2143);
xnor U2488 (N_2488,N_2320,N_2152);
nand U2489 (N_2489,N_2112,N_2244);
xnor U2490 (N_2490,N_2183,N_2279);
and U2491 (N_2491,N_2151,N_2237);
nand U2492 (N_2492,N_2189,N_2149);
xnor U2493 (N_2493,N_2327,N_2316);
xnor U2494 (N_2494,N_2270,N_2203);
and U2495 (N_2495,N_2350,N_2259);
xnor U2496 (N_2496,N_2289,N_2391);
nor U2497 (N_2497,N_2167,N_2144);
nand U2498 (N_2498,N_2341,N_2377);
or U2499 (N_2499,N_2264,N_2122);
xnor U2500 (N_2500,N_2381,N_2224);
or U2501 (N_2501,N_2282,N_2283);
or U2502 (N_2502,N_2120,N_2100);
and U2503 (N_2503,N_2396,N_2326);
xnor U2504 (N_2504,N_2285,N_2133);
and U2505 (N_2505,N_2148,N_2191);
nand U2506 (N_2506,N_2101,N_2372);
nand U2507 (N_2507,N_2315,N_2230);
xor U2508 (N_2508,N_2218,N_2222);
nor U2509 (N_2509,N_2304,N_2384);
and U2510 (N_2510,N_2137,N_2311);
nand U2511 (N_2511,N_2159,N_2132);
nand U2512 (N_2512,N_2220,N_2255);
and U2513 (N_2513,N_2178,N_2337);
nor U2514 (N_2514,N_2284,N_2344);
or U2515 (N_2515,N_2210,N_2172);
or U2516 (N_2516,N_2158,N_2312);
xor U2517 (N_2517,N_2194,N_2239);
or U2518 (N_2518,N_2161,N_2258);
or U2519 (N_2519,N_2106,N_2303);
xnor U2520 (N_2520,N_2153,N_2105);
nor U2521 (N_2521,N_2395,N_2340);
or U2522 (N_2522,N_2179,N_2157);
nor U2523 (N_2523,N_2336,N_2205);
or U2524 (N_2524,N_2211,N_2329);
xor U2525 (N_2525,N_2166,N_2190);
nand U2526 (N_2526,N_2219,N_2319);
or U2527 (N_2527,N_2225,N_2113);
nor U2528 (N_2528,N_2142,N_2156);
xor U2529 (N_2529,N_2128,N_2236);
xor U2530 (N_2530,N_2348,N_2187);
and U2531 (N_2531,N_2162,N_2322);
nor U2532 (N_2532,N_2392,N_2163);
and U2533 (N_2533,N_2114,N_2252);
nor U2534 (N_2534,N_2221,N_2130);
nor U2535 (N_2535,N_2278,N_2213);
nor U2536 (N_2536,N_2175,N_2235);
nand U2537 (N_2537,N_2111,N_2365);
and U2538 (N_2538,N_2246,N_2394);
xnor U2539 (N_2539,N_2374,N_2214);
nor U2540 (N_2540,N_2269,N_2186);
xor U2541 (N_2541,N_2217,N_2195);
nor U2542 (N_2542,N_2296,N_2109);
and U2543 (N_2543,N_2272,N_2129);
and U2544 (N_2544,N_2243,N_2212);
or U2545 (N_2545,N_2147,N_2332);
nor U2546 (N_2546,N_2263,N_2171);
nand U2547 (N_2547,N_2107,N_2138);
nor U2548 (N_2548,N_2238,N_2380);
nor U2549 (N_2549,N_2177,N_2333);
nand U2550 (N_2550,N_2109,N_2234);
nor U2551 (N_2551,N_2158,N_2341);
and U2552 (N_2552,N_2360,N_2139);
xor U2553 (N_2553,N_2195,N_2230);
nand U2554 (N_2554,N_2234,N_2398);
xnor U2555 (N_2555,N_2358,N_2214);
and U2556 (N_2556,N_2101,N_2364);
nand U2557 (N_2557,N_2251,N_2273);
or U2558 (N_2558,N_2236,N_2339);
nand U2559 (N_2559,N_2316,N_2295);
or U2560 (N_2560,N_2287,N_2123);
or U2561 (N_2561,N_2284,N_2355);
and U2562 (N_2562,N_2304,N_2334);
nor U2563 (N_2563,N_2281,N_2323);
or U2564 (N_2564,N_2224,N_2341);
and U2565 (N_2565,N_2104,N_2149);
xor U2566 (N_2566,N_2119,N_2390);
nand U2567 (N_2567,N_2397,N_2259);
nand U2568 (N_2568,N_2219,N_2332);
or U2569 (N_2569,N_2204,N_2187);
and U2570 (N_2570,N_2323,N_2388);
or U2571 (N_2571,N_2324,N_2293);
nand U2572 (N_2572,N_2302,N_2259);
and U2573 (N_2573,N_2333,N_2172);
nor U2574 (N_2574,N_2326,N_2279);
and U2575 (N_2575,N_2358,N_2352);
xnor U2576 (N_2576,N_2211,N_2327);
nor U2577 (N_2577,N_2372,N_2301);
or U2578 (N_2578,N_2334,N_2204);
nor U2579 (N_2579,N_2365,N_2243);
nor U2580 (N_2580,N_2349,N_2187);
or U2581 (N_2581,N_2294,N_2285);
and U2582 (N_2582,N_2187,N_2199);
and U2583 (N_2583,N_2224,N_2273);
xnor U2584 (N_2584,N_2166,N_2398);
xor U2585 (N_2585,N_2332,N_2226);
and U2586 (N_2586,N_2285,N_2323);
nand U2587 (N_2587,N_2383,N_2153);
or U2588 (N_2588,N_2212,N_2324);
or U2589 (N_2589,N_2102,N_2357);
nor U2590 (N_2590,N_2341,N_2324);
nand U2591 (N_2591,N_2261,N_2221);
or U2592 (N_2592,N_2272,N_2253);
xnor U2593 (N_2593,N_2211,N_2356);
and U2594 (N_2594,N_2151,N_2372);
or U2595 (N_2595,N_2162,N_2178);
or U2596 (N_2596,N_2168,N_2167);
xor U2597 (N_2597,N_2285,N_2385);
nor U2598 (N_2598,N_2363,N_2295);
or U2599 (N_2599,N_2265,N_2232);
nor U2600 (N_2600,N_2317,N_2352);
nor U2601 (N_2601,N_2386,N_2191);
xor U2602 (N_2602,N_2301,N_2158);
nor U2603 (N_2603,N_2364,N_2398);
nor U2604 (N_2604,N_2370,N_2155);
nor U2605 (N_2605,N_2157,N_2198);
nand U2606 (N_2606,N_2270,N_2129);
nand U2607 (N_2607,N_2366,N_2325);
or U2608 (N_2608,N_2272,N_2356);
nor U2609 (N_2609,N_2377,N_2263);
nor U2610 (N_2610,N_2120,N_2371);
nand U2611 (N_2611,N_2106,N_2168);
xor U2612 (N_2612,N_2210,N_2225);
xor U2613 (N_2613,N_2256,N_2110);
nor U2614 (N_2614,N_2391,N_2229);
nor U2615 (N_2615,N_2263,N_2149);
nand U2616 (N_2616,N_2389,N_2277);
and U2617 (N_2617,N_2149,N_2227);
nor U2618 (N_2618,N_2200,N_2241);
xor U2619 (N_2619,N_2205,N_2195);
or U2620 (N_2620,N_2387,N_2152);
nand U2621 (N_2621,N_2116,N_2374);
or U2622 (N_2622,N_2200,N_2391);
and U2623 (N_2623,N_2253,N_2172);
xnor U2624 (N_2624,N_2173,N_2129);
or U2625 (N_2625,N_2333,N_2146);
nand U2626 (N_2626,N_2144,N_2299);
xnor U2627 (N_2627,N_2302,N_2255);
xor U2628 (N_2628,N_2332,N_2205);
nor U2629 (N_2629,N_2284,N_2196);
nand U2630 (N_2630,N_2172,N_2214);
xor U2631 (N_2631,N_2178,N_2111);
or U2632 (N_2632,N_2326,N_2226);
or U2633 (N_2633,N_2311,N_2321);
xnor U2634 (N_2634,N_2212,N_2308);
or U2635 (N_2635,N_2346,N_2230);
nor U2636 (N_2636,N_2242,N_2337);
nor U2637 (N_2637,N_2189,N_2346);
nand U2638 (N_2638,N_2320,N_2130);
xor U2639 (N_2639,N_2190,N_2249);
nand U2640 (N_2640,N_2316,N_2356);
nand U2641 (N_2641,N_2119,N_2128);
or U2642 (N_2642,N_2271,N_2244);
and U2643 (N_2643,N_2207,N_2266);
or U2644 (N_2644,N_2130,N_2185);
xor U2645 (N_2645,N_2300,N_2379);
or U2646 (N_2646,N_2326,N_2143);
nand U2647 (N_2647,N_2216,N_2236);
nand U2648 (N_2648,N_2133,N_2130);
and U2649 (N_2649,N_2350,N_2267);
nand U2650 (N_2650,N_2272,N_2282);
nand U2651 (N_2651,N_2271,N_2398);
and U2652 (N_2652,N_2243,N_2186);
and U2653 (N_2653,N_2228,N_2331);
and U2654 (N_2654,N_2255,N_2198);
nand U2655 (N_2655,N_2207,N_2361);
or U2656 (N_2656,N_2317,N_2122);
xnor U2657 (N_2657,N_2253,N_2348);
and U2658 (N_2658,N_2365,N_2382);
and U2659 (N_2659,N_2132,N_2213);
xnor U2660 (N_2660,N_2185,N_2198);
or U2661 (N_2661,N_2336,N_2314);
or U2662 (N_2662,N_2119,N_2243);
or U2663 (N_2663,N_2328,N_2184);
nor U2664 (N_2664,N_2111,N_2374);
nand U2665 (N_2665,N_2311,N_2278);
xnor U2666 (N_2666,N_2302,N_2101);
and U2667 (N_2667,N_2101,N_2341);
nor U2668 (N_2668,N_2270,N_2329);
nor U2669 (N_2669,N_2281,N_2320);
or U2670 (N_2670,N_2369,N_2208);
xor U2671 (N_2671,N_2270,N_2147);
or U2672 (N_2672,N_2175,N_2156);
or U2673 (N_2673,N_2241,N_2316);
and U2674 (N_2674,N_2388,N_2347);
nor U2675 (N_2675,N_2124,N_2107);
nand U2676 (N_2676,N_2109,N_2257);
xnor U2677 (N_2677,N_2337,N_2190);
nor U2678 (N_2678,N_2388,N_2252);
nand U2679 (N_2679,N_2178,N_2210);
or U2680 (N_2680,N_2273,N_2223);
and U2681 (N_2681,N_2327,N_2234);
or U2682 (N_2682,N_2264,N_2128);
and U2683 (N_2683,N_2256,N_2131);
nor U2684 (N_2684,N_2112,N_2235);
and U2685 (N_2685,N_2236,N_2198);
or U2686 (N_2686,N_2388,N_2322);
nor U2687 (N_2687,N_2305,N_2273);
and U2688 (N_2688,N_2384,N_2158);
or U2689 (N_2689,N_2218,N_2229);
nor U2690 (N_2690,N_2172,N_2393);
xnor U2691 (N_2691,N_2327,N_2362);
and U2692 (N_2692,N_2227,N_2154);
xnor U2693 (N_2693,N_2290,N_2238);
xnor U2694 (N_2694,N_2131,N_2230);
nand U2695 (N_2695,N_2299,N_2359);
or U2696 (N_2696,N_2170,N_2245);
nor U2697 (N_2697,N_2150,N_2146);
and U2698 (N_2698,N_2342,N_2347);
nor U2699 (N_2699,N_2241,N_2236);
or U2700 (N_2700,N_2517,N_2647);
or U2701 (N_2701,N_2514,N_2583);
xnor U2702 (N_2702,N_2459,N_2485);
or U2703 (N_2703,N_2570,N_2548);
xnor U2704 (N_2704,N_2561,N_2539);
nand U2705 (N_2705,N_2653,N_2424);
and U2706 (N_2706,N_2553,N_2474);
or U2707 (N_2707,N_2496,N_2666);
nor U2708 (N_2708,N_2697,N_2693);
xnor U2709 (N_2709,N_2590,N_2630);
or U2710 (N_2710,N_2623,N_2461);
or U2711 (N_2711,N_2498,N_2420);
or U2712 (N_2712,N_2520,N_2457);
or U2713 (N_2713,N_2426,N_2511);
xnor U2714 (N_2714,N_2476,N_2628);
or U2715 (N_2715,N_2555,N_2542);
nand U2716 (N_2716,N_2413,N_2683);
nor U2717 (N_2717,N_2509,N_2617);
or U2718 (N_2718,N_2422,N_2594);
nand U2719 (N_2719,N_2691,N_2613);
nor U2720 (N_2720,N_2581,N_2421);
nor U2721 (N_2721,N_2659,N_2600);
nor U2722 (N_2722,N_2437,N_2680);
nor U2723 (N_2723,N_2547,N_2560);
nor U2724 (N_2724,N_2460,N_2602);
nand U2725 (N_2725,N_2595,N_2534);
nand U2726 (N_2726,N_2592,N_2569);
nor U2727 (N_2727,N_2652,N_2552);
or U2728 (N_2728,N_2451,N_2625);
and U2729 (N_2729,N_2657,N_2449);
xor U2730 (N_2730,N_2638,N_2528);
and U2731 (N_2731,N_2551,N_2438);
nand U2732 (N_2732,N_2502,N_2521);
or U2733 (N_2733,N_2470,N_2490);
and U2734 (N_2734,N_2486,N_2455);
or U2735 (N_2735,N_2417,N_2650);
or U2736 (N_2736,N_2596,N_2489);
nor U2737 (N_2737,N_2453,N_2563);
nor U2738 (N_2738,N_2444,N_2627);
and U2739 (N_2739,N_2436,N_2611);
or U2740 (N_2740,N_2448,N_2566);
nor U2741 (N_2741,N_2684,N_2546);
nor U2742 (N_2742,N_2568,N_2587);
nand U2743 (N_2743,N_2559,N_2523);
nor U2744 (N_2744,N_2504,N_2495);
and U2745 (N_2745,N_2649,N_2631);
xor U2746 (N_2746,N_2678,N_2688);
nor U2747 (N_2747,N_2527,N_2614);
nor U2748 (N_2748,N_2533,N_2440);
nand U2749 (N_2749,N_2400,N_2667);
and U2750 (N_2750,N_2624,N_2535);
and U2751 (N_2751,N_2418,N_2562);
nor U2752 (N_2752,N_2427,N_2526);
or U2753 (N_2753,N_2503,N_2419);
xor U2754 (N_2754,N_2501,N_2639);
nand U2755 (N_2755,N_2471,N_2519);
or U2756 (N_2756,N_2478,N_2597);
xnor U2757 (N_2757,N_2622,N_2513);
and U2758 (N_2758,N_2685,N_2518);
xnor U2759 (N_2759,N_2605,N_2441);
nor U2760 (N_2760,N_2468,N_2416);
and U2761 (N_2761,N_2507,N_2609);
nand U2762 (N_2762,N_2656,N_2598);
nor U2763 (N_2763,N_2682,N_2505);
and U2764 (N_2764,N_2512,N_2642);
xor U2765 (N_2765,N_2475,N_2402);
xnor U2766 (N_2766,N_2578,N_2644);
nor U2767 (N_2767,N_2607,N_2616);
nand U2768 (N_2768,N_2525,N_2536);
xor U2769 (N_2769,N_2557,N_2604);
nand U2770 (N_2770,N_2403,N_2465);
nand U2771 (N_2771,N_2589,N_2654);
and U2772 (N_2772,N_2698,N_2506);
nor U2773 (N_2773,N_2655,N_2425);
xnor U2774 (N_2774,N_2538,N_2483);
xnor U2775 (N_2775,N_2580,N_2433);
nand U2776 (N_2776,N_2524,N_2567);
nor U2777 (N_2777,N_2491,N_2549);
nor U2778 (N_2778,N_2544,N_2677);
xor U2779 (N_2779,N_2537,N_2522);
nor U2780 (N_2780,N_2577,N_2515);
or U2781 (N_2781,N_2676,N_2540);
nand U2782 (N_2782,N_2405,N_2637);
and U2783 (N_2783,N_2530,N_2477);
nor U2784 (N_2784,N_2550,N_2660);
or U2785 (N_2785,N_2454,N_2692);
or U2786 (N_2786,N_2414,N_2469);
and U2787 (N_2787,N_2482,N_2479);
nor U2788 (N_2788,N_2588,N_2410);
or U2789 (N_2789,N_2621,N_2447);
xor U2790 (N_2790,N_2634,N_2665);
and U2791 (N_2791,N_2442,N_2612);
nor U2792 (N_2792,N_2618,N_2664);
xnor U2793 (N_2793,N_2651,N_2599);
or U2794 (N_2794,N_2575,N_2565);
nor U2795 (N_2795,N_2584,N_2412);
nor U2796 (N_2796,N_2629,N_2661);
and U2797 (N_2797,N_2670,N_2432);
nor U2798 (N_2798,N_2543,N_2434);
or U2799 (N_2799,N_2593,N_2443);
or U2800 (N_2800,N_2579,N_2696);
and U2801 (N_2801,N_2462,N_2671);
and U2802 (N_2802,N_2669,N_2586);
or U2803 (N_2803,N_2699,N_2487);
and U2804 (N_2804,N_2480,N_2679);
or U2805 (N_2805,N_2633,N_2687);
nor U2806 (N_2806,N_2545,N_2508);
or U2807 (N_2807,N_2675,N_2658);
xor U2808 (N_2808,N_2641,N_2576);
nand U2809 (N_2809,N_2672,N_2632);
nand U2810 (N_2810,N_2415,N_2601);
and U2811 (N_2811,N_2564,N_2463);
nor U2812 (N_2812,N_2466,N_2408);
and U2813 (N_2813,N_2648,N_2431);
and U2814 (N_2814,N_2674,N_2686);
and U2815 (N_2815,N_2423,N_2516);
xor U2816 (N_2816,N_2406,N_2662);
nor U2817 (N_2817,N_2608,N_2429);
xor U2818 (N_2818,N_2481,N_2635);
xnor U2819 (N_2819,N_2458,N_2558);
or U2820 (N_2820,N_2493,N_2404);
or U2821 (N_2821,N_2541,N_2473);
nor U2822 (N_2822,N_2456,N_2556);
or U2823 (N_2823,N_2673,N_2554);
xnor U2824 (N_2824,N_2445,N_2467);
xor U2825 (N_2825,N_2572,N_2603);
xor U2826 (N_2826,N_2695,N_2446);
and U2827 (N_2827,N_2582,N_2636);
nor U2828 (N_2828,N_2407,N_2610);
or U2829 (N_2829,N_2439,N_2531);
xnor U2830 (N_2830,N_2646,N_2409);
or U2831 (N_2831,N_2573,N_2499);
xnor U2832 (N_2832,N_2450,N_2668);
nand U2833 (N_2833,N_2435,N_2497);
or U2834 (N_2834,N_2690,N_2452);
nor U2835 (N_2835,N_2500,N_2488);
and U2836 (N_2836,N_2472,N_2681);
nand U2837 (N_2837,N_2689,N_2529);
and U2838 (N_2838,N_2585,N_2619);
and U2839 (N_2839,N_2484,N_2492);
nand U2840 (N_2840,N_2620,N_2645);
or U2841 (N_2841,N_2615,N_2464);
nand U2842 (N_2842,N_2694,N_2643);
and U2843 (N_2843,N_2606,N_2428);
and U2844 (N_2844,N_2574,N_2430);
nor U2845 (N_2845,N_2401,N_2411);
xor U2846 (N_2846,N_2494,N_2663);
and U2847 (N_2847,N_2532,N_2626);
and U2848 (N_2848,N_2571,N_2510);
xnor U2849 (N_2849,N_2640,N_2591);
xor U2850 (N_2850,N_2627,N_2545);
nor U2851 (N_2851,N_2521,N_2699);
nor U2852 (N_2852,N_2401,N_2650);
nor U2853 (N_2853,N_2577,N_2459);
nand U2854 (N_2854,N_2523,N_2425);
or U2855 (N_2855,N_2645,N_2441);
and U2856 (N_2856,N_2578,N_2608);
xor U2857 (N_2857,N_2461,N_2666);
xnor U2858 (N_2858,N_2481,N_2515);
nor U2859 (N_2859,N_2593,N_2494);
nand U2860 (N_2860,N_2425,N_2466);
or U2861 (N_2861,N_2643,N_2696);
nor U2862 (N_2862,N_2626,N_2573);
nand U2863 (N_2863,N_2516,N_2402);
and U2864 (N_2864,N_2402,N_2473);
xor U2865 (N_2865,N_2490,N_2668);
or U2866 (N_2866,N_2433,N_2496);
xnor U2867 (N_2867,N_2431,N_2530);
nor U2868 (N_2868,N_2690,N_2417);
and U2869 (N_2869,N_2613,N_2417);
nor U2870 (N_2870,N_2596,N_2495);
nor U2871 (N_2871,N_2483,N_2404);
xor U2872 (N_2872,N_2407,N_2563);
and U2873 (N_2873,N_2483,N_2574);
or U2874 (N_2874,N_2533,N_2637);
or U2875 (N_2875,N_2676,N_2495);
nand U2876 (N_2876,N_2472,N_2582);
xnor U2877 (N_2877,N_2534,N_2696);
nand U2878 (N_2878,N_2646,N_2424);
xor U2879 (N_2879,N_2590,N_2466);
nand U2880 (N_2880,N_2465,N_2464);
and U2881 (N_2881,N_2405,N_2634);
nand U2882 (N_2882,N_2460,N_2628);
nand U2883 (N_2883,N_2465,N_2623);
and U2884 (N_2884,N_2623,N_2512);
nand U2885 (N_2885,N_2628,N_2411);
and U2886 (N_2886,N_2510,N_2472);
xnor U2887 (N_2887,N_2664,N_2686);
nor U2888 (N_2888,N_2545,N_2499);
or U2889 (N_2889,N_2404,N_2590);
and U2890 (N_2890,N_2528,N_2678);
nor U2891 (N_2891,N_2423,N_2575);
nand U2892 (N_2892,N_2550,N_2422);
xor U2893 (N_2893,N_2476,N_2620);
nor U2894 (N_2894,N_2488,N_2513);
and U2895 (N_2895,N_2625,N_2683);
and U2896 (N_2896,N_2552,N_2645);
and U2897 (N_2897,N_2627,N_2417);
xor U2898 (N_2898,N_2570,N_2544);
or U2899 (N_2899,N_2427,N_2698);
nor U2900 (N_2900,N_2583,N_2488);
nor U2901 (N_2901,N_2486,N_2438);
and U2902 (N_2902,N_2430,N_2485);
nand U2903 (N_2903,N_2507,N_2515);
and U2904 (N_2904,N_2536,N_2629);
nor U2905 (N_2905,N_2520,N_2518);
xnor U2906 (N_2906,N_2477,N_2417);
and U2907 (N_2907,N_2584,N_2426);
and U2908 (N_2908,N_2556,N_2526);
xnor U2909 (N_2909,N_2613,N_2693);
and U2910 (N_2910,N_2406,N_2413);
and U2911 (N_2911,N_2683,N_2470);
and U2912 (N_2912,N_2606,N_2645);
nor U2913 (N_2913,N_2571,N_2545);
and U2914 (N_2914,N_2465,N_2543);
nand U2915 (N_2915,N_2414,N_2470);
nand U2916 (N_2916,N_2631,N_2691);
xor U2917 (N_2917,N_2410,N_2632);
or U2918 (N_2918,N_2408,N_2422);
nand U2919 (N_2919,N_2569,N_2693);
xnor U2920 (N_2920,N_2416,N_2667);
xor U2921 (N_2921,N_2524,N_2534);
xor U2922 (N_2922,N_2543,N_2517);
nand U2923 (N_2923,N_2641,N_2637);
nor U2924 (N_2924,N_2615,N_2625);
xor U2925 (N_2925,N_2420,N_2688);
nor U2926 (N_2926,N_2529,N_2566);
and U2927 (N_2927,N_2670,N_2593);
nand U2928 (N_2928,N_2623,N_2631);
and U2929 (N_2929,N_2557,N_2418);
nor U2930 (N_2930,N_2478,N_2675);
xor U2931 (N_2931,N_2563,N_2693);
nor U2932 (N_2932,N_2446,N_2636);
nor U2933 (N_2933,N_2497,N_2489);
nor U2934 (N_2934,N_2552,N_2686);
xor U2935 (N_2935,N_2592,N_2482);
and U2936 (N_2936,N_2582,N_2584);
nand U2937 (N_2937,N_2628,N_2444);
nor U2938 (N_2938,N_2405,N_2669);
nor U2939 (N_2939,N_2667,N_2547);
xnor U2940 (N_2940,N_2582,N_2560);
nor U2941 (N_2941,N_2503,N_2671);
nor U2942 (N_2942,N_2433,N_2685);
nand U2943 (N_2943,N_2650,N_2469);
xnor U2944 (N_2944,N_2687,N_2497);
nand U2945 (N_2945,N_2425,N_2519);
nand U2946 (N_2946,N_2538,N_2641);
nand U2947 (N_2947,N_2538,N_2616);
xnor U2948 (N_2948,N_2563,N_2501);
or U2949 (N_2949,N_2470,N_2510);
xnor U2950 (N_2950,N_2656,N_2625);
xnor U2951 (N_2951,N_2522,N_2584);
and U2952 (N_2952,N_2448,N_2460);
nor U2953 (N_2953,N_2452,N_2683);
xnor U2954 (N_2954,N_2417,N_2656);
xor U2955 (N_2955,N_2695,N_2443);
nor U2956 (N_2956,N_2424,N_2633);
nor U2957 (N_2957,N_2579,N_2511);
xor U2958 (N_2958,N_2536,N_2550);
xnor U2959 (N_2959,N_2414,N_2661);
nor U2960 (N_2960,N_2666,N_2552);
or U2961 (N_2961,N_2695,N_2628);
and U2962 (N_2962,N_2668,N_2661);
nand U2963 (N_2963,N_2692,N_2539);
or U2964 (N_2964,N_2492,N_2698);
nor U2965 (N_2965,N_2526,N_2638);
xor U2966 (N_2966,N_2635,N_2461);
xnor U2967 (N_2967,N_2527,N_2699);
or U2968 (N_2968,N_2592,N_2559);
nor U2969 (N_2969,N_2637,N_2686);
nand U2970 (N_2970,N_2519,N_2537);
and U2971 (N_2971,N_2611,N_2497);
and U2972 (N_2972,N_2661,N_2691);
xnor U2973 (N_2973,N_2426,N_2452);
and U2974 (N_2974,N_2501,N_2445);
xnor U2975 (N_2975,N_2461,N_2427);
and U2976 (N_2976,N_2623,N_2581);
nand U2977 (N_2977,N_2491,N_2446);
xor U2978 (N_2978,N_2465,N_2606);
nand U2979 (N_2979,N_2647,N_2681);
nor U2980 (N_2980,N_2488,N_2609);
nor U2981 (N_2981,N_2650,N_2677);
and U2982 (N_2982,N_2674,N_2545);
nand U2983 (N_2983,N_2440,N_2415);
nand U2984 (N_2984,N_2664,N_2584);
xor U2985 (N_2985,N_2442,N_2647);
and U2986 (N_2986,N_2657,N_2560);
xor U2987 (N_2987,N_2448,N_2507);
or U2988 (N_2988,N_2553,N_2533);
or U2989 (N_2989,N_2404,N_2649);
nand U2990 (N_2990,N_2639,N_2554);
or U2991 (N_2991,N_2437,N_2635);
nor U2992 (N_2992,N_2427,N_2612);
nand U2993 (N_2993,N_2418,N_2682);
nand U2994 (N_2994,N_2682,N_2600);
and U2995 (N_2995,N_2579,N_2595);
and U2996 (N_2996,N_2670,N_2614);
or U2997 (N_2997,N_2469,N_2591);
xor U2998 (N_2998,N_2423,N_2612);
or U2999 (N_2999,N_2553,N_2531);
nand U3000 (N_3000,N_2798,N_2775);
nand U3001 (N_3001,N_2879,N_2981);
nand U3002 (N_3002,N_2866,N_2997);
nand U3003 (N_3003,N_2767,N_2794);
nor U3004 (N_3004,N_2954,N_2906);
and U3005 (N_3005,N_2855,N_2887);
nor U3006 (N_3006,N_2845,N_2863);
nor U3007 (N_3007,N_2894,N_2918);
or U3008 (N_3008,N_2849,N_2868);
nor U3009 (N_3009,N_2987,N_2967);
nand U3010 (N_3010,N_2992,N_2925);
or U3011 (N_3011,N_2742,N_2813);
xor U3012 (N_3012,N_2793,N_2755);
nor U3013 (N_3013,N_2764,N_2832);
or U3014 (N_3014,N_2938,N_2709);
xnor U3015 (N_3015,N_2984,N_2939);
nor U3016 (N_3016,N_2738,N_2723);
xnor U3017 (N_3017,N_2873,N_2920);
xor U3018 (N_3018,N_2808,N_2989);
and U3019 (N_3019,N_2715,N_2791);
or U3020 (N_3020,N_2747,N_2802);
nand U3021 (N_3021,N_2757,N_2736);
xnor U3022 (N_3022,N_2853,N_2896);
or U3023 (N_3023,N_2781,N_2864);
nand U3024 (N_3024,N_2702,N_2985);
nor U3025 (N_3025,N_2947,N_2986);
or U3026 (N_3026,N_2994,N_2842);
and U3027 (N_3027,N_2799,N_2850);
nand U3028 (N_3028,N_2903,N_2877);
xnor U3029 (N_3029,N_2725,N_2933);
xnor U3030 (N_3030,N_2858,N_2843);
xnor U3031 (N_3031,N_2979,N_2942);
nor U3032 (N_3032,N_2727,N_2988);
or U3033 (N_3033,N_2854,N_2834);
and U3034 (N_3034,N_2953,N_2885);
nand U3035 (N_3035,N_2883,N_2833);
or U3036 (N_3036,N_2905,N_2910);
xnor U3037 (N_3037,N_2851,N_2831);
or U3038 (N_3038,N_2932,N_2705);
nor U3039 (N_3039,N_2713,N_2810);
nor U3040 (N_3040,N_2991,N_2719);
nand U3041 (N_3041,N_2812,N_2968);
and U3042 (N_3042,N_2974,N_2919);
or U3043 (N_3043,N_2874,N_2957);
nand U3044 (N_3044,N_2745,N_2819);
nor U3045 (N_3045,N_2960,N_2839);
nand U3046 (N_3046,N_2733,N_2724);
and U3047 (N_3047,N_2941,N_2825);
nor U3048 (N_3048,N_2928,N_2912);
nand U3049 (N_3049,N_2886,N_2814);
nor U3050 (N_3050,N_2895,N_2970);
and U3051 (N_3051,N_2824,N_2720);
and U3052 (N_3052,N_2728,N_2703);
or U3053 (N_3053,N_2917,N_2870);
nor U3054 (N_3054,N_2800,N_2787);
and U3055 (N_3055,N_2721,N_2714);
nor U3056 (N_3056,N_2862,N_2948);
and U3057 (N_3057,N_2930,N_2888);
nand U3058 (N_3058,N_2935,N_2783);
and U3059 (N_3059,N_2828,N_2789);
nand U3060 (N_3060,N_2982,N_2878);
xnor U3061 (N_3061,N_2978,N_2993);
xor U3062 (N_3062,N_2766,N_2951);
xor U3063 (N_3063,N_2762,N_2729);
or U3064 (N_3064,N_2983,N_2712);
and U3065 (N_3065,N_2711,N_2772);
xor U3066 (N_3066,N_2759,N_2904);
nor U3067 (N_3067,N_2884,N_2803);
xnor U3068 (N_3068,N_2750,N_2922);
or U3069 (N_3069,N_2881,N_2990);
nor U3070 (N_3070,N_2784,N_2797);
xor U3071 (N_3071,N_2805,N_2893);
or U3072 (N_3072,N_2804,N_2908);
or U3073 (N_3073,N_2914,N_2734);
or U3074 (N_3074,N_2796,N_2753);
nor U3075 (N_3075,N_2934,N_2722);
and U3076 (N_3076,N_2786,N_2707);
nand U3077 (N_3077,N_2773,N_2963);
nor U3078 (N_3078,N_2741,N_2913);
and U3079 (N_3079,N_2717,N_2769);
nand U3080 (N_3080,N_2731,N_2876);
xor U3081 (N_3081,N_2859,N_2946);
nor U3082 (N_3082,N_2704,N_2971);
and U3083 (N_3083,N_2761,N_2836);
or U3084 (N_3084,N_2875,N_2861);
or U3085 (N_3085,N_2867,N_2763);
xor U3086 (N_3086,N_2776,N_2716);
nor U3087 (N_3087,N_2726,N_2902);
nand U3088 (N_3088,N_2737,N_2823);
xor U3089 (N_3089,N_2929,N_2980);
nor U3090 (N_3090,N_2740,N_2756);
nor U3091 (N_3091,N_2754,N_2923);
and U3092 (N_3092,N_2872,N_2785);
and U3093 (N_3093,N_2840,N_2961);
xnor U3094 (N_3094,N_2811,N_2846);
or U3095 (N_3095,N_2706,N_2901);
nor U3096 (N_3096,N_2771,N_2739);
nand U3097 (N_3097,N_2765,N_2807);
nor U3098 (N_3098,N_2749,N_2936);
xor U3099 (N_3099,N_2899,N_2860);
nand U3100 (N_3100,N_2848,N_2999);
nand U3101 (N_3101,N_2841,N_2826);
or U3102 (N_3102,N_2926,N_2821);
nand U3103 (N_3103,N_2829,N_2927);
nor U3104 (N_3104,N_2900,N_2950);
nor U3105 (N_3105,N_2897,N_2777);
xnor U3106 (N_3106,N_2952,N_2827);
nor U3107 (N_3107,N_2955,N_2898);
nor U3108 (N_3108,N_2795,N_2907);
and U3109 (N_3109,N_2958,N_2730);
or U3110 (N_3110,N_2890,N_2732);
and U3111 (N_3111,N_2998,N_2743);
nor U3112 (N_3112,N_2944,N_2820);
nor U3113 (N_3113,N_2931,N_2751);
xor U3114 (N_3114,N_2768,N_2770);
or U3115 (N_3115,N_2977,N_2915);
nor U3116 (N_3116,N_2882,N_2782);
or U3117 (N_3117,N_2937,N_2816);
nand U3118 (N_3118,N_2815,N_2744);
or U3119 (N_3119,N_2949,N_2966);
nand U3120 (N_3120,N_2889,N_2844);
xor U3121 (N_3121,N_2995,N_2774);
nand U3122 (N_3122,N_2809,N_2924);
xnor U3123 (N_3123,N_2973,N_2909);
nand U3124 (N_3124,N_2806,N_2700);
nor U3125 (N_3125,N_2801,N_2940);
nand U3126 (N_3126,N_2969,N_2911);
nand U3127 (N_3127,N_2838,N_2718);
and U3128 (N_3128,N_2792,N_2830);
xnor U3129 (N_3129,N_2943,N_2701);
xnor U3130 (N_3130,N_2778,N_2871);
and U3131 (N_3131,N_2964,N_2780);
or U3132 (N_3132,N_2972,N_2735);
and U3133 (N_3133,N_2996,N_2865);
nor U3134 (N_3134,N_2956,N_2760);
nor U3135 (N_3135,N_2891,N_2962);
xnor U3136 (N_3136,N_2746,N_2857);
nor U3137 (N_3137,N_2976,N_2869);
or U3138 (N_3138,N_2710,N_2758);
nor U3139 (N_3139,N_2880,N_2837);
xnor U3140 (N_3140,N_2965,N_2822);
xor U3141 (N_3141,N_2921,N_2847);
xor U3142 (N_3142,N_2817,N_2708);
or U3143 (N_3143,N_2945,N_2748);
or U3144 (N_3144,N_2779,N_2818);
nand U3145 (N_3145,N_2916,N_2892);
xnor U3146 (N_3146,N_2959,N_2835);
nor U3147 (N_3147,N_2790,N_2852);
nor U3148 (N_3148,N_2856,N_2788);
nand U3149 (N_3149,N_2752,N_2975);
nand U3150 (N_3150,N_2942,N_2927);
nand U3151 (N_3151,N_2896,N_2731);
and U3152 (N_3152,N_2905,N_2940);
xor U3153 (N_3153,N_2819,N_2843);
nand U3154 (N_3154,N_2993,N_2753);
or U3155 (N_3155,N_2770,N_2941);
nor U3156 (N_3156,N_2908,N_2917);
nand U3157 (N_3157,N_2907,N_2730);
and U3158 (N_3158,N_2813,N_2864);
xnor U3159 (N_3159,N_2999,N_2752);
and U3160 (N_3160,N_2825,N_2853);
nor U3161 (N_3161,N_2930,N_2882);
or U3162 (N_3162,N_2710,N_2986);
and U3163 (N_3163,N_2786,N_2884);
and U3164 (N_3164,N_2983,N_2706);
nor U3165 (N_3165,N_2855,N_2961);
nor U3166 (N_3166,N_2797,N_2973);
nand U3167 (N_3167,N_2979,N_2955);
and U3168 (N_3168,N_2947,N_2809);
nor U3169 (N_3169,N_2750,N_2943);
and U3170 (N_3170,N_2896,N_2707);
and U3171 (N_3171,N_2804,N_2894);
nand U3172 (N_3172,N_2868,N_2703);
or U3173 (N_3173,N_2939,N_2704);
xor U3174 (N_3174,N_2847,N_2976);
or U3175 (N_3175,N_2956,N_2994);
or U3176 (N_3176,N_2716,N_2919);
nor U3177 (N_3177,N_2761,N_2804);
nand U3178 (N_3178,N_2730,N_2879);
nand U3179 (N_3179,N_2948,N_2922);
nand U3180 (N_3180,N_2729,N_2960);
or U3181 (N_3181,N_2981,N_2702);
nor U3182 (N_3182,N_2885,N_2786);
xnor U3183 (N_3183,N_2924,N_2723);
or U3184 (N_3184,N_2748,N_2795);
and U3185 (N_3185,N_2839,N_2763);
nand U3186 (N_3186,N_2814,N_2859);
nand U3187 (N_3187,N_2728,N_2940);
or U3188 (N_3188,N_2768,N_2987);
nor U3189 (N_3189,N_2908,N_2820);
nand U3190 (N_3190,N_2751,N_2945);
or U3191 (N_3191,N_2982,N_2708);
or U3192 (N_3192,N_2896,N_2791);
nor U3193 (N_3193,N_2774,N_2904);
nand U3194 (N_3194,N_2747,N_2753);
nand U3195 (N_3195,N_2924,N_2738);
nand U3196 (N_3196,N_2795,N_2925);
and U3197 (N_3197,N_2718,N_2928);
or U3198 (N_3198,N_2899,N_2837);
nor U3199 (N_3199,N_2912,N_2926);
xor U3200 (N_3200,N_2924,N_2705);
and U3201 (N_3201,N_2956,N_2738);
or U3202 (N_3202,N_2787,N_2878);
nor U3203 (N_3203,N_2836,N_2913);
nor U3204 (N_3204,N_2958,N_2734);
xor U3205 (N_3205,N_2828,N_2826);
xor U3206 (N_3206,N_2859,N_2899);
nor U3207 (N_3207,N_2919,N_2918);
or U3208 (N_3208,N_2941,N_2821);
and U3209 (N_3209,N_2951,N_2787);
and U3210 (N_3210,N_2821,N_2831);
nor U3211 (N_3211,N_2913,N_2763);
nor U3212 (N_3212,N_2715,N_2894);
xnor U3213 (N_3213,N_2823,N_2769);
and U3214 (N_3214,N_2863,N_2892);
xor U3215 (N_3215,N_2883,N_2979);
or U3216 (N_3216,N_2840,N_2897);
xor U3217 (N_3217,N_2976,N_2767);
and U3218 (N_3218,N_2709,N_2846);
xor U3219 (N_3219,N_2893,N_2862);
and U3220 (N_3220,N_2861,N_2800);
and U3221 (N_3221,N_2887,N_2875);
nand U3222 (N_3222,N_2905,N_2760);
xor U3223 (N_3223,N_2761,N_2890);
nor U3224 (N_3224,N_2818,N_2874);
and U3225 (N_3225,N_2926,N_2814);
nor U3226 (N_3226,N_2932,N_2714);
nor U3227 (N_3227,N_2740,N_2963);
or U3228 (N_3228,N_2935,N_2752);
or U3229 (N_3229,N_2903,N_2825);
nor U3230 (N_3230,N_2876,N_2942);
nand U3231 (N_3231,N_2947,N_2888);
and U3232 (N_3232,N_2885,N_2715);
and U3233 (N_3233,N_2991,N_2718);
nor U3234 (N_3234,N_2860,N_2882);
or U3235 (N_3235,N_2963,N_2766);
and U3236 (N_3236,N_2973,N_2847);
nand U3237 (N_3237,N_2802,N_2955);
xor U3238 (N_3238,N_2862,N_2767);
nand U3239 (N_3239,N_2728,N_2878);
nor U3240 (N_3240,N_2890,N_2965);
nand U3241 (N_3241,N_2756,N_2822);
or U3242 (N_3242,N_2993,N_2844);
or U3243 (N_3243,N_2703,N_2918);
or U3244 (N_3244,N_2965,N_2776);
xor U3245 (N_3245,N_2783,N_2914);
xor U3246 (N_3246,N_2959,N_2853);
and U3247 (N_3247,N_2997,N_2776);
and U3248 (N_3248,N_2835,N_2838);
or U3249 (N_3249,N_2781,N_2825);
and U3250 (N_3250,N_2909,N_2819);
nand U3251 (N_3251,N_2927,N_2806);
and U3252 (N_3252,N_2724,N_2753);
nor U3253 (N_3253,N_2708,N_2921);
nor U3254 (N_3254,N_2839,N_2861);
and U3255 (N_3255,N_2826,N_2820);
xor U3256 (N_3256,N_2848,N_2995);
nand U3257 (N_3257,N_2907,N_2914);
or U3258 (N_3258,N_2752,N_2921);
or U3259 (N_3259,N_2804,N_2964);
nand U3260 (N_3260,N_2950,N_2815);
and U3261 (N_3261,N_2848,N_2812);
nor U3262 (N_3262,N_2883,N_2925);
nor U3263 (N_3263,N_2708,N_2991);
and U3264 (N_3264,N_2747,N_2995);
xor U3265 (N_3265,N_2763,N_2951);
nand U3266 (N_3266,N_2906,N_2828);
nor U3267 (N_3267,N_2842,N_2940);
nand U3268 (N_3268,N_2768,N_2810);
or U3269 (N_3269,N_2828,N_2712);
nor U3270 (N_3270,N_2944,N_2744);
nand U3271 (N_3271,N_2808,N_2735);
and U3272 (N_3272,N_2931,N_2747);
or U3273 (N_3273,N_2729,N_2935);
nand U3274 (N_3274,N_2991,N_2833);
or U3275 (N_3275,N_2933,N_2821);
nand U3276 (N_3276,N_2823,N_2879);
xor U3277 (N_3277,N_2701,N_2791);
xor U3278 (N_3278,N_2951,N_2781);
xnor U3279 (N_3279,N_2712,N_2744);
or U3280 (N_3280,N_2888,N_2966);
or U3281 (N_3281,N_2761,N_2992);
xor U3282 (N_3282,N_2839,N_2902);
nor U3283 (N_3283,N_2779,N_2702);
xor U3284 (N_3284,N_2865,N_2783);
xnor U3285 (N_3285,N_2965,N_2708);
or U3286 (N_3286,N_2968,N_2836);
xnor U3287 (N_3287,N_2714,N_2997);
xnor U3288 (N_3288,N_2744,N_2930);
nand U3289 (N_3289,N_2733,N_2722);
nand U3290 (N_3290,N_2846,N_2768);
nand U3291 (N_3291,N_2987,N_2900);
nor U3292 (N_3292,N_2861,N_2817);
nor U3293 (N_3293,N_2891,N_2814);
and U3294 (N_3294,N_2786,N_2952);
nor U3295 (N_3295,N_2747,N_2919);
nor U3296 (N_3296,N_2704,N_2739);
and U3297 (N_3297,N_2714,N_2788);
and U3298 (N_3298,N_2786,N_2767);
or U3299 (N_3299,N_2826,N_2726);
nor U3300 (N_3300,N_3038,N_3212);
and U3301 (N_3301,N_3261,N_3194);
or U3302 (N_3302,N_3168,N_3266);
nor U3303 (N_3303,N_3272,N_3230);
nand U3304 (N_3304,N_3264,N_3015);
and U3305 (N_3305,N_3258,N_3162);
nand U3306 (N_3306,N_3145,N_3196);
and U3307 (N_3307,N_3222,N_3044);
and U3308 (N_3308,N_3132,N_3218);
xor U3309 (N_3309,N_3270,N_3110);
xor U3310 (N_3310,N_3282,N_3062);
xor U3311 (N_3311,N_3241,N_3112);
xor U3312 (N_3312,N_3078,N_3281);
xor U3313 (N_3313,N_3036,N_3239);
xnor U3314 (N_3314,N_3126,N_3021);
nor U3315 (N_3315,N_3150,N_3224);
xnor U3316 (N_3316,N_3004,N_3048);
or U3317 (N_3317,N_3250,N_3231);
and U3318 (N_3318,N_3103,N_3170);
xor U3319 (N_3319,N_3268,N_3051);
nor U3320 (N_3320,N_3067,N_3167);
and U3321 (N_3321,N_3243,N_3041);
nand U3322 (N_3322,N_3293,N_3244);
and U3323 (N_3323,N_3101,N_3122);
xnor U3324 (N_3324,N_3057,N_3135);
and U3325 (N_3325,N_3013,N_3107);
nor U3326 (N_3326,N_3260,N_3269);
or U3327 (N_3327,N_3134,N_3081);
nor U3328 (N_3328,N_3257,N_3275);
xor U3329 (N_3329,N_3207,N_3031);
or U3330 (N_3330,N_3007,N_3087);
and U3331 (N_3331,N_3117,N_3287);
nor U3332 (N_3332,N_3032,N_3164);
nor U3333 (N_3333,N_3027,N_3128);
or U3334 (N_3334,N_3156,N_3193);
or U3335 (N_3335,N_3034,N_3129);
or U3336 (N_3336,N_3183,N_3157);
xnor U3337 (N_3337,N_3095,N_3137);
xnor U3338 (N_3338,N_3277,N_3182);
nor U3339 (N_3339,N_3197,N_3178);
or U3340 (N_3340,N_3200,N_3173);
and U3341 (N_3341,N_3104,N_3166);
xnor U3342 (N_3342,N_3047,N_3221);
nor U3343 (N_3343,N_3203,N_3232);
nand U3344 (N_3344,N_3094,N_3001);
nor U3345 (N_3345,N_3151,N_3235);
and U3346 (N_3346,N_3210,N_3071);
or U3347 (N_3347,N_3248,N_3204);
xor U3348 (N_3348,N_3090,N_3070);
nor U3349 (N_3349,N_3003,N_3100);
and U3350 (N_3350,N_3080,N_3017);
or U3351 (N_3351,N_3180,N_3050);
or U3352 (N_3352,N_3000,N_3160);
and U3353 (N_3353,N_3278,N_3176);
xnor U3354 (N_3354,N_3147,N_3082);
and U3355 (N_3355,N_3109,N_3133);
nor U3356 (N_3356,N_3064,N_3143);
xor U3357 (N_3357,N_3014,N_3102);
xnor U3358 (N_3358,N_3208,N_3121);
nor U3359 (N_3359,N_3296,N_3020);
nand U3360 (N_3360,N_3083,N_3024);
and U3361 (N_3361,N_3019,N_3002);
xnor U3362 (N_3362,N_3063,N_3115);
nor U3363 (N_3363,N_3053,N_3079);
nor U3364 (N_3364,N_3220,N_3215);
or U3365 (N_3365,N_3255,N_3025);
and U3366 (N_3366,N_3205,N_3219);
nor U3367 (N_3367,N_3273,N_3154);
nand U3368 (N_3368,N_3245,N_3238);
or U3369 (N_3369,N_3247,N_3012);
and U3370 (N_3370,N_3234,N_3276);
nor U3371 (N_3371,N_3185,N_3075);
and U3372 (N_3372,N_3256,N_3184);
and U3373 (N_3373,N_3190,N_3165);
xor U3374 (N_3374,N_3130,N_3259);
nand U3375 (N_3375,N_3213,N_3052);
and U3376 (N_3376,N_3280,N_3141);
or U3377 (N_3377,N_3274,N_3123);
xor U3378 (N_3378,N_3199,N_3227);
and U3379 (N_3379,N_3285,N_3217);
xor U3380 (N_3380,N_3005,N_3120);
xnor U3381 (N_3381,N_3069,N_3127);
xnor U3382 (N_3382,N_3174,N_3061);
or U3383 (N_3383,N_3189,N_3091);
nand U3384 (N_3384,N_3265,N_3073);
xor U3385 (N_3385,N_3179,N_3116);
or U3386 (N_3386,N_3253,N_3099);
and U3387 (N_3387,N_3271,N_3295);
or U3388 (N_3388,N_3254,N_3225);
nand U3389 (N_3389,N_3049,N_3098);
nand U3390 (N_3390,N_3028,N_3035);
nand U3391 (N_3391,N_3169,N_3089);
xor U3392 (N_3392,N_3092,N_3066);
and U3393 (N_3393,N_3148,N_3186);
nand U3394 (N_3394,N_3125,N_3009);
nand U3395 (N_3395,N_3188,N_3046);
nor U3396 (N_3396,N_3022,N_3142);
xor U3397 (N_3397,N_3093,N_3131);
and U3398 (N_3398,N_3292,N_3263);
or U3399 (N_3399,N_3056,N_3010);
xor U3400 (N_3400,N_3045,N_3113);
xor U3401 (N_3401,N_3290,N_3267);
or U3402 (N_3402,N_3201,N_3140);
or U3403 (N_3403,N_3262,N_3175);
and U3404 (N_3404,N_3181,N_3202);
nor U3405 (N_3405,N_3139,N_3249);
nand U3406 (N_3406,N_3136,N_3055);
nor U3407 (N_3407,N_3018,N_3153);
nor U3408 (N_3408,N_3294,N_3054);
nand U3409 (N_3409,N_3299,N_3237);
and U3410 (N_3410,N_3223,N_3240);
nand U3411 (N_3411,N_3086,N_3043);
nand U3412 (N_3412,N_3172,N_3152);
xor U3413 (N_3413,N_3298,N_3008);
xnor U3414 (N_3414,N_3149,N_3072);
nand U3415 (N_3415,N_3233,N_3088);
and U3416 (N_3416,N_3216,N_3029);
nand U3417 (N_3417,N_3195,N_3163);
xor U3418 (N_3418,N_3096,N_3059);
nand U3419 (N_3419,N_3037,N_3206);
and U3420 (N_3420,N_3108,N_3286);
xnor U3421 (N_3421,N_3279,N_3026);
xor U3422 (N_3422,N_3283,N_3144);
and U3423 (N_3423,N_3191,N_3118);
xor U3424 (N_3424,N_3074,N_3119);
nor U3425 (N_3425,N_3161,N_3146);
and U3426 (N_3426,N_3016,N_3097);
xnor U3427 (N_3427,N_3209,N_3229);
or U3428 (N_3428,N_3158,N_3284);
and U3429 (N_3429,N_3011,N_3077);
or U3430 (N_3430,N_3076,N_3006);
nand U3431 (N_3431,N_3171,N_3060);
and U3432 (N_3432,N_3023,N_3068);
nor U3433 (N_3433,N_3040,N_3198);
nor U3434 (N_3434,N_3033,N_3030);
nand U3435 (N_3435,N_3251,N_3106);
nand U3436 (N_3436,N_3288,N_3114);
nor U3437 (N_3437,N_3246,N_3226);
or U3438 (N_3438,N_3042,N_3211);
nor U3439 (N_3439,N_3291,N_3177);
xnor U3440 (N_3440,N_3192,N_3105);
nand U3441 (N_3441,N_3155,N_3058);
xnor U3442 (N_3442,N_3236,N_3084);
xnor U3443 (N_3443,N_3039,N_3138);
or U3444 (N_3444,N_3228,N_3159);
xnor U3445 (N_3445,N_3252,N_3297);
or U3446 (N_3446,N_3124,N_3085);
nand U3447 (N_3447,N_3242,N_3065);
or U3448 (N_3448,N_3111,N_3187);
nand U3449 (N_3449,N_3214,N_3289);
and U3450 (N_3450,N_3286,N_3123);
or U3451 (N_3451,N_3142,N_3260);
nand U3452 (N_3452,N_3290,N_3093);
or U3453 (N_3453,N_3145,N_3107);
xor U3454 (N_3454,N_3287,N_3064);
nand U3455 (N_3455,N_3042,N_3012);
xnor U3456 (N_3456,N_3102,N_3222);
nor U3457 (N_3457,N_3105,N_3274);
and U3458 (N_3458,N_3233,N_3108);
nand U3459 (N_3459,N_3231,N_3090);
nor U3460 (N_3460,N_3081,N_3128);
and U3461 (N_3461,N_3251,N_3228);
and U3462 (N_3462,N_3256,N_3143);
nor U3463 (N_3463,N_3126,N_3230);
and U3464 (N_3464,N_3039,N_3008);
nand U3465 (N_3465,N_3274,N_3159);
nand U3466 (N_3466,N_3256,N_3158);
and U3467 (N_3467,N_3108,N_3064);
or U3468 (N_3468,N_3096,N_3252);
xnor U3469 (N_3469,N_3213,N_3084);
nand U3470 (N_3470,N_3162,N_3077);
nand U3471 (N_3471,N_3035,N_3007);
nor U3472 (N_3472,N_3088,N_3105);
and U3473 (N_3473,N_3011,N_3203);
nand U3474 (N_3474,N_3074,N_3030);
and U3475 (N_3475,N_3011,N_3279);
xor U3476 (N_3476,N_3184,N_3043);
nor U3477 (N_3477,N_3232,N_3010);
nand U3478 (N_3478,N_3093,N_3281);
nand U3479 (N_3479,N_3025,N_3159);
nor U3480 (N_3480,N_3131,N_3288);
nor U3481 (N_3481,N_3051,N_3176);
and U3482 (N_3482,N_3214,N_3201);
xnor U3483 (N_3483,N_3056,N_3120);
xor U3484 (N_3484,N_3114,N_3220);
and U3485 (N_3485,N_3095,N_3132);
or U3486 (N_3486,N_3197,N_3082);
or U3487 (N_3487,N_3048,N_3231);
nor U3488 (N_3488,N_3286,N_3107);
and U3489 (N_3489,N_3103,N_3048);
nand U3490 (N_3490,N_3144,N_3258);
or U3491 (N_3491,N_3083,N_3264);
nand U3492 (N_3492,N_3232,N_3032);
and U3493 (N_3493,N_3191,N_3207);
xnor U3494 (N_3494,N_3001,N_3083);
nor U3495 (N_3495,N_3151,N_3089);
xor U3496 (N_3496,N_3090,N_3216);
or U3497 (N_3497,N_3003,N_3259);
nand U3498 (N_3498,N_3011,N_3228);
xnor U3499 (N_3499,N_3187,N_3019);
nand U3500 (N_3500,N_3128,N_3133);
and U3501 (N_3501,N_3072,N_3008);
nor U3502 (N_3502,N_3001,N_3037);
xnor U3503 (N_3503,N_3084,N_3297);
xnor U3504 (N_3504,N_3192,N_3110);
nor U3505 (N_3505,N_3118,N_3088);
and U3506 (N_3506,N_3205,N_3188);
or U3507 (N_3507,N_3181,N_3211);
or U3508 (N_3508,N_3111,N_3186);
nand U3509 (N_3509,N_3115,N_3200);
or U3510 (N_3510,N_3053,N_3138);
nor U3511 (N_3511,N_3105,N_3082);
or U3512 (N_3512,N_3125,N_3169);
nand U3513 (N_3513,N_3233,N_3186);
nor U3514 (N_3514,N_3232,N_3062);
and U3515 (N_3515,N_3168,N_3293);
nor U3516 (N_3516,N_3161,N_3277);
and U3517 (N_3517,N_3074,N_3070);
nor U3518 (N_3518,N_3149,N_3123);
nand U3519 (N_3519,N_3048,N_3023);
and U3520 (N_3520,N_3271,N_3299);
xnor U3521 (N_3521,N_3064,N_3025);
or U3522 (N_3522,N_3233,N_3289);
nor U3523 (N_3523,N_3005,N_3231);
xor U3524 (N_3524,N_3120,N_3161);
or U3525 (N_3525,N_3255,N_3121);
and U3526 (N_3526,N_3295,N_3134);
or U3527 (N_3527,N_3022,N_3146);
and U3528 (N_3528,N_3019,N_3026);
nand U3529 (N_3529,N_3087,N_3105);
or U3530 (N_3530,N_3283,N_3009);
or U3531 (N_3531,N_3013,N_3102);
nor U3532 (N_3532,N_3197,N_3188);
nor U3533 (N_3533,N_3295,N_3133);
or U3534 (N_3534,N_3158,N_3244);
xnor U3535 (N_3535,N_3288,N_3111);
nor U3536 (N_3536,N_3017,N_3031);
nor U3537 (N_3537,N_3289,N_3222);
or U3538 (N_3538,N_3214,N_3117);
and U3539 (N_3539,N_3027,N_3257);
nand U3540 (N_3540,N_3165,N_3293);
or U3541 (N_3541,N_3186,N_3273);
nand U3542 (N_3542,N_3284,N_3087);
and U3543 (N_3543,N_3033,N_3247);
and U3544 (N_3544,N_3126,N_3242);
or U3545 (N_3545,N_3150,N_3270);
nand U3546 (N_3546,N_3201,N_3114);
xor U3547 (N_3547,N_3186,N_3045);
and U3548 (N_3548,N_3249,N_3050);
nor U3549 (N_3549,N_3186,N_3150);
and U3550 (N_3550,N_3198,N_3144);
or U3551 (N_3551,N_3212,N_3297);
nor U3552 (N_3552,N_3195,N_3024);
and U3553 (N_3553,N_3098,N_3162);
nor U3554 (N_3554,N_3145,N_3186);
xnor U3555 (N_3555,N_3237,N_3137);
or U3556 (N_3556,N_3213,N_3002);
nand U3557 (N_3557,N_3216,N_3260);
or U3558 (N_3558,N_3183,N_3166);
or U3559 (N_3559,N_3126,N_3223);
nor U3560 (N_3560,N_3211,N_3216);
nand U3561 (N_3561,N_3239,N_3133);
and U3562 (N_3562,N_3160,N_3133);
xnor U3563 (N_3563,N_3030,N_3295);
nand U3564 (N_3564,N_3174,N_3027);
nand U3565 (N_3565,N_3107,N_3293);
xor U3566 (N_3566,N_3231,N_3108);
nand U3567 (N_3567,N_3290,N_3040);
nand U3568 (N_3568,N_3256,N_3157);
and U3569 (N_3569,N_3162,N_3209);
and U3570 (N_3570,N_3192,N_3156);
nor U3571 (N_3571,N_3083,N_3106);
xnor U3572 (N_3572,N_3032,N_3203);
nor U3573 (N_3573,N_3108,N_3201);
nand U3574 (N_3574,N_3131,N_3272);
and U3575 (N_3575,N_3234,N_3055);
and U3576 (N_3576,N_3009,N_3274);
nor U3577 (N_3577,N_3269,N_3156);
or U3578 (N_3578,N_3273,N_3112);
nor U3579 (N_3579,N_3145,N_3073);
nand U3580 (N_3580,N_3213,N_3189);
xor U3581 (N_3581,N_3067,N_3187);
and U3582 (N_3582,N_3095,N_3029);
nand U3583 (N_3583,N_3221,N_3248);
and U3584 (N_3584,N_3025,N_3253);
or U3585 (N_3585,N_3123,N_3053);
and U3586 (N_3586,N_3254,N_3196);
nand U3587 (N_3587,N_3080,N_3185);
nor U3588 (N_3588,N_3157,N_3004);
and U3589 (N_3589,N_3058,N_3174);
or U3590 (N_3590,N_3170,N_3276);
or U3591 (N_3591,N_3055,N_3264);
and U3592 (N_3592,N_3171,N_3102);
and U3593 (N_3593,N_3147,N_3228);
and U3594 (N_3594,N_3064,N_3268);
and U3595 (N_3595,N_3285,N_3229);
and U3596 (N_3596,N_3263,N_3190);
or U3597 (N_3597,N_3002,N_3158);
and U3598 (N_3598,N_3272,N_3196);
xor U3599 (N_3599,N_3168,N_3260);
and U3600 (N_3600,N_3325,N_3446);
xor U3601 (N_3601,N_3508,N_3456);
nor U3602 (N_3602,N_3420,N_3386);
nand U3603 (N_3603,N_3582,N_3462);
nor U3604 (N_3604,N_3577,N_3583);
and U3605 (N_3605,N_3348,N_3337);
and U3606 (N_3606,N_3564,N_3320);
nand U3607 (N_3607,N_3436,N_3532);
nand U3608 (N_3608,N_3485,N_3306);
xnor U3609 (N_3609,N_3424,N_3598);
nand U3610 (N_3610,N_3563,N_3355);
nand U3611 (N_3611,N_3599,N_3341);
xor U3612 (N_3612,N_3472,N_3552);
nand U3613 (N_3613,N_3385,N_3499);
nand U3614 (N_3614,N_3498,N_3595);
and U3615 (N_3615,N_3489,N_3407);
xnor U3616 (N_3616,N_3584,N_3486);
or U3617 (N_3617,N_3468,N_3345);
nor U3618 (N_3618,N_3309,N_3321);
and U3619 (N_3619,N_3349,N_3529);
xnor U3620 (N_3620,N_3568,N_3570);
xnor U3621 (N_3621,N_3578,N_3557);
or U3622 (N_3622,N_3562,N_3537);
and U3623 (N_3623,N_3504,N_3482);
nor U3624 (N_3624,N_3470,N_3343);
nand U3625 (N_3625,N_3512,N_3413);
nand U3626 (N_3626,N_3567,N_3402);
and U3627 (N_3627,N_3412,N_3597);
nand U3628 (N_3628,N_3364,N_3590);
and U3629 (N_3629,N_3330,N_3459);
nor U3630 (N_3630,N_3387,N_3332);
or U3631 (N_3631,N_3594,N_3353);
nor U3632 (N_3632,N_3319,N_3535);
or U3633 (N_3633,N_3440,N_3521);
nor U3634 (N_3634,N_3558,N_3536);
nor U3635 (N_3635,N_3515,N_3315);
xor U3636 (N_3636,N_3447,N_3548);
and U3637 (N_3637,N_3547,N_3333);
xnor U3638 (N_3638,N_3403,N_3464);
and U3639 (N_3639,N_3494,N_3352);
nand U3640 (N_3640,N_3488,N_3540);
nor U3641 (N_3641,N_3369,N_3549);
nor U3642 (N_3642,N_3399,N_3372);
or U3643 (N_3643,N_3560,N_3452);
nor U3644 (N_3644,N_3383,N_3373);
and U3645 (N_3645,N_3398,N_3401);
xnor U3646 (N_3646,N_3382,N_3551);
or U3647 (N_3647,N_3493,N_3334);
nand U3648 (N_3648,N_3395,N_3545);
or U3649 (N_3649,N_3307,N_3469);
or U3650 (N_3650,N_3565,N_3311);
or U3651 (N_3651,N_3411,N_3396);
nor U3652 (N_3652,N_3408,N_3495);
nand U3653 (N_3653,N_3439,N_3342);
or U3654 (N_3654,N_3528,N_3581);
or U3655 (N_3655,N_3335,N_3429);
xor U3656 (N_3656,N_3478,N_3410);
and U3657 (N_3657,N_3354,N_3514);
and U3658 (N_3658,N_3454,N_3326);
and U3659 (N_3659,N_3397,N_3517);
and U3660 (N_3660,N_3390,N_3530);
nor U3661 (N_3661,N_3338,N_3520);
nand U3662 (N_3662,N_3585,N_3487);
and U3663 (N_3663,N_3465,N_3384);
and U3664 (N_3664,N_3592,N_3451);
nor U3665 (N_3665,N_3400,N_3308);
xor U3666 (N_3666,N_3448,N_3550);
nand U3667 (N_3667,N_3365,N_3575);
xor U3668 (N_3668,N_3531,N_3339);
nor U3669 (N_3669,N_3303,N_3479);
nor U3670 (N_3670,N_3589,N_3357);
nor U3671 (N_3671,N_3449,N_3404);
nor U3672 (N_3672,N_3414,N_3313);
nor U3673 (N_3673,N_3358,N_3432);
nand U3674 (N_3674,N_3300,N_3302);
or U3675 (N_3675,N_3458,N_3490);
and U3676 (N_3676,N_3476,N_3546);
nand U3677 (N_3677,N_3324,N_3501);
nor U3678 (N_3678,N_3569,N_3511);
or U3679 (N_3679,N_3572,N_3375);
nor U3680 (N_3680,N_3463,N_3312);
nand U3681 (N_3681,N_3496,N_3561);
and U3682 (N_3682,N_3559,N_3474);
nand U3683 (N_3683,N_3331,N_3393);
nand U3684 (N_3684,N_3327,N_3344);
and U3685 (N_3685,N_3427,N_3475);
and U3686 (N_3686,N_3450,N_3444);
xor U3687 (N_3687,N_3510,N_3576);
nand U3688 (N_3688,N_3310,N_3428);
and U3689 (N_3689,N_3418,N_3363);
and U3690 (N_3690,N_3359,N_3519);
or U3691 (N_3691,N_3457,N_3322);
xnor U3692 (N_3692,N_3417,N_3502);
xnor U3693 (N_3693,N_3588,N_3347);
or U3694 (N_3694,N_3571,N_3461);
and U3695 (N_3695,N_3453,N_3316);
or U3696 (N_3696,N_3527,N_3368);
xor U3697 (N_3697,N_3361,N_3574);
or U3698 (N_3698,N_3304,N_3433);
and U3699 (N_3699,N_3522,N_3591);
nand U3700 (N_3700,N_3544,N_3445);
or U3701 (N_3701,N_3409,N_3497);
and U3702 (N_3702,N_3441,N_3370);
or U3703 (N_3703,N_3430,N_3534);
or U3704 (N_3704,N_3415,N_3467);
xnor U3705 (N_3705,N_3329,N_3518);
nor U3706 (N_3706,N_3406,N_3305);
nand U3707 (N_3707,N_3523,N_3351);
or U3708 (N_3708,N_3380,N_3513);
nor U3709 (N_3709,N_3422,N_3481);
xnor U3710 (N_3710,N_3438,N_3500);
nand U3711 (N_3711,N_3483,N_3317);
and U3712 (N_3712,N_3538,N_3516);
xnor U3713 (N_3713,N_3503,N_3477);
nor U3714 (N_3714,N_3423,N_3466);
and U3715 (N_3715,N_3542,N_3376);
nor U3716 (N_3716,N_3431,N_3471);
nor U3717 (N_3717,N_3573,N_3323);
and U3718 (N_3718,N_3378,N_3318);
and U3719 (N_3719,N_3533,N_3555);
xor U3720 (N_3720,N_3443,N_3377);
nor U3721 (N_3721,N_3426,N_3491);
and U3722 (N_3722,N_3596,N_3525);
and U3723 (N_3723,N_3526,N_3336);
nor U3724 (N_3724,N_3371,N_3541);
nor U3725 (N_3725,N_3435,N_3473);
or U3726 (N_3726,N_3379,N_3374);
and U3727 (N_3727,N_3593,N_3346);
nor U3728 (N_3728,N_3460,N_3442);
nor U3729 (N_3729,N_3554,N_3566);
xor U3730 (N_3730,N_3492,N_3389);
xnor U3731 (N_3731,N_3362,N_3553);
and U3732 (N_3732,N_3437,N_3421);
or U3733 (N_3733,N_3419,N_3580);
xnor U3734 (N_3734,N_3509,N_3350);
nor U3735 (N_3735,N_3328,N_3556);
xor U3736 (N_3736,N_3586,N_3301);
nor U3737 (N_3737,N_3484,N_3366);
xnor U3738 (N_3738,N_3367,N_3434);
nand U3739 (N_3739,N_3425,N_3507);
or U3740 (N_3740,N_3405,N_3506);
or U3741 (N_3741,N_3381,N_3480);
and U3742 (N_3742,N_3360,N_3579);
and U3743 (N_3743,N_3340,N_3356);
nor U3744 (N_3744,N_3524,N_3416);
or U3745 (N_3745,N_3394,N_3391);
xor U3746 (N_3746,N_3587,N_3392);
nor U3747 (N_3747,N_3314,N_3539);
nand U3748 (N_3748,N_3543,N_3505);
xnor U3749 (N_3749,N_3455,N_3388);
and U3750 (N_3750,N_3598,N_3495);
xor U3751 (N_3751,N_3344,N_3490);
or U3752 (N_3752,N_3462,N_3571);
or U3753 (N_3753,N_3464,N_3314);
nand U3754 (N_3754,N_3446,N_3566);
xor U3755 (N_3755,N_3338,N_3570);
xor U3756 (N_3756,N_3567,N_3541);
xnor U3757 (N_3757,N_3385,N_3527);
nand U3758 (N_3758,N_3471,N_3487);
and U3759 (N_3759,N_3470,N_3477);
nand U3760 (N_3760,N_3435,N_3320);
xnor U3761 (N_3761,N_3546,N_3459);
nor U3762 (N_3762,N_3542,N_3397);
and U3763 (N_3763,N_3524,N_3430);
or U3764 (N_3764,N_3564,N_3538);
nand U3765 (N_3765,N_3511,N_3490);
xnor U3766 (N_3766,N_3465,N_3588);
xor U3767 (N_3767,N_3594,N_3503);
xnor U3768 (N_3768,N_3428,N_3412);
xnor U3769 (N_3769,N_3557,N_3370);
nand U3770 (N_3770,N_3434,N_3411);
nor U3771 (N_3771,N_3557,N_3416);
nor U3772 (N_3772,N_3406,N_3434);
xnor U3773 (N_3773,N_3484,N_3461);
xor U3774 (N_3774,N_3323,N_3597);
or U3775 (N_3775,N_3421,N_3354);
nor U3776 (N_3776,N_3584,N_3525);
or U3777 (N_3777,N_3372,N_3520);
nor U3778 (N_3778,N_3381,N_3405);
nand U3779 (N_3779,N_3451,N_3535);
nand U3780 (N_3780,N_3595,N_3592);
and U3781 (N_3781,N_3552,N_3582);
nor U3782 (N_3782,N_3419,N_3538);
xnor U3783 (N_3783,N_3472,N_3316);
and U3784 (N_3784,N_3586,N_3380);
nand U3785 (N_3785,N_3309,N_3395);
nor U3786 (N_3786,N_3371,N_3544);
nor U3787 (N_3787,N_3556,N_3592);
or U3788 (N_3788,N_3363,N_3515);
and U3789 (N_3789,N_3542,N_3379);
xor U3790 (N_3790,N_3462,N_3452);
nor U3791 (N_3791,N_3489,N_3402);
nor U3792 (N_3792,N_3519,N_3598);
or U3793 (N_3793,N_3364,N_3435);
or U3794 (N_3794,N_3371,N_3376);
xnor U3795 (N_3795,N_3456,N_3534);
xnor U3796 (N_3796,N_3456,N_3495);
or U3797 (N_3797,N_3495,N_3376);
xnor U3798 (N_3798,N_3439,N_3583);
or U3799 (N_3799,N_3395,N_3317);
or U3800 (N_3800,N_3412,N_3457);
xnor U3801 (N_3801,N_3306,N_3378);
xnor U3802 (N_3802,N_3343,N_3349);
nand U3803 (N_3803,N_3371,N_3460);
xor U3804 (N_3804,N_3423,N_3551);
xnor U3805 (N_3805,N_3369,N_3337);
or U3806 (N_3806,N_3346,N_3483);
nor U3807 (N_3807,N_3409,N_3359);
nand U3808 (N_3808,N_3414,N_3394);
nor U3809 (N_3809,N_3414,N_3508);
or U3810 (N_3810,N_3360,N_3387);
nor U3811 (N_3811,N_3568,N_3545);
xor U3812 (N_3812,N_3328,N_3586);
nor U3813 (N_3813,N_3353,N_3517);
nand U3814 (N_3814,N_3345,N_3406);
xnor U3815 (N_3815,N_3438,N_3451);
nand U3816 (N_3816,N_3559,N_3511);
and U3817 (N_3817,N_3381,N_3439);
or U3818 (N_3818,N_3479,N_3383);
and U3819 (N_3819,N_3436,N_3447);
or U3820 (N_3820,N_3551,N_3507);
and U3821 (N_3821,N_3323,N_3318);
nor U3822 (N_3822,N_3557,N_3434);
or U3823 (N_3823,N_3451,N_3567);
nor U3824 (N_3824,N_3381,N_3308);
or U3825 (N_3825,N_3404,N_3498);
or U3826 (N_3826,N_3338,N_3425);
nand U3827 (N_3827,N_3364,N_3588);
or U3828 (N_3828,N_3545,N_3323);
nor U3829 (N_3829,N_3557,N_3430);
nand U3830 (N_3830,N_3485,N_3379);
or U3831 (N_3831,N_3549,N_3578);
or U3832 (N_3832,N_3370,N_3412);
or U3833 (N_3833,N_3399,N_3453);
xnor U3834 (N_3834,N_3573,N_3328);
nand U3835 (N_3835,N_3597,N_3319);
nor U3836 (N_3836,N_3448,N_3405);
or U3837 (N_3837,N_3554,N_3557);
or U3838 (N_3838,N_3574,N_3496);
nand U3839 (N_3839,N_3408,N_3566);
and U3840 (N_3840,N_3427,N_3365);
xor U3841 (N_3841,N_3448,N_3592);
nor U3842 (N_3842,N_3408,N_3400);
and U3843 (N_3843,N_3524,N_3323);
nand U3844 (N_3844,N_3534,N_3356);
nor U3845 (N_3845,N_3573,N_3415);
xor U3846 (N_3846,N_3370,N_3533);
xor U3847 (N_3847,N_3328,N_3352);
or U3848 (N_3848,N_3414,N_3554);
xnor U3849 (N_3849,N_3443,N_3312);
or U3850 (N_3850,N_3479,N_3373);
or U3851 (N_3851,N_3575,N_3490);
nor U3852 (N_3852,N_3526,N_3556);
nand U3853 (N_3853,N_3549,N_3349);
nand U3854 (N_3854,N_3318,N_3322);
or U3855 (N_3855,N_3486,N_3501);
xor U3856 (N_3856,N_3321,N_3513);
nor U3857 (N_3857,N_3376,N_3406);
xnor U3858 (N_3858,N_3356,N_3391);
xnor U3859 (N_3859,N_3423,N_3427);
xnor U3860 (N_3860,N_3498,N_3362);
or U3861 (N_3861,N_3475,N_3546);
and U3862 (N_3862,N_3450,N_3386);
and U3863 (N_3863,N_3308,N_3399);
and U3864 (N_3864,N_3574,N_3422);
nor U3865 (N_3865,N_3474,N_3588);
xnor U3866 (N_3866,N_3433,N_3400);
nor U3867 (N_3867,N_3429,N_3501);
or U3868 (N_3868,N_3500,N_3394);
or U3869 (N_3869,N_3402,N_3510);
xor U3870 (N_3870,N_3327,N_3477);
nor U3871 (N_3871,N_3488,N_3318);
nand U3872 (N_3872,N_3346,N_3343);
or U3873 (N_3873,N_3353,N_3323);
xnor U3874 (N_3874,N_3468,N_3572);
xor U3875 (N_3875,N_3511,N_3459);
nand U3876 (N_3876,N_3324,N_3407);
and U3877 (N_3877,N_3532,N_3313);
or U3878 (N_3878,N_3401,N_3400);
or U3879 (N_3879,N_3518,N_3599);
nor U3880 (N_3880,N_3476,N_3344);
and U3881 (N_3881,N_3458,N_3370);
and U3882 (N_3882,N_3577,N_3303);
nor U3883 (N_3883,N_3430,N_3409);
and U3884 (N_3884,N_3586,N_3426);
nand U3885 (N_3885,N_3451,N_3320);
or U3886 (N_3886,N_3467,N_3469);
and U3887 (N_3887,N_3375,N_3465);
or U3888 (N_3888,N_3474,N_3406);
or U3889 (N_3889,N_3559,N_3398);
xor U3890 (N_3890,N_3428,N_3306);
xnor U3891 (N_3891,N_3397,N_3592);
and U3892 (N_3892,N_3351,N_3353);
or U3893 (N_3893,N_3539,N_3519);
nand U3894 (N_3894,N_3376,N_3490);
and U3895 (N_3895,N_3467,N_3395);
nand U3896 (N_3896,N_3502,N_3409);
or U3897 (N_3897,N_3421,N_3463);
nand U3898 (N_3898,N_3409,N_3448);
nor U3899 (N_3899,N_3535,N_3399);
xnor U3900 (N_3900,N_3707,N_3608);
xnor U3901 (N_3901,N_3771,N_3831);
or U3902 (N_3902,N_3739,N_3672);
and U3903 (N_3903,N_3688,N_3708);
or U3904 (N_3904,N_3788,N_3700);
and U3905 (N_3905,N_3809,N_3897);
and U3906 (N_3906,N_3892,N_3818);
xnor U3907 (N_3907,N_3732,N_3746);
nand U3908 (N_3908,N_3713,N_3886);
nand U3909 (N_3909,N_3874,N_3813);
nor U3910 (N_3910,N_3738,N_3881);
nor U3911 (N_3911,N_3662,N_3778);
nor U3912 (N_3912,N_3797,N_3763);
and U3913 (N_3913,N_3824,N_3604);
xor U3914 (N_3914,N_3721,N_3876);
nor U3915 (N_3915,N_3849,N_3751);
nand U3916 (N_3916,N_3845,N_3804);
and U3917 (N_3917,N_3833,N_3650);
xor U3918 (N_3918,N_3684,N_3769);
nand U3919 (N_3919,N_3836,N_3622);
or U3920 (N_3920,N_3756,N_3642);
nand U3921 (N_3921,N_3726,N_3750);
or U3922 (N_3922,N_3776,N_3605);
xnor U3923 (N_3923,N_3888,N_3737);
xor U3924 (N_3924,N_3693,N_3657);
and U3925 (N_3925,N_3618,N_3795);
or U3926 (N_3926,N_3733,N_3743);
nand U3927 (N_3927,N_3861,N_3865);
xnor U3928 (N_3928,N_3641,N_3759);
and U3929 (N_3929,N_3663,N_3819);
or U3930 (N_3930,N_3667,N_3669);
or U3931 (N_3931,N_3855,N_3723);
nand U3932 (N_3932,N_3682,N_3649);
xnor U3933 (N_3933,N_3614,N_3864);
nor U3934 (N_3934,N_3815,N_3821);
xor U3935 (N_3935,N_3734,N_3617);
nand U3936 (N_3936,N_3810,N_3757);
nand U3937 (N_3937,N_3696,N_3814);
and U3938 (N_3938,N_3600,N_3890);
xor U3939 (N_3939,N_3882,N_3867);
nor U3940 (N_3940,N_3764,N_3725);
and U3941 (N_3941,N_3740,N_3727);
or U3942 (N_3942,N_3654,N_3841);
and U3943 (N_3943,N_3875,N_3638);
or U3944 (N_3944,N_3811,N_3630);
nand U3945 (N_3945,N_3646,N_3767);
xnor U3946 (N_3946,N_3679,N_3619);
xnor U3947 (N_3947,N_3636,N_3893);
nand U3948 (N_3948,N_3703,N_3632);
nor U3949 (N_3949,N_3768,N_3828);
and U3950 (N_3950,N_3678,N_3798);
xnor U3951 (N_3951,N_3747,N_3782);
or U3952 (N_3952,N_3668,N_3774);
and U3953 (N_3953,N_3644,N_3629);
nor U3954 (N_3954,N_3710,N_3611);
or U3955 (N_3955,N_3698,N_3854);
and U3956 (N_3956,N_3832,N_3887);
xnor U3957 (N_3957,N_3772,N_3862);
xor U3958 (N_3958,N_3722,N_3752);
nand U3959 (N_3959,N_3883,N_3791);
nor U3960 (N_3960,N_3775,N_3607);
nor U3961 (N_3961,N_3633,N_3820);
nor U3962 (N_3962,N_3834,N_3784);
nand U3963 (N_3963,N_3623,N_3896);
xnor U3964 (N_3964,N_3805,N_3616);
or U3965 (N_3965,N_3749,N_3706);
and U3966 (N_3966,N_3685,N_3736);
xnor U3967 (N_3967,N_3694,N_3793);
nor U3968 (N_3968,N_3885,N_3871);
nor U3969 (N_3969,N_3785,N_3635);
nand U3970 (N_3970,N_3786,N_3661);
nor U3971 (N_3971,N_3844,N_3826);
nand U3972 (N_3972,N_3655,N_3856);
or U3973 (N_3973,N_3760,N_3891);
and U3974 (N_3974,N_3762,N_3877);
nor U3975 (N_3975,N_3626,N_3730);
nor U3976 (N_3976,N_3806,N_3651);
or U3977 (N_3977,N_3719,N_3643);
and U3978 (N_3978,N_3660,N_3825);
and U3979 (N_3979,N_3753,N_3603);
nand U3980 (N_3980,N_3794,N_3899);
and U3981 (N_3981,N_3701,N_3724);
xor U3982 (N_3982,N_3823,N_3777);
xnor U3983 (N_3983,N_3691,N_3681);
or U3984 (N_3984,N_3859,N_3838);
and U3985 (N_3985,N_3683,N_3714);
nor U3986 (N_3986,N_3677,N_3610);
nor U3987 (N_3987,N_3673,N_3686);
or U3988 (N_3988,N_3658,N_3695);
nor U3989 (N_3989,N_3674,N_3731);
and U3990 (N_3990,N_3748,N_3816);
nand U3991 (N_3991,N_3766,N_3742);
xnor U3992 (N_3992,N_3601,N_3689);
nor U3993 (N_3993,N_3645,N_3853);
or U3994 (N_3994,N_3755,N_3758);
xor U3995 (N_3995,N_3884,N_3664);
and U3996 (N_3996,N_3640,N_3781);
nor U3997 (N_3997,N_3652,N_3624);
or U3998 (N_3998,N_3666,N_3676);
and U3999 (N_3999,N_3835,N_3829);
and U4000 (N_4000,N_3858,N_3843);
nand U4001 (N_4001,N_3720,N_3789);
nand U4002 (N_4002,N_3765,N_3709);
xor U4003 (N_4003,N_3680,N_3830);
nand U4004 (N_4004,N_3656,N_3799);
and U4005 (N_4005,N_3827,N_3729);
xor U4006 (N_4006,N_3648,N_3741);
or U4007 (N_4007,N_3615,N_3704);
or U4008 (N_4008,N_3889,N_3625);
xor U4009 (N_4009,N_3898,N_3606);
nand U4010 (N_4010,N_3697,N_3852);
nand U4011 (N_4011,N_3671,N_3773);
or U4012 (N_4012,N_3705,N_3894);
and U4013 (N_4013,N_3792,N_3602);
or U4014 (N_4014,N_3808,N_3728);
xnor U4015 (N_4015,N_3873,N_3863);
nand U4016 (N_4016,N_3860,N_3647);
nor U4017 (N_4017,N_3639,N_3780);
nand U4018 (N_4018,N_3612,N_3879);
or U4019 (N_4019,N_3754,N_3807);
nor U4020 (N_4020,N_3620,N_3692);
and U4021 (N_4021,N_3880,N_3761);
or U4022 (N_4022,N_3735,N_3839);
nand U4023 (N_4023,N_3631,N_3857);
xor U4024 (N_4024,N_3803,N_3817);
nand U4025 (N_4025,N_3822,N_3665);
nor U4026 (N_4026,N_3840,N_3670);
and U4027 (N_4027,N_3868,N_3770);
or U4028 (N_4028,N_3846,N_3718);
nand U4029 (N_4029,N_3716,N_3800);
or U4030 (N_4030,N_3715,N_3790);
nand U4031 (N_4031,N_3628,N_3711);
and U4032 (N_4032,N_3783,N_3801);
xor U4033 (N_4033,N_3717,N_3699);
or U4034 (N_4034,N_3802,N_3779);
nor U4035 (N_4035,N_3675,N_3872);
or U4036 (N_4036,N_3812,N_3627);
and U4037 (N_4037,N_3687,N_3837);
and U4038 (N_4038,N_3745,N_3744);
and U4039 (N_4039,N_3869,N_3653);
and U4040 (N_4040,N_3842,N_3609);
or U4041 (N_4041,N_3870,N_3796);
and U4042 (N_4042,N_3850,N_3878);
nand U4043 (N_4043,N_3848,N_3895);
nand U4044 (N_4044,N_3634,N_3702);
nand U4045 (N_4045,N_3613,N_3659);
and U4046 (N_4046,N_3690,N_3712);
xor U4047 (N_4047,N_3851,N_3866);
nor U4048 (N_4048,N_3621,N_3787);
xor U4049 (N_4049,N_3637,N_3847);
nand U4050 (N_4050,N_3650,N_3821);
xor U4051 (N_4051,N_3705,N_3635);
and U4052 (N_4052,N_3771,N_3803);
or U4053 (N_4053,N_3756,N_3760);
xnor U4054 (N_4054,N_3715,N_3672);
and U4055 (N_4055,N_3877,N_3866);
nor U4056 (N_4056,N_3712,N_3615);
nand U4057 (N_4057,N_3618,N_3669);
and U4058 (N_4058,N_3601,N_3754);
nor U4059 (N_4059,N_3882,N_3699);
xnor U4060 (N_4060,N_3863,N_3619);
xor U4061 (N_4061,N_3789,N_3890);
xor U4062 (N_4062,N_3868,N_3755);
nand U4063 (N_4063,N_3859,N_3833);
xor U4064 (N_4064,N_3719,N_3689);
nor U4065 (N_4065,N_3675,N_3711);
xor U4066 (N_4066,N_3805,N_3798);
or U4067 (N_4067,N_3729,N_3848);
or U4068 (N_4068,N_3689,N_3803);
nor U4069 (N_4069,N_3800,N_3669);
and U4070 (N_4070,N_3893,N_3814);
or U4071 (N_4071,N_3872,N_3890);
or U4072 (N_4072,N_3666,N_3689);
nand U4073 (N_4073,N_3665,N_3897);
nor U4074 (N_4074,N_3898,N_3708);
nor U4075 (N_4075,N_3771,N_3736);
nor U4076 (N_4076,N_3617,N_3632);
xnor U4077 (N_4077,N_3710,N_3758);
xnor U4078 (N_4078,N_3824,N_3686);
nand U4079 (N_4079,N_3679,N_3782);
xor U4080 (N_4080,N_3681,N_3866);
nand U4081 (N_4081,N_3821,N_3827);
xor U4082 (N_4082,N_3736,N_3880);
nand U4083 (N_4083,N_3898,N_3640);
nor U4084 (N_4084,N_3627,N_3745);
nor U4085 (N_4085,N_3605,N_3838);
nand U4086 (N_4086,N_3810,N_3823);
or U4087 (N_4087,N_3753,N_3670);
and U4088 (N_4088,N_3872,N_3895);
or U4089 (N_4089,N_3622,N_3810);
nor U4090 (N_4090,N_3796,N_3628);
or U4091 (N_4091,N_3857,N_3826);
xnor U4092 (N_4092,N_3669,N_3842);
and U4093 (N_4093,N_3724,N_3603);
or U4094 (N_4094,N_3879,N_3823);
xnor U4095 (N_4095,N_3669,N_3831);
or U4096 (N_4096,N_3704,N_3698);
nor U4097 (N_4097,N_3660,N_3704);
or U4098 (N_4098,N_3805,N_3815);
nor U4099 (N_4099,N_3876,N_3747);
and U4100 (N_4100,N_3876,N_3754);
nand U4101 (N_4101,N_3836,N_3863);
nand U4102 (N_4102,N_3801,N_3624);
or U4103 (N_4103,N_3794,N_3723);
nand U4104 (N_4104,N_3878,N_3644);
xor U4105 (N_4105,N_3730,N_3769);
nand U4106 (N_4106,N_3766,N_3836);
nor U4107 (N_4107,N_3769,N_3746);
and U4108 (N_4108,N_3895,N_3608);
or U4109 (N_4109,N_3802,N_3669);
xor U4110 (N_4110,N_3602,N_3699);
nor U4111 (N_4111,N_3660,N_3857);
xor U4112 (N_4112,N_3602,N_3633);
xnor U4113 (N_4113,N_3858,N_3777);
and U4114 (N_4114,N_3839,N_3899);
nand U4115 (N_4115,N_3792,N_3786);
nand U4116 (N_4116,N_3867,N_3647);
nor U4117 (N_4117,N_3753,N_3673);
xnor U4118 (N_4118,N_3888,N_3832);
or U4119 (N_4119,N_3811,N_3774);
nand U4120 (N_4120,N_3604,N_3601);
nor U4121 (N_4121,N_3779,N_3798);
or U4122 (N_4122,N_3883,N_3641);
xnor U4123 (N_4123,N_3613,N_3892);
xor U4124 (N_4124,N_3822,N_3886);
xnor U4125 (N_4125,N_3706,N_3713);
xnor U4126 (N_4126,N_3896,N_3698);
xor U4127 (N_4127,N_3610,N_3878);
or U4128 (N_4128,N_3719,N_3797);
nand U4129 (N_4129,N_3727,N_3834);
nor U4130 (N_4130,N_3647,N_3899);
and U4131 (N_4131,N_3739,N_3674);
nand U4132 (N_4132,N_3833,N_3792);
nor U4133 (N_4133,N_3786,N_3714);
or U4134 (N_4134,N_3701,N_3640);
or U4135 (N_4135,N_3783,N_3648);
nand U4136 (N_4136,N_3628,N_3622);
nand U4137 (N_4137,N_3789,N_3730);
nor U4138 (N_4138,N_3681,N_3740);
nand U4139 (N_4139,N_3675,N_3692);
xor U4140 (N_4140,N_3610,N_3763);
nor U4141 (N_4141,N_3861,N_3777);
or U4142 (N_4142,N_3612,N_3666);
nand U4143 (N_4143,N_3772,N_3882);
or U4144 (N_4144,N_3630,N_3680);
nor U4145 (N_4145,N_3856,N_3659);
nand U4146 (N_4146,N_3731,N_3737);
xnor U4147 (N_4147,N_3771,N_3679);
and U4148 (N_4148,N_3689,N_3672);
or U4149 (N_4149,N_3778,N_3840);
nor U4150 (N_4150,N_3822,N_3720);
or U4151 (N_4151,N_3819,N_3645);
nand U4152 (N_4152,N_3743,N_3614);
and U4153 (N_4153,N_3836,N_3776);
and U4154 (N_4154,N_3828,N_3667);
nand U4155 (N_4155,N_3839,N_3834);
nor U4156 (N_4156,N_3886,N_3878);
nand U4157 (N_4157,N_3701,N_3860);
or U4158 (N_4158,N_3827,N_3825);
xnor U4159 (N_4159,N_3747,N_3758);
xor U4160 (N_4160,N_3721,N_3680);
xor U4161 (N_4161,N_3639,N_3717);
and U4162 (N_4162,N_3676,N_3687);
or U4163 (N_4163,N_3736,N_3625);
and U4164 (N_4164,N_3733,N_3739);
or U4165 (N_4165,N_3874,N_3606);
and U4166 (N_4166,N_3684,N_3739);
and U4167 (N_4167,N_3682,N_3764);
and U4168 (N_4168,N_3751,N_3750);
or U4169 (N_4169,N_3839,N_3796);
nor U4170 (N_4170,N_3841,N_3805);
and U4171 (N_4171,N_3633,N_3737);
nor U4172 (N_4172,N_3716,N_3684);
nand U4173 (N_4173,N_3871,N_3793);
nand U4174 (N_4174,N_3621,N_3831);
nor U4175 (N_4175,N_3867,N_3828);
xor U4176 (N_4176,N_3652,N_3764);
and U4177 (N_4177,N_3723,N_3825);
and U4178 (N_4178,N_3704,N_3622);
and U4179 (N_4179,N_3848,N_3623);
or U4180 (N_4180,N_3860,N_3633);
and U4181 (N_4181,N_3813,N_3852);
nand U4182 (N_4182,N_3888,N_3692);
or U4183 (N_4183,N_3741,N_3694);
nand U4184 (N_4184,N_3674,N_3795);
nor U4185 (N_4185,N_3662,N_3736);
and U4186 (N_4186,N_3733,N_3686);
xor U4187 (N_4187,N_3893,N_3682);
and U4188 (N_4188,N_3663,N_3754);
or U4189 (N_4189,N_3839,N_3812);
or U4190 (N_4190,N_3605,N_3733);
or U4191 (N_4191,N_3754,N_3847);
nor U4192 (N_4192,N_3633,N_3793);
nand U4193 (N_4193,N_3749,N_3621);
or U4194 (N_4194,N_3874,N_3846);
xor U4195 (N_4195,N_3828,N_3674);
or U4196 (N_4196,N_3710,N_3767);
xnor U4197 (N_4197,N_3748,N_3698);
nand U4198 (N_4198,N_3613,N_3788);
or U4199 (N_4199,N_3767,N_3774);
nor U4200 (N_4200,N_3997,N_4061);
nor U4201 (N_4201,N_4160,N_4041);
nor U4202 (N_4202,N_4166,N_3947);
and U4203 (N_4203,N_3966,N_4118);
and U4204 (N_4204,N_4198,N_4152);
nand U4205 (N_4205,N_4101,N_3968);
nor U4206 (N_4206,N_4057,N_4018);
nand U4207 (N_4207,N_4171,N_4058);
xnor U4208 (N_4208,N_4167,N_4093);
or U4209 (N_4209,N_4053,N_4019);
nor U4210 (N_4210,N_4078,N_4007);
nand U4211 (N_4211,N_4134,N_4001);
xor U4212 (N_4212,N_4131,N_4047);
and U4213 (N_4213,N_3978,N_4073);
nand U4214 (N_4214,N_4147,N_4179);
and U4215 (N_4215,N_4157,N_3915);
and U4216 (N_4216,N_4128,N_4129);
or U4217 (N_4217,N_4066,N_4153);
nor U4218 (N_4218,N_4027,N_3986);
nor U4219 (N_4219,N_4062,N_4105);
nand U4220 (N_4220,N_4127,N_3937);
nand U4221 (N_4221,N_3957,N_4145);
xnor U4222 (N_4222,N_4032,N_4056);
and U4223 (N_4223,N_3903,N_3995);
xor U4224 (N_4224,N_4136,N_4138);
nand U4225 (N_4225,N_4035,N_4170);
nor U4226 (N_4226,N_4126,N_3972);
or U4227 (N_4227,N_3921,N_4119);
and U4228 (N_4228,N_3965,N_4072);
nand U4229 (N_4229,N_3949,N_3991);
xor U4230 (N_4230,N_4089,N_4184);
and U4231 (N_4231,N_4199,N_3927);
xor U4232 (N_4232,N_4196,N_4055);
nor U4233 (N_4233,N_4059,N_4017);
and U4234 (N_4234,N_4109,N_4162);
xor U4235 (N_4235,N_4005,N_3993);
nor U4236 (N_4236,N_3930,N_4130);
or U4237 (N_4237,N_4116,N_3979);
xnor U4238 (N_4238,N_4025,N_3918);
xnor U4239 (N_4239,N_3950,N_3974);
nand U4240 (N_4240,N_4183,N_4068);
and U4241 (N_4241,N_4188,N_4192);
nor U4242 (N_4242,N_3938,N_4120);
nor U4243 (N_4243,N_3945,N_4177);
nor U4244 (N_4244,N_4037,N_3964);
xor U4245 (N_4245,N_4150,N_4180);
nor U4246 (N_4246,N_4121,N_4030);
and U4247 (N_4247,N_3967,N_3943);
xor U4248 (N_4248,N_3923,N_4046);
and U4249 (N_4249,N_3929,N_4139);
and U4250 (N_4250,N_4115,N_3900);
nor U4251 (N_4251,N_4094,N_4125);
xor U4252 (N_4252,N_3911,N_4028);
nand U4253 (N_4253,N_4043,N_3955);
or U4254 (N_4254,N_4023,N_4155);
nor U4255 (N_4255,N_4067,N_4107);
and U4256 (N_4256,N_4029,N_4176);
xor U4257 (N_4257,N_4190,N_3926);
nor U4258 (N_4258,N_4106,N_3984);
or U4259 (N_4259,N_3917,N_4151);
nor U4260 (N_4260,N_4174,N_4172);
or U4261 (N_4261,N_3922,N_4102);
xnor U4262 (N_4262,N_4051,N_4175);
nor U4263 (N_4263,N_3941,N_4050);
xnor U4264 (N_4264,N_4108,N_4012);
xnor U4265 (N_4265,N_4158,N_4079);
nand U4266 (N_4266,N_3956,N_4069);
and U4267 (N_4267,N_3901,N_4006);
nand U4268 (N_4268,N_4004,N_4140);
and U4269 (N_4269,N_4112,N_3994);
xor U4270 (N_4270,N_3931,N_3952);
and U4271 (N_4271,N_4026,N_4084);
or U4272 (N_4272,N_4161,N_3944);
and U4273 (N_4273,N_4081,N_4137);
nand U4274 (N_4274,N_4049,N_4142);
nand U4275 (N_4275,N_3948,N_4022);
and U4276 (N_4276,N_4194,N_4163);
nor U4277 (N_4277,N_3958,N_3914);
nor U4278 (N_4278,N_4100,N_4169);
nor U4279 (N_4279,N_3913,N_3999);
xnor U4280 (N_4280,N_3988,N_3940);
or U4281 (N_4281,N_3925,N_4091);
nor U4282 (N_4282,N_4103,N_3932);
and U4283 (N_4283,N_4031,N_4090);
or U4284 (N_4284,N_3971,N_4016);
nor U4285 (N_4285,N_4168,N_4191);
or U4286 (N_4286,N_4076,N_4164);
and U4287 (N_4287,N_3992,N_3910);
or U4288 (N_4288,N_3902,N_4086);
and U4289 (N_4289,N_4034,N_3977);
nand U4290 (N_4290,N_4141,N_4020);
nand U4291 (N_4291,N_4114,N_4111);
nor U4292 (N_4292,N_4186,N_3906);
and U4293 (N_4293,N_4077,N_3912);
nor U4294 (N_4294,N_3939,N_4187);
or U4295 (N_4295,N_4098,N_4124);
or U4296 (N_4296,N_4080,N_4133);
nor U4297 (N_4297,N_3976,N_4045);
xor U4298 (N_4298,N_3953,N_4193);
or U4299 (N_4299,N_3924,N_4064);
and U4300 (N_4300,N_4185,N_4146);
xor U4301 (N_4301,N_4099,N_3936);
or U4302 (N_4302,N_4173,N_3970);
or U4303 (N_4303,N_4063,N_4039);
and U4304 (N_4304,N_4144,N_3983);
xnor U4305 (N_4305,N_4033,N_4095);
xnor U4306 (N_4306,N_4065,N_3987);
nand U4307 (N_4307,N_3989,N_3934);
nand U4308 (N_4308,N_3907,N_3982);
or U4309 (N_4309,N_3916,N_3935);
and U4310 (N_4310,N_4014,N_4011);
and U4311 (N_4311,N_4156,N_4048);
nor U4312 (N_4312,N_3946,N_4038);
and U4313 (N_4313,N_4054,N_3985);
nand U4314 (N_4314,N_4052,N_3908);
xor U4315 (N_4315,N_4075,N_4104);
or U4316 (N_4316,N_4113,N_4117);
xor U4317 (N_4317,N_3954,N_4000);
and U4318 (N_4318,N_4021,N_4159);
xor U4319 (N_4319,N_4060,N_3963);
nand U4320 (N_4320,N_3981,N_3905);
and U4321 (N_4321,N_3933,N_3990);
nor U4322 (N_4322,N_3996,N_4040);
or U4323 (N_4323,N_4036,N_4135);
nor U4324 (N_4324,N_3962,N_4132);
and U4325 (N_4325,N_4110,N_4013);
xnor U4326 (N_4326,N_4085,N_3919);
nor U4327 (N_4327,N_3928,N_4002);
or U4328 (N_4328,N_3961,N_3909);
nor U4329 (N_4329,N_4123,N_4088);
xor U4330 (N_4330,N_3998,N_4044);
xnor U4331 (N_4331,N_4165,N_4181);
nand U4332 (N_4332,N_4178,N_4154);
nand U4333 (N_4333,N_3980,N_4042);
nor U4334 (N_4334,N_4070,N_4197);
nand U4335 (N_4335,N_4143,N_4009);
xor U4336 (N_4336,N_4071,N_3920);
nand U4337 (N_4337,N_4148,N_4010);
xor U4338 (N_4338,N_4096,N_4015);
nand U4339 (N_4339,N_4097,N_3960);
nor U4340 (N_4340,N_4149,N_4092);
or U4341 (N_4341,N_4195,N_4074);
xor U4342 (N_4342,N_3951,N_4082);
nor U4343 (N_4343,N_4003,N_4182);
xor U4344 (N_4344,N_4024,N_3973);
and U4345 (N_4345,N_4122,N_4189);
and U4346 (N_4346,N_3904,N_4083);
xnor U4347 (N_4347,N_4008,N_3975);
nand U4348 (N_4348,N_3942,N_4087);
or U4349 (N_4349,N_3969,N_3959);
xor U4350 (N_4350,N_3999,N_4056);
nor U4351 (N_4351,N_3969,N_4034);
nand U4352 (N_4352,N_3913,N_3910);
nand U4353 (N_4353,N_4049,N_4169);
nor U4354 (N_4354,N_3928,N_4173);
nor U4355 (N_4355,N_3927,N_4036);
nand U4356 (N_4356,N_4193,N_3973);
xor U4357 (N_4357,N_3954,N_4008);
nand U4358 (N_4358,N_3988,N_4057);
and U4359 (N_4359,N_4044,N_4172);
nor U4360 (N_4360,N_3949,N_3911);
nand U4361 (N_4361,N_4194,N_3955);
and U4362 (N_4362,N_3944,N_4036);
nor U4363 (N_4363,N_4050,N_3939);
xnor U4364 (N_4364,N_4166,N_4068);
nor U4365 (N_4365,N_4117,N_4072);
nand U4366 (N_4366,N_4149,N_4055);
nand U4367 (N_4367,N_3900,N_4160);
xnor U4368 (N_4368,N_4177,N_4171);
and U4369 (N_4369,N_4086,N_4142);
xnor U4370 (N_4370,N_3923,N_4173);
xor U4371 (N_4371,N_4054,N_4008);
and U4372 (N_4372,N_4105,N_4125);
nor U4373 (N_4373,N_3955,N_4044);
and U4374 (N_4374,N_3942,N_4009);
and U4375 (N_4375,N_4084,N_3929);
nand U4376 (N_4376,N_4168,N_3984);
and U4377 (N_4377,N_4111,N_4015);
xor U4378 (N_4378,N_4181,N_4102);
nand U4379 (N_4379,N_3978,N_3926);
nor U4380 (N_4380,N_3962,N_4117);
and U4381 (N_4381,N_4015,N_4076);
nor U4382 (N_4382,N_4192,N_4195);
and U4383 (N_4383,N_4134,N_3940);
nand U4384 (N_4384,N_4007,N_4037);
and U4385 (N_4385,N_3956,N_4082);
and U4386 (N_4386,N_3925,N_4119);
xor U4387 (N_4387,N_4081,N_3931);
xor U4388 (N_4388,N_4070,N_3923);
nor U4389 (N_4389,N_4099,N_3984);
and U4390 (N_4390,N_3904,N_4132);
nor U4391 (N_4391,N_3905,N_3984);
and U4392 (N_4392,N_3943,N_4097);
nor U4393 (N_4393,N_4007,N_4159);
and U4394 (N_4394,N_4135,N_4044);
nor U4395 (N_4395,N_4105,N_4187);
xnor U4396 (N_4396,N_3910,N_3973);
or U4397 (N_4397,N_4198,N_4068);
nor U4398 (N_4398,N_3919,N_4101);
and U4399 (N_4399,N_3948,N_3959);
nor U4400 (N_4400,N_4128,N_4042);
or U4401 (N_4401,N_3959,N_3972);
or U4402 (N_4402,N_4068,N_4027);
nand U4403 (N_4403,N_4159,N_3914);
or U4404 (N_4404,N_4130,N_3992);
nand U4405 (N_4405,N_4152,N_3974);
and U4406 (N_4406,N_4143,N_3910);
nor U4407 (N_4407,N_4043,N_3965);
nand U4408 (N_4408,N_4191,N_4197);
nor U4409 (N_4409,N_4003,N_3916);
and U4410 (N_4410,N_4055,N_3983);
xor U4411 (N_4411,N_4141,N_4000);
nor U4412 (N_4412,N_4036,N_4088);
xnor U4413 (N_4413,N_4030,N_4120);
and U4414 (N_4414,N_4138,N_3904);
nand U4415 (N_4415,N_4117,N_4173);
and U4416 (N_4416,N_4140,N_4113);
and U4417 (N_4417,N_3980,N_4096);
nor U4418 (N_4418,N_4060,N_4112);
and U4419 (N_4419,N_3932,N_3975);
nor U4420 (N_4420,N_3999,N_3945);
and U4421 (N_4421,N_3993,N_4107);
nand U4422 (N_4422,N_3998,N_4105);
nor U4423 (N_4423,N_4083,N_4113);
xnor U4424 (N_4424,N_3932,N_4171);
nor U4425 (N_4425,N_4172,N_3918);
xor U4426 (N_4426,N_4120,N_4149);
or U4427 (N_4427,N_3923,N_4178);
and U4428 (N_4428,N_3973,N_4098);
xor U4429 (N_4429,N_4167,N_3924);
or U4430 (N_4430,N_4167,N_4195);
nor U4431 (N_4431,N_4046,N_4147);
nor U4432 (N_4432,N_4161,N_4071);
nor U4433 (N_4433,N_4083,N_4055);
or U4434 (N_4434,N_4077,N_3922);
nor U4435 (N_4435,N_4020,N_4068);
nand U4436 (N_4436,N_4007,N_3915);
or U4437 (N_4437,N_4028,N_3936);
and U4438 (N_4438,N_4009,N_4084);
or U4439 (N_4439,N_4084,N_4049);
xnor U4440 (N_4440,N_4017,N_4075);
nand U4441 (N_4441,N_4058,N_3975);
nand U4442 (N_4442,N_4083,N_4111);
nor U4443 (N_4443,N_4045,N_3926);
nor U4444 (N_4444,N_3947,N_4133);
or U4445 (N_4445,N_4169,N_3908);
nor U4446 (N_4446,N_3944,N_3988);
xnor U4447 (N_4447,N_3906,N_3933);
nor U4448 (N_4448,N_3924,N_4145);
nand U4449 (N_4449,N_4097,N_4069);
nand U4450 (N_4450,N_4158,N_3988);
xor U4451 (N_4451,N_4017,N_4116);
and U4452 (N_4452,N_4036,N_4010);
or U4453 (N_4453,N_3985,N_3991);
xor U4454 (N_4454,N_4002,N_4017);
nand U4455 (N_4455,N_4065,N_3947);
or U4456 (N_4456,N_4129,N_4105);
nor U4457 (N_4457,N_3992,N_4105);
nand U4458 (N_4458,N_4013,N_4197);
nor U4459 (N_4459,N_4014,N_3917);
nor U4460 (N_4460,N_4139,N_3951);
nor U4461 (N_4461,N_4179,N_4093);
and U4462 (N_4462,N_3931,N_3979);
nand U4463 (N_4463,N_4114,N_3945);
xnor U4464 (N_4464,N_4067,N_4023);
nand U4465 (N_4465,N_4083,N_4173);
nand U4466 (N_4466,N_3975,N_4002);
xor U4467 (N_4467,N_4076,N_4040);
nor U4468 (N_4468,N_4083,N_3905);
xor U4469 (N_4469,N_3923,N_3933);
nor U4470 (N_4470,N_4182,N_3996);
xnor U4471 (N_4471,N_3987,N_4055);
or U4472 (N_4472,N_3927,N_3989);
and U4473 (N_4473,N_3999,N_3982);
nand U4474 (N_4474,N_3934,N_4004);
nor U4475 (N_4475,N_3944,N_4124);
or U4476 (N_4476,N_3927,N_3994);
or U4477 (N_4477,N_4068,N_3963);
or U4478 (N_4478,N_3944,N_4064);
and U4479 (N_4479,N_4077,N_4100);
nand U4480 (N_4480,N_3902,N_4108);
and U4481 (N_4481,N_3900,N_4089);
xnor U4482 (N_4482,N_4030,N_3915);
nand U4483 (N_4483,N_4014,N_4003);
xor U4484 (N_4484,N_4072,N_3907);
nor U4485 (N_4485,N_4189,N_4044);
xnor U4486 (N_4486,N_4178,N_4189);
nor U4487 (N_4487,N_4067,N_3930);
nand U4488 (N_4488,N_3981,N_4142);
xor U4489 (N_4489,N_4111,N_3991);
or U4490 (N_4490,N_3975,N_3974);
and U4491 (N_4491,N_4150,N_3992);
nor U4492 (N_4492,N_3921,N_3931);
nand U4493 (N_4493,N_4118,N_3913);
and U4494 (N_4494,N_4031,N_4109);
nor U4495 (N_4495,N_4184,N_4168);
nor U4496 (N_4496,N_3928,N_4095);
nand U4497 (N_4497,N_3907,N_3943);
xor U4498 (N_4498,N_4119,N_4092);
nor U4499 (N_4499,N_3901,N_4147);
nor U4500 (N_4500,N_4240,N_4379);
nor U4501 (N_4501,N_4247,N_4348);
and U4502 (N_4502,N_4326,N_4293);
and U4503 (N_4503,N_4301,N_4400);
nor U4504 (N_4504,N_4239,N_4456);
or U4505 (N_4505,N_4487,N_4223);
xor U4506 (N_4506,N_4231,N_4337);
or U4507 (N_4507,N_4334,N_4453);
or U4508 (N_4508,N_4479,N_4288);
nor U4509 (N_4509,N_4366,N_4261);
and U4510 (N_4510,N_4317,N_4286);
xnor U4511 (N_4511,N_4344,N_4258);
nand U4512 (N_4512,N_4346,N_4279);
nand U4513 (N_4513,N_4455,N_4257);
nor U4514 (N_4514,N_4207,N_4322);
xor U4515 (N_4515,N_4458,N_4353);
and U4516 (N_4516,N_4225,N_4454);
or U4517 (N_4517,N_4267,N_4252);
nor U4518 (N_4518,N_4451,N_4265);
and U4519 (N_4519,N_4382,N_4251);
or U4520 (N_4520,N_4367,N_4450);
nand U4521 (N_4521,N_4374,N_4270);
and U4522 (N_4522,N_4206,N_4269);
or U4523 (N_4523,N_4394,N_4427);
or U4524 (N_4524,N_4282,N_4295);
nand U4525 (N_4525,N_4307,N_4368);
nor U4526 (N_4526,N_4484,N_4475);
nor U4527 (N_4527,N_4491,N_4418);
xnor U4528 (N_4528,N_4444,N_4470);
xor U4529 (N_4529,N_4404,N_4228);
nor U4530 (N_4530,N_4417,N_4256);
nand U4531 (N_4531,N_4436,N_4424);
nand U4532 (N_4532,N_4320,N_4280);
xor U4533 (N_4533,N_4481,N_4467);
or U4534 (N_4534,N_4294,N_4312);
nand U4535 (N_4535,N_4290,N_4381);
xnor U4536 (N_4536,N_4416,N_4438);
nor U4537 (N_4537,N_4340,N_4241);
and U4538 (N_4538,N_4216,N_4474);
xnor U4539 (N_4539,N_4237,N_4311);
nand U4540 (N_4540,N_4421,N_4389);
and U4541 (N_4541,N_4242,N_4358);
nor U4542 (N_4542,N_4413,N_4443);
nor U4543 (N_4543,N_4403,N_4375);
nor U4544 (N_4544,N_4328,N_4437);
nor U4545 (N_4545,N_4380,N_4289);
nor U4546 (N_4546,N_4415,N_4472);
nand U4547 (N_4547,N_4271,N_4296);
or U4548 (N_4548,N_4214,N_4325);
xnor U4549 (N_4549,N_4445,N_4492);
or U4550 (N_4550,N_4373,N_4327);
xor U4551 (N_4551,N_4477,N_4468);
xor U4552 (N_4552,N_4278,N_4384);
xor U4553 (N_4553,N_4426,N_4466);
nor U4554 (N_4554,N_4494,N_4496);
nor U4555 (N_4555,N_4230,N_4315);
and U4556 (N_4556,N_4473,N_4341);
nand U4557 (N_4557,N_4245,N_4482);
xor U4558 (N_4558,N_4486,N_4359);
xnor U4559 (N_4559,N_4433,N_4243);
and U4560 (N_4560,N_4365,N_4420);
xnor U4561 (N_4561,N_4268,N_4485);
xnor U4562 (N_4562,N_4330,N_4483);
nor U4563 (N_4563,N_4281,N_4446);
nand U4564 (N_4564,N_4246,N_4407);
nor U4565 (N_4565,N_4305,N_4302);
nor U4566 (N_4566,N_4463,N_4360);
and U4567 (N_4567,N_4499,N_4419);
nand U4568 (N_4568,N_4357,N_4234);
or U4569 (N_4569,N_4277,N_4263);
xnor U4570 (N_4570,N_4332,N_4405);
nand U4571 (N_4571,N_4291,N_4209);
nor U4572 (N_4572,N_4253,N_4319);
xnor U4573 (N_4573,N_4355,N_4428);
xor U4574 (N_4574,N_4387,N_4352);
nor U4575 (N_4575,N_4306,N_4442);
nand U4576 (N_4576,N_4464,N_4298);
nor U4577 (N_4577,N_4390,N_4364);
or U4578 (N_4578,N_4383,N_4210);
nor U4579 (N_4579,N_4412,N_4248);
nand U4580 (N_4580,N_4273,N_4323);
and U4581 (N_4581,N_4410,N_4376);
nand U4582 (N_4582,N_4349,N_4201);
nand U4583 (N_4583,N_4462,N_4314);
nor U4584 (N_4584,N_4249,N_4272);
and U4585 (N_4585,N_4318,N_4222);
nand U4586 (N_4586,N_4498,N_4284);
nand U4587 (N_4587,N_4440,N_4339);
xor U4588 (N_4588,N_4220,N_4211);
and U4589 (N_4589,N_4465,N_4292);
and U4590 (N_4590,N_4287,N_4370);
nand U4591 (N_4591,N_4488,N_4324);
xor U4592 (N_4592,N_4309,N_4274);
or U4593 (N_4593,N_4378,N_4493);
nand U4594 (N_4594,N_4342,N_4304);
and U4595 (N_4595,N_4409,N_4371);
nand U4596 (N_4596,N_4347,N_4449);
nor U4597 (N_4597,N_4208,N_4388);
nor U4598 (N_4598,N_4232,N_4432);
nand U4599 (N_4599,N_4224,N_4264);
and U4600 (N_4600,N_4459,N_4329);
and U4601 (N_4601,N_4435,N_4414);
nor U4602 (N_4602,N_4215,N_4395);
xor U4603 (N_4603,N_4200,N_4350);
nor U4604 (N_4604,N_4354,N_4259);
xor U4605 (N_4605,N_4285,N_4316);
nand U4606 (N_4606,N_4338,N_4351);
and U4607 (N_4607,N_4276,N_4377);
xor U4608 (N_4608,N_4333,N_4227);
or U4609 (N_4609,N_4397,N_4300);
nand U4610 (N_4610,N_4461,N_4429);
nor U4611 (N_4611,N_4489,N_4205);
nand U4612 (N_4612,N_4204,N_4460);
and U4613 (N_4613,N_4452,N_4254);
or U4614 (N_4614,N_4219,N_4310);
xnor U4615 (N_4615,N_4369,N_4434);
or U4616 (N_4616,N_4238,N_4283);
xnor U4617 (N_4617,N_4266,N_4471);
xor U4618 (N_4618,N_4490,N_4423);
or U4619 (N_4619,N_4217,N_4362);
or U4620 (N_4620,N_4299,N_4430);
nor U4621 (N_4621,N_4203,N_4448);
nand U4622 (N_4622,N_4226,N_4235);
or U4623 (N_4623,N_4233,N_4336);
or U4624 (N_4624,N_4345,N_4386);
nor U4625 (N_4625,N_4218,N_4303);
or U4626 (N_4626,N_4308,N_4356);
nor U4627 (N_4627,N_4497,N_4393);
and U4628 (N_4628,N_4313,N_4361);
and U4629 (N_4629,N_4406,N_4250);
nand U4630 (N_4630,N_4335,N_4255);
nor U4631 (N_4631,N_4343,N_4425);
nand U4632 (N_4632,N_4441,N_4495);
xnor U4633 (N_4633,N_4478,N_4275);
or U4634 (N_4634,N_4244,N_4391);
and U4635 (N_4635,N_4221,N_4411);
or U4636 (N_4636,N_4262,N_4476);
nor U4637 (N_4637,N_4297,N_4447);
xor U4638 (N_4638,N_4363,N_4431);
xnor U4639 (N_4639,N_4422,N_4385);
xor U4640 (N_4640,N_4331,N_4212);
nand U4641 (N_4641,N_4469,N_4408);
nor U4642 (N_4642,N_4213,N_4321);
and U4643 (N_4643,N_4202,N_4398);
nor U4644 (N_4644,N_4260,N_4401);
nor U4645 (N_4645,N_4236,N_4480);
and U4646 (N_4646,N_4399,N_4372);
nand U4647 (N_4647,N_4402,N_4396);
nand U4648 (N_4648,N_4439,N_4229);
or U4649 (N_4649,N_4392,N_4457);
and U4650 (N_4650,N_4362,N_4373);
or U4651 (N_4651,N_4476,N_4263);
nand U4652 (N_4652,N_4230,N_4474);
nand U4653 (N_4653,N_4422,N_4387);
and U4654 (N_4654,N_4245,N_4315);
xnor U4655 (N_4655,N_4480,N_4394);
nor U4656 (N_4656,N_4440,N_4378);
nor U4657 (N_4657,N_4378,N_4283);
or U4658 (N_4658,N_4357,N_4335);
and U4659 (N_4659,N_4216,N_4301);
nor U4660 (N_4660,N_4344,N_4342);
or U4661 (N_4661,N_4276,N_4417);
nor U4662 (N_4662,N_4204,N_4484);
nor U4663 (N_4663,N_4347,N_4241);
xnor U4664 (N_4664,N_4343,N_4476);
nand U4665 (N_4665,N_4463,N_4455);
and U4666 (N_4666,N_4313,N_4257);
and U4667 (N_4667,N_4440,N_4226);
nand U4668 (N_4668,N_4361,N_4338);
nand U4669 (N_4669,N_4479,N_4386);
or U4670 (N_4670,N_4465,N_4442);
or U4671 (N_4671,N_4369,N_4295);
and U4672 (N_4672,N_4394,N_4317);
and U4673 (N_4673,N_4449,N_4283);
nand U4674 (N_4674,N_4282,N_4442);
xor U4675 (N_4675,N_4461,N_4423);
nand U4676 (N_4676,N_4368,N_4431);
and U4677 (N_4677,N_4261,N_4226);
nand U4678 (N_4678,N_4375,N_4361);
xnor U4679 (N_4679,N_4230,N_4310);
or U4680 (N_4680,N_4359,N_4388);
nor U4681 (N_4681,N_4480,N_4337);
and U4682 (N_4682,N_4452,N_4334);
nor U4683 (N_4683,N_4321,N_4259);
xor U4684 (N_4684,N_4478,N_4299);
or U4685 (N_4685,N_4360,N_4208);
nand U4686 (N_4686,N_4334,N_4477);
nand U4687 (N_4687,N_4402,N_4255);
nor U4688 (N_4688,N_4325,N_4334);
xnor U4689 (N_4689,N_4289,N_4438);
nor U4690 (N_4690,N_4408,N_4283);
nor U4691 (N_4691,N_4297,N_4274);
or U4692 (N_4692,N_4363,N_4388);
xnor U4693 (N_4693,N_4408,N_4341);
nor U4694 (N_4694,N_4278,N_4489);
or U4695 (N_4695,N_4427,N_4355);
nand U4696 (N_4696,N_4406,N_4478);
xnor U4697 (N_4697,N_4307,N_4324);
xnor U4698 (N_4698,N_4221,N_4218);
xnor U4699 (N_4699,N_4338,N_4459);
nand U4700 (N_4700,N_4338,N_4271);
nand U4701 (N_4701,N_4384,N_4475);
xor U4702 (N_4702,N_4284,N_4459);
and U4703 (N_4703,N_4372,N_4379);
nand U4704 (N_4704,N_4404,N_4448);
or U4705 (N_4705,N_4252,N_4415);
nand U4706 (N_4706,N_4215,N_4208);
or U4707 (N_4707,N_4476,N_4331);
xnor U4708 (N_4708,N_4283,N_4349);
or U4709 (N_4709,N_4288,N_4359);
and U4710 (N_4710,N_4462,N_4491);
nand U4711 (N_4711,N_4407,N_4385);
or U4712 (N_4712,N_4401,N_4321);
nor U4713 (N_4713,N_4441,N_4338);
xor U4714 (N_4714,N_4284,N_4259);
nor U4715 (N_4715,N_4297,N_4279);
nor U4716 (N_4716,N_4253,N_4369);
and U4717 (N_4717,N_4361,N_4291);
and U4718 (N_4718,N_4440,N_4285);
or U4719 (N_4719,N_4479,N_4388);
or U4720 (N_4720,N_4347,N_4216);
or U4721 (N_4721,N_4408,N_4261);
and U4722 (N_4722,N_4313,N_4290);
nand U4723 (N_4723,N_4303,N_4397);
and U4724 (N_4724,N_4359,N_4489);
and U4725 (N_4725,N_4458,N_4339);
nand U4726 (N_4726,N_4491,N_4426);
or U4727 (N_4727,N_4477,N_4385);
nand U4728 (N_4728,N_4238,N_4269);
and U4729 (N_4729,N_4434,N_4307);
or U4730 (N_4730,N_4308,N_4388);
nand U4731 (N_4731,N_4205,N_4467);
xnor U4732 (N_4732,N_4304,N_4437);
nand U4733 (N_4733,N_4225,N_4233);
nor U4734 (N_4734,N_4439,N_4317);
and U4735 (N_4735,N_4445,N_4203);
xor U4736 (N_4736,N_4242,N_4398);
nor U4737 (N_4737,N_4291,N_4277);
xnor U4738 (N_4738,N_4224,N_4415);
xor U4739 (N_4739,N_4230,N_4263);
nand U4740 (N_4740,N_4206,N_4429);
nand U4741 (N_4741,N_4358,N_4465);
nand U4742 (N_4742,N_4225,N_4238);
and U4743 (N_4743,N_4240,N_4253);
and U4744 (N_4744,N_4377,N_4265);
xor U4745 (N_4745,N_4345,N_4302);
and U4746 (N_4746,N_4461,N_4422);
or U4747 (N_4747,N_4242,N_4344);
nand U4748 (N_4748,N_4465,N_4284);
nand U4749 (N_4749,N_4378,N_4340);
and U4750 (N_4750,N_4329,N_4219);
nor U4751 (N_4751,N_4221,N_4432);
or U4752 (N_4752,N_4349,N_4379);
xor U4753 (N_4753,N_4216,N_4445);
and U4754 (N_4754,N_4283,N_4203);
nand U4755 (N_4755,N_4269,N_4421);
and U4756 (N_4756,N_4258,N_4359);
or U4757 (N_4757,N_4332,N_4240);
xor U4758 (N_4758,N_4225,N_4269);
or U4759 (N_4759,N_4355,N_4365);
nand U4760 (N_4760,N_4472,N_4241);
nor U4761 (N_4761,N_4371,N_4389);
or U4762 (N_4762,N_4319,N_4347);
nand U4763 (N_4763,N_4224,N_4232);
and U4764 (N_4764,N_4498,N_4374);
or U4765 (N_4765,N_4333,N_4454);
or U4766 (N_4766,N_4312,N_4398);
nand U4767 (N_4767,N_4270,N_4376);
nor U4768 (N_4768,N_4417,N_4481);
xnor U4769 (N_4769,N_4345,N_4380);
nand U4770 (N_4770,N_4482,N_4240);
xor U4771 (N_4771,N_4489,N_4441);
and U4772 (N_4772,N_4283,N_4499);
nand U4773 (N_4773,N_4238,N_4370);
or U4774 (N_4774,N_4301,N_4353);
nand U4775 (N_4775,N_4484,N_4492);
or U4776 (N_4776,N_4302,N_4425);
and U4777 (N_4777,N_4476,N_4291);
nand U4778 (N_4778,N_4260,N_4235);
xnor U4779 (N_4779,N_4379,N_4275);
nor U4780 (N_4780,N_4375,N_4391);
nor U4781 (N_4781,N_4304,N_4371);
nand U4782 (N_4782,N_4440,N_4262);
or U4783 (N_4783,N_4309,N_4273);
nand U4784 (N_4784,N_4409,N_4475);
nor U4785 (N_4785,N_4223,N_4379);
or U4786 (N_4786,N_4454,N_4487);
and U4787 (N_4787,N_4219,N_4479);
nand U4788 (N_4788,N_4328,N_4393);
xor U4789 (N_4789,N_4452,N_4448);
nor U4790 (N_4790,N_4294,N_4237);
and U4791 (N_4791,N_4305,N_4238);
or U4792 (N_4792,N_4279,N_4416);
or U4793 (N_4793,N_4495,N_4334);
xnor U4794 (N_4794,N_4417,N_4450);
nand U4795 (N_4795,N_4420,N_4279);
nand U4796 (N_4796,N_4377,N_4346);
and U4797 (N_4797,N_4305,N_4315);
nand U4798 (N_4798,N_4434,N_4227);
and U4799 (N_4799,N_4320,N_4322);
xnor U4800 (N_4800,N_4602,N_4660);
or U4801 (N_4801,N_4527,N_4793);
nor U4802 (N_4802,N_4657,N_4753);
or U4803 (N_4803,N_4693,N_4638);
xnor U4804 (N_4804,N_4726,N_4530);
nor U4805 (N_4805,N_4694,N_4731);
or U4806 (N_4806,N_4671,N_4666);
or U4807 (N_4807,N_4648,N_4763);
xor U4808 (N_4808,N_4784,N_4668);
and U4809 (N_4809,N_4709,N_4725);
nor U4810 (N_4810,N_4652,N_4552);
or U4811 (N_4811,N_4600,N_4727);
nand U4812 (N_4812,N_4594,N_4506);
nand U4813 (N_4813,N_4733,N_4697);
or U4814 (N_4814,N_4592,N_4670);
nor U4815 (N_4815,N_4584,N_4569);
nor U4816 (N_4816,N_4661,N_4580);
xor U4817 (N_4817,N_4768,N_4511);
or U4818 (N_4818,N_4729,N_4749);
xnor U4819 (N_4819,N_4528,N_4781);
nor U4820 (N_4820,N_4604,N_4581);
or U4821 (N_4821,N_4656,N_4790);
xnor U4822 (N_4822,N_4675,N_4708);
nand U4823 (N_4823,N_4543,N_4681);
xnor U4824 (N_4824,N_4537,N_4539);
or U4825 (N_4825,N_4767,N_4712);
xor U4826 (N_4826,N_4662,N_4780);
and U4827 (N_4827,N_4651,N_4746);
xor U4828 (N_4828,N_4667,N_4788);
xor U4829 (N_4829,N_4502,N_4514);
xnor U4830 (N_4830,N_4601,N_4633);
xor U4831 (N_4831,N_4717,N_4587);
nor U4832 (N_4832,N_4724,N_4771);
xor U4833 (N_4833,N_4605,N_4560);
or U4834 (N_4834,N_4586,N_4618);
nand U4835 (N_4835,N_4711,N_4567);
nand U4836 (N_4836,N_4553,N_4799);
or U4837 (N_4837,N_4555,N_4642);
xnor U4838 (N_4838,N_4565,N_4748);
nand U4839 (N_4839,N_4597,N_4765);
nor U4840 (N_4840,N_4645,N_4551);
or U4841 (N_4841,N_4625,N_4534);
nand U4842 (N_4842,N_4519,N_4538);
xor U4843 (N_4843,N_4698,N_4680);
or U4844 (N_4844,N_4540,N_4617);
nand U4845 (N_4845,N_4575,N_4745);
and U4846 (N_4846,N_4773,N_4623);
xnor U4847 (N_4847,N_4754,N_4785);
nor U4848 (N_4848,N_4619,N_4734);
or U4849 (N_4849,N_4524,N_4590);
and U4850 (N_4850,N_4732,N_4607);
nor U4851 (N_4851,N_4742,N_4568);
nand U4852 (N_4852,N_4710,N_4620);
nor U4853 (N_4853,N_4778,N_4704);
nand U4854 (N_4854,N_4699,N_4596);
and U4855 (N_4855,N_4783,N_4735);
nor U4856 (N_4856,N_4761,N_4676);
xnor U4857 (N_4857,N_4513,N_4701);
nor U4858 (N_4858,N_4639,N_4593);
and U4859 (N_4859,N_4595,N_4533);
and U4860 (N_4860,N_4603,N_4503);
or U4861 (N_4861,N_4797,N_4673);
or U4862 (N_4862,N_4689,N_4629);
nor U4863 (N_4863,N_4678,N_4787);
and U4864 (N_4864,N_4550,N_4556);
and U4865 (N_4865,N_4665,N_4641);
and U4866 (N_4866,N_4570,N_4792);
or U4867 (N_4867,N_4628,N_4504);
nor U4868 (N_4868,N_4614,N_4541);
and U4869 (N_4869,N_4782,N_4723);
nand U4870 (N_4870,N_4585,N_4544);
nor U4871 (N_4871,N_4624,N_4789);
nor U4872 (N_4872,N_4549,N_4566);
and U4873 (N_4873,N_4627,N_4647);
or U4874 (N_4874,N_4564,N_4622);
nand U4875 (N_4875,N_4578,N_4684);
nor U4876 (N_4876,N_4686,N_4561);
nand U4877 (N_4877,N_4518,N_4703);
and U4878 (N_4878,N_4545,N_4775);
nor U4879 (N_4879,N_4722,N_4509);
nand U4880 (N_4880,N_4598,N_4736);
and U4881 (N_4881,N_4643,N_4720);
nor U4882 (N_4882,N_4500,N_4691);
and U4883 (N_4883,N_4752,N_4571);
nor U4884 (N_4884,N_4547,N_4501);
xor U4885 (N_4885,N_4679,N_4772);
nor U4886 (N_4886,N_4756,N_4508);
xor U4887 (N_4887,N_4791,N_4608);
or U4888 (N_4888,N_4705,N_4616);
xor U4889 (N_4889,N_4672,N_4535);
xnor U4890 (N_4890,N_4505,N_4738);
and U4891 (N_4891,N_4626,N_4794);
and U4892 (N_4892,N_4612,N_4706);
and U4893 (N_4893,N_4589,N_4649);
and U4894 (N_4894,N_4690,N_4659);
and U4895 (N_4895,N_4507,N_4588);
or U4896 (N_4896,N_4515,N_4692);
nand U4897 (N_4897,N_4755,N_4750);
xnor U4898 (N_4898,N_4774,N_4687);
nor U4899 (N_4899,N_4523,N_4532);
xor U4900 (N_4900,N_4702,N_4653);
or U4901 (N_4901,N_4542,N_4522);
nor U4902 (N_4902,N_4635,N_4777);
xnor U4903 (N_4903,N_4707,N_4757);
nor U4904 (N_4904,N_4760,N_4719);
or U4905 (N_4905,N_4741,N_4525);
xnor U4906 (N_4906,N_4526,N_4510);
xnor U4907 (N_4907,N_4658,N_4636);
and U4908 (N_4908,N_4730,N_4721);
or U4909 (N_4909,N_4718,N_4786);
nand U4910 (N_4910,N_4517,N_4688);
and U4911 (N_4911,N_4613,N_4531);
and U4912 (N_4912,N_4737,N_4677);
nor U4913 (N_4913,N_4715,N_4574);
xor U4914 (N_4914,N_4770,N_4728);
and U4915 (N_4915,N_4714,N_4669);
and U4916 (N_4916,N_4512,N_4716);
nand U4917 (N_4917,N_4582,N_4634);
or U4918 (N_4918,N_4762,N_4674);
or U4919 (N_4919,N_4559,N_4536);
nand U4920 (N_4920,N_4664,N_4696);
nand U4921 (N_4921,N_4655,N_4743);
xnor U4922 (N_4922,N_4795,N_4798);
and U4923 (N_4923,N_4685,N_4621);
xnor U4924 (N_4924,N_4591,N_4739);
and U4925 (N_4925,N_4779,N_4529);
or U4926 (N_4926,N_4583,N_4577);
and U4927 (N_4927,N_4776,N_4713);
xnor U4928 (N_4928,N_4573,N_4650);
xnor U4929 (N_4929,N_4548,N_4644);
and U4930 (N_4930,N_4546,N_4599);
and U4931 (N_4931,N_4700,N_4683);
xor U4932 (N_4932,N_4579,N_4637);
nand U4933 (N_4933,N_4562,N_4682);
nand U4934 (N_4934,N_4521,N_4611);
nor U4935 (N_4935,N_4632,N_4747);
and U4936 (N_4936,N_4758,N_4516);
and U4937 (N_4937,N_4663,N_4764);
xnor U4938 (N_4938,N_4576,N_4520);
nand U4939 (N_4939,N_4615,N_4744);
and U4940 (N_4940,N_4796,N_4654);
nor U4941 (N_4941,N_4572,N_4751);
xor U4942 (N_4942,N_4631,N_4606);
or U4943 (N_4943,N_4630,N_4609);
nor U4944 (N_4944,N_4769,N_4558);
nand U4945 (N_4945,N_4640,N_4554);
nand U4946 (N_4946,N_4759,N_4557);
and U4947 (N_4947,N_4740,N_4563);
and U4948 (N_4948,N_4646,N_4695);
or U4949 (N_4949,N_4610,N_4766);
and U4950 (N_4950,N_4733,N_4604);
or U4951 (N_4951,N_4531,N_4514);
and U4952 (N_4952,N_4798,N_4606);
nor U4953 (N_4953,N_4782,N_4511);
or U4954 (N_4954,N_4727,N_4753);
nand U4955 (N_4955,N_4686,N_4527);
nor U4956 (N_4956,N_4741,N_4714);
or U4957 (N_4957,N_4606,N_4504);
or U4958 (N_4958,N_4736,N_4766);
nor U4959 (N_4959,N_4574,N_4655);
nand U4960 (N_4960,N_4579,N_4767);
and U4961 (N_4961,N_4635,N_4598);
and U4962 (N_4962,N_4583,N_4734);
or U4963 (N_4963,N_4514,N_4537);
nor U4964 (N_4964,N_4636,N_4720);
and U4965 (N_4965,N_4613,N_4632);
or U4966 (N_4966,N_4562,N_4600);
nand U4967 (N_4967,N_4675,N_4705);
xor U4968 (N_4968,N_4566,N_4628);
nor U4969 (N_4969,N_4776,N_4662);
and U4970 (N_4970,N_4682,N_4658);
nor U4971 (N_4971,N_4676,N_4726);
or U4972 (N_4972,N_4558,N_4691);
and U4973 (N_4973,N_4653,N_4617);
nor U4974 (N_4974,N_4646,N_4675);
and U4975 (N_4975,N_4735,N_4555);
nor U4976 (N_4976,N_4729,N_4681);
nor U4977 (N_4977,N_4701,N_4629);
xor U4978 (N_4978,N_4553,N_4507);
xor U4979 (N_4979,N_4791,N_4518);
or U4980 (N_4980,N_4652,N_4634);
or U4981 (N_4981,N_4659,N_4639);
and U4982 (N_4982,N_4778,N_4502);
nor U4983 (N_4983,N_4797,N_4550);
and U4984 (N_4984,N_4695,N_4616);
xor U4985 (N_4985,N_4521,N_4753);
nor U4986 (N_4986,N_4663,N_4513);
xnor U4987 (N_4987,N_4746,N_4605);
xnor U4988 (N_4988,N_4776,N_4762);
nand U4989 (N_4989,N_4753,N_4686);
and U4990 (N_4990,N_4654,N_4745);
or U4991 (N_4991,N_4587,N_4575);
or U4992 (N_4992,N_4753,N_4586);
nor U4993 (N_4993,N_4785,N_4631);
nand U4994 (N_4994,N_4613,N_4559);
xor U4995 (N_4995,N_4758,N_4693);
xor U4996 (N_4996,N_4749,N_4585);
xor U4997 (N_4997,N_4750,N_4618);
and U4998 (N_4998,N_4644,N_4507);
and U4999 (N_4999,N_4637,N_4550);
xor U5000 (N_5000,N_4753,N_4761);
or U5001 (N_5001,N_4561,N_4696);
xor U5002 (N_5002,N_4697,N_4705);
and U5003 (N_5003,N_4793,N_4570);
xnor U5004 (N_5004,N_4795,N_4504);
and U5005 (N_5005,N_4501,N_4703);
nand U5006 (N_5006,N_4563,N_4769);
xor U5007 (N_5007,N_4648,N_4716);
xnor U5008 (N_5008,N_4575,N_4549);
or U5009 (N_5009,N_4528,N_4732);
nand U5010 (N_5010,N_4691,N_4779);
nand U5011 (N_5011,N_4714,N_4773);
nor U5012 (N_5012,N_4781,N_4520);
nor U5013 (N_5013,N_4501,N_4573);
nand U5014 (N_5014,N_4698,N_4789);
xor U5015 (N_5015,N_4528,N_4677);
xor U5016 (N_5016,N_4521,N_4642);
or U5017 (N_5017,N_4672,N_4754);
nand U5018 (N_5018,N_4544,N_4573);
nor U5019 (N_5019,N_4596,N_4706);
xor U5020 (N_5020,N_4618,N_4633);
nor U5021 (N_5021,N_4687,N_4727);
nand U5022 (N_5022,N_4748,N_4741);
or U5023 (N_5023,N_4511,N_4523);
nor U5024 (N_5024,N_4566,N_4597);
or U5025 (N_5025,N_4538,N_4653);
xnor U5026 (N_5026,N_4555,N_4540);
nor U5027 (N_5027,N_4548,N_4688);
xnor U5028 (N_5028,N_4678,N_4608);
xnor U5029 (N_5029,N_4678,N_4515);
xnor U5030 (N_5030,N_4698,N_4791);
nand U5031 (N_5031,N_4781,N_4730);
and U5032 (N_5032,N_4575,N_4608);
and U5033 (N_5033,N_4564,N_4769);
or U5034 (N_5034,N_4730,N_4612);
and U5035 (N_5035,N_4657,N_4762);
xnor U5036 (N_5036,N_4628,N_4782);
or U5037 (N_5037,N_4524,N_4694);
nand U5038 (N_5038,N_4605,N_4653);
nand U5039 (N_5039,N_4656,N_4659);
nor U5040 (N_5040,N_4572,N_4726);
nand U5041 (N_5041,N_4791,N_4704);
nor U5042 (N_5042,N_4657,N_4538);
xor U5043 (N_5043,N_4514,N_4715);
or U5044 (N_5044,N_4638,N_4615);
and U5045 (N_5045,N_4772,N_4665);
xnor U5046 (N_5046,N_4534,N_4643);
nor U5047 (N_5047,N_4641,N_4668);
and U5048 (N_5048,N_4602,N_4651);
xor U5049 (N_5049,N_4514,N_4651);
nor U5050 (N_5050,N_4608,N_4562);
nor U5051 (N_5051,N_4718,N_4542);
and U5052 (N_5052,N_4755,N_4657);
nor U5053 (N_5053,N_4584,N_4619);
or U5054 (N_5054,N_4723,N_4687);
xnor U5055 (N_5055,N_4598,N_4535);
or U5056 (N_5056,N_4716,N_4544);
nand U5057 (N_5057,N_4692,N_4786);
nor U5058 (N_5058,N_4675,N_4557);
nand U5059 (N_5059,N_4770,N_4661);
and U5060 (N_5060,N_4572,N_4529);
nand U5061 (N_5061,N_4563,N_4684);
or U5062 (N_5062,N_4742,N_4669);
or U5063 (N_5063,N_4726,N_4668);
or U5064 (N_5064,N_4735,N_4580);
xnor U5065 (N_5065,N_4524,N_4532);
nor U5066 (N_5066,N_4788,N_4612);
xnor U5067 (N_5067,N_4745,N_4664);
or U5068 (N_5068,N_4525,N_4742);
nand U5069 (N_5069,N_4604,N_4555);
nand U5070 (N_5070,N_4644,N_4501);
nor U5071 (N_5071,N_4502,N_4733);
nor U5072 (N_5072,N_4762,N_4707);
nand U5073 (N_5073,N_4511,N_4629);
nor U5074 (N_5074,N_4737,N_4578);
and U5075 (N_5075,N_4636,N_4672);
xnor U5076 (N_5076,N_4776,N_4754);
and U5077 (N_5077,N_4626,N_4520);
nor U5078 (N_5078,N_4628,N_4727);
and U5079 (N_5079,N_4649,N_4795);
nand U5080 (N_5080,N_4540,N_4734);
nor U5081 (N_5081,N_4663,N_4589);
or U5082 (N_5082,N_4677,N_4610);
nand U5083 (N_5083,N_4783,N_4743);
or U5084 (N_5084,N_4562,N_4639);
nand U5085 (N_5085,N_4603,N_4617);
and U5086 (N_5086,N_4605,N_4683);
nor U5087 (N_5087,N_4688,N_4634);
or U5088 (N_5088,N_4534,N_4784);
xnor U5089 (N_5089,N_4552,N_4673);
and U5090 (N_5090,N_4764,N_4509);
nand U5091 (N_5091,N_4765,N_4676);
nor U5092 (N_5092,N_4612,N_4673);
or U5093 (N_5093,N_4758,N_4617);
or U5094 (N_5094,N_4759,N_4769);
or U5095 (N_5095,N_4700,N_4657);
nand U5096 (N_5096,N_4569,N_4505);
nand U5097 (N_5097,N_4626,N_4513);
xnor U5098 (N_5098,N_4736,N_4520);
and U5099 (N_5099,N_4604,N_4738);
nand U5100 (N_5100,N_4984,N_5033);
xnor U5101 (N_5101,N_4938,N_5008);
and U5102 (N_5102,N_4927,N_5056);
nand U5103 (N_5103,N_5070,N_5045);
nor U5104 (N_5104,N_4868,N_5089);
nand U5105 (N_5105,N_4903,N_4853);
nand U5106 (N_5106,N_4866,N_4967);
nor U5107 (N_5107,N_5090,N_5021);
and U5108 (N_5108,N_4851,N_5023);
and U5109 (N_5109,N_4857,N_4964);
xnor U5110 (N_5110,N_4965,N_4827);
nor U5111 (N_5111,N_5050,N_4836);
xnor U5112 (N_5112,N_4976,N_4961);
nand U5113 (N_5113,N_4824,N_5007);
xnor U5114 (N_5114,N_4814,N_5041);
or U5115 (N_5115,N_4915,N_4848);
xor U5116 (N_5116,N_5001,N_4881);
and U5117 (N_5117,N_5061,N_4818);
and U5118 (N_5118,N_5049,N_4820);
nor U5119 (N_5119,N_5003,N_4962);
nand U5120 (N_5120,N_4977,N_5087);
or U5121 (N_5121,N_5043,N_4929);
and U5122 (N_5122,N_5018,N_5011);
and U5123 (N_5123,N_5047,N_4804);
nand U5124 (N_5124,N_4901,N_5097);
and U5125 (N_5125,N_4988,N_4859);
nor U5126 (N_5126,N_4919,N_4801);
nor U5127 (N_5127,N_4909,N_4847);
nand U5128 (N_5128,N_5012,N_5009);
nand U5129 (N_5129,N_5060,N_4870);
xor U5130 (N_5130,N_5088,N_4995);
nand U5131 (N_5131,N_4849,N_4992);
and U5132 (N_5132,N_4913,N_4966);
nand U5133 (N_5133,N_4879,N_4939);
xor U5134 (N_5134,N_5024,N_5067);
nand U5135 (N_5135,N_4987,N_5096);
or U5136 (N_5136,N_4884,N_4980);
or U5137 (N_5137,N_4910,N_4816);
nor U5138 (N_5138,N_4960,N_5081);
and U5139 (N_5139,N_5030,N_4833);
nor U5140 (N_5140,N_5017,N_5057);
xnor U5141 (N_5141,N_4952,N_4872);
nor U5142 (N_5142,N_4994,N_4885);
xor U5143 (N_5143,N_4918,N_4823);
and U5144 (N_5144,N_4930,N_4907);
nor U5145 (N_5145,N_4944,N_4834);
or U5146 (N_5146,N_4817,N_5093);
xnor U5147 (N_5147,N_4946,N_4880);
nor U5148 (N_5148,N_5016,N_4899);
nor U5149 (N_5149,N_5072,N_4902);
or U5150 (N_5150,N_4940,N_4894);
nand U5151 (N_5151,N_4887,N_5055);
and U5152 (N_5152,N_4943,N_4810);
and U5153 (N_5153,N_4948,N_5080);
xor U5154 (N_5154,N_4945,N_5038);
and U5155 (N_5155,N_4972,N_5062);
nand U5156 (N_5156,N_5053,N_4954);
or U5157 (N_5157,N_4832,N_5025);
or U5158 (N_5158,N_5068,N_4809);
xor U5159 (N_5159,N_4921,N_4897);
xor U5160 (N_5160,N_4807,N_4981);
nand U5161 (N_5161,N_5022,N_5032);
nand U5162 (N_5162,N_4999,N_5000);
xnor U5163 (N_5163,N_5066,N_4911);
and U5164 (N_5164,N_4931,N_5034);
nand U5165 (N_5165,N_5054,N_4983);
xnor U5166 (N_5166,N_4850,N_4843);
and U5167 (N_5167,N_4996,N_4941);
or U5168 (N_5168,N_4878,N_4835);
or U5169 (N_5169,N_4861,N_4935);
nor U5170 (N_5170,N_4828,N_4844);
nor U5171 (N_5171,N_4985,N_4854);
or U5172 (N_5172,N_4819,N_4813);
nand U5173 (N_5173,N_4863,N_4989);
nor U5174 (N_5174,N_4974,N_4947);
or U5175 (N_5175,N_4846,N_5079);
or U5176 (N_5176,N_5059,N_4924);
and U5177 (N_5177,N_4963,N_4949);
nand U5178 (N_5178,N_4890,N_5065);
and U5179 (N_5179,N_4958,N_4839);
xor U5180 (N_5180,N_5075,N_4975);
xor U5181 (N_5181,N_4955,N_4803);
nor U5182 (N_5182,N_5014,N_4934);
nor U5183 (N_5183,N_5044,N_4959);
nand U5184 (N_5184,N_4875,N_4825);
xor U5185 (N_5185,N_4860,N_4877);
or U5186 (N_5186,N_5076,N_5082);
or U5187 (N_5187,N_4805,N_5015);
and U5188 (N_5188,N_4991,N_4882);
xnor U5189 (N_5189,N_5013,N_4842);
or U5190 (N_5190,N_4898,N_4971);
xnor U5191 (N_5191,N_5098,N_4951);
nor U5192 (N_5192,N_5095,N_4925);
and U5193 (N_5193,N_4855,N_4993);
nand U5194 (N_5194,N_4841,N_4942);
nand U5195 (N_5195,N_5084,N_4888);
nor U5196 (N_5196,N_4811,N_5029);
xnor U5197 (N_5197,N_4869,N_4908);
nand U5198 (N_5198,N_5036,N_4831);
nor U5199 (N_5199,N_4876,N_4895);
xor U5200 (N_5200,N_5028,N_4871);
and U5201 (N_5201,N_4812,N_5052);
and U5202 (N_5202,N_5051,N_5035);
and U5203 (N_5203,N_5005,N_4852);
or U5204 (N_5204,N_4969,N_4982);
nor U5205 (N_5205,N_4873,N_4891);
or U5206 (N_5206,N_5094,N_4917);
xnor U5207 (N_5207,N_5077,N_5085);
or U5208 (N_5208,N_4822,N_4900);
or U5209 (N_5209,N_4928,N_4874);
and U5210 (N_5210,N_5019,N_5020);
and U5211 (N_5211,N_5048,N_4906);
xnor U5212 (N_5212,N_4933,N_4802);
or U5213 (N_5213,N_4856,N_4916);
and U5214 (N_5214,N_4956,N_4926);
and U5215 (N_5215,N_5092,N_5099);
xnor U5216 (N_5216,N_4920,N_5091);
nor U5217 (N_5217,N_4950,N_5037);
or U5218 (N_5218,N_5010,N_5064);
nand U5219 (N_5219,N_4840,N_4837);
or U5220 (N_5220,N_4867,N_4973);
and U5221 (N_5221,N_4886,N_4829);
and U5222 (N_5222,N_4883,N_5002);
nand U5223 (N_5223,N_4845,N_5071);
or U5224 (N_5224,N_4978,N_4830);
and U5225 (N_5225,N_4970,N_4912);
or U5226 (N_5226,N_4937,N_5031);
nor U5227 (N_5227,N_4957,N_4905);
nand U5228 (N_5228,N_5078,N_4858);
or U5229 (N_5229,N_4986,N_4892);
nand U5230 (N_5230,N_4914,N_4864);
or U5231 (N_5231,N_4896,N_4862);
xnor U5232 (N_5232,N_4893,N_4998);
or U5233 (N_5233,N_5026,N_4923);
nor U5234 (N_5234,N_5058,N_4990);
nand U5235 (N_5235,N_4808,N_4953);
nor U5236 (N_5236,N_4800,N_4904);
xnor U5237 (N_5237,N_5004,N_5042);
or U5238 (N_5238,N_5086,N_4806);
and U5239 (N_5239,N_4815,N_5063);
nor U5240 (N_5240,N_4932,N_4865);
xor U5241 (N_5241,N_5040,N_4979);
nor U5242 (N_5242,N_5039,N_5006);
xor U5243 (N_5243,N_4936,N_5074);
nand U5244 (N_5244,N_4826,N_4968);
nand U5245 (N_5245,N_4838,N_5083);
nor U5246 (N_5246,N_5073,N_4821);
nand U5247 (N_5247,N_4922,N_5046);
or U5248 (N_5248,N_5069,N_4889);
nand U5249 (N_5249,N_4997,N_5027);
or U5250 (N_5250,N_4806,N_5070);
or U5251 (N_5251,N_4800,N_4803);
nand U5252 (N_5252,N_5019,N_5033);
nor U5253 (N_5253,N_5099,N_5097);
nand U5254 (N_5254,N_5090,N_4921);
nor U5255 (N_5255,N_4965,N_5049);
xor U5256 (N_5256,N_4829,N_4834);
nand U5257 (N_5257,N_4930,N_4953);
xor U5258 (N_5258,N_5069,N_4922);
nor U5259 (N_5259,N_5059,N_4943);
and U5260 (N_5260,N_4985,N_4935);
xor U5261 (N_5261,N_5082,N_4953);
nand U5262 (N_5262,N_4947,N_4823);
xnor U5263 (N_5263,N_4979,N_4949);
xnor U5264 (N_5264,N_4871,N_4944);
and U5265 (N_5265,N_4858,N_4901);
and U5266 (N_5266,N_5006,N_5080);
and U5267 (N_5267,N_4972,N_4840);
nand U5268 (N_5268,N_4838,N_4994);
or U5269 (N_5269,N_5062,N_4832);
nor U5270 (N_5270,N_5008,N_4944);
xor U5271 (N_5271,N_4953,N_4931);
nand U5272 (N_5272,N_4975,N_4919);
nand U5273 (N_5273,N_4801,N_5092);
xor U5274 (N_5274,N_4938,N_5024);
xor U5275 (N_5275,N_4910,N_4888);
nand U5276 (N_5276,N_4936,N_4937);
and U5277 (N_5277,N_4845,N_4915);
and U5278 (N_5278,N_4920,N_4978);
xor U5279 (N_5279,N_4844,N_4855);
xnor U5280 (N_5280,N_4896,N_4859);
or U5281 (N_5281,N_4805,N_4962);
nor U5282 (N_5282,N_5084,N_5076);
and U5283 (N_5283,N_5024,N_4875);
and U5284 (N_5284,N_4866,N_4997);
xor U5285 (N_5285,N_5086,N_4944);
nor U5286 (N_5286,N_5003,N_4894);
nor U5287 (N_5287,N_5055,N_4825);
nor U5288 (N_5288,N_5004,N_4919);
or U5289 (N_5289,N_4986,N_5057);
or U5290 (N_5290,N_4995,N_4816);
nand U5291 (N_5291,N_4862,N_4805);
and U5292 (N_5292,N_4976,N_5095);
nand U5293 (N_5293,N_5054,N_4942);
nor U5294 (N_5294,N_4831,N_5047);
or U5295 (N_5295,N_4975,N_4826);
nor U5296 (N_5296,N_5064,N_4850);
xnor U5297 (N_5297,N_4899,N_4904);
xnor U5298 (N_5298,N_5014,N_4948);
and U5299 (N_5299,N_4851,N_4847);
xnor U5300 (N_5300,N_4954,N_5062);
nand U5301 (N_5301,N_4978,N_4827);
nand U5302 (N_5302,N_5029,N_5069);
nand U5303 (N_5303,N_4881,N_4867);
and U5304 (N_5304,N_5029,N_4910);
and U5305 (N_5305,N_4978,N_4890);
and U5306 (N_5306,N_5007,N_4825);
xnor U5307 (N_5307,N_4995,N_4895);
nor U5308 (N_5308,N_5008,N_5049);
nor U5309 (N_5309,N_5038,N_5086);
nor U5310 (N_5310,N_4965,N_4917);
nor U5311 (N_5311,N_5050,N_4940);
or U5312 (N_5312,N_4887,N_5067);
nor U5313 (N_5313,N_4998,N_4915);
nor U5314 (N_5314,N_4903,N_4973);
xor U5315 (N_5315,N_5024,N_5047);
and U5316 (N_5316,N_4969,N_5071);
or U5317 (N_5317,N_5042,N_4831);
nand U5318 (N_5318,N_5021,N_4828);
or U5319 (N_5319,N_4884,N_5068);
xor U5320 (N_5320,N_4845,N_4932);
nor U5321 (N_5321,N_4862,N_4847);
nand U5322 (N_5322,N_5090,N_5020);
and U5323 (N_5323,N_4957,N_4974);
xnor U5324 (N_5324,N_5006,N_4816);
nor U5325 (N_5325,N_5061,N_4925);
xor U5326 (N_5326,N_5048,N_4857);
nor U5327 (N_5327,N_4824,N_5026);
or U5328 (N_5328,N_4820,N_4871);
nand U5329 (N_5329,N_5022,N_4856);
nor U5330 (N_5330,N_5032,N_4871);
and U5331 (N_5331,N_5024,N_4957);
and U5332 (N_5332,N_5048,N_4824);
nand U5333 (N_5333,N_4964,N_4937);
xnor U5334 (N_5334,N_4825,N_4974);
xor U5335 (N_5335,N_4838,N_5027);
nor U5336 (N_5336,N_4994,N_5030);
nor U5337 (N_5337,N_4821,N_4956);
xor U5338 (N_5338,N_4963,N_4986);
or U5339 (N_5339,N_5053,N_5010);
nand U5340 (N_5340,N_4904,N_4870);
or U5341 (N_5341,N_4835,N_4879);
and U5342 (N_5342,N_5046,N_4941);
nor U5343 (N_5343,N_4896,N_4829);
nor U5344 (N_5344,N_5046,N_4891);
or U5345 (N_5345,N_5099,N_4953);
and U5346 (N_5346,N_4883,N_4857);
or U5347 (N_5347,N_5080,N_4953);
or U5348 (N_5348,N_4806,N_5008);
nand U5349 (N_5349,N_4932,N_4968);
and U5350 (N_5350,N_4863,N_4909);
nand U5351 (N_5351,N_4853,N_5011);
nand U5352 (N_5352,N_4801,N_4944);
nor U5353 (N_5353,N_4832,N_4810);
xor U5354 (N_5354,N_4932,N_4870);
nor U5355 (N_5355,N_4813,N_5094);
and U5356 (N_5356,N_5018,N_4898);
and U5357 (N_5357,N_4850,N_4835);
nor U5358 (N_5358,N_4811,N_5096);
or U5359 (N_5359,N_4824,N_4996);
or U5360 (N_5360,N_5035,N_4996);
nor U5361 (N_5361,N_4956,N_4923);
nand U5362 (N_5362,N_5037,N_4842);
xnor U5363 (N_5363,N_5076,N_4899);
nand U5364 (N_5364,N_4827,N_4979);
or U5365 (N_5365,N_4913,N_5013);
xnor U5366 (N_5366,N_4897,N_5084);
nand U5367 (N_5367,N_4827,N_4833);
and U5368 (N_5368,N_5038,N_5025);
or U5369 (N_5369,N_4922,N_4854);
xnor U5370 (N_5370,N_4833,N_4975);
nor U5371 (N_5371,N_4960,N_4894);
or U5372 (N_5372,N_5059,N_5025);
and U5373 (N_5373,N_5062,N_4876);
nor U5374 (N_5374,N_4934,N_4975);
and U5375 (N_5375,N_5035,N_4944);
xor U5376 (N_5376,N_4972,N_4800);
nand U5377 (N_5377,N_4850,N_4976);
nor U5378 (N_5378,N_4948,N_5007);
nand U5379 (N_5379,N_4823,N_4939);
nand U5380 (N_5380,N_4817,N_4993);
and U5381 (N_5381,N_4826,N_4907);
and U5382 (N_5382,N_4896,N_5095);
and U5383 (N_5383,N_5000,N_5092);
or U5384 (N_5384,N_4950,N_5097);
xnor U5385 (N_5385,N_4975,N_4980);
nand U5386 (N_5386,N_4805,N_4819);
xor U5387 (N_5387,N_4895,N_4907);
xnor U5388 (N_5388,N_5049,N_4866);
nand U5389 (N_5389,N_5036,N_4806);
or U5390 (N_5390,N_4853,N_4812);
or U5391 (N_5391,N_5025,N_4852);
and U5392 (N_5392,N_5057,N_4995);
and U5393 (N_5393,N_4905,N_4941);
and U5394 (N_5394,N_4978,N_4941);
xnor U5395 (N_5395,N_5038,N_5096);
xnor U5396 (N_5396,N_4864,N_5064);
xnor U5397 (N_5397,N_5017,N_4896);
xnor U5398 (N_5398,N_5057,N_4801);
nor U5399 (N_5399,N_5041,N_4988);
xor U5400 (N_5400,N_5279,N_5320);
nor U5401 (N_5401,N_5384,N_5179);
nor U5402 (N_5402,N_5308,N_5131);
or U5403 (N_5403,N_5153,N_5157);
or U5404 (N_5404,N_5195,N_5228);
and U5405 (N_5405,N_5167,N_5247);
xor U5406 (N_5406,N_5250,N_5216);
or U5407 (N_5407,N_5102,N_5152);
nand U5408 (N_5408,N_5263,N_5106);
nor U5409 (N_5409,N_5118,N_5252);
nor U5410 (N_5410,N_5222,N_5124);
nand U5411 (N_5411,N_5382,N_5351);
or U5412 (N_5412,N_5150,N_5285);
or U5413 (N_5413,N_5380,N_5161);
nand U5414 (N_5414,N_5290,N_5293);
and U5415 (N_5415,N_5169,N_5260);
and U5416 (N_5416,N_5189,N_5353);
nand U5417 (N_5417,N_5211,N_5230);
nor U5418 (N_5418,N_5149,N_5237);
nor U5419 (N_5419,N_5256,N_5394);
xnor U5420 (N_5420,N_5192,N_5162);
and U5421 (N_5421,N_5392,N_5108);
and U5422 (N_5422,N_5141,N_5229);
and U5423 (N_5423,N_5313,N_5218);
nor U5424 (N_5424,N_5132,N_5205);
nor U5425 (N_5425,N_5369,N_5171);
nand U5426 (N_5426,N_5361,N_5238);
nor U5427 (N_5427,N_5133,N_5310);
and U5428 (N_5428,N_5284,N_5296);
or U5429 (N_5429,N_5219,N_5273);
xor U5430 (N_5430,N_5282,N_5289);
xor U5431 (N_5431,N_5348,N_5120);
and U5432 (N_5432,N_5375,N_5318);
nor U5433 (N_5433,N_5226,N_5220);
and U5434 (N_5434,N_5372,N_5266);
xor U5435 (N_5435,N_5387,N_5116);
nor U5436 (N_5436,N_5200,N_5378);
or U5437 (N_5437,N_5281,N_5350);
and U5438 (N_5438,N_5140,N_5286);
nand U5439 (N_5439,N_5180,N_5344);
and U5440 (N_5440,N_5271,N_5255);
and U5441 (N_5441,N_5213,N_5242);
nand U5442 (N_5442,N_5272,N_5374);
or U5443 (N_5443,N_5335,N_5144);
xnor U5444 (N_5444,N_5364,N_5340);
nor U5445 (N_5445,N_5154,N_5371);
nor U5446 (N_5446,N_5125,N_5101);
xnor U5447 (N_5447,N_5151,N_5166);
and U5448 (N_5448,N_5275,N_5197);
and U5449 (N_5449,N_5182,N_5309);
xnor U5450 (N_5450,N_5241,N_5183);
or U5451 (N_5451,N_5187,N_5277);
xnor U5452 (N_5452,N_5262,N_5323);
nand U5453 (N_5453,N_5163,N_5224);
or U5454 (N_5454,N_5155,N_5297);
nor U5455 (N_5455,N_5388,N_5209);
xor U5456 (N_5456,N_5345,N_5383);
nand U5457 (N_5457,N_5317,N_5215);
and U5458 (N_5458,N_5235,N_5236);
xor U5459 (N_5459,N_5134,N_5299);
or U5460 (N_5460,N_5186,N_5276);
nor U5461 (N_5461,N_5336,N_5304);
or U5462 (N_5462,N_5107,N_5145);
nand U5463 (N_5463,N_5331,N_5212);
nor U5464 (N_5464,N_5326,N_5135);
nor U5465 (N_5465,N_5160,N_5128);
nand U5466 (N_5466,N_5146,N_5334);
nor U5467 (N_5467,N_5324,N_5343);
nor U5468 (N_5468,N_5159,N_5176);
xnor U5469 (N_5469,N_5257,N_5319);
nand U5470 (N_5470,N_5370,N_5341);
nand U5471 (N_5471,N_5165,N_5258);
nor U5472 (N_5472,N_5329,N_5337);
and U5473 (N_5473,N_5253,N_5280);
and U5474 (N_5474,N_5203,N_5113);
or U5475 (N_5475,N_5181,N_5156);
xnor U5476 (N_5476,N_5129,N_5117);
or U5477 (N_5477,N_5349,N_5367);
and U5478 (N_5478,N_5379,N_5231);
and U5479 (N_5479,N_5254,N_5243);
nor U5480 (N_5480,N_5339,N_5190);
nand U5481 (N_5481,N_5201,N_5100);
or U5482 (N_5482,N_5206,N_5127);
nor U5483 (N_5483,N_5357,N_5112);
xor U5484 (N_5484,N_5330,N_5338);
xor U5485 (N_5485,N_5168,N_5245);
xnor U5486 (N_5486,N_5246,N_5325);
and U5487 (N_5487,N_5358,N_5104);
and U5488 (N_5488,N_5239,N_5225);
and U5489 (N_5489,N_5227,N_5223);
and U5490 (N_5490,N_5360,N_5199);
xor U5491 (N_5491,N_5119,N_5232);
nand U5492 (N_5492,N_5269,N_5322);
nor U5493 (N_5493,N_5139,N_5346);
and U5494 (N_5494,N_5312,N_5267);
nor U5495 (N_5495,N_5204,N_5207);
nor U5496 (N_5496,N_5302,N_5240);
xor U5497 (N_5497,N_5397,N_5355);
or U5498 (N_5498,N_5385,N_5158);
nor U5499 (N_5499,N_5311,N_5287);
or U5500 (N_5500,N_5261,N_5121);
or U5501 (N_5501,N_5214,N_5138);
and U5502 (N_5502,N_5178,N_5268);
and U5503 (N_5503,N_5303,N_5347);
or U5504 (N_5504,N_5298,N_5390);
nand U5505 (N_5505,N_5194,N_5115);
nand U5506 (N_5506,N_5359,N_5103);
nor U5507 (N_5507,N_5196,N_5316);
nor U5508 (N_5508,N_5210,N_5288);
and U5509 (N_5509,N_5193,N_5170);
and U5510 (N_5510,N_5399,N_5221);
nand U5511 (N_5511,N_5251,N_5362);
or U5512 (N_5512,N_5191,N_5174);
nor U5513 (N_5513,N_5314,N_5365);
and U5514 (N_5514,N_5185,N_5278);
nor U5515 (N_5515,N_5249,N_5248);
or U5516 (N_5516,N_5136,N_5300);
or U5517 (N_5517,N_5123,N_5109);
or U5518 (N_5518,N_5122,N_5332);
nand U5519 (N_5519,N_5327,N_5173);
xor U5520 (N_5520,N_5202,N_5164);
and U5521 (N_5521,N_5328,N_5377);
and U5522 (N_5522,N_5295,N_5233);
nand U5523 (N_5523,N_5142,N_5356);
and U5524 (N_5524,N_5148,N_5137);
nand U5525 (N_5525,N_5363,N_5175);
nor U5526 (N_5526,N_5188,N_5368);
xnor U5527 (N_5527,N_5147,N_5111);
and U5528 (N_5528,N_5172,N_5398);
and U5529 (N_5529,N_5386,N_5265);
and U5530 (N_5530,N_5315,N_5306);
nor U5531 (N_5531,N_5114,N_5291);
xnor U5532 (N_5532,N_5395,N_5110);
nand U5533 (N_5533,N_5393,N_5270);
nand U5534 (N_5534,N_5208,N_5321);
xor U5535 (N_5535,N_5105,N_5292);
nor U5536 (N_5536,N_5305,N_5294);
or U5537 (N_5537,N_5244,N_5366);
and U5538 (N_5538,N_5283,N_5354);
nor U5539 (N_5539,N_5274,N_5389);
nor U5540 (N_5540,N_5381,N_5217);
or U5541 (N_5541,N_5342,N_5376);
and U5542 (N_5542,N_5373,N_5184);
and U5543 (N_5543,N_5130,N_5301);
xor U5544 (N_5544,N_5177,N_5391);
nor U5545 (N_5545,N_5264,N_5333);
nand U5546 (N_5546,N_5234,N_5396);
nand U5547 (N_5547,N_5259,N_5143);
or U5548 (N_5548,N_5126,N_5307);
and U5549 (N_5549,N_5198,N_5352);
xnor U5550 (N_5550,N_5297,N_5234);
and U5551 (N_5551,N_5262,N_5187);
or U5552 (N_5552,N_5124,N_5259);
nor U5553 (N_5553,N_5109,N_5320);
or U5554 (N_5554,N_5320,N_5134);
nand U5555 (N_5555,N_5320,N_5283);
or U5556 (N_5556,N_5304,N_5133);
xnor U5557 (N_5557,N_5342,N_5110);
or U5558 (N_5558,N_5147,N_5362);
nand U5559 (N_5559,N_5325,N_5335);
and U5560 (N_5560,N_5105,N_5147);
nor U5561 (N_5561,N_5327,N_5365);
nor U5562 (N_5562,N_5195,N_5399);
nor U5563 (N_5563,N_5151,N_5218);
nor U5564 (N_5564,N_5297,N_5318);
and U5565 (N_5565,N_5371,N_5272);
or U5566 (N_5566,N_5375,N_5308);
xor U5567 (N_5567,N_5132,N_5146);
nand U5568 (N_5568,N_5271,N_5292);
xnor U5569 (N_5569,N_5280,N_5365);
and U5570 (N_5570,N_5299,N_5110);
xnor U5571 (N_5571,N_5335,N_5381);
nand U5572 (N_5572,N_5398,N_5315);
nor U5573 (N_5573,N_5360,N_5249);
nor U5574 (N_5574,N_5328,N_5257);
nand U5575 (N_5575,N_5194,N_5341);
nor U5576 (N_5576,N_5386,N_5125);
or U5577 (N_5577,N_5148,N_5273);
or U5578 (N_5578,N_5119,N_5214);
xnor U5579 (N_5579,N_5258,N_5110);
nor U5580 (N_5580,N_5174,N_5288);
nor U5581 (N_5581,N_5369,N_5356);
and U5582 (N_5582,N_5210,N_5372);
and U5583 (N_5583,N_5306,N_5191);
and U5584 (N_5584,N_5275,N_5289);
nor U5585 (N_5585,N_5301,N_5340);
nand U5586 (N_5586,N_5340,N_5240);
or U5587 (N_5587,N_5322,N_5154);
and U5588 (N_5588,N_5292,N_5351);
xor U5589 (N_5589,N_5232,N_5279);
or U5590 (N_5590,N_5236,N_5364);
or U5591 (N_5591,N_5388,N_5112);
or U5592 (N_5592,N_5147,N_5113);
xor U5593 (N_5593,N_5345,N_5316);
and U5594 (N_5594,N_5379,N_5323);
nor U5595 (N_5595,N_5229,N_5278);
nor U5596 (N_5596,N_5223,N_5129);
or U5597 (N_5597,N_5363,N_5145);
or U5598 (N_5598,N_5200,N_5360);
and U5599 (N_5599,N_5306,N_5192);
and U5600 (N_5600,N_5128,N_5201);
or U5601 (N_5601,N_5357,N_5165);
nand U5602 (N_5602,N_5380,N_5125);
nor U5603 (N_5603,N_5345,N_5352);
nor U5604 (N_5604,N_5310,N_5237);
xnor U5605 (N_5605,N_5387,N_5396);
nand U5606 (N_5606,N_5104,N_5387);
and U5607 (N_5607,N_5239,N_5130);
xor U5608 (N_5608,N_5280,N_5316);
nor U5609 (N_5609,N_5250,N_5395);
nand U5610 (N_5610,N_5357,N_5103);
nand U5611 (N_5611,N_5136,N_5258);
nand U5612 (N_5612,N_5282,N_5155);
nand U5613 (N_5613,N_5322,N_5184);
and U5614 (N_5614,N_5289,N_5328);
xnor U5615 (N_5615,N_5290,N_5132);
or U5616 (N_5616,N_5189,N_5110);
nand U5617 (N_5617,N_5187,N_5179);
and U5618 (N_5618,N_5291,N_5380);
xor U5619 (N_5619,N_5137,N_5151);
nand U5620 (N_5620,N_5343,N_5230);
or U5621 (N_5621,N_5281,N_5344);
xnor U5622 (N_5622,N_5114,N_5126);
nand U5623 (N_5623,N_5329,N_5260);
nor U5624 (N_5624,N_5247,N_5279);
xnor U5625 (N_5625,N_5303,N_5337);
and U5626 (N_5626,N_5223,N_5360);
and U5627 (N_5627,N_5174,N_5126);
nand U5628 (N_5628,N_5387,N_5379);
xnor U5629 (N_5629,N_5299,N_5129);
nor U5630 (N_5630,N_5204,N_5319);
and U5631 (N_5631,N_5292,N_5126);
xor U5632 (N_5632,N_5123,N_5378);
and U5633 (N_5633,N_5249,N_5346);
and U5634 (N_5634,N_5361,N_5197);
nor U5635 (N_5635,N_5189,N_5340);
xor U5636 (N_5636,N_5199,N_5354);
xor U5637 (N_5637,N_5123,N_5181);
or U5638 (N_5638,N_5397,N_5202);
or U5639 (N_5639,N_5367,N_5201);
and U5640 (N_5640,N_5391,N_5246);
nor U5641 (N_5641,N_5268,N_5224);
xor U5642 (N_5642,N_5162,N_5228);
or U5643 (N_5643,N_5104,N_5351);
or U5644 (N_5644,N_5280,N_5182);
xnor U5645 (N_5645,N_5226,N_5128);
nand U5646 (N_5646,N_5187,N_5330);
xnor U5647 (N_5647,N_5214,N_5204);
and U5648 (N_5648,N_5372,N_5339);
xnor U5649 (N_5649,N_5357,N_5232);
or U5650 (N_5650,N_5169,N_5275);
xor U5651 (N_5651,N_5106,N_5301);
nand U5652 (N_5652,N_5308,N_5339);
or U5653 (N_5653,N_5239,N_5211);
nand U5654 (N_5654,N_5213,N_5376);
xor U5655 (N_5655,N_5325,N_5181);
and U5656 (N_5656,N_5192,N_5102);
xnor U5657 (N_5657,N_5131,N_5259);
xor U5658 (N_5658,N_5375,N_5331);
xor U5659 (N_5659,N_5389,N_5237);
nor U5660 (N_5660,N_5379,N_5214);
nand U5661 (N_5661,N_5229,N_5174);
nor U5662 (N_5662,N_5367,N_5380);
xor U5663 (N_5663,N_5380,N_5285);
xor U5664 (N_5664,N_5369,N_5314);
and U5665 (N_5665,N_5322,N_5294);
nor U5666 (N_5666,N_5260,N_5314);
xor U5667 (N_5667,N_5220,N_5203);
nor U5668 (N_5668,N_5263,N_5318);
or U5669 (N_5669,N_5151,N_5114);
nand U5670 (N_5670,N_5285,N_5129);
and U5671 (N_5671,N_5382,N_5298);
nor U5672 (N_5672,N_5357,N_5325);
or U5673 (N_5673,N_5354,N_5163);
and U5674 (N_5674,N_5314,N_5391);
and U5675 (N_5675,N_5260,N_5211);
nand U5676 (N_5676,N_5260,N_5270);
nor U5677 (N_5677,N_5296,N_5216);
xor U5678 (N_5678,N_5177,N_5194);
or U5679 (N_5679,N_5100,N_5263);
nand U5680 (N_5680,N_5115,N_5387);
and U5681 (N_5681,N_5362,N_5215);
nor U5682 (N_5682,N_5211,N_5335);
nand U5683 (N_5683,N_5203,N_5157);
xor U5684 (N_5684,N_5322,N_5266);
nand U5685 (N_5685,N_5127,N_5257);
nor U5686 (N_5686,N_5359,N_5180);
and U5687 (N_5687,N_5331,N_5358);
or U5688 (N_5688,N_5148,N_5115);
nor U5689 (N_5689,N_5376,N_5179);
nor U5690 (N_5690,N_5211,N_5113);
and U5691 (N_5691,N_5116,N_5223);
nand U5692 (N_5692,N_5338,N_5198);
or U5693 (N_5693,N_5108,N_5251);
and U5694 (N_5694,N_5201,N_5226);
xor U5695 (N_5695,N_5351,N_5394);
xor U5696 (N_5696,N_5230,N_5183);
or U5697 (N_5697,N_5173,N_5315);
xnor U5698 (N_5698,N_5240,N_5379);
and U5699 (N_5699,N_5105,N_5205);
xor U5700 (N_5700,N_5654,N_5561);
xnor U5701 (N_5701,N_5668,N_5525);
or U5702 (N_5702,N_5593,N_5607);
or U5703 (N_5703,N_5510,N_5573);
nand U5704 (N_5704,N_5553,N_5449);
and U5705 (N_5705,N_5647,N_5436);
and U5706 (N_5706,N_5485,N_5591);
xnor U5707 (N_5707,N_5699,N_5680);
or U5708 (N_5708,N_5592,N_5685);
xnor U5709 (N_5709,N_5651,N_5583);
nand U5710 (N_5710,N_5434,N_5418);
xnor U5711 (N_5711,N_5567,N_5667);
or U5712 (N_5712,N_5536,N_5474);
and U5713 (N_5713,N_5601,N_5401);
nand U5714 (N_5714,N_5446,N_5657);
nor U5715 (N_5715,N_5422,N_5440);
nor U5716 (N_5716,N_5585,N_5495);
nor U5717 (N_5717,N_5546,N_5427);
or U5718 (N_5718,N_5649,N_5619);
and U5719 (N_5719,N_5673,N_5484);
or U5720 (N_5720,N_5527,N_5499);
and U5721 (N_5721,N_5448,N_5479);
or U5722 (N_5722,N_5468,N_5686);
or U5723 (N_5723,N_5611,N_5432);
or U5724 (N_5724,N_5571,N_5570);
nor U5725 (N_5725,N_5490,N_5429);
and U5726 (N_5726,N_5403,N_5450);
xnor U5727 (N_5727,N_5535,N_5617);
xor U5728 (N_5728,N_5579,N_5463);
nor U5729 (N_5729,N_5635,N_5589);
and U5730 (N_5730,N_5626,N_5497);
or U5731 (N_5731,N_5530,N_5698);
and U5732 (N_5732,N_5603,N_5409);
xnor U5733 (N_5733,N_5478,N_5400);
nor U5734 (N_5734,N_5564,N_5636);
xor U5735 (N_5735,N_5594,N_5630);
xor U5736 (N_5736,N_5684,N_5665);
nand U5737 (N_5737,N_5582,N_5671);
or U5738 (N_5738,N_5531,N_5565);
xnor U5739 (N_5739,N_5662,N_5599);
xnor U5740 (N_5740,N_5454,N_5445);
xor U5741 (N_5741,N_5515,N_5494);
nor U5742 (N_5742,N_5470,N_5595);
and U5743 (N_5743,N_5683,N_5508);
nand U5744 (N_5744,N_5580,N_5618);
or U5745 (N_5745,N_5509,N_5581);
nor U5746 (N_5746,N_5653,N_5514);
nor U5747 (N_5747,N_5419,N_5696);
xnor U5748 (N_5748,N_5614,N_5545);
nor U5749 (N_5749,N_5493,N_5458);
and U5750 (N_5750,N_5512,N_5532);
nand U5751 (N_5751,N_5424,N_5615);
or U5752 (N_5752,N_5669,N_5502);
and U5753 (N_5753,N_5522,N_5562);
nor U5754 (N_5754,N_5578,N_5656);
nand U5755 (N_5755,N_5690,N_5648);
nor U5756 (N_5756,N_5444,N_5439);
nor U5757 (N_5757,N_5623,N_5610);
or U5758 (N_5758,N_5670,N_5620);
nor U5759 (N_5759,N_5459,N_5542);
nand U5760 (N_5760,N_5658,N_5574);
xnor U5761 (N_5761,N_5586,N_5455);
nor U5762 (N_5762,N_5505,N_5628);
and U5763 (N_5763,N_5691,N_5412);
nand U5764 (N_5764,N_5489,N_5642);
or U5765 (N_5765,N_5451,N_5616);
xnor U5766 (N_5766,N_5520,N_5641);
nand U5767 (N_5767,N_5491,N_5661);
or U5768 (N_5768,N_5410,N_5548);
and U5769 (N_5769,N_5606,N_5472);
nand U5770 (N_5770,N_5576,N_5677);
or U5771 (N_5771,N_5694,N_5597);
or U5772 (N_5772,N_5453,N_5467);
xor U5773 (N_5773,N_5676,N_5513);
or U5774 (N_5774,N_5456,N_5442);
nand U5775 (N_5775,N_5693,N_5646);
or U5776 (N_5776,N_5469,N_5511);
xnor U5777 (N_5777,N_5621,N_5644);
or U5778 (N_5778,N_5689,N_5487);
xor U5779 (N_5779,N_5404,N_5645);
and U5780 (N_5780,N_5687,N_5602);
or U5781 (N_5781,N_5627,N_5678);
or U5782 (N_5782,N_5559,N_5555);
xor U5783 (N_5783,N_5584,N_5547);
nand U5784 (N_5784,N_5402,N_5457);
xor U5785 (N_5785,N_5550,N_5558);
nand U5786 (N_5786,N_5541,N_5568);
nand U5787 (N_5787,N_5590,N_5528);
and U5788 (N_5788,N_5475,N_5417);
nor U5789 (N_5789,N_5675,N_5416);
or U5790 (N_5790,N_5481,N_5435);
nand U5791 (N_5791,N_5441,N_5413);
xnor U5792 (N_5792,N_5486,N_5426);
nor U5793 (N_5793,N_5554,N_5517);
nand U5794 (N_5794,N_5674,N_5543);
nand U5795 (N_5795,N_5560,N_5544);
nand U5796 (N_5796,N_5430,N_5498);
xnor U5797 (N_5797,N_5516,N_5431);
nor U5798 (N_5798,N_5504,N_5697);
nor U5799 (N_5799,N_5428,N_5681);
nor U5800 (N_5800,N_5534,N_5643);
nand U5801 (N_5801,N_5473,N_5679);
or U5802 (N_5802,N_5682,N_5629);
and U5803 (N_5803,N_5652,N_5423);
xor U5804 (N_5804,N_5660,N_5462);
nand U5805 (N_5805,N_5460,N_5464);
and U5806 (N_5806,N_5538,N_5569);
nand U5807 (N_5807,N_5465,N_5411);
nor U5808 (N_5808,N_5443,N_5466);
xor U5809 (N_5809,N_5631,N_5414);
or U5810 (N_5810,N_5624,N_5471);
or U5811 (N_5811,N_5549,N_5612);
xor U5812 (N_5812,N_5655,N_5650);
xnor U5813 (N_5813,N_5526,N_5552);
and U5814 (N_5814,N_5604,N_5507);
or U5815 (N_5815,N_5421,N_5447);
and U5816 (N_5816,N_5577,N_5425);
and U5817 (N_5817,N_5625,N_5613);
and U5818 (N_5818,N_5663,N_5503);
nand U5819 (N_5819,N_5688,N_5537);
or U5820 (N_5820,N_5605,N_5415);
nor U5821 (N_5821,N_5608,N_5523);
nor U5822 (N_5822,N_5477,N_5540);
or U5823 (N_5823,N_5672,N_5461);
or U5824 (N_5824,N_5566,N_5407);
nand U5825 (N_5825,N_5488,N_5420);
and U5826 (N_5826,N_5588,N_5476);
nand U5827 (N_5827,N_5406,N_5695);
nor U5828 (N_5828,N_5632,N_5492);
nand U5829 (N_5829,N_5521,N_5533);
nand U5830 (N_5830,N_5572,N_5437);
nand U5831 (N_5831,N_5518,N_5557);
and U5832 (N_5832,N_5408,N_5452);
nor U5833 (N_5833,N_5539,N_5496);
or U5834 (N_5834,N_5634,N_5638);
and U5835 (N_5835,N_5405,N_5529);
and U5836 (N_5836,N_5563,N_5482);
xnor U5837 (N_5837,N_5633,N_5664);
and U5838 (N_5838,N_5501,N_5587);
nand U5839 (N_5839,N_5666,N_5692);
nand U5840 (N_5840,N_5596,N_5524);
nand U5841 (N_5841,N_5600,N_5659);
nand U5842 (N_5842,N_5483,N_5551);
and U5843 (N_5843,N_5575,N_5519);
and U5844 (N_5844,N_5480,N_5622);
or U5845 (N_5845,N_5433,N_5609);
nand U5846 (N_5846,N_5506,N_5637);
and U5847 (N_5847,N_5556,N_5500);
or U5848 (N_5848,N_5598,N_5640);
nor U5849 (N_5849,N_5438,N_5639);
and U5850 (N_5850,N_5679,N_5423);
or U5851 (N_5851,N_5437,N_5644);
xor U5852 (N_5852,N_5478,N_5693);
nand U5853 (N_5853,N_5667,N_5543);
xor U5854 (N_5854,N_5664,N_5551);
or U5855 (N_5855,N_5425,N_5669);
xor U5856 (N_5856,N_5663,N_5673);
or U5857 (N_5857,N_5423,N_5692);
and U5858 (N_5858,N_5577,N_5532);
and U5859 (N_5859,N_5615,N_5594);
or U5860 (N_5860,N_5573,N_5474);
and U5861 (N_5861,N_5572,N_5579);
nor U5862 (N_5862,N_5641,N_5600);
or U5863 (N_5863,N_5606,N_5639);
xor U5864 (N_5864,N_5429,N_5572);
xor U5865 (N_5865,N_5495,N_5689);
xor U5866 (N_5866,N_5411,N_5587);
nand U5867 (N_5867,N_5526,N_5600);
or U5868 (N_5868,N_5543,N_5425);
xor U5869 (N_5869,N_5524,N_5549);
or U5870 (N_5870,N_5410,N_5665);
and U5871 (N_5871,N_5490,N_5669);
nand U5872 (N_5872,N_5455,N_5539);
and U5873 (N_5873,N_5488,N_5425);
nor U5874 (N_5874,N_5486,N_5668);
nor U5875 (N_5875,N_5555,N_5542);
and U5876 (N_5876,N_5562,N_5594);
nand U5877 (N_5877,N_5593,N_5639);
nand U5878 (N_5878,N_5422,N_5415);
nand U5879 (N_5879,N_5538,N_5603);
and U5880 (N_5880,N_5471,N_5571);
nand U5881 (N_5881,N_5600,N_5537);
or U5882 (N_5882,N_5537,N_5579);
xor U5883 (N_5883,N_5406,N_5602);
xor U5884 (N_5884,N_5506,N_5517);
nor U5885 (N_5885,N_5455,N_5609);
xor U5886 (N_5886,N_5625,N_5566);
and U5887 (N_5887,N_5597,N_5640);
and U5888 (N_5888,N_5665,N_5661);
or U5889 (N_5889,N_5619,N_5691);
and U5890 (N_5890,N_5473,N_5491);
and U5891 (N_5891,N_5607,N_5566);
or U5892 (N_5892,N_5470,N_5685);
nand U5893 (N_5893,N_5610,N_5474);
nand U5894 (N_5894,N_5607,N_5606);
xor U5895 (N_5895,N_5477,N_5416);
nor U5896 (N_5896,N_5545,N_5523);
nor U5897 (N_5897,N_5512,N_5613);
xnor U5898 (N_5898,N_5445,N_5409);
nand U5899 (N_5899,N_5684,N_5500);
nand U5900 (N_5900,N_5634,N_5421);
and U5901 (N_5901,N_5427,N_5662);
nand U5902 (N_5902,N_5547,N_5616);
and U5903 (N_5903,N_5486,N_5504);
or U5904 (N_5904,N_5599,N_5541);
or U5905 (N_5905,N_5574,N_5569);
or U5906 (N_5906,N_5541,N_5504);
xor U5907 (N_5907,N_5655,N_5592);
nand U5908 (N_5908,N_5454,N_5658);
nor U5909 (N_5909,N_5699,N_5625);
or U5910 (N_5910,N_5519,N_5428);
or U5911 (N_5911,N_5482,N_5675);
xnor U5912 (N_5912,N_5659,N_5462);
xor U5913 (N_5913,N_5666,N_5459);
xnor U5914 (N_5914,N_5410,N_5540);
xnor U5915 (N_5915,N_5625,N_5444);
nand U5916 (N_5916,N_5411,N_5665);
nand U5917 (N_5917,N_5639,N_5507);
or U5918 (N_5918,N_5464,N_5658);
and U5919 (N_5919,N_5407,N_5485);
nor U5920 (N_5920,N_5577,N_5520);
and U5921 (N_5921,N_5528,N_5411);
or U5922 (N_5922,N_5660,N_5457);
or U5923 (N_5923,N_5486,N_5465);
xor U5924 (N_5924,N_5627,N_5409);
nor U5925 (N_5925,N_5545,N_5575);
nand U5926 (N_5926,N_5623,N_5657);
xnor U5927 (N_5927,N_5403,N_5580);
xnor U5928 (N_5928,N_5452,N_5573);
or U5929 (N_5929,N_5633,N_5533);
and U5930 (N_5930,N_5592,N_5484);
xnor U5931 (N_5931,N_5508,N_5433);
xnor U5932 (N_5932,N_5669,N_5555);
and U5933 (N_5933,N_5617,N_5661);
or U5934 (N_5934,N_5564,N_5541);
xor U5935 (N_5935,N_5543,N_5648);
xor U5936 (N_5936,N_5611,N_5464);
nand U5937 (N_5937,N_5607,N_5554);
nand U5938 (N_5938,N_5576,N_5681);
nand U5939 (N_5939,N_5409,N_5486);
or U5940 (N_5940,N_5520,N_5428);
nor U5941 (N_5941,N_5409,N_5544);
or U5942 (N_5942,N_5432,N_5677);
xor U5943 (N_5943,N_5542,N_5587);
nor U5944 (N_5944,N_5454,N_5408);
xnor U5945 (N_5945,N_5515,N_5416);
nor U5946 (N_5946,N_5574,N_5442);
nor U5947 (N_5947,N_5565,N_5456);
nor U5948 (N_5948,N_5612,N_5412);
nand U5949 (N_5949,N_5596,N_5667);
and U5950 (N_5950,N_5423,N_5412);
and U5951 (N_5951,N_5648,N_5445);
or U5952 (N_5952,N_5415,N_5513);
and U5953 (N_5953,N_5492,N_5566);
nand U5954 (N_5954,N_5688,N_5582);
and U5955 (N_5955,N_5533,N_5526);
and U5956 (N_5956,N_5603,N_5623);
xnor U5957 (N_5957,N_5698,N_5582);
and U5958 (N_5958,N_5632,N_5401);
nor U5959 (N_5959,N_5657,N_5616);
or U5960 (N_5960,N_5669,N_5607);
or U5961 (N_5961,N_5446,N_5426);
xnor U5962 (N_5962,N_5644,N_5588);
or U5963 (N_5963,N_5453,N_5406);
nor U5964 (N_5964,N_5433,N_5412);
nor U5965 (N_5965,N_5405,N_5583);
nand U5966 (N_5966,N_5526,N_5698);
and U5967 (N_5967,N_5684,N_5412);
nand U5968 (N_5968,N_5604,N_5564);
and U5969 (N_5969,N_5521,N_5436);
nor U5970 (N_5970,N_5545,N_5557);
xnor U5971 (N_5971,N_5559,N_5651);
xor U5972 (N_5972,N_5503,N_5427);
or U5973 (N_5973,N_5499,N_5623);
nand U5974 (N_5974,N_5575,N_5576);
and U5975 (N_5975,N_5570,N_5688);
or U5976 (N_5976,N_5615,N_5535);
or U5977 (N_5977,N_5526,N_5559);
nor U5978 (N_5978,N_5426,N_5650);
or U5979 (N_5979,N_5419,N_5421);
nor U5980 (N_5980,N_5578,N_5690);
nor U5981 (N_5981,N_5443,N_5664);
and U5982 (N_5982,N_5593,N_5598);
and U5983 (N_5983,N_5483,N_5630);
and U5984 (N_5984,N_5635,N_5549);
nor U5985 (N_5985,N_5634,N_5605);
xor U5986 (N_5986,N_5454,N_5554);
nand U5987 (N_5987,N_5423,N_5603);
xor U5988 (N_5988,N_5589,N_5699);
xnor U5989 (N_5989,N_5415,N_5568);
or U5990 (N_5990,N_5497,N_5538);
nor U5991 (N_5991,N_5585,N_5689);
or U5992 (N_5992,N_5637,N_5573);
or U5993 (N_5993,N_5456,N_5552);
nor U5994 (N_5994,N_5500,N_5480);
or U5995 (N_5995,N_5549,N_5609);
and U5996 (N_5996,N_5602,N_5563);
or U5997 (N_5997,N_5458,N_5401);
xnor U5998 (N_5998,N_5639,N_5681);
nor U5999 (N_5999,N_5517,N_5677);
xor U6000 (N_6000,N_5757,N_5994);
xor U6001 (N_6001,N_5988,N_5919);
nor U6002 (N_6002,N_5808,N_5874);
xnor U6003 (N_6003,N_5794,N_5811);
and U6004 (N_6004,N_5899,N_5873);
xor U6005 (N_6005,N_5776,N_5922);
xnor U6006 (N_6006,N_5796,N_5967);
nor U6007 (N_6007,N_5876,N_5774);
and U6008 (N_6008,N_5840,N_5886);
and U6009 (N_6009,N_5805,N_5845);
or U6010 (N_6010,N_5906,N_5832);
nand U6011 (N_6011,N_5931,N_5755);
nor U6012 (N_6012,N_5768,N_5918);
nor U6013 (N_6013,N_5907,N_5861);
nor U6014 (N_6014,N_5885,N_5712);
and U6015 (N_6015,N_5834,N_5766);
or U6016 (N_6016,N_5702,N_5833);
or U6017 (N_6017,N_5820,N_5891);
or U6018 (N_6018,N_5705,N_5802);
or U6019 (N_6019,N_5955,N_5842);
nand U6020 (N_6020,N_5806,N_5835);
nor U6021 (N_6021,N_5784,N_5945);
and U6022 (N_6022,N_5814,N_5782);
or U6023 (N_6023,N_5828,N_5844);
nor U6024 (N_6024,N_5853,N_5930);
xor U6025 (N_6025,N_5941,N_5747);
or U6026 (N_6026,N_5859,N_5979);
nand U6027 (N_6027,N_5895,N_5708);
or U6028 (N_6028,N_5860,N_5713);
nand U6029 (N_6029,N_5872,N_5952);
and U6030 (N_6030,N_5875,N_5966);
nand U6031 (N_6031,N_5924,N_5803);
nor U6032 (N_6032,N_5710,N_5908);
nor U6033 (N_6033,N_5877,N_5937);
and U6034 (N_6034,N_5946,N_5850);
and U6035 (N_6035,N_5778,N_5737);
xor U6036 (N_6036,N_5790,N_5995);
nor U6037 (N_6037,N_5986,N_5881);
and U6038 (N_6038,N_5989,N_5734);
nor U6039 (N_6039,N_5750,N_5838);
xor U6040 (N_6040,N_5701,N_5973);
or U6041 (N_6041,N_5735,N_5741);
nand U6042 (N_6042,N_5867,N_5816);
and U6043 (N_6043,N_5723,N_5773);
or U6044 (N_6044,N_5781,N_5731);
or U6045 (N_6045,N_5788,N_5926);
nand U6046 (N_6046,N_5896,N_5836);
and U6047 (N_6047,N_5999,N_5948);
xor U6048 (N_6048,N_5746,N_5754);
and U6049 (N_6049,N_5901,N_5958);
or U6050 (N_6050,N_5884,N_5717);
and U6051 (N_6051,N_5911,N_5865);
or U6052 (N_6052,N_5887,N_5858);
xnor U6053 (N_6053,N_5711,N_5951);
and U6054 (N_6054,N_5764,N_5954);
and U6055 (N_6055,N_5730,N_5719);
xor U6056 (N_6056,N_5866,N_5933);
nor U6057 (N_6057,N_5940,N_5990);
or U6058 (N_6058,N_5914,N_5787);
and U6059 (N_6059,N_5852,N_5943);
and U6060 (N_6060,N_5793,N_5785);
or U6061 (N_6061,N_5724,N_5831);
or U6062 (N_6062,N_5935,N_5738);
nor U6063 (N_6063,N_5942,N_5792);
nor U6064 (N_6064,N_5956,N_5978);
xor U6065 (N_6065,N_5976,N_5862);
nor U6066 (N_6066,N_5718,N_5917);
xor U6067 (N_6067,N_5704,N_5932);
xnor U6068 (N_6068,N_5703,N_5991);
xor U6069 (N_6069,N_5912,N_5900);
nand U6070 (N_6070,N_5714,N_5799);
nand U6071 (N_6071,N_5758,N_5936);
nor U6072 (N_6072,N_5759,N_5916);
xor U6073 (N_6073,N_5998,N_5837);
nor U6074 (N_6074,N_5753,N_5798);
nand U6075 (N_6075,N_5984,N_5733);
xor U6076 (N_6076,N_5771,N_5997);
nand U6077 (N_6077,N_5721,N_5846);
and U6078 (N_6078,N_5857,N_5920);
xor U6079 (N_6079,N_5740,N_5957);
nand U6080 (N_6080,N_5810,N_5789);
nand U6081 (N_6081,N_5934,N_5763);
xor U6082 (N_6082,N_5807,N_5851);
xnor U6083 (N_6083,N_5824,N_5909);
and U6084 (N_6084,N_5849,N_5826);
nor U6085 (N_6085,N_5823,N_5879);
or U6086 (N_6086,N_5728,N_5868);
nor U6087 (N_6087,N_5927,N_5707);
xor U6088 (N_6088,N_5777,N_5729);
xnor U6089 (N_6089,N_5751,N_5950);
and U6090 (N_6090,N_5791,N_5987);
and U6091 (N_6091,N_5739,N_5736);
nand U6092 (N_6092,N_5971,N_5812);
nor U6093 (N_6093,N_5725,N_5847);
xnor U6094 (N_6094,N_5970,N_5709);
or U6095 (N_6095,N_5779,N_5726);
and U6096 (N_6096,N_5815,N_5938);
nor U6097 (N_6097,N_5915,N_5897);
nor U6098 (N_6098,N_5761,N_5925);
or U6099 (N_6099,N_5921,N_5745);
xor U6100 (N_6100,N_5827,N_5821);
or U6101 (N_6101,N_5964,N_5928);
xnor U6102 (N_6102,N_5880,N_5772);
and U6103 (N_6103,N_5795,N_5818);
nand U6104 (N_6104,N_5848,N_5974);
and U6105 (N_6105,N_5817,N_5830);
nor U6106 (N_6106,N_5762,N_5720);
and U6107 (N_6107,N_5882,N_5975);
nor U6108 (N_6108,N_5947,N_5985);
or U6109 (N_6109,N_5904,N_5883);
nor U6110 (N_6110,N_5939,N_5804);
or U6111 (N_6111,N_5742,N_5786);
or U6112 (N_6112,N_5813,N_5983);
nand U6113 (N_6113,N_5890,N_5892);
xnor U6114 (N_6114,N_5878,N_5765);
nand U6115 (N_6115,N_5822,N_5825);
xnor U6116 (N_6116,N_5905,N_5962);
xor U6117 (N_6117,N_5749,N_5864);
nor U6118 (N_6118,N_5923,N_5969);
nand U6119 (N_6119,N_5929,N_5855);
and U6120 (N_6120,N_5700,N_5961);
and U6121 (N_6121,N_5902,N_5913);
xor U6122 (N_6122,N_5944,N_5727);
nand U6123 (N_6123,N_5870,N_5949);
or U6124 (N_6124,N_5769,N_5953);
xnor U6125 (N_6125,N_5841,N_5809);
xor U6126 (N_6126,N_5775,N_5843);
nand U6127 (N_6127,N_5722,N_5854);
nor U6128 (N_6128,N_5993,N_5992);
nand U6129 (N_6129,N_5819,N_5780);
nor U6130 (N_6130,N_5856,N_5888);
xnor U6131 (N_6131,N_5963,N_5871);
or U6132 (N_6132,N_5829,N_5903);
xor U6133 (N_6133,N_5715,N_5732);
nand U6134 (N_6134,N_5980,N_5839);
and U6135 (N_6135,N_5910,N_5756);
xor U6136 (N_6136,N_5960,N_5760);
nand U6137 (N_6137,N_5965,N_5863);
nor U6138 (N_6138,N_5959,N_5977);
nand U6139 (N_6139,N_5800,N_5706);
or U6140 (N_6140,N_5869,N_5797);
nand U6141 (N_6141,N_5968,N_5783);
and U6142 (N_6142,N_5748,N_5893);
nand U6143 (N_6143,N_5996,N_5898);
or U6144 (N_6144,N_5752,N_5889);
xor U6145 (N_6145,N_5982,N_5981);
or U6146 (N_6146,N_5972,N_5767);
nand U6147 (N_6147,N_5743,N_5770);
and U6148 (N_6148,N_5801,N_5744);
nor U6149 (N_6149,N_5716,N_5894);
or U6150 (N_6150,N_5994,N_5966);
or U6151 (N_6151,N_5855,N_5983);
xor U6152 (N_6152,N_5814,N_5775);
and U6153 (N_6153,N_5909,N_5713);
nand U6154 (N_6154,N_5886,N_5819);
nand U6155 (N_6155,N_5811,N_5786);
and U6156 (N_6156,N_5905,N_5921);
and U6157 (N_6157,N_5738,N_5927);
nand U6158 (N_6158,N_5897,N_5745);
nor U6159 (N_6159,N_5906,N_5861);
nand U6160 (N_6160,N_5823,N_5810);
or U6161 (N_6161,N_5926,N_5770);
and U6162 (N_6162,N_5841,N_5786);
or U6163 (N_6163,N_5922,N_5735);
nand U6164 (N_6164,N_5963,N_5902);
nand U6165 (N_6165,N_5727,N_5872);
xnor U6166 (N_6166,N_5754,N_5703);
and U6167 (N_6167,N_5866,N_5883);
nor U6168 (N_6168,N_5974,N_5834);
xor U6169 (N_6169,N_5782,N_5837);
or U6170 (N_6170,N_5866,N_5703);
or U6171 (N_6171,N_5938,N_5744);
xor U6172 (N_6172,N_5841,N_5924);
or U6173 (N_6173,N_5807,N_5968);
xnor U6174 (N_6174,N_5829,N_5948);
nor U6175 (N_6175,N_5862,N_5758);
and U6176 (N_6176,N_5975,N_5895);
nor U6177 (N_6177,N_5835,N_5863);
and U6178 (N_6178,N_5893,N_5773);
nand U6179 (N_6179,N_5807,N_5839);
nor U6180 (N_6180,N_5873,N_5856);
nor U6181 (N_6181,N_5861,N_5787);
xnor U6182 (N_6182,N_5729,N_5891);
nand U6183 (N_6183,N_5724,N_5960);
nand U6184 (N_6184,N_5988,N_5908);
nand U6185 (N_6185,N_5855,N_5718);
or U6186 (N_6186,N_5767,N_5834);
nand U6187 (N_6187,N_5713,N_5918);
nor U6188 (N_6188,N_5856,N_5726);
nand U6189 (N_6189,N_5852,N_5964);
nand U6190 (N_6190,N_5709,N_5743);
xor U6191 (N_6191,N_5704,N_5993);
nand U6192 (N_6192,N_5869,N_5912);
nor U6193 (N_6193,N_5757,N_5943);
xnor U6194 (N_6194,N_5749,N_5701);
xnor U6195 (N_6195,N_5833,N_5821);
xor U6196 (N_6196,N_5940,N_5917);
xor U6197 (N_6197,N_5938,N_5886);
or U6198 (N_6198,N_5969,N_5976);
nand U6199 (N_6199,N_5967,N_5753);
nand U6200 (N_6200,N_5971,N_5786);
and U6201 (N_6201,N_5821,N_5953);
or U6202 (N_6202,N_5762,N_5840);
nand U6203 (N_6203,N_5885,N_5807);
or U6204 (N_6204,N_5793,N_5797);
xor U6205 (N_6205,N_5709,N_5824);
nand U6206 (N_6206,N_5999,N_5858);
or U6207 (N_6207,N_5878,N_5736);
xnor U6208 (N_6208,N_5828,N_5929);
nand U6209 (N_6209,N_5910,N_5847);
nor U6210 (N_6210,N_5962,N_5779);
or U6211 (N_6211,N_5974,N_5962);
xnor U6212 (N_6212,N_5734,N_5744);
nand U6213 (N_6213,N_5799,N_5966);
or U6214 (N_6214,N_5764,N_5754);
xnor U6215 (N_6215,N_5759,N_5721);
nand U6216 (N_6216,N_5934,N_5841);
nor U6217 (N_6217,N_5874,N_5730);
nand U6218 (N_6218,N_5986,N_5783);
and U6219 (N_6219,N_5956,N_5761);
nand U6220 (N_6220,N_5899,N_5729);
nor U6221 (N_6221,N_5928,N_5783);
nor U6222 (N_6222,N_5770,N_5761);
nand U6223 (N_6223,N_5879,N_5933);
nand U6224 (N_6224,N_5862,N_5895);
or U6225 (N_6225,N_5808,N_5920);
nor U6226 (N_6226,N_5786,N_5720);
xnor U6227 (N_6227,N_5836,N_5845);
and U6228 (N_6228,N_5994,N_5852);
nand U6229 (N_6229,N_5995,N_5744);
nand U6230 (N_6230,N_5960,N_5998);
or U6231 (N_6231,N_5888,N_5869);
and U6232 (N_6232,N_5734,N_5713);
xor U6233 (N_6233,N_5836,N_5872);
nor U6234 (N_6234,N_5909,N_5703);
or U6235 (N_6235,N_5929,N_5909);
nor U6236 (N_6236,N_5756,N_5806);
nand U6237 (N_6237,N_5989,N_5772);
xnor U6238 (N_6238,N_5901,N_5847);
nor U6239 (N_6239,N_5735,N_5871);
nor U6240 (N_6240,N_5943,N_5889);
xnor U6241 (N_6241,N_5938,N_5860);
nand U6242 (N_6242,N_5873,N_5807);
xor U6243 (N_6243,N_5769,N_5820);
or U6244 (N_6244,N_5742,N_5968);
nor U6245 (N_6245,N_5761,N_5862);
and U6246 (N_6246,N_5845,N_5724);
nand U6247 (N_6247,N_5795,N_5727);
or U6248 (N_6248,N_5890,N_5853);
or U6249 (N_6249,N_5927,N_5897);
nand U6250 (N_6250,N_5866,N_5797);
xor U6251 (N_6251,N_5731,N_5772);
nand U6252 (N_6252,N_5936,N_5819);
or U6253 (N_6253,N_5987,N_5964);
and U6254 (N_6254,N_5854,N_5919);
nand U6255 (N_6255,N_5700,N_5771);
nand U6256 (N_6256,N_5799,N_5977);
nand U6257 (N_6257,N_5894,N_5943);
nand U6258 (N_6258,N_5823,N_5974);
or U6259 (N_6259,N_5812,N_5734);
xor U6260 (N_6260,N_5811,N_5947);
xor U6261 (N_6261,N_5947,N_5790);
xnor U6262 (N_6262,N_5797,N_5785);
nor U6263 (N_6263,N_5963,N_5992);
nor U6264 (N_6264,N_5804,N_5877);
or U6265 (N_6265,N_5930,N_5867);
or U6266 (N_6266,N_5858,N_5807);
xnor U6267 (N_6267,N_5906,N_5860);
nor U6268 (N_6268,N_5705,N_5764);
nand U6269 (N_6269,N_5792,N_5969);
nand U6270 (N_6270,N_5934,N_5837);
or U6271 (N_6271,N_5872,N_5931);
xnor U6272 (N_6272,N_5736,N_5703);
xor U6273 (N_6273,N_5827,N_5708);
or U6274 (N_6274,N_5960,N_5916);
xnor U6275 (N_6275,N_5833,N_5700);
xor U6276 (N_6276,N_5709,N_5732);
nor U6277 (N_6277,N_5744,N_5900);
xnor U6278 (N_6278,N_5883,N_5897);
nand U6279 (N_6279,N_5717,N_5834);
or U6280 (N_6280,N_5724,N_5957);
nor U6281 (N_6281,N_5789,N_5821);
xor U6282 (N_6282,N_5822,N_5900);
nor U6283 (N_6283,N_5933,N_5849);
and U6284 (N_6284,N_5718,N_5955);
xnor U6285 (N_6285,N_5770,N_5842);
nand U6286 (N_6286,N_5982,N_5866);
nor U6287 (N_6287,N_5712,N_5877);
nand U6288 (N_6288,N_5784,N_5771);
or U6289 (N_6289,N_5964,N_5974);
xor U6290 (N_6290,N_5881,N_5849);
or U6291 (N_6291,N_5979,N_5856);
and U6292 (N_6292,N_5926,N_5999);
nor U6293 (N_6293,N_5892,N_5973);
nor U6294 (N_6294,N_5798,N_5886);
nor U6295 (N_6295,N_5980,N_5708);
xor U6296 (N_6296,N_5933,N_5957);
nand U6297 (N_6297,N_5946,N_5761);
nand U6298 (N_6298,N_5904,N_5709);
nor U6299 (N_6299,N_5900,N_5884);
nor U6300 (N_6300,N_6110,N_6214);
or U6301 (N_6301,N_6235,N_6024);
nand U6302 (N_6302,N_6289,N_6074);
or U6303 (N_6303,N_6103,N_6100);
or U6304 (N_6304,N_6246,N_6185);
xor U6305 (N_6305,N_6046,N_6051);
nor U6306 (N_6306,N_6273,N_6233);
and U6307 (N_6307,N_6287,N_6044);
and U6308 (N_6308,N_6066,N_6174);
or U6309 (N_6309,N_6261,N_6231);
and U6310 (N_6310,N_6173,N_6114);
and U6311 (N_6311,N_6148,N_6128);
xnor U6312 (N_6312,N_6230,N_6172);
nand U6313 (N_6313,N_6236,N_6071);
nand U6314 (N_6314,N_6138,N_6149);
nor U6315 (N_6315,N_6256,N_6279);
nor U6316 (N_6316,N_6067,N_6035);
nand U6317 (N_6317,N_6033,N_6210);
nor U6318 (N_6318,N_6019,N_6225);
xor U6319 (N_6319,N_6107,N_6120);
xnor U6320 (N_6320,N_6147,N_6218);
and U6321 (N_6321,N_6018,N_6140);
or U6322 (N_6322,N_6102,N_6058);
nor U6323 (N_6323,N_6183,N_6027);
xnor U6324 (N_6324,N_6077,N_6284);
xor U6325 (N_6325,N_6178,N_6265);
nand U6326 (N_6326,N_6108,N_6157);
nand U6327 (N_6327,N_6245,N_6171);
nand U6328 (N_6328,N_6286,N_6132);
nor U6329 (N_6329,N_6264,N_6288);
or U6330 (N_6330,N_6168,N_6196);
nand U6331 (N_6331,N_6060,N_6032);
xor U6332 (N_6332,N_6091,N_6129);
or U6333 (N_6333,N_6179,N_6117);
or U6334 (N_6334,N_6036,N_6180);
and U6335 (N_6335,N_6283,N_6276);
or U6336 (N_6336,N_6099,N_6293);
nor U6337 (N_6337,N_6269,N_6258);
and U6338 (N_6338,N_6039,N_6251);
or U6339 (N_6339,N_6189,N_6270);
xor U6340 (N_6340,N_6267,N_6255);
and U6341 (N_6341,N_6104,N_6224);
nor U6342 (N_6342,N_6192,N_6041);
nand U6343 (N_6343,N_6217,N_6154);
nand U6344 (N_6344,N_6298,N_6134);
or U6345 (N_6345,N_6215,N_6026);
xnor U6346 (N_6346,N_6075,N_6028);
and U6347 (N_6347,N_6175,N_6169);
or U6348 (N_6348,N_6294,N_6199);
and U6349 (N_6349,N_6242,N_6042);
nor U6350 (N_6350,N_6228,N_6029);
and U6351 (N_6351,N_6112,N_6010);
nand U6352 (N_6352,N_6078,N_6272);
nor U6353 (N_6353,N_6278,N_6271);
and U6354 (N_6354,N_6291,N_6084);
or U6355 (N_6355,N_6054,N_6232);
or U6356 (N_6356,N_6122,N_6166);
and U6357 (N_6357,N_6127,N_6204);
and U6358 (N_6358,N_6106,N_6203);
xnor U6359 (N_6359,N_6249,N_6275);
and U6360 (N_6360,N_6038,N_6259);
nand U6361 (N_6361,N_6181,N_6105);
nand U6362 (N_6362,N_6266,N_6012);
nand U6363 (N_6363,N_6295,N_6186);
or U6364 (N_6364,N_6151,N_6123);
xor U6365 (N_6365,N_6088,N_6253);
nand U6366 (N_6366,N_6087,N_6167);
or U6367 (N_6367,N_6188,N_6119);
or U6368 (N_6368,N_6109,N_6197);
nand U6369 (N_6369,N_6222,N_6238);
xor U6370 (N_6370,N_6137,N_6263);
nor U6371 (N_6371,N_6209,N_6045);
or U6372 (N_6372,N_6096,N_6239);
and U6373 (N_6373,N_6205,N_6202);
or U6374 (N_6374,N_6011,N_6003);
nand U6375 (N_6375,N_6001,N_6195);
nand U6376 (N_6376,N_6257,N_6031);
and U6377 (N_6377,N_6097,N_6125);
nand U6378 (N_6378,N_6141,N_6290);
xnor U6379 (N_6379,N_6146,N_6130);
or U6380 (N_6380,N_6159,N_6229);
or U6381 (N_6381,N_6016,N_6143);
or U6382 (N_6382,N_6126,N_6030);
or U6383 (N_6383,N_6009,N_6206);
nand U6384 (N_6384,N_6013,N_6281);
nor U6385 (N_6385,N_6101,N_6017);
xor U6386 (N_6386,N_6144,N_6177);
nor U6387 (N_6387,N_6049,N_6182);
xnor U6388 (N_6388,N_6086,N_6212);
or U6389 (N_6389,N_6048,N_6296);
nand U6390 (N_6390,N_6111,N_6133);
and U6391 (N_6391,N_6135,N_6158);
xor U6392 (N_6392,N_6252,N_6007);
or U6393 (N_6393,N_6162,N_6082);
nor U6394 (N_6394,N_6247,N_6059);
nor U6395 (N_6395,N_6299,N_6220);
or U6396 (N_6396,N_6052,N_6150);
nand U6397 (N_6397,N_6089,N_6070);
xor U6398 (N_6398,N_6113,N_6211);
nor U6399 (N_6399,N_6098,N_6248);
nand U6400 (N_6400,N_6194,N_6040);
or U6401 (N_6401,N_6131,N_6241);
nor U6402 (N_6402,N_6223,N_6160);
xnor U6403 (N_6403,N_6201,N_6050);
or U6404 (N_6404,N_6187,N_6164);
xnor U6405 (N_6405,N_6118,N_6037);
nand U6406 (N_6406,N_6020,N_6240);
or U6407 (N_6407,N_6090,N_6093);
nor U6408 (N_6408,N_6285,N_6047);
nor U6409 (N_6409,N_6095,N_6083);
nand U6410 (N_6410,N_6190,N_6208);
xor U6411 (N_6411,N_6260,N_6002);
and U6412 (N_6412,N_6221,N_6092);
and U6413 (N_6413,N_6055,N_6081);
nand U6414 (N_6414,N_6142,N_6226);
or U6415 (N_6415,N_6065,N_6250);
nand U6416 (N_6416,N_6161,N_6198);
nand U6417 (N_6417,N_6085,N_6139);
nor U6418 (N_6418,N_6193,N_6080);
and U6419 (N_6419,N_6008,N_6282);
nor U6420 (N_6420,N_6297,N_6277);
and U6421 (N_6421,N_6163,N_6234);
or U6422 (N_6422,N_6227,N_6000);
or U6423 (N_6423,N_6219,N_6116);
xnor U6424 (N_6424,N_6237,N_6200);
and U6425 (N_6425,N_6053,N_6064);
nor U6426 (N_6426,N_6068,N_6184);
or U6427 (N_6427,N_6056,N_6170);
and U6428 (N_6428,N_6034,N_6274);
and U6429 (N_6429,N_6216,N_6262);
and U6430 (N_6430,N_6268,N_6244);
or U6431 (N_6431,N_6023,N_6156);
or U6432 (N_6432,N_6213,N_6165);
xnor U6433 (N_6433,N_6152,N_6004);
xor U6434 (N_6434,N_6025,N_6153);
and U6435 (N_6435,N_6014,N_6115);
xor U6436 (N_6436,N_6254,N_6292);
and U6437 (N_6437,N_6005,N_6072);
xnor U6438 (N_6438,N_6022,N_6076);
nor U6439 (N_6439,N_6121,N_6062);
nor U6440 (N_6440,N_6207,N_6043);
nor U6441 (N_6441,N_6136,N_6006);
and U6442 (N_6442,N_6057,N_6079);
or U6443 (N_6443,N_6061,N_6145);
or U6444 (N_6444,N_6094,N_6073);
nor U6445 (N_6445,N_6021,N_6069);
xor U6446 (N_6446,N_6191,N_6124);
nor U6447 (N_6447,N_6015,N_6243);
nand U6448 (N_6448,N_6063,N_6176);
xnor U6449 (N_6449,N_6155,N_6280);
and U6450 (N_6450,N_6216,N_6078);
xor U6451 (N_6451,N_6100,N_6166);
nand U6452 (N_6452,N_6163,N_6070);
nand U6453 (N_6453,N_6141,N_6006);
nor U6454 (N_6454,N_6241,N_6150);
nand U6455 (N_6455,N_6012,N_6066);
nor U6456 (N_6456,N_6120,N_6117);
xnor U6457 (N_6457,N_6145,N_6246);
and U6458 (N_6458,N_6093,N_6117);
or U6459 (N_6459,N_6299,N_6151);
xnor U6460 (N_6460,N_6129,N_6044);
nand U6461 (N_6461,N_6128,N_6243);
and U6462 (N_6462,N_6163,N_6039);
or U6463 (N_6463,N_6066,N_6094);
xnor U6464 (N_6464,N_6098,N_6043);
nor U6465 (N_6465,N_6110,N_6285);
or U6466 (N_6466,N_6109,N_6226);
and U6467 (N_6467,N_6118,N_6006);
and U6468 (N_6468,N_6181,N_6270);
nand U6469 (N_6469,N_6085,N_6206);
nand U6470 (N_6470,N_6198,N_6168);
or U6471 (N_6471,N_6254,N_6299);
xnor U6472 (N_6472,N_6092,N_6156);
xnor U6473 (N_6473,N_6018,N_6197);
and U6474 (N_6474,N_6101,N_6008);
xnor U6475 (N_6475,N_6222,N_6050);
xor U6476 (N_6476,N_6118,N_6244);
or U6477 (N_6477,N_6284,N_6259);
or U6478 (N_6478,N_6080,N_6272);
or U6479 (N_6479,N_6281,N_6138);
and U6480 (N_6480,N_6224,N_6098);
and U6481 (N_6481,N_6210,N_6271);
or U6482 (N_6482,N_6219,N_6051);
nand U6483 (N_6483,N_6163,N_6264);
and U6484 (N_6484,N_6072,N_6282);
or U6485 (N_6485,N_6234,N_6024);
nor U6486 (N_6486,N_6011,N_6135);
or U6487 (N_6487,N_6062,N_6264);
nor U6488 (N_6488,N_6046,N_6205);
xnor U6489 (N_6489,N_6150,N_6189);
nand U6490 (N_6490,N_6267,N_6061);
xnor U6491 (N_6491,N_6108,N_6125);
xor U6492 (N_6492,N_6055,N_6130);
and U6493 (N_6493,N_6143,N_6214);
nand U6494 (N_6494,N_6076,N_6079);
or U6495 (N_6495,N_6021,N_6033);
or U6496 (N_6496,N_6149,N_6014);
nand U6497 (N_6497,N_6022,N_6150);
or U6498 (N_6498,N_6098,N_6011);
nor U6499 (N_6499,N_6271,N_6012);
nand U6500 (N_6500,N_6015,N_6090);
nand U6501 (N_6501,N_6189,N_6297);
nand U6502 (N_6502,N_6262,N_6122);
and U6503 (N_6503,N_6223,N_6056);
or U6504 (N_6504,N_6092,N_6181);
and U6505 (N_6505,N_6206,N_6120);
or U6506 (N_6506,N_6137,N_6013);
xor U6507 (N_6507,N_6046,N_6066);
or U6508 (N_6508,N_6120,N_6103);
nand U6509 (N_6509,N_6173,N_6258);
and U6510 (N_6510,N_6057,N_6111);
nor U6511 (N_6511,N_6125,N_6191);
nand U6512 (N_6512,N_6227,N_6166);
nor U6513 (N_6513,N_6207,N_6257);
and U6514 (N_6514,N_6292,N_6112);
nand U6515 (N_6515,N_6124,N_6063);
nand U6516 (N_6516,N_6216,N_6179);
and U6517 (N_6517,N_6148,N_6298);
and U6518 (N_6518,N_6140,N_6032);
and U6519 (N_6519,N_6261,N_6284);
or U6520 (N_6520,N_6284,N_6124);
xnor U6521 (N_6521,N_6041,N_6053);
xor U6522 (N_6522,N_6213,N_6118);
or U6523 (N_6523,N_6264,N_6120);
or U6524 (N_6524,N_6193,N_6200);
nor U6525 (N_6525,N_6077,N_6282);
nor U6526 (N_6526,N_6050,N_6019);
nand U6527 (N_6527,N_6053,N_6267);
or U6528 (N_6528,N_6028,N_6195);
xor U6529 (N_6529,N_6035,N_6044);
or U6530 (N_6530,N_6095,N_6112);
nand U6531 (N_6531,N_6285,N_6208);
nor U6532 (N_6532,N_6010,N_6111);
or U6533 (N_6533,N_6265,N_6247);
nand U6534 (N_6534,N_6079,N_6129);
nor U6535 (N_6535,N_6084,N_6161);
nor U6536 (N_6536,N_6070,N_6063);
xnor U6537 (N_6537,N_6225,N_6179);
nand U6538 (N_6538,N_6138,N_6229);
xor U6539 (N_6539,N_6135,N_6064);
and U6540 (N_6540,N_6254,N_6141);
nand U6541 (N_6541,N_6048,N_6229);
xnor U6542 (N_6542,N_6117,N_6152);
and U6543 (N_6543,N_6249,N_6212);
or U6544 (N_6544,N_6189,N_6111);
nand U6545 (N_6545,N_6042,N_6135);
nand U6546 (N_6546,N_6082,N_6122);
or U6547 (N_6547,N_6087,N_6072);
nor U6548 (N_6548,N_6033,N_6194);
or U6549 (N_6549,N_6204,N_6034);
nor U6550 (N_6550,N_6025,N_6001);
nand U6551 (N_6551,N_6079,N_6040);
xor U6552 (N_6552,N_6105,N_6034);
nand U6553 (N_6553,N_6022,N_6237);
xnor U6554 (N_6554,N_6236,N_6264);
nor U6555 (N_6555,N_6154,N_6278);
xor U6556 (N_6556,N_6095,N_6285);
nand U6557 (N_6557,N_6254,N_6296);
and U6558 (N_6558,N_6115,N_6269);
nor U6559 (N_6559,N_6148,N_6065);
or U6560 (N_6560,N_6212,N_6141);
nand U6561 (N_6561,N_6049,N_6096);
nor U6562 (N_6562,N_6264,N_6278);
or U6563 (N_6563,N_6104,N_6027);
and U6564 (N_6564,N_6057,N_6141);
nand U6565 (N_6565,N_6267,N_6242);
xor U6566 (N_6566,N_6158,N_6252);
nor U6567 (N_6567,N_6223,N_6063);
or U6568 (N_6568,N_6046,N_6234);
nor U6569 (N_6569,N_6262,N_6157);
or U6570 (N_6570,N_6230,N_6040);
xnor U6571 (N_6571,N_6166,N_6051);
xor U6572 (N_6572,N_6231,N_6124);
and U6573 (N_6573,N_6267,N_6191);
nand U6574 (N_6574,N_6128,N_6289);
nand U6575 (N_6575,N_6047,N_6057);
or U6576 (N_6576,N_6114,N_6005);
nor U6577 (N_6577,N_6042,N_6083);
nor U6578 (N_6578,N_6037,N_6206);
or U6579 (N_6579,N_6252,N_6010);
or U6580 (N_6580,N_6152,N_6279);
nand U6581 (N_6581,N_6231,N_6008);
nor U6582 (N_6582,N_6203,N_6219);
or U6583 (N_6583,N_6020,N_6062);
nand U6584 (N_6584,N_6074,N_6144);
xor U6585 (N_6585,N_6083,N_6046);
nand U6586 (N_6586,N_6207,N_6195);
xnor U6587 (N_6587,N_6003,N_6088);
nand U6588 (N_6588,N_6244,N_6032);
xor U6589 (N_6589,N_6040,N_6224);
nor U6590 (N_6590,N_6053,N_6192);
nand U6591 (N_6591,N_6035,N_6127);
nor U6592 (N_6592,N_6134,N_6119);
or U6593 (N_6593,N_6041,N_6229);
and U6594 (N_6594,N_6046,N_6239);
xor U6595 (N_6595,N_6212,N_6275);
or U6596 (N_6596,N_6003,N_6117);
nand U6597 (N_6597,N_6166,N_6069);
xnor U6598 (N_6598,N_6014,N_6183);
and U6599 (N_6599,N_6042,N_6066);
nor U6600 (N_6600,N_6352,N_6328);
xnor U6601 (N_6601,N_6577,N_6310);
xnor U6602 (N_6602,N_6516,N_6460);
or U6603 (N_6603,N_6321,N_6312);
nor U6604 (N_6604,N_6594,N_6424);
nor U6605 (N_6605,N_6379,N_6375);
or U6606 (N_6606,N_6332,N_6430);
and U6607 (N_6607,N_6329,N_6392);
or U6608 (N_6608,N_6389,N_6349);
xnor U6609 (N_6609,N_6523,N_6432);
and U6610 (N_6610,N_6400,N_6452);
xnor U6611 (N_6611,N_6562,N_6308);
nand U6612 (N_6612,N_6489,N_6590);
xor U6613 (N_6613,N_6341,N_6428);
nand U6614 (N_6614,N_6313,N_6412);
or U6615 (N_6615,N_6326,N_6527);
nor U6616 (N_6616,N_6451,N_6592);
nor U6617 (N_6617,N_6338,N_6364);
and U6618 (N_6618,N_6539,N_6476);
nand U6619 (N_6619,N_6462,N_6355);
nand U6620 (N_6620,N_6384,N_6547);
xnor U6621 (N_6621,N_6518,N_6455);
and U6622 (N_6622,N_6560,N_6427);
or U6623 (N_6623,N_6550,N_6533);
xor U6624 (N_6624,N_6359,N_6507);
nand U6625 (N_6625,N_6433,N_6413);
and U6626 (N_6626,N_6382,N_6463);
xnor U6627 (N_6627,N_6544,N_6549);
nor U6628 (N_6628,N_6464,N_6469);
and U6629 (N_6629,N_6598,N_6351);
nor U6630 (N_6630,N_6457,N_6568);
xnor U6631 (N_6631,N_6512,N_6571);
nor U6632 (N_6632,N_6579,N_6330);
or U6633 (N_6633,N_6435,N_6542);
xnor U6634 (N_6634,N_6362,N_6487);
nor U6635 (N_6635,N_6481,N_6555);
and U6636 (N_6636,N_6575,N_6587);
nor U6637 (N_6637,N_6361,N_6311);
xnor U6638 (N_6638,N_6448,N_6509);
nand U6639 (N_6639,N_6365,N_6561);
or U6640 (N_6640,N_6386,N_6580);
nor U6641 (N_6641,N_6371,N_6459);
and U6642 (N_6642,N_6327,N_6565);
and U6643 (N_6643,N_6322,N_6508);
nor U6644 (N_6644,N_6342,N_6535);
xnor U6645 (N_6645,N_6445,N_6485);
xnor U6646 (N_6646,N_6343,N_6353);
and U6647 (N_6647,N_6356,N_6324);
or U6648 (N_6648,N_6500,N_6515);
and U6649 (N_6649,N_6395,N_6385);
and U6650 (N_6650,N_6543,N_6466);
nand U6651 (N_6651,N_6369,N_6490);
or U6652 (N_6652,N_6388,N_6554);
nor U6653 (N_6653,N_6557,N_6531);
xor U6654 (N_6654,N_6429,N_6537);
xor U6655 (N_6655,N_6406,N_6530);
nor U6656 (N_6656,N_6477,N_6563);
nor U6657 (N_6657,N_6529,N_6425);
and U6658 (N_6658,N_6446,N_6499);
xnor U6659 (N_6659,N_6434,N_6346);
xnor U6660 (N_6660,N_6556,N_6437);
nor U6661 (N_6661,N_6519,N_6569);
or U6662 (N_6662,N_6373,N_6378);
nor U6663 (N_6663,N_6447,N_6300);
and U6664 (N_6664,N_6407,N_6302);
nand U6665 (N_6665,N_6454,N_6528);
nor U6666 (N_6666,N_6586,N_6393);
xnor U6667 (N_6667,N_6301,N_6405);
xor U6668 (N_6668,N_6572,N_6478);
xor U6669 (N_6669,N_6497,N_6504);
or U6670 (N_6670,N_6370,N_6409);
or U6671 (N_6671,N_6410,N_6488);
or U6672 (N_6672,N_6416,N_6576);
and U6673 (N_6673,N_6304,N_6503);
or U6674 (N_6674,N_6599,N_6415);
xnor U6675 (N_6675,N_6306,N_6559);
or U6676 (N_6676,N_6414,N_6450);
nor U6677 (N_6677,N_6491,N_6525);
nor U6678 (N_6678,N_6468,N_6501);
or U6679 (N_6679,N_6502,N_6358);
nand U6680 (N_6680,N_6418,N_6588);
or U6681 (N_6681,N_6426,N_6540);
or U6682 (N_6682,N_6458,N_6526);
nor U6683 (N_6683,N_6408,N_6583);
nand U6684 (N_6684,N_6398,N_6517);
xor U6685 (N_6685,N_6484,N_6366);
xor U6686 (N_6686,N_6318,N_6381);
or U6687 (N_6687,N_6551,N_6335);
or U6688 (N_6688,N_6337,N_6316);
and U6689 (N_6689,N_6475,N_6474);
nor U6690 (N_6690,N_6564,N_6574);
xor U6691 (N_6691,N_6320,N_6354);
or U6692 (N_6692,N_6520,N_6506);
nor U6693 (N_6693,N_6566,N_6511);
nor U6694 (N_6694,N_6480,N_6431);
and U6695 (N_6695,N_6470,N_6585);
nor U6696 (N_6696,N_6548,N_6495);
nor U6697 (N_6697,N_6317,N_6441);
or U6698 (N_6698,N_6344,N_6319);
nor U6699 (N_6699,N_6394,N_6325);
or U6700 (N_6700,N_6545,N_6350);
and U6701 (N_6701,N_6348,N_6403);
or U6702 (N_6702,N_6305,N_6391);
xnor U6703 (N_6703,N_6496,N_6536);
and U6704 (N_6704,N_6376,N_6473);
xor U6705 (N_6705,N_6380,N_6584);
xor U6706 (N_6706,N_6315,N_6534);
nand U6707 (N_6707,N_6417,N_6510);
xor U6708 (N_6708,N_6336,N_6593);
or U6709 (N_6709,N_6493,N_6582);
nor U6710 (N_6710,N_6479,N_6422);
or U6711 (N_6711,N_6595,N_6521);
and U6712 (N_6712,N_6423,N_6461);
or U6713 (N_6713,N_6339,N_6513);
and U6714 (N_6714,N_6401,N_6390);
xor U6715 (N_6715,N_6522,N_6372);
and U6716 (N_6716,N_6442,N_6387);
and U6717 (N_6717,N_6333,N_6597);
and U6718 (N_6718,N_6449,N_6570);
nor U6719 (N_6719,N_6397,N_6314);
nor U6720 (N_6720,N_6552,N_6309);
and U6721 (N_6721,N_6363,N_6581);
or U6722 (N_6722,N_6472,N_6483);
or U6723 (N_6723,N_6402,N_6546);
xnor U6724 (N_6724,N_6347,N_6443);
xor U6725 (N_6725,N_6492,N_6368);
nand U6726 (N_6726,N_6399,N_6383);
or U6727 (N_6727,N_6538,N_6334);
nor U6728 (N_6728,N_6573,N_6465);
xnor U6729 (N_6729,N_6486,N_6360);
nand U6730 (N_6730,N_6420,N_6553);
or U6731 (N_6731,N_6456,N_6331);
and U6732 (N_6732,N_6377,N_6357);
xor U6733 (N_6733,N_6421,N_6567);
xnor U6734 (N_6734,N_6578,N_6411);
nor U6735 (N_6735,N_6367,N_6453);
xor U6736 (N_6736,N_6498,N_6438);
or U6737 (N_6737,N_6396,N_6345);
nor U6738 (N_6738,N_6482,N_6323);
xor U6739 (N_6739,N_6558,N_6591);
nand U6740 (N_6740,N_6596,N_6436);
and U6741 (N_6741,N_6444,N_6467);
nor U6742 (N_6742,N_6532,N_6471);
and U6743 (N_6743,N_6514,N_6340);
xor U6744 (N_6744,N_6589,N_6439);
nand U6745 (N_6745,N_6374,N_6419);
and U6746 (N_6746,N_6303,N_6494);
nor U6747 (N_6747,N_6440,N_6505);
nor U6748 (N_6748,N_6541,N_6307);
nor U6749 (N_6749,N_6404,N_6524);
xnor U6750 (N_6750,N_6567,N_6586);
or U6751 (N_6751,N_6567,N_6442);
and U6752 (N_6752,N_6548,N_6563);
and U6753 (N_6753,N_6335,N_6583);
nor U6754 (N_6754,N_6304,N_6494);
nor U6755 (N_6755,N_6304,N_6303);
or U6756 (N_6756,N_6305,N_6399);
and U6757 (N_6757,N_6433,N_6363);
xnor U6758 (N_6758,N_6304,N_6448);
nand U6759 (N_6759,N_6452,N_6354);
nor U6760 (N_6760,N_6314,N_6480);
and U6761 (N_6761,N_6558,N_6355);
or U6762 (N_6762,N_6483,N_6587);
and U6763 (N_6763,N_6303,N_6300);
nand U6764 (N_6764,N_6585,N_6477);
nor U6765 (N_6765,N_6456,N_6504);
and U6766 (N_6766,N_6451,N_6522);
and U6767 (N_6767,N_6544,N_6588);
nor U6768 (N_6768,N_6306,N_6372);
and U6769 (N_6769,N_6555,N_6491);
and U6770 (N_6770,N_6599,N_6442);
and U6771 (N_6771,N_6574,N_6386);
or U6772 (N_6772,N_6335,N_6488);
nor U6773 (N_6773,N_6385,N_6536);
xor U6774 (N_6774,N_6351,N_6360);
nor U6775 (N_6775,N_6446,N_6452);
nor U6776 (N_6776,N_6595,N_6465);
nor U6777 (N_6777,N_6416,N_6580);
xnor U6778 (N_6778,N_6580,N_6379);
nand U6779 (N_6779,N_6567,N_6367);
nand U6780 (N_6780,N_6332,N_6566);
and U6781 (N_6781,N_6595,N_6377);
and U6782 (N_6782,N_6413,N_6556);
or U6783 (N_6783,N_6585,N_6302);
xnor U6784 (N_6784,N_6580,N_6381);
xor U6785 (N_6785,N_6562,N_6399);
or U6786 (N_6786,N_6323,N_6405);
nand U6787 (N_6787,N_6380,N_6395);
nand U6788 (N_6788,N_6342,N_6596);
xor U6789 (N_6789,N_6486,N_6477);
nand U6790 (N_6790,N_6388,N_6359);
nand U6791 (N_6791,N_6402,N_6447);
or U6792 (N_6792,N_6554,N_6347);
and U6793 (N_6793,N_6522,N_6325);
or U6794 (N_6794,N_6302,N_6354);
xor U6795 (N_6795,N_6372,N_6361);
nor U6796 (N_6796,N_6400,N_6325);
nor U6797 (N_6797,N_6471,N_6594);
nand U6798 (N_6798,N_6365,N_6520);
or U6799 (N_6799,N_6340,N_6391);
nor U6800 (N_6800,N_6541,N_6358);
xor U6801 (N_6801,N_6432,N_6395);
or U6802 (N_6802,N_6428,N_6440);
nor U6803 (N_6803,N_6386,N_6495);
xor U6804 (N_6804,N_6352,N_6565);
nor U6805 (N_6805,N_6513,N_6549);
or U6806 (N_6806,N_6591,N_6522);
and U6807 (N_6807,N_6312,N_6450);
xnor U6808 (N_6808,N_6463,N_6551);
xnor U6809 (N_6809,N_6346,N_6478);
nor U6810 (N_6810,N_6444,N_6385);
and U6811 (N_6811,N_6480,N_6570);
and U6812 (N_6812,N_6593,N_6457);
xnor U6813 (N_6813,N_6485,N_6570);
xnor U6814 (N_6814,N_6449,N_6536);
or U6815 (N_6815,N_6594,N_6590);
nand U6816 (N_6816,N_6310,N_6389);
nor U6817 (N_6817,N_6341,N_6505);
xnor U6818 (N_6818,N_6355,N_6544);
nor U6819 (N_6819,N_6357,N_6522);
xor U6820 (N_6820,N_6315,N_6551);
nand U6821 (N_6821,N_6315,N_6429);
nor U6822 (N_6822,N_6377,N_6445);
or U6823 (N_6823,N_6413,N_6563);
nor U6824 (N_6824,N_6406,N_6439);
nor U6825 (N_6825,N_6598,N_6560);
nand U6826 (N_6826,N_6547,N_6507);
nand U6827 (N_6827,N_6364,N_6464);
or U6828 (N_6828,N_6513,N_6331);
nand U6829 (N_6829,N_6367,N_6396);
or U6830 (N_6830,N_6399,N_6302);
nand U6831 (N_6831,N_6302,N_6520);
xnor U6832 (N_6832,N_6322,N_6455);
and U6833 (N_6833,N_6550,N_6596);
or U6834 (N_6834,N_6309,N_6331);
xnor U6835 (N_6835,N_6364,N_6579);
nand U6836 (N_6836,N_6584,N_6401);
xnor U6837 (N_6837,N_6438,N_6584);
nor U6838 (N_6838,N_6452,N_6487);
nand U6839 (N_6839,N_6497,N_6451);
nor U6840 (N_6840,N_6484,N_6398);
or U6841 (N_6841,N_6573,N_6413);
nand U6842 (N_6842,N_6316,N_6489);
xnor U6843 (N_6843,N_6427,N_6483);
nand U6844 (N_6844,N_6334,N_6412);
and U6845 (N_6845,N_6488,N_6381);
nor U6846 (N_6846,N_6498,N_6415);
xnor U6847 (N_6847,N_6360,N_6539);
or U6848 (N_6848,N_6304,N_6405);
nor U6849 (N_6849,N_6326,N_6398);
or U6850 (N_6850,N_6477,N_6364);
nand U6851 (N_6851,N_6414,N_6572);
and U6852 (N_6852,N_6587,N_6361);
nor U6853 (N_6853,N_6472,N_6575);
nand U6854 (N_6854,N_6534,N_6339);
xnor U6855 (N_6855,N_6344,N_6367);
nand U6856 (N_6856,N_6337,N_6462);
and U6857 (N_6857,N_6391,N_6576);
or U6858 (N_6858,N_6356,N_6466);
or U6859 (N_6859,N_6471,N_6416);
and U6860 (N_6860,N_6384,N_6372);
xnor U6861 (N_6861,N_6343,N_6594);
and U6862 (N_6862,N_6578,N_6475);
or U6863 (N_6863,N_6355,N_6512);
nor U6864 (N_6864,N_6331,N_6595);
nand U6865 (N_6865,N_6568,N_6561);
or U6866 (N_6866,N_6593,N_6530);
nor U6867 (N_6867,N_6502,N_6354);
or U6868 (N_6868,N_6444,N_6402);
or U6869 (N_6869,N_6306,N_6355);
and U6870 (N_6870,N_6393,N_6322);
and U6871 (N_6871,N_6501,N_6557);
and U6872 (N_6872,N_6384,N_6312);
nor U6873 (N_6873,N_6590,N_6525);
nand U6874 (N_6874,N_6510,N_6546);
nand U6875 (N_6875,N_6581,N_6509);
and U6876 (N_6876,N_6517,N_6411);
nor U6877 (N_6877,N_6574,N_6317);
xor U6878 (N_6878,N_6524,N_6426);
and U6879 (N_6879,N_6542,N_6362);
or U6880 (N_6880,N_6554,N_6478);
nand U6881 (N_6881,N_6499,N_6400);
nor U6882 (N_6882,N_6406,N_6550);
xnor U6883 (N_6883,N_6461,N_6394);
nand U6884 (N_6884,N_6482,N_6458);
nor U6885 (N_6885,N_6538,N_6593);
and U6886 (N_6886,N_6548,N_6345);
nand U6887 (N_6887,N_6350,N_6335);
xnor U6888 (N_6888,N_6533,N_6367);
nor U6889 (N_6889,N_6300,N_6409);
and U6890 (N_6890,N_6505,N_6527);
and U6891 (N_6891,N_6589,N_6534);
nor U6892 (N_6892,N_6598,N_6366);
nand U6893 (N_6893,N_6522,N_6467);
nor U6894 (N_6894,N_6565,N_6308);
xnor U6895 (N_6895,N_6467,N_6441);
and U6896 (N_6896,N_6584,N_6317);
nand U6897 (N_6897,N_6568,N_6555);
xor U6898 (N_6898,N_6382,N_6542);
or U6899 (N_6899,N_6401,N_6530);
or U6900 (N_6900,N_6855,N_6812);
nor U6901 (N_6901,N_6691,N_6898);
or U6902 (N_6902,N_6840,N_6872);
nand U6903 (N_6903,N_6636,N_6697);
nand U6904 (N_6904,N_6686,N_6658);
xor U6905 (N_6905,N_6749,N_6874);
nand U6906 (N_6906,N_6716,N_6663);
and U6907 (N_6907,N_6746,N_6837);
and U6908 (N_6908,N_6611,N_6679);
and U6909 (N_6909,N_6865,N_6635);
and U6910 (N_6910,N_6754,N_6878);
and U6911 (N_6911,N_6876,N_6816);
nor U6912 (N_6912,N_6677,N_6825);
xor U6913 (N_6913,N_6850,N_6775);
nor U6914 (N_6914,N_6701,N_6639);
or U6915 (N_6915,N_6700,N_6612);
and U6916 (N_6916,N_6732,N_6610);
xor U6917 (N_6917,N_6854,N_6879);
or U6918 (N_6918,N_6648,N_6653);
nand U6919 (N_6919,N_6651,N_6613);
xor U6920 (N_6920,N_6801,N_6852);
nand U6921 (N_6921,N_6631,N_6678);
xor U6922 (N_6922,N_6827,N_6818);
nand U6923 (N_6923,N_6699,N_6861);
nor U6924 (N_6924,N_6731,N_6877);
and U6925 (N_6925,N_6622,N_6790);
nand U6926 (N_6926,N_6673,N_6712);
and U6927 (N_6927,N_6643,N_6765);
or U6928 (N_6928,N_6873,N_6682);
nand U6929 (N_6929,N_6762,N_6871);
or U6930 (N_6930,N_6674,N_6751);
xnor U6931 (N_6931,N_6843,N_6761);
xnor U6932 (N_6932,N_6836,N_6784);
or U6933 (N_6933,N_6721,N_6778);
xor U6934 (N_6934,N_6766,N_6817);
and U6935 (N_6935,N_6806,N_6623);
xor U6936 (N_6936,N_6769,N_6884);
nor U6937 (N_6937,N_6758,N_6605);
and U6938 (N_6938,N_6846,N_6655);
nand U6939 (N_6939,N_6767,N_6857);
and U6940 (N_6940,N_6710,N_6747);
xor U6941 (N_6941,N_6882,N_6708);
or U6942 (N_6942,N_6860,N_6616);
or U6943 (N_6943,N_6844,N_6634);
or U6944 (N_6944,N_6689,N_6608);
nor U6945 (N_6945,N_6795,N_6880);
nand U6946 (N_6946,N_6890,N_6798);
xnor U6947 (N_6947,N_6828,N_6654);
nand U6948 (N_6948,N_6780,N_6870);
or U6949 (N_6949,N_6803,N_6811);
xnor U6950 (N_6950,N_6647,N_6681);
or U6951 (N_6951,N_6789,N_6845);
and U6952 (N_6952,N_6630,N_6786);
or U6953 (N_6953,N_6834,N_6740);
or U6954 (N_6954,N_6617,N_6723);
or U6955 (N_6955,N_6742,N_6864);
xor U6956 (N_6956,N_6722,N_6680);
nor U6957 (N_6957,N_6771,N_6842);
nor U6958 (N_6958,N_6602,N_6665);
nor U6959 (N_6959,N_6764,N_6727);
xnor U6960 (N_6960,N_6640,N_6619);
or U6961 (N_6961,N_6847,N_6695);
and U6962 (N_6962,N_6802,N_6604);
and U6963 (N_6963,N_6897,N_6744);
and U6964 (N_6964,N_6776,N_6683);
or U6965 (N_6965,N_6796,N_6787);
or U6966 (N_6966,N_6848,N_6614);
or U6967 (N_6967,N_6807,N_6813);
or U6968 (N_6968,N_6675,N_6704);
nand U6969 (N_6969,N_6753,N_6885);
xnor U6970 (N_6970,N_6756,N_6777);
or U6971 (N_6971,N_6821,N_6706);
nor U6972 (N_6972,N_6735,N_6607);
xor U6973 (N_6973,N_6649,N_6759);
nor U6974 (N_6974,N_6814,N_6692);
or U6975 (N_6975,N_6737,N_6646);
or U6976 (N_6976,N_6650,N_6738);
and U6977 (N_6977,N_6815,N_6830);
xnor U6978 (N_6978,N_6626,N_6615);
and U6979 (N_6979,N_6698,N_6863);
xnor U6980 (N_6980,N_6770,N_6601);
or U6981 (N_6981,N_6808,N_6791);
nor U6982 (N_6982,N_6660,N_6831);
xnor U6983 (N_6983,N_6755,N_6819);
or U6984 (N_6984,N_6833,N_6892);
or U6985 (N_6985,N_6750,N_6888);
nor U6986 (N_6986,N_6606,N_6866);
and U6987 (N_6987,N_6661,N_6868);
nor U6988 (N_6988,N_6886,N_6662);
nor U6989 (N_6989,N_6652,N_6748);
and U6990 (N_6990,N_6720,N_6693);
nor U6991 (N_6991,N_6734,N_6633);
and U6992 (N_6992,N_6671,N_6781);
or U6993 (N_6993,N_6656,N_6768);
or U6994 (N_6994,N_6881,N_6718);
and U6995 (N_6995,N_6687,N_6858);
nand U6996 (N_6996,N_6822,N_6659);
nand U6997 (N_6997,N_6797,N_6688);
nand U6998 (N_6998,N_6869,N_6672);
or U6999 (N_6999,N_6618,N_6637);
and U7000 (N_7000,N_6609,N_6730);
nor U7001 (N_7001,N_6707,N_6785);
xor U7002 (N_7002,N_6887,N_6794);
nand U7003 (N_7003,N_6728,N_6745);
and U7004 (N_7004,N_6703,N_6670);
nand U7005 (N_7005,N_6853,N_6895);
nor U7006 (N_7006,N_6896,N_6713);
nand U7007 (N_7007,N_6625,N_6835);
xor U7008 (N_7008,N_6724,N_6711);
nand U7009 (N_7009,N_6774,N_6641);
nand U7010 (N_7010,N_6829,N_6757);
xnor U7011 (N_7011,N_6841,N_6743);
nor U7012 (N_7012,N_6824,N_6603);
and U7013 (N_7013,N_6627,N_6719);
xnor U7014 (N_7014,N_6709,N_6705);
nand U7015 (N_7015,N_6600,N_6760);
or U7016 (N_7016,N_6899,N_6823);
nor U7017 (N_7017,N_6729,N_6717);
nand U7018 (N_7018,N_6668,N_6736);
or U7019 (N_7019,N_6891,N_6838);
nand U7020 (N_7020,N_6893,N_6859);
xnor U7021 (N_7021,N_6638,N_6792);
and U7022 (N_7022,N_6799,N_6676);
nor U7023 (N_7023,N_6694,N_6862);
xnor U7024 (N_7024,N_6629,N_6667);
or U7025 (N_7025,N_6642,N_6894);
xor U7026 (N_7026,N_6883,N_6804);
nor U7027 (N_7027,N_6733,N_6810);
nor U7028 (N_7028,N_6644,N_6669);
xor U7029 (N_7029,N_6690,N_6875);
nand U7030 (N_7030,N_6809,N_6826);
and U7031 (N_7031,N_6684,N_6800);
and U7032 (N_7032,N_6779,N_6666);
xnor U7033 (N_7033,N_6725,N_6763);
nor U7034 (N_7034,N_6867,N_6849);
nor U7035 (N_7035,N_6856,N_6726);
xor U7036 (N_7036,N_6714,N_6772);
nor U7037 (N_7037,N_6752,N_6620);
nor U7038 (N_7038,N_6685,N_6851);
and U7039 (N_7039,N_6739,N_6793);
or U7040 (N_7040,N_6889,N_6696);
nand U7041 (N_7041,N_6805,N_6632);
nor U7042 (N_7042,N_6621,N_6741);
nand U7043 (N_7043,N_6783,N_6788);
xor U7044 (N_7044,N_6664,N_6773);
nand U7045 (N_7045,N_6702,N_6832);
xor U7046 (N_7046,N_6715,N_6624);
nor U7047 (N_7047,N_6657,N_6820);
xor U7048 (N_7048,N_6839,N_6628);
nor U7049 (N_7049,N_6645,N_6782);
xnor U7050 (N_7050,N_6729,N_6752);
nand U7051 (N_7051,N_6768,N_6879);
xnor U7052 (N_7052,N_6839,N_6870);
or U7053 (N_7053,N_6704,N_6862);
and U7054 (N_7054,N_6790,N_6834);
and U7055 (N_7055,N_6853,N_6631);
nor U7056 (N_7056,N_6749,N_6830);
and U7057 (N_7057,N_6733,N_6618);
nand U7058 (N_7058,N_6627,N_6623);
nand U7059 (N_7059,N_6849,N_6627);
or U7060 (N_7060,N_6699,N_6637);
xor U7061 (N_7061,N_6740,N_6626);
nor U7062 (N_7062,N_6844,N_6715);
and U7063 (N_7063,N_6737,N_6728);
xor U7064 (N_7064,N_6659,N_6681);
nand U7065 (N_7065,N_6774,N_6703);
xnor U7066 (N_7066,N_6649,N_6658);
xnor U7067 (N_7067,N_6667,N_6797);
xnor U7068 (N_7068,N_6656,N_6879);
xor U7069 (N_7069,N_6657,N_6830);
xnor U7070 (N_7070,N_6783,N_6641);
nor U7071 (N_7071,N_6607,N_6793);
and U7072 (N_7072,N_6760,N_6832);
xor U7073 (N_7073,N_6720,N_6859);
nor U7074 (N_7074,N_6891,N_6894);
and U7075 (N_7075,N_6890,N_6804);
and U7076 (N_7076,N_6808,N_6613);
and U7077 (N_7077,N_6749,N_6621);
nor U7078 (N_7078,N_6868,N_6765);
nor U7079 (N_7079,N_6645,N_6826);
and U7080 (N_7080,N_6854,N_6824);
nor U7081 (N_7081,N_6629,N_6634);
or U7082 (N_7082,N_6758,N_6644);
xnor U7083 (N_7083,N_6695,N_6645);
nor U7084 (N_7084,N_6618,N_6604);
nand U7085 (N_7085,N_6883,N_6643);
nor U7086 (N_7086,N_6708,N_6686);
and U7087 (N_7087,N_6693,N_6853);
xnor U7088 (N_7088,N_6732,N_6775);
and U7089 (N_7089,N_6715,N_6761);
or U7090 (N_7090,N_6842,N_6714);
xnor U7091 (N_7091,N_6718,N_6814);
nor U7092 (N_7092,N_6862,N_6775);
and U7093 (N_7093,N_6897,N_6839);
nand U7094 (N_7094,N_6614,N_6743);
nand U7095 (N_7095,N_6676,N_6611);
and U7096 (N_7096,N_6876,N_6622);
nor U7097 (N_7097,N_6789,N_6679);
nor U7098 (N_7098,N_6868,N_6865);
or U7099 (N_7099,N_6644,N_6786);
and U7100 (N_7100,N_6761,N_6620);
xnor U7101 (N_7101,N_6781,N_6621);
xor U7102 (N_7102,N_6715,N_6855);
nor U7103 (N_7103,N_6635,N_6608);
and U7104 (N_7104,N_6688,N_6834);
nor U7105 (N_7105,N_6762,N_6834);
or U7106 (N_7106,N_6674,N_6681);
nand U7107 (N_7107,N_6890,N_6749);
nand U7108 (N_7108,N_6602,N_6899);
nand U7109 (N_7109,N_6611,N_6613);
xnor U7110 (N_7110,N_6844,N_6720);
nor U7111 (N_7111,N_6784,N_6787);
or U7112 (N_7112,N_6885,N_6805);
nor U7113 (N_7113,N_6677,N_6887);
nor U7114 (N_7114,N_6653,N_6808);
xnor U7115 (N_7115,N_6857,N_6628);
or U7116 (N_7116,N_6657,N_6643);
nand U7117 (N_7117,N_6892,N_6869);
xor U7118 (N_7118,N_6820,N_6647);
or U7119 (N_7119,N_6782,N_6773);
or U7120 (N_7120,N_6613,N_6678);
or U7121 (N_7121,N_6643,N_6607);
nand U7122 (N_7122,N_6714,N_6690);
and U7123 (N_7123,N_6724,N_6784);
nand U7124 (N_7124,N_6742,N_6867);
nand U7125 (N_7125,N_6640,N_6795);
or U7126 (N_7126,N_6833,N_6898);
and U7127 (N_7127,N_6763,N_6817);
xor U7128 (N_7128,N_6729,N_6817);
and U7129 (N_7129,N_6714,N_6631);
nand U7130 (N_7130,N_6730,N_6727);
nor U7131 (N_7131,N_6814,N_6633);
nor U7132 (N_7132,N_6807,N_6681);
nor U7133 (N_7133,N_6638,N_6657);
nor U7134 (N_7134,N_6812,N_6731);
nand U7135 (N_7135,N_6643,N_6706);
xnor U7136 (N_7136,N_6662,N_6796);
nand U7137 (N_7137,N_6742,N_6774);
xnor U7138 (N_7138,N_6832,N_6793);
and U7139 (N_7139,N_6684,N_6832);
and U7140 (N_7140,N_6857,N_6740);
or U7141 (N_7141,N_6674,N_6893);
or U7142 (N_7142,N_6894,N_6721);
nand U7143 (N_7143,N_6779,N_6799);
nor U7144 (N_7144,N_6632,N_6688);
xor U7145 (N_7145,N_6724,N_6742);
or U7146 (N_7146,N_6632,N_6861);
nand U7147 (N_7147,N_6732,N_6787);
or U7148 (N_7148,N_6684,N_6813);
nor U7149 (N_7149,N_6796,N_6746);
nand U7150 (N_7150,N_6791,N_6632);
xor U7151 (N_7151,N_6620,N_6648);
and U7152 (N_7152,N_6750,N_6625);
or U7153 (N_7153,N_6645,N_6690);
nand U7154 (N_7154,N_6609,N_6616);
or U7155 (N_7155,N_6810,N_6719);
xor U7156 (N_7156,N_6687,N_6874);
xnor U7157 (N_7157,N_6625,N_6731);
and U7158 (N_7158,N_6873,N_6846);
and U7159 (N_7159,N_6729,N_6618);
and U7160 (N_7160,N_6848,N_6738);
nand U7161 (N_7161,N_6812,N_6895);
xor U7162 (N_7162,N_6713,N_6852);
and U7163 (N_7163,N_6612,N_6782);
and U7164 (N_7164,N_6613,N_6851);
nand U7165 (N_7165,N_6741,N_6877);
xor U7166 (N_7166,N_6710,N_6780);
nor U7167 (N_7167,N_6691,N_6655);
nor U7168 (N_7168,N_6822,N_6887);
nand U7169 (N_7169,N_6725,N_6861);
xnor U7170 (N_7170,N_6756,N_6665);
nand U7171 (N_7171,N_6612,N_6817);
nand U7172 (N_7172,N_6860,N_6883);
nand U7173 (N_7173,N_6664,N_6682);
nor U7174 (N_7174,N_6702,N_6835);
nand U7175 (N_7175,N_6771,N_6735);
nor U7176 (N_7176,N_6790,N_6754);
or U7177 (N_7177,N_6643,N_6646);
nor U7178 (N_7178,N_6725,N_6752);
nand U7179 (N_7179,N_6649,N_6872);
or U7180 (N_7180,N_6717,N_6783);
xnor U7181 (N_7181,N_6742,N_6708);
and U7182 (N_7182,N_6612,N_6708);
xor U7183 (N_7183,N_6804,N_6727);
or U7184 (N_7184,N_6724,N_6612);
and U7185 (N_7185,N_6887,N_6771);
or U7186 (N_7186,N_6651,N_6665);
or U7187 (N_7187,N_6765,N_6798);
and U7188 (N_7188,N_6757,N_6628);
nor U7189 (N_7189,N_6803,N_6768);
nand U7190 (N_7190,N_6872,N_6650);
nor U7191 (N_7191,N_6604,N_6849);
or U7192 (N_7192,N_6717,N_6689);
and U7193 (N_7193,N_6867,N_6769);
xor U7194 (N_7194,N_6669,N_6640);
or U7195 (N_7195,N_6754,N_6628);
nand U7196 (N_7196,N_6691,N_6780);
or U7197 (N_7197,N_6622,N_6895);
nor U7198 (N_7198,N_6760,N_6752);
and U7199 (N_7199,N_6864,N_6679);
and U7200 (N_7200,N_6962,N_7113);
xor U7201 (N_7201,N_7043,N_7013);
xor U7202 (N_7202,N_6929,N_7006);
nand U7203 (N_7203,N_7162,N_7023);
or U7204 (N_7204,N_6999,N_7193);
or U7205 (N_7205,N_7117,N_7109);
xor U7206 (N_7206,N_6955,N_7041);
xnor U7207 (N_7207,N_7167,N_7081);
nand U7208 (N_7208,N_7087,N_6931);
xor U7209 (N_7209,N_6916,N_7010);
and U7210 (N_7210,N_7079,N_7085);
xnor U7211 (N_7211,N_7105,N_7021);
xor U7212 (N_7212,N_7172,N_6963);
nand U7213 (N_7213,N_6978,N_7042);
nand U7214 (N_7214,N_7178,N_7086);
and U7215 (N_7215,N_7082,N_6944);
nor U7216 (N_7216,N_6950,N_6924);
xnor U7217 (N_7217,N_6956,N_7030);
nor U7218 (N_7218,N_7099,N_6968);
or U7219 (N_7219,N_7094,N_6977);
nand U7220 (N_7220,N_6988,N_7019);
or U7221 (N_7221,N_7179,N_7139);
or U7222 (N_7222,N_7046,N_6943);
nor U7223 (N_7223,N_7029,N_7176);
nand U7224 (N_7224,N_7131,N_7054);
xor U7225 (N_7225,N_6948,N_7148);
and U7226 (N_7226,N_6938,N_7025);
and U7227 (N_7227,N_6935,N_7173);
xor U7228 (N_7228,N_7145,N_7050);
xor U7229 (N_7229,N_6930,N_7101);
and U7230 (N_7230,N_6995,N_7002);
xnor U7231 (N_7231,N_7038,N_6970);
or U7232 (N_7232,N_6985,N_7133);
nand U7233 (N_7233,N_6957,N_6980);
or U7234 (N_7234,N_7044,N_7191);
and U7235 (N_7235,N_7014,N_6966);
and U7236 (N_7236,N_7161,N_7115);
nand U7237 (N_7237,N_6920,N_7015);
nand U7238 (N_7238,N_6953,N_6902);
nor U7239 (N_7239,N_7022,N_7197);
or U7240 (N_7240,N_7152,N_7008);
or U7241 (N_7241,N_7166,N_6909);
nor U7242 (N_7242,N_6925,N_6933);
nand U7243 (N_7243,N_7140,N_6951);
xnor U7244 (N_7244,N_6994,N_7096);
and U7245 (N_7245,N_7088,N_6934);
and U7246 (N_7246,N_7111,N_7174);
or U7247 (N_7247,N_6997,N_6915);
nor U7248 (N_7248,N_6937,N_6984);
nand U7249 (N_7249,N_7104,N_7063);
and U7250 (N_7250,N_7159,N_7137);
xor U7251 (N_7251,N_7092,N_6958);
and U7252 (N_7252,N_6993,N_7070);
and U7253 (N_7253,N_7003,N_7129);
nor U7254 (N_7254,N_6964,N_7199);
nand U7255 (N_7255,N_7160,N_7141);
nand U7256 (N_7256,N_6965,N_7169);
nor U7257 (N_7257,N_7034,N_7151);
xor U7258 (N_7258,N_7000,N_7190);
and U7259 (N_7259,N_7058,N_6996);
or U7260 (N_7260,N_7168,N_7114);
or U7261 (N_7261,N_7187,N_7156);
xor U7262 (N_7262,N_6945,N_7112);
and U7263 (N_7263,N_7031,N_7138);
nand U7264 (N_7264,N_6961,N_7067);
and U7265 (N_7265,N_7163,N_7149);
xor U7266 (N_7266,N_6976,N_6912);
and U7267 (N_7267,N_7126,N_7007);
or U7268 (N_7268,N_7180,N_7055);
and U7269 (N_7269,N_6911,N_7078);
or U7270 (N_7270,N_7170,N_7072);
or U7271 (N_7271,N_7186,N_7011);
or U7272 (N_7272,N_6910,N_7116);
nor U7273 (N_7273,N_7153,N_7147);
or U7274 (N_7274,N_6982,N_7061);
xor U7275 (N_7275,N_6901,N_7090);
and U7276 (N_7276,N_6991,N_6960);
nor U7277 (N_7277,N_6983,N_6903);
or U7278 (N_7278,N_7069,N_7150);
nand U7279 (N_7279,N_7033,N_7047);
nor U7280 (N_7280,N_7028,N_7051);
xor U7281 (N_7281,N_7049,N_6959);
nor U7282 (N_7282,N_7056,N_6919);
nor U7283 (N_7283,N_7142,N_6967);
nand U7284 (N_7284,N_7017,N_7089);
nand U7285 (N_7285,N_6954,N_6987);
nor U7286 (N_7286,N_6986,N_7060);
xor U7287 (N_7287,N_7135,N_6975);
and U7288 (N_7288,N_7144,N_7183);
nand U7289 (N_7289,N_7040,N_7052);
nand U7290 (N_7290,N_7004,N_7074);
nand U7291 (N_7291,N_6947,N_7073);
and U7292 (N_7292,N_7084,N_7018);
and U7293 (N_7293,N_6941,N_6921);
or U7294 (N_7294,N_6990,N_7110);
nand U7295 (N_7295,N_6974,N_7185);
and U7296 (N_7296,N_6917,N_7122);
xnor U7297 (N_7297,N_6989,N_7128);
xor U7298 (N_7298,N_7076,N_6936);
or U7299 (N_7299,N_7005,N_6981);
and U7300 (N_7300,N_7102,N_7154);
xor U7301 (N_7301,N_6923,N_6949);
and U7302 (N_7302,N_7103,N_7016);
nor U7303 (N_7303,N_7136,N_7125);
nand U7304 (N_7304,N_6942,N_7035);
nor U7305 (N_7305,N_6998,N_7066);
or U7306 (N_7306,N_6927,N_7098);
xor U7307 (N_7307,N_6932,N_7188);
nand U7308 (N_7308,N_6946,N_7009);
nand U7309 (N_7309,N_6928,N_7196);
nor U7310 (N_7310,N_7107,N_7130);
or U7311 (N_7311,N_6969,N_7134);
nor U7312 (N_7312,N_7075,N_6971);
nor U7313 (N_7313,N_7012,N_7001);
xnor U7314 (N_7314,N_7192,N_7182);
or U7315 (N_7315,N_7146,N_7097);
or U7316 (N_7316,N_7143,N_7181);
xnor U7317 (N_7317,N_6922,N_7157);
xnor U7318 (N_7318,N_7175,N_7194);
xor U7319 (N_7319,N_7155,N_7080);
xnor U7320 (N_7320,N_7064,N_7048);
xnor U7321 (N_7321,N_7198,N_7039);
xor U7322 (N_7322,N_7164,N_6918);
nand U7323 (N_7323,N_6992,N_7093);
and U7324 (N_7324,N_7158,N_7068);
nor U7325 (N_7325,N_7124,N_6973);
xor U7326 (N_7326,N_7059,N_7108);
xnor U7327 (N_7327,N_7177,N_7127);
and U7328 (N_7328,N_6908,N_7077);
nand U7329 (N_7329,N_7106,N_7120);
nor U7330 (N_7330,N_7119,N_6906);
nor U7331 (N_7331,N_7095,N_6926);
nor U7332 (N_7332,N_7026,N_7032);
or U7333 (N_7333,N_7020,N_6907);
nand U7334 (N_7334,N_7189,N_6913);
and U7335 (N_7335,N_7071,N_7037);
or U7336 (N_7336,N_6979,N_7171);
xor U7337 (N_7337,N_7132,N_6900);
or U7338 (N_7338,N_7027,N_6972);
or U7339 (N_7339,N_7053,N_7091);
nor U7340 (N_7340,N_7065,N_6914);
or U7341 (N_7341,N_7184,N_7100);
xor U7342 (N_7342,N_6905,N_7118);
and U7343 (N_7343,N_6904,N_7083);
xor U7344 (N_7344,N_7045,N_7024);
or U7345 (N_7345,N_7036,N_7121);
xor U7346 (N_7346,N_7123,N_7062);
nor U7347 (N_7347,N_6939,N_7165);
or U7348 (N_7348,N_7195,N_7057);
or U7349 (N_7349,N_6952,N_6940);
xnor U7350 (N_7350,N_7032,N_7042);
nand U7351 (N_7351,N_7036,N_6997);
or U7352 (N_7352,N_7000,N_7161);
or U7353 (N_7353,N_7194,N_6971);
and U7354 (N_7354,N_7110,N_7040);
xor U7355 (N_7355,N_6931,N_7012);
nor U7356 (N_7356,N_6969,N_6954);
nand U7357 (N_7357,N_6987,N_7000);
nor U7358 (N_7358,N_6997,N_7012);
nand U7359 (N_7359,N_7038,N_6953);
or U7360 (N_7360,N_7100,N_7048);
and U7361 (N_7361,N_7157,N_7114);
xnor U7362 (N_7362,N_7170,N_6940);
nor U7363 (N_7363,N_7131,N_7169);
nor U7364 (N_7364,N_6924,N_7137);
nor U7365 (N_7365,N_7026,N_6955);
xor U7366 (N_7366,N_7169,N_7022);
nor U7367 (N_7367,N_6965,N_7080);
nand U7368 (N_7368,N_7017,N_7018);
or U7369 (N_7369,N_7068,N_7084);
and U7370 (N_7370,N_7044,N_7166);
and U7371 (N_7371,N_6986,N_7149);
nand U7372 (N_7372,N_6997,N_7072);
nand U7373 (N_7373,N_6963,N_7075);
and U7374 (N_7374,N_7162,N_7006);
nand U7375 (N_7375,N_7023,N_7152);
or U7376 (N_7376,N_7101,N_7043);
or U7377 (N_7377,N_7078,N_6900);
xor U7378 (N_7378,N_6963,N_7089);
or U7379 (N_7379,N_7171,N_7031);
xor U7380 (N_7380,N_6914,N_7101);
nand U7381 (N_7381,N_7155,N_7183);
or U7382 (N_7382,N_6962,N_6914);
xor U7383 (N_7383,N_6956,N_7162);
nor U7384 (N_7384,N_7039,N_7139);
and U7385 (N_7385,N_6962,N_7115);
or U7386 (N_7386,N_7140,N_7077);
and U7387 (N_7387,N_6962,N_6937);
and U7388 (N_7388,N_7156,N_7071);
nor U7389 (N_7389,N_7105,N_7002);
or U7390 (N_7390,N_7012,N_7192);
and U7391 (N_7391,N_7106,N_7160);
nand U7392 (N_7392,N_7124,N_7133);
or U7393 (N_7393,N_7077,N_6919);
nand U7394 (N_7394,N_6946,N_6929);
nand U7395 (N_7395,N_7166,N_7138);
nor U7396 (N_7396,N_6996,N_7071);
xor U7397 (N_7397,N_6970,N_7074);
or U7398 (N_7398,N_7083,N_7140);
xor U7399 (N_7399,N_7069,N_6901);
nor U7400 (N_7400,N_6953,N_6973);
and U7401 (N_7401,N_7164,N_7095);
xor U7402 (N_7402,N_7113,N_6985);
nand U7403 (N_7403,N_7159,N_7023);
nand U7404 (N_7404,N_6940,N_6927);
or U7405 (N_7405,N_7069,N_6930);
nand U7406 (N_7406,N_6959,N_6901);
xor U7407 (N_7407,N_7102,N_6967);
xor U7408 (N_7408,N_7086,N_6948);
or U7409 (N_7409,N_6946,N_7039);
xor U7410 (N_7410,N_7147,N_7181);
nor U7411 (N_7411,N_7161,N_7060);
xor U7412 (N_7412,N_7119,N_7189);
xnor U7413 (N_7413,N_7085,N_6923);
nand U7414 (N_7414,N_7000,N_7026);
and U7415 (N_7415,N_7033,N_6985);
nor U7416 (N_7416,N_6994,N_7119);
xnor U7417 (N_7417,N_7084,N_7064);
and U7418 (N_7418,N_7112,N_6920);
xnor U7419 (N_7419,N_7110,N_6923);
xnor U7420 (N_7420,N_7075,N_6948);
xnor U7421 (N_7421,N_7134,N_7049);
nor U7422 (N_7422,N_6989,N_6978);
nand U7423 (N_7423,N_7182,N_7046);
and U7424 (N_7424,N_7068,N_6931);
nand U7425 (N_7425,N_7066,N_7196);
and U7426 (N_7426,N_6962,N_6991);
nand U7427 (N_7427,N_6993,N_7141);
nand U7428 (N_7428,N_7052,N_7003);
and U7429 (N_7429,N_7032,N_7166);
nor U7430 (N_7430,N_7137,N_7115);
or U7431 (N_7431,N_7160,N_7190);
xnor U7432 (N_7432,N_7021,N_7166);
nand U7433 (N_7433,N_7122,N_6936);
nand U7434 (N_7434,N_7172,N_7058);
nor U7435 (N_7435,N_7111,N_7121);
and U7436 (N_7436,N_7061,N_6969);
and U7437 (N_7437,N_6906,N_7081);
xor U7438 (N_7438,N_7019,N_6986);
nor U7439 (N_7439,N_7195,N_7030);
nand U7440 (N_7440,N_6996,N_7118);
nand U7441 (N_7441,N_7138,N_6912);
nor U7442 (N_7442,N_7132,N_7088);
xnor U7443 (N_7443,N_7087,N_6990);
xor U7444 (N_7444,N_7198,N_6973);
and U7445 (N_7445,N_7013,N_6977);
xnor U7446 (N_7446,N_7166,N_7111);
and U7447 (N_7447,N_7075,N_7107);
xnor U7448 (N_7448,N_7113,N_7097);
nand U7449 (N_7449,N_7053,N_7138);
xor U7450 (N_7450,N_6926,N_7174);
xnor U7451 (N_7451,N_7036,N_7015);
nand U7452 (N_7452,N_6959,N_7082);
and U7453 (N_7453,N_7130,N_6972);
nand U7454 (N_7454,N_6993,N_7006);
and U7455 (N_7455,N_7049,N_7051);
and U7456 (N_7456,N_6931,N_7115);
xor U7457 (N_7457,N_7108,N_7109);
or U7458 (N_7458,N_7026,N_6960);
and U7459 (N_7459,N_7153,N_7036);
or U7460 (N_7460,N_7073,N_6922);
or U7461 (N_7461,N_6930,N_7118);
and U7462 (N_7462,N_7061,N_7050);
nand U7463 (N_7463,N_6950,N_6952);
nor U7464 (N_7464,N_7127,N_7123);
xnor U7465 (N_7465,N_6936,N_7064);
nor U7466 (N_7466,N_6940,N_7047);
nor U7467 (N_7467,N_6903,N_7057);
or U7468 (N_7468,N_7102,N_7184);
xnor U7469 (N_7469,N_7139,N_6994);
nor U7470 (N_7470,N_7060,N_6997);
xnor U7471 (N_7471,N_7083,N_6995);
or U7472 (N_7472,N_7045,N_6961);
or U7473 (N_7473,N_6992,N_7097);
or U7474 (N_7474,N_7168,N_6962);
nor U7475 (N_7475,N_7125,N_6976);
nand U7476 (N_7476,N_6945,N_7015);
nand U7477 (N_7477,N_6914,N_7001);
nor U7478 (N_7478,N_7016,N_6900);
xnor U7479 (N_7479,N_7003,N_7099);
or U7480 (N_7480,N_6915,N_6958);
nand U7481 (N_7481,N_7107,N_6950);
nand U7482 (N_7482,N_7109,N_6996);
or U7483 (N_7483,N_6921,N_7082);
nand U7484 (N_7484,N_7049,N_7080);
nand U7485 (N_7485,N_6944,N_7020);
nor U7486 (N_7486,N_7195,N_7052);
and U7487 (N_7487,N_7114,N_7099);
and U7488 (N_7488,N_7019,N_7023);
xor U7489 (N_7489,N_7027,N_6982);
nand U7490 (N_7490,N_7049,N_7014);
or U7491 (N_7491,N_6903,N_6924);
nand U7492 (N_7492,N_6930,N_7002);
xnor U7493 (N_7493,N_6962,N_7157);
or U7494 (N_7494,N_6958,N_7179);
nand U7495 (N_7495,N_6964,N_7174);
nor U7496 (N_7496,N_6938,N_7011);
or U7497 (N_7497,N_6941,N_7139);
nor U7498 (N_7498,N_7101,N_7185);
nor U7499 (N_7499,N_7196,N_7067);
or U7500 (N_7500,N_7236,N_7346);
nor U7501 (N_7501,N_7360,N_7244);
nand U7502 (N_7502,N_7427,N_7245);
nor U7503 (N_7503,N_7399,N_7242);
nand U7504 (N_7504,N_7309,N_7248);
and U7505 (N_7505,N_7293,N_7285);
xor U7506 (N_7506,N_7376,N_7214);
nand U7507 (N_7507,N_7365,N_7478);
or U7508 (N_7508,N_7370,N_7385);
or U7509 (N_7509,N_7257,N_7276);
and U7510 (N_7510,N_7382,N_7468);
and U7511 (N_7511,N_7284,N_7423);
nand U7512 (N_7512,N_7348,N_7436);
or U7513 (N_7513,N_7356,N_7444);
or U7514 (N_7514,N_7218,N_7233);
xnor U7515 (N_7515,N_7495,N_7331);
nand U7516 (N_7516,N_7221,N_7339);
nand U7517 (N_7517,N_7475,N_7234);
nor U7518 (N_7518,N_7440,N_7315);
or U7519 (N_7519,N_7393,N_7231);
nor U7520 (N_7520,N_7347,N_7390);
nor U7521 (N_7521,N_7483,N_7206);
nand U7522 (N_7522,N_7352,N_7232);
nor U7523 (N_7523,N_7251,N_7493);
or U7524 (N_7524,N_7490,N_7354);
or U7525 (N_7525,N_7380,N_7417);
and U7526 (N_7526,N_7419,N_7458);
and U7527 (N_7527,N_7292,N_7303);
or U7528 (N_7528,N_7268,N_7246);
and U7529 (N_7529,N_7326,N_7249);
xor U7530 (N_7530,N_7469,N_7396);
and U7531 (N_7531,N_7388,N_7443);
nor U7532 (N_7532,N_7484,N_7461);
nand U7533 (N_7533,N_7366,N_7256);
nand U7534 (N_7534,N_7486,N_7305);
or U7535 (N_7535,N_7448,N_7266);
or U7536 (N_7536,N_7404,N_7391);
nand U7537 (N_7537,N_7379,N_7273);
or U7538 (N_7538,N_7263,N_7405);
and U7539 (N_7539,N_7216,N_7464);
nor U7540 (N_7540,N_7397,N_7479);
nor U7541 (N_7541,N_7334,N_7219);
and U7542 (N_7542,N_7431,N_7491);
xor U7543 (N_7543,N_7407,N_7301);
nand U7544 (N_7544,N_7361,N_7375);
nand U7545 (N_7545,N_7480,N_7269);
or U7546 (N_7546,N_7314,N_7373);
and U7547 (N_7547,N_7445,N_7439);
nor U7548 (N_7548,N_7384,N_7368);
xnor U7549 (N_7549,N_7435,N_7333);
and U7550 (N_7550,N_7497,N_7243);
and U7551 (N_7551,N_7302,N_7306);
nand U7552 (N_7552,N_7310,N_7212);
xnor U7553 (N_7553,N_7330,N_7332);
and U7554 (N_7554,N_7317,N_7406);
nor U7555 (N_7555,N_7278,N_7204);
nand U7556 (N_7556,N_7449,N_7470);
or U7557 (N_7557,N_7386,N_7498);
nand U7558 (N_7558,N_7261,N_7222);
or U7559 (N_7559,N_7447,N_7424);
and U7560 (N_7560,N_7259,N_7327);
or U7561 (N_7561,N_7455,N_7372);
nand U7562 (N_7562,N_7316,N_7297);
xor U7563 (N_7563,N_7325,N_7336);
or U7564 (N_7564,N_7451,N_7320);
and U7565 (N_7565,N_7494,N_7477);
nand U7566 (N_7566,N_7254,N_7355);
nor U7567 (N_7567,N_7255,N_7217);
nor U7568 (N_7568,N_7398,N_7350);
nor U7569 (N_7569,N_7476,N_7446);
nor U7570 (N_7570,N_7296,N_7202);
nor U7571 (N_7571,N_7338,N_7323);
xor U7572 (N_7572,N_7413,N_7430);
nand U7573 (N_7573,N_7415,N_7462);
or U7574 (N_7574,N_7299,N_7262);
and U7575 (N_7575,N_7241,N_7342);
or U7576 (N_7576,N_7459,N_7279);
nor U7577 (N_7577,N_7329,N_7357);
xnor U7578 (N_7578,N_7207,N_7416);
nor U7579 (N_7579,N_7369,N_7265);
xor U7580 (N_7580,N_7275,N_7358);
nor U7581 (N_7581,N_7422,N_7453);
or U7582 (N_7582,N_7272,N_7438);
and U7583 (N_7583,N_7211,N_7496);
or U7584 (N_7584,N_7337,N_7465);
xor U7585 (N_7585,N_7240,N_7247);
or U7586 (N_7586,N_7313,N_7238);
nand U7587 (N_7587,N_7425,N_7281);
and U7588 (N_7588,N_7291,N_7230);
and U7589 (N_7589,N_7270,N_7203);
and U7590 (N_7590,N_7288,N_7377);
or U7591 (N_7591,N_7298,N_7304);
or U7592 (N_7592,N_7457,N_7400);
xor U7593 (N_7593,N_7414,N_7488);
or U7594 (N_7594,N_7201,N_7383);
or U7595 (N_7595,N_7412,N_7253);
and U7596 (N_7596,N_7467,N_7229);
or U7597 (N_7597,N_7353,N_7434);
nor U7598 (N_7598,N_7374,N_7437);
xnor U7599 (N_7599,N_7324,N_7289);
nand U7600 (N_7600,N_7274,N_7441);
or U7601 (N_7601,N_7466,N_7267);
and U7602 (N_7602,N_7228,N_7426);
or U7603 (N_7603,N_7286,N_7210);
nor U7604 (N_7604,N_7349,N_7271);
and U7605 (N_7605,N_7409,N_7220);
and U7606 (N_7606,N_7223,N_7307);
xor U7607 (N_7607,N_7237,N_7280);
nor U7608 (N_7608,N_7226,N_7472);
xor U7609 (N_7609,N_7321,N_7208);
and U7610 (N_7610,N_7225,N_7258);
xnor U7611 (N_7611,N_7344,N_7454);
xor U7612 (N_7612,N_7295,N_7308);
nand U7613 (N_7613,N_7312,N_7319);
or U7614 (N_7614,N_7362,N_7456);
xnor U7615 (N_7615,N_7387,N_7411);
nand U7616 (N_7616,N_7481,N_7489);
or U7617 (N_7617,N_7287,N_7487);
and U7618 (N_7618,N_7200,N_7290);
nand U7619 (N_7619,N_7335,N_7410);
and U7620 (N_7620,N_7460,N_7224);
nand U7621 (N_7621,N_7418,N_7239);
nand U7622 (N_7622,N_7215,N_7300);
nand U7623 (N_7623,N_7294,N_7378);
xor U7624 (N_7624,N_7205,N_7264);
and U7625 (N_7625,N_7442,N_7408);
xnor U7626 (N_7626,N_7252,N_7213);
and U7627 (N_7627,N_7474,N_7322);
or U7628 (N_7628,N_7394,N_7452);
and U7629 (N_7629,N_7359,N_7499);
and U7630 (N_7630,N_7471,N_7328);
nor U7631 (N_7631,N_7485,N_7429);
nand U7632 (N_7632,N_7363,N_7402);
and U7633 (N_7633,N_7463,N_7420);
or U7634 (N_7634,N_7318,N_7450);
xor U7635 (N_7635,N_7209,N_7364);
nor U7636 (N_7636,N_7227,N_7482);
nand U7637 (N_7637,N_7235,N_7282);
or U7638 (N_7638,N_7389,N_7395);
nand U7639 (N_7639,N_7351,N_7311);
nand U7640 (N_7640,N_7250,N_7381);
xor U7641 (N_7641,N_7392,N_7341);
xor U7642 (N_7642,N_7428,N_7260);
and U7643 (N_7643,N_7367,N_7343);
or U7644 (N_7644,N_7492,N_7277);
xor U7645 (N_7645,N_7403,N_7345);
nor U7646 (N_7646,N_7473,N_7433);
nand U7647 (N_7647,N_7401,N_7340);
nand U7648 (N_7648,N_7421,N_7432);
and U7649 (N_7649,N_7371,N_7283);
and U7650 (N_7650,N_7495,N_7389);
xnor U7651 (N_7651,N_7499,N_7217);
nand U7652 (N_7652,N_7212,N_7227);
xor U7653 (N_7653,N_7383,N_7387);
or U7654 (N_7654,N_7295,N_7490);
or U7655 (N_7655,N_7347,N_7428);
and U7656 (N_7656,N_7418,N_7208);
nand U7657 (N_7657,N_7242,N_7495);
and U7658 (N_7658,N_7350,N_7264);
xnor U7659 (N_7659,N_7308,N_7369);
xor U7660 (N_7660,N_7410,N_7290);
or U7661 (N_7661,N_7314,N_7385);
nand U7662 (N_7662,N_7335,N_7441);
nand U7663 (N_7663,N_7364,N_7287);
or U7664 (N_7664,N_7333,N_7441);
xnor U7665 (N_7665,N_7210,N_7491);
or U7666 (N_7666,N_7288,N_7413);
and U7667 (N_7667,N_7372,N_7404);
and U7668 (N_7668,N_7484,N_7436);
nand U7669 (N_7669,N_7443,N_7352);
nand U7670 (N_7670,N_7410,N_7392);
nor U7671 (N_7671,N_7264,N_7351);
and U7672 (N_7672,N_7450,N_7329);
or U7673 (N_7673,N_7360,N_7433);
and U7674 (N_7674,N_7353,N_7305);
nor U7675 (N_7675,N_7405,N_7425);
nor U7676 (N_7676,N_7420,N_7402);
or U7677 (N_7677,N_7292,N_7347);
nor U7678 (N_7678,N_7210,N_7216);
nand U7679 (N_7679,N_7460,N_7269);
xnor U7680 (N_7680,N_7381,N_7316);
and U7681 (N_7681,N_7380,N_7404);
xnor U7682 (N_7682,N_7475,N_7492);
nor U7683 (N_7683,N_7490,N_7324);
nor U7684 (N_7684,N_7306,N_7230);
nor U7685 (N_7685,N_7474,N_7355);
or U7686 (N_7686,N_7480,N_7431);
or U7687 (N_7687,N_7330,N_7277);
nand U7688 (N_7688,N_7415,N_7396);
nand U7689 (N_7689,N_7220,N_7432);
nor U7690 (N_7690,N_7343,N_7281);
or U7691 (N_7691,N_7334,N_7450);
nand U7692 (N_7692,N_7415,N_7372);
xnor U7693 (N_7693,N_7342,N_7213);
nor U7694 (N_7694,N_7452,N_7321);
and U7695 (N_7695,N_7368,N_7442);
and U7696 (N_7696,N_7437,N_7315);
and U7697 (N_7697,N_7427,N_7445);
nor U7698 (N_7698,N_7380,N_7472);
nand U7699 (N_7699,N_7330,N_7474);
or U7700 (N_7700,N_7489,N_7290);
xor U7701 (N_7701,N_7412,N_7352);
and U7702 (N_7702,N_7408,N_7204);
or U7703 (N_7703,N_7450,N_7315);
nand U7704 (N_7704,N_7469,N_7257);
nor U7705 (N_7705,N_7325,N_7492);
or U7706 (N_7706,N_7388,N_7299);
and U7707 (N_7707,N_7410,N_7201);
xnor U7708 (N_7708,N_7226,N_7468);
or U7709 (N_7709,N_7422,N_7406);
xor U7710 (N_7710,N_7405,N_7462);
xnor U7711 (N_7711,N_7256,N_7379);
and U7712 (N_7712,N_7347,N_7404);
and U7713 (N_7713,N_7372,N_7233);
nor U7714 (N_7714,N_7425,N_7292);
nor U7715 (N_7715,N_7459,N_7242);
and U7716 (N_7716,N_7254,N_7200);
xnor U7717 (N_7717,N_7427,N_7470);
or U7718 (N_7718,N_7346,N_7366);
xnor U7719 (N_7719,N_7427,N_7286);
xnor U7720 (N_7720,N_7491,N_7224);
or U7721 (N_7721,N_7266,N_7291);
xor U7722 (N_7722,N_7369,N_7458);
or U7723 (N_7723,N_7418,N_7431);
xnor U7724 (N_7724,N_7371,N_7248);
nand U7725 (N_7725,N_7436,N_7250);
or U7726 (N_7726,N_7249,N_7380);
and U7727 (N_7727,N_7254,N_7340);
xnor U7728 (N_7728,N_7471,N_7304);
nor U7729 (N_7729,N_7264,N_7289);
and U7730 (N_7730,N_7445,N_7217);
nor U7731 (N_7731,N_7416,N_7466);
nor U7732 (N_7732,N_7362,N_7259);
or U7733 (N_7733,N_7360,N_7435);
or U7734 (N_7734,N_7282,N_7418);
nand U7735 (N_7735,N_7338,N_7480);
nor U7736 (N_7736,N_7443,N_7334);
and U7737 (N_7737,N_7308,N_7422);
nand U7738 (N_7738,N_7399,N_7281);
nand U7739 (N_7739,N_7327,N_7422);
xnor U7740 (N_7740,N_7422,N_7466);
and U7741 (N_7741,N_7495,N_7237);
and U7742 (N_7742,N_7201,N_7488);
and U7743 (N_7743,N_7212,N_7362);
or U7744 (N_7744,N_7279,N_7353);
nor U7745 (N_7745,N_7378,N_7462);
xor U7746 (N_7746,N_7238,N_7321);
or U7747 (N_7747,N_7368,N_7374);
xnor U7748 (N_7748,N_7257,N_7348);
nor U7749 (N_7749,N_7240,N_7275);
nand U7750 (N_7750,N_7443,N_7367);
or U7751 (N_7751,N_7255,N_7437);
or U7752 (N_7752,N_7200,N_7238);
and U7753 (N_7753,N_7241,N_7487);
and U7754 (N_7754,N_7331,N_7238);
nand U7755 (N_7755,N_7449,N_7367);
and U7756 (N_7756,N_7222,N_7419);
nand U7757 (N_7757,N_7317,N_7215);
xor U7758 (N_7758,N_7474,N_7428);
or U7759 (N_7759,N_7273,N_7264);
xnor U7760 (N_7760,N_7404,N_7213);
nor U7761 (N_7761,N_7363,N_7224);
xnor U7762 (N_7762,N_7447,N_7327);
and U7763 (N_7763,N_7382,N_7232);
and U7764 (N_7764,N_7365,N_7352);
xnor U7765 (N_7765,N_7283,N_7333);
nand U7766 (N_7766,N_7442,N_7205);
nor U7767 (N_7767,N_7284,N_7353);
xor U7768 (N_7768,N_7331,N_7305);
xnor U7769 (N_7769,N_7407,N_7330);
xnor U7770 (N_7770,N_7453,N_7204);
and U7771 (N_7771,N_7437,N_7263);
nor U7772 (N_7772,N_7379,N_7344);
or U7773 (N_7773,N_7413,N_7464);
nor U7774 (N_7774,N_7316,N_7255);
or U7775 (N_7775,N_7334,N_7360);
and U7776 (N_7776,N_7273,N_7363);
nand U7777 (N_7777,N_7351,N_7425);
and U7778 (N_7778,N_7276,N_7443);
nand U7779 (N_7779,N_7447,N_7259);
nand U7780 (N_7780,N_7313,N_7372);
nor U7781 (N_7781,N_7303,N_7410);
nand U7782 (N_7782,N_7394,N_7418);
nand U7783 (N_7783,N_7394,N_7473);
and U7784 (N_7784,N_7206,N_7495);
nor U7785 (N_7785,N_7379,N_7442);
or U7786 (N_7786,N_7438,N_7347);
or U7787 (N_7787,N_7386,N_7340);
and U7788 (N_7788,N_7367,N_7254);
or U7789 (N_7789,N_7455,N_7407);
nand U7790 (N_7790,N_7207,N_7464);
nor U7791 (N_7791,N_7394,N_7378);
and U7792 (N_7792,N_7208,N_7289);
xor U7793 (N_7793,N_7299,N_7307);
nand U7794 (N_7794,N_7330,N_7254);
and U7795 (N_7795,N_7498,N_7345);
and U7796 (N_7796,N_7431,N_7305);
xnor U7797 (N_7797,N_7316,N_7246);
nand U7798 (N_7798,N_7446,N_7411);
and U7799 (N_7799,N_7437,N_7379);
nand U7800 (N_7800,N_7593,N_7762);
or U7801 (N_7801,N_7580,N_7642);
nor U7802 (N_7802,N_7616,N_7790);
or U7803 (N_7803,N_7624,N_7722);
nand U7804 (N_7804,N_7670,N_7599);
xor U7805 (N_7805,N_7797,N_7535);
and U7806 (N_7806,N_7667,N_7559);
nand U7807 (N_7807,N_7613,N_7777);
xnor U7808 (N_7808,N_7786,N_7774);
and U7809 (N_7809,N_7606,N_7765);
nor U7810 (N_7810,N_7779,N_7603);
and U7811 (N_7811,N_7677,N_7618);
xnor U7812 (N_7812,N_7770,N_7748);
and U7813 (N_7813,N_7671,N_7706);
or U7814 (N_7814,N_7731,N_7585);
xor U7815 (N_7815,N_7697,N_7761);
or U7816 (N_7816,N_7652,N_7569);
xnor U7817 (N_7817,N_7752,N_7699);
nand U7818 (N_7818,N_7653,N_7771);
and U7819 (N_7819,N_7750,N_7622);
nor U7820 (N_7820,N_7772,N_7525);
and U7821 (N_7821,N_7773,N_7620);
nand U7822 (N_7822,N_7510,N_7798);
and U7823 (N_7823,N_7675,N_7693);
nor U7824 (N_7824,N_7723,N_7742);
xnor U7825 (N_7825,N_7789,N_7720);
xor U7826 (N_7826,N_7565,N_7547);
xor U7827 (N_7827,N_7610,N_7778);
nand U7828 (N_7828,N_7702,N_7649);
nor U7829 (N_7829,N_7726,N_7733);
and U7830 (N_7830,N_7554,N_7645);
nand U7831 (N_7831,N_7621,N_7544);
or U7832 (N_7832,N_7792,N_7632);
xnor U7833 (N_7833,N_7586,N_7517);
nor U7834 (N_7834,N_7734,N_7740);
nand U7835 (N_7835,N_7515,N_7781);
nand U7836 (N_7836,N_7692,N_7721);
nor U7837 (N_7837,N_7615,N_7567);
nor U7838 (N_7838,N_7531,N_7636);
and U7839 (N_7839,N_7678,N_7719);
nand U7840 (N_7840,N_7540,N_7738);
nor U7841 (N_7841,N_7764,N_7795);
or U7842 (N_7842,N_7638,N_7766);
nor U7843 (N_7843,N_7573,N_7756);
xor U7844 (N_7844,N_7662,N_7572);
nand U7845 (N_7845,N_7658,N_7551);
or U7846 (N_7846,N_7711,N_7700);
nand U7847 (N_7847,N_7717,N_7509);
or U7848 (N_7848,N_7537,N_7614);
nand U7849 (N_7849,N_7579,N_7788);
nand U7850 (N_7850,N_7663,N_7555);
nor U7851 (N_7851,N_7617,N_7791);
nand U7852 (N_7852,N_7793,N_7557);
nor U7853 (N_7853,N_7688,N_7698);
and U7854 (N_7854,N_7524,N_7602);
and U7855 (N_7855,N_7628,N_7534);
nand U7856 (N_7856,N_7665,N_7705);
or U7857 (N_7857,N_7589,N_7631);
nor U7858 (N_7858,N_7528,N_7595);
or U7859 (N_7859,N_7527,N_7785);
nor U7860 (N_7860,N_7558,N_7657);
nand U7861 (N_7861,N_7577,N_7560);
nor U7862 (N_7862,N_7716,N_7685);
nor U7863 (N_7863,N_7594,N_7530);
nor U7864 (N_7864,N_7550,N_7584);
nand U7865 (N_7865,N_7647,N_7767);
nor U7866 (N_7866,N_7783,N_7598);
nor U7867 (N_7867,N_7536,N_7541);
or U7868 (N_7868,N_7533,N_7566);
and U7869 (N_7869,N_7591,N_7745);
nor U7870 (N_7870,N_7576,N_7582);
nand U7871 (N_7871,N_7501,N_7600);
and U7872 (N_7872,N_7590,N_7741);
or U7873 (N_7873,N_7597,N_7629);
and U7874 (N_7874,N_7763,N_7757);
or U7875 (N_7875,N_7609,N_7633);
nand U7876 (N_7876,N_7732,N_7523);
xor U7877 (N_7877,N_7648,N_7759);
and U7878 (N_7878,N_7561,N_7680);
nor U7879 (N_7879,N_7686,N_7506);
nor U7880 (N_7880,N_7782,N_7730);
nand U7881 (N_7881,N_7736,N_7562);
and U7882 (N_7882,N_7660,N_7707);
nor U7883 (N_7883,N_7511,N_7634);
xor U7884 (N_7884,N_7760,N_7724);
nand U7885 (N_7885,N_7701,N_7507);
or U7886 (N_7886,N_7502,N_7556);
and U7887 (N_7887,N_7529,N_7625);
and U7888 (N_7888,N_7753,N_7626);
and U7889 (N_7889,N_7521,N_7553);
nor U7890 (N_7890,N_7718,N_7713);
or U7891 (N_7891,N_7651,N_7635);
or U7892 (N_7892,N_7604,N_7708);
xnor U7893 (N_7893,N_7564,N_7520);
xor U7894 (N_7894,N_7640,N_7668);
nand U7895 (N_7895,N_7543,N_7681);
xor U7896 (N_7896,N_7674,N_7592);
nor U7897 (N_7897,N_7746,N_7780);
nand U7898 (N_7898,N_7644,N_7690);
and U7899 (N_7899,N_7650,N_7666);
nor U7900 (N_7900,N_7794,N_7545);
nor U7901 (N_7901,N_7776,N_7571);
xnor U7902 (N_7902,N_7601,N_7715);
xor U7903 (N_7903,N_7710,N_7695);
or U7904 (N_7904,N_7641,N_7575);
nand U7905 (N_7905,N_7587,N_7519);
nand U7906 (N_7906,N_7596,N_7784);
nor U7907 (N_7907,N_7608,N_7754);
and U7908 (N_7908,N_7751,N_7578);
xor U7909 (N_7909,N_7548,N_7643);
or U7910 (N_7910,N_7743,N_7691);
nor U7911 (N_7911,N_7522,N_7725);
nor U7912 (N_7912,N_7505,N_7612);
nor U7913 (N_7913,N_7539,N_7714);
nand U7914 (N_7914,N_7669,N_7549);
nor U7915 (N_7915,N_7664,N_7758);
and U7916 (N_7916,N_7694,N_7683);
xnor U7917 (N_7917,N_7611,N_7563);
nand U7918 (N_7918,N_7735,N_7696);
nor U7919 (N_7919,N_7588,N_7687);
xnor U7920 (N_7920,N_7682,N_7538);
or U7921 (N_7921,N_7775,N_7526);
nor U7922 (N_7922,N_7656,N_7583);
and U7923 (N_7923,N_7796,N_7676);
nor U7924 (N_7924,N_7542,N_7513);
nand U7925 (N_7925,N_7737,N_7503);
or U7926 (N_7926,N_7532,N_7574);
nor U7927 (N_7927,N_7768,N_7546);
xnor U7928 (N_7928,N_7727,N_7769);
nor U7929 (N_7929,N_7799,N_7581);
nor U7930 (N_7930,N_7755,N_7605);
or U7931 (N_7931,N_7747,N_7500);
xor U7932 (N_7932,N_7739,N_7508);
xnor U7933 (N_7933,N_7679,N_7654);
xor U7934 (N_7934,N_7646,N_7518);
and U7935 (N_7935,N_7637,N_7787);
nor U7936 (N_7936,N_7661,N_7516);
nand U7937 (N_7937,N_7689,N_7709);
xor U7938 (N_7938,N_7570,N_7512);
and U7939 (N_7939,N_7607,N_7639);
nor U7940 (N_7940,N_7655,N_7504);
and U7941 (N_7941,N_7749,N_7568);
or U7942 (N_7942,N_7619,N_7672);
or U7943 (N_7943,N_7729,N_7703);
or U7944 (N_7944,N_7630,N_7684);
nor U7945 (N_7945,N_7712,N_7552);
nor U7946 (N_7946,N_7514,N_7623);
nor U7947 (N_7947,N_7627,N_7728);
or U7948 (N_7948,N_7704,N_7659);
xor U7949 (N_7949,N_7673,N_7744);
and U7950 (N_7950,N_7780,N_7768);
or U7951 (N_7951,N_7598,N_7671);
or U7952 (N_7952,N_7558,N_7597);
or U7953 (N_7953,N_7758,N_7693);
nor U7954 (N_7954,N_7682,N_7546);
or U7955 (N_7955,N_7786,N_7602);
and U7956 (N_7956,N_7691,N_7756);
and U7957 (N_7957,N_7644,N_7700);
xor U7958 (N_7958,N_7714,N_7625);
nand U7959 (N_7959,N_7767,N_7702);
and U7960 (N_7960,N_7666,N_7607);
or U7961 (N_7961,N_7615,N_7724);
nor U7962 (N_7962,N_7514,N_7709);
xor U7963 (N_7963,N_7750,N_7752);
nand U7964 (N_7964,N_7561,N_7658);
xor U7965 (N_7965,N_7725,N_7745);
or U7966 (N_7966,N_7700,N_7572);
xor U7967 (N_7967,N_7569,N_7724);
or U7968 (N_7968,N_7655,N_7681);
and U7969 (N_7969,N_7593,N_7652);
and U7970 (N_7970,N_7584,N_7660);
or U7971 (N_7971,N_7592,N_7736);
and U7972 (N_7972,N_7575,N_7743);
nand U7973 (N_7973,N_7605,N_7577);
nor U7974 (N_7974,N_7621,N_7593);
nor U7975 (N_7975,N_7761,N_7602);
xor U7976 (N_7976,N_7510,N_7518);
xor U7977 (N_7977,N_7615,N_7534);
nand U7978 (N_7978,N_7625,N_7745);
nand U7979 (N_7979,N_7768,N_7757);
nand U7980 (N_7980,N_7591,N_7710);
xor U7981 (N_7981,N_7575,N_7748);
nor U7982 (N_7982,N_7680,N_7610);
nand U7983 (N_7983,N_7591,N_7505);
nor U7984 (N_7984,N_7793,N_7778);
nand U7985 (N_7985,N_7500,N_7586);
nand U7986 (N_7986,N_7724,N_7554);
xnor U7987 (N_7987,N_7618,N_7793);
nand U7988 (N_7988,N_7733,N_7613);
and U7989 (N_7989,N_7626,N_7527);
nor U7990 (N_7990,N_7787,N_7546);
nand U7991 (N_7991,N_7730,N_7544);
or U7992 (N_7992,N_7682,N_7643);
xnor U7993 (N_7993,N_7619,N_7723);
or U7994 (N_7994,N_7548,N_7714);
nor U7995 (N_7995,N_7532,N_7587);
nor U7996 (N_7996,N_7543,N_7702);
nand U7997 (N_7997,N_7582,N_7799);
or U7998 (N_7998,N_7764,N_7551);
nor U7999 (N_7999,N_7556,N_7788);
xor U8000 (N_8000,N_7583,N_7647);
or U8001 (N_8001,N_7712,N_7508);
xnor U8002 (N_8002,N_7672,N_7732);
nand U8003 (N_8003,N_7651,N_7576);
xnor U8004 (N_8004,N_7629,N_7647);
nor U8005 (N_8005,N_7505,N_7636);
and U8006 (N_8006,N_7650,N_7762);
or U8007 (N_8007,N_7634,N_7636);
nor U8008 (N_8008,N_7639,N_7594);
xor U8009 (N_8009,N_7793,N_7580);
or U8010 (N_8010,N_7798,N_7732);
nand U8011 (N_8011,N_7636,N_7641);
nor U8012 (N_8012,N_7664,N_7714);
nor U8013 (N_8013,N_7744,N_7536);
and U8014 (N_8014,N_7668,N_7709);
or U8015 (N_8015,N_7739,N_7571);
and U8016 (N_8016,N_7544,N_7798);
or U8017 (N_8017,N_7524,N_7552);
xor U8018 (N_8018,N_7719,N_7662);
or U8019 (N_8019,N_7718,N_7519);
xor U8020 (N_8020,N_7597,N_7533);
and U8021 (N_8021,N_7636,N_7573);
xor U8022 (N_8022,N_7568,N_7592);
xnor U8023 (N_8023,N_7515,N_7697);
nor U8024 (N_8024,N_7739,N_7592);
xor U8025 (N_8025,N_7743,N_7626);
xnor U8026 (N_8026,N_7763,N_7556);
and U8027 (N_8027,N_7605,N_7566);
nand U8028 (N_8028,N_7667,N_7555);
xnor U8029 (N_8029,N_7599,N_7549);
or U8030 (N_8030,N_7501,N_7508);
nor U8031 (N_8031,N_7534,N_7609);
nand U8032 (N_8032,N_7565,N_7652);
or U8033 (N_8033,N_7623,N_7657);
nand U8034 (N_8034,N_7594,N_7651);
nand U8035 (N_8035,N_7666,N_7536);
nand U8036 (N_8036,N_7752,N_7536);
nor U8037 (N_8037,N_7543,N_7713);
nand U8038 (N_8038,N_7793,N_7518);
nor U8039 (N_8039,N_7747,N_7640);
and U8040 (N_8040,N_7737,N_7666);
xnor U8041 (N_8041,N_7559,N_7510);
xor U8042 (N_8042,N_7750,N_7567);
and U8043 (N_8043,N_7774,N_7552);
nor U8044 (N_8044,N_7556,N_7728);
nand U8045 (N_8045,N_7607,N_7668);
nor U8046 (N_8046,N_7729,N_7659);
xnor U8047 (N_8047,N_7785,N_7598);
xnor U8048 (N_8048,N_7506,N_7540);
nand U8049 (N_8049,N_7572,N_7623);
or U8050 (N_8050,N_7772,N_7685);
nor U8051 (N_8051,N_7562,N_7522);
or U8052 (N_8052,N_7768,N_7787);
nand U8053 (N_8053,N_7613,N_7665);
and U8054 (N_8054,N_7650,N_7508);
or U8055 (N_8055,N_7714,N_7622);
nor U8056 (N_8056,N_7747,N_7505);
or U8057 (N_8057,N_7529,N_7556);
nor U8058 (N_8058,N_7544,N_7576);
nand U8059 (N_8059,N_7652,N_7661);
or U8060 (N_8060,N_7664,N_7580);
and U8061 (N_8061,N_7508,N_7600);
xnor U8062 (N_8062,N_7683,N_7748);
nor U8063 (N_8063,N_7604,N_7521);
nand U8064 (N_8064,N_7782,N_7793);
or U8065 (N_8065,N_7658,N_7742);
nor U8066 (N_8066,N_7633,N_7737);
or U8067 (N_8067,N_7641,N_7749);
nor U8068 (N_8068,N_7515,N_7514);
nor U8069 (N_8069,N_7717,N_7572);
nand U8070 (N_8070,N_7782,N_7598);
xor U8071 (N_8071,N_7701,N_7658);
and U8072 (N_8072,N_7773,N_7618);
or U8073 (N_8073,N_7797,N_7505);
and U8074 (N_8074,N_7772,N_7554);
nor U8075 (N_8075,N_7516,N_7726);
nand U8076 (N_8076,N_7692,N_7671);
or U8077 (N_8077,N_7788,N_7572);
nor U8078 (N_8078,N_7520,N_7753);
or U8079 (N_8079,N_7667,N_7687);
and U8080 (N_8080,N_7683,N_7681);
nand U8081 (N_8081,N_7779,N_7576);
nand U8082 (N_8082,N_7731,N_7532);
xnor U8083 (N_8083,N_7551,N_7545);
and U8084 (N_8084,N_7703,N_7604);
nand U8085 (N_8085,N_7754,N_7698);
and U8086 (N_8086,N_7552,N_7558);
and U8087 (N_8087,N_7614,N_7713);
nor U8088 (N_8088,N_7676,N_7530);
nor U8089 (N_8089,N_7788,N_7620);
nand U8090 (N_8090,N_7548,N_7585);
nor U8091 (N_8091,N_7789,N_7766);
and U8092 (N_8092,N_7653,N_7643);
xor U8093 (N_8093,N_7612,N_7689);
and U8094 (N_8094,N_7537,N_7758);
and U8095 (N_8095,N_7747,N_7658);
and U8096 (N_8096,N_7663,N_7550);
xor U8097 (N_8097,N_7756,N_7749);
and U8098 (N_8098,N_7784,N_7732);
xor U8099 (N_8099,N_7727,N_7542);
or U8100 (N_8100,N_7838,N_7813);
nor U8101 (N_8101,N_7962,N_7960);
nor U8102 (N_8102,N_7973,N_7819);
nor U8103 (N_8103,N_7829,N_7992);
xnor U8104 (N_8104,N_8067,N_7818);
nand U8105 (N_8105,N_7832,N_7821);
nor U8106 (N_8106,N_7948,N_7870);
and U8107 (N_8107,N_7814,N_8023);
xor U8108 (N_8108,N_7990,N_7892);
nor U8109 (N_8109,N_7862,N_7817);
nor U8110 (N_8110,N_8072,N_8074);
xnor U8111 (N_8111,N_8063,N_8020);
and U8112 (N_8112,N_7909,N_7911);
nor U8113 (N_8113,N_7884,N_7897);
or U8114 (N_8114,N_7834,N_7947);
xnor U8115 (N_8115,N_8098,N_7855);
nor U8116 (N_8116,N_7878,N_8053);
and U8117 (N_8117,N_8009,N_7859);
xor U8118 (N_8118,N_7972,N_7856);
and U8119 (N_8119,N_7954,N_7957);
nor U8120 (N_8120,N_8057,N_7865);
xor U8121 (N_8121,N_7995,N_7842);
xnor U8122 (N_8122,N_7847,N_7854);
and U8123 (N_8123,N_8078,N_7934);
nand U8124 (N_8124,N_7807,N_7905);
and U8125 (N_8125,N_7853,N_7946);
nor U8126 (N_8126,N_8019,N_7841);
or U8127 (N_8127,N_8000,N_8056);
xnor U8128 (N_8128,N_7949,N_7866);
and U8129 (N_8129,N_8016,N_8086);
and U8130 (N_8130,N_8005,N_8007);
nor U8131 (N_8131,N_7888,N_7997);
nand U8132 (N_8132,N_7966,N_8047);
and U8133 (N_8133,N_7978,N_7925);
nor U8134 (N_8134,N_7915,N_7881);
and U8135 (N_8135,N_7858,N_7981);
nand U8136 (N_8136,N_7820,N_8075);
or U8137 (N_8137,N_8064,N_7950);
nor U8138 (N_8138,N_8002,N_8094);
nor U8139 (N_8139,N_7874,N_7920);
or U8140 (N_8140,N_7969,N_8024);
nand U8141 (N_8141,N_7898,N_8071);
nand U8142 (N_8142,N_7805,N_8046);
nor U8143 (N_8143,N_8093,N_7851);
xor U8144 (N_8144,N_8076,N_8012);
xor U8145 (N_8145,N_7823,N_8058);
nand U8146 (N_8146,N_8082,N_7882);
nor U8147 (N_8147,N_8040,N_8022);
and U8148 (N_8148,N_7968,N_7837);
xor U8149 (N_8149,N_7991,N_7809);
nand U8150 (N_8150,N_7886,N_7956);
nand U8151 (N_8151,N_7937,N_7986);
or U8152 (N_8152,N_7875,N_7891);
nor U8153 (N_8153,N_7831,N_7951);
nor U8154 (N_8154,N_8079,N_7811);
or U8155 (N_8155,N_7923,N_8014);
or U8156 (N_8156,N_7952,N_7993);
xor U8157 (N_8157,N_7926,N_7974);
nor U8158 (N_8158,N_7955,N_8025);
and U8159 (N_8159,N_8003,N_7835);
and U8160 (N_8160,N_7980,N_7977);
and U8161 (N_8161,N_7877,N_7945);
nor U8162 (N_8162,N_7979,N_7996);
nor U8163 (N_8163,N_8081,N_7907);
nand U8164 (N_8164,N_7861,N_8089);
nor U8165 (N_8165,N_7885,N_7876);
xnor U8166 (N_8166,N_7903,N_8080);
and U8167 (N_8167,N_8044,N_7822);
nand U8168 (N_8168,N_7836,N_7916);
nand U8169 (N_8169,N_7815,N_8090);
or U8170 (N_8170,N_8055,N_7840);
and U8171 (N_8171,N_7827,N_7963);
nand U8172 (N_8172,N_7887,N_8029);
nor U8173 (N_8173,N_8097,N_8099);
or U8174 (N_8174,N_7816,N_7967);
xor U8175 (N_8175,N_7924,N_8087);
and U8176 (N_8176,N_8095,N_7850);
nor U8177 (N_8177,N_8039,N_7958);
or U8178 (N_8178,N_7932,N_7918);
nand U8179 (N_8179,N_8049,N_7806);
and U8180 (N_8180,N_8018,N_8054);
nand U8181 (N_8181,N_7879,N_7944);
or U8182 (N_8182,N_7860,N_8037);
and U8183 (N_8183,N_7998,N_8021);
or U8184 (N_8184,N_7825,N_7913);
xor U8185 (N_8185,N_7988,N_7894);
or U8186 (N_8186,N_8048,N_8062);
and U8187 (N_8187,N_7953,N_7872);
or U8188 (N_8188,N_7919,N_8034);
nand U8189 (N_8189,N_7873,N_7930);
or U8190 (N_8190,N_8041,N_7843);
nand U8191 (N_8191,N_8008,N_8038);
and U8192 (N_8192,N_7961,N_8070);
and U8193 (N_8193,N_7889,N_7801);
and U8194 (N_8194,N_8083,N_7984);
nor U8195 (N_8195,N_8011,N_7939);
xor U8196 (N_8196,N_7824,N_8065);
or U8197 (N_8197,N_7857,N_7910);
xnor U8198 (N_8198,N_7931,N_7959);
and U8199 (N_8199,N_7846,N_8092);
or U8200 (N_8200,N_7810,N_7871);
and U8201 (N_8201,N_7936,N_8059);
xor U8202 (N_8202,N_8042,N_7985);
nand U8203 (N_8203,N_8096,N_8085);
and U8204 (N_8204,N_7994,N_7971);
or U8205 (N_8205,N_7864,N_7845);
xnor U8206 (N_8206,N_8077,N_7804);
and U8207 (N_8207,N_7928,N_7942);
xor U8208 (N_8208,N_7901,N_7868);
or U8209 (N_8209,N_7800,N_7808);
or U8210 (N_8210,N_7975,N_8060);
xnor U8211 (N_8211,N_8032,N_8061);
or U8212 (N_8212,N_8017,N_7965);
nor U8213 (N_8213,N_7830,N_8051);
nor U8214 (N_8214,N_8006,N_8073);
nand U8215 (N_8215,N_7906,N_7989);
nand U8216 (N_8216,N_8052,N_7929);
nand U8217 (N_8217,N_8069,N_7983);
nor U8218 (N_8218,N_7812,N_7839);
nand U8219 (N_8219,N_8036,N_7912);
or U8220 (N_8220,N_7863,N_7848);
or U8221 (N_8221,N_8091,N_7922);
nand U8222 (N_8222,N_7902,N_7849);
or U8223 (N_8223,N_8033,N_7833);
xnor U8224 (N_8224,N_8027,N_7883);
nand U8225 (N_8225,N_8013,N_7943);
or U8226 (N_8226,N_8088,N_7896);
and U8227 (N_8227,N_7921,N_7899);
and U8228 (N_8228,N_7938,N_7927);
xnor U8229 (N_8229,N_7982,N_8010);
xor U8230 (N_8230,N_7895,N_7900);
nand U8231 (N_8231,N_7867,N_7852);
xnor U8232 (N_8232,N_7826,N_8028);
nand U8233 (N_8233,N_7869,N_7917);
xnor U8234 (N_8234,N_8030,N_7970);
nor U8235 (N_8235,N_7880,N_7802);
nor U8236 (N_8236,N_7940,N_8031);
nand U8237 (N_8237,N_8050,N_7890);
and U8238 (N_8238,N_7844,N_7904);
nor U8239 (N_8239,N_7914,N_8066);
nand U8240 (N_8240,N_8001,N_7828);
xor U8241 (N_8241,N_8004,N_8015);
nand U8242 (N_8242,N_7941,N_7908);
nor U8243 (N_8243,N_8043,N_7987);
or U8244 (N_8244,N_7964,N_7976);
nor U8245 (N_8245,N_7893,N_7803);
nand U8246 (N_8246,N_7933,N_7999);
or U8247 (N_8247,N_8084,N_7935);
nand U8248 (N_8248,N_8035,N_8068);
nand U8249 (N_8249,N_8045,N_8026);
or U8250 (N_8250,N_7847,N_8087);
nand U8251 (N_8251,N_8064,N_7907);
xnor U8252 (N_8252,N_7941,N_7911);
xor U8253 (N_8253,N_7808,N_7855);
nand U8254 (N_8254,N_7939,N_7918);
xnor U8255 (N_8255,N_7916,N_7936);
or U8256 (N_8256,N_7929,N_7804);
or U8257 (N_8257,N_8020,N_7943);
or U8258 (N_8258,N_7917,N_7857);
or U8259 (N_8259,N_7806,N_7887);
xor U8260 (N_8260,N_7901,N_8086);
or U8261 (N_8261,N_7965,N_8090);
nand U8262 (N_8262,N_8002,N_7822);
xor U8263 (N_8263,N_7836,N_7911);
and U8264 (N_8264,N_7989,N_7974);
and U8265 (N_8265,N_7970,N_7942);
and U8266 (N_8266,N_8028,N_8079);
and U8267 (N_8267,N_7898,N_7970);
nor U8268 (N_8268,N_7941,N_7800);
or U8269 (N_8269,N_8046,N_7944);
nor U8270 (N_8270,N_7982,N_7918);
or U8271 (N_8271,N_8012,N_7970);
nor U8272 (N_8272,N_8078,N_8004);
nor U8273 (N_8273,N_7970,N_7805);
or U8274 (N_8274,N_7944,N_7881);
and U8275 (N_8275,N_7990,N_7823);
xor U8276 (N_8276,N_7869,N_7876);
and U8277 (N_8277,N_7975,N_8028);
nor U8278 (N_8278,N_7867,N_7912);
nor U8279 (N_8279,N_7879,N_8047);
nand U8280 (N_8280,N_7995,N_7979);
or U8281 (N_8281,N_7832,N_7825);
or U8282 (N_8282,N_7914,N_8045);
and U8283 (N_8283,N_8012,N_7852);
nor U8284 (N_8284,N_7968,N_8073);
or U8285 (N_8285,N_7989,N_7851);
or U8286 (N_8286,N_7917,N_7934);
or U8287 (N_8287,N_7879,N_7913);
nor U8288 (N_8288,N_7958,N_7836);
or U8289 (N_8289,N_7926,N_7803);
or U8290 (N_8290,N_8004,N_8095);
and U8291 (N_8291,N_7873,N_8090);
or U8292 (N_8292,N_7852,N_7887);
nor U8293 (N_8293,N_7808,N_7858);
nand U8294 (N_8294,N_7908,N_7929);
and U8295 (N_8295,N_8004,N_7942);
xnor U8296 (N_8296,N_7954,N_7830);
nand U8297 (N_8297,N_7890,N_7825);
nand U8298 (N_8298,N_8036,N_7864);
or U8299 (N_8299,N_7920,N_7857);
and U8300 (N_8300,N_8086,N_8090);
xnor U8301 (N_8301,N_7847,N_7899);
xor U8302 (N_8302,N_7973,N_7956);
xor U8303 (N_8303,N_7981,N_8057);
xor U8304 (N_8304,N_8091,N_8078);
xnor U8305 (N_8305,N_8090,N_8007);
nand U8306 (N_8306,N_7974,N_7961);
xnor U8307 (N_8307,N_7972,N_7947);
xnor U8308 (N_8308,N_7850,N_7921);
or U8309 (N_8309,N_7876,N_8094);
and U8310 (N_8310,N_7953,N_8036);
xor U8311 (N_8311,N_8051,N_8027);
nor U8312 (N_8312,N_8031,N_7853);
nand U8313 (N_8313,N_7809,N_8033);
nor U8314 (N_8314,N_7956,N_8065);
and U8315 (N_8315,N_8088,N_7999);
or U8316 (N_8316,N_7922,N_7923);
nor U8317 (N_8317,N_8007,N_8066);
and U8318 (N_8318,N_8025,N_7828);
and U8319 (N_8319,N_8030,N_8054);
nor U8320 (N_8320,N_7859,N_8061);
and U8321 (N_8321,N_7958,N_7987);
or U8322 (N_8322,N_8019,N_8080);
xnor U8323 (N_8323,N_8010,N_7846);
xor U8324 (N_8324,N_7978,N_7872);
nand U8325 (N_8325,N_7882,N_7893);
and U8326 (N_8326,N_7996,N_7891);
or U8327 (N_8327,N_8078,N_8064);
nand U8328 (N_8328,N_7891,N_7988);
xnor U8329 (N_8329,N_8000,N_8064);
xor U8330 (N_8330,N_8040,N_8085);
xnor U8331 (N_8331,N_7846,N_7905);
or U8332 (N_8332,N_7859,N_7901);
xor U8333 (N_8333,N_8056,N_8041);
or U8334 (N_8334,N_7950,N_7840);
nand U8335 (N_8335,N_8076,N_7965);
xnor U8336 (N_8336,N_7999,N_7855);
nand U8337 (N_8337,N_7816,N_8071);
and U8338 (N_8338,N_8085,N_7988);
and U8339 (N_8339,N_7814,N_7988);
or U8340 (N_8340,N_7881,N_8053);
xnor U8341 (N_8341,N_7860,N_8007);
nor U8342 (N_8342,N_8036,N_7965);
nand U8343 (N_8343,N_7845,N_8091);
nor U8344 (N_8344,N_7825,N_7812);
xnor U8345 (N_8345,N_7857,N_7976);
xor U8346 (N_8346,N_7924,N_7882);
or U8347 (N_8347,N_8087,N_7904);
or U8348 (N_8348,N_7950,N_7801);
or U8349 (N_8349,N_7916,N_7815);
xor U8350 (N_8350,N_7878,N_7914);
and U8351 (N_8351,N_7930,N_7917);
nor U8352 (N_8352,N_7858,N_7861);
xor U8353 (N_8353,N_7884,N_7994);
nor U8354 (N_8354,N_7950,N_7975);
nor U8355 (N_8355,N_7805,N_8081);
nand U8356 (N_8356,N_8000,N_7919);
or U8357 (N_8357,N_8083,N_7928);
nor U8358 (N_8358,N_7952,N_7860);
xnor U8359 (N_8359,N_8008,N_7956);
or U8360 (N_8360,N_8070,N_8095);
or U8361 (N_8361,N_7963,N_7867);
or U8362 (N_8362,N_7840,N_7841);
nand U8363 (N_8363,N_7996,N_7845);
nand U8364 (N_8364,N_8089,N_7834);
or U8365 (N_8365,N_7842,N_8061);
nor U8366 (N_8366,N_7933,N_8099);
or U8367 (N_8367,N_7987,N_7863);
or U8368 (N_8368,N_7927,N_7895);
or U8369 (N_8369,N_7943,N_8003);
nor U8370 (N_8370,N_7827,N_7838);
nor U8371 (N_8371,N_7931,N_8023);
and U8372 (N_8372,N_7843,N_8075);
xnor U8373 (N_8373,N_7896,N_8064);
and U8374 (N_8374,N_8068,N_7992);
nor U8375 (N_8375,N_8010,N_7934);
nand U8376 (N_8376,N_7904,N_8072);
nand U8377 (N_8377,N_7882,N_7985);
nor U8378 (N_8378,N_7971,N_7830);
and U8379 (N_8379,N_7998,N_8043);
xnor U8380 (N_8380,N_8027,N_7860);
xor U8381 (N_8381,N_7805,N_7827);
nor U8382 (N_8382,N_7865,N_7880);
and U8383 (N_8383,N_8071,N_8027);
xnor U8384 (N_8384,N_8059,N_7960);
xor U8385 (N_8385,N_8018,N_8091);
and U8386 (N_8386,N_8021,N_7911);
and U8387 (N_8387,N_7955,N_7991);
or U8388 (N_8388,N_8018,N_7842);
or U8389 (N_8389,N_7896,N_7858);
and U8390 (N_8390,N_7821,N_8098);
nor U8391 (N_8391,N_7979,N_7814);
xnor U8392 (N_8392,N_7895,N_8036);
and U8393 (N_8393,N_7900,N_8078);
xnor U8394 (N_8394,N_7928,N_8053);
nand U8395 (N_8395,N_7958,N_7839);
and U8396 (N_8396,N_8053,N_8081);
or U8397 (N_8397,N_7990,N_8000);
xor U8398 (N_8398,N_8076,N_7954);
nor U8399 (N_8399,N_8031,N_7985);
xor U8400 (N_8400,N_8364,N_8383);
xor U8401 (N_8401,N_8256,N_8189);
and U8402 (N_8402,N_8353,N_8248);
nand U8403 (N_8403,N_8314,N_8266);
or U8404 (N_8404,N_8111,N_8394);
xor U8405 (N_8405,N_8182,N_8140);
nand U8406 (N_8406,N_8113,N_8347);
nor U8407 (N_8407,N_8270,N_8144);
and U8408 (N_8408,N_8183,N_8222);
nand U8409 (N_8409,N_8318,N_8294);
nand U8410 (N_8410,N_8213,N_8168);
xnor U8411 (N_8411,N_8199,N_8355);
nand U8412 (N_8412,N_8231,N_8336);
or U8413 (N_8413,N_8103,N_8350);
or U8414 (N_8414,N_8267,N_8203);
and U8415 (N_8415,N_8263,N_8186);
or U8416 (N_8416,N_8329,N_8250);
or U8417 (N_8417,N_8181,N_8292);
xnor U8418 (N_8418,N_8370,N_8133);
or U8419 (N_8419,N_8385,N_8138);
xor U8420 (N_8420,N_8377,N_8200);
nor U8421 (N_8421,N_8220,N_8191);
nand U8422 (N_8422,N_8110,N_8163);
or U8423 (N_8423,N_8348,N_8324);
and U8424 (N_8424,N_8239,N_8255);
xnor U8425 (N_8425,N_8384,N_8160);
and U8426 (N_8426,N_8262,N_8376);
xnor U8427 (N_8427,N_8300,N_8321);
or U8428 (N_8428,N_8169,N_8346);
nor U8429 (N_8429,N_8121,N_8178);
nor U8430 (N_8430,N_8349,N_8315);
or U8431 (N_8431,N_8386,N_8293);
xnor U8432 (N_8432,N_8141,N_8257);
nor U8433 (N_8433,N_8284,N_8332);
nor U8434 (N_8434,N_8151,N_8225);
xor U8435 (N_8435,N_8130,N_8221);
or U8436 (N_8436,N_8393,N_8149);
nand U8437 (N_8437,N_8108,N_8165);
xnor U8438 (N_8438,N_8193,N_8340);
nor U8439 (N_8439,N_8125,N_8287);
and U8440 (N_8440,N_8190,N_8396);
nor U8441 (N_8441,N_8148,N_8312);
and U8442 (N_8442,N_8127,N_8338);
nor U8443 (N_8443,N_8155,N_8143);
nand U8444 (N_8444,N_8304,N_8253);
and U8445 (N_8445,N_8275,N_8245);
nand U8446 (N_8446,N_8123,N_8279);
nor U8447 (N_8447,N_8299,N_8237);
and U8448 (N_8448,N_8156,N_8274);
xor U8449 (N_8449,N_8295,N_8378);
xnor U8450 (N_8450,N_8136,N_8387);
or U8451 (N_8451,N_8362,N_8214);
and U8452 (N_8452,N_8351,N_8205);
or U8453 (N_8453,N_8322,N_8271);
or U8454 (N_8454,N_8210,N_8335);
xnor U8455 (N_8455,N_8184,N_8195);
nand U8456 (N_8456,N_8217,N_8337);
or U8457 (N_8457,N_8341,N_8211);
nor U8458 (N_8458,N_8372,N_8235);
or U8459 (N_8459,N_8283,N_8281);
nand U8460 (N_8460,N_8249,N_8319);
and U8461 (N_8461,N_8202,N_8244);
and U8462 (N_8462,N_8154,N_8260);
and U8463 (N_8463,N_8258,N_8309);
xnor U8464 (N_8464,N_8219,N_8166);
nand U8465 (N_8465,N_8259,N_8180);
nor U8466 (N_8466,N_8152,N_8146);
or U8467 (N_8467,N_8242,N_8176);
and U8468 (N_8468,N_8280,N_8101);
and U8469 (N_8469,N_8162,N_8288);
nand U8470 (N_8470,N_8192,N_8323);
or U8471 (N_8471,N_8331,N_8252);
or U8472 (N_8472,N_8261,N_8230);
and U8473 (N_8473,N_8187,N_8109);
nand U8474 (N_8474,N_8236,N_8356);
xnor U8475 (N_8475,N_8398,N_8254);
nor U8476 (N_8476,N_8296,N_8273);
nor U8477 (N_8477,N_8358,N_8159);
and U8478 (N_8478,N_8354,N_8172);
nand U8479 (N_8479,N_8373,N_8291);
or U8480 (N_8480,N_8313,N_8161);
xor U8481 (N_8481,N_8269,N_8171);
nand U8482 (N_8482,N_8104,N_8158);
nand U8483 (N_8483,N_8302,N_8390);
nor U8484 (N_8484,N_8212,N_8164);
nor U8485 (N_8485,N_8366,N_8129);
xnor U8486 (N_8486,N_8115,N_8363);
nand U8487 (N_8487,N_8301,N_8157);
or U8488 (N_8488,N_8174,N_8114);
xor U8489 (N_8489,N_8228,N_8328);
nand U8490 (N_8490,N_8188,N_8179);
and U8491 (N_8491,N_8264,N_8122);
nor U8492 (N_8492,N_8311,N_8352);
or U8493 (N_8493,N_8277,N_8128);
xnor U8494 (N_8494,N_8117,N_8360);
or U8495 (N_8495,N_8126,N_8102);
and U8496 (N_8496,N_8381,N_8310);
nand U8497 (N_8497,N_8147,N_8170);
xnor U8498 (N_8498,N_8142,N_8241);
nor U8499 (N_8499,N_8204,N_8265);
xnor U8500 (N_8500,N_8326,N_8391);
xnor U8501 (N_8501,N_8333,N_8112);
and U8502 (N_8502,N_8345,N_8361);
and U8503 (N_8503,N_8175,N_8368);
or U8504 (N_8504,N_8224,N_8196);
xor U8505 (N_8505,N_8298,N_8238);
nand U8506 (N_8506,N_8290,N_8107);
xor U8507 (N_8507,N_8388,N_8397);
or U8508 (N_8508,N_8207,N_8272);
and U8509 (N_8509,N_8375,N_8106);
nand U8510 (N_8510,N_8206,N_8227);
nor U8511 (N_8511,N_8197,N_8139);
and U8512 (N_8512,N_8289,N_8276);
and U8513 (N_8513,N_8240,N_8137);
nand U8514 (N_8514,N_8100,N_8208);
xor U8515 (N_8515,N_8215,N_8177);
nor U8516 (N_8516,N_8359,N_8119);
nor U8517 (N_8517,N_8307,N_8120);
nor U8518 (N_8518,N_8167,N_8216);
xor U8519 (N_8519,N_8232,N_8374);
nand U8520 (N_8520,N_8369,N_8342);
or U8521 (N_8521,N_8395,N_8367);
nand U8522 (N_8522,N_8153,N_8135);
xnor U8523 (N_8523,N_8389,N_8124);
or U8524 (N_8524,N_8131,N_8382);
nor U8525 (N_8525,N_8218,N_8282);
and U8526 (N_8526,N_8223,N_8251);
nand U8527 (N_8527,N_8132,N_8306);
nand U8528 (N_8528,N_8286,N_8343);
nor U8529 (N_8529,N_8233,N_8234);
or U8530 (N_8530,N_8134,N_8379);
and U8531 (N_8531,N_8371,N_8198);
or U8532 (N_8532,N_8330,N_8194);
nor U8533 (N_8533,N_8317,N_8303);
nand U8534 (N_8534,N_8334,N_8268);
xnor U8535 (N_8535,N_8380,N_8316);
or U8536 (N_8536,N_8392,N_8209);
nor U8537 (N_8537,N_8344,N_8226);
nor U8538 (N_8538,N_8246,N_8308);
nand U8539 (N_8539,N_8145,N_8185);
and U8540 (N_8540,N_8297,N_8339);
or U8541 (N_8541,N_8105,N_8116);
and U8542 (N_8542,N_8118,N_8243);
nor U8543 (N_8543,N_8173,N_8247);
and U8544 (N_8544,N_8278,N_8365);
nand U8545 (N_8545,N_8305,N_8150);
or U8546 (N_8546,N_8357,N_8399);
nand U8547 (N_8547,N_8320,N_8325);
xnor U8548 (N_8548,N_8285,N_8201);
or U8549 (N_8549,N_8229,N_8327);
xnor U8550 (N_8550,N_8247,N_8346);
nand U8551 (N_8551,N_8241,N_8188);
xnor U8552 (N_8552,N_8210,N_8251);
or U8553 (N_8553,N_8280,N_8124);
nand U8554 (N_8554,N_8330,N_8130);
nand U8555 (N_8555,N_8355,N_8101);
xor U8556 (N_8556,N_8372,N_8257);
or U8557 (N_8557,N_8183,N_8281);
xnor U8558 (N_8558,N_8232,N_8229);
and U8559 (N_8559,N_8195,N_8126);
and U8560 (N_8560,N_8225,N_8311);
nand U8561 (N_8561,N_8384,N_8325);
nor U8562 (N_8562,N_8331,N_8351);
nand U8563 (N_8563,N_8347,N_8281);
and U8564 (N_8564,N_8300,N_8399);
nand U8565 (N_8565,N_8310,N_8187);
nand U8566 (N_8566,N_8178,N_8335);
xor U8567 (N_8567,N_8379,N_8237);
and U8568 (N_8568,N_8177,N_8238);
or U8569 (N_8569,N_8141,N_8306);
or U8570 (N_8570,N_8100,N_8204);
xnor U8571 (N_8571,N_8290,N_8286);
xor U8572 (N_8572,N_8276,N_8383);
or U8573 (N_8573,N_8302,N_8247);
xnor U8574 (N_8574,N_8174,N_8154);
nor U8575 (N_8575,N_8359,N_8301);
or U8576 (N_8576,N_8155,N_8280);
xnor U8577 (N_8577,N_8103,N_8168);
or U8578 (N_8578,N_8229,N_8325);
and U8579 (N_8579,N_8362,N_8381);
nor U8580 (N_8580,N_8109,N_8362);
xnor U8581 (N_8581,N_8144,N_8337);
or U8582 (N_8582,N_8201,N_8281);
or U8583 (N_8583,N_8188,N_8126);
nand U8584 (N_8584,N_8230,N_8239);
and U8585 (N_8585,N_8172,N_8251);
and U8586 (N_8586,N_8186,N_8130);
xnor U8587 (N_8587,N_8117,N_8334);
and U8588 (N_8588,N_8319,N_8307);
and U8589 (N_8589,N_8172,N_8201);
and U8590 (N_8590,N_8104,N_8135);
nor U8591 (N_8591,N_8386,N_8213);
nor U8592 (N_8592,N_8214,N_8171);
or U8593 (N_8593,N_8328,N_8244);
and U8594 (N_8594,N_8299,N_8398);
and U8595 (N_8595,N_8326,N_8124);
and U8596 (N_8596,N_8283,N_8151);
and U8597 (N_8597,N_8366,N_8380);
or U8598 (N_8598,N_8322,N_8308);
nand U8599 (N_8599,N_8363,N_8209);
nand U8600 (N_8600,N_8375,N_8334);
nand U8601 (N_8601,N_8178,N_8257);
nor U8602 (N_8602,N_8174,N_8228);
and U8603 (N_8603,N_8241,N_8248);
and U8604 (N_8604,N_8105,N_8333);
and U8605 (N_8605,N_8309,N_8301);
nor U8606 (N_8606,N_8105,N_8373);
xor U8607 (N_8607,N_8344,N_8220);
xor U8608 (N_8608,N_8264,N_8351);
or U8609 (N_8609,N_8374,N_8215);
or U8610 (N_8610,N_8194,N_8112);
nor U8611 (N_8611,N_8376,N_8116);
nor U8612 (N_8612,N_8293,N_8138);
nand U8613 (N_8613,N_8147,N_8295);
nand U8614 (N_8614,N_8249,N_8185);
nand U8615 (N_8615,N_8157,N_8100);
or U8616 (N_8616,N_8338,N_8164);
xnor U8617 (N_8617,N_8334,N_8330);
nand U8618 (N_8618,N_8346,N_8319);
xor U8619 (N_8619,N_8168,N_8362);
nor U8620 (N_8620,N_8278,N_8155);
or U8621 (N_8621,N_8113,N_8167);
xor U8622 (N_8622,N_8216,N_8353);
and U8623 (N_8623,N_8394,N_8182);
or U8624 (N_8624,N_8157,N_8136);
and U8625 (N_8625,N_8316,N_8223);
xor U8626 (N_8626,N_8376,N_8313);
nor U8627 (N_8627,N_8172,N_8100);
or U8628 (N_8628,N_8128,N_8138);
nand U8629 (N_8629,N_8166,N_8365);
nand U8630 (N_8630,N_8299,N_8243);
or U8631 (N_8631,N_8205,N_8226);
or U8632 (N_8632,N_8337,N_8172);
nand U8633 (N_8633,N_8259,N_8167);
nand U8634 (N_8634,N_8215,N_8337);
and U8635 (N_8635,N_8285,N_8157);
and U8636 (N_8636,N_8185,N_8347);
nand U8637 (N_8637,N_8291,N_8325);
xor U8638 (N_8638,N_8315,N_8334);
nor U8639 (N_8639,N_8374,N_8321);
or U8640 (N_8640,N_8275,N_8165);
nand U8641 (N_8641,N_8187,N_8374);
nor U8642 (N_8642,N_8263,N_8377);
nor U8643 (N_8643,N_8387,N_8160);
and U8644 (N_8644,N_8329,N_8252);
xor U8645 (N_8645,N_8149,N_8304);
nand U8646 (N_8646,N_8343,N_8315);
nor U8647 (N_8647,N_8218,N_8313);
and U8648 (N_8648,N_8243,N_8133);
nand U8649 (N_8649,N_8240,N_8142);
xnor U8650 (N_8650,N_8298,N_8331);
and U8651 (N_8651,N_8364,N_8111);
nand U8652 (N_8652,N_8293,N_8305);
or U8653 (N_8653,N_8163,N_8103);
nand U8654 (N_8654,N_8294,N_8317);
nor U8655 (N_8655,N_8257,N_8180);
xnor U8656 (N_8656,N_8363,N_8327);
or U8657 (N_8657,N_8366,N_8254);
and U8658 (N_8658,N_8390,N_8230);
nor U8659 (N_8659,N_8369,N_8236);
or U8660 (N_8660,N_8212,N_8347);
nand U8661 (N_8661,N_8168,N_8286);
nand U8662 (N_8662,N_8328,N_8250);
xor U8663 (N_8663,N_8336,N_8148);
nor U8664 (N_8664,N_8144,N_8152);
or U8665 (N_8665,N_8169,N_8371);
nand U8666 (N_8666,N_8345,N_8159);
or U8667 (N_8667,N_8264,N_8380);
nand U8668 (N_8668,N_8267,N_8395);
nand U8669 (N_8669,N_8134,N_8341);
xnor U8670 (N_8670,N_8251,N_8222);
nor U8671 (N_8671,N_8316,N_8262);
or U8672 (N_8672,N_8155,N_8390);
and U8673 (N_8673,N_8326,N_8117);
xnor U8674 (N_8674,N_8216,N_8168);
and U8675 (N_8675,N_8164,N_8184);
nor U8676 (N_8676,N_8186,N_8163);
nand U8677 (N_8677,N_8246,N_8300);
or U8678 (N_8678,N_8347,N_8155);
and U8679 (N_8679,N_8181,N_8314);
nand U8680 (N_8680,N_8293,N_8290);
and U8681 (N_8681,N_8174,N_8190);
and U8682 (N_8682,N_8261,N_8307);
or U8683 (N_8683,N_8232,N_8272);
nor U8684 (N_8684,N_8179,N_8271);
nand U8685 (N_8685,N_8106,N_8228);
or U8686 (N_8686,N_8137,N_8129);
and U8687 (N_8687,N_8159,N_8348);
or U8688 (N_8688,N_8272,N_8318);
and U8689 (N_8689,N_8115,N_8138);
nand U8690 (N_8690,N_8245,N_8202);
nand U8691 (N_8691,N_8396,N_8266);
nor U8692 (N_8692,N_8239,N_8138);
xnor U8693 (N_8693,N_8239,N_8399);
xor U8694 (N_8694,N_8289,N_8323);
nand U8695 (N_8695,N_8360,N_8320);
xnor U8696 (N_8696,N_8176,N_8346);
and U8697 (N_8697,N_8264,N_8299);
xnor U8698 (N_8698,N_8123,N_8221);
nor U8699 (N_8699,N_8259,N_8388);
nand U8700 (N_8700,N_8467,N_8604);
xor U8701 (N_8701,N_8549,N_8627);
or U8702 (N_8702,N_8502,N_8527);
nor U8703 (N_8703,N_8555,N_8656);
and U8704 (N_8704,N_8464,N_8667);
xor U8705 (N_8705,N_8426,N_8475);
and U8706 (N_8706,N_8674,N_8658);
and U8707 (N_8707,N_8542,N_8439);
nor U8708 (N_8708,N_8420,N_8451);
nand U8709 (N_8709,N_8414,N_8480);
or U8710 (N_8710,N_8533,N_8629);
nand U8711 (N_8711,N_8589,N_8540);
or U8712 (N_8712,N_8400,N_8639);
and U8713 (N_8713,N_8575,N_8406);
nor U8714 (N_8714,N_8423,N_8504);
or U8715 (N_8715,N_8476,N_8413);
nand U8716 (N_8716,N_8570,N_8671);
xor U8717 (N_8717,N_8500,N_8568);
and U8718 (N_8718,N_8490,N_8453);
and U8719 (N_8719,N_8548,N_8431);
nand U8720 (N_8720,N_8634,N_8421);
nand U8721 (N_8721,N_8447,N_8651);
or U8722 (N_8722,N_8507,N_8695);
xor U8723 (N_8723,N_8481,N_8586);
nor U8724 (N_8724,N_8641,N_8486);
nor U8725 (N_8725,N_8636,N_8443);
xor U8726 (N_8726,N_8583,N_8588);
or U8727 (N_8727,N_8638,N_8672);
or U8728 (N_8728,N_8498,N_8544);
or U8729 (N_8729,N_8462,N_8566);
and U8730 (N_8730,N_8644,N_8587);
xor U8731 (N_8731,N_8608,N_8428);
xnor U8732 (N_8732,N_8620,N_8687);
xor U8733 (N_8733,N_8492,N_8561);
or U8734 (N_8734,N_8622,N_8471);
or U8735 (N_8735,N_8616,N_8522);
or U8736 (N_8736,N_8433,N_8404);
nand U8737 (N_8737,N_8430,N_8693);
or U8738 (N_8738,N_8519,N_8485);
and U8739 (N_8739,N_8681,N_8611);
xor U8740 (N_8740,N_8654,N_8576);
xor U8741 (N_8741,N_8669,N_8553);
nand U8742 (N_8742,N_8605,N_8600);
xor U8743 (N_8743,N_8601,N_8624);
nand U8744 (N_8744,N_8596,N_8652);
xnor U8745 (N_8745,N_8625,N_8633);
and U8746 (N_8746,N_8528,N_8683);
xor U8747 (N_8747,N_8662,N_8455);
or U8748 (N_8748,N_8559,N_8469);
nand U8749 (N_8749,N_8564,N_8461);
and U8750 (N_8750,N_8456,N_8665);
or U8751 (N_8751,N_8673,N_8689);
or U8752 (N_8752,N_8445,N_8512);
or U8753 (N_8753,N_8440,N_8424);
nand U8754 (N_8754,N_8460,N_8621);
nor U8755 (N_8755,N_8686,N_8599);
and U8756 (N_8756,N_8628,N_8536);
nor U8757 (N_8757,N_8463,N_8554);
or U8758 (N_8758,N_8678,N_8403);
or U8759 (N_8759,N_8562,N_8525);
nand U8760 (N_8760,N_8594,N_8410);
or U8761 (N_8761,N_8565,N_8552);
nor U8762 (N_8762,N_8581,N_8493);
nor U8763 (N_8763,N_8432,N_8523);
xnor U8764 (N_8764,N_8541,N_8526);
and U8765 (N_8765,N_8574,N_8405);
xnor U8766 (N_8766,N_8524,N_8609);
and U8767 (N_8767,N_8670,N_8496);
nor U8768 (N_8768,N_8613,N_8535);
xor U8769 (N_8769,N_8545,N_8546);
xnor U8770 (N_8770,N_8560,N_8516);
and U8771 (N_8771,N_8450,N_8477);
or U8772 (N_8772,N_8547,N_8614);
and U8773 (N_8773,N_8680,N_8661);
or U8774 (N_8774,N_8513,N_8698);
nor U8775 (N_8775,N_8446,N_8538);
nand U8776 (N_8776,N_8408,N_8648);
xnor U8777 (N_8777,N_8517,N_8643);
or U8778 (N_8778,N_8473,N_8488);
nor U8779 (N_8779,N_8676,N_8584);
and U8780 (N_8780,N_8696,N_8598);
nor U8781 (N_8781,N_8466,N_8539);
nor U8782 (N_8782,N_8692,N_8407);
and U8783 (N_8783,N_8470,N_8556);
nor U8784 (N_8784,N_8657,N_8521);
and U8785 (N_8785,N_8697,N_8448);
nand U8786 (N_8786,N_8677,N_8646);
nor U8787 (N_8787,N_8663,N_8438);
xor U8788 (N_8788,N_8416,N_8543);
and U8789 (N_8789,N_8606,N_8690);
xor U8790 (N_8790,N_8412,N_8558);
or U8791 (N_8791,N_8664,N_8402);
nand U8792 (N_8792,N_8444,N_8623);
xor U8793 (N_8793,N_8573,N_8495);
and U8794 (N_8794,N_8668,N_8457);
nand U8795 (N_8795,N_8551,N_8579);
nor U8796 (N_8796,N_8452,N_8659);
nand U8797 (N_8797,N_8499,N_8653);
nor U8798 (N_8798,N_8422,N_8567);
and U8799 (N_8799,N_8691,N_8458);
and U8800 (N_8800,N_8617,N_8482);
nor U8801 (N_8801,N_8645,N_8563);
or U8802 (N_8802,N_8484,N_8637);
or U8803 (N_8803,N_8449,N_8590);
and U8804 (N_8804,N_8572,N_8468);
nand U8805 (N_8805,N_8514,N_8580);
nand U8806 (N_8806,N_8465,N_8497);
and U8807 (N_8807,N_8441,N_8427);
xor U8808 (N_8808,N_8534,N_8585);
nand U8809 (N_8809,N_8632,N_8603);
or U8810 (N_8810,N_8531,N_8626);
and U8811 (N_8811,N_8436,N_8635);
nor U8812 (N_8812,N_8532,N_8610);
xor U8813 (N_8813,N_8682,N_8592);
xnor U8814 (N_8814,N_8688,N_8655);
xnor U8815 (N_8815,N_8642,N_8518);
xor U8816 (N_8816,N_8631,N_8582);
nand U8817 (N_8817,N_8472,N_8602);
nand U8818 (N_8818,N_8649,N_8474);
xnor U8819 (N_8819,N_8675,N_8537);
xnor U8820 (N_8820,N_8515,N_8647);
nor U8821 (N_8821,N_8429,N_8607);
and U8822 (N_8822,N_8411,N_8684);
and U8823 (N_8823,N_8530,N_8419);
nor U8824 (N_8824,N_8415,N_8401);
or U8825 (N_8825,N_8501,N_8510);
nand U8826 (N_8826,N_8630,N_8694);
xnor U8827 (N_8827,N_8506,N_8434);
xor U8828 (N_8828,N_8494,N_8618);
nand U8829 (N_8829,N_8487,N_8550);
nand U8830 (N_8830,N_8511,N_8615);
and U8831 (N_8831,N_8520,N_8491);
and U8832 (N_8832,N_8578,N_8425);
xor U8833 (N_8833,N_8437,N_8509);
xor U8834 (N_8834,N_8666,N_8409);
or U8835 (N_8835,N_8612,N_8557);
nor U8836 (N_8836,N_8619,N_8529);
nand U8837 (N_8837,N_8505,N_8571);
nand U8838 (N_8838,N_8679,N_8597);
nand U8839 (N_8839,N_8685,N_8699);
and U8840 (N_8840,N_8640,N_8577);
nand U8841 (N_8841,N_8417,N_8478);
and U8842 (N_8842,N_8503,N_8660);
or U8843 (N_8843,N_8591,N_8459);
xor U8844 (N_8844,N_8479,N_8595);
xor U8845 (N_8845,N_8483,N_8442);
nand U8846 (N_8846,N_8508,N_8454);
xnor U8847 (N_8847,N_8435,N_8593);
or U8848 (N_8848,N_8569,N_8650);
and U8849 (N_8849,N_8418,N_8489);
nand U8850 (N_8850,N_8606,N_8500);
or U8851 (N_8851,N_8673,N_8685);
xor U8852 (N_8852,N_8647,N_8580);
nand U8853 (N_8853,N_8467,N_8582);
and U8854 (N_8854,N_8541,N_8559);
and U8855 (N_8855,N_8474,N_8647);
nand U8856 (N_8856,N_8621,N_8677);
and U8857 (N_8857,N_8500,N_8686);
nand U8858 (N_8858,N_8512,N_8562);
and U8859 (N_8859,N_8620,N_8632);
nand U8860 (N_8860,N_8515,N_8552);
nor U8861 (N_8861,N_8695,N_8669);
and U8862 (N_8862,N_8652,N_8416);
nand U8863 (N_8863,N_8642,N_8667);
nor U8864 (N_8864,N_8634,N_8438);
or U8865 (N_8865,N_8629,N_8633);
or U8866 (N_8866,N_8639,N_8446);
xnor U8867 (N_8867,N_8522,N_8573);
or U8868 (N_8868,N_8437,N_8598);
and U8869 (N_8869,N_8605,N_8653);
nor U8870 (N_8870,N_8489,N_8691);
xnor U8871 (N_8871,N_8550,N_8547);
and U8872 (N_8872,N_8518,N_8693);
and U8873 (N_8873,N_8513,N_8408);
nand U8874 (N_8874,N_8669,N_8401);
and U8875 (N_8875,N_8632,N_8462);
xnor U8876 (N_8876,N_8564,N_8522);
or U8877 (N_8877,N_8540,N_8485);
nand U8878 (N_8878,N_8683,N_8465);
or U8879 (N_8879,N_8472,N_8585);
xor U8880 (N_8880,N_8498,N_8508);
xor U8881 (N_8881,N_8537,N_8622);
nand U8882 (N_8882,N_8577,N_8486);
and U8883 (N_8883,N_8645,N_8531);
or U8884 (N_8884,N_8645,N_8480);
nand U8885 (N_8885,N_8644,N_8566);
nand U8886 (N_8886,N_8516,N_8639);
nor U8887 (N_8887,N_8530,N_8648);
nor U8888 (N_8888,N_8534,N_8681);
or U8889 (N_8889,N_8404,N_8487);
nor U8890 (N_8890,N_8482,N_8608);
and U8891 (N_8891,N_8450,N_8465);
nand U8892 (N_8892,N_8439,N_8409);
nor U8893 (N_8893,N_8453,N_8629);
and U8894 (N_8894,N_8623,N_8558);
and U8895 (N_8895,N_8430,N_8595);
nand U8896 (N_8896,N_8462,N_8515);
nor U8897 (N_8897,N_8602,N_8587);
nand U8898 (N_8898,N_8422,N_8698);
xor U8899 (N_8899,N_8687,N_8627);
nor U8900 (N_8900,N_8522,N_8407);
or U8901 (N_8901,N_8538,N_8449);
and U8902 (N_8902,N_8500,N_8459);
nor U8903 (N_8903,N_8527,N_8663);
xor U8904 (N_8904,N_8520,N_8576);
nand U8905 (N_8905,N_8457,N_8667);
xnor U8906 (N_8906,N_8402,N_8501);
nor U8907 (N_8907,N_8486,N_8633);
or U8908 (N_8908,N_8499,N_8519);
nor U8909 (N_8909,N_8691,N_8676);
nand U8910 (N_8910,N_8644,N_8511);
xor U8911 (N_8911,N_8676,N_8407);
and U8912 (N_8912,N_8563,N_8580);
or U8913 (N_8913,N_8404,N_8459);
or U8914 (N_8914,N_8568,N_8698);
nand U8915 (N_8915,N_8430,N_8538);
nor U8916 (N_8916,N_8451,N_8667);
nand U8917 (N_8917,N_8481,N_8695);
or U8918 (N_8918,N_8506,N_8419);
nor U8919 (N_8919,N_8474,N_8694);
xnor U8920 (N_8920,N_8459,N_8641);
nor U8921 (N_8921,N_8588,N_8599);
or U8922 (N_8922,N_8694,N_8665);
nor U8923 (N_8923,N_8683,N_8552);
or U8924 (N_8924,N_8643,N_8669);
or U8925 (N_8925,N_8401,N_8544);
or U8926 (N_8926,N_8427,N_8472);
and U8927 (N_8927,N_8401,N_8537);
or U8928 (N_8928,N_8662,N_8535);
and U8929 (N_8929,N_8490,N_8416);
xor U8930 (N_8930,N_8678,N_8499);
nand U8931 (N_8931,N_8543,N_8461);
or U8932 (N_8932,N_8551,N_8507);
and U8933 (N_8933,N_8400,N_8490);
nor U8934 (N_8934,N_8425,N_8641);
nor U8935 (N_8935,N_8688,N_8675);
nor U8936 (N_8936,N_8488,N_8408);
and U8937 (N_8937,N_8599,N_8600);
nand U8938 (N_8938,N_8678,N_8569);
xor U8939 (N_8939,N_8541,N_8699);
nor U8940 (N_8940,N_8669,N_8563);
nand U8941 (N_8941,N_8647,N_8694);
or U8942 (N_8942,N_8617,N_8650);
xor U8943 (N_8943,N_8550,N_8656);
nor U8944 (N_8944,N_8427,N_8521);
and U8945 (N_8945,N_8424,N_8427);
and U8946 (N_8946,N_8636,N_8621);
nand U8947 (N_8947,N_8583,N_8654);
nor U8948 (N_8948,N_8634,N_8612);
and U8949 (N_8949,N_8550,N_8494);
or U8950 (N_8950,N_8528,N_8565);
nor U8951 (N_8951,N_8413,N_8430);
xor U8952 (N_8952,N_8695,N_8483);
nor U8953 (N_8953,N_8432,N_8539);
or U8954 (N_8954,N_8476,N_8522);
nand U8955 (N_8955,N_8592,N_8414);
and U8956 (N_8956,N_8494,N_8579);
and U8957 (N_8957,N_8477,N_8572);
xor U8958 (N_8958,N_8624,N_8614);
nand U8959 (N_8959,N_8418,N_8650);
or U8960 (N_8960,N_8476,N_8617);
and U8961 (N_8961,N_8553,N_8442);
or U8962 (N_8962,N_8635,N_8677);
and U8963 (N_8963,N_8617,N_8571);
or U8964 (N_8964,N_8565,N_8419);
nand U8965 (N_8965,N_8566,N_8410);
and U8966 (N_8966,N_8449,N_8646);
nor U8967 (N_8967,N_8488,N_8555);
or U8968 (N_8968,N_8471,N_8406);
or U8969 (N_8969,N_8475,N_8545);
nand U8970 (N_8970,N_8646,N_8436);
xnor U8971 (N_8971,N_8571,N_8472);
nor U8972 (N_8972,N_8687,N_8500);
or U8973 (N_8973,N_8428,N_8678);
xnor U8974 (N_8974,N_8588,N_8641);
or U8975 (N_8975,N_8497,N_8541);
and U8976 (N_8976,N_8463,N_8581);
xnor U8977 (N_8977,N_8516,N_8481);
nand U8978 (N_8978,N_8511,N_8600);
xnor U8979 (N_8979,N_8437,N_8651);
and U8980 (N_8980,N_8508,N_8571);
nor U8981 (N_8981,N_8517,N_8510);
nand U8982 (N_8982,N_8402,N_8652);
and U8983 (N_8983,N_8645,N_8621);
or U8984 (N_8984,N_8539,N_8533);
nor U8985 (N_8985,N_8609,N_8552);
and U8986 (N_8986,N_8571,N_8698);
or U8987 (N_8987,N_8461,N_8482);
xnor U8988 (N_8988,N_8460,N_8401);
or U8989 (N_8989,N_8656,N_8542);
nor U8990 (N_8990,N_8559,N_8548);
and U8991 (N_8991,N_8612,N_8429);
xor U8992 (N_8992,N_8420,N_8640);
nor U8993 (N_8993,N_8639,N_8683);
nor U8994 (N_8994,N_8597,N_8510);
or U8995 (N_8995,N_8467,N_8436);
nor U8996 (N_8996,N_8480,N_8616);
or U8997 (N_8997,N_8469,N_8576);
or U8998 (N_8998,N_8615,N_8460);
nand U8999 (N_8999,N_8675,N_8666);
nand U9000 (N_9000,N_8830,N_8890);
or U9001 (N_9001,N_8978,N_8759);
xnor U9002 (N_9002,N_8885,N_8758);
nand U9003 (N_9003,N_8960,N_8993);
nor U9004 (N_9004,N_8748,N_8703);
or U9005 (N_9005,N_8826,N_8939);
nand U9006 (N_9006,N_8930,N_8980);
xnor U9007 (N_9007,N_8818,N_8805);
or U9008 (N_9008,N_8832,N_8743);
and U9009 (N_9009,N_8860,N_8902);
or U9010 (N_9010,N_8824,N_8907);
and U9011 (N_9011,N_8858,N_8976);
or U9012 (N_9012,N_8829,N_8793);
or U9013 (N_9013,N_8712,N_8956);
xor U9014 (N_9014,N_8945,N_8742);
or U9015 (N_9015,N_8903,N_8745);
nand U9016 (N_9016,N_8937,N_8822);
xor U9017 (N_9017,N_8773,N_8854);
and U9018 (N_9018,N_8875,N_8856);
nand U9019 (N_9019,N_8908,N_8869);
and U9020 (N_9020,N_8938,N_8844);
xnor U9021 (N_9021,N_8765,N_8861);
xor U9022 (N_9022,N_8749,N_8768);
nand U9023 (N_9023,N_8734,N_8896);
xor U9024 (N_9024,N_8986,N_8876);
xor U9025 (N_9025,N_8761,N_8819);
or U9026 (N_9026,N_8878,N_8729);
or U9027 (N_9027,N_8846,N_8931);
nor U9028 (N_9028,N_8925,N_8851);
xnor U9029 (N_9029,N_8871,N_8760);
nand U9030 (N_9030,N_8798,N_8811);
xnor U9031 (N_9031,N_8766,N_8927);
nor U9032 (N_9032,N_8895,N_8750);
or U9033 (N_9033,N_8794,N_8998);
nand U9034 (N_9034,N_8797,N_8840);
nand U9035 (N_9035,N_8954,N_8946);
and U9036 (N_9036,N_8736,N_8953);
or U9037 (N_9037,N_8916,N_8928);
and U9038 (N_9038,N_8912,N_8724);
xor U9039 (N_9039,N_8727,N_8800);
or U9040 (N_9040,N_8899,N_8834);
xnor U9041 (N_9041,N_8911,N_8786);
nor U9042 (N_9042,N_8702,N_8837);
or U9043 (N_9043,N_8877,N_8762);
xnor U9044 (N_9044,N_8725,N_8807);
nor U9045 (N_9045,N_8892,N_8873);
and U9046 (N_9046,N_8949,N_8728);
xnor U9047 (N_9047,N_8841,N_8905);
nand U9048 (N_9048,N_8988,N_8754);
and U9049 (N_9049,N_8992,N_8771);
nor U9050 (N_9050,N_8808,N_8792);
xnor U9051 (N_9051,N_8772,N_8733);
and U9052 (N_9052,N_8970,N_8744);
and U9053 (N_9053,N_8936,N_8780);
and U9054 (N_9054,N_8973,N_8842);
xor U9055 (N_9055,N_8801,N_8731);
xnor U9056 (N_9056,N_8787,N_8815);
or U9057 (N_9057,N_8906,N_8984);
nand U9058 (N_9058,N_8812,N_8955);
nor U9059 (N_9059,N_8894,N_8763);
xnor U9060 (N_9060,N_8884,N_8940);
nor U9061 (N_9061,N_8726,N_8710);
or U9062 (N_9062,N_8926,N_8962);
xor U9063 (N_9063,N_8747,N_8880);
nand U9064 (N_9064,N_8923,N_8828);
and U9065 (N_9065,N_8838,N_8823);
and U9066 (N_9066,N_8974,N_8806);
nand U9067 (N_9067,N_8817,N_8847);
nand U9068 (N_9068,N_8757,N_8722);
nand U9069 (N_9069,N_8782,N_8755);
nor U9070 (N_9070,N_8967,N_8879);
nand U9071 (N_9071,N_8803,N_8966);
nand U9072 (N_9072,N_8713,N_8735);
and U9073 (N_9073,N_8843,N_8770);
nor U9074 (N_9074,N_8999,N_8900);
nand U9075 (N_9075,N_8882,N_8752);
nand U9076 (N_9076,N_8715,N_8718);
and U9077 (N_9077,N_8711,N_8987);
or U9078 (N_9078,N_8738,N_8746);
and U9079 (N_9079,N_8705,N_8972);
nor U9080 (N_9080,N_8753,N_8975);
nand U9081 (N_9081,N_8917,N_8821);
xnor U9082 (N_9082,N_8985,N_8950);
nor U9083 (N_9083,N_8891,N_8933);
xor U9084 (N_9084,N_8741,N_8921);
nor U9085 (N_9085,N_8706,N_8716);
xor U9086 (N_9086,N_8827,N_8951);
or U9087 (N_9087,N_8957,N_8901);
nor U9088 (N_9088,N_8979,N_8810);
nand U9089 (N_9089,N_8932,N_8717);
nor U9090 (N_9090,N_8777,N_8935);
and U9091 (N_9091,N_8839,N_8971);
nand U9092 (N_9092,N_8996,N_8784);
nand U9093 (N_9093,N_8790,N_8701);
nor U9094 (N_9094,N_8835,N_8852);
nor U9095 (N_9095,N_8809,N_8989);
nor U9096 (N_9096,N_8977,N_8994);
or U9097 (N_9097,N_8789,N_8751);
nand U9098 (N_9098,N_8934,N_8774);
and U9099 (N_9099,N_8816,N_8796);
nor U9100 (N_9100,N_8700,N_8963);
nand U9101 (N_9101,N_8920,N_8732);
nor U9102 (N_9102,N_8874,N_8922);
nor U9103 (N_9103,N_8775,N_8855);
and U9104 (N_9104,N_8862,N_8886);
nand U9105 (N_9105,N_8866,N_8850);
and U9106 (N_9106,N_8959,N_8958);
or U9107 (N_9107,N_8943,N_8785);
and U9108 (N_9108,N_8929,N_8991);
nand U9109 (N_9109,N_8888,N_8964);
xor U9110 (N_9110,N_8941,N_8825);
xor U9111 (N_9111,N_8887,N_8769);
xor U9112 (N_9112,N_8864,N_8981);
nand U9113 (N_9113,N_8863,N_8969);
nand U9114 (N_9114,N_8883,N_8730);
xnor U9115 (N_9115,N_8704,N_8948);
nand U9116 (N_9116,N_8898,N_8952);
or U9117 (N_9117,N_8804,N_8914);
and U9118 (N_9118,N_8776,N_8719);
nor U9119 (N_9119,N_8942,N_8791);
nand U9120 (N_9120,N_8709,N_8767);
xnor U9121 (N_9121,N_8965,N_8737);
nand U9122 (N_9122,N_8783,N_8918);
xnor U9123 (N_9123,N_8919,N_8802);
or U9124 (N_9124,N_8995,N_8909);
xor U9125 (N_9125,N_8947,N_8764);
xor U9126 (N_9126,N_8788,N_8814);
nand U9127 (N_9127,N_8756,N_8961);
nor U9128 (N_9128,N_8872,N_8913);
and U9129 (N_9129,N_8868,N_8848);
and U9130 (N_9130,N_8897,N_8833);
nand U9131 (N_9131,N_8723,N_8795);
nand U9132 (N_9132,N_8849,N_8720);
or U9133 (N_9133,N_8857,N_8944);
and U9134 (N_9134,N_8831,N_8910);
xnor U9135 (N_9135,N_8836,N_8997);
or U9136 (N_9136,N_8740,N_8721);
xor U9137 (N_9137,N_8982,N_8904);
xnor U9138 (N_9138,N_8708,N_8845);
or U9139 (N_9139,N_8865,N_8853);
nor U9140 (N_9140,N_8739,N_8781);
and U9141 (N_9141,N_8924,N_8983);
nor U9142 (N_9142,N_8813,N_8859);
nand U9143 (N_9143,N_8799,N_8867);
nand U9144 (N_9144,N_8820,N_8889);
nand U9145 (N_9145,N_8870,N_8778);
and U9146 (N_9146,N_8779,N_8968);
nor U9147 (N_9147,N_8714,N_8881);
xor U9148 (N_9148,N_8707,N_8915);
nand U9149 (N_9149,N_8893,N_8990);
nand U9150 (N_9150,N_8943,N_8981);
and U9151 (N_9151,N_8895,N_8837);
and U9152 (N_9152,N_8876,N_8702);
and U9153 (N_9153,N_8810,N_8977);
nor U9154 (N_9154,N_8993,N_8974);
and U9155 (N_9155,N_8927,N_8850);
and U9156 (N_9156,N_8975,N_8978);
xor U9157 (N_9157,N_8882,N_8721);
nor U9158 (N_9158,N_8746,N_8986);
or U9159 (N_9159,N_8873,N_8742);
nor U9160 (N_9160,N_8776,N_8892);
nand U9161 (N_9161,N_8919,N_8984);
xnor U9162 (N_9162,N_8826,N_8914);
or U9163 (N_9163,N_8932,N_8732);
xor U9164 (N_9164,N_8701,N_8853);
nor U9165 (N_9165,N_8847,N_8905);
and U9166 (N_9166,N_8821,N_8905);
nand U9167 (N_9167,N_8863,N_8774);
nand U9168 (N_9168,N_8809,N_8992);
nand U9169 (N_9169,N_8898,N_8853);
nand U9170 (N_9170,N_8793,N_8710);
xor U9171 (N_9171,N_8806,N_8885);
or U9172 (N_9172,N_8710,N_8873);
nor U9173 (N_9173,N_8757,N_8763);
nand U9174 (N_9174,N_8821,N_8877);
nor U9175 (N_9175,N_8803,N_8937);
xor U9176 (N_9176,N_8771,N_8884);
and U9177 (N_9177,N_8777,N_8797);
or U9178 (N_9178,N_8867,N_8986);
xor U9179 (N_9179,N_8731,N_8977);
nor U9180 (N_9180,N_8754,N_8862);
xor U9181 (N_9181,N_8742,N_8906);
or U9182 (N_9182,N_8845,N_8978);
nand U9183 (N_9183,N_8838,N_8958);
nor U9184 (N_9184,N_8763,N_8884);
and U9185 (N_9185,N_8854,N_8772);
nor U9186 (N_9186,N_8946,N_8957);
or U9187 (N_9187,N_8740,N_8851);
nor U9188 (N_9188,N_8979,N_8877);
nor U9189 (N_9189,N_8822,N_8740);
xor U9190 (N_9190,N_8852,N_8952);
xnor U9191 (N_9191,N_8773,N_8903);
xnor U9192 (N_9192,N_8994,N_8870);
and U9193 (N_9193,N_8792,N_8813);
and U9194 (N_9194,N_8789,N_8730);
nand U9195 (N_9195,N_8906,N_8779);
nand U9196 (N_9196,N_8837,N_8950);
or U9197 (N_9197,N_8892,N_8934);
xor U9198 (N_9198,N_8830,N_8889);
nor U9199 (N_9199,N_8777,N_8773);
xor U9200 (N_9200,N_8708,N_8871);
nand U9201 (N_9201,N_8702,N_8940);
xor U9202 (N_9202,N_8925,N_8939);
xnor U9203 (N_9203,N_8781,N_8810);
nor U9204 (N_9204,N_8723,N_8729);
nand U9205 (N_9205,N_8847,N_8881);
or U9206 (N_9206,N_8955,N_8859);
xnor U9207 (N_9207,N_8872,N_8935);
or U9208 (N_9208,N_8767,N_8944);
nand U9209 (N_9209,N_8902,N_8976);
xor U9210 (N_9210,N_8924,N_8885);
nor U9211 (N_9211,N_8755,N_8839);
and U9212 (N_9212,N_8943,N_8845);
or U9213 (N_9213,N_8943,N_8862);
and U9214 (N_9214,N_8851,N_8845);
nand U9215 (N_9215,N_8706,N_8714);
xor U9216 (N_9216,N_8716,N_8974);
xor U9217 (N_9217,N_8751,N_8772);
nor U9218 (N_9218,N_8915,N_8929);
or U9219 (N_9219,N_8866,N_8795);
xnor U9220 (N_9220,N_8840,N_8806);
xnor U9221 (N_9221,N_8833,N_8966);
and U9222 (N_9222,N_8836,N_8760);
or U9223 (N_9223,N_8895,N_8774);
xnor U9224 (N_9224,N_8846,N_8705);
xor U9225 (N_9225,N_8906,N_8989);
nor U9226 (N_9226,N_8949,N_8930);
xor U9227 (N_9227,N_8725,N_8822);
xnor U9228 (N_9228,N_8898,N_8928);
and U9229 (N_9229,N_8757,N_8884);
nand U9230 (N_9230,N_8934,N_8867);
xnor U9231 (N_9231,N_8768,N_8799);
xor U9232 (N_9232,N_8747,N_8785);
and U9233 (N_9233,N_8832,N_8993);
nand U9234 (N_9234,N_8901,N_8966);
nor U9235 (N_9235,N_8705,N_8865);
and U9236 (N_9236,N_8747,N_8958);
and U9237 (N_9237,N_8963,N_8892);
or U9238 (N_9238,N_8842,N_8805);
or U9239 (N_9239,N_8773,N_8747);
and U9240 (N_9240,N_8776,N_8782);
or U9241 (N_9241,N_8888,N_8946);
or U9242 (N_9242,N_8730,N_8722);
and U9243 (N_9243,N_8752,N_8869);
or U9244 (N_9244,N_8928,N_8750);
or U9245 (N_9245,N_8992,N_8792);
xnor U9246 (N_9246,N_8728,N_8901);
and U9247 (N_9247,N_8729,N_8788);
nand U9248 (N_9248,N_8822,N_8715);
or U9249 (N_9249,N_8794,N_8744);
and U9250 (N_9250,N_8875,N_8721);
and U9251 (N_9251,N_8801,N_8916);
xnor U9252 (N_9252,N_8972,N_8939);
nor U9253 (N_9253,N_8745,N_8774);
or U9254 (N_9254,N_8899,N_8869);
nor U9255 (N_9255,N_8909,N_8931);
nand U9256 (N_9256,N_8962,N_8985);
xor U9257 (N_9257,N_8766,N_8861);
nand U9258 (N_9258,N_8894,N_8837);
nor U9259 (N_9259,N_8944,N_8973);
nand U9260 (N_9260,N_8920,N_8996);
or U9261 (N_9261,N_8827,N_8784);
or U9262 (N_9262,N_8990,N_8756);
nand U9263 (N_9263,N_8991,N_8833);
nor U9264 (N_9264,N_8792,N_8727);
xnor U9265 (N_9265,N_8809,N_8751);
and U9266 (N_9266,N_8731,N_8743);
nand U9267 (N_9267,N_8913,N_8778);
nor U9268 (N_9268,N_8733,N_8763);
and U9269 (N_9269,N_8820,N_8702);
and U9270 (N_9270,N_8872,N_8714);
or U9271 (N_9271,N_8915,N_8837);
xor U9272 (N_9272,N_8739,N_8925);
xnor U9273 (N_9273,N_8898,N_8706);
nor U9274 (N_9274,N_8744,N_8844);
xnor U9275 (N_9275,N_8892,N_8832);
nand U9276 (N_9276,N_8880,N_8864);
and U9277 (N_9277,N_8978,N_8797);
or U9278 (N_9278,N_8864,N_8906);
nor U9279 (N_9279,N_8725,N_8730);
xor U9280 (N_9280,N_8971,N_8906);
nand U9281 (N_9281,N_8862,N_8728);
and U9282 (N_9282,N_8879,N_8736);
xor U9283 (N_9283,N_8867,N_8742);
or U9284 (N_9284,N_8904,N_8743);
xnor U9285 (N_9285,N_8927,N_8750);
nor U9286 (N_9286,N_8717,N_8747);
nand U9287 (N_9287,N_8886,N_8721);
and U9288 (N_9288,N_8898,N_8870);
xnor U9289 (N_9289,N_8932,N_8982);
or U9290 (N_9290,N_8930,N_8928);
nand U9291 (N_9291,N_8774,N_8770);
xnor U9292 (N_9292,N_8796,N_8766);
or U9293 (N_9293,N_8783,N_8724);
nand U9294 (N_9294,N_8838,N_8700);
nor U9295 (N_9295,N_8841,N_8896);
nor U9296 (N_9296,N_8880,N_8995);
nand U9297 (N_9297,N_8789,N_8967);
nand U9298 (N_9298,N_8878,N_8726);
nor U9299 (N_9299,N_8796,N_8895);
nand U9300 (N_9300,N_9101,N_9075);
or U9301 (N_9301,N_9264,N_9218);
or U9302 (N_9302,N_9076,N_9277);
and U9303 (N_9303,N_9027,N_9220);
or U9304 (N_9304,N_9250,N_9071);
and U9305 (N_9305,N_9169,N_9286);
xor U9306 (N_9306,N_9179,N_9156);
nor U9307 (N_9307,N_9193,N_9161);
and U9308 (N_9308,N_9280,N_9049);
nor U9309 (N_9309,N_9154,N_9162);
or U9310 (N_9310,N_9257,N_9092);
nor U9311 (N_9311,N_9270,N_9108);
or U9312 (N_9312,N_9096,N_9068);
nand U9313 (N_9313,N_9039,N_9278);
or U9314 (N_9314,N_9177,N_9145);
and U9315 (N_9315,N_9007,N_9082);
and U9316 (N_9316,N_9000,N_9202);
nand U9317 (N_9317,N_9015,N_9104);
nor U9318 (N_9318,N_9139,N_9146);
nand U9319 (N_9319,N_9002,N_9237);
nor U9320 (N_9320,N_9234,N_9091);
nor U9321 (N_9321,N_9095,N_9038);
or U9322 (N_9322,N_9013,N_9080);
nor U9323 (N_9323,N_9230,N_9070);
nor U9324 (N_9324,N_9133,N_9191);
nand U9325 (N_9325,N_9040,N_9164);
xnor U9326 (N_9326,N_9273,N_9026);
xnor U9327 (N_9327,N_9229,N_9131);
xor U9328 (N_9328,N_9195,N_9119);
nand U9329 (N_9329,N_9276,N_9054);
and U9330 (N_9330,N_9217,N_9248);
nand U9331 (N_9331,N_9186,N_9142);
or U9332 (N_9332,N_9099,N_9228);
or U9333 (N_9333,N_9214,N_9023);
nand U9334 (N_9334,N_9051,N_9223);
nor U9335 (N_9335,N_9028,N_9106);
xnor U9336 (N_9336,N_9135,N_9100);
or U9337 (N_9337,N_9073,N_9094);
xor U9338 (N_9338,N_9261,N_9034);
nand U9339 (N_9339,N_9182,N_9287);
and U9340 (N_9340,N_9187,N_9019);
xor U9341 (N_9341,N_9173,N_9282);
nor U9342 (N_9342,N_9134,N_9235);
and U9343 (N_9343,N_9275,N_9102);
xnor U9344 (N_9344,N_9140,N_9292);
nor U9345 (N_9345,N_9188,N_9215);
xnor U9346 (N_9346,N_9009,N_9242);
xor U9347 (N_9347,N_9160,N_9246);
and U9348 (N_9348,N_9059,N_9090);
xor U9349 (N_9349,N_9231,N_9258);
xor U9350 (N_9350,N_9152,N_9114);
xor U9351 (N_9351,N_9201,N_9239);
nand U9352 (N_9352,N_9232,N_9016);
xnor U9353 (N_9353,N_9065,N_9003);
xnor U9354 (N_9354,N_9299,N_9168);
xor U9355 (N_9355,N_9115,N_9124);
xnor U9356 (N_9356,N_9185,N_9022);
or U9357 (N_9357,N_9271,N_9151);
and U9358 (N_9358,N_9132,N_9253);
or U9359 (N_9359,N_9021,N_9204);
and U9360 (N_9360,N_9172,N_9005);
and U9361 (N_9361,N_9233,N_9084);
or U9362 (N_9362,N_9128,N_9295);
and U9363 (N_9363,N_9254,N_9057);
nand U9364 (N_9364,N_9157,N_9180);
xor U9365 (N_9365,N_9098,N_9171);
or U9366 (N_9366,N_9155,N_9196);
xor U9367 (N_9367,N_9066,N_9121);
or U9368 (N_9368,N_9285,N_9159);
or U9369 (N_9369,N_9227,N_9127);
nand U9370 (N_9370,N_9004,N_9208);
nor U9371 (N_9371,N_9052,N_9263);
or U9372 (N_9372,N_9024,N_9194);
and U9373 (N_9373,N_9032,N_9060);
or U9374 (N_9374,N_9093,N_9089);
nand U9375 (N_9375,N_9291,N_9043);
or U9376 (N_9376,N_9141,N_9125);
xnor U9377 (N_9377,N_9031,N_9249);
and U9378 (N_9378,N_9211,N_9033);
and U9379 (N_9379,N_9255,N_9297);
xnor U9380 (N_9380,N_9126,N_9298);
nand U9381 (N_9381,N_9199,N_9097);
nand U9382 (N_9382,N_9018,N_9283);
xor U9383 (N_9383,N_9206,N_9175);
and U9384 (N_9384,N_9165,N_9219);
and U9385 (N_9385,N_9063,N_9259);
xnor U9386 (N_9386,N_9281,N_9158);
or U9387 (N_9387,N_9107,N_9244);
and U9388 (N_9388,N_9147,N_9025);
nor U9389 (N_9389,N_9120,N_9269);
or U9390 (N_9390,N_9061,N_9110);
or U9391 (N_9391,N_9224,N_9085);
and U9392 (N_9392,N_9113,N_9045);
or U9393 (N_9393,N_9176,N_9088);
xor U9394 (N_9394,N_9267,N_9056);
or U9395 (N_9395,N_9279,N_9138);
xor U9396 (N_9396,N_9086,N_9046);
nor U9397 (N_9397,N_9037,N_9178);
or U9398 (N_9398,N_9190,N_9137);
or U9399 (N_9399,N_9247,N_9011);
or U9400 (N_9400,N_9166,N_9130);
or U9401 (N_9401,N_9055,N_9200);
or U9402 (N_9402,N_9198,N_9243);
nor U9403 (N_9403,N_9036,N_9014);
and U9404 (N_9404,N_9058,N_9163);
nand U9405 (N_9405,N_9020,N_9077);
and U9406 (N_9406,N_9212,N_9112);
and U9407 (N_9407,N_9296,N_9047);
nand U9408 (N_9408,N_9221,N_9245);
nor U9409 (N_9409,N_9150,N_9167);
xor U9410 (N_9410,N_9064,N_9029);
nor U9411 (N_9411,N_9111,N_9213);
and U9412 (N_9412,N_9240,N_9181);
or U9413 (N_9413,N_9251,N_9222);
or U9414 (N_9414,N_9216,N_9050);
nor U9415 (N_9415,N_9153,N_9048);
nor U9416 (N_9416,N_9262,N_9288);
and U9417 (N_9417,N_9226,N_9174);
xnor U9418 (N_9418,N_9017,N_9256);
and U9419 (N_9419,N_9192,N_9122);
or U9420 (N_9420,N_9260,N_9268);
nand U9421 (N_9421,N_9207,N_9197);
xor U9422 (N_9422,N_9083,N_9143);
nand U9423 (N_9423,N_9241,N_9044);
nor U9424 (N_9424,N_9118,N_9284);
nor U9425 (N_9425,N_9236,N_9105);
and U9426 (N_9426,N_9148,N_9069);
or U9427 (N_9427,N_9203,N_9074);
or U9428 (N_9428,N_9274,N_9144);
or U9429 (N_9429,N_9170,N_9081);
nand U9430 (N_9430,N_9129,N_9006);
or U9431 (N_9431,N_9189,N_9184);
or U9432 (N_9432,N_9290,N_9205);
and U9433 (N_9433,N_9008,N_9252);
nor U9434 (N_9434,N_9001,N_9010);
and U9435 (N_9435,N_9012,N_9289);
or U9436 (N_9436,N_9272,N_9136);
xor U9437 (N_9437,N_9067,N_9078);
nor U9438 (N_9438,N_9103,N_9293);
nand U9439 (N_9439,N_9238,N_9035);
xnor U9440 (N_9440,N_9117,N_9210);
nand U9441 (N_9441,N_9116,N_9225);
and U9442 (N_9442,N_9109,N_9079);
or U9443 (N_9443,N_9209,N_9072);
nor U9444 (N_9444,N_9294,N_9041);
nor U9445 (N_9445,N_9265,N_9087);
and U9446 (N_9446,N_9123,N_9149);
xor U9447 (N_9447,N_9183,N_9030);
and U9448 (N_9448,N_9042,N_9053);
or U9449 (N_9449,N_9062,N_9266);
and U9450 (N_9450,N_9295,N_9229);
or U9451 (N_9451,N_9136,N_9199);
and U9452 (N_9452,N_9131,N_9270);
nand U9453 (N_9453,N_9020,N_9002);
or U9454 (N_9454,N_9184,N_9088);
nor U9455 (N_9455,N_9260,N_9067);
or U9456 (N_9456,N_9104,N_9094);
or U9457 (N_9457,N_9199,N_9180);
xor U9458 (N_9458,N_9048,N_9160);
and U9459 (N_9459,N_9050,N_9232);
xnor U9460 (N_9460,N_9075,N_9256);
or U9461 (N_9461,N_9145,N_9091);
xnor U9462 (N_9462,N_9200,N_9075);
nand U9463 (N_9463,N_9068,N_9027);
or U9464 (N_9464,N_9129,N_9192);
or U9465 (N_9465,N_9242,N_9257);
xnor U9466 (N_9466,N_9283,N_9095);
xor U9467 (N_9467,N_9096,N_9026);
and U9468 (N_9468,N_9092,N_9128);
and U9469 (N_9469,N_9108,N_9050);
nand U9470 (N_9470,N_9082,N_9103);
xor U9471 (N_9471,N_9218,N_9128);
nor U9472 (N_9472,N_9036,N_9025);
or U9473 (N_9473,N_9195,N_9086);
xor U9474 (N_9474,N_9036,N_9227);
xor U9475 (N_9475,N_9098,N_9130);
xnor U9476 (N_9476,N_9243,N_9212);
and U9477 (N_9477,N_9113,N_9013);
nor U9478 (N_9478,N_9115,N_9056);
and U9479 (N_9479,N_9212,N_9211);
and U9480 (N_9480,N_9127,N_9067);
nand U9481 (N_9481,N_9230,N_9196);
and U9482 (N_9482,N_9082,N_9116);
nor U9483 (N_9483,N_9196,N_9142);
nand U9484 (N_9484,N_9195,N_9112);
or U9485 (N_9485,N_9059,N_9120);
or U9486 (N_9486,N_9059,N_9263);
xnor U9487 (N_9487,N_9215,N_9220);
or U9488 (N_9488,N_9162,N_9101);
or U9489 (N_9489,N_9182,N_9216);
and U9490 (N_9490,N_9223,N_9065);
nor U9491 (N_9491,N_9029,N_9066);
nor U9492 (N_9492,N_9012,N_9097);
nand U9493 (N_9493,N_9271,N_9040);
nand U9494 (N_9494,N_9013,N_9150);
or U9495 (N_9495,N_9221,N_9125);
and U9496 (N_9496,N_9024,N_9079);
nand U9497 (N_9497,N_9092,N_9262);
or U9498 (N_9498,N_9102,N_9020);
nand U9499 (N_9499,N_9028,N_9110);
and U9500 (N_9500,N_9116,N_9198);
or U9501 (N_9501,N_9164,N_9193);
and U9502 (N_9502,N_9033,N_9206);
or U9503 (N_9503,N_9090,N_9227);
nand U9504 (N_9504,N_9100,N_9143);
and U9505 (N_9505,N_9254,N_9003);
and U9506 (N_9506,N_9171,N_9177);
or U9507 (N_9507,N_9150,N_9027);
xor U9508 (N_9508,N_9283,N_9035);
nor U9509 (N_9509,N_9179,N_9029);
and U9510 (N_9510,N_9212,N_9244);
or U9511 (N_9511,N_9182,N_9154);
nor U9512 (N_9512,N_9196,N_9182);
nand U9513 (N_9513,N_9003,N_9242);
nor U9514 (N_9514,N_9009,N_9127);
nor U9515 (N_9515,N_9194,N_9157);
xor U9516 (N_9516,N_9236,N_9220);
xor U9517 (N_9517,N_9032,N_9274);
or U9518 (N_9518,N_9041,N_9229);
nor U9519 (N_9519,N_9069,N_9255);
or U9520 (N_9520,N_9049,N_9228);
nor U9521 (N_9521,N_9104,N_9156);
and U9522 (N_9522,N_9207,N_9185);
or U9523 (N_9523,N_9091,N_9131);
xor U9524 (N_9524,N_9065,N_9157);
and U9525 (N_9525,N_9141,N_9151);
or U9526 (N_9526,N_9227,N_9254);
xor U9527 (N_9527,N_9267,N_9106);
nor U9528 (N_9528,N_9208,N_9225);
xnor U9529 (N_9529,N_9282,N_9012);
nor U9530 (N_9530,N_9183,N_9128);
nand U9531 (N_9531,N_9181,N_9019);
nand U9532 (N_9532,N_9145,N_9016);
nand U9533 (N_9533,N_9152,N_9288);
nor U9534 (N_9534,N_9065,N_9218);
nand U9535 (N_9535,N_9261,N_9019);
xor U9536 (N_9536,N_9235,N_9260);
nand U9537 (N_9537,N_9082,N_9061);
or U9538 (N_9538,N_9155,N_9098);
and U9539 (N_9539,N_9189,N_9188);
nor U9540 (N_9540,N_9224,N_9076);
and U9541 (N_9541,N_9201,N_9025);
xor U9542 (N_9542,N_9206,N_9204);
or U9543 (N_9543,N_9104,N_9288);
or U9544 (N_9544,N_9296,N_9227);
and U9545 (N_9545,N_9192,N_9185);
nand U9546 (N_9546,N_9240,N_9270);
xor U9547 (N_9547,N_9176,N_9201);
nor U9548 (N_9548,N_9062,N_9269);
xnor U9549 (N_9549,N_9219,N_9262);
xnor U9550 (N_9550,N_9246,N_9182);
xor U9551 (N_9551,N_9154,N_9221);
xnor U9552 (N_9552,N_9214,N_9120);
nor U9553 (N_9553,N_9042,N_9265);
or U9554 (N_9554,N_9097,N_9294);
or U9555 (N_9555,N_9273,N_9099);
xnor U9556 (N_9556,N_9120,N_9083);
nor U9557 (N_9557,N_9265,N_9145);
nand U9558 (N_9558,N_9101,N_9079);
nand U9559 (N_9559,N_9296,N_9157);
and U9560 (N_9560,N_9097,N_9237);
xor U9561 (N_9561,N_9251,N_9288);
nor U9562 (N_9562,N_9029,N_9156);
or U9563 (N_9563,N_9093,N_9256);
xnor U9564 (N_9564,N_9090,N_9165);
xor U9565 (N_9565,N_9065,N_9214);
and U9566 (N_9566,N_9067,N_9002);
or U9567 (N_9567,N_9280,N_9256);
and U9568 (N_9568,N_9146,N_9135);
and U9569 (N_9569,N_9222,N_9215);
nor U9570 (N_9570,N_9234,N_9220);
xor U9571 (N_9571,N_9008,N_9042);
xnor U9572 (N_9572,N_9218,N_9099);
xnor U9573 (N_9573,N_9271,N_9028);
nor U9574 (N_9574,N_9027,N_9241);
and U9575 (N_9575,N_9224,N_9075);
nor U9576 (N_9576,N_9012,N_9075);
nor U9577 (N_9577,N_9151,N_9205);
or U9578 (N_9578,N_9233,N_9149);
nor U9579 (N_9579,N_9109,N_9184);
xor U9580 (N_9580,N_9161,N_9113);
xnor U9581 (N_9581,N_9183,N_9113);
or U9582 (N_9582,N_9131,N_9288);
nand U9583 (N_9583,N_9267,N_9166);
or U9584 (N_9584,N_9191,N_9233);
or U9585 (N_9585,N_9089,N_9196);
nor U9586 (N_9586,N_9238,N_9275);
and U9587 (N_9587,N_9025,N_9285);
xnor U9588 (N_9588,N_9161,N_9145);
and U9589 (N_9589,N_9040,N_9112);
nor U9590 (N_9590,N_9289,N_9117);
nor U9591 (N_9591,N_9163,N_9293);
or U9592 (N_9592,N_9040,N_9169);
and U9593 (N_9593,N_9132,N_9284);
or U9594 (N_9594,N_9209,N_9071);
and U9595 (N_9595,N_9044,N_9141);
nand U9596 (N_9596,N_9235,N_9158);
and U9597 (N_9597,N_9088,N_9121);
nor U9598 (N_9598,N_9269,N_9282);
nor U9599 (N_9599,N_9189,N_9243);
xor U9600 (N_9600,N_9309,N_9484);
nor U9601 (N_9601,N_9599,N_9576);
or U9602 (N_9602,N_9594,N_9445);
nor U9603 (N_9603,N_9429,N_9418);
or U9604 (N_9604,N_9520,N_9427);
or U9605 (N_9605,N_9317,N_9305);
xnor U9606 (N_9606,N_9479,N_9423);
nand U9607 (N_9607,N_9453,N_9425);
xnor U9608 (N_9608,N_9416,N_9442);
nand U9609 (N_9609,N_9395,N_9568);
xnor U9610 (N_9610,N_9478,N_9308);
and U9611 (N_9611,N_9525,N_9513);
and U9612 (N_9612,N_9476,N_9336);
nor U9613 (N_9613,N_9417,N_9539);
nor U9614 (N_9614,N_9583,N_9311);
or U9615 (N_9615,N_9567,N_9443);
xor U9616 (N_9616,N_9329,N_9388);
nand U9617 (N_9617,N_9385,N_9335);
xnor U9618 (N_9618,N_9447,N_9468);
xnor U9619 (N_9619,N_9566,N_9362);
or U9620 (N_9620,N_9565,N_9350);
nand U9621 (N_9621,N_9454,N_9545);
nor U9622 (N_9622,N_9538,N_9482);
nor U9623 (N_9623,N_9526,N_9592);
nor U9624 (N_9624,N_9507,N_9521);
nand U9625 (N_9625,N_9316,N_9352);
nor U9626 (N_9626,N_9575,N_9561);
nor U9627 (N_9627,N_9318,N_9499);
xor U9628 (N_9628,N_9422,N_9304);
nand U9629 (N_9629,N_9370,N_9574);
or U9630 (N_9630,N_9589,N_9436);
and U9631 (N_9631,N_9483,N_9344);
nand U9632 (N_9632,N_9456,N_9477);
and U9633 (N_9633,N_9300,N_9364);
or U9634 (N_9634,N_9307,N_9514);
nand U9635 (N_9635,N_9532,N_9371);
nor U9636 (N_9636,N_9383,N_9314);
xnor U9637 (N_9637,N_9377,N_9597);
and U9638 (N_9638,N_9387,N_9508);
or U9639 (N_9639,N_9480,N_9515);
or U9640 (N_9640,N_9459,N_9342);
nand U9641 (N_9641,N_9426,N_9518);
nand U9642 (N_9642,N_9376,N_9501);
or U9643 (N_9643,N_9503,N_9546);
nor U9644 (N_9644,N_9455,N_9366);
nand U9645 (N_9645,N_9412,N_9558);
nor U9646 (N_9646,N_9319,N_9542);
nor U9647 (N_9647,N_9461,N_9560);
and U9648 (N_9648,N_9348,N_9509);
xnor U9649 (N_9649,N_9511,N_9487);
xor U9650 (N_9650,N_9524,N_9504);
xor U9651 (N_9651,N_9301,N_9533);
nand U9652 (N_9652,N_9552,N_9578);
or U9653 (N_9653,N_9506,N_9323);
nor U9654 (N_9654,N_9465,N_9406);
nor U9655 (N_9655,N_9421,N_9384);
nand U9656 (N_9656,N_9523,N_9531);
xor U9657 (N_9657,N_9580,N_9378);
xnor U9658 (N_9658,N_9500,N_9302);
nand U9659 (N_9659,N_9351,N_9355);
or U9660 (N_9660,N_9457,N_9534);
xnor U9661 (N_9661,N_9375,N_9555);
or U9662 (N_9662,N_9448,N_9363);
nand U9663 (N_9663,N_9333,N_9581);
nand U9664 (N_9664,N_9550,N_9595);
and U9665 (N_9665,N_9530,N_9451);
and U9666 (N_9666,N_9571,N_9463);
nor U9667 (N_9667,N_9432,N_9497);
and U9668 (N_9668,N_9494,N_9391);
and U9669 (N_9669,N_9593,N_9389);
xnor U9670 (N_9670,N_9549,N_9343);
or U9671 (N_9671,N_9324,N_9392);
nand U9672 (N_9672,N_9419,N_9430);
xor U9673 (N_9673,N_9536,N_9381);
and U9674 (N_9674,N_9393,N_9372);
and U9675 (N_9675,N_9347,N_9466);
xor U9676 (N_9676,N_9559,N_9379);
xnor U9677 (N_9677,N_9481,N_9556);
nand U9678 (N_9678,N_9462,N_9553);
or U9679 (N_9679,N_9439,N_9441);
nor U9680 (N_9680,N_9413,N_9306);
nand U9681 (N_9681,N_9554,N_9386);
nand U9682 (N_9682,N_9492,N_9402);
or U9683 (N_9683,N_9598,N_9321);
nand U9684 (N_9684,N_9510,N_9390);
nand U9685 (N_9685,N_9359,N_9397);
and U9686 (N_9686,N_9334,N_9354);
nand U9687 (N_9687,N_9428,N_9407);
nor U9688 (N_9688,N_9572,N_9368);
or U9689 (N_9689,N_9410,N_9475);
nor U9690 (N_9690,N_9367,N_9472);
nand U9691 (N_9691,N_9548,N_9398);
xor U9692 (N_9692,N_9551,N_9331);
xnor U9693 (N_9693,N_9327,N_9361);
nand U9694 (N_9694,N_9471,N_9440);
and U9695 (N_9695,N_9541,N_9544);
xnor U9696 (N_9696,N_9338,N_9540);
nand U9697 (N_9697,N_9433,N_9313);
nor U9698 (N_9698,N_9473,N_9341);
nor U9699 (N_9699,N_9562,N_9529);
or U9700 (N_9700,N_9431,N_9345);
nor U9701 (N_9701,N_9435,N_9339);
and U9702 (N_9702,N_9415,N_9325);
nand U9703 (N_9703,N_9467,N_9373);
xor U9704 (N_9704,N_9585,N_9458);
nor U9705 (N_9705,N_9519,N_9516);
xor U9706 (N_9706,N_9332,N_9315);
nand U9707 (N_9707,N_9438,N_9587);
nor U9708 (N_9708,N_9517,N_9444);
or U9709 (N_9709,N_9596,N_9353);
and U9710 (N_9710,N_9486,N_9564);
nor U9711 (N_9711,N_9586,N_9340);
xor U9712 (N_9712,N_9535,N_9312);
or U9713 (N_9713,N_9450,N_9394);
nor U9714 (N_9714,N_9577,N_9464);
or U9715 (N_9715,N_9349,N_9396);
or U9716 (N_9716,N_9401,N_9330);
nor U9717 (N_9717,N_9403,N_9505);
xnor U9718 (N_9718,N_9337,N_9414);
or U9719 (N_9719,N_9446,N_9502);
xor U9720 (N_9720,N_9573,N_9328);
xor U9721 (N_9721,N_9358,N_9320);
or U9722 (N_9722,N_9360,N_9303);
nor U9723 (N_9723,N_9557,N_9489);
or U9724 (N_9724,N_9322,N_9380);
or U9725 (N_9725,N_9491,N_9582);
nand U9726 (N_9726,N_9356,N_9570);
and U9727 (N_9727,N_9496,N_9357);
or U9728 (N_9728,N_9399,N_9563);
nand U9729 (N_9729,N_9528,N_9522);
nor U9730 (N_9730,N_9409,N_9569);
xnor U9731 (N_9731,N_9405,N_9512);
nor U9732 (N_9732,N_9527,N_9310);
nand U9733 (N_9733,N_9420,N_9346);
nor U9734 (N_9734,N_9547,N_9374);
xor U9735 (N_9735,N_9470,N_9449);
and U9736 (N_9736,N_9537,N_9326);
nor U9737 (N_9737,N_9591,N_9579);
nand U9738 (N_9738,N_9437,N_9365);
and U9739 (N_9739,N_9382,N_9411);
nand U9740 (N_9740,N_9488,N_9584);
nand U9741 (N_9741,N_9460,N_9495);
and U9742 (N_9742,N_9452,N_9485);
nand U9743 (N_9743,N_9474,N_9400);
nor U9744 (N_9744,N_9543,N_9493);
and U9745 (N_9745,N_9434,N_9498);
or U9746 (N_9746,N_9469,N_9408);
xnor U9747 (N_9747,N_9490,N_9369);
nor U9748 (N_9748,N_9590,N_9424);
and U9749 (N_9749,N_9404,N_9588);
and U9750 (N_9750,N_9315,N_9492);
and U9751 (N_9751,N_9315,N_9537);
or U9752 (N_9752,N_9444,N_9407);
xnor U9753 (N_9753,N_9334,N_9391);
or U9754 (N_9754,N_9356,N_9530);
xor U9755 (N_9755,N_9578,N_9571);
xor U9756 (N_9756,N_9326,N_9504);
nor U9757 (N_9757,N_9596,N_9411);
nor U9758 (N_9758,N_9365,N_9591);
xor U9759 (N_9759,N_9532,N_9548);
nand U9760 (N_9760,N_9586,N_9418);
nor U9761 (N_9761,N_9572,N_9556);
and U9762 (N_9762,N_9513,N_9478);
nor U9763 (N_9763,N_9505,N_9512);
or U9764 (N_9764,N_9322,N_9533);
nor U9765 (N_9765,N_9500,N_9513);
and U9766 (N_9766,N_9413,N_9415);
nand U9767 (N_9767,N_9463,N_9407);
and U9768 (N_9768,N_9378,N_9415);
xor U9769 (N_9769,N_9582,N_9556);
nand U9770 (N_9770,N_9585,N_9347);
nor U9771 (N_9771,N_9514,N_9521);
and U9772 (N_9772,N_9553,N_9435);
and U9773 (N_9773,N_9519,N_9456);
nor U9774 (N_9774,N_9363,N_9372);
or U9775 (N_9775,N_9321,N_9564);
nor U9776 (N_9776,N_9381,N_9583);
xor U9777 (N_9777,N_9357,N_9465);
nand U9778 (N_9778,N_9411,N_9444);
xor U9779 (N_9779,N_9367,N_9400);
nand U9780 (N_9780,N_9554,N_9517);
and U9781 (N_9781,N_9432,N_9347);
nand U9782 (N_9782,N_9497,N_9317);
nor U9783 (N_9783,N_9496,N_9464);
xnor U9784 (N_9784,N_9563,N_9342);
nor U9785 (N_9785,N_9585,N_9571);
xnor U9786 (N_9786,N_9537,N_9581);
nor U9787 (N_9787,N_9379,N_9525);
xnor U9788 (N_9788,N_9460,N_9549);
xor U9789 (N_9789,N_9356,N_9350);
and U9790 (N_9790,N_9352,N_9541);
or U9791 (N_9791,N_9555,N_9513);
and U9792 (N_9792,N_9504,N_9543);
nand U9793 (N_9793,N_9400,N_9439);
xor U9794 (N_9794,N_9444,N_9386);
or U9795 (N_9795,N_9314,N_9560);
nand U9796 (N_9796,N_9427,N_9352);
and U9797 (N_9797,N_9410,N_9547);
nand U9798 (N_9798,N_9437,N_9302);
nor U9799 (N_9799,N_9328,N_9559);
xor U9800 (N_9800,N_9412,N_9342);
nor U9801 (N_9801,N_9407,N_9561);
nor U9802 (N_9802,N_9326,N_9533);
and U9803 (N_9803,N_9422,N_9328);
and U9804 (N_9804,N_9408,N_9549);
and U9805 (N_9805,N_9346,N_9560);
nand U9806 (N_9806,N_9332,N_9511);
xor U9807 (N_9807,N_9314,N_9340);
and U9808 (N_9808,N_9323,N_9404);
nor U9809 (N_9809,N_9449,N_9383);
nor U9810 (N_9810,N_9509,N_9356);
xnor U9811 (N_9811,N_9553,N_9582);
and U9812 (N_9812,N_9433,N_9315);
and U9813 (N_9813,N_9526,N_9553);
and U9814 (N_9814,N_9329,N_9325);
or U9815 (N_9815,N_9543,N_9352);
or U9816 (N_9816,N_9306,N_9420);
or U9817 (N_9817,N_9506,N_9373);
nor U9818 (N_9818,N_9513,N_9300);
or U9819 (N_9819,N_9366,N_9304);
nor U9820 (N_9820,N_9393,N_9324);
and U9821 (N_9821,N_9580,N_9478);
or U9822 (N_9822,N_9332,N_9525);
and U9823 (N_9823,N_9568,N_9575);
nor U9824 (N_9824,N_9359,N_9461);
xor U9825 (N_9825,N_9578,N_9414);
xor U9826 (N_9826,N_9365,N_9521);
nor U9827 (N_9827,N_9490,N_9435);
nand U9828 (N_9828,N_9373,N_9470);
nand U9829 (N_9829,N_9562,N_9436);
nor U9830 (N_9830,N_9591,N_9484);
or U9831 (N_9831,N_9368,N_9481);
nor U9832 (N_9832,N_9592,N_9339);
or U9833 (N_9833,N_9495,N_9361);
xnor U9834 (N_9834,N_9403,N_9561);
and U9835 (N_9835,N_9463,N_9553);
and U9836 (N_9836,N_9379,N_9534);
nand U9837 (N_9837,N_9419,N_9580);
or U9838 (N_9838,N_9388,N_9431);
and U9839 (N_9839,N_9464,N_9428);
nor U9840 (N_9840,N_9564,N_9365);
or U9841 (N_9841,N_9324,N_9540);
and U9842 (N_9842,N_9398,N_9359);
xnor U9843 (N_9843,N_9428,N_9438);
or U9844 (N_9844,N_9565,N_9420);
xor U9845 (N_9845,N_9583,N_9476);
xnor U9846 (N_9846,N_9575,N_9567);
or U9847 (N_9847,N_9410,N_9416);
xnor U9848 (N_9848,N_9599,N_9481);
nor U9849 (N_9849,N_9488,N_9314);
nand U9850 (N_9850,N_9546,N_9599);
xor U9851 (N_9851,N_9554,N_9595);
xnor U9852 (N_9852,N_9438,N_9522);
xor U9853 (N_9853,N_9463,N_9539);
and U9854 (N_9854,N_9315,N_9552);
xnor U9855 (N_9855,N_9382,N_9568);
nor U9856 (N_9856,N_9362,N_9442);
xnor U9857 (N_9857,N_9302,N_9546);
or U9858 (N_9858,N_9565,N_9407);
nand U9859 (N_9859,N_9332,N_9336);
and U9860 (N_9860,N_9333,N_9496);
nand U9861 (N_9861,N_9390,N_9366);
nand U9862 (N_9862,N_9393,N_9379);
or U9863 (N_9863,N_9413,N_9420);
or U9864 (N_9864,N_9462,N_9444);
or U9865 (N_9865,N_9425,N_9456);
or U9866 (N_9866,N_9558,N_9408);
or U9867 (N_9867,N_9466,N_9437);
xnor U9868 (N_9868,N_9512,N_9500);
and U9869 (N_9869,N_9324,N_9488);
xnor U9870 (N_9870,N_9325,N_9333);
nand U9871 (N_9871,N_9549,N_9428);
xnor U9872 (N_9872,N_9550,N_9379);
nor U9873 (N_9873,N_9527,N_9526);
nor U9874 (N_9874,N_9526,N_9379);
nand U9875 (N_9875,N_9360,N_9570);
and U9876 (N_9876,N_9330,N_9425);
and U9877 (N_9877,N_9536,N_9312);
nand U9878 (N_9878,N_9539,N_9501);
nand U9879 (N_9879,N_9422,N_9510);
xor U9880 (N_9880,N_9500,N_9301);
or U9881 (N_9881,N_9375,N_9440);
xnor U9882 (N_9882,N_9317,N_9440);
nor U9883 (N_9883,N_9575,N_9403);
nand U9884 (N_9884,N_9599,N_9342);
or U9885 (N_9885,N_9493,N_9396);
nor U9886 (N_9886,N_9440,N_9447);
xor U9887 (N_9887,N_9441,N_9313);
nor U9888 (N_9888,N_9330,N_9421);
nor U9889 (N_9889,N_9301,N_9597);
nand U9890 (N_9890,N_9408,N_9533);
xnor U9891 (N_9891,N_9342,N_9329);
and U9892 (N_9892,N_9576,N_9305);
or U9893 (N_9893,N_9389,N_9379);
nand U9894 (N_9894,N_9428,N_9490);
nand U9895 (N_9895,N_9431,N_9362);
nand U9896 (N_9896,N_9435,N_9485);
nor U9897 (N_9897,N_9390,N_9455);
xnor U9898 (N_9898,N_9531,N_9482);
nand U9899 (N_9899,N_9560,N_9476);
xnor U9900 (N_9900,N_9613,N_9825);
and U9901 (N_9901,N_9889,N_9620);
nand U9902 (N_9902,N_9644,N_9899);
nor U9903 (N_9903,N_9891,N_9831);
xor U9904 (N_9904,N_9788,N_9654);
and U9905 (N_9905,N_9679,N_9822);
and U9906 (N_9906,N_9854,N_9705);
nor U9907 (N_9907,N_9779,N_9638);
nor U9908 (N_9908,N_9643,N_9751);
xor U9909 (N_9909,N_9699,N_9816);
xnor U9910 (N_9910,N_9856,N_9604);
or U9911 (N_9911,N_9782,N_9748);
xor U9912 (N_9912,N_9676,N_9651);
and U9913 (N_9913,N_9871,N_9785);
nor U9914 (N_9914,N_9645,N_9830);
xor U9915 (N_9915,N_9750,N_9778);
or U9916 (N_9916,N_9684,N_9635);
or U9917 (N_9917,N_9708,N_9802);
and U9918 (N_9918,N_9660,N_9797);
and U9919 (N_9919,N_9832,N_9895);
xor U9920 (N_9920,N_9823,N_9617);
or U9921 (N_9921,N_9893,N_9622);
or U9922 (N_9922,N_9861,N_9695);
and U9923 (N_9923,N_9612,N_9636);
and U9924 (N_9924,N_9682,N_9824);
xor U9925 (N_9925,N_9650,N_9809);
xnor U9926 (N_9926,N_9698,N_9719);
nor U9927 (N_9927,N_9611,N_9688);
nor U9928 (N_9928,N_9789,N_9659);
and U9929 (N_9929,N_9729,N_9640);
or U9930 (N_9930,N_9722,N_9641);
and U9931 (N_9931,N_9806,N_9717);
xnor U9932 (N_9932,N_9655,N_9857);
and U9933 (N_9933,N_9671,N_9632);
nand U9934 (N_9934,N_9800,N_9714);
nand U9935 (N_9935,N_9639,N_9852);
nand U9936 (N_9936,N_9828,N_9656);
and U9937 (N_9937,N_9880,N_9775);
or U9938 (N_9938,N_9793,N_9602);
nand U9939 (N_9939,N_9675,N_9850);
and U9940 (N_9940,N_9637,N_9711);
nand U9941 (N_9941,N_9787,N_9710);
or U9942 (N_9942,N_9653,N_9601);
or U9943 (N_9943,N_9606,N_9702);
or U9944 (N_9944,N_9746,N_9736);
and U9945 (N_9945,N_9855,N_9795);
nand U9946 (N_9946,N_9725,N_9847);
and U9947 (N_9947,N_9885,N_9759);
nor U9948 (N_9948,N_9777,N_9649);
and U9949 (N_9949,N_9745,N_9815);
xnor U9950 (N_9950,N_9683,N_9799);
nand U9951 (N_9951,N_9603,N_9737);
nand U9952 (N_9952,N_9624,N_9694);
xnor U9953 (N_9953,N_9890,N_9887);
nand U9954 (N_9954,N_9741,N_9819);
and U9955 (N_9955,N_9860,N_9886);
or U9956 (N_9956,N_9668,N_9662);
nand U9957 (N_9957,N_9680,N_9703);
nand U9958 (N_9958,N_9869,N_9619);
nor U9959 (N_9959,N_9820,N_9652);
nor U9960 (N_9960,N_9833,N_9739);
and U9961 (N_9961,N_9701,N_9721);
or U9962 (N_9962,N_9625,N_9757);
and U9963 (N_9963,N_9672,N_9616);
nor U9964 (N_9964,N_9858,N_9866);
nand U9965 (N_9965,N_9811,N_9600);
and U9966 (N_9966,N_9844,N_9826);
and U9967 (N_9967,N_9813,N_9874);
or U9968 (N_9968,N_9744,N_9692);
nand U9969 (N_9969,N_9877,N_9898);
or U9970 (N_9970,N_9661,N_9609);
and U9971 (N_9971,N_9634,N_9756);
and U9972 (N_9972,N_9827,N_9864);
and U9973 (N_9973,N_9818,N_9839);
xor U9974 (N_9974,N_9881,N_9837);
or U9975 (N_9975,N_9657,N_9642);
and U9976 (N_9976,N_9853,N_9628);
nand U9977 (N_9977,N_9726,N_9631);
xor U9978 (N_9978,N_9753,N_9674);
nand U9979 (N_9979,N_9768,N_9704);
nand U9980 (N_9980,N_9665,N_9770);
or U9981 (N_9981,N_9859,N_9846);
xor U9982 (N_9982,N_9670,N_9673);
xor U9983 (N_9983,N_9687,N_9879);
nor U9984 (N_9984,N_9865,N_9892);
and U9985 (N_9985,N_9614,N_9713);
and U9986 (N_9986,N_9872,N_9786);
or U9987 (N_9987,N_9771,N_9664);
nor U9988 (N_9988,N_9740,N_9766);
xor U9989 (N_9989,N_9834,N_9715);
nor U9990 (N_9990,N_9790,N_9758);
or U9991 (N_9991,N_9730,N_9734);
nor U9992 (N_9992,N_9618,N_9761);
nor U9993 (N_9993,N_9621,N_9772);
nor U9994 (N_9994,N_9851,N_9685);
xor U9995 (N_9995,N_9728,N_9623);
nand U9996 (N_9996,N_9848,N_9629);
or U9997 (N_9997,N_9798,N_9700);
or U9998 (N_9998,N_9681,N_9842);
or U9999 (N_9999,N_9838,N_9610);
nor U10000 (N_10000,N_9720,N_9735);
nor U10001 (N_10001,N_9817,N_9810);
nor U10002 (N_10002,N_9882,N_9884);
or U10003 (N_10003,N_9696,N_9663);
nor U10004 (N_10004,N_9707,N_9731);
xnor U10005 (N_10005,N_9808,N_9686);
nand U10006 (N_10006,N_9780,N_9845);
and U10007 (N_10007,N_9883,N_9697);
nor U10008 (N_10008,N_9862,N_9646);
nor U10009 (N_10009,N_9607,N_9615);
xor U10010 (N_10010,N_9723,N_9767);
nand U10011 (N_10011,N_9803,N_9841);
xor U10012 (N_10012,N_9706,N_9773);
xnor U10013 (N_10013,N_9693,N_9829);
nor U10014 (N_10014,N_9749,N_9863);
xor U10015 (N_10015,N_9801,N_9689);
or U10016 (N_10016,N_9763,N_9807);
xnor U10017 (N_10017,N_9765,N_9605);
or U10018 (N_10018,N_9796,N_9804);
and U10019 (N_10019,N_9691,N_9752);
or U10020 (N_10020,N_9849,N_9888);
nor U10021 (N_10021,N_9783,N_9876);
xor U10022 (N_10022,N_9727,N_9627);
nor U10023 (N_10023,N_9781,N_9626);
nand U10024 (N_10024,N_9738,N_9769);
nand U10025 (N_10025,N_9836,N_9667);
or U10026 (N_10026,N_9677,N_9678);
nand U10027 (N_10027,N_9608,N_9762);
or U10028 (N_10028,N_9754,N_9760);
nand U10029 (N_10029,N_9633,N_9718);
xnor U10030 (N_10030,N_9742,N_9878);
nand U10031 (N_10031,N_9896,N_9868);
or U10032 (N_10032,N_9658,N_9709);
or U10033 (N_10033,N_9894,N_9690);
xor U10034 (N_10034,N_9774,N_9755);
xor U10035 (N_10035,N_9764,N_9835);
and U10036 (N_10036,N_9743,N_9732);
or U10037 (N_10037,N_9814,N_9843);
or U10038 (N_10038,N_9776,N_9821);
nor U10039 (N_10039,N_9630,N_9784);
or U10040 (N_10040,N_9812,N_9724);
xor U10041 (N_10041,N_9897,N_9648);
nor U10042 (N_10042,N_9733,N_9747);
nand U10043 (N_10043,N_9805,N_9712);
nand U10044 (N_10044,N_9647,N_9867);
or U10045 (N_10045,N_9791,N_9875);
nor U10046 (N_10046,N_9873,N_9870);
nor U10047 (N_10047,N_9716,N_9669);
nand U10048 (N_10048,N_9666,N_9794);
or U10049 (N_10049,N_9840,N_9792);
nor U10050 (N_10050,N_9788,N_9655);
or U10051 (N_10051,N_9738,N_9893);
nor U10052 (N_10052,N_9829,N_9865);
and U10053 (N_10053,N_9666,N_9806);
nand U10054 (N_10054,N_9766,N_9833);
and U10055 (N_10055,N_9786,N_9627);
and U10056 (N_10056,N_9643,N_9702);
or U10057 (N_10057,N_9716,N_9881);
xor U10058 (N_10058,N_9749,N_9631);
xnor U10059 (N_10059,N_9657,N_9655);
xor U10060 (N_10060,N_9810,N_9653);
and U10061 (N_10061,N_9722,N_9757);
nand U10062 (N_10062,N_9895,N_9867);
or U10063 (N_10063,N_9624,N_9770);
nand U10064 (N_10064,N_9656,N_9829);
xnor U10065 (N_10065,N_9709,N_9855);
xor U10066 (N_10066,N_9671,N_9674);
nor U10067 (N_10067,N_9854,N_9636);
or U10068 (N_10068,N_9836,N_9705);
or U10069 (N_10069,N_9600,N_9751);
or U10070 (N_10070,N_9687,N_9855);
nand U10071 (N_10071,N_9843,N_9879);
xnor U10072 (N_10072,N_9755,N_9819);
xnor U10073 (N_10073,N_9783,N_9666);
nand U10074 (N_10074,N_9751,N_9631);
nand U10075 (N_10075,N_9673,N_9629);
and U10076 (N_10076,N_9876,N_9853);
nand U10077 (N_10077,N_9774,N_9634);
or U10078 (N_10078,N_9790,N_9895);
nor U10079 (N_10079,N_9830,N_9703);
or U10080 (N_10080,N_9882,N_9691);
nor U10081 (N_10081,N_9801,N_9659);
nor U10082 (N_10082,N_9854,N_9658);
or U10083 (N_10083,N_9690,N_9887);
nand U10084 (N_10084,N_9617,N_9838);
nand U10085 (N_10085,N_9709,N_9711);
nand U10086 (N_10086,N_9852,N_9615);
xnor U10087 (N_10087,N_9674,N_9740);
and U10088 (N_10088,N_9625,N_9784);
or U10089 (N_10089,N_9665,N_9610);
and U10090 (N_10090,N_9743,N_9758);
or U10091 (N_10091,N_9667,N_9818);
xnor U10092 (N_10092,N_9781,N_9751);
nand U10093 (N_10093,N_9853,N_9600);
xor U10094 (N_10094,N_9846,N_9685);
or U10095 (N_10095,N_9771,N_9623);
nor U10096 (N_10096,N_9718,N_9634);
xor U10097 (N_10097,N_9888,N_9698);
nand U10098 (N_10098,N_9660,N_9711);
or U10099 (N_10099,N_9716,N_9785);
nand U10100 (N_10100,N_9891,N_9897);
nand U10101 (N_10101,N_9695,N_9678);
xor U10102 (N_10102,N_9722,N_9622);
nand U10103 (N_10103,N_9615,N_9624);
or U10104 (N_10104,N_9861,N_9625);
nor U10105 (N_10105,N_9794,N_9833);
nor U10106 (N_10106,N_9637,N_9676);
or U10107 (N_10107,N_9643,N_9864);
or U10108 (N_10108,N_9809,N_9832);
or U10109 (N_10109,N_9635,N_9648);
and U10110 (N_10110,N_9696,N_9788);
or U10111 (N_10111,N_9828,N_9771);
or U10112 (N_10112,N_9658,N_9861);
nand U10113 (N_10113,N_9845,N_9798);
nand U10114 (N_10114,N_9655,N_9634);
nand U10115 (N_10115,N_9635,N_9791);
and U10116 (N_10116,N_9876,N_9823);
and U10117 (N_10117,N_9823,N_9664);
nand U10118 (N_10118,N_9670,N_9617);
or U10119 (N_10119,N_9604,N_9828);
nand U10120 (N_10120,N_9804,N_9743);
xnor U10121 (N_10121,N_9630,N_9840);
nand U10122 (N_10122,N_9757,N_9715);
nor U10123 (N_10123,N_9682,N_9607);
or U10124 (N_10124,N_9863,N_9607);
nand U10125 (N_10125,N_9635,N_9717);
nand U10126 (N_10126,N_9755,N_9853);
nor U10127 (N_10127,N_9788,N_9857);
nor U10128 (N_10128,N_9644,N_9826);
xnor U10129 (N_10129,N_9645,N_9793);
xnor U10130 (N_10130,N_9704,N_9835);
xnor U10131 (N_10131,N_9757,N_9686);
xor U10132 (N_10132,N_9831,N_9716);
or U10133 (N_10133,N_9601,N_9648);
nand U10134 (N_10134,N_9768,N_9707);
xnor U10135 (N_10135,N_9766,N_9741);
or U10136 (N_10136,N_9844,N_9741);
nor U10137 (N_10137,N_9746,N_9801);
and U10138 (N_10138,N_9631,N_9759);
nor U10139 (N_10139,N_9707,N_9711);
xnor U10140 (N_10140,N_9768,N_9897);
or U10141 (N_10141,N_9854,N_9778);
or U10142 (N_10142,N_9780,N_9681);
xor U10143 (N_10143,N_9616,N_9695);
xnor U10144 (N_10144,N_9706,N_9607);
and U10145 (N_10145,N_9690,N_9750);
nor U10146 (N_10146,N_9618,N_9665);
xor U10147 (N_10147,N_9863,N_9729);
nand U10148 (N_10148,N_9736,N_9726);
nor U10149 (N_10149,N_9619,N_9657);
xor U10150 (N_10150,N_9614,N_9679);
nand U10151 (N_10151,N_9802,N_9678);
xnor U10152 (N_10152,N_9770,N_9757);
and U10153 (N_10153,N_9842,N_9665);
and U10154 (N_10154,N_9788,N_9626);
nand U10155 (N_10155,N_9891,N_9797);
xor U10156 (N_10156,N_9607,N_9610);
and U10157 (N_10157,N_9775,N_9861);
nand U10158 (N_10158,N_9874,N_9808);
nand U10159 (N_10159,N_9854,N_9830);
and U10160 (N_10160,N_9788,N_9728);
nor U10161 (N_10161,N_9626,N_9848);
or U10162 (N_10162,N_9708,N_9862);
and U10163 (N_10163,N_9619,N_9715);
xnor U10164 (N_10164,N_9802,N_9628);
nor U10165 (N_10165,N_9685,N_9878);
or U10166 (N_10166,N_9662,N_9709);
nand U10167 (N_10167,N_9895,N_9626);
nand U10168 (N_10168,N_9866,N_9763);
xnor U10169 (N_10169,N_9652,N_9842);
or U10170 (N_10170,N_9701,N_9806);
xor U10171 (N_10171,N_9888,N_9731);
nand U10172 (N_10172,N_9762,N_9869);
xnor U10173 (N_10173,N_9779,N_9716);
nand U10174 (N_10174,N_9721,N_9689);
or U10175 (N_10175,N_9818,N_9640);
nor U10176 (N_10176,N_9625,N_9858);
and U10177 (N_10177,N_9753,N_9803);
xor U10178 (N_10178,N_9615,N_9640);
nand U10179 (N_10179,N_9682,N_9671);
nand U10180 (N_10180,N_9799,N_9876);
xor U10181 (N_10181,N_9604,N_9602);
xor U10182 (N_10182,N_9784,N_9659);
nand U10183 (N_10183,N_9883,N_9738);
nand U10184 (N_10184,N_9782,N_9881);
and U10185 (N_10185,N_9711,N_9810);
and U10186 (N_10186,N_9749,N_9657);
nor U10187 (N_10187,N_9713,N_9843);
xor U10188 (N_10188,N_9853,N_9736);
xor U10189 (N_10189,N_9711,N_9684);
xnor U10190 (N_10190,N_9683,N_9654);
nand U10191 (N_10191,N_9607,N_9668);
and U10192 (N_10192,N_9874,N_9730);
nand U10193 (N_10193,N_9801,N_9705);
nand U10194 (N_10194,N_9807,N_9869);
nor U10195 (N_10195,N_9701,N_9707);
nor U10196 (N_10196,N_9752,N_9826);
nor U10197 (N_10197,N_9838,N_9822);
and U10198 (N_10198,N_9614,N_9842);
xor U10199 (N_10199,N_9804,N_9619);
xor U10200 (N_10200,N_9976,N_10144);
xnor U10201 (N_10201,N_10092,N_10093);
and U10202 (N_10202,N_10129,N_10167);
or U10203 (N_10203,N_10185,N_10098);
and U10204 (N_10204,N_9916,N_10004);
or U10205 (N_10205,N_9987,N_9998);
and U10206 (N_10206,N_10070,N_9919);
nand U10207 (N_10207,N_10106,N_9974);
and U10208 (N_10208,N_10044,N_9904);
or U10209 (N_10209,N_10154,N_10149);
nand U10210 (N_10210,N_9951,N_10166);
nand U10211 (N_10211,N_10029,N_10023);
and U10212 (N_10212,N_10010,N_9970);
or U10213 (N_10213,N_10035,N_9901);
nand U10214 (N_10214,N_9906,N_10078);
xor U10215 (N_10215,N_10071,N_10081);
nand U10216 (N_10216,N_10137,N_10189);
xor U10217 (N_10217,N_10155,N_9942);
nand U10218 (N_10218,N_9903,N_10125);
and U10219 (N_10219,N_10158,N_10022);
and U10220 (N_10220,N_9994,N_9940);
xor U10221 (N_10221,N_10183,N_10009);
and U10222 (N_10222,N_9937,N_10053);
nor U10223 (N_10223,N_10136,N_10055);
or U10224 (N_10224,N_9945,N_10096);
xnor U10225 (N_10225,N_9985,N_9996);
nand U10226 (N_10226,N_10019,N_9947);
nor U10227 (N_10227,N_9991,N_10174);
or U10228 (N_10228,N_10073,N_10181);
and U10229 (N_10229,N_9978,N_10140);
nor U10230 (N_10230,N_10057,N_10061);
xor U10231 (N_10231,N_10087,N_10094);
and U10232 (N_10232,N_9953,N_10198);
nand U10233 (N_10233,N_10095,N_9932);
or U10234 (N_10234,N_9988,N_9948);
or U10235 (N_10235,N_10016,N_10134);
xor U10236 (N_10236,N_10188,N_10021);
or U10237 (N_10237,N_10082,N_10164);
nor U10238 (N_10238,N_10039,N_9949);
and U10239 (N_10239,N_10091,N_10162);
nor U10240 (N_10240,N_10005,N_9911);
and U10241 (N_10241,N_10177,N_10182);
and U10242 (N_10242,N_10145,N_10049);
or U10243 (N_10243,N_9924,N_10123);
or U10244 (N_10244,N_10160,N_10028);
xnor U10245 (N_10245,N_10020,N_10064);
xor U10246 (N_10246,N_9923,N_9905);
and U10247 (N_10247,N_9984,N_10088);
and U10248 (N_10248,N_10027,N_10015);
nand U10249 (N_10249,N_10191,N_10157);
nor U10250 (N_10250,N_9900,N_10052);
nand U10251 (N_10251,N_9961,N_9943);
xor U10252 (N_10252,N_10018,N_9902);
and U10253 (N_10253,N_10141,N_10058);
and U10254 (N_10254,N_10068,N_10146);
nor U10255 (N_10255,N_9959,N_10056);
or U10256 (N_10256,N_10006,N_9990);
or U10257 (N_10257,N_9912,N_10197);
xnor U10258 (N_10258,N_10163,N_9989);
nor U10259 (N_10259,N_9980,N_9914);
and U10260 (N_10260,N_10037,N_10178);
nor U10261 (N_10261,N_9986,N_10076);
or U10262 (N_10262,N_10050,N_9913);
nor U10263 (N_10263,N_10063,N_9997);
or U10264 (N_10264,N_10017,N_9921);
and U10265 (N_10265,N_10175,N_9927);
nor U10266 (N_10266,N_10043,N_10024);
nand U10267 (N_10267,N_9983,N_9929);
xnor U10268 (N_10268,N_10047,N_10135);
xor U10269 (N_10269,N_10173,N_10051);
or U10270 (N_10270,N_10194,N_9972);
and U10271 (N_10271,N_9909,N_9995);
or U10272 (N_10272,N_9955,N_10003);
and U10273 (N_10273,N_10090,N_10131);
nand U10274 (N_10274,N_10120,N_10179);
nor U10275 (N_10275,N_10180,N_9939);
nor U10276 (N_10276,N_10169,N_9958);
nand U10277 (N_10277,N_10121,N_9954);
nand U10278 (N_10278,N_9992,N_10109);
and U10279 (N_10279,N_9931,N_10040);
and U10280 (N_10280,N_9999,N_10085);
or U10281 (N_10281,N_9950,N_10042);
nor U10282 (N_10282,N_10030,N_10139);
nand U10283 (N_10283,N_10147,N_9963);
and U10284 (N_10284,N_9946,N_10007);
nor U10285 (N_10285,N_10036,N_10186);
xnor U10286 (N_10286,N_10080,N_9910);
nor U10287 (N_10287,N_10115,N_9982);
or U10288 (N_10288,N_10083,N_10187);
nor U10289 (N_10289,N_9966,N_10195);
or U10290 (N_10290,N_10001,N_10199);
nor U10291 (N_10291,N_10156,N_10034);
xor U10292 (N_10292,N_10045,N_10190);
and U10293 (N_10293,N_9993,N_10152);
and U10294 (N_10294,N_10127,N_10104);
and U10295 (N_10295,N_10110,N_10126);
and U10296 (N_10296,N_10165,N_10105);
or U10297 (N_10297,N_10012,N_9973);
and U10298 (N_10298,N_10072,N_9981);
nor U10299 (N_10299,N_9926,N_10084);
nor U10300 (N_10300,N_10048,N_10128);
nor U10301 (N_10301,N_9920,N_10000);
and U10302 (N_10302,N_9915,N_10008);
nand U10303 (N_10303,N_10114,N_10002);
and U10304 (N_10304,N_10046,N_10193);
and U10305 (N_10305,N_10171,N_9956);
xnor U10306 (N_10306,N_10143,N_9962);
nand U10307 (N_10307,N_10132,N_10079);
and U10308 (N_10308,N_10161,N_10196);
and U10309 (N_10309,N_10159,N_10038);
nor U10310 (N_10310,N_10089,N_10118);
nor U10311 (N_10311,N_10138,N_9941);
and U10312 (N_10312,N_10142,N_10025);
xor U10313 (N_10313,N_10112,N_10086);
nand U10314 (N_10314,N_9908,N_9957);
nor U10315 (N_10315,N_10032,N_9918);
and U10316 (N_10316,N_10184,N_9907);
or U10317 (N_10317,N_10059,N_10133);
nor U10318 (N_10318,N_9975,N_10011);
nor U10319 (N_10319,N_10103,N_10130);
or U10320 (N_10320,N_10116,N_9938);
or U10321 (N_10321,N_10031,N_9934);
nor U10322 (N_10322,N_10170,N_10041);
nand U10323 (N_10323,N_9922,N_10124);
nand U10324 (N_10324,N_9928,N_10102);
nor U10325 (N_10325,N_9964,N_9917);
nor U10326 (N_10326,N_10192,N_10075);
or U10327 (N_10327,N_10099,N_10060);
nor U10328 (N_10328,N_10026,N_10097);
xnor U10329 (N_10329,N_9965,N_10066);
nand U10330 (N_10330,N_10100,N_9960);
nand U10331 (N_10331,N_10113,N_10151);
xnor U10332 (N_10332,N_9935,N_9925);
nand U10333 (N_10333,N_10067,N_10033);
or U10334 (N_10334,N_10054,N_10101);
nor U10335 (N_10335,N_10119,N_10122);
nor U10336 (N_10336,N_10117,N_9952);
and U10337 (N_10337,N_10111,N_9936);
nor U10338 (N_10338,N_10153,N_10107);
xor U10339 (N_10339,N_10014,N_10069);
nor U10340 (N_10340,N_9969,N_10077);
xnor U10341 (N_10341,N_10172,N_10062);
nor U10342 (N_10342,N_9977,N_10065);
or U10343 (N_10343,N_9968,N_9971);
nand U10344 (N_10344,N_10108,N_10150);
or U10345 (N_10345,N_10168,N_9933);
nand U10346 (N_10346,N_10148,N_9944);
xor U10347 (N_10347,N_10074,N_10013);
xor U10348 (N_10348,N_10176,N_9979);
nor U10349 (N_10349,N_9930,N_9967);
and U10350 (N_10350,N_10092,N_9970);
nor U10351 (N_10351,N_9949,N_10191);
nand U10352 (N_10352,N_9911,N_10077);
nand U10353 (N_10353,N_10181,N_10185);
nor U10354 (N_10354,N_9998,N_10013);
and U10355 (N_10355,N_10124,N_10036);
nor U10356 (N_10356,N_9976,N_10193);
nor U10357 (N_10357,N_9990,N_9938);
or U10358 (N_10358,N_10052,N_10119);
nand U10359 (N_10359,N_9958,N_10005);
and U10360 (N_10360,N_10040,N_10174);
xor U10361 (N_10361,N_10027,N_10198);
and U10362 (N_10362,N_10049,N_9935);
or U10363 (N_10363,N_10097,N_10092);
xnor U10364 (N_10364,N_10096,N_9990);
nor U10365 (N_10365,N_10148,N_9990);
and U10366 (N_10366,N_10159,N_9989);
and U10367 (N_10367,N_10161,N_10136);
nor U10368 (N_10368,N_9967,N_10185);
nand U10369 (N_10369,N_10026,N_9912);
nand U10370 (N_10370,N_9964,N_9979);
and U10371 (N_10371,N_10038,N_10095);
nand U10372 (N_10372,N_9928,N_10110);
nand U10373 (N_10373,N_10022,N_10102);
nand U10374 (N_10374,N_10098,N_10187);
nand U10375 (N_10375,N_9999,N_10124);
or U10376 (N_10376,N_10179,N_10055);
nor U10377 (N_10377,N_10154,N_10031);
or U10378 (N_10378,N_9936,N_10114);
nand U10379 (N_10379,N_10199,N_9914);
nand U10380 (N_10380,N_10104,N_9905);
and U10381 (N_10381,N_10055,N_10126);
xor U10382 (N_10382,N_9981,N_10042);
xnor U10383 (N_10383,N_10138,N_10049);
and U10384 (N_10384,N_9911,N_10142);
or U10385 (N_10385,N_10193,N_9950);
and U10386 (N_10386,N_9945,N_10120);
xnor U10387 (N_10387,N_10039,N_10074);
and U10388 (N_10388,N_10087,N_10038);
and U10389 (N_10389,N_10010,N_9996);
or U10390 (N_10390,N_10143,N_9916);
and U10391 (N_10391,N_9994,N_9904);
and U10392 (N_10392,N_10025,N_10116);
or U10393 (N_10393,N_9916,N_10039);
and U10394 (N_10394,N_10192,N_9906);
xor U10395 (N_10395,N_10151,N_10153);
nor U10396 (N_10396,N_10165,N_10015);
and U10397 (N_10397,N_10138,N_10101);
or U10398 (N_10398,N_9984,N_10144);
and U10399 (N_10399,N_9934,N_10143);
or U10400 (N_10400,N_10155,N_10097);
and U10401 (N_10401,N_10104,N_10173);
or U10402 (N_10402,N_10017,N_9995);
or U10403 (N_10403,N_10149,N_9909);
nand U10404 (N_10404,N_10197,N_9918);
nand U10405 (N_10405,N_10161,N_10090);
xor U10406 (N_10406,N_10136,N_9938);
nor U10407 (N_10407,N_10004,N_10026);
xnor U10408 (N_10408,N_9958,N_10058);
nor U10409 (N_10409,N_10106,N_10018);
and U10410 (N_10410,N_10173,N_10176);
xor U10411 (N_10411,N_10160,N_10031);
nand U10412 (N_10412,N_10131,N_10024);
or U10413 (N_10413,N_10100,N_10026);
nor U10414 (N_10414,N_10023,N_10107);
xnor U10415 (N_10415,N_9900,N_10078);
xor U10416 (N_10416,N_10010,N_10150);
or U10417 (N_10417,N_10145,N_9951);
nor U10418 (N_10418,N_10163,N_10083);
nand U10419 (N_10419,N_9962,N_10005);
or U10420 (N_10420,N_9956,N_10155);
nor U10421 (N_10421,N_10139,N_10167);
or U10422 (N_10422,N_10180,N_9902);
or U10423 (N_10423,N_10165,N_10181);
and U10424 (N_10424,N_10063,N_9931);
nor U10425 (N_10425,N_9942,N_10191);
nand U10426 (N_10426,N_10084,N_9971);
nand U10427 (N_10427,N_10090,N_9905);
and U10428 (N_10428,N_10129,N_10138);
xnor U10429 (N_10429,N_9974,N_10167);
nand U10430 (N_10430,N_10150,N_9986);
and U10431 (N_10431,N_10033,N_9964);
nand U10432 (N_10432,N_10036,N_10165);
or U10433 (N_10433,N_9920,N_9984);
xnor U10434 (N_10434,N_10030,N_10171);
nand U10435 (N_10435,N_9913,N_9960);
nor U10436 (N_10436,N_10021,N_9912);
nand U10437 (N_10437,N_10052,N_10185);
nor U10438 (N_10438,N_9943,N_9963);
xor U10439 (N_10439,N_9968,N_10131);
and U10440 (N_10440,N_9917,N_9923);
xor U10441 (N_10441,N_9960,N_10002);
nor U10442 (N_10442,N_10093,N_9987);
nor U10443 (N_10443,N_10025,N_10067);
and U10444 (N_10444,N_10151,N_10168);
nor U10445 (N_10445,N_10170,N_9938);
nor U10446 (N_10446,N_10151,N_9980);
nand U10447 (N_10447,N_10109,N_10124);
or U10448 (N_10448,N_10071,N_10182);
and U10449 (N_10449,N_9935,N_10043);
nor U10450 (N_10450,N_9957,N_9974);
nor U10451 (N_10451,N_10119,N_10039);
nand U10452 (N_10452,N_9936,N_10020);
and U10453 (N_10453,N_9997,N_9998);
or U10454 (N_10454,N_10039,N_10108);
nor U10455 (N_10455,N_9977,N_10150);
or U10456 (N_10456,N_10087,N_10126);
and U10457 (N_10457,N_9945,N_10038);
xor U10458 (N_10458,N_10163,N_9949);
or U10459 (N_10459,N_10199,N_10033);
or U10460 (N_10460,N_10173,N_10006);
and U10461 (N_10461,N_10082,N_10163);
xnor U10462 (N_10462,N_9990,N_9947);
nor U10463 (N_10463,N_10198,N_9968);
nand U10464 (N_10464,N_10147,N_10127);
or U10465 (N_10465,N_9919,N_10166);
nand U10466 (N_10466,N_10065,N_10069);
xnor U10467 (N_10467,N_10165,N_10188);
nor U10468 (N_10468,N_10075,N_9909);
xor U10469 (N_10469,N_10028,N_9961);
nand U10470 (N_10470,N_10132,N_9977);
nor U10471 (N_10471,N_10125,N_10002);
or U10472 (N_10472,N_9935,N_9987);
or U10473 (N_10473,N_10084,N_10154);
or U10474 (N_10474,N_10011,N_10154);
and U10475 (N_10475,N_10146,N_10091);
nor U10476 (N_10476,N_10016,N_9929);
or U10477 (N_10477,N_9934,N_10140);
or U10478 (N_10478,N_9945,N_9996);
nor U10479 (N_10479,N_10127,N_10051);
or U10480 (N_10480,N_9922,N_10159);
or U10481 (N_10481,N_9918,N_10069);
xnor U10482 (N_10482,N_10084,N_10095);
and U10483 (N_10483,N_10042,N_9998);
or U10484 (N_10484,N_10110,N_10191);
nand U10485 (N_10485,N_10070,N_10169);
and U10486 (N_10486,N_10183,N_9959);
nand U10487 (N_10487,N_10066,N_10040);
nand U10488 (N_10488,N_10179,N_9924);
nor U10489 (N_10489,N_10049,N_9987);
nor U10490 (N_10490,N_9968,N_10054);
xnor U10491 (N_10491,N_10086,N_10032);
and U10492 (N_10492,N_9939,N_9924);
or U10493 (N_10493,N_9979,N_10028);
or U10494 (N_10494,N_9991,N_10168);
xnor U10495 (N_10495,N_10005,N_9906);
xnor U10496 (N_10496,N_10074,N_10093);
or U10497 (N_10497,N_9954,N_10119);
nand U10498 (N_10498,N_10029,N_9973);
nand U10499 (N_10499,N_10081,N_10150);
and U10500 (N_10500,N_10322,N_10372);
nor U10501 (N_10501,N_10351,N_10496);
and U10502 (N_10502,N_10200,N_10359);
nand U10503 (N_10503,N_10212,N_10380);
nand U10504 (N_10504,N_10203,N_10464);
nor U10505 (N_10505,N_10442,N_10488);
nand U10506 (N_10506,N_10354,N_10264);
and U10507 (N_10507,N_10345,N_10392);
or U10508 (N_10508,N_10315,N_10455);
xnor U10509 (N_10509,N_10469,N_10438);
xnor U10510 (N_10510,N_10422,N_10299);
xnor U10511 (N_10511,N_10478,N_10445);
and U10512 (N_10512,N_10314,N_10361);
and U10513 (N_10513,N_10435,N_10397);
or U10514 (N_10514,N_10470,N_10326);
nand U10515 (N_10515,N_10337,N_10495);
and U10516 (N_10516,N_10208,N_10403);
or U10517 (N_10517,N_10382,N_10207);
and U10518 (N_10518,N_10268,N_10350);
or U10519 (N_10519,N_10233,N_10221);
nand U10520 (N_10520,N_10320,N_10325);
or U10521 (N_10521,N_10269,N_10405);
or U10522 (N_10522,N_10311,N_10241);
xor U10523 (N_10523,N_10352,N_10296);
nor U10524 (N_10524,N_10390,N_10305);
xor U10525 (N_10525,N_10290,N_10228);
nor U10526 (N_10526,N_10347,N_10301);
nand U10527 (N_10527,N_10260,N_10249);
or U10528 (N_10528,N_10238,N_10224);
nand U10529 (N_10529,N_10338,N_10419);
xnor U10530 (N_10530,N_10294,N_10246);
nor U10531 (N_10531,N_10291,N_10493);
nand U10532 (N_10532,N_10202,N_10379);
and U10533 (N_10533,N_10467,N_10358);
or U10534 (N_10534,N_10420,N_10417);
xor U10535 (N_10535,N_10414,N_10477);
xnor U10536 (N_10536,N_10210,N_10211);
nand U10537 (N_10537,N_10370,N_10277);
xor U10538 (N_10538,N_10329,N_10432);
nand U10539 (N_10539,N_10279,N_10218);
and U10540 (N_10540,N_10385,N_10313);
and U10541 (N_10541,N_10446,N_10273);
and U10542 (N_10542,N_10402,N_10250);
or U10543 (N_10543,N_10215,N_10276);
and U10544 (N_10544,N_10307,N_10460);
nor U10545 (N_10545,N_10374,N_10349);
xnor U10546 (N_10546,N_10317,N_10484);
nand U10547 (N_10547,N_10466,N_10366);
nor U10548 (N_10548,N_10365,N_10209);
nand U10549 (N_10549,N_10258,N_10275);
nor U10550 (N_10550,N_10281,N_10408);
and U10551 (N_10551,N_10312,N_10286);
nand U10552 (N_10552,N_10458,N_10214);
nor U10553 (N_10553,N_10259,N_10426);
nor U10554 (N_10554,N_10447,N_10453);
or U10555 (N_10555,N_10243,N_10318);
or U10556 (N_10556,N_10292,N_10398);
nor U10557 (N_10557,N_10356,N_10284);
xnor U10558 (N_10558,N_10425,N_10295);
and U10559 (N_10559,N_10232,N_10413);
xnor U10560 (N_10560,N_10396,N_10375);
or U10561 (N_10561,N_10234,N_10239);
xor U10562 (N_10562,N_10491,N_10404);
nand U10563 (N_10563,N_10452,N_10482);
and U10564 (N_10564,N_10334,N_10483);
nor U10565 (N_10565,N_10437,N_10407);
nand U10566 (N_10566,N_10383,N_10450);
nand U10567 (N_10567,N_10457,N_10297);
or U10568 (N_10568,N_10499,N_10306);
nor U10569 (N_10569,N_10401,N_10223);
and U10570 (N_10570,N_10216,N_10267);
nor U10571 (N_10571,N_10471,N_10377);
nor U10572 (N_10572,N_10309,N_10368);
nor U10573 (N_10573,N_10409,N_10436);
and U10574 (N_10574,N_10247,N_10391);
xor U10575 (N_10575,N_10384,N_10415);
nor U10576 (N_10576,N_10308,N_10360);
nor U10577 (N_10577,N_10271,N_10348);
xnor U10578 (N_10578,N_10448,N_10245);
or U10579 (N_10579,N_10327,N_10490);
nand U10580 (N_10580,N_10480,N_10244);
or U10581 (N_10581,N_10310,N_10463);
nand U10582 (N_10582,N_10400,N_10346);
nor U10583 (N_10583,N_10430,N_10266);
and U10584 (N_10584,N_10433,N_10353);
nor U10585 (N_10585,N_10248,N_10459);
nand U10586 (N_10586,N_10231,N_10222);
or U10587 (N_10587,N_10412,N_10220);
and U10588 (N_10588,N_10381,N_10479);
nor U10589 (N_10589,N_10323,N_10237);
nor U10590 (N_10590,N_10336,N_10240);
or U10591 (N_10591,N_10369,N_10304);
or U10592 (N_10592,N_10461,N_10319);
xor U10593 (N_10593,N_10363,N_10283);
nor U10594 (N_10594,N_10321,N_10387);
or U10595 (N_10595,N_10300,N_10205);
and U10596 (N_10596,N_10395,N_10230);
nor U10597 (N_10597,N_10406,N_10252);
nand U10598 (N_10598,N_10262,N_10474);
xnor U10599 (N_10599,N_10439,N_10465);
and U10600 (N_10600,N_10217,N_10242);
or U10601 (N_10601,N_10434,N_10272);
nand U10602 (N_10602,N_10399,N_10204);
or U10603 (N_10603,N_10206,N_10421);
and U10604 (N_10604,N_10378,N_10293);
nor U10605 (N_10605,N_10362,N_10364);
nor U10606 (N_10606,N_10298,N_10394);
or U10607 (N_10607,N_10226,N_10344);
or U10608 (N_10608,N_10454,N_10257);
xnor U10609 (N_10609,N_10481,N_10441);
and U10610 (N_10610,N_10303,N_10431);
and U10611 (N_10611,N_10373,N_10340);
nor U10612 (N_10612,N_10330,N_10254);
or U10613 (N_10613,N_10324,N_10339);
or U10614 (N_10614,N_10333,N_10411);
xor U10615 (N_10615,N_10468,N_10427);
nor U10616 (N_10616,N_10393,N_10274);
and U10617 (N_10617,N_10487,N_10440);
and U10618 (N_10618,N_10255,N_10416);
or U10619 (N_10619,N_10201,N_10475);
xnor U10620 (N_10620,N_10219,N_10270);
xnor U10621 (N_10621,N_10443,N_10355);
nor U10622 (N_10622,N_10251,N_10449);
or U10623 (N_10623,N_10476,N_10424);
and U10624 (N_10624,N_10444,N_10489);
and U10625 (N_10625,N_10376,N_10388);
and U10626 (N_10626,N_10280,N_10472);
and U10627 (N_10627,N_10265,N_10335);
nand U10628 (N_10628,N_10282,N_10462);
nand U10629 (N_10629,N_10328,N_10451);
or U10630 (N_10630,N_10410,N_10429);
nor U10631 (N_10631,N_10367,N_10263);
and U10632 (N_10632,N_10497,N_10492);
nand U10633 (N_10633,N_10287,N_10357);
or U10634 (N_10634,N_10423,N_10278);
or U10635 (N_10635,N_10225,N_10342);
nor U10636 (N_10636,N_10498,N_10485);
nand U10637 (N_10637,N_10288,N_10302);
nor U10638 (N_10638,N_10227,N_10428);
or U10639 (N_10639,N_10473,N_10285);
xnor U10640 (N_10640,N_10235,N_10343);
or U10641 (N_10641,N_10456,N_10494);
and U10642 (N_10642,N_10316,N_10331);
nand U10643 (N_10643,N_10332,N_10418);
and U10644 (N_10644,N_10289,N_10253);
nand U10645 (N_10645,N_10386,N_10486);
and U10646 (N_10646,N_10213,N_10236);
and U10647 (N_10647,N_10229,N_10261);
xnor U10648 (N_10648,N_10341,N_10256);
or U10649 (N_10649,N_10371,N_10389);
or U10650 (N_10650,N_10357,N_10398);
xnor U10651 (N_10651,N_10306,N_10459);
xor U10652 (N_10652,N_10413,N_10314);
or U10653 (N_10653,N_10397,N_10236);
nor U10654 (N_10654,N_10363,N_10382);
nor U10655 (N_10655,N_10229,N_10268);
and U10656 (N_10656,N_10366,N_10218);
or U10657 (N_10657,N_10266,N_10470);
xor U10658 (N_10658,N_10494,N_10318);
nor U10659 (N_10659,N_10354,N_10454);
nand U10660 (N_10660,N_10473,N_10356);
nand U10661 (N_10661,N_10489,N_10346);
or U10662 (N_10662,N_10288,N_10386);
xnor U10663 (N_10663,N_10258,N_10358);
nand U10664 (N_10664,N_10330,N_10444);
nor U10665 (N_10665,N_10244,N_10306);
xor U10666 (N_10666,N_10487,N_10248);
or U10667 (N_10667,N_10404,N_10331);
or U10668 (N_10668,N_10441,N_10277);
nand U10669 (N_10669,N_10250,N_10337);
and U10670 (N_10670,N_10245,N_10437);
nor U10671 (N_10671,N_10422,N_10249);
or U10672 (N_10672,N_10252,N_10426);
or U10673 (N_10673,N_10489,N_10342);
nand U10674 (N_10674,N_10381,N_10285);
or U10675 (N_10675,N_10440,N_10481);
nor U10676 (N_10676,N_10339,N_10338);
nand U10677 (N_10677,N_10436,N_10315);
nand U10678 (N_10678,N_10375,N_10398);
and U10679 (N_10679,N_10342,N_10206);
nor U10680 (N_10680,N_10280,N_10414);
or U10681 (N_10681,N_10401,N_10305);
nor U10682 (N_10682,N_10357,N_10460);
and U10683 (N_10683,N_10448,N_10442);
and U10684 (N_10684,N_10398,N_10351);
nand U10685 (N_10685,N_10418,N_10405);
or U10686 (N_10686,N_10402,N_10343);
nand U10687 (N_10687,N_10463,N_10456);
xor U10688 (N_10688,N_10354,N_10450);
and U10689 (N_10689,N_10470,N_10251);
and U10690 (N_10690,N_10451,N_10309);
nand U10691 (N_10691,N_10384,N_10496);
and U10692 (N_10692,N_10492,N_10242);
nand U10693 (N_10693,N_10366,N_10238);
xnor U10694 (N_10694,N_10421,N_10283);
xor U10695 (N_10695,N_10485,N_10307);
nor U10696 (N_10696,N_10294,N_10450);
nor U10697 (N_10697,N_10320,N_10247);
xor U10698 (N_10698,N_10357,N_10239);
nand U10699 (N_10699,N_10463,N_10497);
nand U10700 (N_10700,N_10450,N_10266);
nand U10701 (N_10701,N_10274,N_10220);
and U10702 (N_10702,N_10480,N_10245);
nor U10703 (N_10703,N_10345,N_10453);
xnor U10704 (N_10704,N_10432,N_10368);
nor U10705 (N_10705,N_10262,N_10471);
and U10706 (N_10706,N_10286,N_10464);
and U10707 (N_10707,N_10477,N_10453);
nor U10708 (N_10708,N_10446,N_10272);
or U10709 (N_10709,N_10498,N_10314);
nand U10710 (N_10710,N_10447,N_10337);
and U10711 (N_10711,N_10400,N_10263);
or U10712 (N_10712,N_10307,N_10216);
nand U10713 (N_10713,N_10249,N_10412);
nor U10714 (N_10714,N_10283,N_10255);
nor U10715 (N_10715,N_10325,N_10315);
and U10716 (N_10716,N_10221,N_10491);
nand U10717 (N_10717,N_10488,N_10373);
or U10718 (N_10718,N_10395,N_10306);
and U10719 (N_10719,N_10461,N_10299);
nand U10720 (N_10720,N_10203,N_10365);
xor U10721 (N_10721,N_10470,N_10226);
nand U10722 (N_10722,N_10319,N_10355);
nor U10723 (N_10723,N_10419,N_10340);
xnor U10724 (N_10724,N_10401,N_10329);
and U10725 (N_10725,N_10390,N_10269);
and U10726 (N_10726,N_10481,N_10447);
xnor U10727 (N_10727,N_10261,N_10372);
nand U10728 (N_10728,N_10402,N_10470);
nand U10729 (N_10729,N_10477,N_10267);
nor U10730 (N_10730,N_10261,N_10289);
or U10731 (N_10731,N_10463,N_10459);
and U10732 (N_10732,N_10248,N_10402);
or U10733 (N_10733,N_10369,N_10361);
nor U10734 (N_10734,N_10435,N_10393);
nor U10735 (N_10735,N_10348,N_10398);
or U10736 (N_10736,N_10407,N_10459);
and U10737 (N_10737,N_10274,N_10425);
xnor U10738 (N_10738,N_10321,N_10372);
nor U10739 (N_10739,N_10494,N_10341);
nor U10740 (N_10740,N_10410,N_10277);
nor U10741 (N_10741,N_10271,N_10289);
nor U10742 (N_10742,N_10250,N_10280);
nand U10743 (N_10743,N_10311,N_10396);
nor U10744 (N_10744,N_10418,N_10487);
nor U10745 (N_10745,N_10395,N_10436);
nand U10746 (N_10746,N_10494,N_10229);
and U10747 (N_10747,N_10291,N_10441);
nor U10748 (N_10748,N_10288,N_10346);
and U10749 (N_10749,N_10357,N_10406);
nor U10750 (N_10750,N_10470,N_10202);
and U10751 (N_10751,N_10474,N_10456);
xnor U10752 (N_10752,N_10305,N_10374);
xnor U10753 (N_10753,N_10313,N_10201);
and U10754 (N_10754,N_10442,N_10369);
xor U10755 (N_10755,N_10375,N_10289);
and U10756 (N_10756,N_10394,N_10268);
xnor U10757 (N_10757,N_10438,N_10221);
nand U10758 (N_10758,N_10401,N_10455);
nor U10759 (N_10759,N_10425,N_10250);
and U10760 (N_10760,N_10378,N_10475);
and U10761 (N_10761,N_10315,N_10257);
nor U10762 (N_10762,N_10334,N_10212);
and U10763 (N_10763,N_10255,N_10210);
xor U10764 (N_10764,N_10337,N_10327);
xor U10765 (N_10765,N_10405,N_10309);
and U10766 (N_10766,N_10337,N_10369);
nor U10767 (N_10767,N_10287,N_10200);
nor U10768 (N_10768,N_10316,N_10281);
nor U10769 (N_10769,N_10234,N_10490);
nor U10770 (N_10770,N_10461,N_10232);
nand U10771 (N_10771,N_10246,N_10207);
or U10772 (N_10772,N_10482,N_10317);
and U10773 (N_10773,N_10307,N_10413);
xnor U10774 (N_10774,N_10452,N_10449);
or U10775 (N_10775,N_10277,N_10465);
or U10776 (N_10776,N_10248,N_10490);
nand U10777 (N_10777,N_10291,N_10277);
nor U10778 (N_10778,N_10220,N_10242);
xor U10779 (N_10779,N_10371,N_10281);
nor U10780 (N_10780,N_10487,N_10211);
nor U10781 (N_10781,N_10357,N_10236);
xnor U10782 (N_10782,N_10451,N_10331);
nor U10783 (N_10783,N_10305,N_10290);
xor U10784 (N_10784,N_10372,N_10234);
xnor U10785 (N_10785,N_10272,N_10494);
nor U10786 (N_10786,N_10484,N_10369);
and U10787 (N_10787,N_10283,N_10473);
and U10788 (N_10788,N_10319,N_10464);
xor U10789 (N_10789,N_10320,N_10337);
nor U10790 (N_10790,N_10240,N_10335);
and U10791 (N_10791,N_10418,N_10344);
nand U10792 (N_10792,N_10288,N_10383);
or U10793 (N_10793,N_10430,N_10447);
nand U10794 (N_10794,N_10334,N_10372);
and U10795 (N_10795,N_10428,N_10374);
and U10796 (N_10796,N_10227,N_10288);
xnor U10797 (N_10797,N_10375,N_10480);
xnor U10798 (N_10798,N_10490,N_10205);
or U10799 (N_10799,N_10471,N_10323);
or U10800 (N_10800,N_10789,N_10737);
nor U10801 (N_10801,N_10703,N_10621);
or U10802 (N_10802,N_10712,N_10577);
nor U10803 (N_10803,N_10582,N_10507);
and U10804 (N_10804,N_10641,N_10516);
nor U10805 (N_10805,N_10740,N_10739);
nor U10806 (N_10806,N_10607,N_10731);
nor U10807 (N_10807,N_10661,N_10776);
nor U10808 (N_10808,N_10609,N_10706);
nor U10809 (N_10809,N_10514,N_10671);
and U10810 (N_10810,N_10742,N_10688);
nor U10811 (N_10811,N_10658,N_10748);
xor U10812 (N_10812,N_10560,N_10669);
xnor U10813 (N_10813,N_10612,N_10628);
or U10814 (N_10814,N_10747,N_10713);
and U10815 (N_10815,N_10589,N_10623);
and U10816 (N_10816,N_10639,N_10636);
or U10817 (N_10817,N_10627,N_10633);
and U10818 (N_10818,N_10724,N_10777);
xnor U10819 (N_10819,N_10592,N_10734);
or U10820 (N_10820,N_10644,N_10642);
and U10821 (N_10821,N_10538,N_10537);
xnor U10822 (N_10822,N_10542,N_10652);
nand U10823 (N_10823,N_10565,N_10718);
and U10824 (N_10824,N_10517,N_10610);
and U10825 (N_10825,N_10505,N_10526);
or U10826 (N_10826,N_10753,N_10611);
or U10827 (N_10827,N_10561,N_10599);
nand U10828 (N_10828,N_10751,N_10735);
or U10829 (N_10829,N_10668,N_10567);
nand U10830 (N_10830,N_10778,N_10660);
and U10831 (N_10831,N_10637,N_10667);
nand U10832 (N_10832,N_10760,N_10682);
or U10833 (N_10833,N_10521,N_10529);
nor U10834 (N_10834,N_10580,N_10763);
nor U10835 (N_10835,N_10715,N_10757);
nand U10836 (N_10836,N_10525,N_10775);
or U10837 (N_10837,N_10579,N_10566);
and U10838 (N_10838,N_10512,N_10531);
nor U10839 (N_10839,N_10646,N_10683);
and U10840 (N_10840,N_10519,N_10794);
or U10841 (N_10841,N_10768,N_10587);
nor U10842 (N_10842,N_10695,N_10554);
and U10843 (N_10843,N_10532,N_10750);
xor U10844 (N_10844,N_10557,N_10745);
or U10845 (N_10845,N_10595,N_10593);
or U10846 (N_10846,N_10543,N_10569);
nand U10847 (N_10847,N_10733,N_10720);
nand U10848 (N_10848,N_10602,N_10769);
xor U10849 (N_10849,N_10727,N_10536);
nor U10850 (N_10850,N_10506,N_10618);
nand U10851 (N_10851,N_10786,N_10701);
or U10852 (N_10852,N_10551,N_10544);
and U10853 (N_10853,N_10691,N_10766);
nand U10854 (N_10854,N_10600,N_10511);
nor U10855 (N_10855,N_10732,N_10620);
and U10856 (N_10856,N_10702,N_10550);
and U10857 (N_10857,N_10509,N_10736);
nor U10858 (N_10858,N_10522,N_10603);
xor U10859 (N_10859,N_10524,N_10541);
nor U10860 (N_10860,N_10500,N_10705);
and U10861 (N_10861,N_10788,N_10635);
nor U10862 (N_10862,N_10534,N_10616);
or U10863 (N_10863,N_10685,N_10651);
xor U10864 (N_10864,N_10798,N_10722);
or U10865 (N_10865,N_10749,N_10594);
nand U10866 (N_10866,N_10773,N_10717);
xor U10867 (N_10867,N_10648,N_10547);
and U10868 (N_10868,N_10540,N_10795);
nor U10869 (N_10869,N_10649,N_10570);
and U10870 (N_10870,N_10729,N_10704);
nand U10871 (N_10871,N_10694,N_10555);
and U10872 (N_10872,N_10546,N_10634);
or U10873 (N_10873,N_10614,N_10656);
xnor U10874 (N_10874,N_10679,N_10548);
nand U10875 (N_10875,N_10608,N_10689);
xor U10876 (N_10876,N_10772,N_10533);
or U10877 (N_10877,N_10674,N_10755);
or U10878 (N_10878,N_10640,N_10714);
or U10879 (N_10879,N_10663,N_10692);
xor U10880 (N_10880,N_10723,N_10698);
nor U10881 (N_10881,N_10782,N_10559);
and U10882 (N_10882,N_10665,N_10508);
and U10883 (N_10883,N_10764,N_10647);
nor U10884 (N_10884,N_10796,N_10588);
nor U10885 (N_10885,N_10711,N_10619);
and U10886 (N_10886,N_10553,N_10575);
xnor U10887 (N_10887,N_10662,N_10653);
and U10888 (N_10888,N_10571,N_10716);
xor U10889 (N_10889,N_10791,N_10693);
nand U10890 (N_10890,N_10754,N_10684);
nor U10891 (N_10891,N_10774,N_10686);
or U10892 (N_10892,N_10539,N_10770);
nor U10893 (N_10893,N_10549,N_10576);
xor U10894 (N_10894,N_10672,N_10645);
xor U10895 (N_10895,N_10578,N_10622);
nor U10896 (N_10896,N_10585,N_10767);
xor U10897 (N_10897,N_10598,N_10676);
nor U10898 (N_10898,N_10564,N_10629);
nand U10899 (N_10899,N_10756,N_10655);
or U10900 (N_10900,N_10743,N_10591);
nand U10901 (N_10901,N_10708,N_10518);
xor U10902 (N_10902,N_10503,N_10624);
xor U10903 (N_10903,N_10631,N_10730);
nand U10904 (N_10904,N_10527,N_10697);
xnor U10905 (N_10905,N_10659,N_10530);
nor U10906 (N_10906,N_10523,N_10677);
nand U10907 (N_10907,N_10752,N_10746);
nand U10908 (N_10908,N_10545,N_10586);
and U10909 (N_10909,N_10574,N_10573);
nor U10910 (N_10910,N_10759,N_10707);
nor U10911 (N_10911,N_10654,N_10625);
nor U10912 (N_10912,N_10687,N_10613);
and U10913 (N_10913,N_10630,N_10785);
nand U10914 (N_10914,N_10710,N_10681);
or U10915 (N_10915,N_10792,N_10657);
xor U10916 (N_10916,N_10673,N_10728);
nand U10917 (N_10917,N_10699,N_10604);
nor U10918 (N_10918,N_10581,N_10556);
nand U10919 (N_10919,N_10784,N_10605);
nand U10920 (N_10920,N_10725,N_10562);
and U10921 (N_10921,N_10513,N_10558);
nor U10922 (N_10922,N_10762,N_10583);
xnor U10923 (N_10923,N_10596,N_10590);
nor U10924 (N_10924,N_10738,N_10680);
nor U10925 (N_10925,N_10700,N_10790);
nand U10926 (N_10926,N_10563,N_10765);
nand U10927 (N_10927,N_10568,N_10799);
xnor U10928 (N_10928,N_10678,N_10510);
and U10929 (N_10929,N_10719,N_10601);
nor U10930 (N_10930,N_10626,N_10780);
xor U10931 (N_10931,N_10721,N_10572);
nor U10932 (N_10932,N_10781,N_10638);
xnor U10933 (N_10933,N_10528,N_10535);
nor U10934 (N_10934,N_10666,N_10709);
and U10935 (N_10935,N_10650,N_10584);
nand U10936 (N_10936,N_10771,N_10664);
nor U10937 (N_10937,N_10779,N_10758);
nand U10938 (N_10938,N_10632,N_10787);
nand U10939 (N_10939,N_10552,N_10643);
and U10940 (N_10940,N_10690,N_10783);
nand U10941 (N_10941,N_10597,N_10726);
nand U10942 (N_10942,N_10744,N_10617);
nand U10943 (N_10943,N_10615,N_10793);
or U10944 (N_10944,N_10696,N_10501);
nand U10945 (N_10945,N_10797,N_10515);
and U10946 (N_10946,N_10670,N_10741);
or U10947 (N_10947,N_10502,N_10504);
xor U10948 (N_10948,N_10675,N_10761);
or U10949 (N_10949,N_10520,N_10606);
xor U10950 (N_10950,N_10556,N_10500);
nor U10951 (N_10951,N_10688,N_10768);
nand U10952 (N_10952,N_10621,N_10697);
nor U10953 (N_10953,N_10707,N_10531);
nor U10954 (N_10954,N_10767,N_10772);
or U10955 (N_10955,N_10692,N_10586);
and U10956 (N_10956,N_10653,N_10737);
or U10957 (N_10957,N_10607,N_10702);
or U10958 (N_10958,N_10535,N_10506);
xnor U10959 (N_10959,N_10663,N_10657);
xor U10960 (N_10960,N_10748,N_10583);
xnor U10961 (N_10961,N_10598,N_10570);
nand U10962 (N_10962,N_10570,N_10642);
xor U10963 (N_10963,N_10765,N_10742);
xor U10964 (N_10964,N_10687,N_10757);
or U10965 (N_10965,N_10706,N_10662);
xnor U10966 (N_10966,N_10618,N_10740);
or U10967 (N_10967,N_10604,N_10524);
xnor U10968 (N_10968,N_10742,N_10781);
xor U10969 (N_10969,N_10724,N_10683);
and U10970 (N_10970,N_10723,N_10779);
or U10971 (N_10971,N_10510,N_10659);
nand U10972 (N_10972,N_10710,N_10651);
xnor U10973 (N_10973,N_10513,N_10502);
or U10974 (N_10974,N_10522,N_10716);
nor U10975 (N_10975,N_10662,N_10590);
nor U10976 (N_10976,N_10675,N_10572);
xnor U10977 (N_10977,N_10658,N_10666);
xor U10978 (N_10978,N_10541,N_10550);
or U10979 (N_10979,N_10650,N_10603);
or U10980 (N_10980,N_10712,N_10626);
or U10981 (N_10981,N_10734,N_10637);
nand U10982 (N_10982,N_10558,N_10777);
or U10983 (N_10983,N_10756,N_10779);
or U10984 (N_10984,N_10626,N_10741);
xor U10985 (N_10985,N_10536,N_10718);
and U10986 (N_10986,N_10715,N_10580);
nor U10987 (N_10987,N_10697,N_10783);
and U10988 (N_10988,N_10713,N_10796);
nand U10989 (N_10989,N_10797,N_10505);
nor U10990 (N_10990,N_10705,N_10681);
and U10991 (N_10991,N_10661,N_10779);
nand U10992 (N_10992,N_10512,N_10625);
nor U10993 (N_10993,N_10709,N_10702);
or U10994 (N_10994,N_10650,N_10680);
nand U10995 (N_10995,N_10537,N_10524);
nand U10996 (N_10996,N_10610,N_10510);
or U10997 (N_10997,N_10767,N_10675);
and U10998 (N_10998,N_10647,N_10743);
xor U10999 (N_10999,N_10792,N_10669);
and U11000 (N_11000,N_10798,N_10503);
nor U11001 (N_11001,N_10622,N_10694);
nor U11002 (N_11002,N_10785,N_10561);
or U11003 (N_11003,N_10545,N_10673);
or U11004 (N_11004,N_10579,N_10510);
nor U11005 (N_11005,N_10614,N_10680);
and U11006 (N_11006,N_10777,N_10705);
nor U11007 (N_11007,N_10765,N_10510);
xor U11008 (N_11008,N_10612,N_10615);
or U11009 (N_11009,N_10746,N_10535);
nand U11010 (N_11010,N_10769,N_10523);
xor U11011 (N_11011,N_10715,N_10712);
or U11012 (N_11012,N_10565,N_10518);
xnor U11013 (N_11013,N_10541,N_10644);
and U11014 (N_11014,N_10628,N_10721);
or U11015 (N_11015,N_10784,N_10690);
or U11016 (N_11016,N_10789,N_10724);
xor U11017 (N_11017,N_10729,N_10617);
and U11018 (N_11018,N_10689,N_10543);
nor U11019 (N_11019,N_10590,N_10598);
nand U11020 (N_11020,N_10771,N_10651);
and U11021 (N_11021,N_10701,N_10572);
nand U11022 (N_11022,N_10564,N_10668);
or U11023 (N_11023,N_10561,N_10731);
nor U11024 (N_11024,N_10744,N_10612);
nand U11025 (N_11025,N_10751,N_10749);
nand U11026 (N_11026,N_10632,N_10647);
and U11027 (N_11027,N_10616,N_10542);
or U11028 (N_11028,N_10616,N_10564);
nand U11029 (N_11029,N_10573,N_10682);
xor U11030 (N_11030,N_10758,N_10788);
xnor U11031 (N_11031,N_10511,N_10767);
nor U11032 (N_11032,N_10700,N_10514);
and U11033 (N_11033,N_10649,N_10636);
nor U11034 (N_11034,N_10774,N_10521);
and U11035 (N_11035,N_10667,N_10788);
xor U11036 (N_11036,N_10584,N_10640);
xnor U11037 (N_11037,N_10742,N_10768);
nand U11038 (N_11038,N_10731,N_10620);
nand U11039 (N_11039,N_10673,N_10657);
nor U11040 (N_11040,N_10623,N_10564);
and U11041 (N_11041,N_10689,N_10632);
nand U11042 (N_11042,N_10662,N_10710);
nor U11043 (N_11043,N_10664,N_10787);
and U11044 (N_11044,N_10747,N_10622);
nand U11045 (N_11045,N_10570,N_10700);
or U11046 (N_11046,N_10640,N_10537);
nor U11047 (N_11047,N_10689,N_10532);
xor U11048 (N_11048,N_10685,N_10769);
nor U11049 (N_11049,N_10555,N_10623);
or U11050 (N_11050,N_10727,N_10527);
nor U11051 (N_11051,N_10797,N_10511);
or U11052 (N_11052,N_10566,N_10611);
or U11053 (N_11053,N_10681,N_10798);
xnor U11054 (N_11054,N_10525,N_10524);
xor U11055 (N_11055,N_10720,N_10558);
or U11056 (N_11056,N_10761,N_10520);
and U11057 (N_11057,N_10564,N_10775);
nand U11058 (N_11058,N_10765,N_10626);
xnor U11059 (N_11059,N_10533,N_10635);
or U11060 (N_11060,N_10566,N_10581);
and U11061 (N_11061,N_10681,N_10598);
and U11062 (N_11062,N_10766,N_10695);
and U11063 (N_11063,N_10756,N_10732);
nor U11064 (N_11064,N_10787,N_10743);
and U11065 (N_11065,N_10796,N_10631);
or U11066 (N_11066,N_10796,N_10596);
and U11067 (N_11067,N_10688,N_10750);
nor U11068 (N_11068,N_10611,N_10619);
and U11069 (N_11069,N_10587,N_10630);
and U11070 (N_11070,N_10762,N_10679);
and U11071 (N_11071,N_10599,N_10623);
xor U11072 (N_11072,N_10706,N_10773);
nand U11073 (N_11073,N_10566,N_10649);
or U11074 (N_11074,N_10768,N_10526);
and U11075 (N_11075,N_10640,N_10746);
and U11076 (N_11076,N_10666,N_10743);
xor U11077 (N_11077,N_10509,N_10726);
nor U11078 (N_11078,N_10715,N_10563);
nor U11079 (N_11079,N_10645,N_10667);
xnor U11080 (N_11080,N_10781,N_10532);
or U11081 (N_11081,N_10752,N_10506);
nand U11082 (N_11082,N_10737,N_10761);
nor U11083 (N_11083,N_10787,N_10736);
and U11084 (N_11084,N_10792,N_10642);
nand U11085 (N_11085,N_10510,N_10615);
and U11086 (N_11086,N_10783,N_10767);
nor U11087 (N_11087,N_10621,N_10701);
nand U11088 (N_11088,N_10767,N_10520);
or U11089 (N_11089,N_10670,N_10514);
nor U11090 (N_11090,N_10777,N_10595);
nand U11091 (N_11091,N_10790,N_10654);
or U11092 (N_11092,N_10612,N_10643);
nand U11093 (N_11093,N_10587,N_10536);
nor U11094 (N_11094,N_10523,N_10560);
nor U11095 (N_11095,N_10510,N_10723);
or U11096 (N_11096,N_10514,N_10690);
nand U11097 (N_11097,N_10602,N_10538);
or U11098 (N_11098,N_10595,N_10727);
xor U11099 (N_11099,N_10647,N_10694);
xor U11100 (N_11100,N_11080,N_10897);
xnor U11101 (N_11101,N_10986,N_11030);
nand U11102 (N_11102,N_11067,N_10831);
xnor U11103 (N_11103,N_10956,N_10950);
or U11104 (N_11104,N_10812,N_11081);
xnor U11105 (N_11105,N_10889,N_10911);
nand U11106 (N_11106,N_11066,N_10962);
nand U11107 (N_11107,N_11050,N_10876);
nor U11108 (N_11108,N_10825,N_11077);
xnor U11109 (N_11109,N_11005,N_11059);
xor U11110 (N_11110,N_11038,N_10830);
nand U11111 (N_11111,N_10861,N_11032);
or U11112 (N_11112,N_10912,N_10909);
and U11113 (N_11113,N_11099,N_10864);
nor U11114 (N_11114,N_10822,N_10824);
nand U11115 (N_11115,N_10965,N_10899);
xnor U11116 (N_11116,N_10934,N_10903);
xor U11117 (N_11117,N_11016,N_11092);
nor U11118 (N_11118,N_10910,N_11095);
nand U11119 (N_11119,N_11057,N_11088);
or U11120 (N_11120,N_10813,N_10845);
and U11121 (N_11121,N_11048,N_10804);
nor U11122 (N_11122,N_11078,N_10891);
nor U11123 (N_11123,N_10960,N_11022);
or U11124 (N_11124,N_11021,N_10916);
xor U11125 (N_11125,N_11097,N_10963);
or U11126 (N_11126,N_10945,N_10947);
and U11127 (N_11127,N_10905,N_11046);
xor U11128 (N_11128,N_11051,N_10879);
and U11129 (N_11129,N_10811,N_10875);
or U11130 (N_11130,N_11075,N_11056);
xnor U11131 (N_11131,N_11012,N_11049);
and U11132 (N_11132,N_11083,N_10959);
nand U11133 (N_11133,N_10968,N_10955);
and U11134 (N_11134,N_10829,N_10842);
nand U11135 (N_11135,N_10866,N_10840);
nand U11136 (N_11136,N_10940,N_10838);
nor U11137 (N_11137,N_10800,N_10852);
and U11138 (N_11138,N_11070,N_10856);
and U11139 (N_11139,N_11089,N_11074);
nor U11140 (N_11140,N_10874,N_10832);
nor U11141 (N_11141,N_10890,N_11020);
or U11142 (N_11142,N_11031,N_10884);
nor U11143 (N_11143,N_10805,N_10818);
and U11144 (N_11144,N_11062,N_10966);
nor U11145 (N_11145,N_10898,N_10894);
nand U11146 (N_11146,N_11076,N_10815);
nand U11147 (N_11147,N_10953,N_10877);
or U11148 (N_11148,N_10993,N_10855);
nand U11149 (N_11149,N_11042,N_10821);
and U11150 (N_11150,N_11018,N_11069);
xnor U11151 (N_11151,N_11064,N_11043);
xnor U11152 (N_11152,N_10979,N_10974);
nor U11153 (N_11153,N_11011,N_10814);
xor U11154 (N_11154,N_11055,N_10972);
xnor U11155 (N_11155,N_10941,N_10990);
xnor U11156 (N_11156,N_10902,N_10881);
or U11157 (N_11157,N_11065,N_10843);
xnor U11158 (N_11158,N_10850,N_11096);
and U11159 (N_11159,N_10980,N_10844);
or U11160 (N_11160,N_10983,N_10969);
nand U11161 (N_11161,N_10878,N_11007);
xnor U11162 (N_11162,N_10998,N_11029);
nand U11163 (N_11163,N_10927,N_11037);
nand U11164 (N_11164,N_10937,N_11094);
nand U11165 (N_11165,N_10924,N_10883);
and U11166 (N_11166,N_10802,N_10808);
or U11167 (N_11167,N_11009,N_10880);
xnor U11168 (N_11168,N_10833,N_11024);
xor U11169 (N_11169,N_11028,N_11002);
nand U11170 (N_11170,N_10939,N_10904);
or U11171 (N_11171,N_11045,N_10892);
and U11172 (N_11172,N_10893,N_10801);
nor U11173 (N_11173,N_10989,N_10920);
nand U11174 (N_11174,N_10870,N_11026);
nor U11175 (N_11175,N_10846,N_10847);
and U11176 (N_11176,N_10922,N_10834);
nand U11177 (N_11177,N_10865,N_10828);
nor U11178 (N_11178,N_10970,N_10896);
xnor U11179 (N_11179,N_10849,N_10987);
nor U11180 (N_11180,N_10809,N_11041);
xnor U11181 (N_11181,N_11040,N_10913);
nand U11182 (N_11182,N_10984,N_11093);
nand U11183 (N_11183,N_11033,N_10938);
xor U11184 (N_11184,N_10976,N_10997);
and U11185 (N_11185,N_11098,N_11025);
xor U11186 (N_11186,N_11087,N_10826);
and U11187 (N_11187,N_10949,N_10961);
nand U11188 (N_11188,N_10820,N_10851);
and U11189 (N_11189,N_10857,N_11061);
and U11190 (N_11190,N_10895,N_11039);
and U11191 (N_11191,N_10819,N_10917);
or U11192 (N_11192,N_10853,N_10873);
and U11193 (N_11193,N_10836,N_10914);
and U11194 (N_11194,N_10839,N_10928);
nor U11195 (N_11195,N_10887,N_10869);
nor U11196 (N_11196,N_10872,N_11023);
nor U11197 (N_11197,N_10988,N_11063);
and U11198 (N_11198,N_10816,N_10933);
or U11199 (N_11199,N_11003,N_11017);
and U11200 (N_11200,N_10868,N_10803);
nand U11201 (N_11201,N_10823,N_10995);
nand U11202 (N_11202,N_10867,N_11044);
and U11203 (N_11203,N_11004,N_11082);
nand U11204 (N_11204,N_11013,N_10944);
nor U11205 (N_11205,N_10952,N_10994);
nor U11206 (N_11206,N_11091,N_10992);
and U11207 (N_11207,N_10921,N_11036);
nor U11208 (N_11208,N_10919,N_10935);
or U11209 (N_11209,N_10837,N_10859);
or U11210 (N_11210,N_11071,N_11072);
and U11211 (N_11211,N_10977,N_10982);
or U11212 (N_11212,N_10951,N_11027);
and U11213 (N_11213,N_11008,N_11001);
nor U11214 (N_11214,N_10973,N_10888);
and U11215 (N_11215,N_10848,N_11010);
nor U11216 (N_11216,N_11068,N_10918);
and U11217 (N_11217,N_10907,N_10835);
nor U11218 (N_11218,N_10810,N_11073);
or U11219 (N_11219,N_10862,N_10981);
nor U11220 (N_11220,N_11090,N_11015);
and U11221 (N_11221,N_10943,N_10871);
or U11222 (N_11222,N_10948,N_10908);
xnor U11223 (N_11223,N_10858,N_10885);
xnor U11224 (N_11224,N_10996,N_11060);
xor U11225 (N_11225,N_10900,N_10860);
nor U11226 (N_11226,N_11035,N_10936);
xnor U11227 (N_11227,N_11079,N_11019);
or U11228 (N_11228,N_11000,N_10806);
nand U11229 (N_11229,N_10985,N_10999);
xnor U11230 (N_11230,N_10991,N_11034);
nor U11231 (N_11231,N_10931,N_11006);
nand U11232 (N_11232,N_10971,N_11047);
xor U11233 (N_11233,N_10932,N_10923);
nor U11234 (N_11234,N_10978,N_10942);
xor U11235 (N_11235,N_10827,N_10925);
nand U11236 (N_11236,N_10967,N_10817);
and U11237 (N_11237,N_10854,N_10915);
or U11238 (N_11238,N_11084,N_10926);
and U11239 (N_11239,N_11053,N_10958);
nor U11240 (N_11240,N_10901,N_10975);
nor U11241 (N_11241,N_11014,N_10954);
xor U11242 (N_11242,N_11054,N_10957);
nor U11243 (N_11243,N_10929,N_10946);
or U11244 (N_11244,N_11086,N_11058);
and U11245 (N_11245,N_11085,N_10906);
and U11246 (N_11246,N_10886,N_10863);
nor U11247 (N_11247,N_10930,N_10882);
nor U11248 (N_11248,N_11052,N_10807);
and U11249 (N_11249,N_10841,N_10964);
nand U11250 (N_11250,N_11029,N_10843);
and U11251 (N_11251,N_10853,N_10861);
nand U11252 (N_11252,N_11053,N_10893);
nand U11253 (N_11253,N_10939,N_10943);
and U11254 (N_11254,N_10944,N_11090);
nand U11255 (N_11255,N_10896,N_11086);
nor U11256 (N_11256,N_10823,N_10950);
or U11257 (N_11257,N_10965,N_10872);
xor U11258 (N_11258,N_11093,N_10943);
nand U11259 (N_11259,N_11038,N_11089);
nor U11260 (N_11260,N_11098,N_11070);
nand U11261 (N_11261,N_10847,N_10934);
and U11262 (N_11262,N_11097,N_10886);
or U11263 (N_11263,N_11017,N_10977);
xor U11264 (N_11264,N_11087,N_11076);
or U11265 (N_11265,N_11003,N_10983);
nand U11266 (N_11266,N_10895,N_10801);
and U11267 (N_11267,N_10972,N_10869);
or U11268 (N_11268,N_10919,N_10995);
nor U11269 (N_11269,N_10914,N_10956);
and U11270 (N_11270,N_10933,N_10835);
nor U11271 (N_11271,N_10929,N_10858);
xor U11272 (N_11272,N_11067,N_10855);
xnor U11273 (N_11273,N_10822,N_11040);
or U11274 (N_11274,N_10935,N_10973);
or U11275 (N_11275,N_10990,N_10932);
nand U11276 (N_11276,N_10853,N_10908);
xor U11277 (N_11277,N_10973,N_10906);
nor U11278 (N_11278,N_10925,N_11026);
nand U11279 (N_11279,N_10869,N_11062);
nand U11280 (N_11280,N_10947,N_10981);
nor U11281 (N_11281,N_10801,N_11044);
xor U11282 (N_11282,N_10858,N_10939);
or U11283 (N_11283,N_10968,N_11025);
or U11284 (N_11284,N_10926,N_11080);
nand U11285 (N_11285,N_11011,N_10803);
or U11286 (N_11286,N_10819,N_11067);
and U11287 (N_11287,N_11012,N_11078);
xor U11288 (N_11288,N_11003,N_10985);
nand U11289 (N_11289,N_10929,N_11057);
nor U11290 (N_11290,N_10930,N_10978);
nand U11291 (N_11291,N_11034,N_10864);
nand U11292 (N_11292,N_11090,N_11071);
or U11293 (N_11293,N_10883,N_10953);
or U11294 (N_11294,N_10864,N_11018);
or U11295 (N_11295,N_10821,N_10827);
or U11296 (N_11296,N_10866,N_11023);
or U11297 (N_11297,N_10850,N_10870);
nor U11298 (N_11298,N_10907,N_10979);
xnor U11299 (N_11299,N_10921,N_11022);
nand U11300 (N_11300,N_10975,N_10962);
or U11301 (N_11301,N_10941,N_10804);
and U11302 (N_11302,N_11012,N_11016);
nor U11303 (N_11303,N_11088,N_10816);
nand U11304 (N_11304,N_10871,N_11087);
xor U11305 (N_11305,N_10853,N_10995);
or U11306 (N_11306,N_10836,N_10874);
and U11307 (N_11307,N_10849,N_11081);
and U11308 (N_11308,N_11098,N_10870);
or U11309 (N_11309,N_10804,N_10813);
nor U11310 (N_11310,N_10917,N_10899);
xnor U11311 (N_11311,N_11093,N_11088);
or U11312 (N_11312,N_10907,N_11036);
or U11313 (N_11313,N_11030,N_10953);
nand U11314 (N_11314,N_10982,N_10858);
nand U11315 (N_11315,N_11002,N_10957);
nor U11316 (N_11316,N_10941,N_11007);
or U11317 (N_11317,N_10986,N_10833);
nand U11318 (N_11318,N_10852,N_10856);
or U11319 (N_11319,N_11019,N_10972);
xnor U11320 (N_11320,N_10916,N_10919);
and U11321 (N_11321,N_10960,N_10810);
xor U11322 (N_11322,N_10803,N_11090);
and U11323 (N_11323,N_11010,N_10959);
nor U11324 (N_11324,N_10961,N_10852);
xnor U11325 (N_11325,N_10940,N_11050);
nor U11326 (N_11326,N_10980,N_10930);
and U11327 (N_11327,N_10893,N_10815);
nand U11328 (N_11328,N_11008,N_10954);
xor U11329 (N_11329,N_10865,N_11035);
or U11330 (N_11330,N_10916,N_10974);
nand U11331 (N_11331,N_11029,N_10949);
nor U11332 (N_11332,N_10945,N_11025);
xor U11333 (N_11333,N_11034,N_10998);
or U11334 (N_11334,N_11069,N_10963);
or U11335 (N_11335,N_10815,N_10850);
nand U11336 (N_11336,N_11061,N_11054);
xnor U11337 (N_11337,N_11049,N_10980);
or U11338 (N_11338,N_10847,N_10894);
nand U11339 (N_11339,N_10834,N_10849);
and U11340 (N_11340,N_10927,N_10901);
xnor U11341 (N_11341,N_10916,N_10868);
nand U11342 (N_11342,N_10954,N_10892);
or U11343 (N_11343,N_10923,N_11047);
nor U11344 (N_11344,N_11074,N_11042);
nand U11345 (N_11345,N_10955,N_11060);
or U11346 (N_11346,N_10975,N_10807);
nor U11347 (N_11347,N_10838,N_10843);
and U11348 (N_11348,N_10945,N_10901);
nor U11349 (N_11349,N_11050,N_10843);
or U11350 (N_11350,N_10868,N_10995);
xor U11351 (N_11351,N_11014,N_10807);
and U11352 (N_11352,N_11015,N_10915);
or U11353 (N_11353,N_11065,N_10988);
or U11354 (N_11354,N_10835,N_11020);
nor U11355 (N_11355,N_11058,N_11063);
nand U11356 (N_11356,N_10838,N_10830);
and U11357 (N_11357,N_10942,N_11073);
nor U11358 (N_11358,N_11040,N_10987);
nor U11359 (N_11359,N_10801,N_11091);
or U11360 (N_11360,N_11083,N_11024);
or U11361 (N_11361,N_10850,N_10884);
nand U11362 (N_11362,N_10883,N_10976);
xor U11363 (N_11363,N_10841,N_11091);
nor U11364 (N_11364,N_11066,N_11016);
or U11365 (N_11365,N_11007,N_10881);
nor U11366 (N_11366,N_11079,N_11058);
and U11367 (N_11367,N_11054,N_10870);
nor U11368 (N_11368,N_10889,N_10807);
nor U11369 (N_11369,N_11003,N_11029);
and U11370 (N_11370,N_11041,N_11083);
nor U11371 (N_11371,N_10941,N_10949);
nor U11372 (N_11372,N_10847,N_11088);
xnor U11373 (N_11373,N_11028,N_11096);
and U11374 (N_11374,N_10904,N_10820);
or U11375 (N_11375,N_11004,N_10902);
and U11376 (N_11376,N_10834,N_10848);
or U11377 (N_11377,N_10983,N_10952);
or U11378 (N_11378,N_10979,N_10807);
or U11379 (N_11379,N_10863,N_11035);
xnor U11380 (N_11380,N_11037,N_11023);
and U11381 (N_11381,N_11060,N_10888);
and U11382 (N_11382,N_11011,N_11045);
xor U11383 (N_11383,N_11049,N_11010);
or U11384 (N_11384,N_10923,N_10866);
and U11385 (N_11385,N_10938,N_10923);
or U11386 (N_11386,N_10894,N_10977);
xor U11387 (N_11387,N_10967,N_10915);
xnor U11388 (N_11388,N_10952,N_11084);
xnor U11389 (N_11389,N_10934,N_10945);
nor U11390 (N_11390,N_10902,N_11057);
nand U11391 (N_11391,N_10814,N_10988);
or U11392 (N_11392,N_10824,N_10924);
nand U11393 (N_11393,N_11020,N_10960);
or U11394 (N_11394,N_10924,N_10956);
xnor U11395 (N_11395,N_10891,N_11031);
xor U11396 (N_11396,N_10845,N_10935);
and U11397 (N_11397,N_11081,N_11070);
and U11398 (N_11398,N_10938,N_10882);
and U11399 (N_11399,N_10900,N_11018);
nor U11400 (N_11400,N_11196,N_11138);
nand U11401 (N_11401,N_11160,N_11308);
nand U11402 (N_11402,N_11128,N_11314);
or U11403 (N_11403,N_11258,N_11276);
xor U11404 (N_11404,N_11312,N_11140);
xnor U11405 (N_11405,N_11331,N_11235);
and U11406 (N_11406,N_11391,N_11365);
and U11407 (N_11407,N_11233,N_11379);
nor U11408 (N_11408,N_11168,N_11121);
and U11409 (N_11409,N_11161,N_11373);
nand U11410 (N_11410,N_11100,N_11164);
nand U11411 (N_11411,N_11209,N_11337);
xor U11412 (N_11412,N_11377,N_11122);
xor U11413 (N_11413,N_11252,N_11107);
xor U11414 (N_11414,N_11204,N_11368);
nand U11415 (N_11415,N_11399,N_11364);
nand U11416 (N_11416,N_11201,N_11398);
xnor U11417 (N_11417,N_11305,N_11354);
nor U11418 (N_11418,N_11386,N_11321);
or U11419 (N_11419,N_11306,N_11264);
nand U11420 (N_11420,N_11370,N_11147);
or U11421 (N_11421,N_11260,N_11342);
and U11422 (N_11422,N_11246,N_11385);
nand U11423 (N_11423,N_11299,N_11101);
nor U11424 (N_11424,N_11292,N_11175);
nor U11425 (N_11425,N_11126,N_11110);
nand U11426 (N_11426,N_11125,N_11149);
nand U11427 (N_11427,N_11394,N_11350);
xnor U11428 (N_11428,N_11120,N_11150);
nor U11429 (N_11429,N_11389,N_11270);
and U11430 (N_11430,N_11297,N_11111);
xor U11431 (N_11431,N_11349,N_11363);
nor U11432 (N_11432,N_11152,N_11362);
nand U11433 (N_11433,N_11341,N_11369);
or U11434 (N_11434,N_11181,N_11115);
and U11435 (N_11435,N_11248,N_11287);
or U11436 (N_11436,N_11145,N_11295);
and U11437 (N_11437,N_11375,N_11320);
and U11438 (N_11438,N_11393,N_11214);
and U11439 (N_11439,N_11199,N_11281);
nor U11440 (N_11440,N_11189,N_11234);
or U11441 (N_11441,N_11244,N_11279);
nor U11442 (N_11442,N_11253,N_11268);
xnor U11443 (N_11443,N_11374,N_11351);
xor U11444 (N_11444,N_11294,N_11262);
or U11445 (N_11445,N_11177,N_11219);
nand U11446 (N_11446,N_11289,N_11272);
xor U11447 (N_11447,N_11284,N_11136);
xnor U11448 (N_11448,N_11215,N_11153);
or U11449 (N_11449,N_11293,N_11275);
and U11450 (N_11450,N_11170,N_11242);
xnor U11451 (N_11451,N_11129,N_11302);
nor U11452 (N_11452,N_11166,N_11203);
nand U11453 (N_11453,N_11271,N_11213);
nand U11454 (N_11454,N_11344,N_11217);
or U11455 (N_11455,N_11301,N_11176);
or U11456 (N_11456,N_11243,N_11266);
or U11457 (N_11457,N_11134,N_11356);
xnor U11458 (N_11458,N_11334,N_11114);
and U11459 (N_11459,N_11208,N_11307);
nand U11460 (N_11460,N_11395,N_11171);
and U11461 (N_11461,N_11240,N_11232);
nor U11462 (N_11462,N_11193,N_11291);
or U11463 (N_11463,N_11322,N_11227);
nand U11464 (N_11464,N_11104,N_11282);
or U11465 (N_11465,N_11113,N_11194);
or U11466 (N_11466,N_11135,N_11187);
xnor U11467 (N_11467,N_11367,N_11336);
nor U11468 (N_11468,N_11165,N_11323);
xor U11469 (N_11469,N_11250,N_11202);
nor U11470 (N_11470,N_11223,N_11315);
or U11471 (N_11471,N_11159,N_11188);
nand U11472 (N_11472,N_11303,N_11340);
nand U11473 (N_11473,N_11130,N_11296);
nand U11474 (N_11474,N_11155,N_11283);
nand U11475 (N_11475,N_11298,N_11222);
nor U11476 (N_11476,N_11206,N_11387);
nand U11477 (N_11477,N_11180,N_11238);
or U11478 (N_11478,N_11324,N_11257);
nand U11479 (N_11479,N_11178,N_11247);
nand U11480 (N_11480,N_11182,N_11127);
nand U11481 (N_11481,N_11319,N_11259);
xnor U11482 (N_11482,N_11346,N_11361);
nand U11483 (N_11483,N_11383,N_11157);
nor U11484 (N_11484,N_11133,N_11117);
and U11485 (N_11485,N_11195,N_11185);
or U11486 (N_11486,N_11143,N_11142);
xnor U11487 (N_11487,N_11237,N_11263);
or U11488 (N_11488,N_11265,N_11317);
nor U11489 (N_11489,N_11343,N_11141);
or U11490 (N_11490,N_11277,N_11224);
or U11491 (N_11491,N_11137,N_11173);
xor U11492 (N_11492,N_11191,N_11357);
nor U11493 (N_11493,N_11328,N_11216);
nor U11494 (N_11494,N_11278,N_11304);
nor U11495 (N_11495,N_11348,N_11359);
nor U11496 (N_11496,N_11392,N_11192);
or U11497 (N_11497,N_11288,N_11229);
nor U11498 (N_11498,N_11186,N_11261);
nor U11499 (N_11499,N_11347,N_11197);
or U11500 (N_11500,N_11378,N_11118);
and U11501 (N_11501,N_11184,N_11332);
or U11502 (N_11502,N_11112,N_11146);
or U11503 (N_11503,N_11116,N_11274);
xor U11504 (N_11504,N_11353,N_11335);
xor U11505 (N_11505,N_11105,N_11300);
nor U11506 (N_11506,N_11231,N_11211);
xor U11507 (N_11507,N_11154,N_11108);
nand U11508 (N_11508,N_11139,N_11388);
or U11509 (N_11509,N_11124,N_11327);
xor U11510 (N_11510,N_11280,N_11251);
nand U11511 (N_11511,N_11169,N_11355);
or U11512 (N_11512,N_11109,N_11167);
xnor U11513 (N_11513,N_11239,N_11352);
nor U11514 (N_11514,N_11221,N_11198);
nand U11515 (N_11515,N_11119,N_11325);
or U11516 (N_11516,N_11255,N_11372);
xor U11517 (N_11517,N_11200,N_11390);
or U11518 (N_11518,N_11339,N_11384);
nand U11519 (N_11519,N_11158,N_11360);
xor U11520 (N_11520,N_11156,N_11382);
nor U11521 (N_11521,N_11163,N_11212);
or U11522 (N_11522,N_11254,N_11226);
xnor U11523 (N_11523,N_11151,N_11381);
nor U11524 (N_11524,N_11162,N_11236);
and U11525 (N_11525,N_11330,N_11220);
or U11526 (N_11526,N_11207,N_11333);
nor U11527 (N_11527,N_11205,N_11269);
and U11528 (N_11528,N_11102,N_11190);
nand U11529 (N_11529,N_11371,N_11329);
nand U11530 (N_11530,N_11311,N_11318);
nand U11531 (N_11531,N_11228,N_11123);
nor U11532 (N_11532,N_11358,N_11249);
nor U11533 (N_11533,N_11313,N_11245);
and U11534 (N_11534,N_11241,N_11310);
nor U11535 (N_11535,N_11103,N_11267);
and U11536 (N_11536,N_11366,N_11106);
nand U11537 (N_11537,N_11376,N_11345);
xnor U11538 (N_11538,N_11210,N_11285);
nand U11539 (N_11539,N_11316,N_11144);
nand U11540 (N_11540,N_11183,N_11148);
xor U11541 (N_11541,N_11131,N_11273);
xnor U11542 (N_11542,N_11338,N_11380);
nand U11543 (N_11543,N_11256,N_11174);
nor U11544 (N_11544,N_11290,N_11309);
nand U11545 (N_11545,N_11132,N_11218);
or U11546 (N_11546,N_11230,N_11172);
xor U11547 (N_11547,N_11396,N_11179);
and U11548 (N_11548,N_11397,N_11225);
xnor U11549 (N_11549,N_11326,N_11286);
nor U11550 (N_11550,N_11273,N_11356);
or U11551 (N_11551,N_11244,N_11313);
nand U11552 (N_11552,N_11261,N_11195);
nand U11553 (N_11553,N_11138,N_11387);
nand U11554 (N_11554,N_11202,N_11248);
and U11555 (N_11555,N_11163,N_11309);
xnor U11556 (N_11556,N_11361,N_11158);
nor U11557 (N_11557,N_11228,N_11244);
nor U11558 (N_11558,N_11139,N_11338);
and U11559 (N_11559,N_11161,N_11250);
nor U11560 (N_11560,N_11178,N_11326);
or U11561 (N_11561,N_11205,N_11252);
nand U11562 (N_11562,N_11315,N_11250);
nor U11563 (N_11563,N_11136,N_11109);
xor U11564 (N_11564,N_11305,N_11396);
xnor U11565 (N_11565,N_11182,N_11203);
nor U11566 (N_11566,N_11346,N_11102);
or U11567 (N_11567,N_11310,N_11127);
and U11568 (N_11568,N_11125,N_11117);
nor U11569 (N_11569,N_11295,N_11123);
or U11570 (N_11570,N_11386,N_11197);
nand U11571 (N_11571,N_11248,N_11167);
nor U11572 (N_11572,N_11224,N_11164);
or U11573 (N_11573,N_11152,N_11293);
nand U11574 (N_11574,N_11358,N_11112);
nor U11575 (N_11575,N_11398,N_11359);
or U11576 (N_11576,N_11206,N_11348);
or U11577 (N_11577,N_11158,N_11180);
nor U11578 (N_11578,N_11347,N_11221);
xnor U11579 (N_11579,N_11336,N_11369);
nand U11580 (N_11580,N_11145,N_11252);
nand U11581 (N_11581,N_11196,N_11281);
nand U11582 (N_11582,N_11208,N_11116);
xnor U11583 (N_11583,N_11131,N_11277);
nor U11584 (N_11584,N_11127,N_11301);
and U11585 (N_11585,N_11106,N_11302);
nor U11586 (N_11586,N_11229,N_11302);
and U11587 (N_11587,N_11379,N_11265);
nand U11588 (N_11588,N_11255,N_11293);
xor U11589 (N_11589,N_11219,N_11354);
nand U11590 (N_11590,N_11185,N_11332);
and U11591 (N_11591,N_11292,N_11103);
xnor U11592 (N_11592,N_11321,N_11275);
or U11593 (N_11593,N_11278,N_11119);
nor U11594 (N_11594,N_11331,N_11370);
and U11595 (N_11595,N_11361,N_11275);
or U11596 (N_11596,N_11255,N_11106);
xnor U11597 (N_11597,N_11162,N_11322);
or U11598 (N_11598,N_11193,N_11337);
nand U11599 (N_11599,N_11246,N_11165);
nand U11600 (N_11600,N_11175,N_11204);
nand U11601 (N_11601,N_11307,N_11232);
nand U11602 (N_11602,N_11248,N_11336);
nand U11603 (N_11603,N_11198,N_11356);
xor U11604 (N_11604,N_11129,N_11376);
nor U11605 (N_11605,N_11286,N_11202);
or U11606 (N_11606,N_11118,N_11296);
nand U11607 (N_11607,N_11347,N_11228);
nand U11608 (N_11608,N_11309,N_11262);
or U11609 (N_11609,N_11359,N_11295);
and U11610 (N_11610,N_11243,N_11264);
and U11611 (N_11611,N_11114,N_11166);
nor U11612 (N_11612,N_11146,N_11398);
or U11613 (N_11613,N_11170,N_11211);
or U11614 (N_11614,N_11202,N_11334);
xor U11615 (N_11615,N_11370,N_11119);
or U11616 (N_11616,N_11197,N_11269);
or U11617 (N_11617,N_11368,N_11265);
and U11618 (N_11618,N_11298,N_11152);
or U11619 (N_11619,N_11338,N_11337);
and U11620 (N_11620,N_11290,N_11389);
xnor U11621 (N_11621,N_11201,N_11273);
nand U11622 (N_11622,N_11229,N_11121);
xor U11623 (N_11623,N_11393,N_11235);
and U11624 (N_11624,N_11188,N_11195);
nand U11625 (N_11625,N_11217,N_11168);
nand U11626 (N_11626,N_11170,N_11121);
xor U11627 (N_11627,N_11202,N_11310);
nor U11628 (N_11628,N_11309,N_11343);
and U11629 (N_11629,N_11195,N_11271);
nand U11630 (N_11630,N_11233,N_11319);
or U11631 (N_11631,N_11270,N_11277);
and U11632 (N_11632,N_11335,N_11293);
xnor U11633 (N_11633,N_11266,N_11278);
and U11634 (N_11634,N_11235,N_11139);
xnor U11635 (N_11635,N_11154,N_11279);
and U11636 (N_11636,N_11248,N_11239);
xor U11637 (N_11637,N_11111,N_11300);
nor U11638 (N_11638,N_11292,N_11383);
and U11639 (N_11639,N_11380,N_11152);
nor U11640 (N_11640,N_11124,N_11325);
xnor U11641 (N_11641,N_11304,N_11149);
or U11642 (N_11642,N_11314,N_11115);
xnor U11643 (N_11643,N_11326,N_11352);
nor U11644 (N_11644,N_11187,N_11392);
xor U11645 (N_11645,N_11308,N_11207);
nand U11646 (N_11646,N_11253,N_11157);
nor U11647 (N_11647,N_11393,N_11144);
xnor U11648 (N_11648,N_11108,N_11132);
xnor U11649 (N_11649,N_11353,N_11375);
nor U11650 (N_11650,N_11216,N_11293);
nor U11651 (N_11651,N_11187,N_11369);
xor U11652 (N_11652,N_11281,N_11253);
and U11653 (N_11653,N_11329,N_11113);
nor U11654 (N_11654,N_11210,N_11264);
and U11655 (N_11655,N_11342,N_11328);
nor U11656 (N_11656,N_11374,N_11395);
nor U11657 (N_11657,N_11141,N_11193);
or U11658 (N_11658,N_11396,N_11174);
nor U11659 (N_11659,N_11103,N_11225);
nor U11660 (N_11660,N_11361,N_11246);
nor U11661 (N_11661,N_11101,N_11164);
and U11662 (N_11662,N_11312,N_11131);
nand U11663 (N_11663,N_11226,N_11320);
xor U11664 (N_11664,N_11149,N_11378);
or U11665 (N_11665,N_11231,N_11310);
nor U11666 (N_11666,N_11195,N_11320);
xor U11667 (N_11667,N_11146,N_11340);
and U11668 (N_11668,N_11298,N_11176);
or U11669 (N_11669,N_11241,N_11194);
and U11670 (N_11670,N_11344,N_11316);
or U11671 (N_11671,N_11156,N_11286);
xor U11672 (N_11672,N_11335,N_11232);
nor U11673 (N_11673,N_11232,N_11109);
and U11674 (N_11674,N_11330,N_11373);
nand U11675 (N_11675,N_11383,N_11318);
or U11676 (N_11676,N_11255,N_11222);
nor U11677 (N_11677,N_11175,N_11264);
nand U11678 (N_11678,N_11140,N_11114);
and U11679 (N_11679,N_11250,N_11341);
xnor U11680 (N_11680,N_11193,N_11106);
nand U11681 (N_11681,N_11124,N_11329);
and U11682 (N_11682,N_11176,N_11312);
nand U11683 (N_11683,N_11195,N_11116);
nor U11684 (N_11684,N_11225,N_11294);
nor U11685 (N_11685,N_11100,N_11226);
nor U11686 (N_11686,N_11115,N_11173);
nand U11687 (N_11687,N_11259,N_11261);
and U11688 (N_11688,N_11243,N_11384);
or U11689 (N_11689,N_11234,N_11140);
nand U11690 (N_11690,N_11350,N_11358);
xnor U11691 (N_11691,N_11285,N_11192);
nor U11692 (N_11692,N_11130,N_11390);
nand U11693 (N_11693,N_11296,N_11237);
xnor U11694 (N_11694,N_11165,N_11223);
xnor U11695 (N_11695,N_11187,N_11339);
or U11696 (N_11696,N_11306,N_11333);
or U11697 (N_11697,N_11173,N_11306);
or U11698 (N_11698,N_11377,N_11382);
nor U11699 (N_11699,N_11173,N_11337);
and U11700 (N_11700,N_11669,N_11569);
nor U11701 (N_11701,N_11557,N_11577);
and U11702 (N_11702,N_11612,N_11457);
and U11703 (N_11703,N_11451,N_11613);
nor U11704 (N_11704,N_11578,N_11606);
nand U11705 (N_11705,N_11592,N_11506);
xor U11706 (N_11706,N_11473,N_11629);
nor U11707 (N_11707,N_11534,N_11658);
nand U11708 (N_11708,N_11548,N_11401);
and U11709 (N_11709,N_11581,N_11424);
and U11710 (N_11710,N_11545,N_11660);
nor U11711 (N_11711,N_11443,N_11491);
or U11712 (N_11712,N_11617,N_11677);
nor U11713 (N_11713,N_11483,N_11511);
xnor U11714 (N_11714,N_11422,N_11566);
nand U11715 (N_11715,N_11406,N_11410);
nand U11716 (N_11716,N_11648,N_11529);
and U11717 (N_11717,N_11670,N_11697);
and U11718 (N_11718,N_11650,N_11567);
xor U11719 (N_11719,N_11453,N_11607);
and U11720 (N_11720,N_11468,N_11503);
and U11721 (N_11721,N_11447,N_11530);
nor U11722 (N_11722,N_11643,N_11633);
nor U11723 (N_11723,N_11458,N_11667);
and U11724 (N_11724,N_11501,N_11591);
nor U11725 (N_11725,N_11590,N_11425);
xor U11726 (N_11726,N_11456,N_11573);
xnor U11727 (N_11727,N_11652,N_11408);
and U11728 (N_11728,N_11657,N_11549);
and U11729 (N_11729,N_11662,N_11626);
or U11730 (N_11730,N_11693,N_11507);
or U11731 (N_11731,N_11547,N_11498);
or U11732 (N_11732,N_11680,N_11684);
and U11733 (N_11733,N_11464,N_11698);
nand U11734 (N_11734,N_11647,N_11435);
and U11735 (N_11735,N_11686,N_11450);
xnor U11736 (N_11736,N_11655,N_11654);
or U11737 (N_11737,N_11563,N_11687);
nor U11738 (N_11738,N_11430,N_11565);
or U11739 (N_11739,N_11681,N_11604);
nand U11740 (N_11740,N_11514,N_11505);
or U11741 (N_11741,N_11672,N_11575);
or U11742 (N_11742,N_11632,N_11452);
or U11743 (N_11743,N_11585,N_11608);
and U11744 (N_11744,N_11615,N_11555);
nand U11745 (N_11745,N_11520,N_11642);
and U11746 (N_11746,N_11644,N_11560);
nand U11747 (N_11747,N_11470,N_11572);
or U11748 (N_11748,N_11689,N_11409);
nand U11749 (N_11749,N_11683,N_11533);
nor U11750 (N_11750,N_11441,N_11415);
and U11751 (N_11751,N_11546,N_11480);
and U11752 (N_11752,N_11664,N_11517);
and U11753 (N_11753,N_11428,N_11541);
nand U11754 (N_11754,N_11436,N_11500);
xnor U11755 (N_11755,N_11671,N_11544);
nand U11756 (N_11756,N_11571,N_11419);
and U11757 (N_11757,N_11601,N_11513);
and U11758 (N_11758,N_11602,N_11434);
nor U11759 (N_11759,N_11521,N_11597);
or U11760 (N_11760,N_11476,N_11663);
or U11761 (N_11761,N_11414,N_11561);
nor U11762 (N_11762,N_11696,N_11463);
nor U11763 (N_11763,N_11499,N_11487);
nor U11764 (N_11764,N_11600,N_11543);
or U11765 (N_11765,N_11678,N_11484);
nor U11766 (N_11766,N_11651,N_11446);
nand U11767 (N_11767,N_11646,N_11522);
nand U11768 (N_11768,N_11502,N_11694);
or U11769 (N_11769,N_11627,N_11586);
nor U11770 (N_11770,N_11445,N_11466);
or U11771 (N_11771,N_11442,N_11588);
nor U11772 (N_11772,N_11564,N_11595);
or U11773 (N_11773,N_11489,N_11695);
nand U11774 (N_11774,N_11598,N_11417);
xnor U11775 (N_11775,N_11559,N_11661);
nor U11776 (N_11776,N_11637,N_11471);
nand U11777 (N_11777,N_11492,N_11594);
xor U11778 (N_11778,N_11461,N_11550);
nor U11779 (N_11779,N_11455,N_11512);
or U11780 (N_11780,N_11481,N_11459);
nor U11781 (N_11781,N_11411,N_11412);
xnor U11782 (N_11782,N_11616,N_11494);
or U11783 (N_11783,N_11413,N_11485);
or U11784 (N_11784,N_11465,N_11558);
nor U11785 (N_11785,N_11580,N_11416);
and U11786 (N_11786,N_11574,N_11621);
and U11787 (N_11787,N_11508,N_11475);
nor U11788 (N_11788,N_11685,N_11431);
xnor U11789 (N_11789,N_11478,N_11504);
and U11790 (N_11790,N_11582,N_11403);
nor U11791 (N_11791,N_11609,N_11634);
nor U11792 (N_11792,N_11688,N_11493);
nand U11793 (N_11793,N_11407,N_11674);
or U11794 (N_11794,N_11526,N_11649);
and U11795 (N_11795,N_11477,N_11554);
nor U11796 (N_11796,N_11538,N_11474);
and U11797 (N_11797,N_11444,N_11552);
nand U11798 (N_11798,N_11614,N_11659);
or U11799 (N_11799,N_11418,N_11583);
nand U11800 (N_11800,N_11528,N_11625);
or U11801 (N_11801,N_11482,N_11620);
and U11802 (N_11802,N_11535,N_11439);
and U11803 (N_11803,N_11656,N_11469);
xnor U11804 (N_11804,N_11562,N_11635);
nand U11805 (N_11805,N_11449,N_11675);
nor U11806 (N_11806,N_11679,N_11454);
nor U11807 (N_11807,N_11579,N_11427);
or U11808 (N_11808,N_11486,N_11515);
and U11809 (N_11809,N_11542,N_11692);
nand U11810 (N_11810,N_11537,N_11599);
and U11811 (N_11811,N_11699,N_11467);
nand U11812 (N_11812,N_11518,N_11429);
xor U11813 (N_11813,N_11432,N_11666);
and U11814 (N_11814,N_11639,N_11527);
or U11815 (N_11815,N_11532,N_11460);
xor U11816 (N_11816,N_11593,N_11570);
or U11817 (N_11817,N_11653,N_11676);
nand U11818 (N_11818,N_11525,N_11531);
nor U11819 (N_11819,N_11603,N_11400);
xor U11820 (N_11820,N_11519,N_11509);
xor U11821 (N_11821,N_11495,N_11631);
nand U11822 (N_11822,N_11618,N_11553);
nor U11823 (N_11823,N_11691,N_11539);
xor U11824 (N_11824,N_11423,N_11665);
or U11825 (N_11825,N_11540,N_11426);
and U11826 (N_11826,N_11605,N_11623);
and U11827 (N_11827,N_11420,N_11630);
and U11828 (N_11828,N_11433,N_11440);
xnor U11829 (N_11829,N_11437,N_11497);
nand U11830 (N_11830,N_11690,N_11496);
xnor U11831 (N_11831,N_11536,N_11556);
nand U11832 (N_11832,N_11438,N_11472);
nand U11833 (N_11833,N_11584,N_11619);
xor U11834 (N_11834,N_11479,N_11405);
nand U11835 (N_11835,N_11523,N_11462);
xor U11836 (N_11836,N_11589,N_11404);
nor U11837 (N_11837,N_11448,N_11587);
or U11838 (N_11838,N_11524,N_11402);
or U11839 (N_11839,N_11596,N_11610);
and U11840 (N_11840,N_11645,N_11622);
nor U11841 (N_11841,N_11636,N_11488);
xnor U11842 (N_11842,N_11638,N_11421);
nand U11843 (N_11843,N_11673,N_11641);
nand U11844 (N_11844,N_11551,N_11510);
and U11845 (N_11845,N_11568,N_11628);
nor U11846 (N_11846,N_11682,N_11611);
and U11847 (N_11847,N_11640,N_11624);
nor U11848 (N_11848,N_11668,N_11490);
nor U11849 (N_11849,N_11516,N_11576);
xor U11850 (N_11850,N_11414,N_11514);
or U11851 (N_11851,N_11614,N_11552);
nand U11852 (N_11852,N_11425,N_11648);
and U11853 (N_11853,N_11482,N_11543);
nor U11854 (N_11854,N_11671,N_11611);
nand U11855 (N_11855,N_11432,N_11490);
nor U11856 (N_11856,N_11476,N_11622);
or U11857 (N_11857,N_11556,N_11461);
xnor U11858 (N_11858,N_11590,N_11621);
or U11859 (N_11859,N_11538,N_11475);
xor U11860 (N_11860,N_11676,N_11626);
xor U11861 (N_11861,N_11624,N_11539);
and U11862 (N_11862,N_11548,N_11696);
nand U11863 (N_11863,N_11492,N_11482);
or U11864 (N_11864,N_11540,N_11508);
and U11865 (N_11865,N_11573,N_11607);
and U11866 (N_11866,N_11461,N_11641);
nand U11867 (N_11867,N_11669,N_11548);
xnor U11868 (N_11868,N_11637,N_11631);
or U11869 (N_11869,N_11563,N_11537);
or U11870 (N_11870,N_11534,N_11545);
nor U11871 (N_11871,N_11658,N_11432);
nand U11872 (N_11872,N_11431,N_11520);
nor U11873 (N_11873,N_11611,N_11441);
nor U11874 (N_11874,N_11488,N_11635);
nand U11875 (N_11875,N_11429,N_11699);
nor U11876 (N_11876,N_11476,N_11445);
nor U11877 (N_11877,N_11633,N_11618);
xnor U11878 (N_11878,N_11689,N_11537);
xor U11879 (N_11879,N_11678,N_11602);
nand U11880 (N_11880,N_11403,N_11465);
nor U11881 (N_11881,N_11505,N_11691);
nor U11882 (N_11882,N_11668,N_11494);
nand U11883 (N_11883,N_11667,N_11512);
or U11884 (N_11884,N_11418,N_11570);
xnor U11885 (N_11885,N_11586,N_11522);
or U11886 (N_11886,N_11597,N_11617);
or U11887 (N_11887,N_11432,N_11462);
nor U11888 (N_11888,N_11569,N_11457);
nor U11889 (N_11889,N_11469,N_11663);
nand U11890 (N_11890,N_11613,N_11646);
nor U11891 (N_11891,N_11489,N_11531);
and U11892 (N_11892,N_11607,N_11472);
or U11893 (N_11893,N_11541,N_11572);
or U11894 (N_11894,N_11657,N_11615);
and U11895 (N_11895,N_11652,N_11606);
nand U11896 (N_11896,N_11503,N_11553);
or U11897 (N_11897,N_11655,N_11602);
or U11898 (N_11898,N_11428,N_11523);
nor U11899 (N_11899,N_11505,N_11601);
nand U11900 (N_11900,N_11522,N_11470);
and U11901 (N_11901,N_11674,N_11444);
nand U11902 (N_11902,N_11596,N_11698);
xor U11903 (N_11903,N_11435,N_11637);
or U11904 (N_11904,N_11692,N_11442);
nand U11905 (N_11905,N_11567,N_11522);
xor U11906 (N_11906,N_11443,N_11469);
nor U11907 (N_11907,N_11612,N_11429);
nor U11908 (N_11908,N_11483,N_11671);
nor U11909 (N_11909,N_11674,N_11499);
nor U11910 (N_11910,N_11430,N_11543);
nand U11911 (N_11911,N_11628,N_11433);
nor U11912 (N_11912,N_11496,N_11525);
nand U11913 (N_11913,N_11465,N_11421);
and U11914 (N_11914,N_11602,N_11536);
nor U11915 (N_11915,N_11451,N_11531);
or U11916 (N_11916,N_11546,N_11664);
and U11917 (N_11917,N_11675,N_11647);
nand U11918 (N_11918,N_11645,N_11447);
xnor U11919 (N_11919,N_11509,N_11450);
xor U11920 (N_11920,N_11494,N_11651);
xor U11921 (N_11921,N_11420,N_11493);
nand U11922 (N_11922,N_11421,N_11552);
nand U11923 (N_11923,N_11571,N_11690);
or U11924 (N_11924,N_11557,N_11612);
nor U11925 (N_11925,N_11450,N_11530);
nand U11926 (N_11926,N_11598,N_11539);
or U11927 (N_11927,N_11612,N_11588);
nor U11928 (N_11928,N_11523,N_11602);
nand U11929 (N_11929,N_11680,N_11458);
nand U11930 (N_11930,N_11625,N_11437);
xor U11931 (N_11931,N_11544,N_11690);
and U11932 (N_11932,N_11579,N_11432);
and U11933 (N_11933,N_11595,N_11475);
or U11934 (N_11934,N_11644,N_11547);
nor U11935 (N_11935,N_11575,N_11401);
or U11936 (N_11936,N_11428,N_11417);
and U11937 (N_11937,N_11458,N_11677);
nand U11938 (N_11938,N_11447,N_11647);
nor U11939 (N_11939,N_11561,N_11628);
or U11940 (N_11940,N_11440,N_11417);
xnor U11941 (N_11941,N_11658,N_11421);
or U11942 (N_11942,N_11439,N_11401);
or U11943 (N_11943,N_11607,N_11699);
nor U11944 (N_11944,N_11608,N_11450);
or U11945 (N_11945,N_11602,N_11438);
nand U11946 (N_11946,N_11424,N_11567);
or U11947 (N_11947,N_11522,N_11539);
nand U11948 (N_11948,N_11517,N_11641);
nor U11949 (N_11949,N_11552,N_11537);
xnor U11950 (N_11950,N_11421,N_11445);
and U11951 (N_11951,N_11441,N_11462);
xnor U11952 (N_11952,N_11666,N_11572);
nand U11953 (N_11953,N_11648,N_11636);
nand U11954 (N_11954,N_11547,N_11699);
nor U11955 (N_11955,N_11453,N_11447);
or U11956 (N_11956,N_11444,N_11551);
or U11957 (N_11957,N_11444,N_11660);
nor U11958 (N_11958,N_11646,N_11660);
xnor U11959 (N_11959,N_11594,N_11477);
xnor U11960 (N_11960,N_11621,N_11539);
nor U11961 (N_11961,N_11479,N_11415);
xnor U11962 (N_11962,N_11618,N_11467);
and U11963 (N_11963,N_11661,N_11487);
and U11964 (N_11964,N_11466,N_11489);
xor U11965 (N_11965,N_11437,N_11695);
nand U11966 (N_11966,N_11429,N_11459);
or U11967 (N_11967,N_11686,N_11469);
or U11968 (N_11968,N_11600,N_11462);
nand U11969 (N_11969,N_11545,N_11656);
nor U11970 (N_11970,N_11522,N_11690);
or U11971 (N_11971,N_11487,N_11519);
and U11972 (N_11972,N_11476,N_11478);
nand U11973 (N_11973,N_11527,N_11442);
and U11974 (N_11974,N_11656,N_11562);
and U11975 (N_11975,N_11450,N_11572);
nor U11976 (N_11976,N_11437,N_11587);
and U11977 (N_11977,N_11506,N_11523);
and U11978 (N_11978,N_11401,N_11580);
or U11979 (N_11979,N_11558,N_11529);
nand U11980 (N_11980,N_11571,N_11531);
or U11981 (N_11981,N_11489,N_11541);
xor U11982 (N_11982,N_11582,N_11648);
or U11983 (N_11983,N_11608,N_11506);
nor U11984 (N_11984,N_11445,N_11681);
nand U11985 (N_11985,N_11672,N_11509);
or U11986 (N_11986,N_11446,N_11623);
and U11987 (N_11987,N_11689,N_11621);
nor U11988 (N_11988,N_11660,N_11669);
or U11989 (N_11989,N_11679,N_11559);
or U11990 (N_11990,N_11424,N_11646);
and U11991 (N_11991,N_11661,N_11672);
nor U11992 (N_11992,N_11611,N_11657);
nor U11993 (N_11993,N_11672,N_11549);
xor U11994 (N_11994,N_11680,N_11547);
or U11995 (N_11995,N_11444,N_11490);
nor U11996 (N_11996,N_11563,N_11604);
nor U11997 (N_11997,N_11524,N_11426);
and U11998 (N_11998,N_11465,N_11568);
or U11999 (N_11999,N_11604,N_11694);
or U12000 (N_12000,N_11774,N_11837);
nand U12001 (N_12001,N_11757,N_11885);
nor U12002 (N_12002,N_11854,N_11945);
xor U12003 (N_12003,N_11781,N_11735);
nor U12004 (N_12004,N_11943,N_11921);
and U12005 (N_12005,N_11908,N_11881);
and U12006 (N_12006,N_11722,N_11828);
or U12007 (N_12007,N_11800,N_11851);
nor U12008 (N_12008,N_11724,N_11756);
nor U12009 (N_12009,N_11845,N_11790);
and U12010 (N_12010,N_11821,N_11794);
nor U12011 (N_12011,N_11751,N_11743);
nand U12012 (N_12012,N_11916,N_11905);
or U12013 (N_12013,N_11780,N_11817);
xnor U12014 (N_12014,N_11831,N_11806);
nand U12015 (N_12015,N_11720,N_11913);
nor U12016 (N_12016,N_11844,N_11951);
and U12017 (N_12017,N_11996,N_11969);
nand U12018 (N_12018,N_11804,N_11795);
and U12019 (N_12019,N_11852,N_11737);
and U12020 (N_12020,N_11771,N_11787);
or U12021 (N_12021,N_11746,N_11853);
or U12022 (N_12022,N_11857,N_11792);
xnor U12023 (N_12023,N_11727,N_11712);
xor U12024 (N_12024,N_11814,N_11975);
or U12025 (N_12025,N_11865,N_11917);
nand U12026 (N_12026,N_11728,N_11875);
xor U12027 (N_12027,N_11726,N_11891);
nand U12028 (N_12028,N_11923,N_11990);
and U12029 (N_12029,N_11983,N_11822);
nand U12030 (N_12030,N_11938,N_11732);
nand U12031 (N_12031,N_11770,N_11887);
xnor U12032 (N_12032,N_11997,N_11892);
or U12033 (N_12033,N_11898,N_11879);
nand U12034 (N_12034,N_11877,N_11918);
and U12035 (N_12035,N_11717,N_11729);
nand U12036 (N_12036,N_11830,N_11721);
nand U12037 (N_12037,N_11723,N_11848);
or U12038 (N_12038,N_11762,N_11931);
or U12039 (N_12039,N_11902,N_11736);
nand U12040 (N_12040,N_11791,N_11974);
nor U12041 (N_12041,N_11798,N_11953);
xor U12042 (N_12042,N_11840,N_11987);
or U12043 (N_12043,N_11763,N_11827);
nand U12044 (N_12044,N_11705,N_11964);
nand U12045 (N_12045,N_11961,N_11759);
xnor U12046 (N_12046,N_11777,N_11888);
xor U12047 (N_12047,N_11883,N_11928);
xnor U12048 (N_12048,N_11776,N_11930);
nor U12049 (N_12049,N_11878,N_11950);
xor U12050 (N_12050,N_11716,N_11764);
nor U12051 (N_12051,N_11899,N_11977);
nor U12052 (N_12052,N_11909,N_11819);
xor U12053 (N_12053,N_11934,N_11957);
xnor U12054 (N_12054,N_11906,N_11785);
nor U12055 (N_12055,N_11850,N_11940);
or U12056 (N_12056,N_11755,N_11709);
nor U12057 (N_12057,N_11895,N_11733);
nand U12058 (N_12058,N_11882,N_11978);
xnor U12059 (N_12059,N_11788,N_11972);
nand U12060 (N_12060,N_11894,N_11939);
or U12061 (N_12061,N_11784,N_11839);
nor U12062 (N_12062,N_11803,N_11719);
and U12063 (N_12063,N_11861,N_11867);
xor U12064 (N_12064,N_11946,N_11838);
or U12065 (N_12065,N_11775,N_11963);
xnor U12066 (N_12066,N_11872,N_11903);
and U12067 (N_12067,N_11933,N_11980);
or U12068 (N_12068,N_11904,N_11932);
nor U12069 (N_12069,N_11876,N_11749);
and U12070 (N_12070,N_11818,N_11949);
or U12071 (N_12071,N_11842,N_11911);
xor U12072 (N_12072,N_11998,N_11740);
and U12073 (N_12073,N_11710,N_11893);
xnor U12074 (N_12074,N_11741,N_11846);
or U12075 (N_12075,N_11880,N_11968);
nor U12076 (N_12076,N_11952,N_11807);
or U12077 (N_12077,N_11915,N_11772);
nor U12078 (N_12078,N_11907,N_11748);
xor U12079 (N_12079,N_11973,N_11805);
nor U12080 (N_12080,N_11919,N_11707);
nand U12081 (N_12081,N_11948,N_11958);
xor U12082 (N_12082,N_11860,N_11797);
nand U12083 (N_12083,N_11959,N_11991);
xnor U12084 (N_12084,N_11873,N_11808);
nor U12085 (N_12085,N_11912,N_11761);
nand U12086 (N_12086,N_11970,N_11967);
nand U12087 (N_12087,N_11981,N_11855);
nand U12088 (N_12088,N_11793,N_11706);
nand U12089 (N_12089,N_11947,N_11823);
nor U12090 (N_12090,N_11703,N_11896);
or U12091 (N_12091,N_11701,N_11927);
xor U12092 (N_12092,N_11976,N_11809);
and U12093 (N_12093,N_11936,N_11935);
nor U12094 (N_12094,N_11825,N_11941);
nor U12095 (N_12095,N_11779,N_11816);
nor U12096 (N_12096,N_11834,N_11944);
and U12097 (N_12097,N_11783,N_11812);
xnor U12098 (N_12098,N_11955,N_11714);
xor U12099 (N_12099,N_11835,N_11815);
and U12100 (N_12100,N_11868,N_11889);
xnor U12101 (N_12101,N_11826,N_11901);
and U12102 (N_12102,N_11747,N_11989);
and U12103 (N_12103,N_11995,N_11802);
nor U12104 (N_12104,N_11862,N_11739);
and U12105 (N_12105,N_11994,N_11859);
nor U12106 (N_12106,N_11811,N_11965);
nor U12107 (N_12107,N_11897,N_11870);
nand U12108 (N_12108,N_11884,N_11926);
nand U12109 (N_12109,N_11874,N_11786);
and U12110 (N_12110,N_11988,N_11773);
or U12111 (N_12111,N_11758,N_11769);
or U12112 (N_12112,N_11801,N_11864);
and U12113 (N_12113,N_11704,N_11982);
and U12114 (N_12114,N_11843,N_11718);
xnor U12115 (N_12115,N_11760,N_11778);
or U12116 (N_12116,N_11824,N_11954);
xor U12117 (N_12117,N_11734,N_11753);
nand U12118 (N_12118,N_11813,N_11890);
and U12119 (N_12119,N_11922,N_11929);
or U12120 (N_12120,N_11702,N_11979);
nand U12121 (N_12121,N_11789,N_11956);
nand U12122 (N_12122,N_11820,N_11829);
nor U12123 (N_12123,N_11836,N_11715);
nand U12124 (N_12124,N_11925,N_11869);
nand U12125 (N_12125,N_11708,N_11871);
xor U12126 (N_12126,N_11768,N_11832);
nand U12127 (N_12127,N_11752,N_11984);
and U12128 (N_12128,N_11750,N_11900);
or U12129 (N_12129,N_11910,N_11863);
nand U12130 (N_12130,N_11986,N_11742);
nand U12131 (N_12131,N_11847,N_11937);
and U12132 (N_12132,N_11866,N_11886);
nand U12133 (N_12133,N_11914,N_11754);
or U12134 (N_12134,N_11993,N_11731);
nor U12135 (N_12135,N_11744,N_11725);
or U12136 (N_12136,N_11738,N_11810);
nand U12137 (N_12137,N_11730,N_11833);
or U12138 (N_12138,N_11765,N_11858);
nor U12139 (N_12139,N_11942,N_11920);
xnor U12140 (N_12140,N_11856,N_11962);
nor U12141 (N_12141,N_11924,N_11796);
xnor U12142 (N_12142,N_11841,N_11971);
nand U12143 (N_12143,N_11960,N_11985);
nand U12144 (N_12144,N_11766,N_11849);
xnor U12145 (N_12145,N_11799,N_11711);
nor U12146 (N_12146,N_11767,N_11999);
nor U12147 (N_12147,N_11700,N_11713);
nor U12148 (N_12148,N_11782,N_11966);
nor U12149 (N_12149,N_11745,N_11992);
nor U12150 (N_12150,N_11895,N_11841);
xnor U12151 (N_12151,N_11797,N_11904);
nand U12152 (N_12152,N_11893,N_11812);
xor U12153 (N_12153,N_11993,N_11850);
nand U12154 (N_12154,N_11758,N_11892);
and U12155 (N_12155,N_11741,N_11724);
and U12156 (N_12156,N_11745,N_11808);
and U12157 (N_12157,N_11748,N_11988);
or U12158 (N_12158,N_11872,N_11951);
and U12159 (N_12159,N_11868,N_11780);
or U12160 (N_12160,N_11977,N_11805);
xor U12161 (N_12161,N_11926,N_11956);
xnor U12162 (N_12162,N_11706,N_11771);
nor U12163 (N_12163,N_11918,N_11825);
and U12164 (N_12164,N_11894,N_11748);
nand U12165 (N_12165,N_11946,N_11929);
nor U12166 (N_12166,N_11874,N_11776);
nand U12167 (N_12167,N_11928,N_11817);
and U12168 (N_12168,N_11890,N_11771);
xnor U12169 (N_12169,N_11860,N_11710);
nand U12170 (N_12170,N_11952,N_11930);
and U12171 (N_12171,N_11943,N_11746);
and U12172 (N_12172,N_11844,N_11773);
and U12173 (N_12173,N_11837,N_11816);
or U12174 (N_12174,N_11936,N_11755);
nor U12175 (N_12175,N_11927,N_11952);
and U12176 (N_12176,N_11998,N_11761);
nor U12177 (N_12177,N_11707,N_11751);
xor U12178 (N_12178,N_11956,N_11787);
or U12179 (N_12179,N_11830,N_11704);
nor U12180 (N_12180,N_11793,N_11844);
nand U12181 (N_12181,N_11871,N_11918);
or U12182 (N_12182,N_11757,N_11844);
nor U12183 (N_12183,N_11729,N_11993);
or U12184 (N_12184,N_11884,N_11917);
nor U12185 (N_12185,N_11868,N_11878);
nand U12186 (N_12186,N_11760,N_11969);
nand U12187 (N_12187,N_11814,N_11830);
xnor U12188 (N_12188,N_11733,N_11957);
and U12189 (N_12189,N_11753,N_11970);
and U12190 (N_12190,N_11814,N_11957);
and U12191 (N_12191,N_11893,N_11970);
xor U12192 (N_12192,N_11886,N_11732);
nor U12193 (N_12193,N_11730,N_11942);
nor U12194 (N_12194,N_11850,N_11797);
nand U12195 (N_12195,N_11821,N_11925);
nor U12196 (N_12196,N_11994,N_11975);
nor U12197 (N_12197,N_11994,N_11894);
and U12198 (N_12198,N_11830,N_11941);
nor U12199 (N_12199,N_11887,N_11778);
nand U12200 (N_12200,N_11761,N_11749);
or U12201 (N_12201,N_11744,N_11964);
nand U12202 (N_12202,N_11722,N_11959);
nor U12203 (N_12203,N_11988,N_11990);
xor U12204 (N_12204,N_11952,N_11946);
and U12205 (N_12205,N_11786,N_11752);
nand U12206 (N_12206,N_11857,N_11919);
or U12207 (N_12207,N_11795,N_11790);
and U12208 (N_12208,N_11805,N_11817);
and U12209 (N_12209,N_11947,N_11859);
xor U12210 (N_12210,N_11745,N_11836);
xor U12211 (N_12211,N_11718,N_11810);
nand U12212 (N_12212,N_11980,N_11704);
xor U12213 (N_12213,N_11811,N_11890);
and U12214 (N_12214,N_11977,N_11929);
and U12215 (N_12215,N_11935,N_11849);
nor U12216 (N_12216,N_11863,N_11768);
and U12217 (N_12217,N_11723,N_11793);
and U12218 (N_12218,N_11853,N_11986);
and U12219 (N_12219,N_11747,N_11821);
xor U12220 (N_12220,N_11929,N_11913);
nor U12221 (N_12221,N_11919,N_11991);
or U12222 (N_12222,N_11828,N_11909);
and U12223 (N_12223,N_11874,N_11986);
nor U12224 (N_12224,N_11831,N_11985);
xor U12225 (N_12225,N_11719,N_11839);
xor U12226 (N_12226,N_11801,N_11810);
or U12227 (N_12227,N_11731,N_11853);
nand U12228 (N_12228,N_11810,N_11701);
or U12229 (N_12229,N_11929,N_11885);
or U12230 (N_12230,N_11810,N_11958);
nor U12231 (N_12231,N_11849,N_11941);
or U12232 (N_12232,N_11780,N_11933);
or U12233 (N_12233,N_11931,N_11747);
nor U12234 (N_12234,N_11744,N_11915);
xnor U12235 (N_12235,N_11732,N_11891);
xor U12236 (N_12236,N_11889,N_11761);
nand U12237 (N_12237,N_11731,N_11700);
and U12238 (N_12238,N_11794,N_11702);
and U12239 (N_12239,N_11934,N_11917);
and U12240 (N_12240,N_11927,N_11733);
xnor U12241 (N_12241,N_11903,N_11733);
and U12242 (N_12242,N_11870,N_11862);
and U12243 (N_12243,N_11731,N_11918);
nand U12244 (N_12244,N_11864,N_11828);
xor U12245 (N_12245,N_11783,N_11952);
or U12246 (N_12246,N_11798,N_11920);
nand U12247 (N_12247,N_11765,N_11995);
nand U12248 (N_12248,N_11851,N_11947);
and U12249 (N_12249,N_11943,N_11743);
or U12250 (N_12250,N_11843,N_11967);
and U12251 (N_12251,N_11928,N_11891);
and U12252 (N_12252,N_11714,N_11871);
nor U12253 (N_12253,N_11727,N_11902);
nand U12254 (N_12254,N_11839,N_11707);
nor U12255 (N_12255,N_11999,N_11893);
and U12256 (N_12256,N_11992,N_11982);
nand U12257 (N_12257,N_11963,N_11958);
nor U12258 (N_12258,N_11783,N_11928);
xnor U12259 (N_12259,N_11825,N_11998);
or U12260 (N_12260,N_11873,N_11779);
or U12261 (N_12261,N_11757,N_11766);
xor U12262 (N_12262,N_11811,N_11917);
nor U12263 (N_12263,N_11765,N_11799);
xnor U12264 (N_12264,N_11825,N_11880);
xor U12265 (N_12265,N_11700,N_11873);
and U12266 (N_12266,N_11715,N_11725);
nand U12267 (N_12267,N_11777,N_11825);
nor U12268 (N_12268,N_11740,N_11784);
nand U12269 (N_12269,N_11819,N_11740);
and U12270 (N_12270,N_11849,N_11925);
nand U12271 (N_12271,N_11781,N_11918);
xor U12272 (N_12272,N_11885,N_11719);
nand U12273 (N_12273,N_11884,N_11861);
or U12274 (N_12274,N_11721,N_11942);
or U12275 (N_12275,N_11841,N_11972);
nand U12276 (N_12276,N_11740,N_11995);
or U12277 (N_12277,N_11781,N_11772);
or U12278 (N_12278,N_11991,N_11797);
and U12279 (N_12279,N_11754,N_11880);
nor U12280 (N_12280,N_11988,N_11841);
or U12281 (N_12281,N_11937,N_11732);
nor U12282 (N_12282,N_11723,N_11808);
xnor U12283 (N_12283,N_11971,N_11883);
and U12284 (N_12284,N_11886,N_11898);
and U12285 (N_12285,N_11740,N_11746);
nand U12286 (N_12286,N_11907,N_11727);
nand U12287 (N_12287,N_11816,N_11825);
nor U12288 (N_12288,N_11990,N_11780);
or U12289 (N_12289,N_11914,N_11851);
xnor U12290 (N_12290,N_11951,N_11927);
xnor U12291 (N_12291,N_11915,N_11858);
nor U12292 (N_12292,N_11954,N_11706);
nor U12293 (N_12293,N_11728,N_11759);
nor U12294 (N_12294,N_11799,N_11953);
nor U12295 (N_12295,N_11791,N_11793);
nand U12296 (N_12296,N_11764,N_11920);
nand U12297 (N_12297,N_11784,N_11702);
xnor U12298 (N_12298,N_11999,N_11911);
or U12299 (N_12299,N_11928,N_11943);
and U12300 (N_12300,N_12145,N_12213);
nor U12301 (N_12301,N_12017,N_12214);
xor U12302 (N_12302,N_12279,N_12246);
nor U12303 (N_12303,N_12066,N_12171);
and U12304 (N_12304,N_12060,N_12273);
nand U12305 (N_12305,N_12035,N_12108);
or U12306 (N_12306,N_12129,N_12204);
and U12307 (N_12307,N_12100,N_12192);
or U12308 (N_12308,N_12120,N_12174);
nor U12309 (N_12309,N_12103,N_12125);
xnor U12310 (N_12310,N_12218,N_12052);
and U12311 (N_12311,N_12118,N_12201);
or U12312 (N_12312,N_12111,N_12098);
nand U12313 (N_12313,N_12211,N_12028);
xnor U12314 (N_12314,N_12141,N_12297);
xnor U12315 (N_12315,N_12245,N_12123);
xor U12316 (N_12316,N_12269,N_12180);
or U12317 (N_12317,N_12217,N_12185);
and U12318 (N_12318,N_12278,N_12262);
or U12319 (N_12319,N_12264,N_12203);
xor U12320 (N_12320,N_12073,N_12070);
xor U12321 (N_12321,N_12265,N_12105);
nand U12322 (N_12322,N_12075,N_12189);
or U12323 (N_12323,N_12226,N_12092);
nor U12324 (N_12324,N_12164,N_12050);
or U12325 (N_12325,N_12181,N_12222);
and U12326 (N_12326,N_12021,N_12179);
xnor U12327 (N_12327,N_12280,N_12132);
and U12328 (N_12328,N_12078,N_12064);
nor U12329 (N_12329,N_12239,N_12095);
nand U12330 (N_12330,N_12253,N_12063);
and U12331 (N_12331,N_12102,N_12295);
or U12332 (N_12332,N_12133,N_12143);
or U12333 (N_12333,N_12029,N_12061);
nand U12334 (N_12334,N_12209,N_12229);
nor U12335 (N_12335,N_12270,N_12291);
xor U12336 (N_12336,N_12298,N_12151);
or U12337 (N_12337,N_12207,N_12072);
or U12338 (N_12338,N_12008,N_12031);
and U12339 (N_12339,N_12002,N_12137);
or U12340 (N_12340,N_12080,N_12085);
nand U12341 (N_12341,N_12289,N_12210);
and U12342 (N_12342,N_12274,N_12041);
and U12343 (N_12343,N_12160,N_12152);
or U12344 (N_12344,N_12071,N_12172);
nor U12345 (N_12345,N_12161,N_12249);
or U12346 (N_12346,N_12094,N_12110);
nand U12347 (N_12347,N_12112,N_12290);
or U12348 (N_12348,N_12130,N_12099);
nor U12349 (N_12349,N_12169,N_12251);
and U12350 (N_12350,N_12055,N_12142);
or U12351 (N_12351,N_12084,N_12195);
and U12352 (N_12352,N_12022,N_12089);
nor U12353 (N_12353,N_12104,N_12106);
nor U12354 (N_12354,N_12252,N_12275);
nand U12355 (N_12355,N_12288,N_12149);
nor U12356 (N_12356,N_12013,N_12039);
nor U12357 (N_12357,N_12230,N_12173);
xnor U12358 (N_12358,N_12096,N_12233);
xnor U12359 (N_12359,N_12266,N_12244);
and U12360 (N_12360,N_12247,N_12199);
nor U12361 (N_12361,N_12018,N_12260);
nand U12362 (N_12362,N_12101,N_12225);
nor U12363 (N_12363,N_12194,N_12007);
or U12364 (N_12364,N_12258,N_12037);
xor U12365 (N_12365,N_12208,N_12285);
xor U12366 (N_12366,N_12198,N_12016);
nand U12367 (N_12367,N_12126,N_12234);
or U12368 (N_12368,N_12147,N_12042);
nor U12369 (N_12369,N_12184,N_12034);
nor U12370 (N_12370,N_12062,N_12281);
nor U12371 (N_12371,N_12267,N_12032);
nor U12372 (N_12372,N_12020,N_12231);
nand U12373 (N_12373,N_12187,N_12107);
nand U12374 (N_12374,N_12023,N_12003);
and U12375 (N_12375,N_12237,N_12068);
nand U12376 (N_12376,N_12083,N_12122);
and U12377 (N_12377,N_12215,N_12188);
or U12378 (N_12378,N_12248,N_12162);
xnor U12379 (N_12379,N_12144,N_12046);
or U12380 (N_12380,N_12012,N_12116);
xnor U12381 (N_12381,N_12283,N_12119);
nand U12382 (N_12382,N_12284,N_12165);
or U12383 (N_12383,N_12205,N_12190);
xor U12384 (N_12384,N_12044,N_12131);
nor U12385 (N_12385,N_12088,N_12287);
xor U12386 (N_12386,N_12001,N_12158);
or U12387 (N_12387,N_12150,N_12293);
nor U12388 (N_12388,N_12069,N_12256);
xor U12389 (N_12389,N_12182,N_12154);
and U12390 (N_12390,N_12250,N_12134);
nand U12391 (N_12391,N_12036,N_12196);
xnor U12392 (N_12392,N_12065,N_12240);
nor U12393 (N_12393,N_12155,N_12216);
nor U12394 (N_12394,N_12047,N_12059);
or U12395 (N_12395,N_12033,N_12043);
or U12396 (N_12396,N_12236,N_12159);
nand U12397 (N_12397,N_12000,N_12235);
or U12398 (N_12398,N_12051,N_12221);
nor U12399 (N_12399,N_12191,N_12128);
nor U12400 (N_12400,N_12049,N_12079);
or U12401 (N_12401,N_12139,N_12272);
nor U12402 (N_12402,N_12257,N_12170);
nor U12403 (N_12403,N_12058,N_12296);
or U12404 (N_12404,N_12186,N_12014);
xor U12405 (N_12405,N_12136,N_12294);
and U12406 (N_12406,N_12193,N_12299);
nand U12407 (N_12407,N_12027,N_12268);
nand U12408 (N_12408,N_12163,N_12114);
nand U12409 (N_12409,N_12200,N_12153);
or U12410 (N_12410,N_12263,N_12271);
nor U12411 (N_12411,N_12282,N_12081);
xnor U12412 (N_12412,N_12030,N_12220);
and U12413 (N_12413,N_12140,N_12146);
or U12414 (N_12414,N_12025,N_12053);
nand U12415 (N_12415,N_12238,N_12086);
nand U12416 (N_12416,N_12168,N_12261);
and U12417 (N_12417,N_12019,N_12056);
and U12418 (N_12418,N_12045,N_12048);
or U12419 (N_12419,N_12157,N_12135);
or U12420 (N_12420,N_12006,N_12010);
xnor U12421 (N_12421,N_12227,N_12156);
nor U12422 (N_12422,N_12026,N_12219);
nand U12423 (N_12423,N_12166,N_12167);
xnor U12424 (N_12424,N_12024,N_12067);
and U12425 (N_12425,N_12206,N_12183);
nand U12426 (N_12426,N_12243,N_12212);
xnor U12427 (N_12427,N_12255,N_12277);
nand U12428 (N_12428,N_12057,N_12004);
and U12429 (N_12429,N_12109,N_12074);
nor U12430 (N_12430,N_12113,N_12148);
or U12431 (N_12431,N_12259,N_12276);
or U12432 (N_12432,N_12228,N_12090);
nor U12433 (N_12433,N_12009,N_12076);
nand U12434 (N_12434,N_12121,N_12242);
nand U12435 (N_12435,N_12175,N_12011);
nor U12436 (N_12436,N_12087,N_12115);
nand U12437 (N_12437,N_12197,N_12178);
xnor U12438 (N_12438,N_12124,N_12292);
or U12439 (N_12439,N_12176,N_12177);
nand U12440 (N_12440,N_12202,N_12241);
nand U12441 (N_12441,N_12117,N_12286);
xor U12442 (N_12442,N_12097,N_12054);
nor U12443 (N_12443,N_12005,N_12077);
and U12444 (N_12444,N_12223,N_12127);
nand U12445 (N_12445,N_12254,N_12138);
or U12446 (N_12446,N_12082,N_12038);
or U12447 (N_12447,N_12232,N_12015);
nand U12448 (N_12448,N_12093,N_12091);
nand U12449 (N_12449,N_12224,N_12040);
and U12450 (N_12450,N_12224,N_12153);
or U12451 (N_12451,N_12110,N_12237);
xor U12452 (N_12452,N_12036,N_12165);
xnor U12453 (N_12453,N_12106,N_12156);
nor U12454 (N_12454,N_12182,N_12153);
or U12455 (N_12455,N_12162,N_12155);
nor U12456 (N_12456,N_12061,N_12013);
and U12457 (N_12457,N_12107,N_12101);
xnor U12458 (N_12458,N_12204,N_12047);
nor U12459 (N_12459,N_12150,N_12243);
nor U12460 (N_12460,N_12173,N_12062);
xnor U12461 (N_12461,N_12178,N_12174);
nor U12462 (N_12462,N_12192,N_12082);
and U12463 (N_12463,N_12012,N_12020);
nor U12464 (N_12464,N_12140,N_12239);
nand U12465 (N_12465,N_12141,N_12170);
xor U12466 (N_12466,N_12000,N_12150);
and U12467 (N_12467,N_12097,N_12291);
and U12468 (N_12468,N_12186,N_12156);
or U12469 (N_12469,N_12075,N_12130);
or U12470 (N_12470,N_12121,N_12255);
or U12471 (N_12471,N_12289,N_12202);
and U12472 (N_12472,N_12072,N_12270);
and U12473 (N_12473,N_12001,N_12253);
nor U12474 (N_12474,N_12080,N_12160);
or U12475 (N_12475,N_12158,N_12039);
and U12476 (N_12476,N_12259,N_12236);
nor U12477 (N_12477,N_12177,N_12149);
and U12478 (N_12478,N_12221,N_12056);
xnor U12479 (N_12479,N_12217,N_12063);
and U12480 (N_12480,N_12014,N_12051);
nor U12481 (N_12481,N_12177,N_12280);
nand U12482 (N_12482,N_12184,N_12276);
nand U12483 (N_12483,N_12209,N_12153);
or U12484 (N_12484,N_12130,N_12132);
nand U12485 (N_12485,N_12283,N_12273);
nor U12486 (N_12486,N_12180,N_12025);
or U12487 (N_12487,N_12089,N_12257);
nand U12488 (N_12488,N_12003,N_12058);
and U12489 (N_12489,N_12018,N_12072);
or U12490 (N_12490,N_12097,N_12107);
xnor U12491 (N_12491,N_12208,N_12094);
nand U12492 (N_12492,N_12268,N_12189);
nor U12493 (N_12493,N_12231,N_12043);
or U12494 (N_12494,N_12034,N_12264);
and U12495 (N_12495,N_12067,N_12278);
nand U12496 (N_12496,N_12133,N_12238);
or U12497 (N_12497,N_12226,N_12257);
and U12498 (N_12498,N_12125,N_12053);
and U12499 (N_12499,N_12012,N_12208);
or U12500 (N_12500,N_12127,N_12207);
nor U12501 (N_12501,N_12035,N_12111);
nor U12502 (N_12502,N_12086,N_12125);
or U12503 (N_12503,N_12256,N_12210);
and U12504 (N_12504,N_12052,N_12190);
nand U12505 (N_12505,N_12142,N_12180);
nor U12506 (N_12506,N_12061,N_12213);
nand U12507 (N_12507,N_12129,N_12174);
nor U12508 (N_12508,N_12082,N_12054);
or U12509 (N_12509,N_12197,N_12124);
or U12510 (N_12510,N_12283,N_12122);
or U12511 (N_12511,N_12117,N_12238);
nor U12512 (N_12512,N_12013,N_12233);
nand U12513 (N_12513,N_12011,N_12221);
nor U12514 (N_12514,N_12255,N_12167);
nand U12515 (N_12515,N_12280,N_12053);
and U12516 (N_12516,N_12152,N_12271);
nand U12517 (N_12517,N_12231,N_12132);
and U12518 (N_12518,N_12290,N_12161);
xnor U12519 (N_12519,N_12040,N_12199);
or U12520 (N_12520,N_12120,N_12198);
nand U12521 (N_12521,N_12284,N_12207);
or U12522 (N_12522,N_12052,N_12061);
xor U12523 (N_12523,N_12099,N_12086);
or U12524 (N_12524,N_12216,N_12123);
and U12525 (N_12525,N_12210,N_12051);
nand U12526 (N_12526,N_12224,N_12286);
xor U12527 (N_12527,N_12080,N_12059);
or U12528 (N_12528,N_12133,N_12214);
nor U12529 (N_12529,N_12257,N_12268);
nand U12530 (N_12530,N_12124,N_12207);
or U12531 (N_12531,N_12298,N_12288);
xnor U12532 (N_12532,N_12004,N_12021);
nand U12533 (N_12533,N_12284,N_12179);
nor U12534 (N_12534,N_12226,N_12254);
xor U12535 (N_12535,N_12090,N_12221);
and U12536 (N_12536,N_12099,N_12088);
or U12537 (N_12537,N_12148,N_12183);
xor U12538 (N_12538,N_12075,N_12246);
nand U12539 (N_12539,N_12178,N_12017);
nor U12540 (N_12540,N_12089,N_12194);
xnor U12541 (N_12541,N_12225,N_12131);
or U12542 (N_12542,N_12294,N_12081);
or U12543 (N_12543,N_12063,N_12110);
xor U12544 (N_12544,N_12265,N_12078);
or U12545 (N_12545,N_12161,N_12150);
and U12546 (N_12546,N_12129,N_12010);
or U12547 (N_12547,N_12054,N_12288);
nor U12548 (N_12548,N_12028,N_12138);
and U12549 (N_12549,N_12257,N_12098);
xor U12550 (N_12550,N_12234,N_12172);
xor U12551 (N_12551,N_12105,N_12095);
nand U12552 (N_12552,N_12139,N_12173);
nor U12553 (N_12553,N_12186,N_12059);
nor U12554 (N_12554,N_12141,N_12104);
or U12555 (N_12555,N_12185,N_12270);
xnor U12556 (N_12556,N_12093,N_12098);
xor U12557 (N_12557,N_12296,N_12035);
nand U12558 (N_12558,N_12127,N_12171);
xor U12559 (N_12559,N_12163,N_12047);
nor U12560 (N_12560,N_12217,N_12097);
nand U12561 (N_12561,N_12223,N_12049);
or U12562 (N_12562,N_12289,N_12180);
nand U12563 (N_12563,N_12153,N_12045);
nand U12564 (N_12564,N_12056,N_12126);
xnor U12565 (N_12565,N_12222,N_12196);
xnor U12566 (N_12566,N_12072,N_12296);
and U12567 (N_12567,N_12120,N_12002);
xnor U12568 (N_12568,N_12148,N_12193);
and U12569 (N_12569,N_12248,N_12229);
nand U12570 (N_12570,N_12166,N_12159);
and U12571 (N_12571,N_12199,N_12104);
nor U12572 (N_12572,N_12283,N_12159);
and U12573 (N_12573,N_12010,N_12025);
or U12574 (N_12574,N_12019,N_12115);
nand U12575 (N_12575,N_12124,N_12188);
nor U12576 (N_12576,N_12014,N_12231);
xor U12577 (N_12577,N_12221,N_12194);
or U12578 (N_12578,N_12063,N_12208);
nand U12579 (N_12579,N_12103,N_12035);
nor U12580 (N_12580,N_12172,N_12026);
and U12581 (N_12581,N_12205,N_12204);
nor U12582 (N_12582,N_12009,N_12075);
or U12583 (N_12583,N_12019,N_12052);
nand U12584 (N_12584,N_12027,N_12100);
nand U12585 (N_12585,N_12073,N_12020);
and U12586 (N_12586,N_12082,N_12295);
nand U12587 (N_12587,N_12232,N_12251);
or U12588 (N_12588,N_12229,N_12156);
xor U12589 (N_12589,N_12294,N_12064);
nor U12590 (N_12590,N_12189,N_12069);
xor U12591 (N_12591,N_12250,N_12151);
or U12592 (N_12592,N_12144,N_12241);
and U12593 (N_12593,N_12049,N_12173);
nand U12594 (N_12594,N_12197,N_12291);
nor U12595 (N_12595,N_12066,N_12164);
or U12596 (N_12596,N_12057,N_12221);
or U12597 (N_12597,N_12239,N_12154);
nand U12598 (N_12598,N_12278,N_12283);
nand U12599 (N_12599,N_12149,N_12245);
and U12600 (N_12600,N_12579,N_12480);
xor U12601 (N_12601,N_12568,N_12461);
nor U12602 (N_12602,N_12352,N_12322);
and U12603 (N_12603,N_12479,N_12306);
nand U12604 (N_12604,N_12563,N_12391);
and U12605 (N_12605,N_12462,N_12452);
or U12606 (N_12606,N_12587,N_12443);
or U12607 (N_12607,N_12403,N_12485);
and U12608 (N_12608,N_12504,N_12341);
or U12609 (N_12609,N_12456,N_12405);
xnor U12610 (N_12610,N_12440,N_12390);
and U12611 (N_12611,N_12399,N_12408);
nor U12612 (N_12612,N_12376,N_12509);
nor U12613 (N_12613,N_12401,N_12330);
nor U12614 (N_12614,N_12539,N_12372);
nand U12615 (N_12615,N_12374,N_12355);
xor U12616 (N_12616,N_12492,N_12394);
nor U12617 (N_12617,N_12474,N_12549);
and U12618 (N_12618,N_12476,N_12547);
and U12619 (N_12619,N_12418,N_12560);
and U12620 (N_12620,N_12530,N_12422);
or U12621 (N_12621,N_12397,N_12375);
and U12622 (N_12622,N_12531,N_12446);
and U12623 (N_12623,N_12385,N_12337);
xor U12624 (N_12624,N_12455,N_12566);
or U12625 (N_12625,N_12594,N_12545);
and U12626 (N_12626,N_12410,N_12544);
and U12627 (N_12627,N_12536,N_12491);
nand U12628 (N_12628,N_12597,N_12535);
xor U12629 (N_12629,N_12356,N_12570);
and U12630 (N_12630,N_12578,N_12468);
nor U12631 (N_12631,N_12467,N_12518);
nand U12632 (N_12632,N_12522,N_12436);
nand U12633 (N_12633,N_12327,N_12500);
nand U12634 (N_12634,N_12379,N_12409);
or U12635 (N_12635,N_12414,N_12498);
or U12636 (N_12636,N_12321,N_12473);
and U12637 (N_12637,N_12359,N_12325);
xor U12638 (N_12638,N_12438,N_12300);
xor U12639 (N_12639,N_12433,N_12360);
nor U12640 (N_12640,N_12377,N_12373);
and U12641 (N_12641,N_12353,N_12576);
nand U12642 (N_12642,N_12302,N_12329);
and U12643 (N_12643,N_12411,N_12534);
nand U12644 (N_12644,N_12543,N_12551);
or U12645 (N_12645,N_12542,N_12464);
or U12646 (N_12646,N_12524,N_12590);
xor U12647 (N_12647,N_12494,N_12515);
nor U12648 (N_12648,N_12471,N_12582);
xnor U12649 (N_12649,N_12589,N_12523);
or U12650 (N_12650,N_12413,N_12386);
nand U12651 (N_12651,N_12315,N_12525);
or U12652 (N_12652,N_12301,N_12393);
nand U12653 (N_12653,N_12310,N_12529);
nand U12654 (N_12654,N_12585,N_12312);
xnor U12655 (N_12655,N_12361,N_12593);
nor U12656 (N_12656,N_12490,N_12305);
nor U12657 (N_12657,N_12338,N_12351);
nor U12658 (N_12658,N_12477,N_12415);
and U12659 (N_12659,N_12557,N_12437);
xnor U12660 (N_12660,N_12483,N_12388);
or U12661 (N_12661,N_12546,N_12572);
and U12662 (N_12662,N_12526,N_12513);
nand U12663 (N_12663,N_12404,N_12577);
xor U12664 (N_12664,N_12345,N_12482);
or U12665 (N_12665,N_12458,N_12512);
nand U12666 (N_12666,N_12333,N_12307);
nand U12667 (N_12667,N_12407,N_12441);
nor U12668 (N_12668,N_12334,N_12516);
nor U12669 (N_12669,N_12431,N_12478);
or U12670 (N_12670,N_12313,N_12466);
and U12671 (N_12671,N_12571,N_12495);
nand U12672 (N_12672,N_12424,N_12396);
or U12673 (N_12673,N_12517,N_12487);
and U12674 (N_12674,N_12331,N_12430);
or U12675 (N_12675,N_12496,N_12323);
or U12676 (N_12676,N_12412,N_12470);
xnor U12677 (N_12677,N_12506,N_12574);
xor U12678 (N_12678,N_12583,N_12527);
xor U12679 (N_12679,N_12421,N_12335);
nand U12680 (N_12680,N_12488,N_12340);
nor U12681 (N_12681,N_12383,N_12580);
and U12682 (N_12682,N_12416,N_12511);
nand U12683 (N_12683,N_12584,N_12465);
nand U12684 (N_12684,N_12556,N_12540);
nor U12685 (N_12685,N_12548,N_12521);
and U12686 (N_12686,N_12592,N_12532);
or U12687 (N_12687,N_12533,N_12426);
nand U12688 (N_12688,N_12550,N_12309);
and U12689 (N_12689,N_12384,N_12481);
nand U12690 (N_12690,N_12505,N_12469);
nand U12691 (N_12691,N_12514,N_12339);
and U12692 (N_12692,N_12448,N_12559);
nand U12693 (N_12693,N_12567,N_12552);
xor U12694 (N_12694,N_12528,N_12596);
nor U12695 (N_12695,N_12395,N_12304);
xor U12696 (N_12696,N_12303,N_12538);
or U12697 (N_12697,N_12346,N_12499);
or U12698 (N_12698,N_12387,N_12365);
nand U12699 (N_12699,N_12502,N_12595);
and U12700 (N_12700,N_12459,N_12564);
or U12701 (N_12701,N_12308,N_12501);
xor U12702 (N_12702,N_12370,N_12445);
or U12703 (N_12703,N_12439,N_12316);
xnor U12704 (N_12704,N_12588,N_12454);
and U12705 (N_12705,N_12489,N_12573);
nor U12706 (N_12706,N_12555,N_12510);
nand U12707 (N_12707,N_12349,N_12311);
or U12708 (N_12708,N_12475,N_12432);
nand U12709 (N_12709,N_12558,N_12493);
or U12710 (N_12710,N_12347,N_12402);
nor U12711 (N_12711,N_12363,N_12314);
xor U12712 (N_12712,N_12503,N_12581);
or U12713 (N_12713,N_12507,N_12371);
nand U12714 (N_12714,N_12447,N_12423);
and U12715 (N_12715,N_12541,N_12451);
xor U12716 (N_12716,N_12358,N_12324);
nor U12717 (N_12717,N_12434,N_12444);
or U12718 (N_12718,N_12326,N_12317);
nor U12719 (N_12719,N_12598,N_12389);
nand U12720 (N_12720,N_12435,N_12450);
nand U12721 (N_12721,N_12419,N_12519);
or U12722 (N_12722,N_12366,N_12417);
nand U12723 (N_12723,N_12420,N_12591);
nor U12724 (N_12724,N_12328,N_12460);
or U12725 (N_12725,N_12429,N_12553);
xor U12726 (N_12726,N_12449,N_12565);
nor U12727 (N_12727,N_12406,N_12392);
and U12728 (N_12728,N_12368,N_12364);
xor U12729 (N_12729,N_12362,N_12453);
and U12730 (N_12730,N_12320,N_12398);
nor U12731 (N_12731,N_12561,N_12484);
nor U12732 (N_12732,N_12382,N_12343);
xor U12733 (N_12733,N_12562,N_12457);
and U12734 (N_12734,N_12357,N_12427);
and U12735 (N_12735,N_12463,N_12348);
nor U12736 (N_12736,N_12425,N_12554);
and U12737 (N_12737,N_12497,N_12367);
or U12738 (N_12738,N_12442,N_12537);
nor U12739 (N_12739,N_12332,N_12354);
xnor U12740 (N_12740,N_12344,N_12508);
xnor U12741 (N_12741,N_12369,N_12380);
and U12742 (N_12742,N_12586,N_12569);
nor U12743 (N_12743,N_12319,N_12381);
or U12744 (N_12744,N_12575,N_12486);
xnor U12745 (N_12745,N_12350,N_12378);
nand U12746 (N_12746,N_12472,N_12400);
nor U12747 (N_12747,N_12520,N_12342);
nand U12748 (N_12748,N_12336,N_12599);
and U12749 (N_12749,N_12318,N_12428);
nand U12750 (N_12750,N_12438,N_12464);
or U12751 (N_12751,N_12428,N_12394);
nor U12752 (N_12752,N_12568,N_12517);
xor U12753 (N_12753,N_12490,N_12430);
xor U12754 (N_12754,N_12393,N_12413);
nor U12755 (N_12755,N_12441,N_12544);
xnor U12756 (N_12756,N_12473,N_12456);
and U12757 (N_12757,N_12336,N_12486);
and U12758 (N_12758,N_12451,N_12333);
xnor U12759 (N_12759,N_12537,N_12524);
xnor U12760 (N_12760,N_12447,N_12502);
or U12761 (N_12761,N_12431,N_12373);
xor U12762 (N_12762,N_12322,N_12365);
nor U12763 (N_12763,N_12308,N_12471);
and U12764 (N_12764,N_12397,N_12314);
and U12765 (N_12765,N_12505,N_12541);
xnor U12766 (N_12766,N_12325,N_12385);
xor U12767 (N_12767,N_12521,N_12366);
or U12768 (N_12768,N_12528,N_12443);
nand U12769 (N_12769,N_12551,N_12575);
or U12770 (N_12770,N_12404,N_12541);
and U12771 (N_12771,N_12553,N_12525);
nand U12772 (N_12772,N_12360,N_12526);
or U12773 (N_12773,N_12459,N_12494);
nand U12774 (N_12774,N_12348,N_12508);
nor U12775 (N_12775,N_12342,N_12599);
xnor U12776 (N_12776,N_12588,N_12569);
or U12777 (N_12777,N_12449,N_12506);
nand U12778 (N_12778,N_12560,N_12390);
or U12779 (N_12779,N_12468,N_12549);
xor U12780 (N_12780,N_12364,N_12485);
xnor U12781 (N_12781,N_12474,N_12571);
or U12782 (N_12782,N_12414,N_12441);
nor U12783 (N_12783,N_12499,N_12517);
nand U12784 (N_12784,N_12384,N_12327);
nor U12785 (N_12785,N_12486,N_12442);
nor U12786 (N_12786,N_12320,N_12322);
nand U12787 (N_12787,N_12382,N_12566);
nand U12788 (N_12788,N_12362,N_12573);
or U12789 (N_12789,N_12516,N_12492);
nor U12790 (N_12790,N_12381,N_12464);
nor U12791 (N_12791,N_12363,N_12323);
or U12792 (N_12792,N_12489,N_12585);
nor U12793 (N_12793,N_12363,N_12335);
nand U12794 (N_12794,N_12453,N_12363);
xnor U12795 (N_12795,N_12538,N_12498);
nand U12796 (N_12796,N_12429,N_12374);
xnor U12797 (N_12797,N_12466,N_12428);
or U12798 (N_12798,N_12597,N_12372);
and U12799 (N_12799,N_12400,N_12583);
nand U12800 (N_12800,N_12363,N_12407);
xnor U12801 (N_12801,N_12483,N_12392);
nand U12802 (N_12802,N_12327,N_12398);
nor U12803 (N_12803,N_12534,N_12450);
nand U12804 (N_12804,N_12418,N_12391);
xor U12805 (N_12805,N_12376,N_12308);
xor U12806 (N_12806,N_12353,N_12411);
nor U12807 (N_12807,N_12488,N_12368);
xor U12808 (N_12808,N_12520,N_12561);
xnor U12809 (N_12809,N_12594,N_12437);
nand U12810 (N_12810,N_12405,N_12348);
nand U12811 (N_12811,N_12591,N_12434);
nand U12812 (N_12812,N_12329,N_12359);
xor U12813 (N_12813,N_12374,N_12469);
nor U12814 (N_12814,N_12396,N_12564);
xor U12815 (N_12815,N_12484,N_12384);
or U12816 (N_12816,N_12340,N_12406);
xnor U12817 (N_12817,N_12508,N_12451);
nor U12818 (N_12818,N_12429,N_12486);
nand U12819 (N_12819,N_12498,N_12556);
nor U12820 (N_12820,N_12385,N_12321);
or U12821 (N_12821,N_12313,N_12434);
xor U12822 (N_12822,N_12534,N_12507);
or U12823 (N_12823,N_12305,N_12357);
nor U12824 (N_12824,N_12382,N_12481);
and U12825 (N_12825,N_12530,N_12473);
and U12826 (N_12826,N_12482,N_12352);
nand U12827 (N_12827,N_12505,N_12410);
nand U12828 (N_12828,N_12318,N_12350);
or U12829 (N_12829,N_12555,N_12588);
nand U12830 (N_12830,N_12321,N_12312);
nor U12831 (N_12831,N_12457,N_12525);
nor U12832 (N_12832,N_12537,N_12362);
and U12833 (N_12833,N_12323,N_12465);
nor U12834 (N_12834,N_12567,N_12430);
or U12835 (N_12835,N_12580,N_12534);
nand U12836 (N_12836,N_12330,N_12383);
and U12837 (N_12837,N_12591,N_12400);
nor U12838 (N_12838,N_12568,N_12312);
nor U12839 (N_12839,N_12579,N_12464);
or U12840 (N_12840,N_12414,N_12302);
nand U12841 (N_12841,N_12467,N_12586);
xor U12842 (N_12842,N_12398,N_12527);
nor U12843 (N_12843,N_12466,N_12491);
nor U12844 (N_12844,N_12444,N_12342);
or U12845 (N_12845,N_12521,N_12320);
nor U12846 (N_12846,N_12492,N_12520);
nor U12847 (N_12847,N_12475,N_12365);
nor U12848 (N_12848,N_12511,N_12368);
or U12849 (N_12849,N_12540,N_12448);
or U12850 (N_12850,N_12323,N_12335);
nor U12851 (N_12851,N_12320,N_12327);
or U12852 (N_12852,N_12438,N_12528);
and U12853 (N_12853,N_12455,N_12342);
nor U12854 (N_12854,N_12458,N_12454);
nand U12855 (N_12855,N_12335,N_12331);
nor U12856 (N_12856,N_12595,N_12374);
or U12857 (N_12857,N_12495,N_12556);
nand U12858 (N_12858,N_12547,N_12492);
nand U12859 (N_12859,N_12519,N_12599);
nand U12860 (N_12860,N_12383,N_12349);
or U12861 (N_12861,N_12579,N_12458);
or U12862 (N_12862,N_12376,N_12332);
xor U12863 (N_12863,N_12597,N_12499);
nor U12864 (N_12864,N_12366,N_12558);
or U12865 (N_12865,N_12471,N_12323);
or U12866 (N_12866,N_12531,N_12538);
nand U12867 (N_12867,N_12437,N_12303);
xnor U12868 (N_12868,N_12436,N_12555);
nand U12869 (N_12869,N_12515,N_12478);
xor U12870 (N_12870,N_12304,N_12487);
nand U12871 (N_12871,N_12467,N_12473);
nor U12872 (N_12872,N_12569,N_12593);
nor U12873 (N_12873,N_12556,N_12523);
nand U12874 (N_12874,N_12498,N_12402);
and U12875 (N_12875,N_12505,N_12530);
and U12876 (N_12876,N_12432,N_12533);
and U12877 (N_12877,N_12467,N_12370);
nor U12878 (N_12878,N_12381,N_12585);
and U12879 (N_12879,N_12390,N_12526);
and U12880 (N_12880,N_12554,N_12541);
nor U12881 (N_12881,N_12367,N_12363);
or U12882 (N_12882,N_12400,N_12453);
or U12883 (N_12883,N_12389,N_12443);
and U12884 (N_12884,N_12486,N_12481);
xor U12885 (N_12885,N_12535,N_12370);
xor U12886 (N_12886,N_12371,N_12566);
and U12887 (N_12887,N_12308,N_12379);
xnor U12888 (N_12888,N_12519,N_12406);
nor U12889 (N_12889,N_12498,N_12342);
and U12890 (N_12890,N_12467,N_12364);
or U12891 (N_12891,N_12516,N_12485);
and U12892 (N_12892,N_12360,N_12463);
nand U12893 (N_12893,N_12337,N_12359);
xor U12894 (N_12894,N_12382,N_12543);
nand U12895 (N_12895,N_12365,N_12418);
xnor U12896 (N_12896,N_12519,N_12398);
and U12897 (N_12897,N_12592,N_12599);
xnor U12898 (N_12898,N_12489,N_12401);
and U12899 (N_12899,N_12415,N_12427);
xnor U12900 (N_12900,N_12772,N_12761);
or U12901 (N_12901,N_12859,N_12769);
or U12902 (N_12902,N_12605,N_12610);
nand U12903 (N_12903,N_12710,N_12852);
nand U12904 (N_12904,N_12792,N_12887);
and U12905 (N_12905,N_12623,N_12816);
and U12906 (N_12906,N_12817,N_12704);
or U12907 (N_12907,N_12663,N_12835);
xnor U12908 (N_12908,N_12726,N_12602);
nand U12909 (N_12909,N_12874,N_12785);
nand U12910 (N_12910,N_12690,N_12821);
nor U12911 (N_12911,N_12834,N_12654);
xnor U12912 (N_12912,N_12880,N_12642);
and U12913 (N_12913,N_12712,N_12678);
or U12914 (N_12914,N_12809,N_12734);
and U12915 (N_12915,N_12643,N_12853);
nor U12916 (N_12916,N_12850,N_12711);
nand U12917 (N_12917,N_12617,N_12893);
nand U12918 (N_12918,N_12763,N_12742);
nor U12919 (N_12919,N_12640,N_12724);
or U12920 (N_12920,N_12787,N_12864);
nand U12921 (N_12921,N_12773,N_12798);
and U12922 (N_12922,N_12856,N_12713);
or U12923 (N_12923,N_12802,N_12737);
nand U12924 (N_12924,N_12689,N_12766);
nand U12925 (N_12925,N_12784,N_12746);
and U12926 (N_12926,N_12867,N_12825);
xor U12927 (N_12927,N_12677,N_12849);
or U12928 (N_12928,N_12673,N_12843);
nor U12929 (N_12929,N_12645,N_12614);
and U12930 (N_12930,N_12791,N_12636);
nor U12931 (N_12931,N_12708,N_12741);
xnor U12932 (N_12932,N_12679,N_12693);
nor U12933 (N_12933,N_12608,N_12718);
nor U12934 (N_12934,N_12622,N_12877);
nand U12935 (N_12935,N_12664,N_12894);
nor U12936 (N_12936,N_12889,N_12871);
xor U12937 (N_12937,N_12759,N_12793);
and U12938 (N_12938,N_12615,N_12800);
or U12939 (N_12939,N_12870,N_12682);
nand U12940 (N_12940,N_12722,N_12727);
or U12941 (N_12941,N_12669,N_12613);
nand U12942 (N_12942,N_12607,N_12804);
nor U12943 (N_12943,N_12783,N_12875);
nand U12944 (N_12944,N_12803,N_12848);
xnor U12945 (N_12945,N_12659,N_12729);
nor U12946 (N_12946,N_12801,N_12700);
xor U12947 (N_12947,N_12695,N_12829);
xor U12948 (N_12948,N_12748,N_12770);
xor U12949 (N_12949,N_12757,N_12730);
and U12950 (N_12950,N_12705,N_12827);
or U12951 (N_12951,N_12767,N_12707);
or U12952 (N_12952,N_12808,N_12671);
nor U12953 (N_12953,N_12616,N_12750);
or U12954 (N_12954,N_12658,N_12703);
nor U12955 (N_12955,N_12681,N_12650);
or U12956 (N_12956,N_12807,N_12691);
or U12957 (N_12957,N_12777,N_12628);
and U12958 (N_12958,N_12885,N_12858);
nor U12959 (N_12959,N_12812,N_12638);
or U12960 (N_12960,N_12692,N_12768);
or U12961 (N_12961,N_12644,N_12627);
and U12962 (N_12962,N_12863,N_12675);
or U12963 (N_12963,N_12831,N_12841);
xnor U12964 (N_12964,N_12882,N_12866);
xnor U12965 (N_12965,N_12646,N_12666);
and U12966 (N_12966,N_12637,N_12662);
or U12967 (N_12967,N_12779,N_12633);
or U12968 (N_12968,N_12743,N_12655);
nand U12969 (N_12969,N_12876,N_12720);
nor U12970 (N_12970,N_12795,N_12733);
nor U12971 (N_12971,N_12651,N_12665);
or U12972 (N_12972,N_12694,N_12721);
and U12973 (N_12973,N_12696,N_12776);
and U12974 (N_12974,N_12869,N_12625);
xnor U12975 (N_12975,N_12600,N_12680);
nor U12976 (N_12976,N_12714,N_12883);
xor U12977 (N_12977,N_12794,N_12676);
or U12978 (N_12978,N_12838,N_12760);
or U12979 (N_12979,N_12836,N_12815);
xnor U12980 (N_12980,N_12652,N_12753);
nor U12981 (N_12981,N_12896,N_12647);
or U12982 (N_12982,N_12629,N_12701);
nor U12983 (N_12983,N_12824,N_12612);
or U12984 (N_12984,N_12755,N_12752);
xnor U12985 (N_12985,N_12844,N_12878);
nand U12986 (N_12986,N_12745,N_12822);
and U12987 (N_12987,N_12797,N_12649);
nand U12988 (N_12988,N_12683,N_12805);
and U12989 (N_12989,N_12635,N_12846);
nand U12990 (N_12990,N_12765,N_12840);
or U12991 (N_12991,N_12719,N_12725);
nor U12992 (N_12992,N_12747,N_12660);
or U12993 (N_12993,N_12771,N_12790);
xnor U12994 (N_12994,N_12839,N_12820);
nor U12995 (N_12995,N_12728,N_12667);
or U12996 (N_12996,N_12837,N_12813);
nor U12997 (N_12997,N_12736,N_12631);
or U12998 (N_12998,N_12892,N_12786);
or U12999 (N_12999,N_12668,N_12855);
xor U13000 (N_13000,N_12653,N_12788);
nand U13001 (N_13001,N_12723,N_12685);
xnor U13002 (N_13002,N_12672,N_12632);
and U13003 (N_13003,N_12740,N_12604);
or U13004 (N_13004,N_12810,N_12754);
or U13005 (N_13005,N_12731,N_12758);
nor U13006 (N_13006,N_12620,N_12796);
nor U13007 (N_13007,N_12890,N_12897);
xnor U13008 (N_13008,N_12626,N_12670);
or U13009 (N_13009,N_12706,N_12648);
nor U13010 (N_13010,N_12847,N_12634);
nand U13011 (N_13011,N_12789,N_12899);
nand U13012 (N_13012,N_12774,N_12873);
xnor U13013 (N_13013,N_12799,N_12884);
nand U13014 (N_13014,N_12756,N_12854);
nor U13015 (N_13015,N_12661,N_12735);
nor U13016 (N_13016,N_12639,N_12656);
nor U13017 (N_13017,N_12698,N_12715);
xor U13018 (N_13018,N_12709,N_12814);
xor U13019 (N_13019,N_12739,N_12780);
xnor U13020 (N_13020,N_12879,N_12609);
and U13021 (N_13021,N_12891,N_12868);
xor U13022 (N_13022,N_12895,N_12738);
or U13023 (N_13023,N_12819,N_12699);
xor U13024 (N_13024,N_12818,N_12716);
nor U13025 (N_13025,N_12845,N_12621);
or U13026 (N_13026,N_12865,N_12697);
nor U13027 (N_13027,N_12619,N_12857);
or U13028 (N_13028,N_12872,N_12828);
and U13029 (N_13029,N_12881,N_12641);
nor U13030 (N_13030,N_12657,N_12830);
and U13031 (N_13031,N_12888,N_12611);
or U13032 (N_13032,N_12842,N_12688);
xnor U13033 (N_13033,N_12781,N_12811);
nand U13034 (N_13034,N_12832,N_12684);
or U13035 (N_13035,N_12823,N_12749);
nand U13036 (N_13036,N_12686,N_12860);
nor U13037 (N_13037,N_12886,N_12702);
nor U13038 (N_13038,N_12751,N_12833);
and U13039 (N_13039,N_12775,N_12606);
or U13040 (N_13040,N_12806,N_12861);
nor U13041 (N_13041,N_12851,N_12603);
nor U13042 (N_13042,N_12624,N_12630);
and U13043 (N_13043,N_12764,N_12618);
or U13044 (N_13044,N_12744,N_12826);
nor U13045 (N_13045,N_12782,N_12778);
nor U13046 (N_13046,N_12674,N_12898);
nand U13047 (N_13047,N_12687,N_12762);
and U13048 (N_13048,N_12601,N_12732);
xor U13049 (N_13049,N_12717,N_12862);
or U13050 (N_13050,N_12861,N_12685);
or U13051 (N_13051,N_12660,N_12692);
or U13052 (N_13052,N_12808,N_12762);
nor U13053 (N_13053,N_12752,N_12745);
or U13054 (N_13054,N_12827,N_12794);
or U13055 (N_13055,N_12801,N_12856);
xnor U13056 (N_13056,N_12756,N_12629);
nor U13057 (N_13057,N_12721,N_12850);
nor U13058 (N_13058,N_12873,N_12889);
nand U13059 (N_13059,N_12844,N_12603);
or U13060 (N_13060,N_12649,N_12698);
nor U13061 (N_13061,N_12796,N_12811);
or U13062 (N_13062,N_12796,N_12869);
or U13063 (N_13063,N_12619,N_12780);
and U13064 (N_13064,N_12657,N_12866);
nand U13065 (N_13065,N_12777,N_12850);
nand U13066 (N_13066,N_12776,N_12768);
and U13067 (N_13067,N_12637,N_12848);
nand U13068 (N_13068,N_12826,N_12652);
or U13069 (N_13069,N_12622,N_12633);
and U13070 (N_13070,N_12786,N_12689);
and U13071 (N_13071,N_12765,N_12640);
xor U13072 (N_13072,N_12790,N_12741);
nand U13073 (N_13073,N_12780,N_12793);
and U13074 (N_13074,N_12672,N_12650);
and U13075 (N_13075,N_12710,N_12657);
or U13076 (N_13076,N_12851,N_12620);
and U13077 (N_13077,N_12836,N_12715);
xor U13078 (N_13078,N_12701,N_12884);
nand U13079 (N_13079,N_12872,N_12690);
nor U13080 (N_13080,N_12846,N_12831);
nand U13081 (N_13081,N_12721,N_12606);
or U13082 (N_13082,N_12742,N_12792);
and U13083 (N_13083,N_12877,N_12860);
or U13084 (N_13084,N_12832,N_12812);
nand U13085 (N_13085,N_12764,N_12796);
xnor U13086 (N_13086,N_12855,N_12786);
nor U13087 (N_13087,N_12863,N_12652);
or U13088 (N_13088,N_12639,N_12784);
nor U13089 (N_13089,N_12878,N_12803);
xor U13090 (N_13090,N_12672,N_12653);
xnor U13091 (N_13091,N_12750,N_12891);
or U13092 (N_13092,N_12619,N_12603);
nand U13093 (N_13093,N_12816,N_12782);
or U13094 (N_13094,N_12791,N_12819);
and U13095 (N_13095,N_12885,N_12650);
or U13096 (N_13096,N_12825,N_12702);
nor U13097 (N_13097,N_12884,N_12829);
or U13098 (N_13098,N_12722,N_12830);
xor U13099 (N_13099,N_12693,N_12825);
and U13100 (N_13100,N_12781,N_12672);
or U13101 (N_13101,N_12680,N_12716);
or U13102 (N_13102,N_12724,N_12864);
or U13103 (N_13103,N_12780,N_12809);
nand U13104 (N_13104,N_12627,N_12781);
nand U13105 (N_13105,N_12850,N_12817);
nor U13106 (N_13106,N_12780,N_12830);
or U13107 (N_13107,N_12807,N_12776);
and U13108 (N_13108,N_12657,N_12707);
xnor U13109 (N_13109,N_12608,N_12742);
or U13110 (N_13110,N_12637,N_12712);
or U13111 (N_13111,N_12765,N_12760);
xnor U13112 (N_13112,N_12675,N_12745);
nand U13113 (N_13113,N_12642,N_12794);
nor U13114 (N_13114,N_12803,N_12608);
xnor U13115 (N_13115,N_12631,N_12892);
and U13116 (N_13116,N_12704,N_12649);
or U13117 (N_13117,N_12693,N_12602);
or U13118 (N_13118,N_12877,N_12737);
nor U13119 (N_13119,N_12635,N_12788);
nand U13120 (N_13120,N_12641,N_12873);
nand U13121 (N_13121,N_12851,N_12712);
nor U13122 (N_13122,N_12608,N_12776);
and U13123 (N_13123,N_12868,N_12658);
or U13124 (N_13124,N_12842,N_12696);
nand U13125 (N_13125,N_12790,N_12770);
or U13126 (N_13126,N_12751,N_12855);
nor U13127 (N_13127,N_12619,N_12703);
and U13128 (N_13128,N_12860,N_12817);
and U13129 (N_13129,N_12847,N_12709);
nand U13130 (N_13130,N_12871,N_12784);
and U13131 (N_13131,N_12739,N_12747);
nor U13132 (N_13132,N_12803,N_12798);
xnor U13133 (N_13133,N_12603,N_12733);
nand U13134 (N_13134,N_12889,N_12665);
xnor U13135 (N_13135,N_12654,N_12676);
or U13136 (N_13136,N_12776,N_12897);
and U13137 (N_13137,N_12643,N_12610);
or U13138 (N_13138,N_12683,N_12604);
or U13139 (N_13139,N_12791,N_12800);
nand U13140 (N_13140,N_12739,N_12639);
nor U13141 (N_13141,N_12680,N_12819);
xor U13142 (N_13142,N_12631,N_12862);
and U13143 (N_13143,N_12707,N_12893);
nor U13144 (N_13144,N_12736,N_12761);
and U13145 (N_13145,N_12655,N_12683);
or U13146 (N_13146,N_12861,N_12782);
xnor U13147 (N_13147,N_12768,N_12719);
and U13148 (N_13148,N_12862,N_12817);
nand U13149 (N_13149,N_12850,N_12874);
and U13150 (N_13150,N_12828,N_12861);
or U13151 (N_13151,N_12878,N_12653);
or U13152 (N_13152,N_12744,N_12668);
nand U13153 (N_13153,N_12668,N_12648);
and U13154 (N_13154,N_12853,N_12762);
nand U13155 (N_13155,N_12705,N_12685);
nor U13156 (N_13156,N_12808,N_12668);
xnor U13157 (N_13157,N_12674,N_12613);
nor U13158 (N_13158,N_12652,N_12653);
nor U13159 (N_13159,N_12857,N_12697);
nor U13160 (N_13160,N_12751,N_12749);
nor U13161 (N_13161,N_12818,N_12719);
nor U13162 (N_13162,N_12688,N_12749);
or U13163 (N_13163,N_12783,N_12863);
and U13164 (N_13164,N_12850,N_12752);
nor U13165 (N_13165,N_12834,N_12876);
and U13166 (N_13166,N_12676,N_12834);
and U13167 (N_13167,N_12738,N_12749);
or U13168 (N_13168,N_12886,N_12877);
xnor U13169 (N_13169,N_12749,N_12891);
or U13170 (N_13170,N_12893,N_12649);
xor U13171 (N_13171,N_12809,N_12719);
nand U13172 (N_13172,N_12851,N_12864);
or U13173 (N_13173,N_12609,N_12660);
xor U13174 (N_13174,N_12840,N_12838);
nor U13175 (N_13175,N_12626,N_12898);
xnor U13176 (N_13176,N_12888,N_12842);
xor U13177 (N_13177,N_12865,N_12635);
nand U13178 (N_13178,N_12878,N_12701);
nor U13179 (N_13179,N_12685,N_12715);
or U13180 (N_13180,N_12650,N_12667);
xnor U13181 (N_13181,N_12745,N_12840);
nand U13182 (N_13182,N_12704,N_12836);
or U13183 (N_13183,N_12663,N_12693);
xor U13184 (N_13184,N_12862,N_12880);
nor U13185 (N_13185,N_12885,N_12738);
or U13186 (N_13186,N_12747,N_12779);
and U13187 (N_13187,N_12647,N_12857);
xnor U13188 (N_13188,N_12752,N_12865);
and U13189 (N_13189,N_12875,N_12885);
nand U13190 (N_13190,N_12748,N_12675);
nand U13191 (N_13191,N_12855,N_12781);
and U13192 (N_13192,N_12794,N_12645);
xnor U13193 (N_13193,N_12602,N_12722);
and U13194 (N_13194,N_12689,N_12643);
nor U13195 (N_13195,N_12825,N_12647);
nand U13196 (N_13196,N_12712,N_12791);
nand U13197 (N_13197,N_12636,N_12878);
nand U13198 (N_13198,N_12673,N_12707);
nand U13199 (N_13199,N_12740,N_12889);
and U13200 (N_13200,N_12984,N_12945);
nor U13201 (N_13201,N_13005,N_13071);
xnor U13202 (N_13202,N_13149,N_13038);
nand U13203 (N_13203,N_12923,N_13126);
nand U13204 (N_13204,N_13179,N_12907);
and U13205 (N_13205,N_12971,N_13115);
and U13206 (N_13206,N_12944,N_12904);
xor U13207 (N_13207,N_13198,N_13143);
xnor U13208 (N_13208,N_12990,N_13035);
or U13209 (N_13209,N_12962,N_13014);
and U13210 (N_13210,N_13156,N_12977);
or U13211 (N_13211,N_13188,N_12974);
xnor U13212 (N_13212,N_12973,N_12909);
xor U13213 (N_13213,N_12975,N_13095);
and U13214 (N_13214,N_13090,N_13140);
xor U13215 (N_13215,N_13151,N_13022);
nand U13216 (N_13216,N_13167,N_13153);
nor U13217 (N_13217,N_13092,N_13029);
nor U13218 (N_13218,N_13015,N_13002);
or U13219 (N_13219,N_13097,N_13109);
xnor U13220 (N_13220,N_13183,N_13091);
or U13221 (N_13221,N_13073,N_13162);
nor U13222 (N_13222,N_12937,N_13016);
or U13223 (N_13223,N_12938,N_13137);
or U13224 (N_13224,N_13182,N_13021);
nand U13225 (N_13225,N_12925,N_12986);
nor U13226 (N_13226,N_13129,N_13055);
or U13227 (N_13227,N_13174,N_13061);
and U13228 (N_13228,N_13039,N_13047);
and U13229 (N_13229,N_13004,N_13003);
xnor U13230 (N_13230,N_13180,N_13168);
or U13231 (N_13231,N_13121,N_13152);
nand U13232 (N_13232,N_12956,N_13093);
or U13233 (N_13233,N_13108,N_13017);
xor U13234 (N_13234,N_13001,N_12980);
nand U13235 (N_13235,N_13146,N_13127);
nand U13236 (N_13236,N_13112,N_13135);
nor U13237 (N_13237,N_13120,N_13133);
nand U13238 (N_13238,N_13045,N_13099);
or U13239 (N_13239,N_12911,N_13128);
xnor U13240 (N_13240,N_13148,N_13125);
nand U13241 (N_13241,N_12959,N_12966);
and U13242 (N_13242,N_13010,N_12967);
and U13243 (N_13243,N_13052,N_13054);
nor U13244 (N_13244,N_13059,N_12915);
xnor U13245 (N_13245,N_12900,N_13000);
nand U13246 (N_13246,N_12935,N_13142);
nand U13247 (N_13247,N_13088,N_13175);
nor U13248 (N_13248,N_12919,N_13011);
xor U13249 (N_13249,N_13196,N_12901);
nand U13250 (N_13250,N_13170,N_12918);
nand U13251 (N_13251,N_13161,N_13110);
nand U13252 (N_13252,N_13163,N_12983);
nand U13253 (N_13253,N_12978,N_12946);
and U13254 (N_13254,N_13083,N_13104);
nor U13255 (N_13255,N_13060,N_13187);
or U13256 (N_13256,N_13186,N_13043);
or U13257 (N_13257,N_13019,N_12999);
and U13258 (N_13258,N_13193,N_12930);
nand U13259 (N_13259,N_12969,N_13114);
or U13260 (N_13260,N_13041,N_13107);
xor U13261 (N_13261,N_12991,N_12927);
nor U13262 (N_13262,N_12920,N_13036);
nand U13263 (N_13263,N_12933,N_13191);
xnor U13264 (N_13264,N_13027,N_12981);
xor U13265 (N_13265,N_13171,N_12996);
xor U13266 (N_13266,N_12957,N_13178);
xnor U13267 (N_13267,N_13176,N_12979);
nor U13268 (N_13268,N_13070,N_13145);
or U13269 (N_13269,N_12965,N_12917);
or U13270 (N_13270,N_12985,N_13199);
nand U13271 (N_13271,N_13131,N_13008);
nor U13272 (N_13272,N_12968,N_13068);
or U13273 (N_13273,N_12960,N_13119);
and U13274 (N_13274,N_13122,N_13032);
nor U13275 (N_13275,N_13160,N_12947);
nand U13276 (N_13276,N_13136,N_13013);
xor U13277 (N_13277,N_13123,N_13139);
or U13278 (N_13278,N_12972,N_12948);
nor U13279 (N_13279,N_13190,N_13177);
xor U13280 (N_13280,N_13067,N_13164);
xor U13281 (N_13281,N_13028,N_12912);
or U13282 (N_13282,N_13147,N_13165);
xnor U13283 (N_13283,N_13064,N_13025);
and U13284 (N_13284,N_12988,N_12997);
and U13285 (N_13285,N_13084,N_13144);
and U13286 (N_13286,N_13051,N_12952);
xnor U13287 (N_13287,N_13006,N_13124);
xor U13288 (N_13288,N_13081,N_12931);
or U13289 (N_13289,N_13077,N_13103);
and U13290 (N_13290,N_13046,N_13100);
and U13291 (N_13291,N_13194,N_13020);
nand U13292 (N_13292,N_13065,N_12950);
xnor U13293 (N_13293,N_13009,N_12922);
or U13294 (N_13294,N_13058,N_13101);
and U13295 (N_13295,N_12905,N_13102);
nand U13296 (N_13296,N_13111,N_13053);
nand U13297 (N_13297,N_13173,N_12961);
or U13298 (N_13298,N_13159,N_12970);
nand U13299 (N_13299,N_13072,N_13062);
nand U13300 (N_13300,N_13155,N_13057);
and U13301 (N_13301,N_13086,N_12906);
nor U13302 (N_13302,N_13116,N_12936);
nor U13303 (N_13303,N_12903,N_13181);
or U13304 (N_13304,N_13080,N_13192);
nor U13305 (N_13305,N_13158,N_12902);
nor U13306 (N_13306,N_13007,N_12934);
or U13307 (N_13307,N_12995,N_13085);
xnor U13308 (N_13308,N_12949,N_12998);
xor U13309 (N_13309,N_13018,N_12955);
xor U13310 (N_13310,N_13138,N_12908);
nor U13311 (N_13311,N_13184,N_13082);
or U13312 (N_13312,N_12943,N_13033);
or U13313 (N_13313,N_13117,N_13056);
nor U13314 (N_13314,N_13012,N_13141);
and U13315 (N_13315,N_13189,N_12982);
nor U13316 (N_13316,N_13118,N_12939);
nand U13317 (N_13317,N_12987,N_13113);
nand U13318 (N_13318,N_13066,N_13037);
or U13319 (N_13319,N_12951,N_13106);
xnor U13320 (N_13320,N_13076,N_13078);
and U13321 (N_13321,N_13150,N_12994);
and U13322 (N_13322,N_13044,N_13130);
and U13323 (N_13323,N_12954,N_12921);
and U13324 (N_13324,N_12924,N_13030);
or U13325 (N_13325,N_13094,N_12910);
nor U13326 (N_13326,N_12928,N_13048);
or U13327 (N_13327,N_13075,N_13096);
or U13328 (N_13328,N_12958,N_13087);
or U13329 (N_13329,N_12932,N_13063);
xor U13330 (N_13330,N_13105,N_13169);
nor U13331 (N_13331,N_13026,N_12914);
or U13332 (N_13332,N_12976,N_13024);
xnor U13333 (N_13333,N_13157,N_13034);
and U13334 (N_13334,N_12963,N_13074);
nand U13335 (N_13335,N_13154,N_13069);
or U13336 (N_13336,N_12989,N_13166);
and U13337 (N_13337,N_12913,N_12940);
xnor U13338 (N_13338,N_12993,N_12926);
and U13339 (N_13339,N_13049,N_13031);
nand U13340 (N_13340,N_13098,N_13040);
or U13341 (N_13341,N_13197,N_13172);
and U13342 (N_13342,N_13132,N_12992);
nor U13343 (N_13343,N_12942,N_13089);
and U13344 (N_13344,N_13042,N_13079);
xnor U13345 (N_13345,N_12964,N_12929);
or U13346 (N_13346,N_12953,N_13195);
nand U13347 (N_13347,N_13023,N_12916);
or U13348 (N_13348,N_13050,N_13185);
xor U13349 (N_13349,N_13134,N_12941);
xor U13350 (N_13350,N_13078,N_12960);
xor U13351 (N_13351,N_13056,N_13105);
and U13352 (N_13352,N_12914,N_12974);
nand U13353 (N_13353,N_13175,N_13047);
nand U13354 (N_13354,N_13045,N_13118);
nand U13355 (N_13355,N_13009,N_12952);
nand U13356 (N_13356,N_12955,N_13194);
or U13357 (N_13357,N_13041,N_13072);
or U13358 (N_13358,N_12967,N_13053);
nor U13359 (N_13359,N_13074,N_13095);
nor U13360 (N_13360,N_13040,N_13096);
xnor U13361 (N_13361,N_13146,N_13048);
xnor U13362 (N_13362,N_12966,N_13199);
xor U13363 (N_13363,N_12904,N_13114);
nor U13364 (N_13364,N_13015,N_12968);
nand U13365 (N_13365,N_12940,N_13018);
xnor U13366 (N_13366,N_12933,N_12999);
xor U13367 (N_13367,N_12917,N_12968);
nor U13368 (N_13368,N_12985,N_13061);
nand U13369 (N_13369,N_12914,N_13001);
and U13370 (N_13370,N_13089,N_12981);
or U13371 (N_13371,N_12944,N_13024);
or U13372 (N_13372,N_12962,N_13074);
nand U13373 (N_13373,N_13183,N_13076);
xor U13374 (N_13374,N_13043,N_12975);
and U13375 (N_13375,N_13031,N_12958);
nand U13376 (N_13376,N_12915,N_13081);
nor U13377 (N_13377,N_13098,N_13029);
or U13378 (N_13378,N_13096,N_13090);
and U13379 (N_13379,N_13119,N_12907);
xor U13380 (N_13380,N_12959,N_13095);
and U13381 (N_13381,N_13036,N_12988);
nor U13382 (N_13382,N_13008,N_13173);
nand U13383 (N_13383,N_12981,N_13059);
and U13384 (N_13384,N_12912,N_13065);
or U13385 (N_13385,N_13147,N_13194);
or U13386 (N_13386,N_12971,N_13088);
xor U13387 (N_13387,N_13189,N_12994);
nor U13388 (N_13388,N_12924,N_13069);
nand U13389 (N_13389,N_13130,N_13039);
nand U13390 (N_13390,N_12918,N_13126);
xnor U13391 (N_13391,N_13134,N_12950);
nor U13392 (N_13392,N_12966,N_13105);
nand U13393 (N_13393,N_13088,N_13065);
nor U13394 (N_13394,N_12915,N_13017);
nor U13395 (N_13395,N_12914,N_13061);
or U13396 (N_13396,N_12935,N_13033);
or U13397 (N_13397,N_12936,N_13010);
nor U13398 (N_13398,N_13129,N_13052);
xor U13399 (N_13399,N_13148,N_12906);
or U13400 (N_13400,N_13047,N_13032);
nor U13401 (N_13401,N_13131,N_12921);
xor U13402 (N_13402,N_13150,N_13189);
nor U13403 (N_13403,N_12996,N_13039);
nand U13404 (N_13404,N_13151,N_13020);
xnor U13405 (N_13405,N_12989,N_13138);
and U13406 (N_13406,N_13181,N_13134);
nand U13407 (N_13407,N_13187,N_13130);
and U13408 (N_13408,N_13010,N_12951);
nor U13409 (N_13409,N_12983,N_13068);
or U13410 (N_13410,N_13136,N_12976);
nor U13411 (N_13411,N_12985,N_12991);
and U13412 (N_13412,N_13120,N_13192);
nand U13413 (N_13413,N_13007,N_13017);
xor U13414 (N_13414,N_12911,N_12991);
or U13415 (N_13415,N_12973,N_13012);
and U13416 (N_13416,N_13167,N_13088);
xor U13417 (N_13417,N_13186,N_13075);
xnor U13418 (N_13418,N_12987,N_13055);
nor U13419 (N_13419,N_13151,N_13160);
xor U13420 (N_13420,N_13105,N_13092);
nor U13421 (N_13421,N_13193,N_13196);
xnor U13422 (N_13422,N_12934,N_13186);
nand U13423 (N_13423,N_13131,N_12931);
or U13424 (N_13424,N_12953,N_13105);
and U13425 (N_13425,N_12990,N_13026);
nor U13426 (N_13426,N_13100,N_12904);
xor U13427 (N_13427,N_12909,N_13112);
or U13428 (N_13428,N_13045,N_13047);
nor U13429 (N_13429,N_13050,N_12942);
xnor U13430 (N_13430,N_12984,N_13031);
nand U13431 (N_13431,N_13021,N_13193);
nor U13432 (N_13432,N_13064,N_13186);
nor U13433 (N_13433,N_13029,N_13016);
nand U13434 (N_13434,N_12974,N_13098);
nand U13435 (N_13435,N_12947,N_12967);
xnor U13436 (N_13436,N_12922,N_13032);
nor U13437 (N_13437,N_13172,N_13002);
and U13438 (N_13438,N_13157,N_13163);
nand U13439 (N_13439,N_13106,N_12945);
nor U13440 (N_13440,N_13196,N_13198);
nor U13441 (N_13441,N_13189,N_13035);
and U13442 (N_13442,N_13086,N_13199);
nor U13443 (N_13443,N_12935,N_13194);
and U13444 (N_13444,N_13100,N_13050);
nor U13445 (N_13445,N_13187,N_13087);
nor U13446 (N_13446,N_13183,N_13082);
xor U13447 (N_13447,N_13030,N_12956);
nand U13448 (N_13448,N_13127,N_12944);
nand U13449 (N_13449,N_13054,N_13079);
nand U13450 (N_13450,N_12902,N_13065);
and U13451 (N_13451,N_13136,N_12957);
xnor U13452 (N_13452,N_13000,N_13192);
and U13453 (N_13453,N_13086,N_13111);
xor U13454 (N_13454,N_13077,N_13052);
nand U13455 (N_13455,N_12923,N_12946);
and U13456 (N_13456,N_13157,N_12961);
and U13457 (N_13457,N_13190,N_13186);
or U13458 (N_13458,N_13007,N_13126);
and U13459 (N_13459,N_12986,N_13199);
nor U13460 (N_13460,N_12997,N_13017);
or U13461 (N_13461,N_13005,N_13181);
nor U13462 (N_13462,N_13044,N_13012);
xnor U13463 (N_13463,N_13197,N_13117);
xor U13464 (N_13464,N_12900,N_12961);
nand U13465 (N_13465,N_13142,N_13002);
and U13466 (N_13466,N_13088,N_12961);
xnor U13467 (N_13467,N_13145,N_13124);
xnor U13468 (N_13468,N_13031,N_13087);
xor U13469 (N_13469,N_13038,N_13144);
and U13470 (N_13470,N_13184,N_13186);
nor U13471 (N_13471,N_12905,N_13176);
nor U13472 (N_13472,N_13177,N_13030);
nor U13473 (N_13473,N_12975,N_13001);
nor U13474 (N_13474,N_13170,N_13076);
or U13475 (N_13475,N_13056,N_12964);
xor U13476 (N_13476,N_12983,N_12952);
and U13477 (N_13477,N_13083,N_12901);
and U13478 (N_13478,N_13037,N_13028);
and U13479 (N_13479,N_12943,N_13156);
and U13480 (N_13480,N_13122,N_13086);
nor U13481 (N_13481,N_13096,N_13105);
or U13482 (N_13482,N_13178,N_12974);
and U13483 (N_13483,N_13044,N_12967);
or U13484 (N_13484,N_13047,N_12954);
xnor U13485 (N_13485,N_13130,N_13111);
or U13486 (N_13486,N_13059,N_13082);
xnor U13487 (N_13487,N_13018,N_13183);
xnor U13488 (N_13488,N_13197,N_13125);
xnor U13489 (N_13489,N_13152,N_13053);
xor U13490 (N_13490,N_13006,N_13099);
nand U13491 (N_13491,N_13197,N_13074);
nor U13492 (N_13492,N_13114,N_13091);
or U13493 (N_13493,N_13061,N_13071);
nor U13494 (N_13494,N_12965,N_12916);
or U13495 (N_13495,N_13119,N_12980);
and U13496 (N_13496,N_13142,N_13196);
or U13497 (N_13497,N_12980,N_13079);
and U13498 (N_13498,N_13013,N_13139);
nand U13499 (N_13499,N_13146,N_13074);
xor U13500 (N_13500,N_13439,N_13297);
nand U13501 (N_13501,N_13448,N_13338);
nor U13502 (N_13502,N_13484,N_13246);
and U13503 (N_13503,N_13299,N_13485);
nor U13504 (N_13504,N_13455,N_13285);
or U13505 (N_13505,N_13245,N_13248);
and U13506 (N_13506,N_13301,N_13295);
nand U13507 (N_13507,N_13453,N_13426);
nand U13508 (N_13508,N_13280,N_13243);
or U13509 (N_13509,N_13257,N_13298);
and U13510 (N_13510,N_13249,N_13305);
xor U13511 (N_13511,N_13290,N_13483);
nand U13512 (N_13512,N_13364,N_13287);
xor U13513 (N_13513,N_13358,N_13202);
nor U13514 (N_13514,N_13407,N_13411);
or U13515 (N_13515,N_13401,N_13308);
and U13516 (N_13516,N_13362,N_13218);
and U13517 (N_13517,N_13209,N_13462);
and U13518 (N_13518,N_13444,N_13420);
and U13519 (N_13519,N_13342,N_13304);
or U13520 (N_13520,N_13256,N_13208);
or U13521 (N_13521,N_13387,N_13478);
nor U13522 (N_13522,N_13349,N_13355);
nand U13523 (N_13523,N_13219,N_13443);
xor U13524 (N_13524,N_13447,N_13493);
xnor U13525 (N_13525,N_13239,N_13354);
and U13526 (N_13526,N_13469,N_13470);
nor U13527 (N_13527,N_13450,N_13494);
and U13528 (N_13528,N_13212,N_13227);
or U13529 (N_13529,N_13482,N_13427);
xor U13530 (N_13530,N_13386,N_13329);
nor U13531 (N_13531,N_13288,N_13289);
and U13532 (N_13532,N_13398,N_13397);
xor U13533 (N_13533,N_13309,N_13436);
nor U13534 (N_13534,N_13492,N_13382);
xor U13535 (N_13535,N_13344,N_13331);
xor U13536 (N_13536,N_13204,N_13459);
nor U13537 (N_13537,N_13375,N_13432);
nand U13538 (N_13538,N_13381,N_13428);
or U13539 (N_13539,N_13247,N_13441);
nor U13540 (N_13540,N_13413,N_13466);
nor U13541 (N_13541,N_13489,N_13324);
and U13542 (N_13542,N_13233,N_13383);
xnor U13543 (N_13543,N_13306,N_13313);
nor U13544 (N_13544,N_13336,N_13419);
xnor U13545 (N_13545,N_13303,N_13400);
nor U13546 (N_13546,N_13270,N_13487);
nand U13547 (N_13547,N_13254,N_13396);
or U13548 (N_13548,N_13291,N_13235);
or U13549 (N_13549,N_13318,N_13445);
or U13550 (N_13550,N_13405,N_13350);
nor U13551 (N_13551,N_13316,N_13292);
xor U13552 (N_13552,N_13211,N_13451);
nand U13553 (N_13553,N_13498,N_13365);
nor U13554 (N_13554,N_13311,N_13269);
nor U13555 (N_13555,N_13341,N_13230);
nor U13556 (N_13556,N_13471,N_13393);
xnor U13557 (N_13557,N_13391,N_13252);
xnor U13558 (N_13558,N_13363,N_13424);
nand U13559 (N_13559,N_13496,N_13216);
or U13560 (N_13560,N_13353,N_13461);
xor U13561 (N_13561,N_13334,N_13335);
or U13562 (N_13562,N_13317,N_13343);
nor U13563 (N_13563,N_13261,N_13214);
nand U13564 (N_13564,N_13431,N_13213);
or U13565 (N_13565,N_13479,N_13377);
nand U13566 (N_13566,N_13416,N_13378);
xor U13567 (N_13567,N_13374,N_13217);
nor U13568 (N_13568,N_13421,N_13236);
nand U13569 (N_13569,N_13368,N_13449);
nand U13570 (N_13570,N_13370,N_13260);
nand U13571 (N_13571,N_13475,N_13330);
and U13572 (N_13572,N_13224,N_13408);
or U13573 (N_13573,N_13367,N_13380);
nor U13574 (N_13574,N_13433,N_13429);
or U13575 (N_13575,N_13430,N_13481);
and U13576 (N_13576,N_13307,N_13491);
xnor U13577 (N_13577,N_13282,N_13242);
or U13578 (N_13578,N_13480,N_13422);
and U13579 (N_13579,N_13389,N_13222);
or U13580 (N_13580,N_13319,N_13332);
xnor U13581 (N_13581,N_13394,N_13225);
nor U13582 (N_13582,N_13474,N_13238);
and U13583 (N_13583,N_13231,N_13201);
xor U13584 (N_13584,N_13271,N_13220);
nand U13585 (N_13585,N_13279,N_13312);
nand U13586 (N_13586,N_13395,N_13322);
xor U13587 (N_13587,N_13337,N_13497);
xor U13588 (N_13588,N_13296,N_13402);
or U13589 (N_13589,N_13276,N_13361);
nand U13590 (N_13590,N_13442,N_13473);
or U13591 (N_13591,N_13205,N_13275);
or U13592 (N_13592,N_13490,N_13315);
or U13593 (N_13593,N_13265,N_13457);
or U13594 (N_13594,N_13274,N_13438);
and U13595 (N_13595,N_13346,N_13388);
or U13596 (N_13596,N_13300,N_13234);
nand U13597 (N_13597,N_13229,N_13464);
xnor U13598 (N_13598,N_13371,N_13259);
nor U13599 (N_13599,N_13321,N_13384);
and U13600 (N_13600,N_13440,N_13412);
nand U13601 (N_13601,N_13278,N_13294);
nand U13602 (N_13602,N_13452,N_13458);
nor U13603 (N_13603,N_13258,N_13320);
nand U13604 (N_13604,N_13345,N_13446);
and U13605 (N_13605,N_13399,N_13215);
nand U13606 (N_13606,N_13406,N_13244);
nand U13607 (N_13607,N_13356,N_13314);
nor U13608 (N_13608,N_13241,N_13339);
nand U13609 (N_13609,N_13477,N_13460);
nand U13610 (N_13610,N_13323,N_13326);
nor U13611 (N_13611,N_13410,N_13263);
or U13612 (N_13612,N_13251,N_13221);
xnor U13613 (N_13613,N_13200,N_13392);
xnor U13614 (N_13614,N_13390,N_13250);
and U13615 (N_13615,N_13348,N_13454);
or U13616 (N_13616,N_13359,N_13206);
xnor U13617 (N_13617,N_13255,N_13372);
xnor U13618 (N_13618,N_13333,N_13476);
nor U13619 (N_13619,N_13404,N_13379);
nand U13620 (N_13620,N_13403,N_13472);
and U13621 (N_13621,N_13418,N_13228);
and U13622 (N_13622,N_13357,N_13272);
and U13623 (N_13623,N_13488,N_13223);
nor U13624 (N_13624,N_13456,N_13373);
and U13625 (N_13625,N_13253,N_13366);
nor U13626 (N_13626,N_13207,N_13210);
or U13627 (N_13627,N_13327,N_13486);
and U13628 (N_13628,N_13283,N_13286);
nand U13629 (N_13629,N_13266,N_13347);
nand U13630 (N_13630,N_13435,N_13328);
xor U13631 (N_13631,N_13385,N_13293);
and U13632 (N_13632,N_13417,N_13434);
nand U13633 (N_13633,N_13376,N_13360);
and U13634 (N_13634,N_13463,N_13273);
or U13635 (N_13635,N_13495,N_13232);
nand U13636 (N_13636,N_13310,N_13226);
and U13637 (N_13637,N_13264,N_13437);
or U13638 (N_13638,N_13302,N_13203);
nor U13639 (N_13639,N_13409,N_13284);
or U13640 (N_13640,N_13415,N_13277);
or U13641 (N_13641,N_13465,N_13325);
nand U13642 (N_13642,N_13351,N_13237);
and U13643 (N_13643,N_13468,N_13281);
or U13644 (N_13644,N_13352,N_13340);
xnor U13645 (N_13645,N_13499,N_13423);
or U13646 (N_13646,N_13369,N_13262);
nand U13647 (N_13647,N_13240,N_13268);
xor U13648 (N_13648,N_13267,N_13467);
nor U13649 (N_13649,N_13414,N_13425);
and U13650 (N_13650,N_13410,N_13351);
nor U13651 (N_13651,N_13303,N_13444);
or U13652 (N_13652,N_13374,N_13259);
or U13653 (N_13653,N_13341,N_13278);
or U13654 (N_13654,N_13386,N_13481);
xnor U13655 (N_13655,N_13330,N_13306);
nor U13656 (N_13656,N_13307,N_13415);
and U13657 (N_13657,N_13408,N_13415);
xor U13658 (N_13658,N_13296,N_13476);
and U13659 (N_13659,N_13407,N_13260);
xnor U13660 (N_13660,N_13439,N_13493);
nor U13661 (N_13661,N_13239,N_13264);
nand U13662 (N_13662,N_13404,N_13345);
xnor U13663 (N_13663,N_13315,N_13221);
and U13664 (N_13664,N_13244,N_13348);
nand U13665 (N_13665,N_13484,N_13291);
or U13666 (N_13666,N_13238,N_13351);
nand U13667 (N_13667,N_13207,N_13324);
and U13668 (N_13668,N_13493,N_13367);
or U13669 (N_13669,N_13318,N_13394);
nand U13670 (N_13670,N_13470,N_13460);
xnor U13671 (N_13671,N_13200,N_13460);
or U13672 (N_13672,N_13402,N_13384);
nand U13673 (N_13673,N_13483,N_13262);
nand U13674 (N_13674,N_13308,N_13313);
or U13675 (N_13675,N_13229,N_13285);
and U13676 (N_13676,N_13233,N_13264);
xnor U13677 (N_13677,N_13248,N_13288);
nand U13678 (N_13678,N_13446,N_13370);
xor U13679 (N_13679,N_13438,N_13291);
and U13680 (N_13680,N_13460,N_13252);
nand U13681 (N_13681,N_13268,N_13317);
or U13682 (N_13682,N_13394,N_13344);
nor U13683 (N_13683,N_13207,N_13354);
or U13684 (N_13684,N_13239,N_13215);
nor U13685 (N_13685,N_13365,N_13289);
and U13686 (N_13686,N_13282,N_13433);
nor U13687 (N_13687,N_13474,N_13387);
xor U13688 (N_13688,N_13341,N_13237);
and U13689 (N_13689,N_13386,N_13415);
and U13690 (N_13690,N_13289,N_13253);
xnor U13691 (N_13691,N_13429,N_13347);
or U13692 (N_13692,N_13319,N_13334);
nor U13693 (N_13693,N_13234,N_13408);
and U13694 (N_13694,N_13371,N_13212);
xnor U13695 (N_13695,N_13362,N_13265);
nor U13696 (N_13696,N_13388,N_13443);
or U13697 (N_13697,N_13235,N_13260);
nand U13698 (N_13698,N_13241,N_13382);
nand U13699 (N_13699,N_13421,N_13231);
xor U13700 (N_13700,N_13229,N_13330);
nand U13701 (N_13701,N_13413,N_13297);
nand U13702 (N_13702,N_13450,N_13287);
xnor U13703 (N_13703,N_13428,N_13297);
xnor U13704 (N_13704,N_13440,N_13353);
and U13705 (N_13705,N_13466,N_13403);
nor U13706 (N_13706,N_13442,N_13296);
nor U13707 (N_13707,N_13401,N_13297);
nor U13708 (N_13708,N_13243,N_13453);
nand U13709 (N_13709,N_13260,N_13374);
nor U13710 (N_13710,N_13451,N_13310);
and U13711 (N_13711,N_13423,N_13260);
and U13712 (N_13712,N_13230,N_13388);
nor U13713 (N_13713,N_13331,N_13471);
and U13714 (N_13714,N_13247,N_13228);
nand U13715 (N_13715,N_13236,N_13301);
nand U13716 (N_13716,N_13233,N_13353);
or U13717 (N_13717,N_13451,N_13332);
nand U13718 (N_13718,N_13306,N_13222);
or U13719 (N_13719,N_13447,N_13206);
nor U13720 (N_13720,N_13479,N_13324);
nand U13721 (N_13721,N_13426,N_13441);
xnor U13722 (N_13722,N_13307,N_13445);
nand U13723 (N_13723,N_13273,N_13206);
nor U13724 (N_13724,N_13382,N_13234);
nand U13725 (N_13725,N_13228,N_13421);
nand U13726 (N_13726,N_13209,N_13307);
and U13727 (N_13727,N_13325,N_13439);
xnor U13728 (N_13728,N_13257,N_13499);
nor U13729 (N_13729,N_13252,N_13420);
nand U13730 (N_13730,N_13386,N_13451);
and U13731 (N_13731,N_13331,N_13208);
or U13732 (N_13732,N_13488,N_13240);
xor U13733 (N_13733,N_13252,N_13271);
nor U13734 (N_13734,N_13384,N_13480);
and U13735 (N_13735,N_13412,N_13263);
nand U13736 (N_13736,N_13463,N_13417);
nand U13737 (N_13737,N_13345,N_13438);
nand U13738 (N_13738,N_13203,N_13328);
xnor U13739 (N_13739,N_13384,N_13496);
nor U13740 (N_13740,N_13353,N_13429);
xnor U13741 (N_13741,N_13254,N_13409);
nor U13742 (N_13742,N_13450,N_13256);
and U13743 (N_13743,N_13253,N_13499);
xor U13744 (N_13744,N_13448,N_13416);
and U13745 (N_13745,N_13268,N_13303);
nor U13746 (N_13746,N_13235,N_13484);
xnor U13747 (N_13747,N_13460,N_13361);
nor U13748 (N_13748,N_13410,N_13272);
or U13749 (N_13749,N_13269,N_13449);
nand U13750 (N_13750,N_13366,N_13312);
nor U13751 (N_13751,N_13373,N_13281);
and U13752 (N_13752,N_13464,N_13404);
or U13753 (N_13753,N_13367,N_13471);
and U13754 (N_13754,N_13388,N_13372);
nand U13755 (N_13755,N_13334,N_13204);
nand U13756 (N_13756,N_13334,N_13316);
or U13757 (N_13757,N_13405,N_13460);
nand U13758 (N_13758,N_13460,N_13482);
or U13759 (N_13759,N_13497,N_13482);
and U13760 (N_13760,N_13446,N_13255);
or U13761 (N_13761,N_13337,N_13458);
and U13762 (N_13762,N_13335,N_13216);
and U13763 (N_13763,N_13483,N_13367);
or U13764 (N_13764,N_13356,N_13413);
or U13765 (N_13765,N_13215,N_13434);
or U13766 (N_13766,N_13461,N_13384);
nor U13767 (N_13767,N_13369,N_13269);
nor U13768 (N_13768,N_13486,N_13385);
and U13769 (N_13769,N_13277,N_13340);
or U13770 (N_13770,N_13279,N_13239);
xnor U13771 (N_13771,N_13250,N_13367);
nor U13772 (N_13772,N_13208,N_13328);
or U13773 (N_13773,N_13472,N_13212);
or U13774 (N_13774,N_13388,N_13203);
or U13775 (N_13775,N_13437,N_13276);
nor U13776 (N_13776,N_13446,N_13315);
xnor U13777 (N_13777,N_13232,N_13270);
and U13778 (N_13778,N_13361,N_13351);
nand U13779 (N_13779,N_13267,N_13336);
nor U13780 (N_13780,N_13309,N_13467);
and U13781 (N_13781,N_13239,N_13246);
nand U13782 (N_13782,N_13306,N_13206);
nand U13783 (N_13783,N_13265,N_13421);
xor U13784 (N_13784,N_13437,N_13445);
or U13785 (N_13785,N_13316,N_13208);
xnor U13786 (N_13786,N_13388,N_13367);
nand U13787 (N_13787,N_13244,N_13385);
nand U13788 (N_13788,N_13353,N_13432);
or U13789 (N_13789,N_13321,N_13371);
xor U13790 (N_13790,N_13498,N_13422);
and U13791 (N_13791,N_13297,N_13470);
nor U13792 (N_13792,N_13473,N_13345);
xnor U13793 (N_13793,N_13348,N_13350);
nor U13794 (N_13794,N_13403,N_13296);
and U13795 (N_13795,N_13205,N_13356);
nand U13796 (N_13796,N_13363,N_13275);
nor U13797 (N_13797,N_13475,N_13359);
xnor U13798 (N_13798,N_13213,N_13415);
nor U13799 (N_13799,N_13318,N_13286);
or U13800 (N_13800,N_13779,N_13788);
nor U13801 (N_13801,N_13501,N_13738);
or U13802 (N_13802,N_13623,N_13747);
or U13803 (N_13803,N_13641,N_13682);
nand U13804 (N_13804,N_13662,N_13651);
and U13805 (N_13805,N_13759,N_13567);
nor U13806 (N_13806,N_13755,N_13615);
nand U13807 (N_13807,N_13640,N_13661);
nor U13808 (N_13808,N_13584,N_13707);
and U13809 (N_13809,N_13777,N_13503);
nand U13810 (N_13810,N_13711,N_13511);
nor U13811 (N_13811,N_13671,N_13739);
or U13812 (N_13812,N_13602,N_13774);
or U13813 (N_13813,N_13605,N_13581);
nor U13814 (N_13814,N_13644,N_13643);
and U13815 (N_13815,N_13732,N_13734);
and U13816 (N_13816,N_13655,N_13728);
nor U13817 (N_13817,N_13650,N_13758);
xnor U13818 (N_13818,N_13538,N_13798);
or U13819 (N_13819,N_13741,N_13796);
or U13820 (N_13820,N_13514,N_13786);
and U13821 (N_13821,N_13793,N_13789);
nor U13822 (N_13822,N_13575,N_13632);
xor U13823 (N_13823,N_13543,N_13713);
or U13824 (N_13824,N_13613,N_13519);
xnor U13825 (N_13825,N_13723,N_13636);
and U13826 (N_13826,N_13586,N_13545);
and U13827 (N_13827,N_13700,N_13768);
or U13828 (N_13828,N_13599,N_13626);
and U13829 (N_13829,N_13757,N_13525);
or U13830 (N_13830,N_13516,N_13585);
or U13831 (N_13831,N_13724,N_13672);
or U13832 (N_13832,N_13642,N_13630);
or U13833 (N_13833,N_13782,N_13524);
nor U13834 (N_13834,N_13729,N_13520);
or U13835 (N_13835,N_13578,N_13685);
nor U13836 (N_13836,N_13703,N_13557);
and U13837 (N_13837,N_13744,N_13542);
or U13838 (N_13838,N_13528,N_13761);
or U13839 (N_13839,N_13702,N_13548);
or U13840 (N_13840,N_13694,N_13561);
xnor U13841 (N_13841,N_13592,N_13714);
and U13842 (N_13842,N_13648,N_13750);
and U13843 (N_13843,N_13583,N_13577);
nand U13844 (N_13844,N_13763,N_13721);
xnor U13845 (N_13845,N_13760,N_13752);
xor U13846 (N_13846,N_13611,N_13673);
or U13847 (N_13847,N_13725,N_13621);
xor U13848 (N_13848,N_13692,N_13595);
nor U13849 (N_13849,N_13748,N_13507);
and U13850 (N_13850,N_13628,N_13799);
and U13851 (N_13851,N_13550,N_13709);
nand U13852 (N_13852,N_13677,N_13629);
nor U13853 (N_13853,N_13502,N_13710);
or U13854 (N_13854,N_13535,N_13637);
nand U13855 (N_13855,N_13670,N_13784);
xor U13856 (N_13856,N_13510,N_13513);
or U13857 (N_13857,N_13778,N_13743);
or U13858 (N_13858,N_13506,N_13783);
nand U13859 (N_13859,N_13504,N_13791);
nand U13860 (N_13860,N_13610,N_13517);
and U13861 (N_13861,N_13740,N_13580);
or U13862 (N_13862,N_13532,N_13515);
or U13863 (N_13863,N_13722,N_13730);
xor U13864 (N_13864,N_13781,N_13579);
or U13865 (N_13865,N_13555,N_13657);
and U13866 (N_13866,N_13746,N_13609);
or U13867 (N_13867,N_13681,N_13676);
nor U13868 (N_13868,N_13639,N_13731);
xnor U13869 (N_13869,N_13546,N_13770);
nand U13870 (N_13870,N_13565,N_13688);
and U13871 (N_13871,N_13518,N_13772);
nor U13872 (N_13872,N_13697,N_13544);
xor U13873 (N_13873,N_13572,N_13530);
or U13874 (N_13874,N_13556,N_13618);
and U13875 (N_13875,N_13505,N_13753);
xnor U13876 (N_13876,N_13665,N_13653);
and U13877 (N_13877,N_13634,N_13527);
nand U13878 (N_13878,N_13563,N_13736);
or U13879 (N_13879,N_13566,N_13715);
and U13880 (N_13880,N_13547,N_13619);
or U13881 (N_13881,N_13534,N_13596);
nand U13882 (N_13882,N_13716,N_13797);
or U13883 (N_13883,N_13652,N_13658);
xor U13884 (N_13884,N_13591,N_13687);
and U13885 (N_13885,N_13775,N_13666);
nand U13886 (N_13886,N_13604,N_13559);
xor U13887 (N_13887,N_13536,N_13686);
nor U13888 (N_13888,N_13749,N_13601);
nor U13889 (N_13889,N_13574,N_13690);
nand U13890 (N_13890,N_13588,N_13766);
nand U13891 (N_13891,N_13792,N_13624);
and U13892 (N_13892,N_13568,N_13773);
or U13893 (N_13893,N_13668,N_13638);
and U13894 (N_13894,N_13622,N_13616);
and U13895 (N_13895,N_13706,N_13573);
nor U13896 (N_13896,N_13663,N_13659);
nor U13897 (N_13897,N_13521,N_13582);
nand U13898 (N_13898,N_13705,N_13558);
and U13899 (N_13899,N_13593,N_13674);
nor U13900 (N_13900,N_13589,N_13625);
nand U13901 (N_13901,N_13587,N_13656);
xnor U13902 (N_13902,N_13560,N_13508);
xor U13903 (N_13903,N_13603,N_13509);
nand U13904 (N_13904,N_13751,N_13552);
and U13905 (N_13905,N_13606,N_13689);
and U13906 (N_13906,N_13664,N_13612);
xnor U13907 (N_13907,N_13745,N_13533);
nand U13908 (N_13908,N_13701,N_13785);
or U13909 (N_13909,N_13726,N_13717);
or U13910 (N_13910,N_13795,N_13594);
nand U13911 (N_13911,N_13754,N_13667);
or U13912 (N_13912,N_13645,N_13771);
and U13913 (N_13913,N_13780,N_13680);
and U13914 (N_13914,N_13684,N_13600);
nor U13915 (N_13915,N_13696,N_13675);
nor U13916 (N_13916,N_13551,N_13699);
nand U13917 (N_13917,N_13764,N_13554);
nor U13918 (N_13918,N_13737,N_13712);
xor U13919 (N_13919,N_13564,N_13590);
or U13920 (N_13920,N_13762,N_13756);
nand U13921 (N_13921,N_13649,N_13704);
xnor U13922 (N_13922,N_13539,N_13512);
nand U13923 (N_13923,N_13570,N_13733);
xnor U13924 (N_13924,N_13794,N_13742);
nor U13925 (N_13925,N_13562,N_13608);
xnor U13926 (N_13926,N_13597,N_13526);
or U13927 (N_13927,N_13787,N_13531);
or U13928 (N_13928,N_13537,N_13691);
nand U13929 (N_13929,N_13660,N_13719);
xnor U13930 (N_13930,N_13698,N_13576);
and U13931 (N_13931,N_13647,N_13617);
or U13932 (N_13932,N_13669,N_13646);
nor U13933 (N_13933,N_13614,N_13620);
xnor U13934 (N_13934,N_13776,N_13695);
nand U13935 (N_13935,N_13631,N_13529);
nor U13936 (N_13936,N_13569,N_13607);
nand U13937 (N_13937,N_13654,N_13735);
nor U13938 (N_13938,N_13522,N_13540);
nand U13939 (N_13939,N_13720,N_13727);
nand U13940 (N_13940,N_13553,N_13767);
xor U13941 (N_13941,N_13571,N_13598);
or U13942 (N_13942,N_13708,N_13500);
or U13943 (N_13943,N_13765,N_13679);
nand U13944 (N_13944,N_13769,N_13523);
nor U13945 (N_13945,N_13633,N_13549);
or U13946 (N_13946,N_13678,N_13790);
xnor U13947 (N_13947,N_13718,N_13683);
xnor U13948 (N_13948,N_13541,N_13627);
or U13949 (N_13949,N_13693,N_13635);
or U13950 (N_13950,N_13597,N_13529);
xor U13951 (N_13951,N_13556,N_13729);
or U13952 (N_13952,N_13742,N_13629);
or U13953 (N_13953,N_13541,N_13706);
and U13954 (N_13954,N_13741,N_13681);
nand U13955 (N_13955,N_13789,N_13798);
xor U13956 (N_13956,N_13545,N_13656);
xor U13957 (N_13957,N_13708,N_13785);
or U13958 (N_13958,N_13664,N_13739);
or U13959 (N_13959,N_13743,N_13760);
xor U13960 (N_13960,N_13528,N_13560);
and U13961 (N_13961,N_13576,N_13674);
nor U13962 (N_13962,N_13795,N_13533);
or U13963 (N_13963,N_13788,N_13567);
or U13964 (N_13964,N_13706,N_13759);
or U13965 (N_13965,N_13702,N_13651);
or U13966 (N_13966,N_13605,N_13678);
or U13967 (N_13967,N_13772,N_13696);
xnor U13968 (N_13968,N_13512,N_13550);
xor U13969 (N_13969,N_13588,N_13636);
nor U13970 (N_13970,N_13632,N_13597);
xor U13971 (N_13971,N_13639,N_13553);
nand U13972 (N_13972,N_13508,N_13744);
and U13973 (N_13973,N_13701,N_13613);
xnor U13974 (N_13974,N_13557,N_13753);
nand U13975 (N_13975,N_13544,N_13569);
or U13976 (N_13976,N_13788,N_13601);
or U13977 (N_13977,N_13702,N_13722);
nor U13978 (N_13978,N_13576,N_13608);
nand U13979 (N_13979,N_13765,N_13501);
nand U13980 (N_13980,N_13793,N_13626);
and U13981 (N_13981,N_13719,N_13707);
and U13982 (N_13982,N_13553,N_13763);
nor U13983 (N_13983,N_13628,N_13516);
nor U13984 (N_13984,N_13653,N_13780);
xnor U13985 (N_13985,N_13522,N_13660);
and U13986 (N_13986,N_13785,N_13709);
nand U13987 (N_13987,N_13691,N_13761);
and U13988 (N_13988,N_13796,N_13599);
nor U13989 (N_13989,N_13503,N_13727);
or U13990 (N_13990,N_13516,N_13545);
nor U13991 (N_13991,N_13683,N_13627);
or U13992 (N_13992,N_13679,N_13586);
xor U13993 (N_13993,N_13701,N_13578);
or U13994 (N_13994,N_13550,N_13544);
nand U13995 (N_13995,N_13637,N_13660);
or U13996 (N_13996,N_13512,N_13536);
nor U13997 (N_13997,N_13514,N_13587);
nor U13998 (N_13998,N_13784,N_13766);
and U13999 (N_13999,N_13757,N_13759);
nor U14000 (N_14000,N_13559,N_13712);
nand U14001 (N_14001,N_13705,N_13614);
nor U14002 (N_14002,N_13743,N_13614);
nor U14003 (N_14003,N_13525,N_13793);
and U14004 (N_14004,N_13579,N_13774);
nor U14005 (N_14005,N_13609,N_13699);
nand U14006 (N_14006,N_13623,N_13546);
nor U14007 (N_14007,N_13587,N_13650);
nor U14008 (N_14008,N_13568,N_13625);
or U14009 (N_14009,N_13693,N_13591);
or U14010 (N_14010,N_13736,N_13684);
or U14011 (N_14011,N_13681,N_13538);
and U14012 (N_14012,N_13685,N_13782);
nand U14013 (N_14013,N_13694,N_13534);
or U14014 (N_14014,N_13739,N_13710);
nor U14015 (N_14015,N_13740,N_13743);
nand U14016 (N_14016,N_13505,N_13634);
xor U14017 (N_14017,N_13739,N_13716);
nand U14018 (N_14018,N_13725,N_13795);
xor U14019 (N_14019,N_13754,N_13602);
or U14020 (N_14020,N_13698,N_13670);
nand U14021 (N_14021,N_13699,N_13796);
xnor U14022 (N_14022,N_13604,N_13649);
nand U14023 (N_14023,N_13760,N_13623);
xor U14024 (N_14024,N_13674,N_13550);
or U14025 (N_14025,N_13689,N_13743);
nor U14026 (N_14026,N_13660,N_13544);
nor U14027 (N_14027,N_13657,N_13572);
or U14028 (N_14028,N_13619,N_13694);
xnor U14029 (N_14029,N_13687,N_13711);
or U14030 (N_14030,N_13707,N_13725);
nor U14031 (N_14031,N_13770,N_13566);
nand U14032 (N_14032,N_13714,N_13781);
nand U14033 (N_14033,N_13722,N_13587);
nand U14034 (N_14034,N_13770,N_13653);
nor U14035 (N_14035,N_13508,N_13587);
xnor U14036 (N_14036,N_13502,N_13522);
xnor U14037 (N_14037,N_13771,N_13791);
or U14038 (N_14038,N_13547,N_13577);
or U14039 (N_14039,N_13562,N_13542);
nand U14040 (N_14040,N_13582,N_13634);
nor U14041 (N_14041,N_13583,N_13647);
nand U14042 (N_14042,N_13581,N_13686);
nand U14043 (N_14043,N_13660,N_13770);
nor U14044 (N_14044,N_13642,N_13748);
or U14045 (N_14045,N_13649,N_13573);
nor U14046 (N_14046,N_13600,N_13715);
nand U14047 (N_14047,N_13707,N_13602);
nor U14048 (N_14048,N_13575,N_13603);
nand U14049 (N_14049,N_13720,N_13750);
nor U14050 (N_14050,N_13640,N_13534);
nor U14051 (N_14051,N_13602,N_13741);
xnor U14052 (N_14052,N_13643,N_13554);
nor U14053 (N_14053,N_13506,N_13779);
nor U14054 (N_14054,N_13617,N_13759);
nand U14055 (N_14055,N_13594,N_13515);
nand U14056 (N_14056,N_13742,N_13683);
nor U14057 (N_14057,N_13717,N_13546);
and U14058 (N_14058,N_13754,N_13555);
xnor U14059 (N_14059,N_13549,N_13526);
nor U14060 (N_14060,N_13779,N_13768);
nor U14061 (N_14061,N_13679,N_13712);
and U14062 (N_14062,N_13567,N_13552);
and U14063 (N_14063,N_13760,N_13573);
or U14064 (N_14064,N_13500,N_13518);
nand U14065 (N_14065,N_13638,N_13548);
nor U14066 (N_14066,N_13754,N_13712);
xor U14067 (N_14067,N_13773,N_13655);
nor U14068 (N_14068,N_13571,N_13686);
nand U14069 (N_14069,N_13534,N_13570);
nand U14070 (N_14070,N_13696,N_13630);
and U14071 (N_14071,N_13732,N_13694);
and U14072 (N_14072,N_13792,N_13633);
or U14073 (N_14073,N_13783,N_13609);
or U14074 (N_14074,N_13561,N_13654);
nand U14075 (N_14075,N_13556,N_13732);
or U14076 (N_14076,N_13761,N_13596);
xnor U14077 (N_14077,N_13753,N_13595);
or U14078 (N_14078,N_13555,N_13504);
nand U14079 (N_14079,N_13620,N_13622);
nand U14080 (N_14080,N_13715,N_13797);
nor U14081 (N_14081,N_13584,N_13661);
nand U14082 (N_14082,N_13555,N_13645);
and U14083 (N_14083,N_13588,N_13732);
nor U14084 (N_14084,N_13645,N_13741);
and U14085 (N_14085,N_13766,N_13735);
nand U14086 (N_14086,N_13551,N_13688);
and U14087 (N_14087,N_13601,N_13503);
xor U14088 (N_14088,N_13577,N_13711);
or U14089 (N_14089,N_13794,N_13538);
nand U14090 (N_14090,N_13546,N_13550);
or U14091 (N_14091,N_13759,N_13619);
nand U14092 (N_14092,N_13634,N_13784);
or U14093 (N_14093,N_13534,N_13585);
or U14094 (N_14094,N_13772,N_13718);
xor U14095 (N_14095,N_13613,N_13564);
and U14096 (N_14096,N_13701,N_13790);
nand U14097 (N_14097,N_13776,N_13743);
nor U14098 (N_14098,N_13585,N_13546);
nand U14099 (N_14099,N_13561,N_13621);
and U14100 (N_14100,N_13820,N_13816);
and U14101 (N_14101,N_14010,N_13849);
nor U14102 (N_14102,N_13898,N_14013);
or U14103 (N_14103,N_13917,N_14064);
nor U14104 (N_14104,N_14031,N_13939);
nand U14105 (N_14105,N_13942,N_13891);
xnor U14106 (N_14106,N_13997,N_13828);
nor U14107 (N_14107,N_14048,N_14087);
nor U14108 (N_14108,N_13953,N_13843);
nor U14109 (N_14109,N_13860,N_13932);
nand U14110 (N_14110,N_13804,N_13890);
nor U14111 (N_14111,N_13899,N_13934);
and U14112 (N_14112,N_14046,N_13961);
nand U14113 (N_14113,N_14038,N_13980);
and U14114 (N_14114,N_13928,N_13812);
nand U14115 (N_14115,N_13862,N_13952);
nor U14116 (N_14116,N_14039,N_14084);
nand U14117 (N_14117,N_13954,N_13853);
xor U14118 (N_14118,N_13927,N_13805);
and U14119 (N_14119,N_13814,N_13809);
or U14120 (N_14120,N_14054,N_13993);
nor U14121 (N_14121,N_14015,N_13888);
nor U14122 (N_14122,N_13838,N_13996);
nor U14123 (N_14123,N_13977,N_13861);
nand U14124 (N_14124,N_13992,N_13935);
or U14125 (N_14125,N_13964,N_13887);
nand U14126 (N_14126,N_13894,N_13845);
nand U14127 (N_14127,N_13825,N_14029);
xor U14128 (N_14128,N_14003,N_14008);
nand U14129 (N_14129,N_13854,N_13863);
nor U14130 (N_14130,N_13889,N_14006);
xor U14131 (N_14131,N_14002,N_14096);
or U14132 (N_14132,N_13817,N_13811);
nand U14133 (N_14133,N_13986,N_13978);
nand U14134 (N_14134,N_14056,N_13920);
or U14135 (N_14135,N_13835,N_13913);
xor U14136 (N_14136,N_13925,N_13965);
or U14137 (N_14137,N_14052,N_14095);
nor U14138 (N_14138,N_13915,N_13836);
nor U14139 (N_14139,N_13966,N_14035);
and U14140 (N_14140,N_13867,N_13810);
nor U14141 (N_14141,N_13971,N_13822);
nor U14142 (N_14142,N_13803,N_14070);
and U14143 (N_14143,N_13855,N_13950);
or U14144 (N_14144,N_13901,N_13908);
or U14145 (N_14145,N_13995,N_13989);
or U14146 (N_14146,N_14063,N_13984);
nor U14147 (N_14147,N_13823,N_13856);
and U14148 (N_14148,N_13922,N_14024);
and U14149 (N_14149,N_14082,N_14059);
nor U14150 (N_14150,N_13982,N_13970);
nand U14151 (N_14151,N_14071,N_13834);
and U14152 (N_14152,N_13975,N_14027);
nor U14153 (N_14153,N_13981,N_14021);
or U14154 (N_14154,N_13929,N_13903);
nand U14155 (N_14155,N_14018,N_14014);
nor U14156 (N_14156,N_13829,N_13857);
xor U14157 (N_14157,N_13918,N_13990);
and U14158 (N_14158,N_13991,N_13951);
nor U14159 (N_14159,N_14090,N_14000);
or U14160 (N_14160,N_13998,N_13958);
and U14161 (N_14161,N_13831,N_13886);
nand U14162 (N_14162,N_14091,N_13873);
or U14163 (N_14163,N_14042,N_13983);
or U14164 (N_14164,N_14097,N_13957);
nor U14165 (N_14165,N_14068,N_13976);
and U14166 (N_14166,N_14023,N_13912);
xor U14167 (N_14167,N_13844,N_13858);
or U14168 (N_14168,N_14061,N_13833);
xnor U14169 (N_14169,N_14065,N_14086);
or U14170 (N_14170,N_13907,N_14079);
and U14171 (N_14171,N_14007,N_13956);
nor U14172 (N_14172,N_14045,N_13870);
or U14173 (N_14173,N_13842,N_14005);
nor U14174 (N_14174,N_13974,N_13933);
and U14175 (N_14175,N_14055,N_13988);
and U14176 (N_14176,N_14026,N_13900);
and U14177 (N_14177,N_14032,N_13839);
and U14178 (N_14178,N_13876,N_14088);
nand U14179 (N_14179,N_13896,N_13883);
nand U14180 (N_14180,N_13972,N_13938);
nor U14181 (N_14181,N_14073,N_13827);
nand U14182 (N_14182,N_13830,N_13926);
xnor U14183 (N_14183,N_14020,N_13818);
or U14184 (N_14184,N_13945,N_13910);
and U14185 (N_14185,N_14074,N_14022);
xor U14186 (N_14186,N_13808,N_13902);
or U14187 (N_14187,N_13880,N_13924);
or U14188 (N_14188,N_13999,N_13871);
and U14189 (N_14189,N_14078,N_13962);
or U14190 (N_14190,N_13946,N_13837);
or U14191 (N_14191,N_13906,N_13940);
nor U14192 (N_14192,N_13800,N_13846);
and U14193 (N_14193,N_13968,N_13897);
nor U14194 (N_14194,N_13813,N_14036);
xnor U14195 (N_14195,N_13947,N_13960);
or U14196 (N_14196,N_14051,N_13882);
xnor U14197 (N_14197,N_13850,N_14016);
nor U14198 (N_14198,N_13948,N_13815);
nor U14199 (N_14199,N_13893,N_13919);
and U14200 (N_14200,N_14040,N_14019);
or U14201 (N_14201,N_14098,N_13963);
or U14202 (N_14202,N_14076,N_13985);
nand U14203 (N_14203,N_13916,N_13930);
xnor U14204 (N_14204,N_13921,N_13851);
xnor U14205 (N_14205,N_14092,N_13866);
xnor U14206 (N_14206,N_13819,N_13973);
nand U14207 (N_14207,N_13937,N_13852);
and U14208 (N_14208,N_13905,N_13885);
xnor U14209 (N_14209,N_13959,N_13859);
nor U14210 (N_14210,N_14058,N_13931);
and U14211 (N_14211,N_13909,N_14094);
or U14212 (N_14212,N_13869,N_13895);
xor U14213 (N_14213,N_14033,N_13979);
xor U14214 (N_14214,N_14044,N_13879);
or U14215 (N_14215,N_13911,N_14089);
nor U14216 (N_14216,N_13802,N_13848);
nand U14217 (N_14217,N_13878,N_13832);
and U14218 (N_14218,N_13936,N_13806);
or U14219 (N_14219,N_14017,N_14069);
nor U14220 (N_14220,N_14025,N_13840);
nand U14221 (N_14221,N_14077,N_13987);
nand U14222 (N_14222,N_14072,N_14049);
nor U14223 (N_14223,N_13826,N_14062);
or U14224 (N_14224,N_13821,N_14047);
xor U14225 (N_14225,N_13941,N_14012);
nor U14226 (N_14226,N_14067,N_14075);
and U14227 (N_14227,N_14034,N_14083);
or U14228 (N_14228,N_14009,N_13914);
or U14229 (N_14229,N_13841,N_14099);
nand U14230 (N_14230,N_14028,N_14053);
or U14231 (N_14231,N_14037,N_13801);
nor U14232 (N_14232,N_14011,N_14001);
nor U14233 (N_14233,N_13824,N_13967);
nor U14234 (N_14234,N_13868,N_13969);
or U14235 (N_14235,N_14066,N_13877);
and U14236 (N_14236,N_13847,N_13884);
nor U14237 (N_14237,N_13904,N_13881);
xor U14238 (N_14238,N_13944,N_14041);
xor U14239 (N_14239,N_14057,N_13807);
xnor U14240 (N_14240,N_14085,N_13943);
and U14241 (N_14241,N_13864,N_13994);
or U14242 (N_14242,N_13874,N_13875);
nor U14243 (N_14243,N_14093,N_13955);
or U14244 (N_14244,N_14080,N_13865);
and U14245 (N_14245,N_14004,N_14081);
or U14246 (N_14246,N_14060,N_13892);
nand U14247 (N_14247,N_14043,N_14030);
nor U14248 (N_14248,N_13949,N_13923);
or U14249 (N_14249,N_14050,N_13872);
nand U14250 (N_14250,N_13860,N_13809);
and U14251 (N_14251,N_13823,N_14034);
nand U14252 (N_14252,N_13942,N_13906);
or U14253 (N_14253,N_14048,N_13937);
nor U14254 (N_14254,N_13864,N_13993);
nand U14255 (N_14255,N_14044,N_14068);
or U14256 (N_14256,N_14098,N_13996);
and U14257 (N_14257,N_13968,N_14060);
nand U14258 (N_14258,N_13968,N_13891);
nor U14259 (N_14259,N_14086,N_14058);
or U14260 (N_14260,N_13896,N_14056);
nor U14261 (N_14261,N_13959,N_13926);
nor U14262 (N_14262,N_13924,N_14016);
or U14263 (N_14263,N_14020,N_13932);
and U14264 (N_14264,N_13858,N_14039);
nor U14265 (N_14265,N_14053,N_14036);
or U14266 (N_14266,N_14084,N_14088);
nand U14267 (N_14267,N_13920,N_14011);
and U14268 (N_14268,N_14036,N_14020);
nor U14269 (N_14269,N_13841,N_13938);
xor U14270 (N_14270,N_13848,N_14003);
and U14271 (N_14271,N_13816,N_13931);
and U14272 (N_14272,N_13869,N_14014);
and U14273 (N_14273,N_13922,N_13841);
and U14274 (N_14274,N_13981,N_14077);
or U14275 (N_14275,N_14030,N_14074);
nand U14276 (N_14276,N_13975,N_14096);
xnor U14277 (N_14277,N_13815,N_14057);
xnor U14278 (N_14278,N_14040,N_14095);
nor U14279 (N_14279,N_13919,N_14026);
or U14280 (N_14280,N_13893,N_13877);
xnor U14281 (N_14281,N_13937,N_14018);
nor U14282 (N_14282,N_14082,N_13968);
or U14283 (N_14283,N_13999,N_13966);
and U14284 (N_14284,N_13811,N_14058);
nor U14285 (N_14285,N_13826,N_14013);
and U14286 (N_14286,N_14036,N_13969);
and U14287 (N_14287,N_13991,N_14066);
or U14288 (N_14288,N_14048,N_14046);
nor U14289 (N_14289,N_14027,N_13981);
xnor U14290 (N_14290,N_14047,N_13807);
xnor U14291 (N_14291,N_14019,N_13857);
nand U14292 (N_14292,N_13801,N_13940);
xor U14293 (N_14293,N_14082,N_13916);
and U14294 (N_14294,N_14017,N_14025);
and U14295 (N_14295,N_13910,N_13892);
and U14296 (N_14296,N_14020,N_13819);
nand U14297 (N_14297,N_13875,N_13974);
and U14298 (N_14298,N_14055,N_13806);
nor U14299 (N_14299,N_14015,N_13972);
xnor U14300 (N_14300,N_13958,N_13879);
nor U14301 (N_14301,N_14032,N_13814);
xor U14302 (N_14302,N_13922,N_14056);
xnor U14303 (N_14303,N_13958,N_13888);
nor U14304 (N_14304,N_13937,N_14025);
xnor U14305 (N_14305,N_13967,N_14037);
xor U14306 (N_14306,N_13939,N_14007);
and U14307 (N_14307,N_13890,N_13907);
nand U14308 (N_14308,N_14090,N_13930);
and U14309 (N_14309,N_13882,N_13827);
nor U14310 (N_14310,N_14036,N_13865);
nand U14311 (N_14311,N_13822,N_14083);
or U14312 (N_14312,N_14048,N_14088);
and U14313 (N_14313,N_13823,N_14077);
nor U14314 (N_14314,N_14058,N_14034);
nand U14315 (N_14315,N_13941,N_14001);
or U14316 (N_14316,N_13957,N_14050);
xor U14317 (N_14317,N_14044,N_13997);
and U14318 (N_14318,N_13886,N_13958);
nor U14319 (N_14319,N_14014,N_13823);
and U14320 (N_14320,N_13816,N_13807);
xnor U14321 (N_14321,N_13817,N_14046);
nand U14322 (N_14322,N_13944,N_13854);
nor U14323 (N_14323,N_13949,N_14004);
or U14324 (N_14324,N_13855,N_14071);
xor U14325 (N_14325,N_13876,N_14063);
xnor U14326 (N_14326,N_14028,N_13802);
nand U14327 (N_14327,N_14033,N_14004);
xor U14328 (N_14328,N_13891,N_13973);
and U14329 (N_14329,N_13813,N_14009);
nor U14330 (N_14330,N_14042,N_14095);
and U14331 (N_14331,N_13865,N_14050);
xnor U14332 (N_14332,N_13820,N_13857);
xnor U14333 (N_14333,N_14024,N_13996);
nor U14334 (N_14334,N_14007,N_13951);
nor U14335 (N_14335,N_14049,N_14043);
xnor U14336 (N_14336,N_14096,N_14091);
nand U14337 (N_14337,N_13928,N_13916);
or U14338 (N_14338,N_13817,N_13835);
nor U14339 (N_14339,N_14012,N_13942);
nand U14340 (N_14340,N_13904,N_13801);
nor U14341 (N_14341,N_13962,N_14082);
xnor U14342 (N_14342,N_13881,N_14083);
or U14343 (N_14343,N_14079,N_13844);
and U14344 (N_14344,N_13896,N_14007);
nor U14345 (N_14345,N_14070,N_14088);
and U14346 (N_14346,N_13876,N_14059);
nand U14347 (N_14347,N_14092,N_13897);
xnor U14348 (N_14348,N_13913,N_13926);
or U14349 (N_14349,N_14057,N_14011);
nor U14350 (N_14350,N_13844,N_13889);
xnor U14351 (N_14351,N_14095,N_13863);
nand U14352 (N_14352,N_13888,N_13919);
and U14353 (N_14353,N_13949,N_13838);
xnor U14354 (N_14354,N_13932,N_13911);
or U14355 (N_14355,N_14001,N_14098);
nand U14356 (N_14356,N_13933,N_13966);
or U14357 (N_14357,N_14094,N_13818);
nand U14358 (N_14358,N_13936,N_14001);
nor U14359 (N_14359,N_14051,N_13847);
and U14360 (N_14360,N_13930,N_14071);
xor U14361 (N_14361,N_13954,N_14001);
nand U14362 (N_14362,N_13924,N_13872);
xor U14363 (N_14363,N_14050,N_14057);
or U14364 (N_14364,N_13989,N_14095);
xnor U14365 (N_14365,N_14084,N_13904);
or U14366 (N_14366,N_14020,N_14049);
and U14367 (N_14367,N_14078,N_14022);
or U14368 (N_14368,N_13895,N_13862);
or U14369 (N_14369,N_13854,N_14047);
nand U14370 (N_14370,N_14084,N_14076);
nor U14371 (N_14371,N_13866,N_13854);
nor U14372 (N_14372,N_13807,N_14006);
or U14373 (N_14373,N_13867,N_14039);
xor U14374 (N_14374,N_13852,N_13995);
nor U14375 (N_14375,N_14024,N_13845);
or U14376 (N_14376,N_14077,N_14030);
nor U14377 (N_14377,N_14062,N_13843);
nand U14378 (N_14378,N_13906,N_13852);
nor U14379 (N_14379,N_13830,N_14060);
or U14380 (N_14380,N_14084,N_13934);
and U14381 (N_14381,N_13842,N_13861);
xor U14382 (N_14382,N_13880,N_14023);
nand U14383 (N_14383,N_14082,N_13935);
xor U14384 (N_14384,N_14051,N_14064);
and U14385 (N_14385,N_14092,N_13937);
nor U14386 (N_14386,N_13803,N_13933);
nand U14387 (N_14387,N_14053,N_13895);
or U14388 (N_14388,N_13834,N_13924);
nand U14389 (N_14389,N_13909,N_14099);
nor U14390 (N_14390,N_14088,N_13959);
xor U14391 (N_14391,N_13825,N_14077);
or U14392 (N_14392,N_13890,N_13803);
and U14393 (N_14393,N_13887,N_13806);
nand U14394 (N_14394,N_14061,N_13917);
nand U14395 (N_14395,N_14001,N_13995);
or U14396 (N_14396,N_14090,N_13929);
or U14397 (N_14397,N_13966,N_14020);
xnor U14398 (N_14398,N_13929,N_13970);
and U14399 (N_14399,N_13994,N_14060);
xor U14400 (N_14400,N_14115,N_14375);
and U14401 (N_14401,N_14111,N_14117);
nor U14402 (N_14402,N_14388,N_14316);
and U14403 (N_14403,N_14183,N_14379);
nor U14404 (N_14404,N_14135,N_14312);
nand U14405 (N_14405,N_14287,N_14241);
or U14406 (N_14406,N_14180,N_14181);
and U14407 (N_14407,N_14167,N_14325);
xnor U14408 (N_14408,N_14277,N_14200);
nor U14409 (N_14409,N_14357,N_14188);
nand U14410 (N_14410,N_14210,N_14237);
and U14411 (N_14411,N_14259,N_14367);
and U14412 (N_14412,N_14278,N_14128);
nand U14413 (N_14413,N_14219,N_14354);
and U14414 (N_14414,N_14308,N_14398);
nand U14415 (N_14415,N_14220,N_14368);
nand U14416 (N_14416,N_14189,N_14217);
xnor U14417 (N_14417,N_14332,N_14168);
nor U14418 (N_14418,N_14131,N_14154);
nand U14419 (N_14419,N_14336,N_14374);
and U14420 (N_14420,N_14299,N_14184);
nor U14421 (N_14421,N_14132,N_14397);
nand U14422 (N_14422,N_14173,N_14164);
and U14423 (N_14423,N_14344,N_14106);
nand U14424 (N_14424,N_14257,N_14209);
nand U14425 (N_14425,N_14350,N_14395);
or U14426 (N_14426,N_14255,N_14364);
nor U14427 (N_14427,N_14177,N_14347);
xor U14428 (N_14428,N_14162,N_14110);
or U14429 (N_14429,N_14270,N_14273);
and U14430 (N_14430,N_14334,N_14383);
and U14431 (N_14431,N_14384,N_14203);
xor U14432 (N_14432,N_14120,N_14208);
xnor U14433 (N_14433,N_14390,N_14335);
and U14434 (N_14434,N_14235,N_14339);
and U14435 (N_14435,N_14207,N_14391);
and U14436 (N_14436,N_14349,N_14254);
nor U14437 (N_14437,N_14320,N_14360);
nand U14438 (N_14438,N_14366,N_14199);
nor U14439 (N_14439,N_14263,N_14190);
nor U14440 (N_14440,N_14202,N_14348);
nor U14441 (N_14441,N_14317,N_14142);
or U14442 (N_14442,N_14187,N_14365);
nand U14443 (N_14443,N_14280,N_14311);
xnor U14444 (N_14444,N_14371,N_14324);
xor U14445 (N_14445,N_14319,N_14153);
nor U14446 (N_14446,N_14197,N_14330);
nand U14447 (N_14447,N_14288,N_14307);
nand U14448 (N_14448,N_14387,N_14205);
or U14449 (N_14449,N_14138,N_14107);
and U14450 (N_14450,N_14266,N_14256);
or U14451 (N_14451,N_14230,N_14300);
and U14452 (N_14452,N_14340,N_14147);
nand U14453 (N_14453,N_14245,N_14179);
and U14454 (N_14454,N_14216,N_14338);
nor U14455 (N_14455,N_14136,N_14114);
nor U14456 (N_14456,N_14198,N_14314);
or U14457 (N_14457,N_14103,N_14359);
and U14458 (N_14458,N_14313,N_14298);
nor U14459 (N_14459,N_14370,N_14112);
nand U14460 (N_14460,N_14382,N_14396);
nor U14461 (N_14461,N_14294,N_14226);
xor U14462 (N_14462,N_14272,N_14109);
nand U14463 (N_14463,N_14170,N_14105);
or U14464 (N_14464,N_14283,N_14305);
and U14465 (N_14465,N_14356,N_14269);
nor U14466 (N_14466,N_14119,N_14211);
or U14467 (N_14467,N_14137,N_14133);
xor U14468 (N_14468,N_14333,N_14250);
nand U14469 (N_14469,N_14353,N_14303);
or U14470 (N_14470,N_14104,N_14102);
and U14471 (N_14471,N_14149,N_14140);
and U14472 (N_14472,N_14224,N_14373);
and U14473 (N_14473,N_14297,N_14281);
or U14474 (N_14474,N_14125,N_14213);
or U14475 (N_14475,N_14141,N_14157);
xor U14476 (N_14476,N_14186,N_14369);
xor U14477 (N_14477,N_14352,N_14243);
nand U14478 (N_14478,N_14225,N_14399);
or U14479 (N_14479,N_14214,N_14378);
and U14480 (N_14480,N_14232,N_14171);
nor U14481 (N_14481,N_14322,N_14218);
or U14482 (N_14482,N_14304,N_14328);
nor U14483 (N_14483,N_14282,N_14337);
nor U14484 (N_14484,N_14155,N_14108);
or U14485 (N_14485,N_14363,N_14268);
or U14486 (N_14486,N_14151,N_14260);
nand U14487 (N_14487,N_14329,N_14160);
nor U14488 (N_14488,N_14302,N_14234);
and U14489 (N_14489,N_14163,N_14318);
and U14490 (N_14490,N_14295,N_14124);
xnor U14491 (N_14491,N_14385,N_14389);
and U14492 (N_14492,N_14323,N_14315);
xnor U14493 (N_14493,N_14331,N_14301);
nand U14494 (N_14494,N_14293,N_14158);
nor U14495 (N_14495,N_14252,N_14355);
or U14496 (N_14496,N_14166,N_14229);
or U14497 (N_14497,N_14127,N_14345);
nand U14498 (N_14498,N_14172,N_14321);
or U14499 (N_14499,N_14122,N_14285);
nor U14500 (N_14500,N_14247,N_14238);
and U14501 (N_14501,N_14291,N_14244);
nor U14502 (N_14502,N_14326,N_14361);
and U14503 (N_14503,N_14194,N_14386);
nand U14504 (N_14504,N_14195,N_14204);
nor U14505 (N_14505,N_14146,N_14292);
nor U14506 (N_14506,N_14242,N_14246);
nand U14507 (N_14507,N_14286,N_14144);
and U14508 (N_14508,N_14206,N_14215);
xor U14509 (N_14509,N_14342,N_14264);
xnor U14510 (N_14510,N_14143,N_14185);
or U14511 (N_14511,N_14201,N_14327);
and U14512 (N_14512,N_14258,N_14351);
or U14513 (N_14513,N_14276,N_14150);
nand U14514 (N_14514,N_14239,N_14271);
nand U14515 (N_14515,N_14251,N_14152);
or U14516 (N_14516,N_14182,N_14159);
nor U14517 (N_14517,N_14358,N_14196);
or U14518 (N_14518,N_14310,N_14228);
nor U14519 (N_14519,N_14118,N_14267);
or U14520 (N_14520,N_14296,N_14362);
nand U14521 (N_14521,N_14381,N_14126);
nor U14522 (N_14522,N_14231,N_14233);
and U14523 (N_14523,N_14148,N_14341);
nor U14524 (N_14524,N_14262,N_14248);
xnor U14525 (N_14525,N_14393,N_14178);
or U14526 (N_14526,N_14156,N_14123);
and U14527 (N_14527,N_14274,N_14289);
nor U14528 (N_14528,N_14376,N_14227);
xor U14529 (N_14529,N_14343,N_14134);
or U14530 (N_14530,N_14261,N_14306);
nor U14531 (N_14531,N_14139,N_14221);
or U14532 (N_14532,N_14240,N_14394);
or U14533 (N_14533,N_14129,N_14372);
and U14534 (N_14534,N_14191,N_14121);
and U14535 (N_14535,N_14346,N_14174);
and U14536 (N_14536,N_14113,N_14290);
nand U14537 (N_14537,N_14175,N_14275);
and U14538 (N_14538,N_14309,N_14145);
nand U14539 (N_14539,N_14284,N_14253);
nand U14540 (N_14540,N_14192,N_14377);
xnor U14541 (N_14541,N_14161,N_14223);
and U14542 (N_14542,N_14169,N_14101);
xnor U14543 (N_14543,N_14100,N_14176);
or U14544 (N_14544,N_14279,N_14392);
and U14545 (N_14545,N_14130,N_14212);
xor U14546 (N_14546,N_14236,N_14222);
nand U14547 (N_14547,N_14249,N_14165);
or U14548 (N_14548,N_14380,N_14116);
and U14549 (N_14549,N_14265,N_14193);
xor U14550 (N_14550,N_14376,N_14153);
xor U14551 (N_14551,N_14264,N_14297);
or U14552 (N_14552,N_14266,N_14311);
or U14553 (N_14553,N_14126,N_14386);
or U14554 (N_14554,N_14274,N_14110);
and U14555 (N_14555,N_14266,N_14204);
or U14556 (N_14556,N_14251,N_14396);
nand U14557 (N_14557,N_14238,N_14210);
and U14558 (N_14558,N_14161,N_14137);
or U14559 (N_14559,N_14240,N_14300);
nand U14560 (N_14560,N_14314,N_14397);
nor U14561 (N_14561,N_14253,N_14181);
xor U14562 (N_14562,N_14184,N_14223);
nand U14563 (N_14563,N_14214,N_14302);
and U14564 (N_14564,N_14174,N_14134);
nand U14565 (N_14565,N_14367,N_14138);
nand U14566 (N_14566,N_14297,N_14222);
or U14567 (N_14567,N_14101,N_14270);
xor U14568 (N_14568,N_14314,N_14359);
nor U14569 (N_14569,N_14159,N_14327);
xor U14570 (N_14570,N_14323,N_14292);
and U14571 (N_14571,N_14352,N_14151);
nor U14572 (N_14572,N_14315,N_14103);
and U14573 (N_14573,N_14246,N_14311);
xor U14574 (N_14574,N_14222,N_14294);
xor U14575 (N_14575,N_14319,N_14352);
nor U14576 (N_14576,N_14189,N_14175);
and U14577 (N_14577,N_14243,N_14355);
xor U14578 (N_14578,N_14139,N_14321);
xnor U14579 (N_14579,N_14118,N_14382);
or U14580 (N_14580,N_14296,N_14120);
or U14581 (N_14581,N_14236,N_14101);
and U14582 (N_14582,N_14223,N_14149);
nor U14583 (N_14583,N_14162,N_14181);
or U14584 (N_14584,N_14348,N_14203);
and U14585 (N_14585,N_14250,N_14290);
or U14586 (N_14586,N_14230,N_14363);
and U14587 (N_14587,N_14380,N_14399);
xor U14588 (N_14588,N_14324,N_14241);
xor U14589 (N_14589,N_14233,N_14382);
xnor U14590 (N_14590,N_14146,N_14343);
nand U14591 (N_14591,N_14282,N_14366);
nor U14592 (N_14592,N_14334,N_14173);
and U14593 (N_14593,N_14397,N_14109);
nor U14594 (N_14594,N_14326,N_14176);
xor U14595 (N_14595,N_14125,N_14394);
nor U14596 (N_14596,N_14111,N_14235);
nor U14597 (N_14597,N_14301,N_14319);
nand U14598 (N_14598,N_14237,N_14251);
or U14599 (N_14599,N_14103,N_14298);
or U14600 (N_14600,N_14135,N_14261);
xor U14601 (N_14601,N_14361,N_14307);
xor U14602 (N_14602,N_14319,N_14267);
xor U14603 (N_14603,N_14271,N_14117);
nand U14604 (N_14604,N_14304,N_14123);
xnor U14605 (N_14605,N_14141,N_14245);
nand U14606 (N_14606,N_14196,N_14387);
xor U14607 (N_14607,N_14282,N_14255);
or U14608 (N_14608,N_14194,N_14370);
xor U14609 (N_14609,N_14392,N_14266);
xnor U14610 (N_14610,N_14234,N_14236);
xor U14611 (N_14611,N_14116,N_14206);
nand U14612 (N_14612,N_14224,N_14216);
and U14613 (N_14613,N_14339,N_14337);
and U14614 (N_14614,N_14254,N_14332);
nand U14615 (N_14615,N_14202,N_14244);
or U14616 (N_14616,N_14302,N_14245);
xor U14617 (N_14617,N_14276,N_14372);
nand U14618 (N_14618,N_14149,N_14370);
and U14619 (N_14619,N_14259,N_14358);
nand U14620 (N_14620,N_14285,N_14365);
or U14621 (N_14621,N_14340,N_14203);
xor U14622 (N_14622,N_14263,N_14296);
nor U14623 (N_14623,N_14135,N_14117);
or U14624 (N_14624,N_14190,N_14132);
or U14625 (N_14625,N_14159,N_14112);
nor U14626 (N_14626,N_14340,N_14155);
xnor U14627 (N_14627,N_14195,N_14310);
nor U14628 (N_14628,N_14255,N_14355);
nand U14629 (N_14629,N_14136,N_14177);
and U14630 (N_14630,N_14300,N_14243);
nand U14631 (N_14631,N_14240,N_14162);
and U14632 (N_14632,N_14113,N_14285);
nand U14633 (N_14633,N_14160,N_14127);
xor U14634 (N_14634,N_14270,N_14239);
nand U14635 (N_14635,N_14226,N_14237);
xnor U14636 (N_14636,N_14154,N_14212);
nand U14637 (N_14637,N_14287,N_14264);
xnor U14638 (N_14638,N_14179,N_14144);
nand U14639 (N_14639,N_14182,N_14352);
and U14640 (N_14640,N_14387,N_14204);
xnor U14641 (N_14641,N_14382,N_14262);
nor U14642 (N_14642,N_14345,N_14376);
and U14643 (N_14643,N_14372,N_14312);
xor U14644 (N_14644,N_14349,N_14145);
or U14645 (N_14645,N_14234,N_14294);
xnor U14646 (N_14646,N_14129,N_14133);
nor U14647 (N_14647,N_14179,N_14118);
xnor U14648 (N_14648,N_14335,N_14144);
and U14649 (N_14649,N_14354,N_14144);
xor U14650 (N_14650,N_14229,N_14245);
xor U14651 (N_14651,N_14139,N_14122);
and U14652 (N_14652,N_14104,N_14320);
nor U14653 (N_14653,N_14238,N_14361);
nor U14654 (N_14654,N_14234,N_14239);
or U14655 (N_14655,N_14191,N_14268);
nor U14656 (N_14656,N_14159,N_14149);
nand U14657 (N_14657,N_14134,N_14200);
or U14658 (N_14658,N_14315,N_14195);
and U14659 (N_14659,N_14147,N_14163);
and U14660 (N_14660,N_14288,N_14231);
nor U14661 (N_14661,N_14175,N_14330);
nand U14662 (N_14662,N_14101,N_14348);
or U14663 (N_14663,N_14305,N_14165);
nor U14664 (N_14664,N_14159,N_14242);
or U14665 (N_14665,N_14229,N_14140);
nand U14666 (N_14666,N_14298,N_14168);
xor U14667 (N_14667,N_14109,N_14249);
nor U14668 (N_14668,N_14186,N_14206);
or U14669 (N_14669,N_14264,N_14265);
and U14670 (N_14670,N_14354,N_14250);
nand U14671 (N_14671,N_14310,N_14205);
xor U14672 (N_14672,N_14268,N_14299);
and U14673 (N_14673,N_14378,N_14340);
and U14674 (N_14674,N_14234,N_14251);
nand U14675 (N_14675,N_14266,N_14276);
nor U14676 (N_14676,N_14211,N_14103);
and U14677 (N_14677,N_14141,N_14151);
nand U14678 (N_14678,N_14208,N_14258);
or U14679 (N_14679,N_14120,N_14246);
nor U14680 (N_14680,N_14153,N_14130);
nand U14681 (N_14681,N_14312,N_14189);
and U14682 (N_14682,N_14271,N_14345);
nor U14683 (N_14683,N_14309,N_14391);
nor U14684 (N_14684,N_14255,N_14396);
nand U14685 (N_14685,N_14381,N_14383);
or U14686 (N_14686,N_14133,N_14158);
nand U14687 (N_14687,N_14142,N_14323);
and U14688 (N_14688,N_14335,N_14267);
nor U14689 (N_14689,N_14330,N_14178);
nor U14690 (N_14690,N_14172,N_14109);
or U14691 (N_14691,N_14351,N_14398);
or U14692 (N_14692,N_14139,N_14154);
or U14693 (N_14693,N_14168,N_14190);
xor U14694 (N_14694,N_14282,N_14298);
and U14695 (N_14695,N_14324,N_14302);
or U14696 (N_14696,N_14123,N_14391);
xor U14697 (N_14697,N_14329,N_14367);
nor U14698 (N_14698,N_14237,N_14214);
or U14699 (N_14699,N_14193,N_14355);
xor U14700 (N_14700,N_14444,N_14489);
or U14701 (N_14701,N_14664,N_14486);
xor U14702 (N_14702,N_14502,N_14592);
or U14703 (N_14703,N_14557,N_14605);
and U14704 (N_14704,N_14689,N_14448);
or U14705 (N_14705,N_14660,N_14650);
nand U14706 (N_14706,N_14493,N_14602);
xnor U14707 (N_14707,N_14668,N_14694);
nor U14708 (N_14708,N_14413,N_14427);
nor U14709 (N_14709,N_14492,N_14421);
nor U14710 (N_14710,N_14613,N_14560);
and U14711 (N_14711,N_14675,N_14482);
and U14712 (N_14712,N_14666,N_14443);
nor U14713 (N_14713,N_14643,N_14572);
nor U14714 (N_14714,N_14642,N_14523);
and U14715 (N_14715,N_14564,N_14635);
or U14716 (N_14716,N_14428,N_14434);
and U14717 (N_14717,N_14681,N_14546);
and U14718 (N_14718,N_14671,N_14562);
nor U14719 (N_14719,N_14518,N_14497);
or U14720 (N_14720,N_14547,N_14691);
or U14721 (N_14721,N_14683,N_14424);
and U14722 (N_14722,N_14555,N_14699);
xnor U14723 (N_14723,N_14506,N_14563);
nand U14724 (N_14724,N_14690,N_14442);
and U14725 (N_14725,N_14591,N_14447);
xnor U14726 (N_14726,N_14619,N_14475);
xnor U14727 (N_14727,N_14498,N_14400);
nand U14728 (N_14728,N_14617,N_14631);
xor U14729 (N_14729,N_14558,N_14543);
and U14730 (N_14730,N_14623,N_14533);
nor U14731 (N_14731,N_14569,N_14685);
and U14732 (N_14732,N_14640,N_14473);
xnor U14733 (N_14733,N_14577,N_14437);
nor U14734 (N_14734,N_14637,N_14471);
nand U14735 (N_14735,N_14653,N_14522);
nor U14736 (N_14736,N_14624,N_14468);
xnor U14737 (N_14737,N_14404,N_14432);
xor U14738 (N_14738,N_14559,N_14667);
nor U14739 (N_14739,N_14586,N_14512);
or U14740 (N_14740,N_14549,N_14414);
nand U14741 (N_14741,N_14672,N_14536);
nand U14742 (N_14742,N_14670,N_14464);
nor U14743 (N_14743,N_14466,N_14460);
nand U14744 (N_14744,N_14607,N_14500);
nor U14745 (N_14745,N_14589,N_14554);
nor U14746 (N_14746,N_14641,N_14620);
xnor U14747 (N_14747,N_14688,N_14696);
nand U14748 (N_14748,N_14556,N_14467);
nand U14749 (N_14749,N_14611,N_14665);
and U14750 (N_14750,N_14509,N_14545);
nand U14751 (N_14751,N_14638,N_14423);
nand U14752 (N_14752,N_14603,N_14618);
nand U14753 (N_14753,N_14480,N_14584);
xnor U14754 (N_14754,N_14416,N_14580);
xor U14755 (N_14755,N_14573,N_14504);
xor U14756 (N_14756,N_14519,N_14651);
nor U14757 (N_14757,N_14422,N_14438);
xor U14758 (N_14758,N_14657,N_14654);
nand U14759 (N_14759,N_14632,N_14487);
xor U14760 (N_14760,N_14596,N_14590);
xnor U14761 (N_14761,N_14417,N_14658);
nand U14762 (N_14762,N_14679,N_14594);
or U14763 (N_14763,N_14561,N_14410);
nand U14764 (N_14764,N_14494,N_14646);
nor U14765 (N_14765,N_14453,N_14692);
xor U14766 (N_14766,N_14520,N_14540);
and U14767 (N_14767,N_14441,N_14528);
nand U14768 (N_14768,N_14610,N_14526);
nor U14769 (N_14769,N_14604,N_14525);
xnor U14770 (N_14770,N_14571,N_14601);
and U14771 (N_14771,N_14662,N_14581);
xnor U14772 (N_14772,N_14595,N_14541);
or U14773 (N_14773,N_14682,N_14656);
and U14774 (N_14774,N_14508,N_14582);
and U14775 (N_14775,N_14621,N_14588);
nand U14776 (N_14776,N_14503,N_14644);
and U14777 (N_14777,N_14609,N_14659);
xnor U14778 (N_14778,N_14511,N_14578);
nand U14779 (N_14779,N_14538,N_14457);
and U14780 (N_14780,N_14515,N_14614);
nor U14781 (N_14781,N_14472,N_14677);
nor U14782 (N_14782,N_14425,N_14686);
nor U14783 (N_14783,N_14478,N_14627);
nor U14784 (N_14784,N_14474,N_14531);
nand U14785 (N_14785,N_14458,N_14440);
nor U14786 (N_14786,N_14647,N_14450);
and U14787 (N_14787,N_14491,N_14553);
and U14788 (N_14788,N_14575,N_14676);
nor U14789 (N_14789,N_14687,N_14496);
nor U14790 (N_14790,N_14680,N_14465);
xor U14791 (N_14791,N_14663,N_14648);
and U14792 (N_14792,N_14429,N_14435);
nand U14793 (N_14793,N_14456,N_14524);
nand U14794 (N_14794,N_14628,N_14461);
or U14795 (N_14795,N_14587,N_14645);
nor U14796 (N_14796,N_14477,N_14405);
nand U14797 (N_14797,N_14420,N_14583);
nor U14798 (N_14798,N_14418,N_14551);
nand U14799 (N_14799,N_14516,N_14629);
xor U14800 (N_14800,N_14537,N_14579);
or U14801 (N_14801,N_14483,N_14597);
xor U14802 (N_14802,N_14661,N_14552);
nand U14803 (N_14803,N_14535,N_14485);
or U14804 (N_14804,N_14406,N_14499);
nand U14805 (N_14805,N_14513,N_14693);
nand U14806 (N_14806,N_14539,N_14673);
nand U14807 (N_14807,N_14636,N_14445);
xnor U14808 (N_14808,N_14455,N_14530);
xnor U14809 (N_14809,N_14534,N_14439);
nor U14810 (N_14810,N_14470,N_14568);
xor U14811 (N_14811,N_14501,N_14403);
nand U14812 (N_14812,N_14585,N_14436);
or U14813 (N_14813,N_14408,N_14476);
or U14814 (N_14814,N_14625,N_14615);
nor U14815 (N_14815,N_14419,N_14655);
and U14816 (N_14816,N_14599,N_14532);
nor U14817 (N_14817,N_14402,N_14409);
nor U14818 (N_14818,N_14411,N_14459);
and U14819 (N_14819,N_14479,N_14544);
nand U14820 (N_14820,N_14612,N_14505);
xor U14821 (N_14821,N_14566,N_14593);
or U14822 (N_14822,N_14608,N_14426);
nand U14823 (N_14823,N_14517,N_14622);
and U14824 (N_14824,N_14674,N_14514);
nand U14825 (N_14825,N_14697,N_14449);
or U14826 (N_14826,N_14652,N_14678);
nor U14827 (N_14827,N_14431,N_14401);
nor U14828 (N_14828,N_14550,N_14598);
xnor U14829 (N_14829,N_14574,N_14649);
or U14830 (N_14830,N_14412,N_14463);
or U14831 (N_14831,N_14576,N_14510);
xor U14832 (N_14832,N_14415,N_14606);
nand U14833 (N_14833,N_14600,N_14446);
or U14834 (N_14834,N_14451,N_14542);
nand U14835 (N_14835,N_14567,N_14490);
or U14836 (N_14836,N_14433,N_14495);
or U14837 (N_14837,N_14639,N_14669);
xor U14838 (N_14838,N_14507,N_14452);
xnor U14839 (N_14839,N_14527,N_14529);
and U14840 (N_14840,N_14462,N_14488);
nand U14841 (N_14841,N_14684,N_14633);
and U14842 (N_14842,N_14521,N_14626);
or U14843 (N_14843,N_14548,N_14634);
nand U14844 (N_14844,N_14430,N_14616);
nand U14845 (N_14845,N_14481,N_14695);
or U14846 (N_14846,N_14698,N_14469);
and U14847 (N_14847,N_14565,N_14454);
and U14848 (N_14848,N_14484,N_14570);
or U14849 (N_14849,N_14630,N_14407);
nor U14850 (N_14850,N_14448,N_14555);
nand U14851 (N_14851,N_14691,N_14407);
nand U14852 (N_14852,N_14628,N_14611);
and U14853 (N_14853,N_14550,N_14539);
or U14854 (N_14854,N_14629,N_14496);
xor U14855 (N_14855,N_14558,N_14472);
xor U14856 (N_14856,N_14585,N_14456);
xor U14857 (N_14857,N_14657,N_14505);
xor U14858 (N_14858,N_14429,N_14598);
nor U14859 (N_14859,N_14434,N_14568);
xor U14860 (N_14860,N_14401,N_14466);
xnor U14861 (N_14861,N_14586,N_14539);
xor U14862 (N_14862,N_14627,N_14625);
or U14863 (N_14863,N_14682,N_14543);
or U14864 (N_14864,N_14573,N_14621);
nand U14865 (N_14865,N_14671,N_14631);
nand U14866 (N_14866,N_14629,N_14426);
and U14867 (N_14867,N_14478,N_14401);
xor U14868 (N_14868,N_14507,N_14506);
nand U14869 (N_14869,N_14553,N_14600);
xor U14870 (N_14870,N_14511,N_14680);
nand U14871 (N_14871,N_14582,N_14647);
nand U14872 (N_14872,N_14508,N_14670);
and U14873 (N_14873,N_14665,N_14539);
xor U14874 (N_14874,N_14416,N_14549);
and U14875 (N_14875,N_14429,N_14663);
nor U14876 (N_14876,N_14695,N_14648);
and U14877 (N_14877,N_14650,N_14692);
xor U14878 (N_14878,N_14627,N_14401);
xor U14879 (N_14879,N_14653,N_14683);
or U14880 (N_14880,N_14415,N_14434);
and U14881 (N_14881,N_14438,N_14447);
or U14882 (N_14882,N_14559,N_14585);
or U14883 (N_14883,N_14535,N_14631);
xor U14884 (N_14884,N_14479,N_14594);
and U14885 (N_14885,N_14563,N_14513);
xor U14886 (N_14886,N_14696,N_14692);
or U14887 (N_14887,N_14626,N_14589);
xnor U14888 (N_14888,N_14452,N_14499);
or U14889 (N_14889,N_14612,N_14596);
xor U14890 (N_14890,N_14622,N_14592);
or U14891 (N_14891,N_14520,N_14435);
nor U14892 (N_14892,N_14569,N_14430);
nor U14893 (N_14893,N_14681,N_14624);
nor U14894 (N_14894,N_14446,N_14534);
nand U14895 (N_14895,N_14538,N_14647);
and U14896 (N_14896,N_14462,N_14519);
nand U14897 (N_14897,N_14409,N_14472);
nand U14898 (N_14898,N_14648,N_14543);
xnor U14899 (N_14899,N_14632,N_14463);
nor U14900 (N_14900,N_14497,N_14685);
nor U14901 (N_14901,N_14477,N_14606);
and U14902 (N_14902,N_14515,N_14475);
nand U14903 (N_14903,N_14471,N_14677);
nand U14904 (N_14904,N_14576,N_14456);
nand U14905 (N_14905,N_14697,N_14596);
nand U14906 (N_14906,N_14490,N_14681);
or U14907 (N_14907,N_14527,N_14530);
nand U14908 (N_14908,N_14666,N_14486);
and U14909 (N_14909,N_14542,N_14642);
and U14910 (N_14910,N_14513,N_14660);
or U14911 (N_14911,N_14547,N_14455);
xor U14912 (N_14912,N_14469,N_14598);
nor U14913 (N_14913,N_14553,N_14441);
and U14914 (N_14914,N_14464,N_14413);
and U14915 (N_14915,N_14549,N_14472);
nor U14916 (N_14916,N_14498,N_14524);
xor U14917 (N_14917,N_14558,N_14541);
nand U14918 (N_14918,N_14577,N_14474);
and U14919 (N_14919,N_14445,N_14530);
nand U14920 (N_14920,N_14441,N_14589);
and U14921 (N_14921,N_14407,N_14597);
and U14922 (N_14922,N_14544,N_14416);
or U14923 (N_14923,N_14598,N_14486);
or U14924 (N_14924,N_14624,N_14577);
nand U14925 (N_14925,N_14593,N_14452);
nor U14926 (N_14926,N_14593,N_14416);
nor U14927 (N_14927,N_14607,N_14605);
and U14928 (N_14928,N_14408,N_14518);
nor U14929 (N_14929,N_14565,N_14409);
nor U14930 (N_14930,N_14586,N_14419);
xor U14931 (N_14931,N_14647,N_14626);
xor U14932 (N_14932,N_14600,N_14434);
nand U14933 (N_14933,N_14421,N_14677);
nand U14934 (N_14934,N_14562,N_14558);
xnor U14935 (N_14935,N_14583,N_14606);
or U14936 (N_14936,N_14463,N_14529);
nand U14937 (N_14937,N_14689,N_14609);
nand U14938 (N_14938,N_14583,N_14404);
nand U14939 (N_14939,N_14683,N_14608);
xnor U14940 (N_14940,N_14699,N_14553);
xnor U14941 (N_14941,N_14566,N_14564);
xor U14942 (N_14942,N_14499,N_14551);
nor U14943 (N_14943,N_14622,N_14510);
and U14944 (N_14944,N_14536,N_14657);
nor U14945 (N_14945,N_14471,N_14485);
or U14946 (N_14946,N_14568,N_14509);
or U14947 (N_14947,N_14523,N_14609);
xor U14948 (N_14948,N_14473,N_14427);
or U14949 (N_14949,N_14556,N_14408);
and U14950 (N_14950,N_14484,N_14431);
nand U14951 (N_14951,N_14517,N_14512);
nand U14952 (N_14952,N_14648,N_14599);
nor U14953 (N_14953,N_14432,N_14400);
xnor U14954 (N_14954,N_14573,N_14646);
nand U14955 (N_14955,N_14403,N_14488);
nand U14956 (N_14956,N_14524,N_14520);
nand U14957 (N_14957,N_14637,N_14570);
nor U14958 (N_14958,N_14650,N_14484);
and U14959 (N_14959,N_14664,N_14474);
nor U14960 (N_14960,N_14692,N_14501);
nand U14961 (N_14961,N_14523,N_14571);
or U14962 (N_14962,N_14659,N_14602);
nand U14963 (N_14963,N_14615,N_14614);
nor U14964 (N_14964,N_14630,N_14578);
nand U14965 (N_14965,N_14610,N_14501);
nor U14966 (N_14966,N_14542,N_14449);
nor U14967 (N_14967,N_14675,N_14678);
xnor U14968 (N_14968,N_14430,N_14469);
nand U14969 (N_14969,N_14682,N_14499);
and U14970 (N_14970,N_14699,N_14482);
or U14971 (N_14971,N_14559,N_14660);
nor U14972 (N_14972,N_14470,N_14667);
and U14973 (N_14973,N_14561,N_14535);
nor U14974 (N_14974,N_14439,N_14589);
nor U14975 (N_14975,N_14550,N_14665);
and U14976 (N_14976,N_14530,N_14699);
or U14977 (N_14977,N_14467,N_14524);
nor U14978 (N_14978,N_14578,N_14518);
xor U14979 (N_14979,N_14610,N_14480);
nor U14980 (N_14980,N_14543,N_14480);
nand U14981 (N_14981,N_14427,N_14636);
and U14982 (N_14982,N_14445,N_14450);
and U14983 (N_14983,N_14596,N_14419);
and U14984 (N_14984,N_14619,N_14622);
and U14985 (N_14985,N_14658,N_14428);
and U14986 (N_14986,N_14489,N_14541);
nor U14987 (N_14987,N_14506,N_14585);
xnor U14988 (N_14988,N_14412,N_14439);
nor U14989 (N_14989,N_14435,N_14612);
nand U14990 (N_14990,N_14611,N_14451);
nor U14991 (N_14991,N_14480,N_14468);
nand U14992 (N_14992,N_14534,N_14673);
nor U14993 (N_14993,N_14571,N_14507);
and U14994 (N_14994,N_14603,N_14577);
and U14995 (N_14995,N_14515,N_14454);
nor U14996 (N_14996,N_14431,N_14455);
xor U14997 (N_14997,N_14546,N_14680);
xor U14998 (N_14998,N_14547,N_14696);
nand U14999 (N_14999,N_14624,N_14689);
or UO_0 (O_0,N_14920,N_14977);
or UO_1 (O_1,N_14899,N_14776);
xor UO_2 (O_2,N_14746,N_14931);
nor UO_3 (O_3,N_14880,N_14989);
or UO_4 (O_4,N_14753,N_14855);
nor UO_5 (O_5,N_14806,N_14848);
nor UO_6 (O_6,N_14840,N_14883);
and UO_7 (O_7,N_14978,N_14781);
nor UO_8 (O_8,N_14739,N_14803);
nand UO_9 (O_9,N_14966,N_14956);
xor UO_10 (O_10,N_14711,N_14768);
nor UO_11 (O_11,N_14907,N_14816);
nor UO_12 (O_12,N_14859,N_14707);
xnor UO_13 (O_13,N_14844,N_14999);
nor UO_14 (O_14,N_14972,N_14908);
nand UO_15 (O_15,N_14827,N_14857);
or UO_16 (O_16,N_14773,N_14932);
xnor UO_17 (O_17,N_14981,N_14790);
nor UO_18 (O_18,N_14964,N_14729);
nor UO_19 (O_19,N_14872,N_14865);
and UO_20 (O_20,N_14847,N_14792);
nor UO_21 (O_21,N_14940,N_14846);
nand UO_22 (O_22,N_14703,N_14897);
and UO_23 (O_23,N_14736,N_14716);
or UO_24 (O_24,N_14722,N_14757);
xor UO_25 (O_25,N_14851,N_14946);
and UO_26 (O_26,N_14777,N_14706);
nor UO_27 (O_27,N_14864,N_14743);
or UO_28 (O_28,N_14747,N_14804);
xor UO_29 (O_29,N_14852,N_14950);
nand UO_30 (O_30,N_14766,N_14969);
or UO_31 (O_31,N_14962,N_14879);
xnor UO_32 (O_32,N_14836,N_14723);
xnor UO_33 (O_33,N_14884,N_14957);
xor UO_34 (O_34,N_14903,N_14991);
or UO_35 (O_35,N_14939,N_14927);
and UO_36 (O_36,N_14955,N_14784);
xor UO_37 (O_37,N_14876,N_14916);
nor UO_38 (O_38,N_14967,N_14944);
nor UO_39 (O_39,N_14718,N_14831);
and UO_40 (O_40,N_14982,N_14705);
or UO_41 (O_41,N_14772,N_14901);
or UO_42 (O_42,N_14719,N_14887);
nor UO_43 (O_43,N_14765,N_14724);
and UO_44 (O_44,N_14984,N_14839);
xor UO_45 (O_45,N_14900,N_14702);
xnor UO_46 (O_46,N_14789,N_14819);
xor UO_47 (O_47,N_14935,N_14938);
nor UO_48 (O_48,N_14878,N_14906);
and UO_49 (O_49,N_14821,N_14965);
nand UO_50 (O_50,N_14841,N_14986);
xor UO_51 (O_51,N_14904,N_14735);
and UO_52 (O_52,N_14800,N_14936);
nor UO_53 (O_53,N_14987,N_14814);
nor UO_54 (O_54,N_14783,N_14854);
xnor UO_55 (O_55,N_14763,N_14731);
or UO_56 (O_56,N_14820,N_14796);
and UO_57 (O_57,N_14813,N_14979);
nor UO_58 (O_58,N_14898,N_14959);
nand UO_59 (O_59,N_14912,N_14822);
nand UO_60 (O_60,N_14889,N_14795);
and UO_61 (O_61,N_14756,N_14873);
and UO_62 (O_62,N_14930,N_14874);
nand UO_63 (O_63,N_14801,N_14805);
nand UO_64 (O_64,N_14961,N_14951);
nor UO_65 (O_65,N_14993,N_14941);
and UO_66 (O_66,N_14910,N_14921);
nor UO_67 (O_67,N_14749,N_14922);
nor UO_68 (O_68,N_14885,N_14829);
nand UO_69 (O_69,N_14764,N_14737);
and UO_70 (O_70,N_14701,N_14871);
nor UO_71 (O_71,N_14728,N_14830);
xor UO_72 (O_72,N_14923,N_14849);
or UO_73 (O_73,N_14990,N_14960);
nand UO_74 (O_74,N_14748,N_14759);
nand UO_75 (O_75,N_14767,N_14917);
xnor UO_76 (O_76,N_14925,N_14882);
or UO_77 (O_77,N_14942,N_14755);
xor UO_78 (O_78,N_14905,N_14970);
or UO_79 (O_79,N_14933,N_14963);
and UO_80 (O_80,N_14915,N_14826);
nand UO_81 (O_81,N_14837,N_14771);
and UO_82 (O_82,N_14824,N_14875);
or UO_83 (O_83,N_14866,N_14797);
and UO_84 (O_84,N_14799,N_14947);
xor UO_85 (O_85,N_14863,N_14811);
xnor UO_86 (O_86,N_14919,N_14971);
and UO_87 (O_87,N_14918,N_14815);
nand UO_88 (O_88,N_14968,N_14778);
and UO_89 (O_89,N_14909,N_14850);
xor UO_90 (O_90,N_14785,N_14992);
and UO_91 (O_91,N_14974,N_14725);
or UO_92 (O_92,N_14937,N_14810);
xnor UO_93 (O_93,N_14709,N_14721);
nor UO_94 (O_94,N_14934,N_14998);
nand UO_95 (O_95,N_14708,N_14733);
nand UO_96 (O_96,N_14704,N_14752);
nand UO_97 (O_97,N_14954,N_14858);
or UO_98 (O_98,N_14712,N_14952);
nand UO_99 (O_99,N_14945,N_14754);
or UO_100 (O_100,N_14744,N_14953);
nand UO_101 (O_101,N_14741,N_14843);
or UO_102 (O_102,N_14994,N_14867);
nand UO_103 (O_103,N_14769,N_14761);
xor UO_104 (O_104,N_14845,N_14740);
nand UO_105 (O_105,N_14802,N_14958);
and UO_106 (O_106,N_14832,N_14782);
xnor UO_107 (O_107,N_14834,N_14787);
nand UO_108 (O_108,N_14794,N_14842);
nand UO_109 (O_109,N_14997,N_14988);
and UO_110 (O_110,N_14717,N_14809);
and UO_111 (O_111,N_14780,N_14825);
nand UO_112 (O_112,N_14896,N_14715);
and UO_113 (O_113,N_14877,N_14742);
or UO_114 (O_114,N_14714,N_14713);
or UO_115 (O_115,N_14817,N_14788);
xnor UO_116 (O_116,N_14976,N_14760);
or UO_117 (O_117,N_14975,N_14823);
and UO_118 (O_118,N_14818,N_14856);
or UO_119 (O_119,N_14861,N_14892);
xor UO_120 (O_120,N_14881,N_14996);
xor UO_121 (O_121,N_14774,N_14911);
xnor UO_122 (O_122,N_14983,N_14902);
and UO_123 (O_123,N_14732,N_14751);
nor UO_124 (O_124,N_14758,N_14980);
and UO_125 (O_125,N_14838,N_14828);
and UO_126 (O_126,N_14791,N_14869);
and UO_127 (O_127,N_14860,N_14745);
nor UO_128 (O_128,N_14913,N_14928);
and UO_129 (O_129,N_14973,N_14929);
or UO_130 (O_130,N_14793,N_14835);
nand UO_131 (O_131,N_14895,N_14807);
nor UO_132 (O_132,N_14924,N_14890);
nor UO_133 (O_133,N_14808,N_14886);
and UO_134 (O_134,N_14926,N_14985);
nor UO_135 (O_135,N_14700,N_14893);
nor UO_136 (O_136,N_14891,N_14888);
or UO_137 (O_137,N_14914,N_14779);
nand UO_138 (O_138,N_14738,N_14762);
and UO_139 (O_139,N_14786,N_14720);
nor UO_140 (O_140,N_14770,N_14862);
or UO_141 (O_141,N_14894,N_14949);
or UO_142 (O_142,N_14943,N_14853);
nor UO_143 (O_143,N_14775,N_14710);
nand UO_144 (O_144,N_14870,N_14995);
xor UO_145 (O_145,N_14833,N_14868);
or UO_146 (O_146,N_14726,N_14948);
and UO_147 (O_147,N_14734,N_14750);
nand UO_148 (O_148,N_14727,N_14798);
or UO_149 (O_149,N_14812,N_14730);
xor UO_150 (O_150,N_14906,N_14729);
or UO_151 (O_151,N_14786,N_14859);
nor UO_152 (O_152,N_14948,N_14814);
nor UO_153 (O_153,N_14872,N_14861);
or UO_154 (O_154,N_14984,N_14901);
and UO_155 (O_155,N_14821,N_14974);
and UO_156 (O_156,N_14837,N_14722);
or UO_157 (O_157,N_14706,N_14960);
or UO_158 (O_158,N_14764,N_14784);
nor UO_159 (O_159,N_14796,N_14781);
nand UO_160 (O_160,N_14994,N_14766);
nand UO_161 (O_161,N_14843,N_14836);
nand UO_162 (O_162,N_14904,N_14783);
and UO_163 (O_163,N_14856,N_14770);
nor UO_164 (O_164,N_14753,N_14981);
nand UO_165 (O_165,N_14726,N_14980);
and UO_166 (O_166,N_14988,N_14906);
xnor UO_167 (O_167,N_14931,N_14970);
or UO_168 (O_168,N_14709,N_14840);
and UO_169 (O_169,N_14884,N_14873);
nand UO_170 (O_170,N_14918,N_14844);
or UO_171 (O_171,N_14997,N_14789);
or UO_172 (O_172,N_14939,N_14842);
nand UO_173 (O_173,N_14795,N_14960);
or UO_174 (O_174,N_14810,N_14829);
nor UO_175 (O_175,N_14935,N_14713);
xnor UO_176 (O_176,N_14958,N_14787);
nor UO_177 (O_177,N_14728,N_14937);
or UO_178 (O_178,N_14952,N_14942);
and UO_179 (O_179,N_14805,N_14708);
or UO_180 (O_180,N_14855,N_14741);
nor UO_181 (O_181,N_14758,N_14700);
or UO_182 (O_182,N_14845,N_14808);
xnor UO_183 (O_183,N_14967,N_14753);
or UO_184 (O_184,N_14977,N_14861);
or UO_185 (O_185,N_14968,N_14802);
or UO_186 (O_186,N_14772,N_14728);
xor UO_187 (O_187,N_14825,N_14860);
nor UO_188 (O_188,N_14967,N_14716);
nand UO_189 (O_189,N_14735,N_14783);
and UO_190 (O_190,N_14982,N_14805);
nand UO_191 (O_191,N_14870,N_14912);
and UO_192 (O_192,N_14991,N_14937);
nand UO_193 (O_193,N_14946,N_14780);
and UO_194 (O_194,N_14765,N_14874);
and UO_195 (O_195,N_14981,N_14857);
and UO_196 (O_196,N_14857,N_14821);
nor UO_197 (O_197,N_14975,N_14774);
nand UO_198 (O_198,N_14849,N_14850);
nor UO_199 (O_199,N_14793,N_14784);
nor UO_200 (O_200,N_14852,N_14956);
or UO_201 (O_201,N_14910,N_14707);
nand UO_202 (O_202,N_14834,N_14931);
and UO_203 (O_203,N_14944,N_14734);
or UO_204 (O_204,N_14774,N_14714);
nand UO_205 (O_205,N_14781,N_14873);
nor UO_206 (O_206,N_14897,N_14879);
nor UO_207 (O_207,N_14955,N_14950);
xnor UO_208 (O_208,N_14940,N_14964);
or UO_209 (O_209,N_14946,N_14833);
and UO_210 (O_210,N_14779,N_14906);
nor UO_211 (O_211,N_14895,N_14754);
nand UO_212 (O_212,N_14886,N_14745);
xnor UO_213 (O_213,N_14921,N_14838);
xor UO_214 (O_214,N_14708,N_14756);
or UO_215 (O_215,N_14877,N_14823);
nor UO_216 (O_216,N_14942,N_14780);
or UO_217 (O_217,N_14850,N_14712);
and UO_218 (O_218,N_14880,N_14838);
or UO_219 (O_219,N_14767,N_14860);
nor UO_220 (O_220,N_14983,N_14811);
xnor UO_221 (O_221,N_14812,N_14930);
nor UO_222 (O_222,N_14987,N_14714);
nor UO_223 (O_223,N_14985,N_14872);
and UO_224 (O_224,N_14849,N_14936);
xor UO_225 (O_225,N_14705,N_14873);
and UO_226 (O_226,N_14985,N_14936);
xor UO_227 (O_227,N_14803,N_14984);
or UO_228 (O_228,N_14892,N_14760);
or UO_229 (O_229,N_14828,N_14735);
nor UO_230 (O_230,N_14882,N_14865);
or UO_231 (O_231,N_14700,N_14932);
xnor UO_232 (O_232,N_14731,N_14961);
and UO_233 (O_233,N_14866,N_14900);
and UO_234 (O_234,N_14718,N_14862);
xnor UO_235 (O_235,N_14757,N_14887);
and UO_236 (O_236,N_14860,N_14873);
nor UO_237 (O_237,N_14977,N_14772);
xnor UO_238 (O_238,N_14735,N_14728);
nand UO_239 (O_239,N_14867,N_14809);
nand UO_240 (O_240,N_14840,N_14926);
and UO_241 (O_241,N_14972,N_14742);
nand UO_242 (O_242,N_14862,N_14761);
or UO_243 (O_243,N_14737,N_14934);
or UO_244 (O_244,N_14977,N_14712);
nor UO_245 (O_245,N_14802,N_14947);
xnor UO_246 (O_246,N_14751,N_14968);
or UO_247 (O_247,N_14824,N_14848);
and UO_248 (O_248,N_14879,N_14912);
nor UO_249 (O_249,N_14836,N_14876);
nand UO_250 (O_250,N_14803,N_14712);
xor UO_251 (O_251,N_14740,N_14783);
nor UO_252 (O_252,N_14838,N_14751);
nor UO_253 (O_253,N_14749,N_14958);
or UO_254 (O_254,N_14774,N_14802);
nor UO_255 (O_255,N_14986,N_14817);
nand UO_256 (O_256,N_14812,N_14927);
nor UO_257 (O_257,N_14868,N_14736);
nand UO_258 (O_258,N_14887,N_14836);
nor UO_259 (O_259,N_14865,N_14943);
nor UO_260 (O_260,N_14956,N_14814);
nor UO_261 (O_261,N_14826,N_14769);
nand UO_262 (O_262,N_14946,N_14857);
nand UO_263 (O_263,N_14998,N_14752);
xor UO_264 (O_264,N_14748,N_14708);
or UO_265 (O_265,N_14923,N_14952);
xor UO_266 (O_266,N_14943,N_14838);
nand UO_267 (O_267,N_14711,N_14773);
nor UO_268 (O_268,N_14789,N_14909);
and UO_269 (O_269,N_14914,N_14805);
nor UO_270 (O_270,N_14846,N_14742);
nand UO_271 (O_271,N_14844,N_14743);
or UO_272 (O_272,N_14816,N_14752);
and UO_273 (O_273,N_14727,N_14728);
and UO_274 (O_274,N_14775,N_14903);
and UO_275 (O_275,N_14984,N_14931);
and UO_276 (O_276,N_14809,N_14775);
or UO_277 (O_277,N_14759,N_14955);
or UO_278 (O_278,N_14841,N_14897);
xor UO_279 (O_279,N_14873,N_14842);
and UO_280 (O_280,N_14767,N_14865);
nand UO_281 (O_281,N_14773,N_14822);
nor UO_282 (O_282,N_14730,N_14951);
nor UO_283 (O_283,N_14775,N_14788);
and UO_284 (O_284,N_14890,N_14829);
nand UO_285 (O_285,N_14828,N_14864);
nand UO_286 (O_286,N_14792,N_14848);
xor UO_287 (O_287,N_14909,N_14966);
or UO_288 (O_288,N_14874,N_14784);
nand UO_289 (O_289,N_14876,N_14933);
xor UO_290 (O_290,N_14884,N_14986);
nor UO_291 (O_291,N_14827,N_14745);
and UO_292 (O_292,N_14757,N_14894);
or UO_293 (O_293,N_14743,N_14929);
xor UO_294 (O_294,N_14858,N_14815);
or UO_295 (O_295,N_14778,N_14883);
or UO_296 (O_296,N_14835,N_14813);
xor UO_297 (O_297,N_14792,N_14787);
and UO_298 (O_298,N_14935,N_14970);
xor UO_299 (O_299,N_14795,N_14799);
xor UO_300 (O_300,N_14744,N_14924);
or UO_301 (O_301,N_14739,N_14898);
xor UO_302 (O_302,N_14781,N_14798);
nand UO_303 (O_303,N_14799,N_14753);
nand UO_304 (O_304,N_14971,N_14704);
nand UO_305 (O_305,N_14793,N_14944);
xnor UO_306 (O_306,N_14909,N_14937);
xor UO_307 (O_307,N_14929,N_14739);
xor UO_308 (O_308,N_14832,N_14920);
nand UO_309 (O_309,N_14946,N_14951);
nand UO_310 (O_310,N_14809,N_14721);
xor UO_311 (O_311,N_14912,N_14784);
xor UO_312 (O_312,N_14954,N_14822);
nand UO_313 (O_313,N_14897,N_14878);
or UO_314 (O_314,N_14747,N_14975);
or UO_315 (O_315,N_14814,N_14838);
or UO_316 (O_316,N_14928,N_14890);
nor UO_317 (O_317,N_14995,N_14881);
nand UO_318 (O_318,N_14793,N_14926);
nand UO_319 (O_319,N_14702,N_14803);
nor UO_320 (O_320,N_14795,N_14706);
xnor UO_321 (O_321,N_14740,N_14805);
xnor UO_322 (O_322,N_14893,N_14991);
xor UO_323 (O_323,N_14705,N_14902);
nand UO_324 (O_324,N_14852,N_14798);
nor UO_325 (O_325,N_14740,N_14879);
or UO_326 (O_326,N_14909,N_14727);
xor UO_327 (O_327,N_14813,N_14780);
or UO_328 (O_328,N_14775,N_14870);
nor UO_329 (O_329,N_14920,N_14913);
nand UO_330 (O_330,N_14792,N_14760);
nor UO_331 (O_331,N_14979,N_14940);
and UO_332 (O_332,N_14838,N_14733);
nor UO_333 (O_333,N_14804,N_14729);
xor UO_334 (O_334,N_14946,N_14895);
xor UO_335 (O_335,N_14829,N_14983);
or UO_336 (O_336,N_14942,N_14773);
and UO_337 (O_337,N_14963,N_14765);
or UO_338 (O_338,N_14864,N_14986);
and UO_339 (O_339,N_14710,N_14993);
nor UO_340 (O_340,N_14962,N_14894);
or UO_341 (O_341,N_14949,N_14877);
or UO_342 (O_342,N_14701,N_14950);
xor UO_343 (O_343,N_14779,N_14871);
xor UO_344 (O_344,N_14803,N_14819);
or UO_345 (O_345,N_14753,N_14750);
nand UO_346 (O_346,N_14778,N_14709);
nand UO_347 (O_347,N_14700,N_14891);
xnor UO_348 (O_348,N_14863,N_14720);
or UO_349 (O_349,N_14748,N_14738);
xnor UO_350 (O_350,N_14979,N_14962);
or UO_351 (O_351,N_14997,N_14828);
and UO_352 (O_352,N_14887,N_14766);
or UO_353 (O_353,N_14714,N_14855);
nand UO_354 (O_354,N_14955,N_14988);
nand UO_355 (O_355,N_14817,N_14949);
nand UO_356 (O_356,N_14977,N_14901);
and UO_357 (O_357,N_14954,N_14738);
or UO_358 (O_358,N_14966,N_14890);
nor UO_359 (O_359,N_14920,N_14711);
nor UO_360 (O_360,N_14831,N_14848);
xnor UO_361 (O_361,N_14848,N_14927);
or UO_362 (O_362,N_14766,N_14942);
or UO_363 (O_363,N_14969,N_14700);
xor UO_364 (O_364,N_14822,N_14942);
nand UO_365 (O_365,N_14969,N_14724);
nand UO_366 (O_366,N_14718,N_14887);
nor UO_367 (O_367,N_14702,N_14875);
or UO_368 (O_368,N_14875,N_14778);
and UO_369 (O_369,N_14870,N_14915);
or UO_370 (O_370,N_14886,N_14948);
nor UO_371 (O_371,N_14964,N_14996);
xor UO_372 (O_372,N_14955,N_14738);
or UO_373 (O_373,N_14766,N_14850);
and UO_374 (O_374,N_14736,N_14897);
nor UO_375 (O_375,N_14966,N_14907);
nand UO_376 (O_376,N_14798,N_14837);
nand UO_377 (O_377,N_14828,N_14800);
and UO_378 (O_378,N_14964,N_14868);
or UO_379 (O_379,N_14729,N_14826);
xor UO_380 (O_380,N_14897,N_14801);
nand UO_381 (O_381,N_14792,N_14767);
xor UO_382 (O_382,N_14707,N_14898);
nand UO_383 (O_383,N_14920,N_14786);
or UO_384 (O_384,N_14795,N_14745);
or UO_385 (O_385,N_14798,N_14850);
nor UO_386 (O_386,N_14785,N_14783);
or UO_387 (O_387,N_14863,N_14950);
or UO_388 (O_388,N_14793,N_14702);
nand UO_389 (O_389,N_14909,N_14849);
nand UO_390 (O_390,N_14932,N_14905);
nor UO_391 (O_391,N_14950,N_14916);
nor UO_392 (O_392,N_14738,N_14871);
nor UO_393 (O_393,N_14809,N_14923);
nor UO_394 (O_394,N_14942,N_14760);
nand UO_395 (O_395,N_14717,N_14744);
and UO_396 (O_396,N_14844,N_14723);
nor UO_397 (O_397,N_14781,N_14732);
nor UO_398 (O_398,N_14825,N_14984);
nor UO_399 (O_399,N_14757,N_14737);
or UO_400 (O_400,N_14832,N_14730);
and UO_401 (O_401,N_14991,N_14790);
and UO_402 (O_402,N_14868,N_14971);
nor UO_403 (O_403,N_14796,N_14895);
and UO_404 (O_404,N_14835,N_14777);
nand UO_405 (O_405,N_14913,N_14798);
and UO_406 (O_406,N_14700,N_14826);
nor UO_407 (O_407,N_14905,N_14980);
xor UO_408 (O_408,N_14844,N_14849);
or UO_409 (O_409,N_14904,N_14818);
xor UO_410 (O_410,N_14824,N_14997);
nand UO_411 (O_411,N_14967,N_14824);
xnor UO_412 (O_412,N_14736,N_14917);
or UO_413 (O_413,N_14830,N_14950);
and UO_414 (O_414,N_14801,N_14710);
xor UO_415 (O_415,N_14999,N_14873);
nand UO_416 (O_416,N_14766,N_14797);
and UO_417 (O_417,N_14972,N_14821);
xor UO_418 (O_418,N_14981,N_14836);
or UO_419 (O_419,N_14924,N_14806);
or UO_420 (O_420,N_14950,N_14911);
nand UO_421 (O_421,N_14718,N_14978);
and UO_422 (O_422,N_14945,N_14785);
nand UO_423 (O_423,N_14931,N_14804);
nor UO_424 (O_424,N_14829,N_14904);
xor UO_425 (O_425,N_14923,N_14991);
or UO_426 (O_426,N_14952,N_14763);
xor UO_427 (O_427,N_14780,N_14811);
nand UO_428 (O_428,N_14868,N_14923);
xnor UO_429 (O_429,N_14978,N_14923);
xnor UO_430 (O_430,N_14998,N_14884);
and UO_431 (O_431,N_14883,N_14757);
nor UO_432 (O_432,N_14712,N_14940);
or UO_433 (O_433,N_14717,N_14848);
and UO_434 (O_434,N_14837,N_14898);
nand UO_435 (O_435,N_14881,N_14747);
or UO_436 (O_436,N_14849,N_14981);
xor UO_437 (O_437,N_14876,N_14814);
nor UO_438 (O_438,N_14993,N_14795);
nor UO_439 (O_439,N_14863,N_14798);
or UO_440 (O_440,N_14834,N_14868);
or UO_441 (O_441,N_14730,N_14946);
nand UO_442 (O_442,N_14971,N_14775);
nand UO_443 (O_443,N_14992,N_14747);
and UO_444 (O_444,N_14954,N_14973);
and UO_445 (O_445,N_14755,N_14913);
and UO_446 (O_446,N_14851,N_14936);
and UO_447 (O_447,N_14851,N_14917);
and UO_448 (O_448,N_14968,N_14846);
nand UO_449 (O_449,N_14948,N_14884);
or UO_450 (O_450,N_14937,N_14971);
nand UO_451 (O_451,N_14745,N_14912);
nor UO_452 (O_452,N_14979,N_14878);
and UO_453 (O_453,N_14914,N_14775);
nor UO_454 (O_454,N_14736,N_14998);
nand UO_455 (O_455,N_14925,N_14885);
nand UO_456 (O_456,N_14790,N_14890);
and UO_457 (O_457,N_14827,N_14879);
nand UO_458 (O_458,N_14811,N_14744);
or UO_459 (O_459,N_14946,N_14885);
xor UO_460 (O_460,N_14908,N_14883);
nor UO_461 (O_461,N_14780,N_14899);
and UO_462 (O_462,N_14987,N_14838);
xor UO_463 (O_463,N_14865,N_14906);
or UO_464 (O_464,N_14738,N_14975);
xor UO_465 (O_465,N_14999,N_14932);
and UO_466 (O_466,N_14859,N_14933);
xnor UO_467 (O_467,N_14784,N_14909);
or UO_468 (O_468,N_14735,N_14901);
nand UO_469 (O_469,N_14765,N_14820);
or UO_470 (O_470,N_14926,N_14954);
xnor UO_471 (O_471,N_14730,N_14964);
xnor UO_472 (O_472,N_14885,N_14775);
xor UO_473 (O_473,N_14705,N_14760);
nand UO_474 (O_474,N_14732,N_14984);
nand UO_475 (O_475,N_14715,N_14841);
xnor UO_476 (O_476,N_14726,N_14911);
xnor UO_477 (O_477,N_14767,N_14758);
xor UO_478 (O_478,N_14760,N_14730);
xor UO_479 (O_479,N_14736,N_14875);
nand UO_480 (O_480,N_14979,N_14786);
or UO_481 (O_481,N_14849,N_14713);
or UO_482 (O_482,N_14966,N_14892);
nand UO_483 (O_483,N_14836,N_14825);
nand UO_484 (O_484,N_14703,N_14738);
nand UO_485 (O_485,N_14800,N_14837);
or UO_486 (O_486,N_14904,N_14985);
and UO_487 (O_487,N_14803,N_14814);
or UO_488 (O_488,N_14768,N_14824);
or UO_489 (O_489,N_14852,N_14793);
or UO_490 (O_490,N_14845,N_14964);
and UO_491 (O_491,N_14860,N_14735);
and UO_492 (O_492,N_14908,N_14807);
or UO_493 (O_493,N_14993,N_14905);
nand UO_494 (O_494,N_14856,N_14922);
nand UO_495 (O_495,N_14720,N_14766);
nand UO_496 (O_496,N_14703,N_14799);
or UO_497 (O_497,N_14893,N_14891);
or UO_498 (O_498,N_14919,N_14894);
or UO_499 (O_499,N_14965,N_14880);
nand UO_500 (O_500,N_14775,N_14980);
or UO_501 (O_501,N_14931,N_14885);
and UO_502 (O_502,N_14736,N_14801);
nand UO_503 (O_503,N_14853,N_14906);
or UO_504 (O_504,N_14811,N_14809);
nand UO_505 (O_505,N_14889,N_14725);
and UO_506 (O_506,N_14910,N_14702);
or UO_507 (O_507,N_14994,N_14797);
or UO_508 (O_508,N_14885,N_14784);
nand UO_509 (O_509,N_14788,N_14725);
nor UO_510 (O_510,N_14974,N_14808);
or UO_511 (O_511,N_14969,N_14867);
nor UO_512 (O_512,N_14778,N_14834);
or UO_513 (O_513,N_14722,N_14820);
nor UO_514 (O_514,N_14794,N_14770);
or UO_515 (O_515,N_14882,N_14714);
or UO_516 (O_516,N_14785,N_14867);
xor UO_517 (O_517,N_14701,N_14807);
xnor UO_518 (O_518,N_14949,N_14707);
or UO_519 (O_519,N_14854,N_14798);
and UO_520 (O_520,N_14873,N_14846);
or UO_521 (O_521,N_14738,N_14741);
or UO_522 (O_522,N_14872,N_14958);
xor UO_523 (O_523,N_14867,N_14998);
and UO_524 (O_524,N_14762,N_14714);
nand UO_525 (O_525,N_14711,N_14967);
nor UO_526 (O_526,N_14988,N_14939);
nor UO_527 (O_527,N_14835,N_14956);
and UO_528 (O_528,N_14959,N_14754);
nor UO_529 (O_529,N_14829,N_14883);
nand UO_530 (O_530,N_14967,N_14960);
nand UO_531 (O_531,N_14923,N_14782);
or UO_532 (O_532,N_14838,N_14715);
and UO_533 (O_533,N_14949,N_14722);
xnor UO_534 (O_534,N_14747,N_14963);
nand UO_535 (O_535,N_14726,N_14876);
xor UO_536 (O_536,N_14894,N_14834);
or UO_537 (O_537,N_14833,N_14952);
and UO_538 (O_538,N_14866,N_14711);
nor UO_539 (O_539,N_14878,N_14999);
or UO_540 (O_540,N_14993,N_14704);
or UO_541 (O_541,N_14750,N_14737);
nand UO_542 (O_542,N_14989,N_14836);
nor UO_543 (O_543,N_14800,N_14991);
or UO_544 (O_544,N_14972,N_14822);
nor UO_545 (O_545,N_14971,N_14715);
xor UO_546 (O_546,N_14881,N_14700);
nor UO_547 (O_547,N_14811,N_14888);
nand UO_548 (O_548,N_14843,N_14940);
nor UO_549 (O_549,N_14886,N_14859);
xor UO_550 (O_550,N_14929,N_14933);
and UO_551 (O_551,N_14993,N_14869);
and UO_552 (O_552,N_14822,N_14936);
xnor UO_553 (O_553,N_14941,N_14928);
nor UO_554 (O_554,N_14719,N_14889);
nor UO_555 (O_555,N_14810,N_14878);
xnor UO_556 (O_556,N_14958,N_14797);
nand UO_557 (O_557,N_14771,N_14871);
nor UO_558 (O_558,N_14906,N_14920);
nor UO_559 (O_559,N_14791,N_14715);
and UO_560 (O_560,N_14916,N_14812);
xor UO_561 (O_561,N_14832,N_14742);
nor UO_562 (O_562,N_14971,N_14819);
xor UO_563 (O_563,N_14729,N_14823);
or UO_564 (O_564,N_14819,N_14809);
or UO_565 (O_565,N_14952,N_14703);
and UO_566 (O_566,N_14957,N_14944);
nor UO_567 (O_567,N_14842,N_14712);
and UO_568 (O_568,N_14827,N_14761);
or UO_569 (O_569,N_14712,N_14942);
nor UO_570 (O_570,N_14738,N_14885);
or UO_571 (O_571,N_14792,N_14968);
nor UO_572 (O_572,N_14972,N_14804);
xor UO_573 (O_573,N_14750,N_14886);
xor UO_574 (O_574,N_14727,N_14784);
xor UO_575 (O_575,N_14903,N_14780);
nor UO_576 (O_576,N_14926,N_14920);
nand UO_577 (O_577,N_14842,N_14764);
and UO_578 (O_578,N_14815,N_14868);
nor UO_579 (O_579,N_14959,N_14903);
xnor UO_580 (O_580,N_14875,N_14752);
nand UO_581 (O_581,N_14744,N_14733);
xor UO_582 (O_582,N_14949,N_14872);
xnor UO_583 (O_583,N_14877,N_14873);
xor UO_584 (O_584,N_14741,N_14962);
or UO_585 (O_585,N_14760,N_14931);
xor UO_586 (O_586,N_14894,N_14797);
xor UO_587 (O_587,N_14769,N_14727);
nor UO_588 (O_588,N_14969,N_14916);
nor UO_589 (O_589,N_14732,N_14975);
xor UO_590 (O_590,N_14979,N_14944);
and UO_591 (O_591,N_14827,N_14833);
and UO_592 (O_592,N_14915,N_14861);
nand UO_593 (O_593,N_14943,N_14887);
xor UO_594 (O_594,N_14814,N_14933);
or UO_595 (O_595,N_14795,N_14861);
and UO_596 (O_596,N_14944,N_14878);
xnor UO_597 (O_597,N_14702,N_14976);
xnor UO_598 (O_598,N_14730,N_14942);
nand UO_599 (O_599,N_14924,N_14766);
and UO_600 (O_600,N_14733,N_14973);
and UO_601 (O_601,N_14713,N_14703);
xor UO_602 (O_602,N_14925,N_14706);
xnor UO_603 (O_603,N_14989,N_14916);
and UO_604 (O_604,N_14834,N_14747);
nand UO_605 (O_605,N_14800,N_14717);
nor UO_606 (O_606,N_14986,N_14870);
nand UO_607 (O_607,N_14888,N_14914);
nand UO_608 (O_608,N_14818,N_14999);
or UO_609 (O_609,N_14916,N_14869);
and UO_610 (O_610,N_14879,N_14987);
xnor UO_611 (O_611,N_14792,N_14757);
and UO_612 (O_612,N_14776,N_14785);
and UO_613 (O_613,N_14988,N_14774);
nand UO_614 (O_614,N_14757,N_14977);
and UO_615 (O_615,N_14725,N_14776);
nand UO_616 (O_616,N_14951,N_14808);
xnor UO_617 (O_617,N_14738,N_14908);
or UO_618 (O_618,N_14991,N_14761);
nand UO_619 (O_619,N_14926,N_14702);
nand UO_620 (O_620,N_14851,N_14803);
nand UO_621 (O_621,N_14798,N_14968);
nand UO_622 (O_622,N_14756,N_14826);
and UO_623 (O_623,N_14817,N_14732);
nand UO_624 (O_624,N_14726,N_14915);
xor UO_625 (O_625,N_14816,N_14709);
and UO_626 (O_626,N_14903,N_14854);
xnor UO_627 (O_627,N_14998,N_14799);
nor UO_628 (O_628,N_14890,N_14700);
nand UO_629 (O_629,N_14724,N_14952);
or UO_630 (O_630,N_14888,N_14978);
xor UO_631 (O_631,N_14782,N_14991);
xnor UO_632 (O_632,N_14883,N_14920);
or UO_633 (O_633,N_14707,N_14959);
nand UO_634 (O_634,N_14845,N_14943);
xnor UO_635 (O_635,N_14825,N_14778);
xor UO_636 (O_636,N_14877,N_14955);
or UO_637 (O_637,N_14891,N_14941);
xor UO_638 (O_638,N_14931,N_14770);
xor UO_639 (O_639,N_14854,N_14864);
nand UO_640 (O_640,N_14703,N_14996);
xor UO_641 (O_641,N_14703,N_14907);
nor UO_642 (O_642,N_14955,N_14743);
or UO_643 (O_643,N_14747,N_14791);
or UO_644 (O_644,N_14904,N_14756);
nor UO_645 (O_645,N_14773,N_14922);
xor UO_646 (O_646,N_14757,N_14920);
xor UO_647 (O_647,N_14878,N_14874);
nand UO_648 (O_648,N_14937,N_14779);
or UO_649 (O_649,N_14795,N_14905);
nand UO_650 (O_650,N_14849,N_14994);
nor UO_651 (O_651,N_14925,N_14906);
and UO_652 (O_652,N_14835,N_14868);
xor UO_653 (O_653,N_14798,N_14731);
or UO_654 (O_654,N_14727,N_14939);
nor UO_655 (O_655,N_14859,N_14944);
xor UO_656 (O_656,N_14787,N_14756);
nand UO_657 (O_657,N_14717,N_14835);
xor UO_658 (O_658,N_14961,N_14902);
nor UO_659 (O_659,N_14735,N_14997);
nand UO_660 (O_660,N_14780,N_14923);
nor UO_661 (O_661,N_14834,N_14925);
nor UO_662 (O_662,N_14921,N_14778);
or UO_663 (O_663,N_14764,N_14712);
nand UO_664 (O_664,N_14832,N_14870);
xor UO_665 (O_665,N_14771,N_14975);
or UO_666 (O_666,N_14953,N_14921);
nand UO_667 (O_667,N_14992,N_14875);
or UO_668 (O_668,N_14848,N_14753);
or UO_669 (O_669,N_14803,N_14858);
xnor UO_670 (O_670,N_14906,N_14889);
xnor UO_671 (O_671,N_14819,N_14805);
xor UO_672 (O_672,N_14936,N_14930);
nor UO_673 (O_673,N_14990,N_14945);
and UO_674 (O_674,N_14793,N_14983);
nand UO_675 (O_675,N_14938,N_14717);
or UO_676 (O_676,N_14861,N_14755);
nand UO_677 (O_677,N_14737,N_14928);
or UO_678 (O_678,N_14783,N_14846);
nor UO_679 (O_679,N_14759,N_14726);
xor UO_680 (O_680,N_14741,N_14998);
and UO_681 (O_681,N_14778,N_14879);
or UO_682 (O_682,N_14865,N_14892);
or UO_683 (O_683,N_14707,N_14711);
nor UO_684 (O_684,N_14985,N_14776);
or UO_685 (O_685,N_14742,N_14734);
nand UO_686 (O_686,N_14788,N_14846);
nor UO_687 (O_687,N_14760,N_14993);
or UO_688 (O_688,N_14972,N_14726);
or UO_689 (O_689,N_14892,N_14744);
and UO_690 (O_690,N_14994,N_14816);
nand UO_691 (O_691,N_14912,N_14917);
and UO_692 (O_692,N_14738,N_14883);
nor UO_693 (O_693,N_14811,N_14817);
nor UO_694 (O_694,N_14996,N_14962);
nand UO_695 (O_695,N_14860,N_14976);
and UO_696 (O_696,N_14828,N_14973);
xor UO_697 (O_697,N_14882,N_14970);
or UO_698 (O_698,N_14892,N_14729);
nor UO_699 (O_699,N_14896,N_14906);
nor UO_700 (O_700,N_14894,N_14968);
and UO_701 (O_701,N_14723,N_14708);
nand UO_702 (O_702,N_14967,N_14982);
nand UO_703 (O_703,N_14744,N_14864);
xor UO_704 (O_704,N_14940,N_14946);
and UO_705 (O_705,N_14889,N_14762);
and UO_706 (O_706,N_14974,N_14786);
nor UO_707 (O_707,N_14833,N_14931);
xnor UO_708 (O_708,N_14872,N_14797);
nand UO_709 (O_709,N_14835,N_14726);
xor UO_710 (O_710,N_14760,N_14700);
xor UO_711 (O_711,N_14897,N_14867);
and UO_712 (O_712,N_14961,N_14754);
or UO_713 (O_713,N_14719,N_14940);
nand UO_714 (O_714,N_14745,N_14911);
and UO_715 (O_715,N_14954,N_14734);
nand UO_716 (O_716,N_14890,N_14917);
nor UO_717 (O_717,N_14751,N_14893);
xnor UO_718 (O_718,N_14944,N_14963);
nand UO_719 (O_719,N_14872,N_14994);
xor UO_720 (O_720,N_14801,N_14746);
or UO_721 (O_721,N_14900,N_14715);
or UO_722 (O_722,N_14918,N_14814);
or UO_723 (O_723,N_14821,N_14786);
nand UO_724 (O_724,N_14819,N_14924);
nand UO_725 (O_725,N_14806,N_14748);
nand UO_726 (O_726,N_14976,N_14900);
or UO_727 (O_727,N_14945,N_14927);
and UO_728 (O_728,N_14856,N_14949);
xor UO_729 (O_729,N_14772,N_14975);
nor UO_730 (O_730,N_14753,N_14931);
xnor UO_731 (O_731,N_14904,N_14738);
xor UO_732 (O_732,N_14751,N_14930);
or UO_733 (O_733,N_14857,N_14954);
nand UO_734 (O_734,N_14735,N_14812);
or UO_735 (O_735,N_14808,N_14724);
xnor UO_736 (O_736,N_14903,N_14850);
and UO_737 (O_737,N_14785,N_14819);
nor UO_738 (O_738,N_14832,N_14940);
nand UO_739 (O_739,N_14842,N_14917);
or UO_740 (O_740,N_14813,N_14791);
xor UO_741 (O_741,N_14981,N_14957);
nor UO_742 (O_742,N_14866,N_14710);
and UO_743 (O_743,N_14754,N_14837);
nor UO_744 (O_744,N_14897,N_14988);
and UO_745 (O_745,N_14834,N_14870);
xor UO_746 (O_746,N_14809,N_14871);
nor UO_747 (O_747,N_14931,N_14737);
or UO_748 (O_748,N_14833,N_14753);
or UO_749 (O_749,N_14868,N_14935);
nor UO_750 (O_750,N_14736,N_14760);
nand UO_751 (O_751,N_14929,N_14709);
or UO_752 (O_752,N_14805,N_14834);
and UO_753 (O_753,N_14801,N_14999);
nor UO_754 (O_754,N_14892,N_14932);
xnor UO_755 (O_755,N_14878,N_14819);
xor UO_756 (O_756,N_14890,N_14782);
nand UO_757 (O_757,N_14739,N_14797);
nand UO_758 (O_758,N_14715,N_14714);
xor UO_759 (O_759,N_14780,N_14995);
xor UO_760 (O_760,N_14897,N_14959);
xor UO_761 (O_761,N_14825,N_14794);
or UO_762 (O_762,N_14787,N_14933);
or UO_763 (O_763,N_14729,N_14893);
or UO_764 (O_764,N_14827,N_14905);
nor UO_765 (O_765,N_14992,N_14760);
nand UO_766 (O_766,N_14946,N_14719);
xnor UO_767 (O_767,N_14811,N_14846);
nor UO_768 (O_768,N_14940,N_14763);
nor UO_769 (O_769,N_14877,N_14799);
xnor UO_770 (O_770,N_14739,N_14853);
and UO_771 (O_771,N_14932,N_14940);
or UO_772 (O_772,N_14860,N_14774);
xnor UO_773 (O_773,N_14761,N_14957);
nor UO_774 (O_774,N_14719,N_14804);
nor UO_775 (O_775,N_14936,N_14997);
nand UO_776 (O_776,N_14715,N_14773);
or UO_777 (O_777,N_14761,N_14773);
and UO_778 (O_778,N_14999,N_14955);
or UO_779 (O_779,N_14935,N_14949);
or UO_780 (O_780,N_14938,N_14986);
or UO_781 (O_781,N_14735,N_14743);
xor UO_782 (O_782,N_14940,N_14986);
nor UO_783 (O_783,N_14965,N_14944);
and UO_784 (O_784,N_14720,N_14715);
nor UO_785 (O_785,N_14720,N_14936);
nand UO_786 (O_786,N_14852,N_14824);
nor UO_787 (O_787,N_14915,N_14827);
xnor UO_788 (O_788,N_14736,N_14754);
nor UO_789 (O_789,N_14851,N_14744);
or UO_790 (O_790,N_14777,N_14788);
nor UO_791 (O_791,N_14985,N_14826);
xnor UO_792 (O_792,N_14955,N_14720);
xor UO_793 (O_793,N_14867,N_14731);
nor UO_794 (O_794,N_14746,N_14788);
or UO_795 (O_795,N_14802,N_14969);
nor UO_796 (O_796,N_14933,N_14865);
and UO_797 (O_797,N_14972,N_14871);
nand UO_798 (O_798,N_14709,N_14739);
and UO_799 (O_799,N_14866,N_14985);
xor UO_800 (O_800,N_14874,N_14899);
nand UO_801 (O_801,N_14823,N_14835);
or UO_802 (O_802,N_14930,N_14784);
and UO_803 (O_803,N_14801,N_14748);
xnor UO_804 (O_804,N_14980,N_14811);
or UO_805 (O_805,N_14802,N_14982);
or UO_806 (O_806,N_14818,N_14898);
and UO_807 (O_807,N_14734,N_14730);
nand UO_808 (O_808,N_14701,N_14801);
nand UO_809 (O_809,N_14884,N_14808);
and UO_810 (O_810,N_14750,N_14934);
nor UO_811 (O_811,N_14955,N_14733);
and UO_812 (O_812,N_14831,N_14924);
nor UO_813 (O_813,N_14750,N_14784);
nand UO_814 (O_814,N_14769,N_14743);
nand UO_815 (O_815,N_14838,N_14992);
or UO_816 (O_816,N_14763,N_14789);
xnor UO_817 (O_817,N_14963,N_14892);
or UO_818 (O_818,N_14971,N_14929);
and UO_819 (O_819,N_14873,N_14764);
or UO_820 (O_820,N_14914,N_14821);
nand UO_821 (O_821,N_14999,N_14970);
nand UO_822 (O_822,N_14828,N_14975);
and UO_823 (O_823,N_14925,N_14755);
nor UO_824 (O_824,N_14717,N_14755);
or UO_825 (O_825,N_14931,N_14742);
xor UO_826 (O_826,N_14771,N_14936);
and UO_827 (O_827,N_14710,N_14880);
or UO_828 (O_828,N_14730,N_14921);
or UO_829 (O_829,N_14722,N_14869);
nor UO_830 (O_830,N_14836,N_14982);
and UO_831 (O_831,N_14922,N_14911);
nor UO_832 (O_832,N_14881,N_14895);
or UO_833 (O_833,N_14735,N_14920);
xor UO_834 (O_834,N_14902,N_14764);
and UO_835 (O_835,N_14762,N_14841);
xnor UO_836 (O_836,N_14785,N_14742);
nand UO_837 (O_837,N_14778,N_14857);
and UO_838 (O_838,N_14992,N_14815);
and UO_839 (O_839,N_14972,N_14792);
or UO_840 (O_840,N_14817,N_14978);
or UO_841 (O_841,N_14973,N_14812);
and UO_842 (O_842,N_14845,N_14709);
and UO_843 (O_843,N_14842,N_14734);
nand UO_844 (O_844,N_14948,N_14706);
or UO_845 (O_845,N_14748,N_14876);
nor UO_846 (O_846,N_14791,N_14863);
nand UO_847 (O_847,N_14760,N_14982);
nand UO_848 (O_848,N_14785,N_14737);
or UO_849 (O_849,N_14790,N_14912);
and UO_850 (O_850,N_14708,N_14961);
xnor UO_851 (O_851,N_14802,N_14905);
or UO_852 (O_852,N_14878,N_14945);
or UO_853 (O_853,N_14702,N_14948);
xnor UO_854 (O_854,N_14904,N_14759);
xor UO_855 (O_855,N_14997,N_14985);
or UO_856 (O_856,N_14864,N_14907);
xor UO_857 (O_857,N_14774,N_14948);
nand UO_858 (O_858,N_14752,N_14932);
nor UO_859 (O_859,N_14745,N_14787);
nand UO_860 (O_860,N_14930,N_14788);
nor UO_861 (O_861,N_14729,N_14999);
nand UO_862 (O_862,N_14831,N_14899);
nand UO_863 (O_863,N_14848,N_14766);
or UO_864 (O_864,N_14999,N_14942);
or UO_865 (O_865,N_14762,N_14733);
xnor UO_866 (O_866,N_14936,N_14913);
xor UO_867 (O_867,N_14892,N_14974);
xor UO_868 (O_868,N_14793,N_14975);
nand UO_869 (O_869,N_14982,N_14720);
and UO_870 (O_870,N_14859,N_14860);
nor UO_871 (O_871,N_14809,N_14768);
nor UO_872 (O_872,N_14813,N_14872);
nor UO_873 (O_873,N_14830,N_14742);
nand UO_874 (O_874,N_14816,N_14906);
or UO_875 (O_875,N_14864,N_14936);
and UO_876 (O_876,N_14831,N_14951);
or UO_877 (O_877,N_14786,N_14817);
xor UO_878 (O_878,N_14753,N_14891);
or UO_879 (O_879,N_14756,N_14796);
nor UO_880 (O_880,N_14850,N_14790);
nor UO_881 (O_881,N_14806,N_14798);
xnor UO_882 (O_882,N_14939,N_14729);
nor UO_883 (O_883,N_14877,N_14874);
xnor UO_884 (O_884,N_14973,N_14841);
nand UO_885 (O_885,N_14952,N_14970);
nand UO_886 (O_886,N_14723,N_14889);
nor UO_887 (O_887,N_14977,N_14924);
and UO_888 (O_888,N_14870,N_14811);
xor UO_889 (O_889,N_14861,N_14907);
nor UO_890 (O_890,N_14985,N_14945);
xnor UO_891 (O_891,N_14701,N_14889);
xor UO_892 (O_892,N_14801,N_14757);
and UO_893 (O_893,N_14920,N_14704);
or UO_894 (O_894,N_14765,N_14726);
and UO_895 (O_895,N_14957,N_14862);
or UO_896 (O_896,N_14762,N_14891);
nand UO_897 (O_897,N_14781,N_14772);
nor UO_898 (O_898,N_14814,N_14887);
xor UO_899 (O_899,N_14755,N_14809);
nand UO_900 (O_900,N_14907,N_14850);
nand UO_901 (O_901,N_14862,N_14880);
nand UO_902 (O_902,N_14704,N_14974);
nand UO_903 (O_903,N_14887,N_14765);
nand UO_904 (O_904,N_14892,N_14717);
nor UO_905 (O_905,N_14983,N_14960);
nand UO_906 (O_906,N_14755,N_14779);
xnor UO_907 (O_907,N_14976,N_14963);
or UO_908 (O_908,N_14887,N_14931);
nor UO_909 (O_909,N_14815,N_14984);
and UO_910 (O_910,N_14979,N_14791);
xor UO_911 (O_911,N_14893,N_14839);
nand UO_912 (O_912,N_14971,N_14832);
nand UO_913 (O_913,N_14728,N_14807);
and UO_914 (O_914,N_14827,N_14997);
xor UO_915 (O_915,N_14712,N_14881);
nand UO_916 (O_916,N_14887,N_14796);
and UO_917 (O_917,N_14750,N_14739);
or UO_918 (O_918,N_14756,N_14958);
or UO_919 (O_919,N_14945,N_14956);
xnor UO_920 (O_920,N_14944,N_14897);
nand UO_921 (O_921,N_14824,N_14982);
xor UO_922 (O_922,N_14852,N_14853);
xnor UO_923 (O_923,N_14939,N_14828);
nand UO_924 (O_924,N_14765,N_14994);
nor UO_925 (O_925,N_14969,N_14740);
and UO_926 (O_926,N_14893,N_14755);
and UO_927 (O_927,N_14754,N_14785);
nand UO_928 (O_928,N_14737,N_14966);
or UO_929 (O_929,N_14998,N_14957);
nor UO_930 (O_930,N_14899,N_14884);
and UO_931 (O_931,N_14898,N_14830);
and UO_932 (O_932,N_14976,N_14812);
nor UO_933 (O_933,N_14765,N_14855);
nor UO_934 (O_934,N_14775,N_14777);
or UO_935 (O_935,N_14962,N_14814);
xor UO_936 (O_936,N_14957,N_14815);
and UO_937 (O_937,N_14886,N_14842);
nor UO_938 (O_938,N_14786,N_14835);
and UO_939 (O_939,N_14857,N_14742);
or UO_940 (O_940,N_14710,N_14809);
and UO_941 (O_941,N_14788,N_14766);
nand UO_942 (O_942,N_14705,N_14877);
and UO_943 (O_943,N_14788,N_14941);
nor UO_944 (O_944,N_14860,N_14708);
or UO_945 (O_945,N_14959,N_14846);
nand UO_946 (O_946,N_14829,N_14882);
and UO_947 (O_947,N_14807,N_14900);
xor UO_948 (O_948,N_14935,N_14871);
nand UO_949 (O_949,N_14858,N_14933);
and UO_950 (O_950,N_14800,N_14887);
or UO_951 (O_951,N_14722,N_14805);
xor UO_952 (O_952,N_14926,N_14809);
and UO_953 (O_953,N_14896,N_14899);
or UO_954 (O_954,N_14845,N_14901);
xor UO_955 (O_955,N_14794,N_14902);
xor UO_956 (O_956,N_14869,N_14878);
or UO_957 (O_957,N_14920,N_14903);
or UO_958 (O_958,N_14818,N_14884);
xor UO_959 (O_959,N_14858,N_14891);
nor UO_960 (O_960,N_14814,N_14926);
and UO_961 (O_961,N_14878,N_14903);
xnor UO_962 (O_962,N_14758,N_14893);
nand UO_963 (O_963,N_14846,N_14701);
nand UO_964 (O_964,N_14974,N_14942);
or UO_965 (O_965,N_14721,N_14964);
nand UO_966 (O_966,N_14859,N_14836);
and UO_967 (O_967,N_14875,N_14876);
nor UO_968 (O_968,N_14873,N_14893);
or UO_969 (O_969,N_14889,N_14877);
or UO_970 (O_970,N_14915,N_14886);
xnor UO_971 (O_971,N_14860,N_14945);
and UO_972 (O_972,N_14786,N_14842);
and UO_973 (O_973,N_14846,N_14807);
nor UO_974 (O_974,N_14701,N_14946);
xor UO_975 (O_975,N_14940,N_14990);
nand UO_976 (O_976,N_14981,N_14865);
nor UO_977 (O_977,N_14769,N_14846);
xnor UO_978 (O_978,N_14748,N_14980);
and UO_979 (O_979,N_14950,N_14945);
or UO_980 (O_980,N_14840,N_14992);
nand UO_981 (O_981,N_14713,N_14763);
nor UO_982 (O_982,N_14839,N_14881);
nand UO_983 (O_983,N_14745,N_14801);
xor UO_984 (O_984,N_14724,N_14711);
and UO_985 (O_985,N_14926,N_14907);
nand UO_986 (O_986,N_14768,N_14756);
nor UO_987 (O_987,N_14826,N_14781);
or UO_988 (O_988,N_14910,N_14836);
or UO_989 (O_989,N_14993,N_14802);
and UO_990 (O_990,N_14997,N_14820);
and UO_991 (O_991,N_14870,N_14747);
nor UO_992 (O_992,N_14856,N_14837);
nor UO_993 (O_993,N_14711,N_14976);
and UO_994 (O_994,N_14762,N_14756);
and UO_995 (O_995,N_14831,N_14735);
nor UO_996 (O_996,N_14718,N_14748);
nor UO_997 (O_997,N_14914,N_14977);
nor UO_998 (O_998,N_14914,N_14982);
nand UO_999 (O_999,N_14845,N_14779);
xor UO_1000 (O_1000,N_14826,N_14921);
nand UO_1001 (O_1001,N_14865,N_14843);
nor UO_1002 (O_1002,N_14942,N_14988);
nand UO_1003 (O_1003,N_14878,N_14965);
nor UO_1004 (O_1004,N_14990,N_14981);
and UO_1005 (O_1005,N_14829,N_14970);
nand UO_1006 (O_1006,N_14718,N_14830);
xnor UO_1007 (O_1007,N_14770,N_14917);
and UO_1008 (O_1008,N_14961,N_14774);
and UO_1009 (O_1009,N_14795,N_14963);
or UO_1010 (O_1010,N_14890,N_14820);
xor UO_1011 (O_1011,N_14823,N_14747);
nand UO_1012 (O_1012,N_14746,N_14992);
or UO_1013 (O_1013,N_14986,N_14857);
nand UO_1014 (O_1014,N_14795,N_14733);
and UO_1015 (O_1015,N_14780,N_14932);
nand UO_1016 (O_1016,N_14967,N_14791);
xnor UO_1017 (O_1017,N_14901,N_14805);
or UO_1018 (O_1018,N_14719,N_14911);
nand UO_1019 (O_1019,N_14700,N_14725);
or UO_1020 (O_1020,N_14993,N_14930);
nor UO_1021 (O_1021,N_14773,N_14787);
nor UO_1022 (O_1022,N_14877,N_14944);
xnor UO_1023 (O_1023,N_14950,N_14959);
nor UO_1024 (O_1024,N_14913,N_14757);
and UO_1025 (O_1025,N_14827,N_14843);
xor UO_1026 (O_1026,N_14940,N_14874);
xor UO_1027 (O_1027,N_14995,N_14872);
xnor UO_1028 (O_1028,N_14723,N_14869);
nor UO_1029 (O_1029,N_14724,N_14897);
nand UO_1030 (O_1030,N_14770,N_14898);
nand UO_1031 (O_1031,N_14875,N_14826);
nand UO_1032 (O_1032,N_14730,N_14708);
and UO_1033 (O_1033,N_14753,N_14739);
nor UO_1034 (O_1034,N_14789,N_14886);
nand UO_1035 (O_1035,N_14836,N_14907);
nand UO_1036 (O_1036,N_14995,N_14729);
nor UO_1037 (O_1037,N_14917,N_14844);
or UO_1038 (O_1038,N_14785,N_14877);
xor UO_1039 (O_1039,N_14988,N_14895);
or UO_1040 (O_1040,N_14943,N_14806);
xor UO_1041 (O_1041,N_14767,N_14704);
nand UO_1042 (O_1042,N_14749,N_14820);
or UO_1043 (O_1043,N_14993,N_14848);
xnor UO_1044 (O_1044,N_14851,N_14798);
and UO_1045 (O_1045,N_14760,N_14803);
nand UO_1046 (O_1046,N_14711,N_14726);
xor UO_1047 (O_1047,N_14731,N_14914);
xnor UO_1048 (O_1048,N_14952,N_14974);
or UO_1049 (O_1049,N_14812,N_14942);
nand UO_1050 (O_1050,N_14714,N_14723);
and UO_1051 (O_1051,N_14861,N_14700);
or UO_1052 (O_1052,N_14944,N_14752);
or UO_1053 (O_1053,N_14715,N_14973);
xnor UO_1054 (O_1054,N_14781,N_14716);
xor UO_1055 (O_1055,N_14987,N_14953);
xnor UO_1056 (O_1056,N_14997,N_14809);
or UO_1057 (O_1057,N_14865,N_14946);
nand UO_1058 (O_1058,N_14873,N_14795);
nor UO_1059 (O_1059,N_14934,N_14980);
xor UO_1060 (O_1060,N_14758,N_14753);
nand UO_1061 (O_1061,N_14706,N_14734);
nor UO_1062 (O_1062,N_14800,N_14707);
nor UO_1063 (O_1063,N_14993,N_14722);
nand UO_1064 (O_1064,N_14824,N_14851);
or UO_1065 (O_1065,N_14904,N_14991);
and UO_1066 (O_1066,N_14774,N_14918);
or UO_1067 (O_1067,N_14946,N_14803);
nor UO_1068 (O_1068,N_14844,N_14749);
xor UO_1069 (O_1069,N_14838,N_14796);
or UO_1070 (O_1070,N_14879,N_14863);
nand UO_1071 (O_1071,N_14965,N_14940);
and UO_1072 (O_1072,N_14706,N_14751);
nand UO_1073 (O_1073,N_14943,N_14791);
nand UO_1074 (O_1074,N_14835,N_14841);
xor UO_1075 (O_1075,N_14757,N_14718);
or UO_1076 (O_1076,N_14731,N_14984);
or UO_1077 (O_1077,N_14740,N_14974);
xnor UO_1078 (O_1078,N_14995,N_14889);
nand UO_1079 (O_1079,N_14794,N_14848);
and UO_1080 (O_1080,N_14705,N_14767);
nand UO_1081 (O_1081,N_14816,N_14975);
nor UO_1082 (O_1082,N_14706,N_14852);
and UO_1083 (O_1083,N_14827,N_14982);
or UO_1084 (O_1084,N_14977,N_14932);
xor UO_1085 (O_1085,N_14712,N_14773);
or UO_1086 (O_1086,N_14889,N_14741);
or UO_1087 (O_1087,N_14809,N_14804);
or UO_1088 (O_1088,N_14801,N_14866);
and UO_1089 (O_1089,N_14896,N_14720);
nor UO_1090 (O_1090,N_14868,N_14996);
nor UO_1091 (O_1091,N_14988,N_14786);
or UO_1092 (O_1092,N_14878,N_14779);
nor UO_1093 (O_1093,N_14863,N_14926);
or UO_1094 (O_1094,N_14775,N_14884);
or UO_1095 (O_1095,N_14851,N_14910);
or UO_1096 (O_1096,N_14732,N_14807);
nand UO_1097 (O_1097,N_14703,N_14779);
or UO_1098 (O_1098,N_14814,N_14857);
nor UO_1099 (O_1099,N_14982,N_14715);
and UO_1100 (O_1100,N_14791,N_14898);
nand UO_1101 (O_1101,N_14910,N_14872);
and UO_1102 (O_1102,N_14807,N_14845);
xnor UO_1103 (O_1103,N_14936,N_14717);
and UO_1104 (O_1104,N_14720,N_14835);
nand UO_1105 (O_1105,N_14992,N_14757);
nand UO_1106 (O_1106,N_14776,N_14996);
or UO_1107 (O_1107,N_14866,N_14911);
and UO_1108 (O_1108,N_14969,N_14921);
nand UO_1109 (O_1109,N_14957,N_14879);
and UO_1110 (O_1110,N_14947,N_14858);
and UO_1111 (O_1111,N_14963,N_14796);
xnor UO_1112 (O_1112,N_14896,N_14770);
nor UO_1113 (O_1113,N_14973,N_14820);
and UO_1114 (O_1114,N_14848,N_14739);
or UO_1115 (O_1115,N_14716,N_14871);
nor UO_1116 (O_1116,N_14902,N_14753);
xnor UO_1117 (O_1117,N_14951,N_14727);
nor UO_1118 (O_1118,N_14872,N_14816);
nor UO_1119 (O_1119,N_14844,N_14812);
nor UO_1120 (O_1120,N_14707,N_14817);
or UO_1121 (O_1121,N_14742,N_14813);
or UO_1122 (O_1122,N_14998,N_14790);
nor UO_1123 (O_1123,N_14942,N_14990);
or UO_1124 (O_1124,N_14814,N_14816);
xor UO_1125 (O_1125,N_14903,N_14908);
xnor UO_1126 (O_1126,N_14900,N_14714);
nor UO_1127 (O_1127,N_14949,N_14846);
nand UO_1128 (O_1128,N_14770,N_14924);
or UO_1129 (O_1129,N_14728,N_14878);
nand UO_1130 (O_1130,N_14805,N_14862);
or UO_1131 (O_1131,N_14758,N_14795);
or UO_1132 (O_1132,N_14901,N_14940);
nor UO_1133 (O_1133,N_14713,N_14900);
or UO_1134 (O_1134,N_14722,N_14724);
nor UO_1135 (O_1135,N_14820,N_14716);
nand UO_1136 (O_1136,N_14805,N_14842);
nand UO_1137 (O_1137,N_14800,N_14963);
or UO_1138 (O_1138,N_14954,N_14764);
nor UO_1139 (O_1139,N_14932,N_14723);
nand UO_1140 (O_1140,N_14762,N_14979);
and UO_1141 (O_1141,N_14713,N_14735);
nor UO_1142 (O_1142,N_14778,N_14964);
and UO_1143 (O_1143,N_14788,N_14980);
or UO_1144 (O_1144,N_14885,N_14811);
or UO_1145 (O_1145,N_14798,N_14774);
nand UO_1146 (O_1146,N_14918,N_14984);
xnor UO_1147 (O_1147,N_14701,N_14938);
nor UO_1148 (O_1148,N_14761,N_14826);
nor UO_1149 (O_1149,N_14912,N_14955);
or UO_1150 (O_1150,N_14790,N_14976);
nor UO_1151 (O_1151,N_14960,N_14834);
nor UO_1152 (O_1152,N_14878,N_14919);
or UO_1153 (O_1153,N_14999,N_14943);
or UO_1154 (O_1154,N_14737,N_14819);
xnor UO_1155 (O_1155,N_14898,N_14728);
nand UO_1156 (O_1156,N_14983,N_14955);
or UO_1157 (O_1157,N_14713,N_14771);
xor UO_1158 (O_1158,N_14892,N_14997);
or UO_1159 (O_1159,N_14790,N_14910);
xor UO_1160 (O_1160,N_14868,N_14723);
xnor UO_1161 (O_1161,N_14718,N_14805);
nand UO_1162 (O_1162,N_14862,N_14966);
xnor UO_1163 (O_1163,N_14976,N_14787);
nand UO_1164 (O_1164,N_14792,N_14913);
xnor UO_1165 (O_1165,N_14774,N_14902);
nor UO_1166 (O_1166,N_14947,N_14771);
nor UO_1167 (O_1167,N_14729,N_14718);
xor UO_1168 (O_1168,N_14750,N_14938);
xor UO_1169 (O_1169,N_14740,N_14826);
nor UO_1170 (O_1170,N_14770,N_14800);
nand UO_1171 (O_1171,N_14828,N_14718);
nor UO_1172 (O_1172,N_14867,N_14744);
nand UO_1173 (O_1173,N_14754,N_14979);
nor UO_1174 (O_1174,N_14711,N_14702);
nand UO_1175 (O_1175,N_14942,N_14907);
xor UO_1176 (O_1176,N_14799,N_14896);
nand UO_1177 (O_1177,N_14779,N_14922);
and UO_1178 (O_1178,N_14866,N_14812);
and UO_1179 (O_1179,N_14818,N_14755);
xor UO_1180 (O_1180,N_14987,N_14715);
nand UO_1181 (O_1181,N_14788,N_14738);
or UO_1182 (O_1182,N_14802,N_14816);
or UO_1183 (O_1183,N_14753,N_14961);
nand UO_1184 (O_1184,N_14778,N_14773);
or UO_1185 (O_1185,N_14948,N_14822);
xnor UO_1186 (O_1186,N_14868,N_14883);
and UO_1187 (O_1187,N_14883,N_14965);
nand UO_1188 (O_1188,N_14939,N_14707);
xnor UO_1189 (O_1189,N_14988,N_14740);
xnor UO_1190 (O_1190,N_14716,N_14760);
nor UO_1191 (O_1191,N_14897,N_14713);
and UO_1192 (O_1192,N_14950,N_14874);
nand UO_1193 (O_1193,N_14899,N_14892);
nand UO_1194 (O_1194,N_14841,N_14914);
xnor UO_1195 (O_1195,N_14819,N_14909);
nand UO_1196 (O_1196,N_14983,N_14790);
xor UO_1197 (O_1197,N_14971,N_14884);
nand UO_1198 (O_1198,N_14927,N_14867);
nand UO_1199 (O_1199,N_14950,N_14823);
or UO_1200 (O_1200,N_14932,N_14899);
and UO_1201 (O_1201,N_14712,N_14839);
or UO_1202 (O_1202,N_14915,N_14797);
nand UO_1203 (O_1203,N_14999,N_14977);
and UO_1204 (O_1204,N_14951,N_14995);
nor UO_1205 (O_1205,N_14783,N_14720);
or UO_1206 (O_1206,N_14960,N_14912);
xor UO_1207 (O_1207,N_14913,N_14737);
or UO_1208 (O_1208,N_14792,N_14912);
nand UO_1209 (O_1209,N_14710,N_14728);
xor UO_1210 (O_1210,N_14887,N_14795);
and UO_1211 (O_1211,N_14822,N_14932);
nand UO_1212 (O_1212,N_14774,N_14949);
xnor UO_1213 (O_1213,N_14952,N_14949);
nand UO_1214 (O_1214,N_14894,N_14811);
nand UO_1215 (O_1215,N_14720,N_14879);
nor UO_1216 (O_1216,N_14857,N_14793);
or UO_1217 (O_1217,N_14715,N_14731);
nand UO_1218 (O_1218,N_14809,N_14814);
xor UO_1219 (O_1219,N_14774,N_14965);
nand UO_1220 (O_1220,N_14825,N_14956);
nand UO_1221 (O_1221,N_14836,N_14794);
or UO_1222 (O_1222,N_14841,N_14970);
or UO_1223 (O_1223,N_14835,N_14985);
or UO_1224 (O_1224,N_14989,N_14704);
nand UO_1225 (O_1225,N_14901,N_14834);
nor UO_1226 (O_1226,N_14713,N_14773);
and UO_1227 (O_1227,N_14910,N_14825);
and UO_1228 (O_1228,N_14801,N_14938);
nand UO_1229 (O_1229,N_14932,N_14941);
and UO_1230 (O_1230,N_14727,N_14764);
xor UO_1231 (O_1231,N_14994,N_14777);
or UO_1232 (O_1232,N_14790,N_14963);
nand UO_1233 (O_1233,N_14747,N_14852);
and UO_1234 (O_1234,N_14931,N_14781);
and UO_1235 (O_1235,N_14766,N_14755);
or UO_1236 (O_1236,N_14960,N_14882);
nand UO_1237 (O_1237,N_14788,N_14844);
xnor UO_1238 (O_1238,N_14858,N_14756);
xnor UO_1239 (O_1239,N_14807,N_14748);
nand UO_1240 (O_1240,N_14883,N_14897);
and UO_1241 (O_1241,N_14707,N_14783);
xor UO_1242 (O_1242,N_14739,N_14994);
or UO_1243 (O_1243,N_14725,N_14714);
nor UO_1244 (O_1244,N_14844,N_14800);
xnor UO_1245 (O_1245,N_14967,N_14894);
or UO_1246 (O_1246,N_14751,N_14722);
xor UO_1247 (O_1247,N_14730,N_14723);
and UO_1248 (O_1248,N_14936,N_14955);
nand UO_1249 (O_1249,N_14874,N_14775);
nor UO_1250 (O_1250,N_14972,N_14886);
and UO_1251 (O_1251,N_14981,N_14928);
and UO_1252 (O_1252,N_14728,N_14964);
nor UO_1253 (O_1253,N_14805,N_14787);
nand UO_1254 (O_1254,N_14763,N_14978);
nor UO_1255 (O_1255,N_14876,N_14811);
and UO_1256 (O_1256,N_14902,N_14931);
nor UO_1257 (O_1257,N_14753,N_14922);
or UO_1258 (O_1258,N_14781,N_14735);
xor UO_1259 (O_1259,N_14903,N_14832);
or UO_1260 (O_1260,N_14999,N_14709);
nand UO_1261 (O_1261,N_14711,N_14986);
and UO_1262 (O_1262,N_14990,N_14743);
nand UO_1263 (O_1263,N_14823,N_14783);
nand UO_1264 (O_1264,N_14758,N_14732);
nand UO_1265 (O_1265,N_14975,N_14782);
or UO_1266 (O_1266,N_14768,N_14902);
nor UO_1267 (O_1267,N_14912,N_14854);
nor UO_1268 (O_1268,N_14725,N_14884);
or UO_1269 (O_1269,N_14850,N_14865);
xor UO_1270 (O_1270,N_14977,N_14915);
or UO_1271 (O_1271,N_14868,N_14986);
or UO_1272 (O_1272,N_14932,N_14796);
nand UO_1273 (O_1273,N_14948,N_14723);
and UO_1274 (O_1274,N_14762,N_14951);
nand UO_1275 (O_1275,N_14771,N_14794);
and UO_1276 (O_1276,N_14811,N_14951);
nand UO_1277 (O_1277,N_14753,N_14707);
nand UO_1278 (O_1278,N_14844,N_14820);
and UO_1279 (O_1279,N_14763,N_14986);
nor UO_1280 (O_1280,N_14722,N_14785);
or UO_1281 (O_1281,N_14811,N_14718);
nand UO_1282 (O_1282,N_14797,N_14843);
nand UO_1283 (O_1283,N_14716,N_14847);
nand UO_1284 (O_1284,N_14971,N_14928);
or UO_1285 (O_1285,N_14777,N_14725);
or UO_1286 (O_1286,N_14911,N_14947);
or UO_1287 (O_1287,N_14937,N_14876);
nor UO_1288 (O_1288,N_14763,N_14833);
nor UO_1289 (O_1289,N_14883,N_14885);
and UO_1290 (O_1290,N_14900,N_14935);
nand UO_1291 (O_1291,N_14912,N_14997);
nor UO_1292 (O_1292,N_14839,N_14758);
nand UO_1293 (O_1293,N_14885,N_14812);
xnor UO_1294 (O_1294,N_14946,N_14920);
xor UO_1295 (O_1295,N_14966,N_14916);
nand UO_1296 (O_1296,N_14823,N_14848);
nor UO_1297 (O_1297,N_14749,N_14792);
and UO_1298 (O_1298,N_14708,N_14844);
nand UO_1299 (O_1299,N_14861,N_14830);
or UO_1300 (O_1300,N_14719,N_14890);
and UO_1301 (O_1301,N_14748,N_14863);
or UO_1302 (O_1302,N_14828,N_14748);
xor UO_1303 (O_1303,N_14878,N_14893);
xor UO_1304 (O_1304,N_14856,N_14903);
xor UO_1305 (O_1305,N_14719,N_14999);
nor UO_1306 (O_1306,N_14734,N_14860);
nor UO_1307 (O_1307,N_14783,N_14756);
nand UO_1308 (O_1308,N_14928,N_14832);
nor UO_1309 (O_1309,N_14715,N_14706);
and UO_1310 (O_1310,N_14800,N_14939);
nor UO_1311 (O_1311,N_14938,N_14885);
or UO_1312 (O_1312,N_14864,N_14928);
xnor UO_1313 (O_1313,N_14975,N_14794);
or UO_1314 (O_1314,N_14957,N_14889);
nor UO_1315 (O_1315,N_14884,N_14972);
or UO_1316 (O_1316,N_14885,N_14777);
or UO_1317 (O_1317,N_14891,N_14880);
nand UO_1318 (O_1318,N_14856,N_14793);
xor UO_1319 (O_1319,N_14866,N_14947);
xor UO_1320 (O_1320,N_14869,N_14856);
xnor UO_1321 (O_1321,N_14781,N_14963);
and UO_1322 (O_1322,N_14898,N_14806);
xor UO_1323 (O_1323,N_14846,N_14948);
xor UO_1324 (O_1324,N_14937,N_14709);
xnor UO_1325 (O_1325,N_14787,N_14785);
nor UO_1326 (O_1326,N_14926,N_14870);
nor UO_1327 (O_1327,N_14980,N_14708);
or UO_1328 (O_1328,N_14747,N_14728);
nand UO_1329 (O_1329,N_14738,N_14833);
nor UO_1330 (O_1330,N_14881,N_14835);
and UO_1331 (O_1331,N_14867,N_14702);
or UO_1332 (O_1332,N_14958,N_14913);
nand UO_1333 (O_1333,N_14913,N_14880);
and UO_1334 (O_1334,N_14808,N_14759);
and UO_1335 (O_1335,N_14921,N_14755);
nor UO_1336 (O_1336,N_14719,N_14900);
nor UO_1337 (O_1337,N_14855,N_14867);
nor UO_1338 (O_1338,N_14888,N_14734);
and UO_1339 (O_1339,N_14787,N_14955);
nand UO_1340 (O_1340,N_14819,N_14914);
xor UO_1341 (O_1341,N_14979,N_14854);
nor UO_1342 (O_1342,N_14813,N_14958);
or UO_1343 (O_1343,N_14832,N_14931);
and UO_1344 (O_1344,N_14900,N_14762);
or UO_1345 (O_1345,N_14874,N_14835);
or UO_1346 (O_1346,N_14877,N_14818);
nor UO_1347 (O_1347,N_14985,N_14944);
or UO_1348 (O_1348,N_14740,N_14828);
and UO_1349 (O_1349,N_14984,N_14810);
nand UO_1350 (O_1350,N_14947,N_14710);
and UO_1351 (O_1351,N_14928,N_14990);
and UO_1352 (O_1352,N_14819,N_14715);
nand UO_1353 (O_1353,N_14998,N_14748);
or UO_1354 (O_1354,N_14766,N_14968);
nor UO_1355 (O_1355,N_14844,N_14923);
xnor UO_1356 (O_1356,N_14728,N_14819);
xnor UO_1357 (O_1357,N_14779,N_14753);
and UO_1358 (O_1358,N_14957,N_14892);
nand UO_1359 (O_1359,N_14715,N_14972);
and UO_1360 (O_1360,N_14707,N_14905);
and UO_1361 (O_1361,N_14789,N_14974);
xor UO_1362 (O_1362,N_14990,N_14973);
nand UO_1363 (O_1363,N_14778,N_14972);
and UO_1364 (O_1364,N_14772,N_14966);
nor UO_1365 (O_1365,N_14790,N_14828);
or UO_1366 (O_1366,N_14884,N_14744);
xnor UO_1367 (O_1367,N_14887,N_14973);
or UO_1368 (O_1368,N_14888,N_14849);
or UO_1369 (O_1369,N_14994,N_14907);
and UO_1370 (O_1370,N_14717,N_14843);
nor UO_1371 (O_1371,N_14904,N_14745);
and UO_1372 (O_1372,N_14732,N_14705);
xor UO_1373 (O_1373,N_14951,N_14945);
and UO_1374 (O_1374,N_14905,N_14733);
or UO_1375 (O_1375,N_14963,N_14813);
and UO_1376 (O_1376,N_14856,N_14861);
nand UO_1377 (O_1377,N_14700,N_14859);
or UO_1378 (O_1378,N_14901,N_14942);
nand UO_1379 (O_1379,N_14901,N_14854);
nor UO_1380 (O_1380,N_14723,N_14980);
nor UO_1381 (O_1381,N_14877,N_14863);
nor UO_1382 (O_1382,N_14819,N_14984);
or UO_1383 (O_1383,N_14989,N_14778);
nor UO_1384 (O_1384,N_14832,N_14929);
or UO_1385 (O_1385,N_14928,N_14780);
or UO_1386 (O_1386,N_14779,N_14967);
nand UO_1387 (O_1387,N_14713,N_14792);
xnor UO_1388 (O_1388,N_14724,N_14838);
xor UO_1389 (O_1389,N_14828,N_14719);
xnor UO_1390 (O_1390,N_14773,N_14833);
or UO_1391 (O_1391,N_14845,N_14704);
or UO_1392 (O_1392,N_14841,N_14979);
and UO_1393 (O_1393,N_14789,N_14941);
xnor UO_1394 (O_1394,N_14831,N_14999);
or UO_1395 (O_1395,N_14835,N_14771);
nand UO_1396 (O_1396,N_14877,N_14780);
nand UO_1397 (O_1397,N_14840,N_14950);
nand UO_1398 (O_1398,N_14714,N_14707);
and UO_1399 (O_1399,N_14999,N_14875);
xor UO_1400 (O_1400,N_14754,N_14709);
and UO_1401 (O_1401,N_14845,N_14794);
nor UO_1402 (O_1402,N_14938,N_14709);
nand UO_1403 (O_1403,N_14790,N_14954);
xnor UO_1404 (O_1404,N_14810,N_14873);
xnor UO_1405 (O_1405,N_14828,N_14879);
or UO_1406 (O_1406,N_14727,N_14749);
and UO_1407 (O_1407,N_14924,N_14942);
or UO_1408 (O_1408,N_14917,N_14854);
or UO_1409 (O_1409,N_14796,N_14956);
nand UO_1410 (O_1410,N_14848,N_14890);
nand UO_1411 (O_1411,N_14769,N_14819);
xnor UO_1412 (O_1412,N_14911,N_14729);
nand UO_1413 (O_1413,N_14979,N_14990);
nand UO_1414 (O_1414,N_14728,N_14971);
and UO_1415 (O_1415,N_14961,N_14791);
xor UO_1416 (O_1416,N_14763,N_14839);
nor UO_1417 (O_1417,N_14839,N_14767);
or UO_1418 (O_1418,N_14809,N_14996);
or UO_1419 (O_1419,N_14995,N_14714);
or UO_1420 (O_1420,N_14847,N_14927);
nor UO_1421 (O_1421,N_14734,N_14985);
xnor UO_1422 (O_1422,N_14760,N_14934);
nor UO_1423 (O_1423,N_14828,N_14794);
xnor UO_1424 (O_1424,N_14739,N_14894);
nor UO_1425 (O_1425,N_14852,N_14898);
xor UO_1426 (O_1426,N_14932,N_14787);
xor UO_1427 (O_1427,N_14990,N_14716);
xnor UO_1428 (O_1428,N_14849,N_14808);
nand UO_1429 (O_1429,N_14945,N_14827);
nor UO_1430 (O_1430,N_14862,N_14841);
xor UO_1431 (O_1431,N_14905,N_14814);
nand UO_1432 (O_1432,N_14913,N_14775);
nand UO_1433 (O_1433,N_14819,N_14926);
nor UO_1434 (O_1434,N_14972,N_14952);
and UO_1435 (O_1435,N_14832,N_14866);
and UO_1436 (O_1436,N_14849,N_14726);
xor UO_1437 (O_1437,N_14777,N_14836);
nor UO_1438 (O_1438,N_14982,N_14707);
or UO_1439 (O_1439,N_14903,N_14723);
nor UO_1440 (O_1440,N_14730,N_14805);
nand UO_1441 (O_1441,N_14922,N_14861);
xnor UO_1442 (O_1442,N_14799,N_14777);
or UO_1443 (O_1443,N_14789,N_14804);
nor UO_1444 (O_1444,N_14877,N_14773);
nand UO_1445 (O_1445,N_14820,N_14781);
xor UO_1446 (O_1446,N_14817,N_14880);
xnor UO_1447 (O_1447,N_14862,N_14849);
nand UO_1448 (O_1448,N_14777,N_14813);
nor UO_1449 (O_1449,N_14924,N_14966);
nand UO_1450 (O_1450,N_14796,N_14765);
nor UO_1451 (O_1451,N_14726,N_14738);
and UO_1452 (O_1452,N_14913,N_14723);
nand UO_1453 (O_1453,N_14759,N_14749);
and UO_1454 (O_1454,N_14926,N_14804);
nor UO_1455 (O_1455,N_14792,N_14997);
xnor UO_1456 (O_1456,N_14944,N_14748);
and UO_1457 (O_1457,N_14759,N_14990);
or UO_1458 (O_1458,N_14749,N_14735);
or UO_1459 (O_1459,N_14766,N_14918);
or UO_1460 (O_1460,N_14931,N_14844);
nor UO_1461 (O_1461,N_14708,N_14845);
or UO_1462 (O_1462,N_14896,N_14990);
nor UO_1463 (O_1463,N_14782,N_14708);
or UO_1464 (O_1464,N_14821,N_14852);
or UO_1465 (O_1465,N_14765,N_14790);
or UO_1466 (O_1466,N_14726,N_14732);
nor UO_1467 (O_1467,N_14824,N_14753);
and UO_1468 (O_1468,N_14976,N_14707);
xor UO_1469 (O_1469,N_14771,N_14878);
and UO_1470 (O_1470,N_14985,N_14823);
nand UO_1471 (O_1471,N_14706,N_14790);
nand UO_1472 (O_1472,N_14958,N_14706);
nand UO_1473 (O_1473,N_14825,N_14957);
or UO_1474 (O_1474,N_14852,N_14743);
xor UO_1475 (O_1475,N_14941,N_14817);
and UO_1476 (O_1476,N_14846,N_14816);
or UO_1477 (O_1477,N_14917,N_14759);
xnor UO_1478 (O_1478,N_14938,N_14766);
nor UO_1479 (O_1479,N_14997,N_14962);
xnor UO_1480 (O_1480,N_14873,N_14840);
nand UO_1481 (O_1481,N_14823,N_14923);
nor UO_1482 (O_1482,N_14819,N_14712);
nor UO_1483 (O_1483,N_14911,N_14918);
xnor UO_1484 (O_1484,N_14976,N_14978);
or UO_1485 (O_1485,N_14993,N_14779);
and UO_1486 (O_1486,N_14938,N_14855);
or UO_1487 (O_1487,N_14703,N_14993);
xor UO_1488 (O_1488,N_14813,N_14927);
nor UO_1489 (O_1489,N_14856,N_14784);
xnor UO_1490 (O_1490,N_14760,N_14949);
xnor UO_1491 (O_1491,N_14702,N_14857);
and UO_1492 (O_1492,N_14730,N_14935);
and UO_1493 (O_1493,N_14989,N_14936);
nand UO_1494 (O_1494,N_14925,N_14777);
nor UO_1495 (O_1495,N_14741,N_14909);
nor UO_1496 (O_1496,N_14988,N_14808);
or UO_1497 (O_1497,N_14773,N_14851);
nand UO_1498 (O_1498,N_14718,N_14951);
nand UO_1499 (O_1499,N_14730,N_14875);
xor UO_1500 (O_1500,N_14784,N_14929);
and UO_1501 (O_1501,N_14742,N_14844);
nand UO_1502 (O_1502,N_14809,N_14728);
and UO_1503 (O_1503,N_14963,N_14730);
and UO_1504 (O_1504,N_14787,N_14972);
and UO_1505 (O_1505,N_14936,N_14725);
or UO_1506 (O_1506,N_14842,N_14752);
nand UO_1507 (O_1507,N_14908,N_14811);
xor UO_1508 (O_1508,N_14920,N_14957);
nand UO_1509 (O_1509,N_14895,N_14743);
nor UO_1510 (O_1510,N_14711,N_14991);
xor UO_1511 (O_1511,N_14852,N_14963);
nand UO_1512 (O_1512,N_14791,N_14720);
nand UO_1513 (O_1513,N_14994,N_14869);
or UO_1514 (O_1514,N_14777,N_14825);
nand UO_1515 (O_1515,N_14981,N_14886);
nor UO_1516 (O_1516,N_14781,N_14944);
and UO_1517 (O_1517,N_14889,N_14982);
and UO_1518 (O_1518,N_14986,N_14781);
xnor UO_1519 (O_1519,N_14724,N_14757);
nand UO_1520 (O_1520,N_14831,N_14885);
nor UO_1521 (O_1521,N_14814,N_14839);
and UO_1522 (O_1522,N_14856,N_14759);
nand UO_1523 (O_1523,N_14884,N_14966);
nand UO_1524 (O_1524,N_14833,N_14849);
nand UO_1525 (O_1525,N_14854,N_14711);
nor UO_1526 (O_1526,N_14959,N_14789);
xor UO_1527 (O_1527,N_14867,N_14941);
nor UO_1528 (O_1528,N_14828,N_14795);
nand UO_1529 (O_1529,N_14987,N_14920);
and UO_1530 (O_1530,N_14958,N_14774);
nor UO_1531 (O_1531,N_14983,N_14832);
nand UO_1532 (O_1532,N_14790,N_14787);
nand UO_1533 (O_1533,N_14985,N_14903);
or UO_1534 (O_1534,N_14995,N_14926);
or UO_1535 (O_1535,N_14789,N_14707);
and UO_1536 (O_1536,N_14816,N_14714);
nor UO_1537 (O_1537,N_14800,N_14700);
nand UO_1538 (O_1538,N_14756,N_14966);
nor UO_1539 (O_1539,N_14818,N_14858);
and UO_1540 (O_1540,N_14748,N_14939);
or UO_1541 (O_1541,N_14749,N_14771);
or UO_1542 (O_1542,N_14702,N_14782);
or UO_1543 (O_1543,N_14990,N_14787);
nand UO_1544 (O_1544,N_14969,N_14995);
and UO_1545 (O_1545,N_14978,N_14865);
xor UO_1546 (O_1546,N_14909,N_14723);
or UO_1547 (O_1547,N_14770,N_14797);
xor UO_1548 (O_1548,N_14893,N_14795);
and UO_1549 (O_1549,N_14783,N_14885);
and UO_1550 (O_1550,N_14986,N_14946);
nor UO_1551 (O_1551,N_14930,N_14909);
nand UO_1552 (O_1552,N_14986,N_14875);
xor UO_1553 (O_1553,N_14841,N_14997);
or UO_1554 (O_1554,N_14704,N_14706);
xor UO_1555 (O_1555,N_14855,N_14768);
nor UO_1556 (O_1556,N_14997,N_14999);
nand UO_1557 (O_1557,N_14817,N_14825);
xor UO_1558 (O_1558,N_14797,N_14871);
xnor UO_1559 (O_1559,N_14739,N_14832);
nand UO_1560 (O_1560,N_14867,N_14750);
nand UO_1561 (O_1561,N_14701,N_14901);
xor UO_1562 (O_1562,N_14844,N_14875);
and UO_1563 (O_1563,N_14850,N_14942);
or UO_1564 (O_1564,N_14827,N_14815);
or UO_1565 (O_1565,N_14991,N_14710);
xor UO_1566 (O_1566,N_14809,N_14980);
nand UO_1567 (O_1567,N_14852,N_14773);
nand UO_1568 (O_1568,N_14737,N_14818);
or UO_1569 (O_1569,N_14941,N_14749);
xor UO_1570 (O_1570,N_14718,N_14966);
nor UO_1571 (O_1571,N_14708,N_14971);
nand UO_1572 (O_1572,N_14890,N_14703);
nand UO_1573 (O_1573,N_14743,N_14824);
or UO_1574 (O_1574,N_14760,N_14959);
nor UO_1575 (O_1575,N_14815,N_14917);
xnor UO_1576 (O_1576,N_14969,N_14915);
or UO_1577 (O_1577,N_14819,N_14893);
nand UO_1578 (O_1578,N_14734,N_14722);
xor UO_1579 (O_1579,N_14792,N_14727);
nand UO_1580 (O_1580,N_14707,N_14937);
or UO_1581 (O_1581,N_14714,N_14736);
xnor UO_1582 (O_1582,N_14707,N_14824);
and UO_1583 (O_1583,N_14835,N_14778);
xor UO_1584 (O_1584,N_14924,N_14767);
or UO_1585 (O_1585,N_14838,N_14790);
or UO_1586 (O_1586,N_14949,N_14862);
and UO_1587 (O_1587,N_14709,N_14873);
nand UO_1588 (O_1588,N_14852,N_14713);
nand UO_1589 (O_1589,N_14849,N_14880);
or UO_1590 (O_1590,N_14792,N_14991);
nor UO_1591 (O_1591,N_14808,N_14722);
or UO_1592 (O_1592,N_14958,N_14822);
nor UO_1593 (O_1593,N_14965,N_14954);
or UO_1594 (O_1594,N_14808,N_14858);
nand UO_1595 (O_1595,N_14935,N_14996);
nor UO_1596 (O_1596,N_14725,N_14774);
or UO_1597 (O_1597,N_14996,N_14760);
xor UO_1598 (O_1598,N_14963,N_14988);
nand UO_1599 (O_1599,N_14877,N_14716);
xnor UO_1600 (O_1600,N_14921,N_14917);
and UO_1601 (O_1601,N_14886,N_14922);
and UO_1602 (O_1602,N_14771,N_14998);
or UO_1603 (O_1603,N_14864,N_14861);
nor UO_1604 (O_1604,N_14864,N_14952);
or UO_1605 (O_1605,N_14708,N_14913);
xnor UO_1606 (O_1606,N_14937,N_14934);
and UO_1607 (O_1607,N_14929,N_14729);
xor UO_1608 (O_1608,N_14949,N_14890);
or UO_1609 (O_1609,N_14982,N_14893);
nor UO_1610 (O_1610,N_14707,N_14847);
or UO_1611 (O_1611,N_14904,N_14917);
xor UO_1612 (O_1612,N_14780,N_14974);
nor UO_1613 (O_1613,N_14763,N_14968);
or UO_1614 (O_1614,N_14981,N_14749);
xnor UO_1615 (O_1615,N_14721,N_14847);
or UO_1616 (O_1616,N_14999,N_14780);
or UO_1617 (O_1617,N_14908,N_14799);
or UO_1618 (O_1618,N_14855,N_14769);
nand UO_1619 (O_1619,N_14953,N_14942);
xnor UO_1620 (O_1620,N_14711,N_14926);
and UO_1621 (O_1621,N_14958,N_14876);
and UO_1622 (O_1622,N_14925,N_14959);
and UO_1623 (O_1623,N_14864,N_14731);
nor UO_1624 (O_1624,N_14875,N_14905);
nand UO_1625 (O_1625,N_14753,N_14910);
or UO_1626 (O_1626,N_14719,N_14861);
or UO_1627 (O_1627,N_14957,N_14852);
and UO_1628 (O_1628,N_14931,N_14779);
and UO_1629 (O_1629,N_14939,N_14867);
xnor UO_1630 (O_1630,N_14777,N_14827);
or UO_1631 (O_1631,N_14858,N_14831);
xnor UO_1632 (O_1632,N_14753,N_14725);
nand UO_1633 (O_1633,N_14944,N_14836);
or UO_1634 (O_1634,N_14885,N_14989);
nor UO_1635 (O_1635,N_14876,N_14950);
and UO_1636 (O_1636,N_14778,N_14970);
nand UO_1637 (O_1637,N_14928,N_14756);
xor UO_1638 (O_1638,N_14749,N_14787);
xnor UO_1639 (O_1639,N_14740,N_14864);
nor UO_1640 (O_1640,N_14973,N_14963);
or UO_1641 (O_1641,N_14943,N_14751);
and UO_1642 (O_1642,N_14850,N_14839);
or UO_1643 (O_1643,N_14767,N_14712);
nor UO_1644 (O_1644,N_14944,N_14741);
nor UO_1645 (O_1645,N_14977,N_14964);
nand UO_1646 (O_1646,N_14910,N_14726);
nand UO_1647 (O_1647,N_14859,N_14830);
xor UO_1648 (O_1648,N_14955,N_14869);
xor UO_1649 (O_1649,N_14730,N_14797);
or UO_1650 (O_1650,N_14992,N_14993);
xnor UO_1651 (O_1651,N_14733,N_14989);
nor UO_1652 (O_1652,N_14735,N_14774);
xor UO_1653 (O_1653,N_14823,N_14931);
or UO_1654 (O_1654,N_14788,N_14787);
or UO_1655 (O_1655,N_14958,N_14815);
or UO_1656 (O_1656,N_14982,N_14873);
and UO_1657 (O_1657,N_14944,N_14719);
nor UO_1658 (O_1658,N_14896,N_14768);
xnor UO_1659 (O_1659,N_14812,N_14880);
nand UO_1660 (O_1660,N_14726,N_14731);
nand UO_1661 (O_1661,N_14773,N_14709);
xor UO_1662 (O_1662,N_14702,N_14899);
nand UO_1663 (O_1663,N_14985,N_14761);
nor UO_1664 (O_1664,N_14762,N_14886);
xor UO_1665 (O_1665,N_14951,N_14704);
and UO_1666 (O_1666,N_14895,N_14716);
nand UO_1667 (O_1667,N_14705,N_14858);
and UO_1668 (O_1668,N_14907,N_14908);
or UO_1669 (O_1669,N_14746,N_14927);
xnor UO_1670 (O_1670,N_14878,N_14710);
and UO_1671 (O_1671,N_14702,N_14713);
xnor UO_1672 (O_1672,N_14708,N_14813);
and UO_1673 (O_1673,N_14885,N_14890);
xor UO_1674 (O_1674,N_14801,N_14810);
and UO_1675 (O_1675,N_14976,N_14972);
nand UO_1676 (O_1676,N_14847,N_14912);
xnor UO_1677 (O_1677,N_14855,N_14844);
or UO_1678 (O_1678,N_14756,N_14997);
or UO_1679 (O_1679,N_14818,N_14842);
nand UO_1680 (O_1680,N_14965,N_14758);
xnor UO_1681 (O_1681,N_14724,N_14995);
xnor UO_1682 (O_1682,N_14723,N_14709);
or UO_1683 (O_1683,N_14857,N_14739);
and UO_1684 (O_1684,N_14993,N_14925);
xnor UO_1685 (O_1685,N_14968,N_14991);
xor UO_1686 (O_1686,N_14733,N_14731);
nor UO_1687 (O_1687,N_14724,N_14988);
nor UO_1688 (O_1688,N_14932,N_14928);
nor UO_1689 (O_1689,N_14714,N_14888);
and UO_1690 (O_1690,N_14915,N_14968);
nand UO_1691 (O_1691,N_14856,N_14977);
xnor UO_1692 (O_1692,N_14859,N_14916);
and UO_1693 (O_1693,N_14767,N_14994);
or UO_1694 (O_1694,N_14859,N_14898);
nand UO_1695 (O_1695,N_14835,N_14967);
and UO_1696 (O_1696,N_14877,N_14926);
or UO_1697 (O_1697,N_14725,N_14722);
or UO_1698 (O_1698,N_14863,N_14832);
nor UO_1699 (O_1699,N_14717,N_14720);
and UO_1700 (O_1700,N_14995,N_14748);
and UO_1701 (O_1701,N_14744,N_14782);
or UO_1702 (O_1702,N_14748,N_14798);
nand UO_1703 (O_1703,N_14880,N_14702);
xor UO_1704 (O_1704,N_14781,N_14862);
xor UO_1705 (O_1705,N_14833,N_14741);
xor UO_1706 (O_1706,N_14725,N_14919);
and UO_1707 (O_1707,N_14923,N_14855);
or UO_1708 (O_1708,N_14944,N_14956);
xnor UO_1709 (O_1709,N_14936,N_14967);
nor UO_1710 (O_1710,N_14742,N_14964);
xnor UO_1711 (O_1711,N_14872,N_14793);
nor UO_1712 (O_1712,N_14959,N_14849);
or UO_1713 (O_1713,N_14820,N_14761);
nor UO_1714 (O_1714,N_14737,N_14944);
xor UO_1715 (O_1715,N_14831,N_14822);
xnor UO_1716 (O_1716,N_14992,N_14831);
or UO_1717 (O_1717,N_14934,N_14891);
nor UO_1718 (O_1718,N_14737,N_14875);
and UO_1719 (O_1719,N_14792,N_14741);
xnor UO_1720 (O_1720,N_14893,N_14791);
nor UO_1721 (O_1721,N_14847,N_14773);
xor UO_1722 (O_1722,N_14708,N_14711);
or UO_1723 (O_1723,N_14858,N_14986);
nor UO_1724 (O_1724,N_14715,N_14848);
or UO_1725 (O_1725,N_14922,N_14997);
or UO_1726 (O_1726,N_14785,N_14726);
xor UO_1727 (O_1727,N_14716,N_14738);
and UO_1728 (O_1728,N_14734,N_14986);
nand UO_1729 (O_1729,N_14929,N_14975);
nand UO_1730 (O_1730,N_14806,N_14809);
or UO_1731 (O_1731,N_14710,N_14854);
and UO_1732 (O_1732,N_14999,N_14998);
nand UO_1733 (O_1733,N_14851,N_14942);
nor UO_1734 (O_1734,N_14721,N_14941);
or UO_1735 (O_1735,N_14910,N_14803);
or UO_1736 (O_1736,N_14788,N_14947);
xor UO_1737 (O_1737,N_14894,N_14817);
and UO_1738 (O_1738,N_14928,N_14887);
nand UO_1739 (O_1739,N_14965,N_14715);
nor UO_1740 (O_1740,N_14955,N_14860);
and UO_1741 (O_1741,N_14752,N_14835);
and UO_1742 (O_1742,N_14879,N_14921);
or UO_1743 (O_1743,N_14834,N_14915);
and UO_1744 (O_1744,N_14948,N_14855);
or UO_1745 (O_1745,N_14783,N_14905);
xor UO_1746 (O_1746,N_14852,N_14724);
nand UO_1747 (O_1747,N_14847,N_14888);
or UO_1748 (O_1748,N_14980,N_14969);
or UO_1749 (O_1749,N_14864,N_14914);
nor UO_1750 (O_1750,N_14925,N_14809);
nor UO_1751 (O_1751,N_14959,N_14833);
and UO_1752 (O_1752,N_14841,N_14821);
nor UO_1753 (O_1753,N_14938,N_14946);
xor UO_1754 (O_1754,N_14811,N_14865);
or UO_1755 (O_1755,N_14934,N_14800);
nor UO_1756 (O_1756,N_14964,N_14883);
nor UO_1757 (O_1757,N_14793,N_14971);
xnor UO_1758 (O_1758,N_14713,N_14985);
xor UO_1759 (O_1759,N_14789,N_14772);
xnor UO_1760 (O_1760,N_14814,N_14820);
nor UO_1761 (O_1761,N_14734,N_14798);
or UO_1762 (O_1762,N_14969,N_14994);
or UO_1763 (O_1763,N_14850,N_14886);
xnor UO_1764 (O_1764,N_14879,N_14872);
and UO_1765 (O_1765,N_14872,N_14713);
nor UO_1766 (O_1766,N_14934,N_14879);
xnor UO_1767 (O_1767,N_14977,N_14862);
or UO_1768 (O_1768,N_14908,N_14814);
nor UO_1769 (O_1769,N_14994,N_14874);
nor UO_1770 (O_1770,N_14927,N_14951);
or UO_1771 (O_1771,N_14890,N_14930);
and UO_1772 (O_1772,N_14986,N_14973);
and UO_1773 (O_1773,N_14974,N_14746);
nand UO_1774 (O_1774,N_14845,N_14905);
nor UO_1775 (O_1775,N_14986,N_14904);
nor UO_1776 (O_1776,N_14841,N_14739);
and UO_1777 (O_1777,N_14920,N_14713);
xor UO_1778 (O_1778,N_14731,N_14855);
or UO_1779 (O_1779,N_14859,N_14753);
nand UO_1780 (O_1780,N_14829,N_14738);
xor UO_1781 (O_1781,N_14837,N_14701);
xor UO_1782 (O_1782,N_14934,N_14790);
or UO_1783 (O_1783,N_14824,N_14890);
and UO_1784 (O_1784,N_14790,N_14754);
nand UO_1785 (O_1785,N_14924,N_14913);
xor UO_1786 (O_1786,N_14934,N_14761);
xor UO_1787 (O_1787,N_14783,N_14860);
nor UO_1788 (O_1788,N_14782,N_14892);
and UO_1789 (O_1789,N_14898,N_14808);
xor UO_1790 (O_1790,N_14918,N_14991);
nor UO_1791 (O_1791,N_14813,N_14714);
or UO_1792 (O_1792,N_14828,N_14771);
and UO_1793 (O_1793,N_14857,N_14939);
xor UO_1794 (O_1794,N_14860,N_14795);
and UO_1795 (O_1795,N_14745,N_14818);
nor UO_1796 (O_1796,N_14778,N_14988);
nand UO_1797 (O_1797,N_14832,N_14799);
and UO_1798 (O_1798,N_14901,N_14992);
and UO_1799 (O_1799,N_14984,N_14805);
nand UO_1800 (O_1800,N_14829,N_14898);
nor UO_1801 (O_1801,N_14808,N_14909);
nand UO_1802 (O_1802,N_14747,N_14884);
nor UO_1803 (O_1803,N_14861,N_14941);
nor UO_1804 (O_1804,N_14893,N_14708);
nor UO_1805 (O_1805,N_14992,N_14828);
or UO_1806 (O_1806,N_14760,N_14784);
or UO_1807 (O_1807,N_14843,N_14880);
nor UO_1808 (O_1808,N_14821,N_14743);
or UO_1809 (O_1809,N_14809,N_14972);
and UO_1810 (O_1810,N_14888,N_14981);
or UO_1811 (O_1811,N_14814,N_14894);
and UO_1812 (O_1812,N_14923,N_14917);
and UO_1813 (O_1813,N_14707,N_14924);
xnor UO_1814 (O_1814,N_14868,N_14827);
nor UO_1815 (O_1815,N_14997,N_14808);
or UO_1816 (O_1816,N_14827,N_14955);
or UO_1817 (O_1817,N_14788,N_14904);
or UO_1818 (O_1818,N_14812,N_14763);
and UO_1819 (O_1819,N_14818,N_14823);
or UO_1820 (O_1820,N_14956,N_14926);
and UO_1821 (O_1821,N_14733,N_14924);
or UO_1822 (O_1822,N_14835,N_14988);
or UO_1823 (O_1823,N_14745,N_14833);
nor UO_1824 (O_1824,N_14974,N_14862);
xnor UO_1825 (O_1825,N_14897,N_14814);
nor UO_1826 (O_1826,N_14903,N_14712);
nand UO_1827 (O_1827,N_14909,N_14929);
and UO_1828 (O_1828,N_14880,N_14782);
and UO_1829 (O_1829,N_14832,N_14700);
nand UO_1830 (O_1830,N_14720,N_14947);
nor UO_1831 (O_1831,N_14760,N_14757);
nand UO_1832 (O_1832,N_14890,N_14859);
nor UO_1833 (O_1833,N_14711,N_14709);
xnor UO_1834 (O_1834,N_14945,N_14924);
and UO_1835 (O_1835,N_14901,N_14815);
or UO_1836 (O_1836,N_14952,N_14836);
or UO_1837 (O_1837,N_14938,N_14828);
xnor UO_1838 (O_1838,N_14761,N_14815);
nand UO_1839 (O_1839,N_14915,N_14930);
xor UO_1840 (O_1840,N_14927,N_14758);
nand UO_1841 (O_1841,N_14812,N_14719);
and UO_1842 (O_1842,N_14889,N_14999);
xnor UO_1843 (O_1843,N_14705,N_14764);
and UO_1844 (O_1844,N_14958,N_14974);
nor UO_1845 (O_1845,N_14791,N_14827);
xnor UO_1846 (O_1846,N_14851,N_14838);
nand UO_1847 (O_1847,N_14816,N_14924);
xnor UO_1848 (O_1848,N_14956,N_14774);
and UO_1849 (O_1849,N_14868,N_14848);
and UO_1850 (O_1850,N_14765,N_14979);
and UO_1851 (O_1851,N_14792,N_14995);
and UO_1852 (O_1852,N_14957,N_14779);
nor UO_1853 (O_1853,N_14931,N_14788);
xor UO_1854 (O_1854,N_14807,N_14811);
nor UO_1855 (O_1855,N_14900,N_14912);
nor UO_1856 (O_1856,N_14750,N_14740);
and UO_1857 (O_1857,N_14801,N_14849);
or UO_1858 (O_1858,N_14758,N_14861);
or UO_1859 (O_1859,N_14802,N_14911);
nand UO_1860 (O_1860,N_14804,N_14943);
or UO_1861 (O_1861,N_14802,N_14748);
xor UO_1862 (O_1862,N_14709,N_14737);
nor UO_1863 (O_1863,N_14909,N_14840);
nor UO_1864 (O_1864,N_14972,N_14926);
or UO_1865 (O_1865,N_14930,N_14779);
or UO_1866 (O_1866,N_14877,N_14712);
and UO_1867 (O_1867,N_14751,N_14745);
xnor UO_1868 (O_1868,N_14968,N_14952);
nand UO_1869 (O_1869,N_14865,N_14728);
or UO_1870 (O_1870,N_14702,N_14871);
and UO_1871 (O_1871,N_14988,N_14714);
xor UO_1872 (O_1872,N_14855,N_14930);
nand UO_1873 (O_1873,N_14844,N_14835);
xor UO_1874 (O_1874,N_14782,N_14760);
nor UO_1875 (O_1875,N_14808,N_14777);
nor UO_1876 (O_1876,N_14861,N_14896);
nor UO_1877 (O_1877,N_14768,N_14865);
and UO_1878 (O_1878,N_14759,N_14801);
nand UO_1879 (O_1879,N_14992,N_14709);
xor UO_1880 (O_1880,N_14762,N_14758);
nor UO_1881 (O_1881,N_14877,N_14732);
nor UO_1882 (O_1882,N_14923,N_14763);
nand UO_1883 (O_1883,N_14814,N_14903);
or UO_1884 (O_1884,N_14888,N_14700);
or UO_1885 (O_1885,N_14701,N_14857);
nor UO_1886 (O_1886,N_14958,N_14789);
nand UO_1887 (O_1887,N_14972,N_14850);
nor UO_1888 (O_1888,N_14769,N_14878);
or UO_1889 (O_1889,N_14773,N_14749);
nor UO_1890 (O_1890,N_14760,N_14917);
nand UO_1891 (O_1891,N_14746,N_14782);
or UO_1892 (O_1892,N_14740,N_14809);
and UO_1893 (O_1893,N_14833,N_14771);
xor UO_1894 (O_1894,N_14916,N_14700);
xor UO_1895 (O_1895,N_14793,N_14881);
nand UO_1896 (O_1896,N_14988,N_14809);
or UO_1897 (O_1897,N_14712,N_14909);
xnor UO_1898 (O_1898,N_14773,N_14842);
or UO_1899 (O_1899,N_14719,N_14854);
nor UO_1900 (O_1900,N_14832,N_14899);
or UO_1901 (O_1901,N_14995,N_14742);
nand UO_1902 (O_1902,N_14990,N_14876);
nor UO_1903 (O_1903,N_14737,N_14965);
nand UO_1904 (O_1904,N_14872,N_14740);
nor UO_1905 (O_1905,N_14984,N_14828);
and UO_1906 (O_1906,N_14817,N_14965);
nand UO_1907 (O_1907,N_14827,N_14779);
nand UO_1908 (O_1908,N_14791,N_14799);
or UO_1909 (O_1909,N_14926,N_14976);
nand UO_1910 (O_1910,N_14866,N_14771);
nor UO_1911 (O_1911,N_14885,N_14865);
or UO_1912 (O_1912,N_14991,N_14944);
xnor UO_1913 (O_1913,N_14789,N_14743);
nor UO_1914 (O_1914,N_14863,N_14721);
nor UO_1915 (O_1915,N_14922,N_14968);
nand UO_1916 (O_1916,N_14727,N_14894);
and UO_1917 (O_1917,N_14833,N_14811);
or UO_1918 (O_1918,N_14969,N_14716);
and UO_1919 (O_1919,N_14759,N_14958);
nor UO_1920 (O_1920,N_14967,N_14937);
or UO_1921 (O_1921,N_14916,N_14755);
or UO_1922 (O_1922,N_14812,N_14905);
nand UO_1923 (O_1923,N_14854,N_14720);
xnor UO_1924 (O_1924,N_14974,N_14703);
nand UO_1925 (O_1925,N_14704,N_14757);
nor UO_1926 (O_1926,N_14815,N_14781);
nor UO_1927 (O_1927,N_14990,N_14739);
or UO_1928 (O_1928,N_14819,N_14823);
and UO_1929 (O_1929,N_14933,N_14985);
xnor UO_1930 (O_1930,N_14898,N_14831);
and UO_1931 (O_1931,N_14912,N_14725);
nor UO_1932 (O_1932,N_14807,N_14965);
xor UO_1933 (O_1933,N_14731,N_14827);
nand UO_1934 (O_1934,N_14895,N_14809);
nand UO_1935 (O_1935,N_14808,N_14975);
nor UO_1936 (O_1936,N_14720,N_14758);
nor UO_1937 (O_1937,N_14945,N_14982);
xnor UO_1938 (O_1938,N_14815,N_14711);
nor UO_1939 (O_1939,N_14730,N_14747);
nand UO_1940 (O_1940,N_14736,N_14818);
nand UO_1941 (O_1941,N_14773,N_14967);
nand UO_1942 (O_1942,N_14947,N_14881);
and UO_1943 (O_1943,N_14788,N_14791);
nand UO_1944 (O_1944,N_14740,N_14831);
nor UO_1945 (O_1945,N_14895,N_14897);
or UO_1946 (O_1946,N_14895,N_14903);
and UO_1947 (O_1947,N_14829,N_14703);
nand UO_1948 (O_1948,N_14985,N_14768);
xnor UO_1949 (O_1949,N_14843,N_14762);
nor UO_1950 (O_1950,N_14814,N_14815);
or UO_1951 (O_1951,N_14760,N_14742);
or UO_1952 (O_1952,N_14939,N_14826);
and UO_1953 (O_1953,N_14871,N_14905);
or UO_1954 (O_1954,N_14944,N_14829);
or UO_1955 (O_1955,N_14783,N_14891);
and UO_1956 (O_1956,N_14957,N_14792);
nor UO_1957 (O_1957,N_14948,N_14982);
nor UO_1958 (O_1958,N_14935,N_14904);
nor UO_1959 (O_1959,N_14921,N_14873);
and UO_1960 (O_1960,N_14727,N_14848);
or UO_1961 (O_1961,N_14969,N_14761);
xnor UO_1962 (O_1962,N_14994,N_14830);
and UO_1963 (O_1963,N_14996,N_14862);
nand UO_1964 (O_1964,N_14759,N_14803);
nor UO_1965 (O_1965,N_14857,N_14805);
or UO_1966 (O_1966,N_14855,N_14804);
nor UO_1967 (O_1967,N_14717,N_14850);
and UO_1968 (O_1968,N_14892,N_14705);
xnor UO_1969 (O_1969,N_14775,N_14807);
and UO_1970 (O_1970,N_14800,N_14945);
nor UO_1971 (O_1971,N_14946,N_14707);
nor UO_1972 (O_1972,N_14983,N_14789);
nor UO_1973 (O_1973,N_14951,N_14737);
nand UO_1974 (O_1974,N_14832,N_14813);
and UO_1975 (O_1975,N_14763,N_14859);
xnor UO_1976 (O_1976,N_14965,N_14956);
and UO_1977 (O_1977,N_14918,N_14722);
and UO_1978 (O_1978,N_14964,N_14745);
and UO_1979 (O_1979,N_14784,N_14987);
or UO_1980 (O_1980,N_14725,N_14724);
or UO_1981 (O_1981,N_14975,N_14917);
nor UO_1982 (O_1982,N_14897,N_14818);
or UO_1983 (O_1983,N_14874,N_14749);
xnor UO_1984 (O_1984,N_14747,N_14755);
xnor UO_1985 (O_1985,N_14719,N_14929);
and UO_1986 (O_1986,N_14848,N_14873);
and UO_1987 (O_1987,N_14760,N_14842);
nor UO_1988 (O_1988,N_14939,N_14747);
xor UO_1989 (O_1989,N_14989,N_14707);
nor UO_1990 (O_1990,N_14863,N_14917);
xor UO_1991 (O_1991,N_14836,N_14820);
and UO_1992 (O_1992,N_14766,N_14808);
or UO_1993 (O_1993,N_14948,N_14824);
nand UO_1994 (O_1994,N_14862,N_14716);
or UO_1995 (O_1995,N_14921,N_14744);
and UO_1996 (O_1996,N_14711,N_14778);
xor UO_1997 (O_1997,N_14929,N_14707);
nand UO_1998 (O_1998,N_14925,N_14928);
and UO_1999 (O_1999,N_14789,N_14981);
endmodule