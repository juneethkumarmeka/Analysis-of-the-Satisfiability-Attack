module basic_2500_25000_3000_8_levels_5xor_1(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,In_750,In_751,In_752,In_753,In_754,In_755,In_756,In_757,In_758,In_759,In_760,In_761,In_762,In_763,In_764,In_765,In_766,In_767,In_768,In_769,In_770,In_771,In_772,In_773,In_774,In_775,In_776,In_777,In_778,In_779,In_780,In_781,In_782,In_783,In_784,In_785,In_786,In_787,In_788,In_789,In_790,In_791,In_792,In_793,In_794,In_795,In_796,In_797,In_798,In_799,In_800,In_801,In_802,In_803,In_804,In_805,In_806,In_807,In_808,In_809,In_810,In_811,In_812,In_813,In_814,In_815,In_816,In_817,In_818,In_819,In_820,In_821,In_822,In_823,In_824,In_825,In_826,In_827,In_828,In_829,In_830,In_831,In_832,In_833,In_834,In_835,In_836,In_837,In_838,In_839,In_840,In_841,In_842,In_843,In_844,In_845,In_846,In_847,In_848,In_849,In_850,In_851,In_852,In_853,In_854,In_855,In_856,In_857,In_858,In_859,In_860,In_861,In_862,In_863,In_864,In_865,In_866,In_867,In_868,In_869,In_870,In_871,In_872,In_873,In_874,In_875,In_876,In_877,In_878,In_879,In_880,In_881,In_882,In_883,In_884,In_885,In_886,In_887,In_888,In_889,In_890,In_891,In_892,In_893,In_894,In_895,In_896,In_897,In_898,In_899,In_900,In_901,In_902,In_903,In_904,In_905,In_906,In_907,In_908,In_909,In_910,In_911,In_912,In_913,In_914,In_915,In_916,In_917,In_918,In_919,In_920,In_921,In_922,In_923,In_924,In_925,In_926,In_927,In_928,In_929,In_930,In_931,In_932,In_933,In_934,In_935,In_936,In_937,In_938,In_939,In_940,In_941,In_942,In_943,In_944,In_945,In_946,In_947,In_948,In_949,In_950,In_951,In_952,In_953,In_954,In_955,In_956,In_957,In_958,In_959,In_960,In_961,In_962,In_963,In_964,In_965,In_966,In_967,In_968,In_969,In_970,In_971,In_972,In_973,In_974,In_975,In_976,In_977,In_978,In_979,In_980,In_981,In_982,In_983,In_984,In_985,In_986,In_987,In_988,In_989,In_990,In_991,In_992,In_993,In_994,In_995,In_996,In_997,In_998,In_999,In_1000,In_1001,In_1002,In_1003,In_1004,In_1005,In_1006,In_1007,In_1008,In_1009,In_1010,In_1011,In_1012,In_1013,In_1014,In_1015,In_1016,In_1017,In_1018,In_1019,In_1020,In_1021,In_1022,In_1023,In_1024,In_1025,In_1026,In_1027,In_1028,In_1029,In_1030,In_1031,In_1032,In_1033,In_1034,In_1035,In_1036,In_1037,In_1038,In_1039,In_1040,In_1041,In_1042,In_1043,In_1044,In_1045,In_1046,In_1047,In_1048,In_1049,In_1050,In_1051,In_1052,In_1053,In_1054,In_1055,In_1056,In_1057,In_1058,In_1059,In_1060,In_1061,In_1062,In_1063,In_1064,In_1065,In_1066,In_1067,In_1068,In_1069,In_1070,In_1071,In_1072,In_1073,In_1074,In_1075,In_1076,In_1077,In_1078,In_1079,In_1080,In_1081,In_1082,In_1083,In_1084,In_1085,In_1086,In_1087,In_1088,In_1089,In_1090,In_1091,In_1092,In_1093,In_1094,In_1095,In_1096,In_1097,In_1098,In_1099,In_1100,In_1101,In_1102,In_1103,In_1104,In_1105,In_1106,In_1107,In_1108,In_1109,In_1110,In_1111,In_1112,In_1113,In_1114,In_1115,In_1116,In_1117,In_1118,In_1119,In_1120,In_1121,In_1122,In_1123,In_1124,In_1125,In_1126,In_1127,In_1128,In_1129,In_1130,In_1131,In_1132,In_1133,In_1134,In_1135,In_1136,In_1137,In_1138,In_1139,In_1140,In_1141,In_1142,In_1143,In_1144,In_1145,In_1146,In_1147,In_1148,In_1149,In_1150,In_1151,In_1152,In_1153,In_1154,In_1155,In_1156,In_1157,In_1158,In_1159,In_1160,In_1161,In_1162,In_1163,In_1164,In_1165,In_1166,In_1167,In_1168,In_1169,In_1170,In_1171,In_1172,In_1173,In_1174,In_1175,In_1176,In_1177,In_1178,In_1179,In_1180,In_1181,In_1182,In_1183,In_1184,In_1185,In_1186,In_1187,In_1188,In_1189,In_1190,In_1191,In_1192,In_1193,In_1194,In_1195,In_1196,In_1197,In_1198,In_1199,In_1200,In_1201,In_1202,In_1203,In_1204,In_1205,In_1206,In_1207,In_1208,In_1209,In_1210,In_1211,In_1212,In_1213,In_1214,In_1215,In_1216,In_1217,In_1218,In_1219,In_1220,In_1221,In_1222,In_1223,In_1224,In_1225,In_1226,In_1227,In_1228,In_1229,In_1230,In_1231,In_1232,In_1233,In_1234,In_1235,In_1236,In_1237,In_1238,In_1239,In_1240,In_1241,In_1242,In_1243,In_1244,In_1245,In_1246,In_1247,In_1248,In_1249,In_1250,In_1251,In_1252,In_1253,In_1254,In_1255,In_1256,In_1257,In_1258,In_1259,In_1260,In_1261,In_1262,In_1263,In_1264,In_1265,In_1266,In_1267,In_1268,In_1269,In_1270,In_1271,In_1272,In_1273,In_1274,In_1275,In_1276,In_1277,In_1278,In_1279,In_1280,In_1281,In_1282,In_1283,In_1284,In_1285,In_1286,In_1287,In_1288,In_1289,In_1290,In_1291,In_1292,In_1293,In_1294,In_1295,In_1296,In_1297,In_1298,In_1299,In_1300,In_1301,In_1302,In_1303,In_1304,In_1305,In_1306,In_1307,In_1308,In_1309,In_1310,In_1311,In_1312,In_1313,In_1314,In_1315,In_1316,In_1317,In_1318,In_1319,In_1320,In_1321,In_1322,In_1323,In_1324,In_1325,In_1326,In_1327,In_1328,In_1329,In_1330,In_1331,In_1332,In_1333,In_1334,In_1335,In_1336,In_1337,In_1338,In_1339,In_1340,In_1341,In_1342,In_1343,In_1344,In_1345,In_1346,In_1347,In_1348,In_1349,In_1350,In_1351,In_1352,In_1353,In_1354,In_1355,In_1356,In_1357,In_1358,In_1359,In_1360,In_1361,In_1362,In_1363,In_1364,In_1365,In_1366,In_1367,In_1368,In_1369,In_1370,In_1371,In_1372,In_1373,In_1374,In_1375,In_1376,In_1377,In_1378,In_1379,In_1380,In_1381,In_1382,In_1383,In_1384,In_1385,In_1386,In_1387,In_1388,In_1389,In_1390,In_1391,In_1392,In_1393,In_1394,In_1395,In_1396,In_1397,In_1398,In_1399,In_1400,In_1401,In_1402,In_1403,In_1404,In_1405,In_1406,In_1407,In_1408,In_1409,In_1410,In_1411,In_1412,In_1413,In_1414,In_1415,In_1416,In_1417,In_1418,In_1419,In_1420,In_1421,In_1422,In_1423,In_1424,In_1425,In_1426,In_1427,In_1428,In_1429,In_1430,In_1431,In_1432,In_1433,In_1434,In_1435,In_1436,In_1437,In_1438,In_1439,In_1440,In_1441,In_1442,In_1443,In_1444,In_1445,In_1446,In_1447,In_1448,In_1449,In_1450,In_1451,In_1452,In_1453,In_1454,In_1455,In_1456,In_1457,In_1458,In_1459,In_1460,In_1461,In_1462,In_1463,In_1464,In_1465,In_1466,In_1467,In_1468,In_1469,In_1470,In_1471,In_1472,In_1473,In_1474,In_1475,In_1476,In_1477,In_1478,In_1479,In_1480,In_1481,In_1482,In_1483,In_1484,In_1485,In_1486,In_1487,In_1488,In_1489,In_1490,In_1491,In_1492,In_1493,In_1494,In_1495,In_1496,In_1497,In_1498,In_1499,In_1500,In_1501,In_1502,In_1503,In_1504,In_1505,In_1506,In_1507,In_1508,In_1509,In_1510,In_1511,In_1512,In_1513,In_1514,In_1515,In_1516,In_1517,In_1518,In_1519,In_1520,In_1521,In_1522,In_1523,In_1524,In_1525,In_1526,In_1527,In_1528,In_1529,In_1530,In_1531,In_1532,In_1533,In_1534,In_1535,In_1536,In_1537,In_1538,In_1539,In_1540,In_1541,In_1542,In_1543,In_1544,In_1545,In_1546,In_1547,In_1548,In_1549,In_1550,In_1551,In_1552,In_1553,In_1554,In_1555,In_1556,In_1557,In_1558,In_1559,In_1560,In_1561,In_1562,In_1563,In_1564,In_1565,In_1566,In_1567,In_1568,In_1569,In_1570,In_1571,In_1572,In_1573,In_1574,In_1575,In_1576,In_1577,In_1578,In_1579,In_1580,In_1581,In_1582,In_1583,In_1584,In_1585,In_1586,In_1587,In_1588,In_1589,In_1590,In_1591,In_1592,In_1593,In_1594,In_1595,In_1596,In_1597,In_1598,In_1599,In_1600,In_1601,In_1602,In_1603,In_1604,In_1605,In_1606,In_1607,In_1608,In_1609,In_1610,In_1611,In_1612,In_1613,In_1614,In_1615,In_1616,In_1617,In_1618,In_1619,In_1620,In_1621,In_1622,In_1623,In_1624,In_1625,In_1626,In_1627,In_1628,In_1629,In_1630,In_1631,In_1632,In_1633,In_1634,In_1635,In_1636,In_1637,In_1638,In_1639,In_1640,In_1641,In_1642,In_1643,In_1644,In_1645,In_1646,In_1647,In_1648,In_1649,In_1650,In_1651,In_1652,In_1653,In_1654,In_1655,In_1656,In_1657,In_1658,In_1659,In_1660,In_1661,In_1662,In_1663,In_1664,In_1665,In_1666,In_1667,In_1668,In_1669,In_1670,In_1671,In_1672,In_1673,In_1674,In_1675,In_1676,In_1677,In_1678,In_1679,In_1680,In_1681,In_1682,In_1683,In_1684,In_1685,In_1686,In_1687,In_1688,In_1689,In_1690,In_1691,In_1692,In_1693,In_1694,In_1695,In_1696,In_1697,In_1698,In_1699,In_1700,In_1701,In_1702,In_1703,In_1704,In_1705,In_1706,In_1707,In_1708,In_1709,In_1710,In_1711,In_1712,In_1713,In_1714,In_1715,In_1716,In_1717,In_1718,In_1719,In_1720,In_1721,In_1722,In_1723,In_1724,In_1725,In_1726,In_1727,In_1728,In_1729,In_1730,In_1731,In_1732,In_1733,In_1734,In_1735,In_1736,In_1737,In_1738,In_1739,In_1740,In_1741,In_1742,In_1743,In_1744,In_1745,In_1746,In_1747,In_1748,In_1749,In_1750,In_1751,In_1752,In_1753,In_1754,In_1755,In_1756,In_1757,In_1758,In_1759,In_1760,In_1761,In_1762,In_1763,In_1764,In_1765,In_1766,In_1767,In_1768,In_1769,In_1770,In_1771,In_1772,In_1773,In_1774,In_1775,In_1776,In_1777,In_1778,In_1779,In_1780,In_1781,In_1782,In_1783,In_1784,In_1785,In_1786,In_1787,In_1788,In_1789,In_1790,In_1791,In_1792,In_1793,In_1794,In_1795,In_1796,In_1797,In_1798,In_1799,In_1800,In_1801,In_1802,In_1803,In_1804,In_1805,In_1806,In_1807,In_1808,In_1809,In_1810,In_1811,In_1812,In_1813,In_1814,In_1815,In_1816,In_1817,In_1818,In_1819,In_1820,In_1821,In_1822,In_1823,In_1824,In_1825,In_1826,In_1827,In_1828,In_1829,In_1830,In_1831,In_1832,In_1833,In_1834,In_1835,In_1836,In_1837,In_1838,In_1839,In_1840,In_1841,In_1842,In_1843,In_1844,In_1845,In_1846,In_1847,In_1848,In_1849,In_1850,In_1851,In_1852,In_1853,In_1854,In_1855,In_1856,In_1857,In_1858,In_1859,In_1860,In_1861,In_1862,In_1863,In_1864,In_1865,In_1866,In_1867,In_1868,In_1869,In_1870,In_1871,In_1872,In_1873,In_1874,In_1875,In_1876,In_1877,In_1878,In_1879,In_1880,In_1881,In_1882,In_1883,In_1884,In_1885,In_1886,In_1887,In_1888,In_1889,In_1890,In_1891,In_1892,In_1893,In_1894,In_1895,In_1896,In_1897,In_1898,In_1899,In_1900,In_1901,In_1902,In_1903,In_1904,In_1905,In_1906,In_1907,In_1908,In_1909,In_1910,In_1911,In_1912,In_1913,In_1914,In_1915,In_1916,In_1917,In_1918,In_1919,In_1920,In_1921,In_1922,In_1923,In_1924,In_1925,In_1926,In_1927,In_1928,In_1929,In_1930,In_1931,In_1932,In_1933,In_1934,In_1935,In_1936,In_1937,In_1938,In_1939,In_1940,In_1941,In_1942,In_1943,In_1944,In_1945,In_1946,In_1947,In_1948,In_1949,In_1950,In_1951,In_1952,In_1953,In_1954,In_1955,In_1956,In_1957,In_1958,In_1959,In_1960,In_1961,In_1962,In_1963,In_1964,In_1965,In_1966,In_1967,In_1968,In_1969,In_1970,In_1971,In_1972,In_1973,In_1974,In_1975,In_1976,In_1977,In_1978,In_1979,In_1980,In_1981,In_1982,In_1983,In_1984,In_1985,In_1986,In_1987,In_1988,In_1989,In_1990,In_1991,In_1992,In_1993,In_1994,In_1995,In_1996,In_1997,In_1998,In_1999,In_2000,In_2001,In_2002,In_2003,In_2004,In_2005,In_2006,In_2007,In_2008,In_2009,In_2010,In_2011,In_2012,In_2013,In_2014,In_2015,In_2016,In_2017,In_2018,In_2019,In_2020,In_2021,In_2022,In_2023,In_2024,In_2025,In_2026,In_2027,In_2028,In_2029,In_2030,In_2031,In_2032,In_2033,In_2034,In_2035,In_2036,In_2037,In_2038,In_2039,In_2040,In_2041,In_2042,In_2043,In_2044,In_2045,In_2046,In_2047,In_2048,In_2049,In_2050,In_2051,In_2052,In_2053,In_2054,In_2055,In_2056,In_2057,In_2058,In_2059,In_2060,In_2061,In_2062,In_2063,In_2064,In_2065,In_2066,In_2067,In_2068,In_2069,In_2070,In_2071,In_2072,In_2073,In_2074,In_2075,In_2076,In_2077,In_2078,In_2079,In_2080,In_2081,In_2082,In_2083,In_2084,In_2085,In_2086,In_2087,In_2088,In_2089,In_2090,In_2091,In_2092,In_2093,In_2094,In_2095,In_2096,In_2097,In_2098,In_2099,In_2100,In_2101,In_2102,In_2103,In_2104,In_2105,In_2106,In_2107,In_2108,In_2109,In_2110,In_2111,In_2112,In_2113,In_2114,In_2115,In_2116,In_2117,In_2118,In_2119,In_2120,In_2121,In_2122,In_2123,In_2124,In_2125,In_2126,In_2127,In_2128,In_2129,In_2130,In_2131,In_2132,In_2133,In_2134,In_2135,In_2136,In_2137,In_2138,In_2139,In_2140,In_2141,In_2142,In_2143,In_2144,In_2145,In_2146,In_2147,In_2148,In_2149,In_2150,In_2151,In_2152,In_2153,In_2154,In_2155,In_2156,In_2157,In_2158,In_2159,In_2160,In_2161,In_2162,In_2163,In_2164,In_2165,In_2166,In_2167,In_2168,In_2169,In_2170,In_2171,In_2172,In_2173,In_2174,In_2175,In_2176,In_2177,In_2178,In_2179,In_2180,In_2181,In_2182,In_2183,In_2184,In_2185,In_2186,In_2187,In_2188,In_2189,In_2190,In_2191,In_2192,In_2193,In_2194,In_2195,In_2196,In_2197,In_2198,In_2199,In_2200,In_2201,In_2202,In_2203,In_2204,In_2205,In_2206,In_2207,In_2208,In_2209,In_2210,In_2211,In_2212,In_2213,In_2214,In_2215,In_2216,In_2217,In_2218,In_2219,In_2220,In_2221,In_2222,In_2223,In_2224,In_2225,In_2226,In_2227,In_2228,In_2229,In_2230,In_2231,In_2232,In_2233,In_2234,In_2235,In_2236,In_2237,In_2238,In_2239,In_2240,In_2241,In_2242,In_2243,In_2244,In_2245,In_2246,In_2247,In_2248,In_2249,In_2250,In_2251,In_2252,In_2253,In_2254,In_2255,In_2256,In_2257,In_2258,In_2259,In_2260,In_2261,In_2262,In_2263,In_2264,In_2265,In_2266,In_2267,In_2268,In_2269,In_2270,In_2271,In_2272,In_2273,In_2274,In_2275,In_2276,In_2277,In_2278,In_2279,In_2280,In_2281,In_2282,In_2283,In_2284,In_2285,In_2286,In_2287,In_2288,In_2289,In_2290,In_2291,In_2292,In_2293,In_2294,In_2295,In_2296,In_2297,In_2298,In_2299,In_2300,In_2301,In_2302,In_2303,In_2304,In_2305,In_2306,In_2307,In_2308,In_2309,In_2310,In_2311,In_2312,In_2313,In_2314,In_2315,In_2316,In_2317,In_2318,In_2319,In_2320,In_2321,In_2322,In_2323,In_2324,In_2325,In_2326,In_2327,In_2328,In_2329,In_2330,In_2331,In_2332,In_2333,In_2334,In_2335,In_2336,In_2337,In_2338,In_2339,In_2340,In_2341,In_2342,In_2343,In_2344,In_2345,In_2346,In_2347,In_2348,In_2349,In_2350,In_2351,In_2352,In_2353,In_2354,In_2355,In_2356,In_2357,In_2358,In_2359,In_2360,In_2361,In_2362,In_2363,In_2364,In_2365,In_2366,In_2367,In_2368,In_2369,In_2370,In_2371,In_2372,In_2373,In_2374,In_2375,In_2376,In_2377,In_2378,In_2379,In_2380,In_2381,In_2382,In_2383,In_2384,In_2385,In_2386,In_2387,In_2388,In_2389,In_2390,In_2391,In_2392,In_2393,In_2394,In_2395,In_2396,In_2397,In_2398,In_2399,In_2400,In_2401,In_2402,In_2403,In_2404,In_2405,In_2406,In_2407,In_2408,In_2409,In_2410,In_2411,In_2412,In_2413,In_2414,In_2415,In_2416,In_2417,In_2418,In_2419,In_2420,In_2421,In_2422,In_2423,In_2424,In_2425,In_2426,In_2427,In_2428,In_2429,In_2430,In_2431,In_2432,In_2433,In_2434,In_2435,In_2436,In_2437,In_2438,In_2439,In_2440,In_2441,In_2442,In_2443,In_2444,In_2445,In_2446,In_2447,In_2448,In_2449,In_2450,In_2451,In_2452,In_2453,In_2454,In_2455,In_2456,In_2457,In_2458,In_2459,In_2460,In_2461,In_2462,In_2463,In_2464,In_2465,In_2466,In_2467,In_2468,In_2469,In_2470,In_2471,In_2472,In_2473,In_2474,In_2475,In_2476,In_2477,In_2478,In_2479,In_2480,In_2481,In_2482,In_2483,In_2484,In_2485,In_2486,In_2487,In_2488,In_2489,In_2490,In_2491,In_2492,In_2493,In_2494,In_2495,In_2496,In_2497,In_2498,In_2499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999,O_1000,O_1001,O_1002,O_1003,O_1004,O_1005,O_1006,O_1007,O_1008,O_1009,O_1010,O_1011,O_1012,O_1013,O_1014,O_1015,O_1016,O_1017,O_1018,O_1019,O_1020,O_1021,O_1022,O_1023,O_1024,O_1025,O_1026,O_1027,O_1028,O_1029,O_1030,O_1031,O_1032,O_1033,O_1034,O_1035,O_1036,O_1037,O_1038,O_1039,O_1040,O_1041,O_1042,O_1043,O_1044,O_1045,O_1046,O_1047,O_1048,O_1049,O_1050,O_1051,O_1052,O_1053,O_1054,O_1055,O_1056,O_1057,O_1058,O_1059,O_1060,O_1061,O_1062,O_1063,O_1064,O_1065,O_1066,O_1067,O_1068,O_1069,O_1070,O_1071,O_1072,O_1073,O_1074,O_1075,O_1076,O_1077,O_1078,O_1079,O_1080,O_1081,O_1082,O_1083,O_1084,O_1085,O_1086,O_1087,O_1088,O_1089,O_1090,O_1091,O_1092,O_1093,O_1094,O_1095,O_1096,O_1097,O_1098,O_1099,O_1100,O_1101,O_1102,O_1103,O_1104,O_1105,O_1106,O_1107,O_1108,O_1109,O_1110,O_1111,O_1112,O_1113,O_1114,O_1115,O_1116,O_1117,O_1118,O_1119,O_1120,O_1121,O_1122,O_1123,O_1124,O_1125,O_1126,O_1127,O_1128,O_1129,O_1130,O_1131,O_1132,O_1133,O_1134,O_1135,O_1136,O_1137,O_1138,O_1139,O_1140,O_1141,O_1142,O_1143,O_1144,O_1145,O_1146,O_1147,O_1148,O_1149,O_1150,O_1151,O_1152,O_1153,O_1154,O_1155,O_1156,O_1157,O_1158,O_1159,O_1160,O_1161,O_1162,O_1163,O_1164,O_1165,O_1166,O_1167,O_1168,O_1169,O_1170,O_1171,O_1172,O_1173,O_1174,O_1175,O_1176,O_1177,O_1178,O_1179,O_1180,O_1181,O_1182,O_1183,O_1184,O_1185,O_1186,O_1187,O_1188,O_1189,O_1190,O_1191,O_1192,O_1193,O_1194,O_1195,O_1196,O_1197,O_1198,O_1199,O_1200,O_1201,O_1202,O_1203,O_1204,O_1205,O_1206,O_1207,O_1208,O_1209,O_1210,O_1211,O_1212,O_1213,O_1214,O_1215,O_1216,O_1217,O_1218,O_1219,O_1220,O_1221,O_1222,O_1223,O_1224,O_1225,O_1226,O_1227,O_1228,O_1229,O_1230,O_1231,O_1232,O_1233,O_1234,O_1235,O_1236,O_1237,O_1238,O_1239,O_1240,O_1241,O_1242,O_1243,O_1244,O_1245,O_1246,O_1247,O_1248,O_1249,O_1250,O_1251,O_1252,O_1253,O_1254,O_1255,O_1256,O_1257,O_1258,O_1259,O_1260,O_1261,O_1262,O_1263,O_1264,O_1265,O_1266,O_1267,O_1268,O_1269,O_1270,O_1271,O_1272,O_1273,O_1274,O_1275,O_1276,O_1277,O_1278,O_1279,O_1280,O_1281,O_1282,O_1283,O_1284,O_1285,O_1286,O_1287,O_1288,O_1289,O_1290,O_1291,O_1292,O_1293,O_1294,O_1295,O_1296,O_1297,O_1298,O_1299,O_1300,O_1301,O_1302,O_1303,O_1304,O_1305,O_1306,O_1307,O_1308,O_1309,O_1310,O_1311,O_1312,O_1313,O_1314,O_1315,O_1316,O_1317,O_1318,O_1319,O_1320,O_1321,O_1322,O_1323,O_1324,O_1325,O_1326,O_1327,O_1328,O_1329,O_1330,O_1331,O_1332,O_1333,O_1334,O_1335,O_1336,O_1337,O_1338,O_1339,O_1340,O_1341,O_1342,O_1343,O_1344,O_1345,O_1346,O_1347,O_1348,O_1349,O_1350,O_1351,O_1352,O_1353,O_1354,O_1355,O_1356,O_1357,O_1358,O_1359,O_1360,O_1361,O_1362,O_1363,O_1364,O_1365,O_1366,O_1367,O_1368,O_1369,O_1370,O_1371,O_1372,O_1373,O_1374,O_1375,O_1376,O_1377,O_1378,O_1379,O_1380,O_1381,O_1382,O_1383,O_1384,O_1385,O_1386,O_1387,O_1388,O_1389,O_1390,O_1391,O_1392,O_1393,O_1394,O_1395,O_1396,O_1397,O_1398,O_1399,O_1400,O_1401,O_1402,O_1403,O_1404,O_1405,O_1406,O_1407,O_1408,O_1409,O_1410,O_1411,O_1412,O_1413,O_1414,O_1415,O_1416,O_1417,O_1418,O_1419,O_1420,O_1421,O_1422,O_1423,O_1424,O_1425,O_1426,O_1427,O_1428,O_1429,O_1430,O_1431,O_1432,O_1433,O_1434,O_1435,O_1436,O_1437,O_1438,O_1439,O_1440,O_1441,O_1442,O_1443,O_1444,O_1445,O_1446,O_1447,O_1448,O_1449,O_1450,O_1451,O_1452,O_1453,O_1454,O_1455,O_1456,O_1457,O_1458,O_1459,O_1460,O_1461,O_1462,O_1463,O_1464,O_1465,O_1466,O_1467,O_1468,O_1469,O_1470,O_1471,O_1472,O_1473,O_1474,O_1475,O_1476,O_1477,O_1478,O_1479,O_1480,O_1481,O_1482,O_1483,O_1484,O_1485,O_1486,O_1487,O_1488,O_1489,O_1490,O_1491,O_1492,O_1493,O_1494,O_1495,O_1496,O_1497,O_1498,O_1499,O_1500,O_1501,O_1502,O_1503,O_1504,O_1505,O_1506,O_1507,O_1508,O_1509,O_1510,O_1511,O_1512,O_1513,O_1514,O_1515,O_1516,O_1517,O_1518,O_1519,O_1520,O_1521,O_1522,O_1523,O_1524,O_1525,O_1526,O_1527,O_1528,O_1529,O_1530,O_1531,O_1532,O_1533,O_1534,O_1535,O_1536,O_1537,O_1538,O_1539,O_1540,O_1541,O_1542,O_1543,O_1544,O_1545,O_1546,O_1547,O_1548,O_1549,O_1550,O_1551,O_1552,O_1553,O_1554,O_1555,O_1556,O_1557,O_1558,O_1559,O_1560,O_1561,O_1562,O_1563,O_1564,O_1565,O_1566,O_1567,O_1568,O_1569,O_1570,O_1571,O_1572,O_1573,O_1574,O_1575,O_1576,O_1577,O_1578,O_1579,O_1580,O_1581,O_1582,O_1583,O_1584,O_1585,O_1586,O_1587,O_1588,O_1589,O_1590,O_1591,O_1592,O_1593,O_1594,O_1595,O_1596,O_1597,O_1598,O_1599,O_1600,O_1601,O_1602,O_1603,O_1604,O_1605,O_1606,O_1607,O_1608,O_1609,O_1610,O_1611,O_1612,O_1613,O_1614,O_1615,O_1616,O_1617,O_1618,O_1619,O_1620,O_1621,O_1622,O_1623,O_1624,O_1625,O_1626,O_1627,O_1628,O_1629,O_1630,O_1631,O_1632,O_1633,O_1634,O_1635,O_1636,O_1637,O_1638,O_1639,O_1640,O_1641,O_1642,O_1643,O_1644,O_1645,O_1646,O_1647,O_1648,O_1649,O_1650,O_1651,O_1652,O_1653,O_1654,O_1655,O_1656,O_1657,O_1658,O_1659,O_1660,O_1661,O_1662,O_1663,O_1664,O_1665,O_1666,O_1667,O_1668,O_1669,O_1670,O_1671,O_1672,O_1673,O_1674,O_1675,O_1676,O_1677,O_1678,O_1679,O_1680,O_1681,O_1682,O_1683,O_1684,O_1685,O_1686,O_1687,O_1688,O_1689,O_1690,O_1691,O_1692,O_1693,O_1694,O_1695,O_1696,O_1697,O_1698,O_1699,O_1700,O_1701,O_1702,O_1703,O_1704,O_1705,O_1706,O_1707,O_1708,O_1709,O_1710,O_1711,O_1712,O_1713,O_1714,O_1715,O_1716,O_1717,O_1718,O_1719,O_1720,O_1721,O_1722,O_1723,O_1724,O_1725,O_1726,O_1727,O_1728,O_1729,O_1730,O_1731,O_1732,O_1733,O_1734,O_1735,O_1736,O_1737,O_1738,O_1739,O_1740,O_1741,O_1742,O_1743,O_1744,O_1745,O_1746,O_1747,O_1748,O_1749,O_1750,O_1751,O_1752,O_1753,O_1754,O_1755,O_1756,O_1757,O_1758,O_1759,O_1760,O_1761,O_1762,O_1763,O_1764,O_1765,O_1766,O_1767,O_1768,O_1769,O_1770,O_1771,O_1772,O_1773,O_1774,O_1775,O_1776,O_1777,O_1778,O_1779,O_1780,O_1781,O_1782,O_1783,O_1784,O_1785,O_1786,O_1787,O_1788,O_1789,O_1790,O_1791,O_1792,O_1793,O_1794,O_1795,O_1796,O_1797,O_1798,O_1799,O_1800,O_1801,O_1802,O_1803,O_1804,O_1805,O_1806,O_1807,O_1808,O_1809,O_1810,O_1811,O_1812,O_1813,O_1814,O_1815,O_1816,O_1817,O_1818,O_1819,O_1820,O_1821,O_1822,O_1823,O_1824,O_1825,O_1826,O_1827,O_1828,O_1829,O_1830,O_1831,O_1832,O_1833,O_1834,O_1835,O_1836,O_1837,O_1838,O_1839,O_1840,O_1841,O_1842,O_1843,O_1844,O_1845,O_1846,O_1847,O_1848,O_1849,O_1850,O_1851,O_1852,O_1853,O_1854,O_1855,O_1856,O_1857,O_1858,O_1859,O_1860,O_1861,O_1862,O_1863,O_1864,O_1865,O_1866,O_1867,O_1868,O_1869,O_1870,O_1871,O_1872,O_1873,O_1874,O_1875,O_1876,O_1877,O_1878,O_1879,O_1880,O_1881,O_1882,O_1883,O_1884,O_1885,O_1886,O_1887,O_1888,O_1889,O_1890,O_1891,O_1892,O_1893,O_1894,O_1895,O_1896,O_1897,O_1898,O_1899,O_1900,O_1901,O_1902,O_1903,O_1904,O_1905,O_1906,O_1907,O_1908,O_1909,O_1910,O_1911,O_1912,O_1913,O_1914,O_1915,O_1916,O_1917,O_1918,O_1919,O_1920,O_1921,O_1922,O_1923,O_1924,O_1925,O_1926,O_1927,O_1928,O_1929,O_1930,O_1931,O_1932,O_1933,O_1934,O_1935,O_1936,O_1937,O_1938,O_1939,O_1940,O_1941,O_1942,O_1943,O_1944,O_1945,O_1946,O_1947,O_1948,O_1949,O_1950,O_1951,O_1952,O_1953,O_1954,O_1955,O_1956,O_1957,O_1958,O_1959,O_1960,O_1961,O_1962,O_1963,O_1964,O_1965,O_1966,O_1967,O_1968,O_1969,O_1970,O_1971,O_1972,O_1973,O_1974,O_1975,O_1976,O_1977,O_1978,O_1979,O_1980,O_1981,O_1982,O_1983,O_1984,O_1985,O_1986,O_1987,O_1988,O_1989,O_1990,O_1991,O_1992,O_1993,O_1994,O_1995,O_1996,O_1997,O_1998,O_1999,O_2000,O_2001,O_2002,O_2003,O_2004,O_2005,O_2006,O_2007,O_2008,O_2009,O_2010,O_2011,O_2012,O_2013,O_2014,O_2015,O_2016,O_2017,O_2018,O_2019,O_2020,O_2021,O_2022,O_2023,O_2024,O_2025,O_2026,O_2027,O_2028,O_2029,O_2030,O_2031,O_2032,O_2033,O_2034,O_2035,O_2036,O_2037,O_2038,O_2039,O_2040,O_2041,O_2042,O_2043,O_2044,O_2045,O_2046,O_2047,O_2048,O_2049,O_2050,O_2051,O_2052,O_2053,O_2054,O_2055,O_2056,O_2057,O_2058,O_2059,O_2060,O_2061,O_2062,O_2063,O_2064,O_2065,O_2066,O_2067,O_2068,O_2069,O_2070,O_2071,O_2072,O_2073,O_2074,O_2075,O_2076,O_2077,O_2078,O_2079,O_2080,O_2081,O_2082,O_2083,O_2084,O_2085,O_2086,O_2087,O_2088,O_2089,O_2090,O_2091,O_2092,O_2093,O_2094,O_2095,O_2096,O_2097,O_2098,O_2099,O_2100,O_2101,O_2102,O_2103,O_2104,O_2105,O_2106,O_2107,O_2108,O_2109,O_2110,O_2111,O_2112,O_2113,O_2114,O_2115,O_2116,O_2117,O_2118,O_2119,O_2120,O_2121,O_2122,O_2123,O_2124,O_2125,O_2126,O_2127,O_2128,O_2129,O_2130,O_2131,O_2132,O_2133,O_2134,O_2135,O_2136,O_2137,O_2138,O_2139,O_2140,O_2141,O_2142,O_2143,O_2144,O_2145,O_2146,O_2147,O_2148,O_2149,O_2150,O_2151,O_2152,O_2153,O_2154,O_2155,O_2156,O_2157,O_2158,O_2159,O_2160,O_2161,O_2162,O_2163,O_2164,O_2165,O_2166,O_2167,O_2168,O_2169,O_2170,O_2171,O_2172,O_2173,O_2174,O_2175,O_2176,O_2177,O_2178,O_2179,O_2180,O_2181,O_2182,O_2183,O_2184,O_2185,O_2186,O_2187,O_2188,O_2189,O_2190,O_2191,O_2192,O_2193,O_2194,O_2195,O_2196,O_2197,O_2198,O_2199,O_2200,O_2201,O_2202,O_2203,O_2204,O_2205,O_2206,O_2207,O_2208,O_2209,O_2210,O_2211,O_2212,O_2213,O_2214,O_2215,O_2216,O_2217,O_2218,O_2219,O_2220,O_2221,O_2222,O_2223,O_2224,O_2225,O_2226,O_2227,O_2228,O_2229,O_2230,O_2231,O_2232,O_2233,O_2234,O_2235,O_2236,O_2237,O_2238,O_2239,O_2240,O_2241,O_2242,O_2243,O_2244,O_2245,O_2246,O_2247,O_2248,O_2249,O_2250,O_2251,O_2252,O_2253,O_2254,O_2255,O_2256,O_2257,O_2258,O_2259,O_2260,O_2261,O_2262,O_2263,O_2264,O_2265,O_2266,O_2267,O_2268,O_2269,O_2270,O_2271,O_2272,O_2273,O_2274,O_2275,O_2276,O_2277,O_2278,O_2279,O_2280,O_2281,O_2282,O_2283,O_2284,O_2285,O_2286,O_2287,O_2288,O_2289,O_2290,O_2291,O_2292,O_2293,O_2294,O_2295,O_2296,O_2297,O_2298,O_2299,O_2300,O_2301,O_2302,O_2303,O_2304,O_2305,O_2306,O_2307,O_2308,O_2309,O_2310,O_2311,O_2312,O_2313,O_2314,O_2315,O_2316,O_2317,O_2318,O_2319,O_2320,O_2321,O_2322,O_2323,O_2324,O_2325,O_2326,O_2327,O_2328,O_2329,O_2330,O_2331,O_2332,O_2333,O_2334,O_2335,O_2336,O_2337,O_2338,O_2339,O_2340,O_2341,O_2342,O_2343,O_2344,O_2345,O_2346,O_2347,O_2348,O_2349,O_2350,O_2351,O_2352,O_2353,O_2354,O_2355,O_2356,O_2357,O_2358,O_2359,O_2360,O_2361,O_2362,O_2363,O_2364,O_2365,O_2366,O_2367,O_2368,O_2369,O_2370,O_2371,O_2372,O_2373,O_2374,O_2375,O_2376,O_2377,O_2378,O_2379,O_2380,O_2381,O_2382,O_2383,O_2384,O_2385,O_2386,O_2387,O_2388,O_2389,O_2390,O_2391,O_2392,O_2393,O_2394,O_2395,O_2396,O_2397,O_2398,O_2399,O_2400,O_2401,O_2402,O_2403,O_2404,O_2405,O_2406,O_2407,O_2408,O_2409,O_2410,O_2411,O_2412,O_2413,O_2414,O_2415,O_2416,O_2417,O_2418,O_2419,O_2420,O_2421,O_2422,O_2423,O_2424,O_2425,O_2426,O_2427,O_2428,O_2429,O_2430,O_2431,O_2432,O_2433,O_2434,O_2435,O_2436,O_2437,O_2438,O_2439,O_2440,O_2441,O_2442,O_2443,O_2444,O_2445,O_2446,O_2447,O_2448,O_2449,O_2450,O_2451,O_2452,O_2453,O_2454,O_2455,O_2456,O_2457,O_2458,O_2459,O_2460,O_2461,O_2462,O_2463,O_2464,O_2465,O_2466,O_2467,O_2468,O_2469,O_2470,O_2471,O_2472,O_2473,O_2474,O_2475,O_2476,O_2477,O_2478,O_2479,O_2480,O_2481,O_2482,O_2483,O_2484,O_2485,O_2486,O_2487,O_2488,O_2489,O_2490,O_2491,O_2492,O_2493,O_2494,O_2495,O_2496,O_2497,O_2498,O_2499,O_2500,O_2501,O_2502,O_2503,O_2504,O_2505,O_2506,O_2507,O_2508,O_2509,O_2510,O_2511,O_2512,O_2513,O_2514,O_2515,O_2516,O_2517,O_2518,O_2519,O_2520,O_2521,O_2522,O_2523,O_2524,O_2525,O_2526,O_2527,O_2528,O_2529,O_2530,O_2531,O_2532,O_2533,O_2534,O_2535,O_2536,O_2537,O_2538,O_2539,O_2540,O_2541,O_2542,O_2543,O_2544,O_2545,O_2546,O_2547,O_2548,O_2549,O_2550,O_2551,O_2552,O_2553,O_2554,O_2555,O_2556,O_2557,O_2558,O_2559,O_2560,O_2561,O_2562,O_2563,O_2564,O_2565,O_2566,O_2567,O_2568,O_2569,O_2570,O_2571,O_2572,O_2573,O_2574,O_2575,O_2576,O_2577,O_2578,O_2579,O_2580,O_2581,O_2582,O_2583,O_2584,O_2585,O_2586,O_2587,O_2588,O_2589,O_2590,O_2591,O_2592,O_2593,O_2594,O_2595,O_2596,O_2597,O_2598,O_2599,O_2600,O_2601,O_2602,O_2603,O_2604,O_2605,O_2606,O_2607,O_2608,O_2609,O_2610,O_2611,O_2612,O_2613,O_2614,O_2615,O_2616,O_2617,O_2618,O_2619,O_2620,O_2621,O_2622,O_2623,O_2624,O_2625,O_2626,O_2627,O_2628,O_2629,O_2630,O_2631,O_2632,O_2633,O_2634,O_2635,O_2636,O_2637,O_2638,O_2639,O_2640,O_2641,O_2642,O_2643,O_2644,O_2645,O_2646,O_2647,O_2648,O_2649,O_2650,O_2651,O_2652,O_2653,O_2654,O_2655,O_2656,O_2657,O_2658,O_2659,O_2660,O_2661,O_2662,O_2663,O_2664,O_2665,O_2666,O_2667,O_2668,O_2669,O_2670,O_2671,O_2672,O_2673,O_2674,O_2675,O_2676,O_2677,O_2678,O_2679,O_2680,O_2681,O_2682,O_2683,O_2684,O_2685,O_2686,O_2687,O_2688,O_2689,O_2690,O_2691,O_2692,O_2693,O_2694,O_2695,O_2696,O_2697,O_2698,O_2699,O_2700,O_2701,O_2702,O_2703,O_2704,O_2705,O_2706,O_2707,O_2708,O_2709,O_2710,O_2711,O_2712,O_2713,O_2714,O_2715,O_2716,O_2717,O_2718,O_2719,O_2720,O_2721,O_2722,O_2723,O_2724,O_2725,O_2726,O_2727,O_2728,O_2729,O_2730,O_2731,O_2732,O_2733,O_2734,O_2735,O_2736,O_2737,O_2738,O_2739,O_2740,O_2741,O_2742,O_2743,O_2744,O_2745,O_2746,O_2747,O_2748,O_2749,O_2750,O_2751,O_2752,O_2753,O_2754,O_2755,O_2756,O_2757,O_2758,O_2759,O_2760,O_2761,O_2762,O_2763,O_2764,O_2765,O_2766,O_2767,O_2768,O_2769,O_2770,O_2771,O_2772,O_2773,O_2774,O_2775,O_2776,O_2777,O_2778,O_2779,O_2780,O_2781,O_2782,O_2783,O_2784,O_2785,O_2786,O_2787,O_2788,O_2789,O_2790,O_2791,O_2792,O_2793,O_2794,O_2795,O_2796,O_2797,O_2798,O_2799,O_2800,O_2801,O_2802,O_2803,O_2804,O_2805,O_2806,O_2807,O_2808,O_2809,O_2810,O_2811,O_2812,O_2813,O_2814,O_2815,O_2816,O_2817,O_2818,O_2819,O_2820,O_2821,O_2822,O_2823,O_2824,O_2825,O_2826,O_2827,O_2828,O_2829,O_2830,O_2831,O_2832,O_2833,O_2834,O_2835,O_2836,O_2837,O_2838,O_2839,O_2840,O_2841,O_2842,O_2843,O_2844,O_2845,O_2846,O_2847,O_2848,O_2849,O_2850,O_2851,O_2852,O_2853,O_2854,O_2855,O_2856,O_2857,O_2858,O_2859,O_2860,O_2861,O_2862,O_2863,O_2864,O_2865,O_2866,O_2867,O_2868,O_2869,O_2870,O_2871,O_2872,O_2873,O_2874,O_2875,O_2876,O_2877,O_2878,O_2879,O_2880,O_2881,O_2882,O_2883,O_2884,O_2885,O_2886,O_2887,O_2888,O_2889,O_2890,O_2891,O_2892,O_2893,O_2894,O_2895,O_2896,O_2897,O_2898,O_2899,O_2900,O_2901,O_2902,O_2903,O_2904,O_2905,O_2906,O_2907,O_2908,O_2909,O_2910,O_2911,O_2912,O_2913,O_2914,O_2915,O_2916,O_2917,O_2918,O_2919,O_2920,O_2921,O_2922,O_2923,O_2924,O_2925,O_2926,O_2927,O_2928,O_2929,O_2930,O_2931,O_2932,O_2933,O_2934,O_2935,O_2936,O_2937,O_2938,O_2939,O_2940,O_2941,O_2942,O_2943,O_2944,O_2945,O_2946,O_2947,O_2948,O_2949,O_2950,O_2951,O_2952,O_2953,O_2954,O_2955,O_2956,O_2957,O_2958,O_2959,O_2960,O_2961,O_2962,O_2963,O_2964,O_2965,O_2966,O_2967,O_2968,O_2969,O_2970,O_2971,O_2972,O_2973,O_2974,O_2975,O_2976,O_2977,O_2978,O_2979,O_2980,O_2981,O_2982,O_2983,O_2984,O_2985,O_2986,O_2987,O_2988,O_2989,O_2990,O_2991,O_2992,O_2993,O_2994,O_2995,O_2996,O_2997,O_2998,O_2999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999,N_5000,N_5001,N_5002,N_5003,N_5004,N_5005,N_5006,N_5007,N_5008,N_5009,N_5010,N_5011,N_5012,N_5013,N_5014,N_5015,N_5016,N_5017,N_5018,N_5019,N_5020,N_5021,N_5022,N_5023,N_5024,N_5025,N_5026,N_5027,N_5028,N_5029,N_5030,N_5031,N_5032,N_5033,N_5034,N_5035,N_5036,N_5037,N_5038,N_5039,N_5040,N_5041,N_5042,N_5043,N_5044,N_5045,N_5046,N_5047,N_5048,N_5049,N_5050,N_5051,N_5052,N_5053,N_5054,N_5055,N_5056,N_5057,N_5058,N_5059,N_5060,N_5061,N_5062,N_5063,N_5064,N_5065,N_5066,N_5067,N_5068,N_5069,N_5070,N_5071,N_5072,N_5073,N_5074,N_5075,N_5076,N_5077,N_5078,N_5079,N_5080,N_5081,N_5082,N_5083,N_5084,N_5085,N_5086,N_5087,N_5088,N_5089,N_5090,N_5091,N_5092,N_5093,N_5094,N_5095,N_5096,N_5097,N_5098,N_5099,N_5100,N_5101,N_5102,N_5103,N_5104,N_5105,N_5106,N_5107,N_5108,N_5109,N_5110,N_5111,N_5112,N_5113,N_5114,N_5115,N_5116,N_5117,N_5118,N_5119,N_5120,N_5121,N_5122,N_5123,N_5124,N_5125,N_5126,N_5127,N_5128,N_5129,N_5130,N_5131,N_5132,N_5133,N_5134,N_5135,N_5136,N_5137,N_5138,N_5139,N_5140,N_5141,N_5142,N_5143,N_5144,N_5145,N_5146,N_5147,N_5148,N_5149,N_5150,N_5151,N_5152,N_5153,N_5154,N_5155,N_5156,N_5157,N_5158,N_5159,N_5160,N_5161,N_5162,N_5163,N_5164,N_5165,N_5166,N_5167,N_5168,N_5169,N_5170,N_5171,N_5172,N_5173,N_5174,N_5175,N_5176,N_5177,N_5178,N_5179,N_5180,N_5181,N_5182,N_5183,N_5184,N_5185,N_5186,N_5187,N_5188,N_5189,N_5190,N_5191,N_5192,N_5193,N_5194,N_5195,N_5196,N_5197,N_5198,N_5199,N_5200,N_5201,N_5202,N_5203,N_5204,N_5205,N_5206,N_5207,N_5208,N_5209,N_5210,N_5211,N_5212,N_5213,N_5214,N_5215,N_5216,N_5217,N_5218,N_5219,N_5220,N_5221,N_5222,N_5223,N_5224,N_5225,N_5226,N_5227,N_5228,N_5229,N_5230,N_5231,N_5232,N_5233,N_5234,N_5235,N_5236,N_5237,N_5238,N_5239,N_5240,N_5241,N_5242,N_5243,N_5244,N_5245,N_5246,N_5247,N_5248,N_5249,N_5250,N_5251,N_5252,N_5253,N_5254,N_5255,N_5256,N_5257,N_5258,N_5259,N_5260,N_5261,N_5262,N_5263,N_5264,N_5265,N_5266,N_5267,N_5268,N_5269,N_5270,N_5271,N_5272,N_5273,N_5274,N_5275,N_5276,N_5277,N_5278,N_5279,N_5280,N_5281,N_5282,N_5283,N_5284,N_5285,N_5286,N_5287,N_5288,N_5289,N_5290,N_5291,N_5292,N_5293,N_5294,N_5295,N_5296,N_5297,N_5298,N_5299,N_5300,N_5301,N_5302,N_5303,N_5304,N_5305,N_5306,N_5307,N_5308,N_5309,N_5310,N_5311,N_5312,N_5313,N_5314,N_5315,N_5316,N_5317,N_5318,N_5319,N_5320,N_5321,N_5322,N_5323,N_5324,N_5325,N_5326,N_5327,N_5328,N_5329,N_5330,N_5331,N_5332,N_5333,N_5334,N_5335,N_5336,N_5337,N_5338,N_5339,N_5340,N_5341,N_5342,N_5343,N_5344,N_5345,N_5346,N_5347,N_5348,N_5349,N_5350,N_5351,N_5352,N_5353,N_5354,N_5355,N_5356,N_5357,N_5358,N_5359,N_5360,N_5361,N_5362,N_5363,N_5364,N_5365,N_5366,N_5367,N_5368,N_5369,N_5370,N_5371,N_5372,N_5373,N_5374,N_5375,N_5376,N_5377,N_5378,N_5379,N_5380,N_5381,N_5382,N_5383,N_5384,N_5385,N_5386,N_5387,N_5388,N_5389,N_5390,N_5391,N_5392,N_5393,N_5394,N_5395,N_5396,N_5397,N_5398,N_5399,N_5400,N_5401,N_5402,N_5403,N_5404,N_5405,N_5406,N_5407,N_5408,N_5409,N_5410,N_5411,N_5412,N_5413,N_5414,N_5415,N_5416,N_5417,N_5418,N_5419,N_5420,N_5421,N_5422,N_5423,N_5424,N_5425,N_5426,N_5427,N_5428,N_5429,N_5430,N_5431,N_5432,N_5433,N_5434,N_5435,N_5436,N_5437,N_5438,N_5439,N_5440,N_5441,N_5442,N_5443,N_5444,N_5445,N_5446,N_5447,N_5448,N_5449,N_5450,N_5451,N_5452,N_5453,N_5454,N_5455,N_5456,N_5457,N_5458,N_5459,N_5460,N_5461,N_5462,N_5463,N_5464,N_5465,N_5466,N_5467,N_5468,N_5469,N_5470,N_5471,N_5472,N_5473,N_5474,N_5475,N_5476,N_5477,N_5478,N_5479,N_5480,N_5481,N_5482,N_5483,N_5484,N_5485,N_5486,N_5487,N_5488,N_5489,N_5490,N_5491,N_5492,N_5493,N_5494,N_5495,N_5496,N_5497,N_5498,N_5499,N_5500,N_5501,N_5502,N_5503,N_5504,N_5505,N_5506,N_5507,N_5508,N_5509,N_5510,N_5511,N_5512,N_5513,N_5514,N_5515,N_5516,N_5517,N_5518,N_5519,N_5520,N_5521,N_5522,N_5523,N_5524,N_5525,N_5526,N_5527,N_5528,N_5529,N_5530,N_5531,N_5532,N_5533,N_5534,N_5535,N_5536,N_5537,N_5538,N_5539,N_5540,N_5541,N_5542,N_5543,N_5544,N_5545,N_5546,N_5547,N_5548,N_5549,N_5550,N_5551,N_5552,N_5553,N_5554,N_5555,N_5556,N_5557,N_5558,N_5559,N_5560,N_5561,N_5562,N_5563,N_5564,N_5565,N_5566,N_5567,N_5568,N_5569,N_5570,N_5571,N_5572,N_5573,N_5574,N_5575,N_5576,N_5577,N_5578,N_5579,N_5580,N_5581,N_5582,N_5583,N_5584,N_5585,N_5586,N_5587,N_5588,N_5589,N_5590,N_5591,N_5592,N_5593,N_5594,N_5595,N_5596,N_5597,N_5598,N_5599,N_5600,N_5601,N_5602,N_5603,N_5604,N_5605,N_5606,N_5607,N_5608,N_5609,N_5610,N_5611,N_5612,N_5613,N_5614,N_5615,N_5616,N_5617,N_5618,N_5619,N_5620,N_5621,N_5622,N_5623,N_5624,N_5625,N_5626,N_5627,N_5628,N_5629,N_5630,N_5631,N_5632,N_5633,N_5634,N_5635,N_5636,N_5637,N_5638,N_5639,N_5640,N_5641,N_5642,N_5643,N_5644,N_5645,N_5646,N_5647,N_5648,N_5649,N_5650,N_5651,N_5652,N_5653,N_5654,N_5655,N_5656,N_5657,N_5658,N_5659,N_5660,N_5661,N_5662,N_5663,N_5664,N_5665,N_5666,N_5667,N_5668,N_5669,N_5670,N_5671,N_5672,N_5673,N_5674,N_5675,N_5676,N_5677,N_5678,N_5679,N_5680,N_5681,N_5682,N_5683,N_5684,N_5685,N_5686,N_5687,N_5688,N_5689,N_5690,N_5691,N_5692,N_5693,N_5694,N_5695,N_5696,N_5697,N_5698,N_5699,N_5700,N_5701,N_5702,N_5703,N_5704,N_5705,N_5706,N_5707,N_5708,N_5709,N_5710,N_5711,N_5712,N_5713,N_5714,N_5715,N_5716,N_5717,N_5718,N_5719,N_5720,N_5721,N_5722,N_5723,N_5724,N_5725,N_5726,N_5727,N_5728,N_5729,N_5730,N_5731,N_5732,N_5733,N_5734,N_5735,N_5736,N_5737,N_5738,N_5739,N_5740,N_5741,N_5742,N_5743,N_5744,N_5745,N_5746,N_5747,N_5748,N_5749,N_5750,N_5751,N_5752,N_5753,N_5754,N_5755,N_5756,N_5757,N_5758,N_5759,N_5760,N_5761,N_5762,N_5763,N_5764,N_5765,N_5766,N_5767,N_5768,N_5769,N_5770,N_5771,N_5772,N_5773,N_5774,N_5775,N_5776,N_5777,N_5778,N_5779,N_5780,N_5781,N_5782,N_5783,N_5784,N_5785,N_5786,N_5787,N_5788,N_5789,N_5790,N_5791,N_5792,N_5793,N_5794,N_5795,N_5796,N_5797,N_5798,N_5799,N_5800,N_5801,N_5802,N_5803,N_5804,N_5805,N_5806,N_5807,N_5808,N_5809,N_5810,N_5811,N_5812,N_5813,N_5814,N_5815,N_5816,N_5817,N_5818,N_5819,N_5820,N_5821,N_5822,N_5823,N_5824,N_5825,N_5826,N_5827,N_5828,N_5829,N_5830,N_5831,N_5832,N_5833,N_5834,N_5835,N_5836,N_5837,N_5838,N_5839,N_5840,N_5841,N_5842,N_5843,N_5844,N_5845,N_5846,N_5847,N_5848,N_5849,N_5850,N_5851,N_5852,N_5853,N_5854,N_5855,N_5856,N_5857,N_5858,N_5859,N_5860,N_5861,N_5862,N_5863,N_5864,N_5865,N_5866,N_5867,N_5868,N_5869,N_5870,N_5871,N_5872,N_5873,N_5874,N_5875,N_5876,N_5877,N_5878,N_5879,N_5880,N_5881,N_5882,N_5883,N_5884,N_5885,N_5886,N_5887,N_5888,N_5889,N_5890,N_5891,N_5892,N_5893,N_5894,N_5895,N_5896,N_5897,N_5898,N_5899,N_5900,N_5901,N_5902,N_5903,N_5904,N_5905,N_5906,N_5907,N_5908,N_5909,N_5910,N_5911,N_5912,N_5913,N_5914,N_5915,N_5916,N_5917,N_5918,N_5919,N_5920,N_5921,N_5922,N_5923,N_5924,N_5925,N_5926,N_5927,N_5928,N_5929,N_5930,N_5931,N_5932,N_5933,N_5934,N_5935,N_5936,N_5937,N_5938,N_5939,N_5940,N_5941,N_5942,N_5943,N_5944,N_5945,N_5946,N_5947,N_5948,N_5949,N_5950,N_5951,N_5952,N_5953,N_5954,N_5955,N_5956,N_5957,N_5958,N_5959,N_5960,N_5961,N_5962,N_5963,N_5964,N_5965,N_5966,N_5967,N_5968,N_5969,N_5970,N_5971,N_5972,N_5973,N_5974,N_5975,N_5976,N_5977,N_5978,N_5979,N_5980,N_5981,N_5982,N_5983,N_5984,N_5985,N_5986,N_5987,N_5988,N_5989,N_5990,N_5991,N_5992,N_5993,N_5994,N_5995,N_5996,N_5997,N_5998,N_5999,N_6000,N_6001,N_6002,N_6003,N_6004,N_6005,N_6006,N_6007,N_6008,N_6009,N_6010,N_6011,N_6012,N_6013,N_6014,N_6015,N_6016,N_6017,N_6018,N_6019,N_6020,N_6021,N_6022,N_6023,N_6024,N_6025,N_6026,N_6027,N_6028,N_6029,N_6030,N_6031,N_6032,N_6033,N_6034,N_6035,N_6036,N_6037,N_6038,N_6039,N_6040,N_6041,N_6042,N_6043,N_6044,N_6045,N_6046,N_6047,N_6048,N_6049,N_6050,N_6051,N_6052,N_6053,N_6054,N_6055,N_6056,N_6057,N_6058,N_6059,N_6060,N_6061,N_6062,N_6063,N_6064,N_6065,N_6066,N_6067,N_6068,N_6069,N_6070,N_6071,N_6072,N_6073,N_6074,N_6075,N_6076,N_6077,N_6078,N_6079,N_6080,N_6081,N_6082,N_6083,N_6084,N_6085,N_6086,N_6087,N_6088,N_6089,N_6090,N_6091,N_6092,N_6093,N_6094,N_6095,N_6096,N_6097,N_6098,N_6099,N_6100,N_6101,N_6102,N_6103,N_6104,N_6105,N_6106,N_6107,N_6108,N_6109,N_6110,N_6111,N_6112,N_6113,N_6114,N_6115,N_6116,N_6117,N_6118,N_6119,N_6120,N_6121,N_6122,N_6123,N_6124,N_6125,N_6126,N_6127,N_6128,N_6129,N_6130,N_6131,N_6132,N_6133,N_6134,N_6135,N_6136,N_6137,N_6138,N_6139,N_6140,N_6141,N_6142,N_6143,N_6144,N_6145,N_6146,N_6147,N_6148,N_6149,N_6150,N_6151,N_6152,N_6153,N_6154,N_6155,N_6156,N_6157,N_6158,N_6159,N_6160,N_6161,N_6162,N_6163,N_6164,N_6165,N_6166,N_6167,N_6168,N_6169,N_6170,N_6171,N_6172,N_6173,N_6174,N_6175,N_6176,N_6177,N_6178,N_6179,N_6180,N_6181,N_6182,N_6183,N_6184,N_6185,N_6186,N_6187,N_6188,N_6189,N_6190,N_6191,N_6192,N_6193,N_6194,N_6195,N_6196,N_6197,N_6198,N_6199,N_6200,N_6201,N_6202,N_6203,N_6204,N_6205,N_6206,N_6207,N_6208,N_6209,N_6210,N_6211,N_6212,N_6213,N_6214,N_6215,N_6216,N_6217,N_6218,N_6219,N_6220,N_6221,N_6222,N_6223,N_6224,N_6225,N_6226,N_6227,N_6228,N_6229,N_6230,N_6231,N_6232,N_6233,N_6234,N_6235,N_6236,N_6237,N_6238,N_6239,N_6240,N_6241,N_6242,N_6243,N_6244,N_6245,N_6246,N_6247,N_6248,N_6249,N_6250,N_6251,N_6252,N_6253,N_6254,N_6255,N_6256,N_6257,N_6258,N_6259,N_6260,N_6261,N_6262,N_6263,N_6264,N_6265,N_6266,N_6267,N_6268,N_6269,N_6270,N_6271,N_6272,N_6273,N_6274,N_6275,N_6276,N_6277,N_6278,N_6279,N_6280,N_6281,N_6282,N_6283,N_6284,N_6285,N_6286,N_6287,N_6288,N_6289,N_6290,N_6291,N_6292,N_6293,N_6294,N_6295,N_6296,N_6297,N_6298,N_6299,N_6300,N_6301,N_6302,N_6303,N_6304,N_6305,N_6306,N_6307,N_6308,N_6309,N_6310,N_6311,N_6312,N_6313,N_6314,N_6315,N_6316,N_6317,N_6318,N_6319,N_6320,N_6321,N_6322,N_6323,N_6324,N_6325,N_6326,N_6327,N_6328,N_6329,N_6330,N_6331,N_6332,N_6333,N_6334,N_6335,N_6336,N_6337,N_6338,N_6339,N_6340,N_6341,N_6342,N_6343,N_6344,N_6345,N_6346,N_6347,N_6348,N_6349,N_6350,N_6351,N_6352,N_6353,N_6354,N_6355,N_6356,N_6357,N_6358,N_6359,N_6360,N_6361,N_6362,N_6363,N_6364,N_6365,N_6366,N_6367,N_6368,N_6369,N_6370,N_6371,N_6372,N_6373,N_6374,N_6375,N_6376,N_6377,N_6378,N_6379,N_6380,N_6381,N_6382,N_6383,N_6384,N_6385,N_6386,N_6387,N_6388,N_6389,N_6390,N_6391,N_6392,N_6393,N_6394,N_6395,N_6396,N_6397,N_6398,N_6399,N_6400,N_6401,N_6402,N_6403,N_6404,N_6405,N_6406,N_6407,N_6408,N_6409,N_6410,N_6411,N_6412,N_6413,N_6414,N_6415,N_6416,N_6417,N_6418,N_6419,N_6420,N_6421,N_6422,N_6423,N_6424,N_6425,N_6426,N_6427,N_6428,N_6429,N_6430,N_6431,N_6432,N_6433,N_6434,N_6435,N_6436,N_6437,N_6438,N_6439,N_6440,N_6441,N_6442,N_6443,N_6444,N_6445,N_6446,N_6447,N_6448,N_6449,N_6450,N_6451,N_6452,N_6453,N_6454,N_6455,N_6456,N_6457,N_6458,N_6459,N_6460,N_6461,N_6462,N_6463,N_6464,N_6465,N_6466,N_6467,N_6468,N_6469,N_6470,N_6471,N_6472,N_6473,N_6474,N_6475,N_6476,N_6477,N_6478,N_6479,N_6480,N_6481,N_6482,N_6483,N_6484,N_6485,N_6486,N_6487,N_6488,N_6489,N_6490,N_6491,N_6492,N_6493,N_6494,N_6495,N_6496,N_6497,N_6498,N_6499,N_6500,N_6501,N_6502,N_6503,N_6504,N_6505,N_6506,N_6507,N_6508,N_6509,N_6510,N_6511,N_6512,N_6513,N_6514,N_6515,N_6516,N_6517,N_6518,N_6519,N_6520,N_6521,N_6522,N_6523,N_6524,N_6525,N_6526,N_6527,N_6528,N_6529,N_6530,N_6531,N_6532,N_6533,N_6534,N_6535,N_6536,N_6537,N_6538,N_6539,N_6540,N_6541,N_6542,N_6543,N_6544,N_6545,N_6546,N_6547,N_6548,N_6549,N_6550,N_6551,N_6552,N_6553,N_6554,N_6555,N_6556,N_6557,N_6558,N_6559,N_6560,N_6561,N_6562,N_6563,N_6564,N_6565,N_6566,N_6567,N_6568,N_6569,N_6570,N_6571,N_6572,N_6573,N_6574,N_6575,N_6576,N_6577,N_6578,N_6579,N_6580,N_6581,N_6582,N_6583,N_6584,N_6585,N_6586,N_6587,N_6588,N_6589,N_6590,N_6591,N_6592,N_6593,N_6594,N_6595,N_6596,N_6597,N_6598,N_6599,N_6600,N_6601,N_6602,N_6603,N_6604,N_6605,N_6606,N_6607,N_6608,N_6609,N_6610,N_6611,N_6612,N_6613,N_6614,N_6615,N_6616,N_6617,N_6618,N_6619,N_6620,N_6621,N_6622,N_6623,N_6624,N_6625,N_6626,N_6627,N_6628,N_6629,N_6630,N_6631,N_6632,N_6633,N_6634,N_6635,N_6636,N_6637,N_6638,N_6639,N_6640,N_6641,N_6642,N_6643,N_6644,N_6645,N_6646,N_6647,N_6648,N_6649,N_6650,N_6651,N_6652,N_6653,N_6654,N_6655,N_6656,N_6657,N_6658,N_6659,N_6660,N_6661,N_6662,N_6663,N_6664,N_6665,N_6666,N_6667,N_6668,N_6669,N_6670,N_6671,N_6672,N_6673,N_6674,N_6675,N_6676,N_6677,N_6678,N_6679,N_6680,N_6681,N_6682,N_6683,N_6684,N_6685,N_6686,N_6687,N_6688,N_6689,N_6690,N_6691,N_6692,N_6693,N_6694,N_6695,N_6696,N_6697,N_6698,N_6699,N_6700,N_6701,N_6702,N_6703,N_6704,N_6705,N_6706,N_6707,N_6708,N_6709,N_6710,N_6711,N_6712,N_6713,N_6714,N_6715,N_6716,N_6717,N_6718,N_6719,N_6720,N_6721,N_6722,N_6723,N_6724,N_6725,N_6726,N_6727,N_6728,N_6729,N_6730,N_6731,N_6732,N_6733,N_6734,N_6735,N_6736,N_6737,N_6738,N_6739,N_6740,N_6741,N_6742,N_6743,N_6744,N_6745,N_6746,N_6747,N_6748,N_6749,N_6750,N_6751,N_6752,N_6753,N_6754,N_6755,N_6756,N_6757,N_6758,N_6759,N_6760,N_6761,N_6762,N_6763,N_6764,N_6765,N_6766,N_6767,N_6768,N_6769,N_6770,N_6771,N_6772,N_6773,N_6774,N_6775,N_6776,N_6777,N_6778,N_6779,N_6780,N_6781,N_6782,N_6783,N_6784,N_6785,N_6786,N_6787,N_6788,N_6789,N_6790,N_6791,N_6792,N_6793,N_6794,N_6795,N_6796,N_6797,N_6798,N_6799,N_6800,N_6801,N_6802,N_6803,N_6804,N_6805,N_6806,N_6807,N_6808,N_6809,N_6810,N_6811,N_6812,N_6813,N_6814,N_6815,N_6816,N_6817,N_6818,N_6819,N_6820,N_6821,N_6822,N_6823,N_6824,N_6825,N_6826,N_6827,N_6828,N_6829,N_6830,N_6831,N_6832,N_6833,N_6834,N_6835,N_6836,N_6837,N_6838,N_6839,N_6840,N_6841,N_6842,N_6843,N_6844,N_6845,N_6846,N_6847,N_6848,N_6849,N_6850,N_6851,N_6852,N_6853,N_6854,N_6855,N_6856,N_6857,N_6858,N_6859,N_6860,N_6861,N_6862,N_6863,N_6864,N_6865,N_6866,N_6867,N_6868,N_6869,N_6870,N_6871,N_6872,N_6873,N_6874,N_6875,N_6876,N_6877,N_6878,N_6879,N_6880,N_6881,N_6882,N_6883,N_6884,N_6885,N_6886,N_6887,N_6888,N_6889,N_6890,N_6891,N_6892,N_6893,N_6894,N_6895,N_6896,N_6897,N_6898,N_6899,N_6900,N_6901,N_6902,N_6903,N_6904,N_6905,N_6906,N_6907,N_6908,N_6909,N_6910,N_6911,N_6912,N_6913,N_6914,N_6915,N_6916,N_6917,N_6918,N_6919,N_6920,N_6921,N_6922,N_6923,N_6924,N_6925,N_6926,N_6927,N_6928,N_6929,N_6930,N_6931,N_6932,N_6933,N_6934,N_6935,N_6936,N_6937,N_6938,N_6939,N_6940,N_6941,N_6942,N_6943,N_6944,N_6945,N_6946,N_6947,N_6948,N_6949,N_6950,N_6951,N_6952,N_6953,N_6954,N_6955,N_6956,N_6957,N_6958,N_6959,N_6960,N_6961,N_6962,N_6963,N_6964,N_6965,N_6966,N_6967,N_6968,N_6969,N_6970,N_6971,N_6972,N_6973,N_6974,N_6975,N_6976,N_6977,N_6978,N_6979,N_6980,N_6981,N_6982,N_6983,N_6984,N_6985,N_6986,N_6987,N_6988,N_6989,N_6990,N_6991,N_6992,N_6993,N_6994,N_6995,N_6996,N_6997,N_6998,N_6999,N_7000,N_7001,N_7002,N_7003,N_7004,N_7005,N_7006,N_7007,N_7008,N_7009,N_7010,N_7011,N_7012,N_7013,N_7014,N_7015,N_7016,N_7017,N_7018,N_7019,N_7020,N_7021,N_7022,N_7023,N_7024,N_7025,N_7026,N_7027,N_7028,N_7029,N_7030,N_7031,N_7032,N_7033,N_7034,N_7035,N_7036,N_7037,N_7038,N_7039,N_7040,N_7041,N_7042,N_7043,N_7044,N_7045,N_7046,N_7047,N_7048,N_7049,N_7050,N_7051,N_7052,N_7053,N_7054,N_7055,N_7056,N_7057,N_7058,N_7059,N_7060,N_7061,N_7062,N_7063,N_7064,N_7065,N_7066,N_7067,N_7068,N_7069,N_7070,N_7071,N_7072,N_7073,N_7074,N_7075,N_7076,N_7077,N_7078,N_7079,N_7080,N_7081,N_7082,N_7083,N_7084,N_7085,N_7086,N_7087,N_7088,N_7089,N_7090,N_7091,N_7092,N_7093,N_7094,N_7095,N_7096,N_7097,N_7098,N_7099,N_7100,N_7101,N_7102,N_7103,N_7104,N_7105,N_7106,N_7107,N_7108,N_7109,N_7110,N_7111,N_7112,N_7113,N_7114,N_7115,N_7116,N_7117,N_7118,N_7119,N_7120,N_7121,N_7122,N_7123,N_7124,N_7125,N_7126,N_7127,N_7128,N_7129,N_7130,N_7131,N_7132,N_7133,N_7134,N_7135,N_7136,N_7137,N_7138,N_7139,N_7140,N_7141,N_7142,N_7143,N_7144,N_7145,N_7146,N_7147,N_7148,N_7149,N_7150,N_7151,N_7152,N_7153,N_7154,N_7155,N_7156,N_7157,N_7158,N_7159,N_7160,N_7161,N_7162,N_7163,N_7164,N_7165,N_7166,N_7167,N_7168,N_7169,N_7170,N_7171,N_7172,N_7173,N_7174,N_7175,N_7176,N_7177,N_7178,N_7179,N_7180,N_7181,N_7182,N_7183,N_7184,N_7185,N_7186,N_7187,N_7188,N_7189,N_7190,N_7191,N_7192,N_7193,N_7194,N_7195,N_7196,N_7197,N_7198,N_7199,N_7200,N_7201,N_7202,N_7203,N_7204,N_7205,N_7206,N_7207,N_7208,N_7209,N_7210,N_7211,N_7212,N_7213,N_7214,N_7215,N_7216,N_7217,N_7218,N_7219,N_7220,N_7221,N_7222,N_7223,N_7224,N_7225,N_7226,N_7227,N_7228,N_7229,N_7230,N_7231,N_7232,N_7233,N_7234,N_7235,N_7236,N_7237,N_7238,N_7239,N_7240,N_7241,N_7242,N_7243,N_7244,N_7245,N_7246,N_7247,N_7248,N_7249,N_7250,N_7251,N_7252,N_7253,N_7254,N_7255,N_7256,N_7257,N_7258,N_7259,N_7260,N_7261,N_7262,N_7263,N_7264,N_7265,N_7266,N_7267,N_7268,N_7269,N_7270,N_7271,N_7272,N_7273,N_7274,N_7275,N_7276,N_7277,N_7278,N_7279,N_7280,N_7281,N_7282,N_7283,N_7284,N_7285,N_7286,N_7287,N_7288,N_7289,N_7290,N_7291,N_7292,N_7293,N_7294,N_7295,N_7296,N_7297,N_7298,N_7299,N_7300,N_7301,N_7302,N_7303,N_7304,N_7305,N_7306,N_7307,N_7308,N_7309,N_7310,N_7311,N_7312,N_7313,N_7314,N_7315,N_7316,N_7317,N_7318,N_7319,N_7320,N_7321,N_7322,N_7323,N_7324,N_7325,N_7326,N_7327,N_7328,N_7329,N_7330,N_7331,N_7332,N_7333,N_7334,N_7335,N_7336,N_7337,N_7338,N_7339,N_7340,N_7341,N_7342,N_7343,N_7344,N_7345,N_7346,N_7347,N_7348,N_7349,N_7350,N_7351,N_7352,N_7353,N_7354,N_7355,N_7356,N_7357,N_7358,N_7359,N_7360,N_7361,N_7362,N_7363,N_7364,N_7365,N_7366,N_7367,N_7368,N_7369,N_7370,N_7371,N_7372,N_7373,N_7374,N_7375,N_7376,N_7377,N_7378,N_7379,N_7380,N_7381,N_7382,N_7383,N_7384,N_7385,N_7386,N_7387,N_7388,N_7389,N_7390,N_7391,N_7392,N_7393,N_7394,N_7395,N_7396,N_7397,N_7398,N_7399,N_7400,N_7401,N_7402,N_7403,N_7404,N_7405,N_7406,N_7407,N_7408,N_7409,N_7410,N_7411,N_7412,N_7413,N_7414,N_7415,N_7416,N_7417,N_7418,N_7419,N_7420,N_7421,N_7422,N_7423,N_7424,N_7425,N_7426,N_7427,N_7428,N_7429,N_7430,N_7431,N_7432,N_7433,N_7434,N_7435,N_7436,N_7437,N_7438,N_7439,N_7440,N_7441,N_7442,N_7443,N_7444,N_7445,N_7446,N_7447,N_7448,N_7449,N_7450,N_7451,N_7452,N_7453,N_7454,N_7455,N_7456,N_7457,N_7458,N_7459,N_7460,N_7461,N_7462,N_7463,N_7464,N_7465,N_7466,N_7467,N_7468,N_7469,N_7470,N_7471,N_7472,N_7473,N_7474,N_7475,N_7476,N_7477,N_7478,N_7479,N_7480,N_7481,N_7482,N_7483,N_7484,N_7485,N_7486,N_7487,N_7488,N_7489,N_7490,N_7491,N_7492,N_7493,N_7494,N_7495,N_7496,N_7497,N_7498,N_7499,N_7500,N_7501,N_7502,N_7503,N_7504,N_7505,N_7506,N_7507,N_7508,N_7509,N_7510,N_7511,N_7512,N_7513,N_7514,N_7515,N_7516,N_7517,N_7518,N_7519,N_7520,N_7521,N_7522,N_7523,N_7524,N_7525,N_7526,N_7527,N_7528,N_7529,N_7530,N_7531,N_7532,N_7533,N_7534,N_7535,N_7536,N_7537,N_7538,N_7539,N_7540,N_7541,N_7542,N_7543,N_7544,N_7545,N_7546,N_7547,N_7548,N_7549,N_7550,N_7551,N_7552,N_7553,N_7554,N_7555,N_7556,N_7557,N_7558,N_7559,N_7560,N_7561,N_7562,N_7563,N_7564,N_7565,N_7566,N_7567,N_7568,N_7569,N_7570,N_7571,N_7572,N_7573,N_7574,N_7575,N_7576,N_7577,N_7578,N_7579,N_7580,N_7581,N_7582,N_7583,N_7584,N_7585,N_7586,N_7587,N_7588,N_7589,N_7590,N_7591,N_7592,N_7593,N_7594,N_7595,N_7596,N_7597,N_7598,N_7599,N_7600,N_7601,N_7602,N_7603,N_7604,N_7605,N_7606,N_7607,N_7608,N_7609,N_7610,N_7611,N_7612,N_7613,N_7614,N_7615,N_7616,N_7617,N_7618,N_7619,N_7620,N_7621,N_7622,N_7623,N_7624,N_7625,N_7626,N_7627,N_7628,N_7629,N_7630,N_7631,N_7632,N_7633,N_7634,N_7635,N_7636,N_7637,N_7638,N_7639,N_7640,N_7641,N_7642,N_7643,N_7644,N_7645,N_7646,N_7647,N_7648,N_7649,N_7650,N_7651,N_7652,N_7653,N_7654,N_7655,N_7656,N_7657,N_7658,N_7659,N_7660,N_7661,N_7662,N_7663,N_7664,N_7665,N_7666,N_7667,N_7668,N_7669,N_7670,N_7671,N_7672,N_7673,N_7674,N_7675,N_7676,N_7677,N_7678,N_7679,N_7680,N_7681,N_7682,N_7683,N_7684,N_7685,N_7686,N_7687,N_7688,N_7689,N_7690,N_7691,N_7692,N_7693,N_7694,N_7695,N_7696,N_7697,N_7698,N_7699,N_7700,N_7701,N_7702,N_7703,N_7704,N_7705,N_7706,N_7707,N_7708,N_7709,N_7710,N_7711,N_7712,N_7713,N_7714,N_7715,N_7716,N_7717,N_7718,N_7719,N_7720,N_7721,N_7722,N_7723,N_7724,N_7725,N_7726,N_7727,N_7728,N_7729,N_7730,N_7731,N_7732,N_7733,N_7734,N_7735,N_7736,N_7737,N_7738,N_7739,N_7740,N_7741,N_7742,N_7743,N_7744,N_7745,N_7746,N_7747,N_7748,N_7749,N_7750,N_7751,N_7752,N_7753,N_7754,N_7755,N_7756,N_7757,N_7758,N_7759,N_7760,N_7761,N_7762,N_7763,N_7764,N_7765,N_7766,N_7767,N_7768,N_7769,N_7770,N_7771,N_7772,N_7773,N_7774,N_7775,N_7776,N_7777,N_7778,N_7779,N_7780,N_7781,N_7782,N_7783,N_7784,N_7785,N_7786,N_7787,N_7788,N_7789,N_7790,N_7791,N_7792,N_7793,N_7794,N_7795,N_7796,N_7797,N_7798,N_7799,N_7800,N_7801,N_7802,N_7803,N_7804,N_7805,N_7806,N_7807,N_7808,N_7809,N_7810,N_7811,N_7812,N_7813,N_7814,N_7815,N_7816,N_7817,N_7818,N_7819,N_7820,N_7821,N_7822,N_7823,N_7824,N_7825,N_7826,N_7827,N_7828,N_7829,N_7830,N_7831,N_7832,N_7833,N_7834,N_7835,N_7836,N_7837,N_7838,N_7839,N_7840,N_7841,N_7842,N_7843,N_7844,N_7845,N_7846,N_7847,N_7848,N_7849,N_7850,N_7851,N_7852,N_7853,N_7854,N_7855,N_7856,N_7857,N_7858,N_7859,N_7860,N_7861,N_7862,N_7863,N_7864,N_7865,N_7866,N_7867,N_7868,N_7869,N_7870,N_7871,N_7872,N_7873,N_7874,N_7875,N_7876,N_7877,N_7878,N_7879,N_7880,N_7881,N_7882,N_7883,N_7884,N_7885,N_7886,N_7887,N_7888,N_7889,N_7890,N_7891,N_7892,N_7893,N_7894,N_7895,N_7896,N_7897,N_7898,N_7899,N_7900,N_7901,N_7902,N_7903,N_7904,N_7905,N_7906,N_7907,N_7908,N_7909,N_7910,N_7911,N_7912,N_7913,N_7914,N_7915,N_7916,N_7917,N_7918,N_7919,N_7920,N_7921,N_7922,N_7923,N_7924,N_7925,N_7926,N_7927,N_7928,N_7929,N_7930,N_7931,N_7932,N_7933,N_7934,N_7935,N_7936,N_7937,N_7938,N_7939,N_7940,N_7941,N_7942,N_7943,N_7944,N_7945,N_7946,N_7947,N_7948,N_7949,N_7950,N_7951,N_7952,N_7953,N_7954,N_7955,N_7956,N_7957,N_7958,N_7959,N_7960,N_7961,N_7962,N_7963,N_7964,N_7965,N_7966,N_7967,N_7968,N_7969,N_7970,N_7971,N_7972,N_7973,N_7974,N_7975,N_7976,N_7977,N_7978,N_7979,N_7980,N_7981,N_7982,N_7983,N_7984,N_7985,N_7986,N_7987,N_7988,N_7989,N_7990,N_7991,N_7992,N_7993,N_7994,N_7995,N_7996,N_7997,N_7998,N_7999,N_8000,N_8001,N_8002,N_8003,N_8004,N_8005,N_8006,N_8007,N_8008,N_8009,N_8010,N_8011,N_8012,N_8013,N_8014,N_8015,N_8016,N_8017,N_8018,N_8019,N_8020,N_8021,N_8022,N_8023,N_8024,N_8025,N_8026,N_8027,N_8028,N_8029,N_8030,N_8031,N_8032,N_8033,N_8034,N_8035,N_8036,N_8037,N_8038,N_8039,N_8040,N_8041,N_8042,N_8043,N_8044,N_8045,N_8046,N_8047,N_8048,N_8049,N_8050,N_8051,N_8052,N_8053,N_8054,N_8055,N_8056,N_8057,N_8058,N_8059,N_8060,N_8061,N_8062,N_8063,N_8064,N_8065,N_8066,N_8067,N_8068,N_8069,N_8070,N_8071,N_8072,N_8073,N_8074,N_8075,N_8076,N_8077,N_8078,N_8079,N_8080,N_8081,N_8082,N_8083,N_8084,N_8085,N_8086,N_8087,N_8088,N_8089,N_8090,N_8091,N_8092,N_8093,N_8094,N_8095,N_8096,N_8097,N_8098,N_8099,N_8100,N_8101,N_8102,N_8103,N_8104,N_8105,N_8106,N_8107,N_8108,N_8109,N_8110,N_8111,N_8112,N_8113,N_8114,N_8115,N_8116,N_8117,N_8118,N_8119,N_8120,N_8121,N_8122,N_8123,N_8124,N_8125,N_8126,N_8127,N_8128,N_8129,N_8130,N_8131,N_8132,N_8133,N_8134,N_8135,N_8136,N_8137,N_8138,N_8139,N_8140,N_8141,N_8142,N_8143,N_8144,N_8145,N_8146,N_8147,N_8148,N_8149,N_8150,N_8151,N_8152,N_8153,N_8154,N_8155,N_8156,N_8157,N_8158,N_8159,N_8160,N_8161,N_8162,N_8163,N_8164,N_8165,N_8166,N_8167,N_8168,N_8169,N_8170,N_8171,N_8172,N_8173,N_8174,N_8175,N_8176,N_8177,N_8178,N_8179,N_8180,N_8181,N_8182,N_8183,N_8184,N_8185,N_8186,N_8187,N_8188,N_8189,N_8190,N_8191,N_8192,N_8193,N_8194,N_8195,N_8196,N_8197,N_8198,N_8199,N_8200,N_8201,N_8202,N_8203,N_8204,N_8205,N_8206,N_8207,N_8208,N_8209,N_8210,N_8211,N_8212,N_8213,N_8214,N_8215,N_8216,N_8217,N_8218,N_8219,N_8220,N_8221,N_8222,N_8223,N_8224,N_8225,N_8226,N_8227,N_8228,N_8229,N_8230,N_8231,N_8232,N_8233,N_8234,N_8235,N_8236,N_8237,N_8238,N_8239,N_8240,N_8241,N_8242,N_8243,N_8244,N_8245,N_8246,N_8247,N_8248,N_8249,N_8250,N_8251,N_8252,N_8253,N_8254,N_8255,N_8256,N_8257,N_8258,N_8259,N_8260,N_8261,N_8262,N_8263,N_8264,N_8265,N_8266,N_8267,N_8268,N_8269,N_8270,N_8271,N_8272,N_8273,N_8274,N_8275,N_8276,N_8277,N_8278,N_8279,N_8280,N_8281,N_8282,N_8283,N_8284,N_8285,N_8286,N_8287,N_8288,N_8289,N_8290,N_8291,N_8292,N_8293,N_8294,N_8295,N_8296,N_8297,N_8298,N_8299,N_8300,N_8301,N_8302,N_8303,N_8304,N_8305,N_8306,N_8307,N_8308,N_8309,N_8310,N_8311,N_8312,N_8313,N_8314,N_8315,N_8316,N_8317,N_8318,N_8319,N_8320,N_8321,N_8322,N_8323,N_8324,N_8325,N_8326,N_8327,N_8328,N_8329,N_8330,N_8331,N_8332,N_8333,N_8334,N_8335,N_8336,N_8337,N_8338,N_8339,N_8340,N_8341,N_8342,N_8343,N_8344,N_8345,N_8346,N_8347,N_8348,N_8349,N_8350,N_8351,N_8352,N_8353,N_8354,N_8355,N_8356,N_8357,N_8358,N_8359,N_8360,N_8361,N_8362,N_8363,N_8364,N_8365,N_8366,N_8367,N_8368,N_8369,N_8370,N_8371,N_8372,N_8373,N_8374,N_8375,N_8376,N_8377,N_8378,N_8379,N_8380,N_8381,N_8382,N_8383,N_8384,N_8385,N_8386,N_8387,N_8388,N_8389,N_8390,N_8391,N_8392,N_8393,N_8394,N_8395,N_8396,N_8397,N_8398,N_8399,N_8400,N_8401,N_8402,N_8403,N_8404,N_8405,N_8406,N_8407,N_8408,N_8409,N_8410,N_8411,N_8412,N_8413,N_8414,N_8415,N_8416,N_8417,N_8418,N_8419,N_8420,N_8421,N_8422,N_8423,N_8424,N_8425,N_8426,N_8427,N_8428,N_8429,N_8430,N_8431,N_8432,N_8433,N_8434,N_8435,N_8436,N_8437,N_8438,N_8439,N_8440,N_8441,N_8442,N_8443,N_8444,N_8445,N_8446,N_8447,N_8448,N_8449,N_8450,N_8451,N_8452,N_8453,N_8454,N_8455,N_8456,N_8457,N_8458,N_8459,N_8460,N_8461,N_8462,N_8463,N_8464,N_8465,N_8466,N_8467,N_8468,N_8469,N_8470,N_8471,N_8472,N_8473,N_8474,N_8475,N_8476,N_8477,N_8478,N_8479,N_8480,N_8481,N_8482,N_8483,N_8484,N_8485,N_8486,N_8487,N_8488,N_8489,N_8490,N_8491,N_8492,N_8493,N_8494,N_8495,N_8496,N_8497,N_8498,N_8499,N_8500,N_8501,N_8502,N_8503,N_8504,N_8505,N_8506,N_8507,N_8508,N_8509,N_8510,N_8511,N_8512,N_8513,N_8514,N_8515,N_8516,N_8517,N_8518,N_8519,N_8520,N_8521,N_8522,N_8523,N_8524,N_8525,N_8526,N_8527,N_8528,N_8529,N_8530,N_8531,N_8532,N_8533,N_8534,N_8535,N_8536,N_8537,N_8538,N_8539,N_8540,N_8541,N_8542,N_8543,N_8544,N_8545,N_8546,N_8547,N_8548,N_8549,N_8550,N_8551,N_8552,N_8553,N_8554,N_8555,N_8556,N_8557,N_8558,N_8559,N_8560,N_8561,N_8562,N_8563,N_8564,N_8565,N_8566,N_8567,N_8568,N_8569,N_8570,N_8571,N_8572,N_8573,N_8574,N_8575,N_8576,N_8577,N_8578,N_8579,N_8580,N_8581,N_8582,N_8583,N_8584,N_8585,N_8586,N_8587,N_8588,N_8589,N_8590,N_8591,N_8592,N_8593,N_8594,N_8595,N_8596,N_8597,N_8598,N_8599,N_8600,N_8601,N_8602,N_8603,N_8604,N_8605,N_8606,N_8607,N_8608,N_8609,N_8610,N_8611,N_8612,N_8613,N_8614,N_8615,N_8616,N_8617,N_8618,N_8619,N_8620,N_8621,N_8622,N_8623,N_8624,N_8625,N_8626,N_8627,N_8628,N_8629,N_8630,N_8631,N_8632,N_8633,N_8634,N_8635,N_8636,N_8637,N_8638,N_8639,N_8640,N_8641,N_8642,N_8643,N_8644,N_8645,N_8646,N_8647,N_8648,N_8649,N_8650,N_8651,N_8652,N_8653,N_8654,N_8655,N_8656,N_8657,N_8658,N_8659,N_8660,N_8661,N_8662,N_8663,N_8664,N_8665,N_8666,N_8667,N_8668,N_8669,N_8670,N_8671,N_8672,N_8673,N_8674,N_8675,N_8676,N_8677,N_8678,N_8679,N_8680,N_8681,N_8682,N_8683,N_8684,N_8685,N_8686,N_8687,N_8688,N_8689,N_8690,N_8691,N_8692,N_8693,N_8694,N_8695,N_8696,N_8697,N_8698,N_8699,N_8700,N_8701,N_8702,N_8703,N_8704,N_8705,N_8706,N_8707,N_8708,N_8709,N_8710,N_8711,N_8712,N_8713,N_8714,N_8715,N_8716,N_8717,N_8718,N_8719,N_8720,N_8721,N_8722,N_8723,N_8724,N_8725,N_8726,N_8727,N_8728,N_8729,N_8730,N_8731,N_8732,N_8733,N_8734,N_8735,N_8736,N_8737,N_8738,N_8739,N_8740,N_8741,N_8742,N_8743,N_8744,N_8745,N_8746,N_8747,N_8748,N_8749,N_8750,N_8751,N_8752,N_8753,N_8754,N_8755,N_8756,N_8757,N_8758,N_8759,N_8760,N_8761,N_8762,N_8763,N_8764,N_8765,N_8766,N_8767,N_8768,N_8769,N_8770,N_8771,N_8772,N_8773,N_8774,N_8775,N_8776,N_8777,N_8778,N_8779,N_8780,N_8781,N_8782,N_8783,N_8784,N_8785,N_8786,N_8787,N_8788,N_8789,N_8790,N_8791,N_8792,N_8793,N_8794,N_8795,N_8796,N_8797,N_8798,N_8799,N_8800,N_8801,N_8802,N_8803,N_8804,N_8805,N_8806,N_8807,N_8808,N_8809,N_8810,N_8811,N_8812,N_8813,N_8814,N_8815,N_8816,N_8817,N_8818,N_8819,N_8820,N_8821,N_8822,N_8823,N_8824,N_8825,N_8826,N_8827,N_8828,N_8829,N_8830,N_8831,N_8832,N_8833,N_8834,N_8835,N_8836,N_8837,N_8838,N_8839,N_8840,N_8841,N_8842,N_8843,N_8844,N_8845,N_8846,N_8847,N_8848,N_8849,N_8850,N_8851,N_8852,N_8853,N_8854,N_8855,N_8856,N_8857,N_8858,N_8859,N_8860,N_8861,N_8862,N_8863,N_8864,N_8865,N_8866,N_8867,N_8868,N_8869,N_8870,N_8871,N_8872,N_8873,N_8874,N_8875,N_8876,N_8877,N_8878,N_8879,N_8880,N_8881,N_8882,N_8883,N_8884,N_8885,N_8886,N_8887,N_8888,N_8889,N_8890,N_8891,N_8892,N_8893,N_8894,N_8895,N_8896,N_8897,N_8898,N_8899,N_8900,N_8901,N_8902,N_8903,N_8904,N_8905,N_8906,N_8907,N_8908,N_8909,N_8910,N_8911,N_8912,N_8913,N_8914,N_8915,N_8916,N_8917,N_8918,N_8919,N_8920,N_8921,N_8922,N_8923,N_8924,N_8925,N_8926,N_8927,N_8928,N_8929,N_8930,N_8931,N_8932,N_8933,N_8934,N_8935,N_8936,N_8937,N_8938,N_8939,N_8940,N_8941,N_8942,N_8943,N_8944,N_8945,N_8946,N_8947,N_8948,N_8949,N_8950,N_8951,N_8952,N_8953,N_8954,N_8955,N_8956,N_8957,N_8958,N_8959,N_8960,N_8961,N_8962,N_8963,N_8964,N_8965,N_8966,N_8967,N_8968,N_8969,N_8970,N_8971,N_8972,N_8973,N_8974,N_8975,N_8976,N_8977,N_8978,N_8979,N_8980,N_8981,N_8982,N_8983,N_8984,N_8985,N_8986,N_8987,N_8988,N_8989,N_8990,N_8991,N_8992,N_8993,N_8994,N_8995,N_8996,N_8997,N_8998,N_8999,N_9000,N_9001,N_9002,N_9003,N_9004,N_9005,N_9006,N_9007,N_9008,N_9009,N_9010,N_9011,N_9012,N_9013,N_9014,N_9015,N_9016,N_9017,N_9018,N_9019,N_9020,N_9021,N_9022,N_9023,N_9024,N_9025,N_9026,N_9027,N_9028,N_9029,N_9030,N_9031,N_9032,N_9033,N_9034,N_9035,N_9036,N_9037,N_9038,N_9039,N_9040,N_9041,N_9042,N_9043,N_9044,N_9045,N_9046,N_9047,N_9048,N_9049,N_9050,N_9051,N_9052,N_9053,N_9054,N_9055,N_9056,N_9057,N_9058,N_9059,N_9060,N_9061,N_9062,N_9063,N_9064,N_9065,N_9066,N_9067,N_9068,N_9069,N_9070,N_9071,N_9072,N_9073,N_9074,N_9075,N_9076,N_9077,N_9078,N_9079,N_9080,N_9081,N_9082,N_9083,N_9084,N_9085,N_9086,N_9087,N_9088,N_9089,N_9090,N_9091,N_9092,N_9093,N_9094,N_9095,N_9096,N_9097,N_9098,N_9099,N_9100,N_9101,N_9102,N_9103,N_9104,N_9105,N_9106,N_9107,N_9108,N_9109,N_9110,N_9111,N_9112,N_9113,N_9114,N_9115,N_9116,N_9117,N_9118,N_9119,N_9120,N_9121,N_9122,N_9123,N_9124,N_9125,N_9126,N_9127,N_9128,N_9129,N_9130,N_9131,N_9132,N_9133,N_9134,N_9135,N_9136,N_9137,N_9138,N_9139,N_9140,N_9141,N_9142,N_9143,N_9144,N_9145,N_9146,N_9147,N_9148,N_9149,N_9150,N_9151,N_9152,N_9153,N_9154,N_9155,N_9156,N_9157,N_9158,N_9159,N_9160,N_9161,N_9162,N_9163,N_9164,N_9165,N_9166,N_9167,N_9168,N_9169,N_9170,N_9171,N_9172,N_9173,N_9174,N_9175,N_9176,N_9177,N_9178,N_9179,N_9180,N_9181,N_9182,N_9183,N_9184,N_9185,N_9186,N_9187,N_9188,N_9189,N_9190,N_9191,N_9192,N_9193,N_9194,N_9195,N_9196,N_9197,N_9198,N_9199,N_9200,N_9201,N_9202,N_9203,N_9204,N_9205,N_9206,N_9207,N_9208,N_9209,N_9210,N_9211,N_9212,N_9213,N_9214,N_9215,N_9216,N_9217,N_9218,N_9219,N_9220,N_9221,N_9222,N_9223,N_9224,N_9225,N_9226,N_9227,N_9228,N_9229,N_9230,N_9231,N_9232,N_9233,N_9234,N_9235,N_9236,N_9237,N_9238,N_9239,N_9240,N_9241,N_9242,N_9243,N_9244,N_9245,N_9246,N_9247,N_9248,N_9249,N_9250,N_9251,N_9252,N_9253,N_9254,N_9255,N_9256,N_9257,N_9258,N_9259,N_9260,N_9261,N_9262,N_9263,N_9264,N_9265,N_9266,N_9267,N_9268,N_9269,N_9270,N_9271,N_9272,N_9273,N_9274,N_9275,N_9276,N_9277,N_9278,N_9279,N_9280,N_9281,N_9282,N_9283,N_9284,N_9285,N_9286,N_9287,N_9288,N_9289,N_9290,N_9291,N_9292,N_9293,N_9294,N_9295,N_9296,N_9297,N_9298,N_9299,N_9300,N_9301,N_9302,N_9303,N_9304,N_9305,N_9306,N_9307,N_9308,N_9309,N_9310,N_9311,N_9312,N_9313,N_9314,N_9315,N_9316,N_9317,N_9318,N_9319,N_9320,N_9321,N_9322,N_9323,N_9324,N_9325,N_9326,N_9327,N_9328,N_9329,N_9330,N_9331,N_9332,N_9333,N_9334,N_9335,N_9336,N_9337,N_9338,N_9339,N_9340,N_9341,N_9342,N_9343,N_9344,N_9345,N_9346,N_9347,N_9348,N_9349,N_9350,N_9351,N_9352,N_9353,N_9354,N_9355,N_9356,N_9357,N_9358,N_9359,N_9360,N_9361,N_9362,N_9363,N_9364,N_9365,N_9366,N_9367,N_9368,N_9369,N_9370,N_9371,N_9372,N_9373,N_9374,N_9375,N_9376,N_9377,N_9378,N_9379,N_9380,N_9381,N_9382,N_9383,N_9384,N_9385,N_9386,N_9387,N_9388,N_9389,N_9390,N_9391,N_9392,N_9393,N_9394,N_9395,N_9396,N_9397,N_9398,N_9399,N_9400,N_9401,N_9402,N_9403,N_9404,N_9405,N_9406,N_9407,N_9408,N_9409,N_9410,N_9411,N_9412,N_9413,N_9414,N_9415,N_9416,N_9417,N_9418,N_9419,N_9420,N_9421,N_9422,N_9423,N_9424,N_9425,N_9426,N_9427,N_9428,N_9429,N_9430,N_9431,N_9432,N_9433,N_9434,N_9435,N_9436,N_9437,N_9438,N_9439,N_9440,N_9441,N_9442,N_9443,N_9444,N_9445,N_9446,N_9447,N_9448,N_9449,N_9450,N_9451,N_9452,N_9453,N_9454,N_9455,N_9456,N_9457,N_9458,N_9459,N_9460,N_9461,N_9462,N_9463,N_9464,N_9465,N_9466,N_9467,N_9468,N_9469,N_9470,N_9471,N_9472,N_9473,N_9474,N_9475,N_9476,N_9477,N_9478,N_9479,N_9480,N_9481,N_9482,N_9483,N_9484,N_9485,N_9486,N_9487,N_9488,N_9489,N_9490,N_9491,N_9492,N_9493,N_9494,N_9495,N_9496,N_9497,N_9498,N_9499,N_9500,N_9501,N_9502,N_9503,N_9504,N_9505,N_9506,N_9507,N_9508,N_9509,N_9510,N_9511,N_9512,N_9513,N_9514,N_9515,N_9516,N_9517,N_9518,N_9519,N_9520,N_9521,N_9522,N_9523,N_9524,N_9525,N_9526,N_9527,N_9528,N_9529,N_9530,N_9531,N_9532,N_9533,N_9534,N_9535,N_9536,N_9537,N_9538,N_9539,N_9540,N_9541,N_9542,N_9543,N_9544,N_9545,N_9546,N_9547,N_9548,N_9549,N_9550,N_9551,N_9552,N_9553,N_9554,N_9555,N_9556,N_9557,N_9558,N_9559,N_9560,N_9561,N_9562,N_9563,N_9564,N_9565,N_9566,N_9567,N_9568,N_9569,N_9570,N_9571,N_9572,N_9573,N_9574,N_9575,N_9576,N_9577,N_9578,N_9579,N_9580,N_9581,N_9582,N_9583,N_9584,N_9585,N_9586,N_9587,N_9588,N_9589,N_9590,N_9591,N_9592,N_9593,N_9594,N_9595,N_9596,N_9597,N_9598,N_9599,N_9600,N_9601,N_9602,N_9603,N_9604,N_9605,N_9606,N_9607,N_9608,N_9609,N_9610,N_9611,N_9612,N_9613,N_9614,N_9615,N_9616,N_9617,N_9618,N_9619,N_9620,N_9621,N_9622,N_9623,N_9624,N_9625,N_9626,N_9627,N_9628,N_9629,N_9630,N_9631,N_9632,N_9633,N_9634,N_9635,N_9636,N_9637,N_9638,N_9639,N_9640,N_9641,N_9642,N_9643,N_9644,N_9645,N_9646,N_9647,N_9648,N_9649,N_9650,N_9651,N_9652,N_9653,N_9654,N_9655,N_9656,N_9657,N_9658,N_9659,N_9660,N_9661,N_9662,N_9663,N_9664,N_9665,N_9666,N_9667,N_9668,N_9669,N_9670,N_9671,N_9672,N_9673,N_9674,N_9675,N_9676,N_9677,N_9678,N_9679,N_9680,N_9681,N_9682,N_9683,N_9684,N_9685,N_9686,N_9687,N_9688,N_9689,N_9690,N_9691,N_9692,N_9693,N_9694,N_9695,N_9696,N_9697,N_9698,N_9699,N_9700,N_9701,N_9702,N_9703,N_9704,N_9705,N_9706,N_9707,N_9708,N_9709,N_9710,N_9711,N_9712,N_9713,N_9714,N_9715,N_9716,N_9717,N_9718,N_9719,N_9720,N_9721,N_9722,N_9723,N_9724,N_9725,N_9726,N_9727,N_9728,N_9729,N_9730,N_9731,N_9732,N_9733,N_9734,N_9735,N_9736,N_9737,N_9738,N_9739,N_9740,N_9741,N_9742,N_9743,N_9744,N_9745,N_9746,N_9747,N_9748,N_9749,N_9750,N_9751,N_9752,N_9753,N_9754,N_9755,N_9756,N_9757,N_9758,N_9759,N_9760,N_9761,N_9762,N_9763,N_9764,N_9765,N_9766,N_9767,N_9768,N_9769,N_9770,N_9771,N_9772,N_9773,N_9774,N_9775,N_9776,N_9777,N_9778,N_9779,N_9780,N_9781,N_9782,N_9783,N_9784,N_9785,N_9786,N_9787,N_9788,N_9789,N_9790,N_9791,N_9792,N_9793,N_9794,N_9795,N_9796,N_9797,N_9798,N_9799,N_9800,N_9801,N_9802,N_9803,N_9804,N_9805,N_9806,N_9807,N_9808,N_9809,N_9810,N_9811,N_9812,N_9813,N_9814,N_9815,N_9816,N_9817,N_9818,N_9819,N_9820,N_9821,N_9822,N_9823,N_9824,N_9825,N_9826,N_9827,N_9828,N_9829,N_9830,N_9831,N_9832,N_9833,N_9834,N_9835,N_9836,N_9837,N_9838,N_9839,N_9840,N_9841,N_9842,N_9843,N_9844,N_9845,N_9846,N_9847,N_9848,N_9849,N_9850,N_9851,N_9852,N_9853,N_9854,N_9855,N_9856,N_9857,N_9858,N_9859,N_9860,N_9861,N_9862,N_9863,N_9864,N_9865,N_9866,N_9867,N_9868,N_9869,N_9870,N_9871,N_9872,N_9873,N_9874,N_9875,N_9876,N_9877,N_9878,N_9879,N_9880,N_9881,N_9882,N_9883,N_9884,N_9885,N_9886,N_9887,N_9888,N_9889,N_9890,N_9891,N_9892,N_9893,N_9894,N_9895,N_9896,N_9897,N_9898,N_9899,N_9900,N_9901,N_9902,N_9903,N_9904,N_9905,N_9906,N_9907,N_9908,N_9909,N_9910,N_9911,N_9912,N_9913,N_9914,N_9915,N_9916,N_9917,N_9918,N_9919,N_9920,N_9921,N_9922,N_9923,N_9924,N_9925,N_9926,N_9927,N_9928,N_9929,N_9930,N_9931,N_9932,N_9933,N_9934,N_9935,N_9936,N_9937,N_9938,N_9939,N_9940,N_9941,N_9942,N_9943,N_9944,N_9945,N_9946,N_9947,N_9948,N_9949,N_9950,N_9951,N_9952,N_9953,N_9954,N_9955,N_9956,N_9957,N_9958,N_9959,N_9960,N_9961,N_9962,N_9963,N_9964,N_9965,N_9966,N_9967,N_9968,N_9969,N_9970,N_9971,N_9972,N_9973,N_9974,N_9975,N_9976,N_9977,N_9978,N_9979,N_9980,N_9981,N_9982,N_9983,N_9984,N_9985,N_9986,N_9987,N_9988,N_9989,N_9990,N_9991,N_9992,N_9993,N_9994,N_9995,N_9996,N_9997,N_9998,N_9999,N_10000,N_10001,N_10002,N_10003,N_10004,N_10005,N_10006,N_10007,N_10008,N_10009,N_10010,N_10011,N_10012,N_10013,N_10014,N_10015,N_10016,N_10017,N_10018,N_10019,N_10020,N_10021,N_10022,N_10023,N_10024,N_10025,N_10026,N_10027,N_10028,N_10029,N_10030,N_10031,N_10032,N_10033,N_10034,N_10035,N_10036,N_10037,N_10038,N_10039,N_10040,N_10041,N_10042,N_10043,N_10044,N_10045,N_10046,N_10047,N_10048,N_10049,N_10050,N_10051,N_10052,N_10053,N_10054,N_10055,N_10056,N_10057,N_10058,N_10059,N_10060,N_10061,N_10062,N_10063,N_10064,N_10065,N_10066,N_10067,N_10068,N_10069,N_10070,N_10071,N_10072,N_10073,N_10074,N_10075,N_10076,N_10077,N_10078,N_10079,N_10080,N_10081,N_10082,N_10083,N_10084,N_10085,N_10086,N_10087,N_10088,N_10089,N_10090,N_10091,N_10092,N_10093,N_10094,N_10095,N_10096,N_10097,N_10098,N_10099,N_10100,N_10101,N_10102,N_10103,N_10104,N_10105,N_10106,N_10107,N_10108,N_10109,N_10110,N_10111,N_10112,N_10113,N_10114,N_10115,N_10116,N_10117,N_10118,N_10119,N_10120,N_10121,N_10122,N_10123,N_10124,N_10125,N_10126,N_10127,N_10128,N_10129,N_10130,N_10131,N_10132,N_10133,N_10134,N_10135,N_10136,N_10137,N_10138,N_10139,N_10140,N_10141,N_10142,N_10143,N_10144,N_10145,N_10146,N_10147,N_10148,N_10149,N_10150,N_10151,N_10152,N_10153,N_10154,N_10155,N_10156,N_10157,N_10158,N_10159,N_10160,N_10161,N_10162,N_10163,N_10164,N_10165,N_10166,N_10167,N_10168,N_10169,N_10170,N_10171,N_10172,N_10173,N_10174,N_10175,N_10176,N_10177,N_10178,N_10179,N_10180,N_10181,N_10182,N_10183,N_10184,N_10185,N_10186,N_10187,N_10188,N_10189,N_10190,N_10191,N_10192,N_10193,N_10194,N_10195,N_10196,N_10197,N_10198,N_10199,N_10200,N_10201,N_10202,N_10203,N_10204,N_10205,N_10206,N_10207,N_10208,N_10209,N_10210,N_10211,N_10212,N_10213,N_10214,N_10215,N_10216,N_10217,N_10218,N_10219,N_10220,N_10221,N_10222,N_10223,N_10224,N_10225,N_10226,N_10227,N_10228,N_10229,N_10230,N_10231,N_10232,N_10233,N_10234,N_10235,N_10236,N_10237,N_10238,N_10239,N_10240,N_10241,N_10242,N_10243,N_10244,N_10245,N_10246,N_10247,N_10248,N_10249,N_10250,N_10251,N_10252,N_10253,N_10254,N_10255,N_10256,N_10257,N_10258,N_10259,N_10260,N_10261,N_10262,N_10263,N_10264,N_10265,N_10266,N_10267,N_10268,N_10269,N_10270,N_10271,N_10272,N_10273,N_10274,N_10275,N_10276,N_10277,N_10278,N_10279,N_10280,N_10281,N_10282,N_10283,N_10284,N_10285,N_10286,N_10287,N_10288,N_10289,N_10290,N_10291,N_10292,N_10293,N_10294,N_10295,N_10296,N_10297,N_10298,N_10299,N_10300,N_10301,N_10302,N_10303,N_10304,N_10305,N_10306,N_10307,N_10308,N_10309,N_10310,N_10311,N_10312,N_10313,N_10314,N_10315,N_10316,N_10317,N_10318,N_10319,N_10320,N_10321,N_10322,N_10323,N_10324,N_10325,N_10326,N_10327,N_10328,N_10329,N_10330,N_10331,N_10332,N_10333,N_10334,N_10335,N_10336,N_10337,N_10338,N_10339,N_10340,N_10341,N_10342,N_10343,N_10344,N_10345,N_10346,N_10347,N_10348,N_10349,N_10350,N_10351,N_10352,N_10353,N_10354,N_10355,N_10356,N_10357,N_10358,N_10359,N_10360,N_10361,N_10362,N_10363,N_10364,N_10365,N_10366,N_10367,N_10368,N_10369,N_10370,N_10371,N_10372,N_10373,N_10374,N_10375,N_10376,N_10377,N_10378,N_10379,N_10380,N_10381,N_10382,N_10383,N_10384,N_10385,N_10386,N_10387,N_10388,N_10389,N_10390,N_10391,N_10392,N_10393,N_10394,N_10395,N_10396,N_10397,N_10398,N_10399,N_10400,N_10401,N_10402,N_10403,N_10404,N_10405,N_10406,N_10407,N_10408,N_10409,N_10410,N_10411,N_10412,N_10413,N_10414,N_10415,N_10416,N_10417,N_10418,N_10419,N_10420,N_10421,N_10422,N_10423,N_10424,N_10425,N_10426,N_10427,N_10428,N_10429,N_10430,N_10431,N_10432,N_10433,N_10434,N_10435,N_10436,N_10437,N_10438,N_10439,N_10440,N_10441,N_10442,N_10443,N_10444,N_10445,N_10446,N_10447,N_10448,N_10449,N_10450,N_10451,N_10452,N_10453,N_10454,N_10455,N_10456,N_10457,N_10458,N_10459,N_10460,N_10461,N_10462,N_10463,N_10464,N_10465,N_10466,N_10467,N_10468,N_10469,N_10470,N_10471,N_10472,N_10473,N_10474,N_10475,N_10476,N_10477,N_10478,N_10479,N_10480,N_10481,N_10482,N_10483,N_10484,N_10485,N_10486,N_10487,N_10488,N_10489,N_10490,N_10491,N_10492,N_10493,N_10494,N_10495,N_10496,N_10497,N_10498,N_10499,N_10500,N_10501,N_10502,N_10503,N_10504,N_10505,N_10506,N_10507,N_10508,N_10509,N_10510,N_10511,N_10512,N_10513,N_10514,N_10515,N_10516,N_10517,N_10518,N_10519,N_10520,N_10521,N_10522,N_10523,N_10524,N_10525,N_10526,N_10527,N_10528,N_10529,N_10530,N_10531,N_10532,N_10533,N_10534,N_10535,N_10536,N_10537,N_10538,N_10539,N_10540,N_10541,N_10542,N_10543,N_10544,N_10545,N_10546,N_10547,N_10548,N_10549,N_10550,N_10551,N_10552,N_10553,N_10554,N_10555,N_10556,N_10557,N_10558,N_10559,N_10560,N_10561,N_10562,N_10563,N_10564,N_10565,N_10566,N_10567,N_10568,N_10569,N_10570,N_10571,N_10572,N_10573,N_10574,N_10575,N_10576,N_10577,N_10578,N_10579,N_10580,N_10581,N_10582,N_10583,N_10584,N_10585,N_10586,N_10587,N_10588,N_10589,N_10590,N_10591,N_10592,N_10593,N_10594,N_10595,N_10596,N_10597,N_10598,N_10599,N_10600,N_10601,N_10602,N_10603,N_10604,N_10605,N_10606,N_10607,N_10608,N_10609,N_10610,N_10611,N_10612,N_10613,N_10614,N_10615,N_10616,N_10617,N_10618,N_10619,N_10620,N_10621,N_10622,N_10623,N_10624,N_10625,N_10626,N_10627,N_10628,N_10629,N_10630,N_10631,N_10632,N_10633,N_10634,N_10635,N_10636,N_10637,N_10638,N_10639,N_10640,N_10641,N_10642,N_10643,N_10644,N_10645,N_10646,N_10647,N_10648,N_10649,N_10650,N_10651,N_10652,N_10653,N_10654,N_10655,N_10656,N_10657,N_10658,N_10659,N_10660,N_10661,N_10662,N_10663,N_10664,N_10665,N_10666,N_10667,N_10668,N_10669,N_10670,N_10671,N_10672,N_10673,N_10674,N_10675,N_10676,N_10677,N_10678,N_10679,N_10680,N_10681,N_10682,N_10683,N_10684,N_10685,N_10686,N_10687,N_10688,N_10689,N_10690,N_10691,N_10692,N_10693,N_10694,N_10695,N_10696,N_10697,N_10698,N_10699,N_10700,N_10701,N_10702,N_10703,N_10704,N_10705,N_10706,N_10707,N_10708,N_10709,N_10710,N_10711,N_10712,N_10713,N_10714,N_10715,N_10716,N_10717,N_10718,N_10719,N_10720,N_10721,N_10722,N_10723,N_10724,N_10725,N_10726,N_10727,N_10728,N_10729,N_10730,N_10731,N_10732,N_10733,N_10734,N_10735,N_10736,N_10737,N_10738,N_10739,N_10740,N_10741,N_10742,N_10743,N_10744,N_10745,N_10746,N_10747,N_10748,N_10749,N_10750,N_10751,N_10752,N_10753,N_10754,N_10755,N_10756,N_10757,N_10758,N_10759,N_10760,N_10761,N_10762,N_10763,N_10764,N_10765,N_10766,N_10767,N_10768,N_10769,N_10770,N_10771,N_10772,N_10773,N_10774,N_10775,N_10776,N_10777,N_10778,N_10779,N_10780,N_10781,N_10782,N_10783,N_10784,N_10785,N_10786,N_10787,N_10788,N_10789,N_10790,N_10791,N_10792,N_10793,N_10794,N_10795,N_10796,N_10797,N_10798,N_10799,N_10800,N_10801,N_10802,N_10803,N_10804,N_10805,N_10806,N_10807,N_10808,N_10809,N_10810,N_10811,N_10812,N_10813,N_10814,N_10815,N_10816,N_10817,N_10818,N_10819,N_10820,N_10821,N_10822,N_10823,N_10824,N_10825,N_10826,N_10827,N_10828,N_10829,N_10830,N_10831,N_10832,N_10833,N_10834,N_10835,N_10836,N_10837,N_10838,N_10839,N_10840,N_10841,N_10842,N_10843,N_10844,N_10845,N_10846,N_10847,N_10848,N_10849,N_10850,N_10851,N_10852,N_10853,N_10854,N_10855,N_10856,N_10857,N_10858,N_10859,N_10860,N_10861,N_10862,N_10863,N_10864,N_10865,N_10866,N_10867,N_10868,N_10869,N_10870,N_10871,N_10872,N_10873,N_10874,N_10875,N_10876,N_10877,N_10878,N_10879,N_10880,N_10881,N_10882,N_10883,N_10884,N_10885,N_10886,N_10887,N_10888,N_10889,N_10890,N_10891,N_10892,N_10893,N_10894,N_10895,N_10896,N_10897,N_10898,N_10899,N_10900,N_10901,N_10902,N_10903,N_10904,N_10905,N_10906,N_10907,N_10908,N_10909,N_10910,N_10911,N_10912,N_10913,N_10914,N_10915,N_10916,N_10917,N_10918,N_10919,N_10920,N_10921,N_10922,N_10923,N_10924,N_10925,N_10926,N_10927,N_10928,N_10929,N_10930,N_10931,N_10932,N_10933,N_10934,N_10935,N_10936,N_10937,N_10938,N_10939,N_10940,N_10941,N_10942,N_10943,N_10944,N_10945,N_10946,N_10947,N_10948,N_10949,N_10950,N_10951,N_10952,N_10953,N_10954,N_10955,N_10956,N_10957,N_10958,N_10959,N_10960,N_10961,N_10962,N_10963,N_10964,N_10965,N_10966,N_10967,N_10968,N_10969,N_10970,N_10971,N_10972,N_10973,N_10974,N_10975,N_10976,N_10977,N_10978,N_10979,N_10980,N_10981,N_10982,N_10983,N_10984,N_10985,N_10986,N_10987,N_10988,N_10989,N_10990,N_10991,N_10992,N_10993,N_10994,N_10995,N_10996,N_10997,N_10998,N_10999,N_11000,N_11001,N_11002,N_11003,N_11004,N_11005,N_11006,N_11007,N_11008,N_11009,N_11010,N_11011,N_11012,N_11013,N_11014,N_11015,N_11016,N_11017,N_11018,N_11019,N_11020,N_11021,N_11022,N_11023,N_11024,N_11025,N_11026,N_11027,N_11028,N_11029,N_11030,N_11031,N_11032,N_11033,N_11034,N_11035,N_11036,N_11037,N_11038,N_11039,N_11040,N_11041,N_11042,N_11043,N_11044,N_11045,N_11046,N_11047,N_11048,N_11049,N_11050,N_11051,N_11052,N_11053,N_11054,N_11055,N_11056,N_11057,N_11058,N_11059,N_11060,N_11061,N_11062,N_11063,N_11064,N_11065,N_11066,N_11067,N_11068,N_11069,N_11070,N_11071,N_11072,N_11073,N_11074,N_11075,N_11076,N_11077,N_11078,N_11079,N_11080,N_11081,N_11082,N_11083,N_11084,N_11085,N_11086,N_11087,N_11088,N_11089,N_11090,N_11091,N_11092,N_11093,N_11094,N_11095,N_11096,N_11097,N_11098,N_11099,N_11100,N_11101,N_11102,N_11103,N_11104,N_11105,N_11106,N_11107,N_11108,N_11109,N_11110,N_11111,N_11112,N_11113,N_11114,N_11115,N_11116,N_11117,N_11118,N_11119,N_11120,N_11121,N_11122,N_11123,N_11124,N_11125,N_11126,N_11127,N_11128,N_11129,N_11130,N_11131,N_11132,N_11133,N_11134,N_11135,N_11136,N_11137,N_11138,N_11139,N_11140,N_11141,N_11142,N_11143,N_11144,N_11145,N_11146,N_11147,N_11148,N_11149,N_11150,N_11151,N_11152,N_11153,N_11154,N_11155,N_11156,N_11157,N_11158,N_11159,N_11160,N_11161,N_11162,N_11163,N_11164,N_11165,N_11166,N_11167,N_11168,N_11169,N_11170,N_11171,N_11172,N_11173,N_11174,N_11175,N_11176,N_11177,N_11178,N_11179,N_11180,N_11181,N_11182,N_11183,N_11184,N_11185,N_11186,N_11187,N_11188,N_11189,N_11190,N_11191,N_11192,N_11193,N_11194,N_11195,N_11196,N_11197,N_11198,N_11199,N_11200,N_11201,N_11202,N_11203,N_11204,N_11205,N_11206,N_11207,N_11208,N_11209,N_11210,N_11211,N_11212,N_11213,N_11214,N_11215,N_11216,N_11217,N_11218,N_11219,N_11220,N_11221,N_11222,N_11223,N_11224,N_11225,N_11226,N_11227,N_11228,N_11229,N_11230,N_11231,N_11232,N_11233,N_11234,N_11235,N_11236,N_11237,N_11238,N_11239,N_11240,N_11241,N_11242,N_11243,N_11244,N_11245,N_11246,N_11247,N_11248,N_11249,N_11250,N_11251,N_11252,N_11253,N_11254,N_11255,N_11256,N_11257,N_11258,N_11259,N_11260,N_11261,N_11262,N_11263,N_11264,N_11265,N_11266,N_11267,N_11268,N_11269,N_11270,N_11271,N_11272,N_11273,N_11274,N_11275,N_11276,N_11277,N_11278,N_11279,N_11280,N_11281,N_11282,N_11283,N_11284,N_11285,N_11286,N_11287,N_11288,N_11289,N_11290,N_11291,N_11292,N_11293,N_11294,N_11295,N_11296,N_11297,N_11298,N_11299,N_11300,N_11301,N_11302,N_11303,N_11304,N_11305,N_11306,N_11307,N_11308,N_11309,N_11310,N_11311,N_11312,N_11313,N_11314,N_11315,N_11316,N_11317,N_11318,N_11319,N_11320,N_11321,N_11322,N_11323,N_11324,N_11325,N_11326,N_11327,N_11328,N_11329,N_11330,N_11331,N_11332,N_11333,N_11334,N_11335,N_11336,N_11337,N_11338,N_11339,N_11340,N_11341,N_11342,N_11343,N_11344,N_11345,N_11346,N_11347,N_11348,N_11349,N_11350,N_11351,N_11352,N_11353,N_11354,N_11355,N_11356,N_11357,N_11358,N_11359,N_11360,N_11361,N_11362,N_11363,N_11364,N_11365,N_11366,N_11367,N_11368,N_11369,N_11370,N_11371,N_11372,N_11373,N_11374,N_11375,N_11376,N_11377,N_11378,N_11379,N_11380,N_11381,N_11382,N_11383,N_11384,N_11385,N_11386,N_11387,N_11388,N_11389,N_11390,N_11391,N_11392,N_11393,N_11394,N_11395,N_11396,N_11397,N_11398,N_11399,N_11400,N_11401,N_11402,N_11403,N_11404,N_11405,N_11406,N_11407,N_11408,N_11409,N_11410,N_11411,N_11412,N_11413,N_11414,N_11415,N_11416,N_11417,N_11418,N_11419,N_11420,N_11421,N_11422,N_11423,N_11424,N_11425,N_11426,N_11427,N_11428,N_11429,N_11430,N_11431,N_11432,N_11433,N_11434,N_11435,N_11436,N_11437,N_11438,N_11439,N_11440,N_11441,N_11442,N_11443,N_11444,N_11445,N_11446,N_11447,N_11448,N_11449,N_11450,N_11451,N_11452,N_11453,N_11454,N_11455,N_11456,N_11457,N_11458,N_11459,N_11460,N_11461,N_11462,N_11463,N_11464,N_11465,N_11466,N_11467,N_11468,N_11469,N_11470,N_11471,N_11472,N_11473,N_11474,N_11475,N_11476,N_11477,N_11478,N_11479,N_11480,N_11481,N_11482,N_11483,N_11484,N_11485,N_11486,N_11487,N_11488,N_11489,N_11490,N_11491,N_11492,N_11493,N_11494,N_11495,N_11496,N_11497,N_11498,N_11499,N_11500,N_11501,N_11502,N_11503,N_11504,N_11505,N_11506,N_11507,N_11508,N_11509,N_11510,N_11511,N_11512,N_11513,N_11514,N_11515,N_11516,N_11517,N_11518,N_11519,N_11520,N_11521,N_11522,N_11523,N_11524,N_11525,N_11526,N_11527,N_11528,N_11529,N_11530,N_11531,N_11532,N_11533,N_11534,N_11535,N_11536,N_11537,N_11538,N_11539,N_11540,N_11541,N_11542,N_11543,N_11544,N_11545,N_11546,N_11547,N_11548,N_11549,N_11550,N_11551,N_11552,N_11553,N_11554,N_11555,N_11556,N_11557,N_11558,N_11559,N_11560,N_11561,N_11562,N_11563,N_11564,N_11565,N_11566,N_11567,N_11568,N_11569,N_11570,N_11571,N_11572,N_11573,N_11574,N_11575,N_11576,N_11577,N_11578,N_11579,N_11580,N_11581,N_11582,N_11583,N_11584,N_11585,N_11586,N_11587,N_11588,N_11589,N_11590,N_11591,N_11592,N_11593,N_11594,N_11595,N_11596,N_11597,N_11598,N_11599,N_11600,N_11601,N_11602,N_11603,N_11604,N_11605,N_11606,N_11607,N_11608,N_11609,N_11610,N_11611,N_11612,N_11613,N_11614,N_11615,N_11616,N_11617,N_11618,N_11619,N_11620,N_11621,N_11622,N_11623,N_11624,N_11625,N_11626,N_11627,N_11628,N_11629,N_11630,N_11631,N_11632,N_11633,N_11634,N_11635,N_11636,N_11637,N_11638,N_11639,N_11640,N_11641,N_11642,N_11643,N_11644,N_11645,N_11646,N_11647,N_11648,N_11649,N_11650,N_11651,N_11652,N_11653,N_11654,N_11655,N_11656,N_11657,N_11658,N_11659,N_11660,N_11661,N_11662,N_11663,N_11664,N_11665,N_11666,N_11667,N_11668,N_11669,N_11670,N_11671,N_11672,N_11673,N_11674,N_11675,N_11676,N_11677,N_11678,N_11679,N_11680,N_11681,N_11682,N_11683,N_11684,N_11685,N_11686,N_11687,N_11688,N_11689,N_11690,N_11691,N_11692,N_11693,N_11694,N_11695,N_11696,N_11697,N_11698,N_11699,N_11700,N_11701,N_11702,N_11703,N_11704,N_11705,N_11706,N_11707,N_11708,N_11709,N_11710,N_11711,N_11712,N_11713,N_11714,N_11715,N_11716,N_11717,N_11718,N_11719,N_11720,N_11721,N_11722,N_11723,N_11724,N_11725,N_11726,N_11727,N_11728,N_11729,N_11730,N_11731,N_11732,N_11733,N_11734,N_11735,N_11736,N_11737,N_11738,N_11739,N_11740,N_11741,N_11742,N_11743,N_11744,N_11745,N_11746,N_11747,N_11748,N_11749,N_11750,N_11751,N_11752,N_11753,N_11754,N_11755,N_11756,N_11757,N_11758,N_11759,N_11760,N_11761,N_11762,N_11763,N_11764,N_11765,N_11766,N_11767,N_11768,N_11769,N_11770,N_11771,N_11772,N_11773,N_11774,N_11775,N_11776,N_11777,N_11778,N_11779,N_11780,N_11781,N_11782,N_11783,N_11784,N_11785,N_11786,N_11787,N_11788,N_11789,N_11790,N_11791,N_11792,N_11793,N_11794,N_11795,N_11796,N_11797,N_11798,N_11799,N_11800,N_11801,N_11802,N_11803,N_11804,N_11805,N_11806,N_11807,N_11808,N_11809,N_11810,N_11811,N_11812,N_11813,N_11814,N_11815,N_11816,N_11817,N_11818,N_11819,N_11820,N_11821,N_11822,N_11823,N_11824,N_11825,N_11826,N_11827,N_11828,N_11829,N_11830,N_11831,N_11832,N_11833,N_11834,N_11835,N_11836,N_11837,N_11838,N_11839,N_11840,N_11841,N_11842,N_11843,N_11844,N_11845,N_11846,N_11847,N_11848,N_11849,N_11850,N_11851,N_11852,N_11853,N_11854,N_11855,N_11856,N_11857,N_11858,N_11859,N_11860,N_11861,N_11862,N_11863,N_11864,N_11865,N_11866,N_11867,N_11868,N_11869,N_11870,N_11871,N_11872,N_11873,N_11874,N_11875,N_11876,N_11877,N_11878,N_11879,N_11880,N_11881,N_11882,N_11883,N_11884,N_11885,N_11886,N_11887,N_11888,N_11889,N_11890,N_11891,N_11892,N_11893,N_11894,N_11895,N_11896,N_11897,N_11898,N_11899,N_11900,N_11901,N_11902,N_11903,N_11904,N_11905,N_11906,N_11907,N_11908,N_11909,N_11910,N_11911,N_11912,N_11913,N_11914,N_11915,N_11916,N_11917,N_11918,N_11919,N_11920,N_11921,N_11922,N_11923,N_11924,N_11925,N_11926,N_11927,N_11928,N_11929,N_11930,N_11931,N_11932,N_11933,N_11934,N_11935,N_11936,N_11937,N_11938,N_11939,N_11940,N_11941,N_11942,N_11943,N_11944,N_11945,N_11946,N_11947,N_11948,N_11949,N_11950,N_11951,N_11952,N_11953,N_11954,N_11955,N_11956,N_11957,N_11958,N_11959,N_11960,N_11961,N_11962,N_11963,N_11964,N_11965,N_11966,N_11967,N_11968,N_11969,N_11970,N_11971,N_11972,N_11973,N_11974,N_11975,N_11976,N_11977,N_11978,N_11979,N_11980,N_11981,N_11982,N_11983,N_11984,N_11985,N_11986,N_11987,N_11988,N_11989,N_11990,N_11991,N_11992,N_11993,N_11994,N_11995,N_11996,N_11997,N_11998,N_11999,N_12000,N_12001,N_12002,N_12003,N_12004,N_12005,N_12006,N_12007,N_12008,N_12009,N_12010,N_12011,N_12012,N_12013,N_12014,N_12015,N_12016,N_12017,N_12018,N_12019,N_12020,N_12021,N_12022,N_12023,N_12024,N_12025,N_12026,N_12027,N_12028,N_12029,N_12030,N_12031,N_12032,N_12033,N_12034,N_12035,N_12036,N_12037,N_12038,N_12039,N_12040,N_12041,N_12042,N_12043,N_12044,N_12045,N_12046,N_12047,N_12048,N_12049,N_12050,N_12051,N_12052,N_12053,N_12054,N_12055,N_12056,N_12057,N_12058,N_12059,N_12060,N_12061,N_12062,N_12063,N_12064,N_12065,N_12066,N_12067,N_12068,N_12069,N_12070,N_12071,N_12072,N_12073,N_12074,N_12075,N_12076,N_12077,N_12078,N_12079,N_12080,N_12081,N_12082,N_12083,N_12084,N_12085,N_12086,N_12087,N_12088,N_12089,N_12090,N_12091,N_12092,N_12093,N_12094,N_12095,N_12096,N_12097,N_12098,N_12099,N_12100,N_12101,N_12102,N_12103,N_12104,N_12105,N_12106,N_12107,N_12108,N_12109,N_12110,N_12111,N_12112,N_12113,N_12114,N_12115,N_12116,N_12117,N_12118,N_12119,N_12120,N_12121,N_12122,N_12123,N_12124,N_12125,N_12126,N_12127,N_12128,N_12129,N_12130,N_12131,N_12132,N_12133,N_12134,N_12135,N_12136,N_12137,N_12138,N_12139,N_12140,N_12141,N_12142,N_12143,N_12144,N_12145,N_12146,N_12147,N_12148,N_12149,N_12150,N_12151,N_12152,N_12153,N_12154,N_12155,N_12156,N_12157,N_12158,N_12159,N_12160,N_12161,N_12162,N_12163,N_12164,N_12165,N_12166,N_12167,N_12168,N_12169,N_12170,N_12171,N_12172,N_12173,N_12174,N_12175,N_12176,N_12177,N_12178,N_12179,N_12180,N_12181,N_12182,N_12183,N_12184,N_12185,N_12186,N_12187,N_12188,N_12189,N_12190,N_12191,N_12192,N_12193,N_12194,N_12195,N_12196,N_12197,N_12198,N_12199,N_12200,N_12201,N_12202,N_12203,N_12204,N_12205,N_12206,N_12207,N_12208,N_12209,N_12210,N_12211,N_12212,N_12213,N_12214,N_12215,N_12216,N_12217,N_12218,N_12219,N_12220,N_12221,N_12222,N_12223,N_12224,N_12225,N_12226,N_12227,N_12228,N_12229,N_12230,N_12231,N_12232,N_12233,N_12234,N_12235,N_12236,N_12237,N_12238,N_12239,N_12240,N_12241,N_12242,N_12243,N_12244,N_12245,N_12246,N_12247,N_12248,N_12249,N_12250,N_12251,N_12252,N_12253,N_12254,N_12255,N_12256,N_12257,N_12258,N_12259,N_12260,N_12261,N_12262,N_12263,N_12264,N_12265,N_12266,N_12267,N_12268,N_12269,N_12270,N_12271,N_12272,N_12273,N_12274,N_12275,N_12276,N_12277,N_12278,N_12279,N_12280,N_12281,N_12282,N_12283,N_12284,N_12285,N_12286,N_12287,N_12288,N_12289,N_12290,N_12291,N_12292,N_12293,N_12294,N_12295,N_12296,N_12297,N_12298,N_12299,N_12300,N_12301,N_12302,N_12303,N_12304,N_12305,N_12306,N_12307,N_12308,N_12309,N_12310,N_12311,N_12312,N_12313,N_12314,N_12315,N_12316,N_12317,N_12318,N_12319,N_12320,N_12321,N_12322,N_12323,N_12324,N_12325,N_12326,N_12327,N_12328,N_12329,N_12330,N_12331,N_12332,N_12333,N_12334,N_12335,N_12336,N_12337,N_12338,N_12339,N_12340,N_12341,N_12342,N_12343,N_12344,N_12345,N_12346,N_12347,N_12348,N_12349,N_12350,N_12351,N_12352,N_12353,N_12354,N_12355,N_12356,N_12357,N_12358,N_12359,N_12360,N_12361,N_12362,N_12363,N_12364,N_12365,N_12366,N_12367,N_12368,N_12369,N_12370,N_12371,N_12372,N_12373,N_12374,N_12375,N_12376,N_12377,N_12378,N_12379,N_12380,N_12381,N_12382,N_12383,N_12384,N_12385,N_12386,N_12387,N_12388,N_12389,N_12390,N_12391,N_12392,N_12393,N_12394,N_12395,N_12396,N_12397,N_12398,N_12399,N_12400,N_12401,N_12402,N_12403,N_12404,N_12405,N_12406,N_12407,N_12408,N_12409,N_12410,N_12411,N_12412,N_12413,N_12414,N_12415,N_12416,N_12417,N_12418,N_12419,N_12420,N_12421,N_12422,N_12423,N_12424,N_12425,N_12426,N_12427,N_12428,N_12429,N_12430,N_12431,N_12432,N_12433,N_12434,N_12435,N_12436,N_12437,N_12438,N_12439,N_12440,N_12441,N_12442,N_12443,N_12444,N_12445,N_12446,N_12447,N_12448,N_12449,N_12450,N_12451,N_12452,N_12453,N_12454,N_12455,N_12456,N_12457,N_12458,N_12459,N_12460,N_12461,N_12462,N_12463,N_12464,N_12465,N_12466,N_12467,N_12468,N_12469,N_12470,N_12471,N_12472,N_12473,N_12474,N_12475,N_12476,N_12477,N_12478,N_12479,N_12480,N_12481,N_12482,N_12483,N_12484,N_12485,N_12486,N_12487,N_12488,N_12489,N_12490,N_12491,N_12492,N_12493,N_12494,N_12495,N_12496,N_12497,N_12498,N_12499,N_12500,N_12501,N_12502,N_12503,N_12504,N_12505,N_12506,N_12507,N_12508,N_12509,N_12510,N_12511,N_12512,N_12513,N_12514,N_12515,N_12516,N_12517,N_12518,N_12519,N_12520,N_12521,N_12522,N_12523,N_12524,N_12525,N_12526,N_12527,N_12528,N_12529,N_12530,N_12531,N_12532,N_12533,N_12534,N_12535,N_12536,N_12537,N_12538,N_12539,N_12540,N_12541,N_12542,N_12543,N_12544,N_12545,N_12546,N_12547,N_12548,N_12549,N_12550,N_12551,N_12552,N_12553,N_12554,N_12555,N_12556,N_12557,N_12558,N_12559,N_12560,N_12561,N_12562,N_12563,N_12564,N_12565,N_12566,N_12567,N_12568,N_12569,N_12570,N_12571,N_12572,N_12573,N_12574,N_12575,N_12576,N_12577,N_12578,N_12579,N_12580,N_12581,N_12582,N_12583,N_12584,N_12585,N_12586,N_12587,N_12588,N_12589,N_12590,N_12591,N_12592,N_12593,N_12594,N_12595,N_12596,N_12597,N_12598,N_12599,N_12600,N_12601,N_12602,N_12603,N_12604,N_12605,N_12606,N_12607,N_12608,N_12609,N_12610,N_12611,N_12612,N_12613,N_12614,N_12615,N_12616,N_12617,N_12618,N_12619,N_12620,N_12621,N_12622,N_12623,N_12624,N_12625,N_12626,N_12627,N_12628,N_12629,N_12630,N_12631,N_12632,N_12633,N_12634,N_12635,N_12636,N_12637,N_12638,N_12639,N_12640,N_12641,N_12642,N_12643,N_12644,N_12645,N_12646,N_12647,N_12648,N_12649,N_12650,N_12651,N_12652,N_12653,N_12654,N_12655,N_12656,N_12657,N_12658,N_12659,N_12660,N_12661,N_12662,N_12663,N_12664,N_12665,N_12666,N_12667,N_12668,N_12669,N_12670,N_12671,N_12672,N_12673,N_12674,N_12675,N_12676,N_12677,N_12678,N_12679,N_12680,N_12681,N_12682,N_12683,N_12684,N_12685,N_12686,N_12687,N_12688,N_12689,N_12690,N_12691,N_12692,N_12693,N_12694,N_12695,N_12696,N_12697,N_12698,N_12699,N_12700,N_12701,N_12702,N_12703,N_12704,N_12705,N_12706,N_12707,N_12708,N_12709,N_12710,N_12711,N_12712,N_12713,N_12714,N_12715,N_12716,N_12717,N_12718,N_12719,N_12720,N_12721,N_12722,N_12723,N_12724,N_12725,N_12726,N_12727,N_12728,N_12729,N_12730,N_12731,N_12732,N_12733,N_12734,N_12735,N_12736,N_12737,N_12738,N_12739,N_12740,N_12741,N_12742,N_12743,N_12744,N_12745,N_12746,N_12747,N_12748,N_12749,N_12750,N_12751,N_12752,N_12753,N_12754,N_12755,N_12756,N_12757,N_12758,N_12759,N_12760,N_12761,N_12762,N_12763,N_12764,N_12765,N_12766,N_12767,N_12768,N_12769,N_12770,N_12771,N_12772,N_12773,N_12774,N_12775,N_12776,N_12777,N_12778,N_12779,N_12780,N_12781,N_12782,N_12783,N_12784,N_12785,N_12786,N_12787,N_12788,N_12789,N_12790,N_12791,N_12792,N_12793,N_12794,N_12795,N_12796,N_12797,N_12798,N_12799,N_12800,N_12801,N_12802,N_12803,N_12804,N_12805,N_12806,N_12807,N_12808,N_12809,N_12810,N_12811,N_12812,N_12813,N_12814,N_12815,N_12816,N_12817,N_12818,N_12819,N_12820,N_12821,N_12822,N_12823,N_12824,N_12825,N_12826,N_12827,N_12828,N_12829,N_12830,N_12831,N_12832,N_12833,N_12834,N_12835,N_12836,N_12837,N_12838,N_12839,N_12840,N_12841,N_12842,N_12843,N_12844,N_12845,N_12846,N_12847,N_12848,N_12849,N_12850,N_12851,N_12852,N_12853,N_12854,N_12855,N_12856,N_12857,N_12858,N_12859,N_12860,N_12861,N_12862,N_12863,N_12864,N_12865,N_12866,N_12867,N_12868,N_12869,N_12870,N_12871,N_12872,N_12873,N_12874,N_12875,N_12876,N_12877,N_12878,N_12879,N_12880,N_12881,N_12882,N_12883,N_12884,N_12885,N_12886,N_12887,N_12888,N_12889,N_12890,N_12891,N_12892,N_12893,N_12894,N_12895,N_12896,N_12897,N_12898,N_12899,N_12900,N_12901,N_12902,N_12903,N_12904,N_12905,N_12906,N_12907,N_12908,N_12909,N_12910,N_12911,N_12912,N_12913,N_12914,N_12915,N_12916,N_12917,N_12918,N_12919,N_12920,N_12921,N_12922,N_12923,N_12924,N_12925,N_12926,N_12927,N_12928,N_12929,N_12930,N_12931,N_12932,N_12933,N_12934,N_12935,N_12936,N_12937,N_12938,N_12939,N_12940,N_12941,N_12942,N_12943,N_12944,N_12945,N_12946,N_12947,N_12948,N_12949,N_12950,N_12951,N_12952,N_12953,N_12954,N_12955,N_12956,N_12957,N_12958,N_12959,N_12960,N_12961,N_12962,N_12963,N_12964,N_12965,N_12966,N_12967,N_12968,N_12969,N_12970,N_12971,N_12972,N_12973,N_12974,N_12975,N_12976,N_12977,N_12978,N_12979,N_12980,N_12981,N_12982,N_12983,N_12984,N_12985,N_12986,N_12987,N_12988,N_12989,N_12990,N_12991,N_12992,N_12993,N_12994,N_12995,N_12996,N_12997,N_12998,N_12999,N_13000,N_13001,N_13002,N_13003,N_13004,N_13005,N_13006,N_13007,N_13008,N_13009,N_13010,N_13011,N_13012,N_13013,N_13014,N_13015,N_13016,N_13017,N_13018,N_13019,N_13020,N_13021,N_13022,N_13023,N_13024,N_13025,N_13026,N_13027,N_13028,N_13029,N_13030,N_13031,N_13032,N_13033,N_13034,N_13035,N_13036,N_13037,N_13038,N_13039,N_13040,N_13041,N_13042,N_13043,N_13044,N_13045,N_13046,N_13047,N_13048,N_13049,N_13050,N_13051,N_13052,N_13053,N_13054,N_13055,N_13056,N_13057,N_13058,N_13059,N_13060,N_13061,N_13062,N_13063,N_13064,N_13065,N_13066,N_13067,N_13068,N_13069,N_13070,N_13071,N_13072,N_13073,N_13074,N_13075,N_13076,N_13077,N_13078,N_13079,N_13080,N_13081,N_13082,N_13083,N_13084,N_13085,N_13086,N_13087,N_13088,N_13089,N_13090,N_13091,N_13092,N_13093,N_13094,N_13095,N_13096,N_13097,N_13098,N_13099,N_13100,N_13101,N_13102,N_13103,N_13104,N_13105,N_13106,N_13107,N_13108,N_13109,N_13110,N_13111,N_13112,N_13113,N_13114,N_13115,N_13116,N_13117,N_13118,N_13119,N_13120,N_13121,N_13122,N_13123,N_13124,N_13125,N_13126,N_13127,N_13128,N_13129,N_13130,N_13131,N_13132,N_13133,N_13134,N_13135,N_13136,N_13137,N_13138,N_13139,N_13140,N_13141,N_13142,N_13143,N_13144,N_13145,N_13146,N_13147,N_13148,N_13149,N_13150,N_13151,N_13152,N_13153,N_13154,N_13155,N_13156,N_13157,N_13158,N_13159,N_13160,N_13161,N_13162,N_13163,N_13164,N_13165,N_13166,N_13167,N_13168,N_13169,N_13170,N_13171,N_13172,N_13173,N_13174,N_13175,N_13176,N_13177,N_13178,N_13179,N_13180,N_13181,N_13182,N_13183,N_13184,N_13185,N_13186,N_13187,N_13188,N_13189,N_13190,N_13191,N_13192,N_13193,N_13194,N_13195,N_13196,N_13197,N_13198,N_13199,N_13200,N_13201,N_13202,N_13203,N_13204,N_13205,N_13206,N_13207,N_13208,N_13209,N_13210,N_13211,N_13212,N_13213,N_13214,N_13215,N_13216,N_13217,N_13218,N_13219,N_13220,N_13221,N_13222,N_13223,N_13224,N_13225,N_13226,N_13227,N_13228,N_13229,N_13230,N_13231,N_13232,N_13233,N_13234,N_13235,N_13236,N_13237,N_13238,N_13239,N_13240,N_13241,N_13242,N_13243,N_13244,N_13245,N_13246,N_13247,N_13248,N_13249,N_13250,N_13251,N_13252,N_13253,N_13254,N_13255,N_13256,N_13257,N_13258,N_13259,N_13260,N_13261,N_13262,N_13263,N_13264,N_13265,N_13266,N_13267,N_13268,N_13269,N_13270,N_13271,N_13272,N_13273,N_13274,N_13275,N_13276,N_13277,N_13278,N_13279,N_13280,N_13281,N_13282,N_13283,N_13284,N_13285,N_13286,N_13287,N_13288,N_13289,N_13290,N_13291,N_13292,N_13293,N_13294,N_13295,N_13296,N_13297,N_13298,N_13299,N_13300,N_13301,N_13302,N_13303,N_13304,N_13305,N_13306,N_13307,N_13308,N_13309,N_13310,N_13311,N_13312,N_13313,N_13314,N_13315,N_13316,N_13317,N_13318,N_13319,N_13320,N_13321,N_13322,N_13323,N_13324,N_13325,N_13326,N_13327,N_13328,N_13329,N_13330,N_13331,N_13332,N_13333,N_13334,N_13335,N_13336,N_13337,N_13338,N_13339,N_13340,N_13341,N_13342,N_13343,N_13344,N_13345,N_13346,N_13347,N_13348,N_13349,N_13350,N_13351,N_13352,N_13353,N_13354,N_13355,N_13356,N_13357,N_13358,N_13359,N_13360,N_13361,N_13362,N_13363,N_13364,N_13365,N_13366,N_13367,N_13368,N_13369,N_13370,N_13371,N_13372,N_13373,N_13374,N_13375,N_13376,N_13377,N_13378,N_13379,N_13380,N_13381,N_13382,N_13383,N_13384,N_13385,N_13386,N_13387,N_13388,N_13389,N_13390,N_13391,N_13392,N_13393,N_13394,N_13395,N_13396,N_13397,N_13398,N_13399,N_13400,N_13401,N_13402,N_13403,N_13404,N_13405,N_13406,N_13407,N_13408,N_13409,N_13410,N_13411,N_13412,N_13413,N_13414,N_13415,N_13416,N_13417,N_13418,N_13419,N_13420,N_13421,N_13422,N_13423,N_13424,N_13425,N_13426,N_13427,N_13428,N_13429,N_13430,N_13431,N_13432,N_13433,N_13434,N_13435,N_13436,N_13437,N_13438,N_13439,N_13440,N_13441,N_13442,N_13443,N_13444,N_13445,N_13446,N_13447,N_13448,N_13449,N_13450,N_13451,N_13452,N_13453,N_13454,N_13455,N_13456,N_13457,N_13458,N_13459,N_13460,N_13461,N_13462,N_13463,N_13464,N_13465,N_13466,N_13467,N_13468,N_13469,N_13470,N_13471,N_13472,N_13473,N_13474,N_13475,N_13476,N_13477,N_13478,N_13479,N_13480,N_13481,N_13482,N_13483,N_13484,N_13485,N_13486,N_13487,N_13488,N_13489,N_13490,N_13491,N_13492,N_13493,N_13494,N_13495,N_13496,N_13497,N_13498,N_13499,N_13500,N_13501,N_13502,N_13503,N_13504,N_13505,N_13506,N_13507,N_13508,N_13509,N_13510,N_13511,N_13512,N_13513,N_13514,N_13515,N_13516,N_13517,N_13518,N_13519,N_13520,N_13521,N_13522,N_13523,N_13524,N_13525,N_13526,N_13527,N_13528,N_13529,N_13530,N_13531,N_13532,N_13533,N_13534,N_13535,N_13536,N_13537,N_13538,N_13539,N_13540,N_13541,N_13542,N_13543,N_13544,N_13545,N_13546,N_13547,N_13548,N_13549,N_13550,N_13551,N_13552,N_13553,N_13554,N_13555,N_13556,N_13557,N_13558,N_13559,N_13560,N_13561,N_13562,N_13563,N_13564,N_13565,N_13566,N_13567,N_13568,N_13569,N_13570,N_13571,N_13572,N_13573,N_13574,N_13575,N_13576,N_13577,N_13578,N_13579,N_13580,N_13581,N_13582,N_13583,N_13584,N_13585,N_13586,N_13587,N_13588,N_13589,N_13590,N_13591,N_13592,N_13593,N_13594,N_13595,N_13596,N_13597,N_13598,N_13599,N_13600,N_13601,N_13602,N_13603,N_13604,N_13605,N_13606,N_13607,N_13608,N_13609,N_13610,N_13611,N_13612,N_13613,N_13614,N_13615,N_13616,N_13617,N_13618,N_13619,N_13620,N_13621,N_13622,N_13623,N_13624,N_13625,N_13626,N_13627,N_13628,N_13629,N_13630,N_13631,N_13632,N_13633,N_13634,N_13635,N_13636,N_13637,N_13638,N_13639,N_13640,N_13641,N_13642,N_13643,N_13644,N_13645,N_13646,N_13647,N_13648,N_13649,N_13650,N_13651,N_13652,N_13653,N_13654,N_13655,N_13656,N_13657,N_13658,N_13659,N_13660,N_13661,N_13662,N_13663,N_13664,N_13665,N_13666,N_13667,N_13668,N_13669,N_13670,N_13671,N_13672,N_13673,N_13674,N_13675,N_13676,N_13677,N_13678,N_13679,N_13680,N_13681,N_13682,N_13683,N_13684,N_13685,N_13686,N_13687,N_13688,N_13689,N_13690,N_13691,N_13692,N_13693,N_13694,N_13695,N_13696,N_13697,N_13698,N_13699,N_13700,N_13701,N_13702,N_13703,N_13704,N_13705,N_13706,N_13707,N_13708,N_13709,N_13710,N_13711,N_13712,N_13713,N_13714,N_13715,N_13716,N_13717,N_13718,N_13719,N_13720,N_13721,N_13722,N_13723,N_13724,N_13725,N_13726,N_13727,N_13728,N_13729,N_13730,N_13731,N_13732,N_13733,N_13734,N_13735,N_13736,N_13737,N_13738,N_13739,N_13740,N_13741,N_13742,N_13743,N_13744,N_13745,N_13746,N_13747,N_13748,N_13749,N_13750,N_13751,N_13752,N_13753,N_13754,N_13755,N_13756,N_13757,N_13758,N_13759,N_13760,N_13761,N_13762,N_13763,N_13764,N_13765,N_13766,N_13767,N_13768,N_13769,N_13770,N_13771,N_13772,N_13773,N_13774,N_13775,N_13776,N_13777,N_13778,N_13779,N_13780,N_13781,N_13782,N_13783,N_13784,N_13785,N_13786,N_13787,N_13788,N_13789,N_13790,N_13791,N_13792,N_13793,N_13794,N_13795,N_13796,N_13797,N_13798,N_13799,N_13800,N_13801,N_13802,N_13803,N_13804,N_13805,N_13806,N_13807,N_13808,N_13809,N_13810,N_13811,N_13812,N_13813,N_13814,N_13815,N_13816,N_13817,N_13818,N_13819,N_13820,N_13821,N_13822,N_13823,N_13824,N_13825,N_13826,N_13827,N_13828,N_13829,N_13830,N_13831,N_13832,N_13833,N_13834,N_13835,N_13836,N_13837,N_13838,N_13839,N_13840,N_13841,N_13842,N_13843,N_13844,N_13845,N_13846,N_13847,N_13848,N_13849,N_13850,N_13851,N_13852,N_13853,N_13854,N_13855,N_13856,N_13857,N_13858,N_13859,N_13860,N_13861,N_13862,N_13863,N_13864,N_13865,N_13866,N_13867,N_13868,N_13869,N_13870,N_13871,N_13872,N_13873,N_13874,N_13875,N_13876,N_13877,N_13878,N_13879,N_13880,N_13881,N_13882,N_13883,N_13884,N_13885,N_13886,N_13887,N_13888,N_13889,N_13890,N_13891,N_13892,N_13893,N_13894,N_13895,N_13896,N_13897,N_13898,N_13899,N_13900,N_13901,N_13902,N_13903,N_13904,N_13905,N_13906,N_13907,N_13908,N_13909,N_13910,N_13911,N_13912,N_13913,N_13914,N_13915,N_13916,N_13917,N_13918,N_13919,N_13920,N_13921,N_13922,N_13923,N_13924,N_13925,N_13926,N_13927,N_13928,N_13929,N_13930,N_13931,N_13932,N_13933,N_13934,N_13935,N_13936,N_13937,N_13938,N_13939,N_13940,N_13941,N_13942,N_13943,N_13944,N_13945,N_13946,N_13947,N_13948,N_13949,N_13950,N_13951,N_13952,N_13953,N_13954,N_13955,N_13956,N_13957,N_13958,N_13959,N_13960,N_13961,N_13962,N_13963,N_13964,N_13965,N_13966,N_13967,N_13968,N_13969,N_13970,N_13971,N_13972,N_13973,N_13974,N_13975,N_13976,N_13977,N_13978,N_13979,N_13980,N_13981,N_13982,N_13983,N_13984,N_13985,N_13986,N_13987,N_13988,N_13989,N_13990,N_13991,N_13992,N_13993,N_13994,N_13995,N_13996,N_13997,N_13998,N_13999,N_14000,N_14001,N_14002,N_14003,N_14004,N_14005,N_14006,N_14007,N_14008,N_14009,N_14010,N_14011,N_14012,N_14013,N_14014,N_14015,N_14016,N_14017,N_14018,N_14019,N_14020,N_14021,N_14022,N_14023,N_14024,N_14025,N_14026,N_14027,N_14028,N_14029,N_14030,N_14031,N_14032,N_14033,N_14034,N_14035,N_14036,N_14037,N_14038,N_14039,N_14040,N_14041,N_14042,N_14043,N_14044,N_14045,N_14046,N_14047,N_14048,N_14049,N_14050,N_14051,N_14052,N_14053,N_14054,N_14055,N_14056,N_14057,N_14058,N_14059,N_14060,N_14061,N_14062,N_14063,N_14064,N_14065,N_14066,N_14067,N_14068,N_14069,N_14070,N_14071,N_14072,N_14073,N_14074,N_14075,N_14076,N_14077,N_14078,N_14079,N_14080,N_14081,N_14082,N_14083,N_14084,N_14085,N_14086,N_14087,N_14088,N_14089,N_14090,N_14091,N_14092,N_14093,N_14094,N_14095,N_14096,N_14097,N_14098,N_14099,N_14100,N_14101,N_14102,N_14103,N_14104,N_14105,N_14106,N_14107,N_14108,N_14109,N_14110,N_14111,N_14112,N_14113,N_14114,N_14115,N_14116,N_14117,N_14118,N_14119,N_14120,N_14121,N_14122,N_14123,N_14124,N_14125,N_14126,N_14127,N_14128,N_14129,N_14130,N_14131,N_14132,N_14133,N_14134,N_14135,N_14136,N_14137,N_14138,N_14139,N_14140,N_14141,N_14142,N_14143,N_14144,N_14145,N_14146,N_14147,N_14148,N_14149,N_14150,N_14151,N_14152,N_14153,N_14154,N_14155,N_14156,N_14157,N_14158,N_14159,N_14160,N_14161,N_14162,N_14163,N_14164,N_14165,N_14166,N_14167,N_14168,N_14169,N_14170,N_14171,N_14172,N_14173,N_14174,N_14175,N_14176,N_14177,N_14178,N_14179,N_14180,N_14181,N_14182,N_14183,N_14184,N_14185,N_14186,N_14187,N_14188,N_14189,N_14190,N_14191,N_14192,N_14193,N_14194,N_14195,N_14196,N_14197,N_14198,N_14199,N_14200,N_14201,N_14202,N_14203,N_14204,N_14205,N_14206,N_14207,N_14208,N_14209,N_14210,N_14211,N_14212,N_14213,N_14214,N_14215,N_14216,N_14217,N_14218,N_14219,N_14220,N_14221,N_14222,N_14223,N_14224,N_14225,N_14226,N_14227,N_14228,N_14229,N_14230,N_14231,N_14232,N_14233,N_14234,N_14235,N_14236,N_14237,N_14238,N_14239,N_14240,N_14241,N_14242,N_14243,N_14244,N_14245,N_14246,N_14247,N_14248,N_14249,N_14250,N_14251,N_14252,N_14253,N_14254,N_14255,N_14256,N_14257,N_14258,N_14259,N_14260,N_14261,N_14262,N_14263,N_14264,N_14265,N_14266,N_14267,N_14268,N_14269,N_14270,N_14271,N_14272,N_14273,N_14274,N_14275,N_14276,N_14277,N_14278,N_14279,N_14280,N_14281,N_14282,N_14283,N_14284,N_14285,N_14286,N_14287,N_14288,N_14289,N_14290,N_14291,N_14292,N_14293,N_14294,N_14295,N_14296,N_14297,N_14298,N_14299,N_14300,N_14301,N_14302,N_14303,N_14304,N_14305,N_14306,N_14307,N_14308,N_14309,N_14310,N_14311,N_14312,N_14313,N_14314,N_14315,N_14316,N_14317,N_14318,N_14319,N_14320,N_14321,N_14322,N_14323,N_14324,N_14325,N_14326,N_14327,N_14328,N_14329,N_14330,N_14331,N_14332,N_14333,N_14334,N_14335,N_14336,N_14337,N_14338,N_14339,N_14340,N_14341,N_14342,N_14343,N_14344,N_14345,N_14346,N_14347,N_14348,N_14349,N_14350,N_14351,N_14352,N_14353,N_14354,N_14355,N_14356,N_14357,N_14358,N_14359,N_14360,N_14361,N_14362,N_14363,N_14364,N_14365,N_14366,N_14367,N_14368,N_14369,N_14370,N_14371,N_14372,N_14373,N_14374,N_14375,N_14376,N_14377,N_14378,N_14379,N_14380,N_14381,N_14382,N_14383,N_14384,N_14385,N_14386,N_14387,N_14388,N_14389,N_14390,N_14391,N_14392,N_14393,N_14394,N_14395,N_14396,N_14397,N_14398,N_14399,N_14400,N_14401,N_14402,N_14403,N_14404,N_14405,N_14406,N_14407,N_14408,N_14409,N_14410,N_14411,N_14412,N_14413,N_14414,N_14415,N_14416,N_14417,N_14418,N_14419,N_14420,N_14421,N_14422,N_14423,N_14424,N_14425,N_14426,N_14427,N_14428,N_14429,N_14430,N_14431,N_14432,N_14433,N_14434,N_14435,N_14436,N_14437,N_14438,N_14439,N_14440,N_14441,N_14442,N_14443,N_14444,N_14445,N_14446,N_14447,N_14448,N_14449,N_14450,N_14451,N_14452,N_14453,N_14454,N_14455,N_14456,N_14457,N_14458,N_14459,N_14460,N_14461,N_14462,N_14463,N_14464,N_14465,N_14466,N_14467,N_14468,N_14469,N_14470,N_14471,N_14472,N_14473,N_14474,N_14475,N_14476,N_14477,N_14478,N_14479,N_14480,N_14481,N_14482,N_14483,N_14484,N_14485,N_14486,N_14487,N_14488,N_14489,N_14490,N_14491,N_14492,N_14493,N_14494,N_14495,N_14496,N_14497,N_14498,N_14499,N_14500,N_14501,N_14502,N_14503,N_14504,N_14505,N_14506,N_14507,N_14508,N_14509,N_14510,N_14511,N_14512,N_14513,N_14514,N_14515,N_14516,N_14517,N_14518,N_14519,N_14520,N_14521,N_14522,N_14523,N_14524,N_14525,N_14526,N_14527,N_14528,N_14529,N_14530,N_14531,N_14532,N_14533,N_14534,N_14535,N_14536,N_14537,N_14538,N_14539,N_14540,N_14541,N_14542,N_14543,N_14544,N_14545,N_14546,N_14547,N_14548,N_14549,N_14550,N_14551,N_14552,N_14553,N_14554,N_14555,N_14556,N_14557,N_14558,N_14559,N_14560,N_14561,N_14562,N_14563,N_14564,N_14565,N_14566,N_14567,N_14568,N_14569,N_14570,N_14571,N_14572,N_14573,N_14574,N_14575,N_14576,N_14577,N_14578,N_14579,N_14580,N_14581,N_14582,N_14583,N_14584,N_14585,N_14586,N_14587,N_14588,N_14589,N_14590,N_14591,N_14592,N_14593,N_14594,N_14595,N_14596,N_14597,N_14598,N_14599,N_14600,N_14601,N_14602,N_14603,N_14604,N_14605,N_14606,N_14607,N_14608,N_14609,N_14610,N_14611,N_14612,N_14613,N_14614,N_14615,N_14616,N_14617,N_14618,N_14619,N_14620,N_14621,N_14622,N_14623,N_14624,N_14625,N_14626,N_14627,N_14628,N_14629,N_14630,N_14631,N_14632,N_14633,N_14634,N_14635,N_14636,N_14637,N_14638,N_14639,N_14640,N_14641,N_14642,N_14643,N_14644,N_14645,N_14646,N_14647,N_14648,N_14649,N_14650,N_14651,N_14652,N_14653,N_14654,N_14655,N_14656,N_14657,N_14658,N_14659,N_14660,N_14661,N_14662,N_14663,N_14664,N_14665,N_14666,N_14667,N_14668,N_14669,N_14670,N_14671,N_14672,N_14673,N_14674,N_14675,N_14676,N_14677,N_14678,N_14679,N_14680,N_14681,N_14682,N_14683,N_14684,N_14685,N_14686,N_14687,N_14688,N_14689,N_14690,N_14691,N_14692,N_14693,N_14694,N_14695,N_14696,N_14697,N_14698,N_14699,N_14700,N_14701,N_14702,N_14703,N_14704,N_14705,N_14706,N_14707,N_14708,N_14709,N_14710,N_14711,N_14712,N_14713,N_14714,N_14715,N_14716,N_14717,N_14718,N_14719,N_14720,N_14721,N_14722,N_14723,N_14724,N_14725,N_14726,N_14727,N_14728,N_14729,N_14730,N_14731,N_14732,N_14733,N_14734,N_14735,N_14736,N_14737,N_14738,N_14739,N_14740,N_14741,N_14742,N_14743,N_14744,N_14745,N_14746,N_14747,N_14748,N_14749,N_14750,N_14751,N_14752,N_14753,N_14754,N_14755,N_14756,N_14757,N_14758,N_14759,N_14760,N_14761,N_14762,N_14763,N_14764,N_14765,N_14766,N_14767,N_14768,N_14769,N_14770,N_14771,N_14772,N_14773,N_14774,N_14775,N_14776,N_14777,N_14778,N_14779,N_14780,N_14781,N_14782,N_14783,N_14784,N_14785,N_14786,N_14787,N_14788,N_14789,N_14790,N_14791,N_14792,N_14793,N_14794,N_14795,N_14796,N_14797,N_14798,N_14799,N_14800,N_14801,N_14802,N_14803,N_14804,N_14805,N_14806,N_14807,N_14808,N_14809,N_14810,N_14811,N_14812,N_14813,N_14814,N_14815,N_14816,N_14817,N_14818,N_14819,N_14820,N_14821,N_14822,N_14823,N_14824,N_14825,N_14826,N_14827,N_14828,N_14829,N_14830,N_14831,N_14832,N_14833,N_14834,N_14835,N_14836,N_14837,N_14838,N_14839,N_14840,N_14841,N_14842,N_14843,N_14844,N_14845,N_14846,N_14847,N_14848,N_14849,N_14850,N_14851,N_14852,N_14853,N_14854,N_14855,N_14856,N_14857,N_14858,N_14859,N_14860,N_14861,N_14862,N_14863,N_14864,N_14865,N_14866,N_14867,N_14868,N_14869,N_14870,N_14871,N_14872,N_14873,N_14874,N_14875,N_14876,N_14877,N_14878,N_14879,N_14880,N_14881,N_14882,N_14883,N_14884,N_14885,N_14886,N_14887,N_14888,N_14889,N_14890,N_14891,N_14892,N_14893,N_14894,N_14895,N_14896,N_14897,N_14898,N_14899,N_14900,N_14901,N_14902,N_14903,N_14904,N_14905,N_14906,N_14907,N_14908,N_14909,N_14910,N_14911,N_14912,N_14913,N_14914,N_14915,N_14916,N_14917,N_14918,N_14919,N_14920,N_14921,N_14922,N_14923,N_14924,N_14925,N_14926,N_14927,N_14928,N_14929,N_14930,N_14931,N_14932,N_14933,N_14934,N_14935,N_14936,N_14937,N_14938,N_14939,N_14940,N_14941,N_14942,N_14943,N_14944,N_14945,N_14946,N_14947,N_14948,N_14949,N_14950,N_14951,N_14952,N_14953,N_14954,N_14955,N_14956,N_14957,N_14958,N_14959,N_14960,N_14961,N_14962,N_14963,N_14964,N_14965,N_14966,N_14967,N_14968,N_14969,N_14970,N_14971,N_14972,N_14973,N_14974,N_14975,N_14976,N_14977,N_14978,N_14979,N_14980,N_14981,N_14982,N_14983,N_14984,N_14985,N_14986,N_14987,N_14988,N_14989,N_14990,N_14991,N_14992,N_14993,N_14994,N_14995,N_14996,N_14997,N_14998,N_14999,N_15000,N_15001,N_15002,N_15003,N_15004,N_15005,N_15006,N_15007,N_15008,N_15009,N_15010,N_15011,N_15012,N_15013,N_15014,N_15015,N_15016,N_15017,N_15018,N_15019,N_15020,N_15021,N_15022,N_15023,N_15024,N_15025,N_15026,N_15027,N_15028,N_15029,N_15030,N_15031,N_15032,N_15033,N_15034,N_15035,N_15036,N_15037,N_15038,N_15039,N_15040,N_15041,N_15042,N_15043,N_15044,N_15045,N_15046,N_15047,N_15048,N_15049,N_15050,N_15051,N_15052,N_15053,N_15054,N_15055,N_15056,N_15057,N_15058,N_15059,N_15060,N_15061,N_15062,N_15063,N_15064,N_15065,N_15066,N_15067,N_15068,N_15069,N_15070,N_15071,N_15072,N_15073,N_15074,N_15075,N_15076,N_15077,N_15078,N_15079,N_15080,N_15081,N_15082,N_15083,N_15084,N_15085,N_15086,N_15087,N_15088,N_15089,N_15090,N_15091,N_15092,N_15093,N_15094,N_15095,N_15096,N_15097,N_15098,N_15099,N_15100,N_15101,N_15102,N_15103,N_15104,N_15105,N_15106,N_15107,N_15108,N_15109,N_15110,N_15111,N_15112,N_15113,N_15114,N_15115,N_15116,N_15117,N_15118,N_15119,N_15120,N_15121,N_15122,N_15123,N_15124,N_15125,N_15126,N_15127,N_15128,N_15129,N_15130,N_15131,N_15132,N_15133,N_15134,N_15135,N_15136,N_15137,N_15138,N_15139,N_15140,N_15141,N_15142,N_15143,N_15144,N_15145,N_15146,N_15147,N_15148,N_15149,N_15150,N_15151,N_15152,N_15153,N_15154,N_15155,N_15156,N_15157,N_15158,N_15159,N_15160,N_15161,N_15162,N_15163,N_15164,N_15165,N_15166,N_15167,N_15168,N_15169,N_15170,N_15171,N_15172,N_15173,N_15174,N_15175,N_15176,N_15177,N_15178,N_15179,N_15180,N_15181,N_15182,N_15183,N_15184,N_15185,N_15186,N_15187,N_15188,N_15189,N_15190,N_15191,N_15192,N_15193,N_15194,N_15195,N_15196,N_15197,N_15198,N_15199,N_15200,N_15201,N_15202,N_15203,N_15204,N_15205,N_15206,N_15207,N_15208,N_15209,N_15210,N_15211,N_15212,N_15213,N_15214,N_15215,N_15216,N_15217,N_15218,N_15219,N_15220,N_15221,N_15222,N_15223,N_15224,N_15225,N_15226,N_15227,N_15228,N_15229,N_15230,N_15231,N_15232,N_15233,N_15234,N_15235,N_15236,N_15237,N_15238,N_15239,N_15240,N_15241,N_15242,N_15243,N_15244,N_15245,N_15246,N_15247,N_15248,N_15249,N_15250,N_15251,N_15252,N_15253,N_15254,N_15255,N_15256,N_15257,N_15258,N_15259,N_15260,N_15261,N_15262,N_15263,N_15264,N_15265,N_15266,N_15267,N_15268,N_15269,N_15270,N_15271,N_15272,N_15273,N_15274,N_15275,N_15276,N_15277,N_15278,N_15279,N_15280,N_15281,N_15282,N_15283,N_15284,N_15285,N_15286,N_15287,N_15288,N_15289,N_15290,N_15291,N_15292,N_15293,N_15294,N_15295,N_15296,N_15297,N_15298,N_15299,N_15300,N_15301,N_15302,N_15303,N_15304,N_15305,N_15306,N_15307,N_15308,N_15309,N_15310,N_15311,N_15312,N_15313,N_15314,N_15315,N_15316,N_15317,N_15318,N_15319,N_15320,N_15321,N_15322,N_15323,N_15324,N_15325,N_15326,N_15327,N_15328,N_15329,N_15330,N_15331,N_15332,N_15333,N_15334,N_15335,N_15336,N_15337,N_15338,N_15339,N_15340,N_15341,N_15342,N_15343,N_15344,N_15345,N_15346,N_15347,N_15348,N_15349,N_15350,N_15351,N_15352,N_15353,N_15354,N_15355,N_15356,N_15357,N_15358,N_15359,N_15360,N_15361,N_15362,N_15363,N_15364,N_15365,N_15366,N_15367,N_15368,N_15369,N_15370,N_15371,N_15372,N_15373,N_15374,N_15375,N_15376,N_15377,N_15378,N_15379,N_15380,N_15381,N_15382,N_15383,N_15384,N_15385,N_15386,N_15387,N_15388,N_15389,N_15390,N_15391,N_15392,N_15393,N_15394,N_15395,N_15396,N_15397,N_15398,N_15399,N_15400,N_15401,N_15402,N_15403,N_15404,N_15405,N_15406,N_15407,N_15408,N_15409,N_15410,N_15411,N_15412,N_15413,N_15414,N_15415,N_15416,N_15417,N_15418,N_15419,N_15420,N_15421,N_15422,N_15423,N_15424,N_15425,N_15426,N_15427,N_15428,N_15429,N_15430,N_15431,N_15432,N_15433,N_15434,N_15435,N_15436,N_15437,N_15438,N_15439,N_15440,N_15441,N_15442,N_15443,N_15444,N_15445,N_15446,N_15447,N_15448,N_15449,N_15450,N_15451,N_15452,N_15453,N_15454,N_15455,N_15456,N_15457,N_15458,N_15459,N_15460,N_15461,N_15462,N_15463,N_15464,N_15465,N_15466,N_15467,N_15468,N_15469,N_15470,N_15471,N_15472,N_15473,N_15474,N_15475,N_15476,N_15477,N_15478,N_15479,N_15480,N_15481,N_15482,N_15483,N_15484,N_15485,N_15486,N_15487,N_15488,N_15489,N_15490,N_15491,N_15492,N_15493,N_15494,N_15495,N_15496,N_15497,N_15498,N_15499,N_15500,N_15501,N_15502,N_15503,N_15504,N_15505,N_15506,N_15507,N_15508,N_15509,N_15510,N_15511,N_15512,N_15513,N_15514,N_15515,N_15516,N_15517,N_15518,N_15519,N_15520,N_15521,N_15522,N_15523,N_15524,N_15525,N_15526,N_15527,N_15528,N_15529,N_15530,N_15531,N_15532,N_15533,N_15534,N_15535,N_15536,N_15537,N_15538,N_15539,N_15540,N_15541,N_15542,N_15543,N_15544,N_15545,N_15546,N_15547,N_15548,N_15549,N_15550,N_15551,N_15552,N_15553,N_15554,N_15555,N_15556,N_15557,N_15558,N_15559,N_15560,N_15561,N_15562,N_15563,N_15564,N_15565,N_15566,N_15567,N_15568,N_15569,N_15570,N_15571,N_15572,N_15573,N_15574,N_15575,N_15576,N_15577,N_15578,N_15579,N_15580,N_15581,N_15582,N_15583,N_15584,N_15585,N_15586,N_15587,N_15588,N_15589,N_15590,N_15591,N_15592,N_15593,N_15594,N_15595,N_15596,N_15597,N_15598,N_15599,N_15600,N_15601,N_15602,N_15603,N_15604,N_15605,N_15606,N_15607,N_15608,N_15609,N_15610,N_15611,N_15612,N_15613,N_15614,N_15615,N_15616,N_15617,N_15618,N_15619,N_15620,N_15621,N_15622,N_15623,N_15624,N_15625,N_15626,N_15627,N_15628,N_15629,N_15630,N_15631,N_15632,N_15633,N_15634,N_15635,N_15636,N_15637,N_15638,N_15639,N_15640,N_15641,N_15642,N_15643,N_15644,N_15645,N_15646,N_15647,N_15648,N_15649,N_15650,N_15651,N_15652,N_15653,N_15654,N_15655,N_15656,N_15657,N_15658,N_15659,N_15660,N_15661,N_15662,N_15663,N_15664,N_15665,N_15666,N_15667,N_15668,N_15669,N_15670,N_15671,N_15672,N_15673,N_15674,N_15675,N_15676,N_15677,N_15678,N_15679,N_15680,N_15681,N_15682,N_15683,N_15684,N_15685,N_15686,N_15687,N_15688,N_15689,N_15690,N_15691,N_15692,N_15693,N_15694,N_15695,N_15696,N_15697,N_15698,N_15699,N_15700,N_15701,N_15702,N_15703,N_15704,N_15705,N_15706,N_15707,N_15708,N_15709,N_15710,N_15711,N_15712,N_15713,N_15714,N_15715,N_15716,N_15717,N_15718,N_15719,N_15720,N_15721,N_15722,N_15723,N_15724,N_15725,N_15726,N_15727,N_15728,N_15729,N_15730,N_15731,N_15732,N_15733,N_15734,N_15735,N_15736,N_15737,N_15738,N_15739,N_15740,N_15741,N_15742,N_15743,N_15744,N_15745,N_15746,N_15747,N_15748,N_15749,N_15750,N_15751,N_15752,N_15753,N_15754,N_15755,N_15756,N_15757,N_15758,N_15759,N_15760,N_15761,N_15762,N_15763,N_15764,N_15765,N_15766,N_15767,N_15768,N_15769,N_15770,N_15771,N_15772,N_15773,N_15774,N_15775,N_15776,N_15777,N_15778,N_15779,N_15780,N_15781,N_15782,N_15783,N_15784,N_15785,N_15786,N_15787,N_15788,N_15789,N_15790,N_15791,N_15792,N_15793,N_15794,N_15795,N_15796,N_15797,N_15798,N_15799,N_15800,N_15801,N_15802,N_15803,N_15804,N_15805,N_15806,N_15807,N_15808,N_15809,N_15810,N_15811,N_15812,N_15813,N_15814,N_15815,N_15816,N_15817,N_15818,N_15819,N_15820,N_15821,N_15822,N_15823,N_15824,N_15825,N_15826,N_15827,N_15828,N_15829,N_15830,N_15831,N_15832,N_15833,N_15834,N_15835,N_15836,N_15837,N_15838,N_15839,N_15840,N_15841,N_15842,N_15843,N_15844,N_15845,N_15846,N_15847,N_15848,N_15849,N_15850,N_15851,N_15852,N_15853,N_15854,N_15855,N_15856,N_15857,N_15858,N_15859,N_15860,N_15861,N_15862,N_15863,N_15864,N_15865,N_15866,N_15867,N_15868,N_15869,N_15870,N_15871,N_15872,N_15873,N_15874,N_15875,N_15876,N_15877,N_15878,N_15879,N_15880,N_15881,N_15882,N_15883,N_15884,N_15885,N_15886,N_15887,N_15888,N_15889,N_15890,N_15891,N_15892,N_15893,N_15894,N_15895,N_15896,N_15897,N_15898,N_15899,N_15900,N_15901,N_15902,N_15903,N_15904,N_15905,N_15906,N_15907,N_15908,N_15909,N_15910,N_15911,N_15912,N_15913,N_15914,N_15915,N_15916,N_15917,N_15918,N_15919,N_15920,N_15921,N_15922,N_15923,N_15924,N_15925,N_15926,N_15927,N_15928,N_15929,N_15930,N_15931,N_15932,N_15933,N_15934,N_15935,N_15936,N_15937,N_15938,N_15939,N_15940,N_15941,N_15942,N_15943,N_15944,N_15945,N_15946,N_15947,N_15948,N_15949,N_15950,N_15951,N_15952,N_15953,N_15954,N_15955,N_15956,N_15957,N_15958,N_15959,N_15960,N_15961,N_15962,N_15963,N_15964,N_15965,N_15966,N_15967,N_15968,N_15969,N_15970,N_15971,N_15972,N_15973,N_15974,N_15975,N_15976,N_15977,N_15978,N_15979,N_15980,N_15981,N_15982,N_15983,N_15984,N_15985,N_15986,N_15987,N_15988,N_15989,N_15990,N_15991,N_15992,N_15993,N_15994,N_15995,N_15996,N_15997,N_15998,N_15999,N_16000,N_16001,N_16002,N_16003,N_16004,N_16005,N_16006,N_16007,N_16008,N_16009,N_16010,N_16011,N_16012,N_16013,N_16014,N_16015,N_16016,N_16017,N_16018,N_16019,N_16020,N_16021,N_16022,N_16023,N_16024,N_16025,N_16026,N_16027,N_16028,N_16029,N_16030,N_16031,N_16032,N_16033,N_16034,N_16035,N_16036,N_16037,N_16038,N_16039,N_16040,N_16041,N_16042,N_16043,N_16044,N_16045,N_16046,N_16047,N_16048,N_16049,N_16050,N_16051,N_16052,N_16053,N_16054,N_16055,N_16056,N_16057,N_16058,N_16059,N_16060,N_16061,N_16062,N_16063,N_16064,N_16065,N_16066,N_16067,N_16068,N_16069,N_16070,N_16071,N_16072,N_16073,N_16074,N_16075,N_16076,N_16077,N_16078,N_16079,N_16080,N_16081,N_16082,N_16083,N_16084,N_16085,N_16086,N_16087,N_16088,N_16089,N_16090,N_16091,N_16092,N_16093,N_16094,N_16095,N_16096,N_16097,N_16098,N_16099,N_16100,N_16101,N_16102,N_16103,N_16104,N_16105,N_16106,N_16107,N_16108,N_16109,N_16110,N_16111,N_16112,N_16113,N_16114,N_16115,N_16116,N_16117,N_16118,N_16119,N_16120,N_16121,N_16122,N_16123,N_16124,N_16125,N_16126,N_16127,N_16128,N_16129,N_16130,N_16131,N_16132,N_16133,N_16134,N_16135,N_16136,N_16137,N_16138,N_16139,N_16140,N_16141,N_16142,N_16143,N_16144,N_16145,N_16146,N_16147,N_16148,N_16149,N_16150,N_16151,N_16152,N_16153,N_16154,N_16155,N_16156,N_16157,N_16158,N_16159,N_16160,N_16161,N_16162,N_16163,N_16164,N_16165,N_16166,N_16167,N_16168,N_16169,N_16170,N_16171,N_16172,N_16173,N_16174,N_16175,N_16176,N_16177,N_16178,N_16179,N_16180,N_16181,N_16182,N_16183,N_16184,N_16185,N_16186,N_16187,N_16188,N_16189,N_16190,N_16191,N_16192,N_16193,N_16194,N_16195,N_16196,N_16197,N_16198,N_16199,N_16200,N_16201,N_16202,N_16203,N_16204,N_16205,N_16206,N_16207,N_16208,N_16209,N_16210,N_16211,N_16212,N_16213,N_16214,N_16215,N_16216,N_16217,N_16218,N_16219,N_16220,N_16221,N_16222,N_16223,N_16224,N_16225,N_16226,N_16227,N_16228,N_16229,N_16230,N_16231,N_16232,N_16233,N_16234,N_16235,N_16236,N_16237,N_16238,N_16239,N_16240,N_16241,N_16242,N_16243,N_16244,N_16245,N_16246,N_16247,N_16248,N_16249,N_16250,N_16251,N_16252,N_16253,N_16254,N_16255,N_16256,N_16257,N_16258,N_16259,N_16260,N_16261,N_16262,N_16263,N_16264,N_16265,N_16266,N_16267,N_16268,N_16269,N_16270,N_16271,N_16272,N_16273,N_16274,N_16275,N_16276,N_16277,N_16278,N_16279,N_16280,N_16281,N_16282,N_16283,N_16284,N_16285,N_16286,N_16287,N_16288,N_16289,N_16290,N_16291,N_16292,N_16293,N_16294,N_16295,N_16296,N_16297,N_16298,N_16299,N_16300,N_16301,N_16302,N_16303,N_16304,N_16305,N_16306,N_16307,N_16308,N_16309,N_16310,N_16311,N_16312,N_16313,N_16314,N_16315,N_16316,N_16317,N_16318,N_16319,N_16320,N_16321,N_16322,N_16323,N_16324,N_16325,N_16326,N_16327,N_16328,N_16329,N_16330,N_16331,N_16332,N_16333,N_16334,N_16335,N_16336,N_16337,N_16338,N_16339,N_16340,N_16341,N_16342,N_16343,N_16344,N_16345,N_16346,N_16347,N_16348,N_16349,N_16350,N_16351,N_16352,N_16353,N_16354,N_16355,N_16356,N_16357,N_16358,N_16359,N_16360,N_16361,N_16362,N_16363,N_16364,N_16365,N_16366,N_16367,N_16368,N_16369,N_16370,N_16371,N_16372,N_16373,N_16374,N_16375,N_16376,N_16377,N_16378,N_16379,N_16380,N_16381,N_16382,N_16383,N_16384,N_16385,N_16386,N_16387,N_16388,N_16389,N_16390,N_16391,N_16392,N_16393,N_16394,N_16395,N_16396,N_16397,N_16398,N_16399,N_16400,N_16401,N_16402,N_16403,N_16404,N_16405,N_16406,N_16407,N_16408,N_16409,N_16410,N_16411,N_16412,N_16413,N_16414,N_16415,N_16416,N_16417,N_16418,N_16419,N_16420,N_16421,N_16422,N_16423,N_16424,N_16425,N_16426,N_16427,N_16428,N_16429,N_16430,N_16431,N_16432,N_16433,N_16434,N_16435,N_16436,N_16437,N_16438,N_16439,N_16440,N_16441,N_16442,N_16443,N_16444,N_16445,N_16446,N_16447,N_16448,N_16449,N_16450,N_16451,N_16452,N_16453,N_16454,N_16455,N_16456,N_16457,N_16458,N_16459,N_16460,N_16461,N_16462,N_16463,N_16464,N_16465,N_16466,N_16467,N_16468,N_16469,N_16470,N_16471,N_16472,N_16473,N_16474,N_16475,N_16476,N_16477,N_16478,N_16479,N_16480,N_16481,N_16482,N_16483,N_16484,N_16485,N_16486,N_16487,N_16488,N_16489,N_16490,N_16491,N_16492,N_16493,N_16494,N_16495,N_16496,N_16497,N_16498,N_16499,N_16500,N_16501,N_16502,N_16503,N_16504,N_16505,N_16506,N_16507,N_16508,N_16509,N_16510,N_16511,N_16512,N_16513,N_16514,N_16515,N_16516,N_16517,N_16518,N_16519,N_16520,N_16521,N_16522,N_16523,N_16524,N_16525,N_16526,N_16527,N_16528,N_16529,N_16530,N_16531,N_16532,N_16533,N_16534,N_16535,N_16536,N_16537,N_16538,N_16539,N_16540,N_16541,N_16542,N_16543,N_16544,N_16545,N_16546,N_16547,N_16548,N_16549,N_16550,N_16551,N_16552,N_16553,N_16554,N_16555,N_16556,N_16557,N_16558,N_16559,N_16560,N_16561,N_16562,N_16563,N_16564,N_16565,N_16566,N_16567,N_16568,N_16569,N_16570,N_16571,N_16572,N_16573,N_16574,N_16575,N_16576,N_16577,N_16578,N_16579,N_16580,N_16581,N_16582,N_16583,N_16584,N_16585,N_16586,N_16587,N_16588,N_16589,N_16590,N_16591,N_16592,N_16593,N_16594,N_16595,N_16596,N_16597,N_16598,N_16599,N_16600,N_16601,N_16602,N_16603,N_16604,N_16605,N_16606,N_16607,N_16608,N_16609,N_16610,N_16611,N_16612,N_16613,N_16614,N_16615,N_16616,N_16617,N_16618,N_16619,N_16620,N_16621,N_16622,N_16623,N_16624,N_16625,N_16626,N_16627,N_16628,N_16629,N_16630,N_16631,N_16632,N_16633,N_16634,N_16635,N_16636,N_16637,N_16638,N_16639,N_16640,N_16641,N_16642,N_16643,N_16644,N_16645,N_16646,N_16647,N_16648,N_16649,N_16650,N_16651,N_16652,N_16653,N_16654,N_16655,N_16656,N_16657,N_16658,N_16659,N_16660,N_16661,N_16662,N_16663,N_16664,N_16665,N_16666,N_16667,N_16668,N_16669,N_16670,N_16671,N_16672,N_16673,N_16674,N_16675,N_16676,N_16677,N_16678,N_16679,N_16680,N_16681,N_16682,N_16683,N_16684,N_16685,N_16686,N_16687,N_16688,N_16689,N_16690,N_16691,N_16692,N_16693,N_16694,N_16695,N_16696,N_16697,N_16698,N_16699,N_16700,N_16701,N_16702,N_16703,N_16704,N_16705,N_16706,N_16707,N_16708,N_16709,N_16710,N_16711,N_16712,N_16713,N_16714,N_16715,N_16716,N_16717,N_16718,N_16719,N_16720,N_16721,N_16722,N_16723,N_16724,N_16725,N_16726,N_16727,N_16728,N_16729,N_16730,N_16731,N_16732,N_16733,N_16734,N_16735,N_16736,N_16737,N_16738,N_16739,N_16740,N_16741,N_16742,N_16743,N_16744,N_16745,N_16746,N_16747,N_16748,N_16749,N_16750,N_16751,N_16752,N_16753,N_16754,N_16755,N_16756,N_16757,N_16758,N_16759,N_16760,N_16761,N_16762,N_16763,N_16764,N_16765,N_16766,N_16767,N_16768,N_16769,N_16770,N_16771,N_16772,N_16773,N_16774,N_16775,N_16776,N_16777,N_16778,N_16779,N_16780,N_16781,N_16782,N_16783,N_16784,N_16785,N_16786,N_16787,N_16788,N_16789,N_16790,N_16791,N_16792,N_16793,N_16794,N_16795,N_16796,N_16797,N_16798,N_16799,N_16800,N_16801,N_16802,N_16803,N_16804,N_16805,N_16806,N_16807,N_16808,N_16809,N_16810,N_16811,N_16812,N_16813,N_16814,N_16815,N_16816,N_16817,N_16818,N_16819,N_16820,N_16821,N_16822,N_16823,N_16824,N_16825,N_16826,N_16827,N_16828,N_16829,N_16830,N_16831,N_16832,N_16833,N_16834,N_16835,N_16836,N_16837,N_16838,N_16839,N_16840,N_16841,N_16842,N_16843,N_16844,N_16845,N_16846,N_16847,N_16848,N_16849,N_16850,N_16851,N_16852,N_16853,N_16854,N_16855,N_16856,N_16857,N_16858,N_16859,N_16860,N_16861,N_16862,N_16863,N_16864,N_16865,N_16866,N_16867,N_16868,N_16869,N_16870,N_16871,N_16872,N_16873,N_16874,N_16875,N_16876,N_16877,N_16878,N_16879,N_16880,N_16881,N_16882,N_16883,N_16884,N_16885,N_16886,N_16887,N_16888,N_16889,N_16890,N_16891,N_16892,N_16893,N_16894,N_16895,N_16896,N_16897,N_16898,N_16899,N_16900,N_16901,N_16902,N_16903,N_16904,N_16905,N_16906,N_16907,N_16908,N_16909,N_16910,N_16911,N_16912,N_16913,N_16914,N_16915,N_16916,N_16917,N_16918,N_16919,N_16920,N_16921,N_16922,N_16923,N_16924,N_16925,N_16926,N_16927,N_16928,N_16929,N_16930,N_16931,N_16932,N_16933,N_16934,N_16935,N_16936,N_16937,N_16938,N_16939,N_16940,N_16941,N_16942,N_16943,N_16944,N_16945,N_16946,N_16947,N_16948,N_16949,N_16950,N_16951,N_16952,N_16953,N_16954,N_16955,N_16956,N_16957,N_16958,N_16959,N_16960,N_16961,N_16962,N_16963,N_16964,N_16965,N_16966,N_16967,N_16968,N_16969,N_16970,N_16971,N_16972,N_16973,N_16974,N_16975,N_16976,N_16977,N_16978,N_16979,N_16980,N_16981,N_16982,N_16983,N_16984,N_16985,N_16986,N_16987,N_16988,N_16989,N_16990,N_16991,N_16992,N_16993,N_16994,N_16995,N_16996,N_16997,N_16998,N_16999,N_17000,N_17001,N_17002,N_17003,N_17004,N_17005,N_17006,N_17007,N_17008,N_17009,N_17010,N_17011,N_17012,N_17013,N_17014,N_17015,N_17016,N_17017,N_17018,N_17019,N_17020,N_17021,N_17022,N_17023,N_17024,N_17025,N_17026,N_17027,N_17028,N_17029,N_17030,N_17031,N_17032,N_17033,N_17034,N_17035,N_17036,N_17037,N_17038,N_17039,N_17040,N_17041,N_17042,N_17043,N_17044,N_17045,N_17046,N_17047,N_17048,N_17049,N_17050,N_17051,N_17052,N_17053,N_17054,N_17055,N_17056,N_17057,N_17058,N_17059,N_17060,N_17061,N_17062,N_17063,N_17064,N_17065,N_17066,N_17067,N_17068,N_17069,N_17070,N_17071,N_17072,N_17073,N_17074,N_17075,N_17076,N_17077,N_17078,N_17079,N_17080,N_17081,N_17082,N_17083,N_17084,N_17085,N_17086,N_17087,N_17088,N_17089,N_17090,N_17091,N_17092,N_17093,N_17094,N_17095,N_17096,N_17097,N_17098,N_17099,N_17100,N_17101,N_17102,N_17103,N_17104,N_17105,N_17106,N_17107,N_17108,N_17109,N_17110,N_17111,N_17112,N_17113,N_17114,N_17115,N_17116,N_17117,N_17118,N_17119,N_17120,N_17121,N_17122,N_17123,N_17124,N_17125,N_17126,N_17127,N_17128,N_17129,N_17130,N_17131,N_17132,N_17133,N_17134,N_17135,N_17136,N_17137,N_17138,N_17139,N_17140,N_17141,N_17142,N_17143,N_17144,N_17145,N_17146,N_17147,N_17148,N_17149,N_17150,N_17151,N_17152,N_17153,N_17154,N_17155,N_17156,N_17157,N_17158,N_17159,N_17160,N_17161,N_17162,N_17163,N_17164,N_17165,N_17166,N_17167,N_17168,N_17169,N_17170,N_17171,N_17172,N_17173,N_17174,N_17175,N_17176,N_17177,N_17178,N_17179,N_17180,N_17181,N_17182,N_17183,N_17184,N_17185,N_17186,N_17187,N_17188,N_17189,N_17190,N_17191,N_17192,N_17193,N_17194,N_17195,N_17196,N_17197,N_17198,N_17199,N_17200,N_17201,N_17202,N_17203,N_17204,N_17205,N_17206,N_17207,N_17208,N_17209,N_17210,N_17211,N_17212,N_17213,N_17214,N_17215,N_17216,N_17217,N_17218,N_17219,N_17220,N_17221,N_17222,N_17223,N_17224,N_17225,N_17226,N_17227,N_17228,N_17229,N_17230,N_17231,N_17232,N_17233,N_17234,N_17235,N_17236,N_17237,N_17238,N_17239,N_17240,N_17241,N_17242,N_17243,N_17244,N_17245,N_17246,N_17247,N_17248,N_17249,N_17250,N_17251,N_17252,N_17253,N_17254,N_17255,N_17256,N_17257,N_17258,N_17259,N_17260,N_17261,N_17262,N_17263,N_17264,N_17265,N_17266,N_17267,N_17268,N_17269,N_17270,N_17271,N_17272,N_17273,N_17274,N_17275,N_17276,N_17277,N_17278,N_17279,N_17280,N_17281,N_17282,N_17283,N_17284,N_17285,N_17286,N_17287,N_17288,N_17289,N_17290,N_17291,N_17292,N_17293,N_17294,N_17295,N_17296,N_17297,N_17298,N_17299,N_17300,N_17301,N_17302,N_17303,N_17304,N_17305,N_17306,N_17307,N_17308,N_17309,N_17310,N_17311,N_17312,N_17313,N_17314,N_17315,N_17316,N_17317,N_17318,N_17319,N_17320,N_17321,N_17322,N_17323,N_17324,N_17325,N_17326,N_17327,N_17328,N_17329,N_17330,N_17331,N_17332,N_17333,N_17334,N_17335,N_17336,N_17337,N_17338,N_17339,N_17340,N_17341,N_17342,N_17343,N_17344,N_17345,N_17346,N_17347,N_17348,N_17349,N_17350,N_17351,N_17352,N_17353,N_17354,N_17355,N_17356,N_17357,N_17358,N_17359,N_17360,N_17361,N_17362,N_17363,N_17364,N_17365,N_17366,N_17367,N_17368,N_17369,N_17370,N_17371,N_17372,N_17373,N_17374,N_17375,N_17376,N_17377,N_17378,N_17379,N_17380,N_17381,N_17382,N_17383,N_17384,N_17385,N_17386,N_17387,N_17388,N_17389,N_17390,N_17391,N_17392,N_17393,N_17394,N_17395,N_17396,N_17397,N_17398,N_17399,N_17400,N_17401,N_17402,N_17403,N_17404,N_17405,N_17406,N_17407,N_17408,N_17409,N_17410,N_17411,N_17412,N_17413,N_17414,N_17415,N_17416,N_17417,N_17418,N_17419,N_17420,N_17421,N_17422,N_17423,N_17424,N_17425,N_17426,N_17427,N_17428,N_17429,N_17430,N_17431,N_17432,N_17433,N_17434,N_17435,N_17436,N_17437,N_17438,N_17439,N_17440,N_17441,N_17442,N_17443,N_17444,N_17445,N_17446,N_17447,N_17448,N_17449,N_17450,N_17451,N_17452,N_17453,N_17454,N_17455,N_17456,N_17457,N_17458,N_17459,N_17460,N_17461,N_17462,N_17463,N_17464,N_17465,N_17466,N_17467,N_17468,N_17469,N_17470,N_17471,N_17472,N_17473,N_17474,N_17475,N_17476,N_17477,N_17478,N_17479,N_17480,N_17481,N_17482,N_17483,N_17484,N_17485,N_17486,N_17487,N_17488,N_17489,N_17490,N_17491,N_17492,N_17493,N_17494,N_17495,N_17496,N_17497,N_17498,N_17499,N_17500,N_17501,N_17502,N_17503,N_17504,N_17505,N_17506,N_17507,N_17508,N_17509,N_17510,N_17511,N_17512,N_17513,N_17514,N_17515,N_17516,N_17517,N_17518,N_17519,N_17520,N_17521,N_17522,N_17523,N_17524,N_17525,N_17526,N_17527,N_17528,N_17529,N_17530,N_17531,N_17532,N_17533,N_17534,N_17535,N_17536,N_17537,N_17538,N_17539,N_17540,N_17541,N_17542,N_17543,N_17544,N_17545,N_17546,N_17547,N_17548,N_17549,N_17550,N_17551,N_17552,N_17553,N_17554,N_17555,N_17556,N_17557,N_17558,N_17559,N_17560,N_17561,N_17562,N_17563,N_17564,N_17565,N_17566,N_17567,N_17568,N_17569,N_17570,N_17571,N_17572,N_17573,N_17574,N_17575,N_17576,N_17577,N_17578,N_17579,N_17580,N_17581,N_17582,N_17583,N_17584,N_17585,N_17586,N_17587,N_17588,N_17589,N_17590,N_17591,N_17592,N_17593,N_17594,N_17595,N_17596,N_17597,N_17598,N_17599,N_17600,N_17601,N_17602,N_17603,N_17604,N_17605,N_17606,N_17607,N_17608,N_17609,N_17610,N_17611,N_17612,N_17613,N_17614,N_17615,N_17616,N_17617,N_17618,N_17619,N_17620,N_17621,N_17622,N_17623,N_17624,N_17625,N_17626,N_17627,N_17628,N_17629,N_17630,N_17631,N_17632,N_17633,N_17634,N_17635,N_17636,N_17637,N_17638,N_17639,N_17640,N_17641,N_17642,N_17643,N_17644,N_17645,N_17646,N_17647,N_17648,N_17649,N_17650,N_17651,N_17652,N_17653,N_17654,N_17655,N_17656,N_17657,N_17658,N_17659,N_17660,N_17661,N_17662,N_17663,N_17664,N_17665,N_17666,N_17667,N_17668,N_17669,N_17670,N_17671,N_17672,N_17673,N_17674,N_17675,N_17676,N_17677,N_17678,N_17679,N_17680,N_17681,N_17682,N_17683,N_17684,N_17685,N_17686,N_17687,N_17688,N_17689,N_17690,N_17691,N_17692,N_17693,N_17694,N_17695,N_17696,N_17697,N_17698,N_17699,N_17700,N_17701,N_17702,N_17703,N_17704,N_17705,N_17706,N_17707,N_17708,N_17709,N_17710,N_17711,N_17712,N_17713,N_17714,N_17715,N_17716,N_17717,N_17718,N_17719,N_17720,N_17721,N_17722,N_17723,N_17724,N_17725,N_17726,N_17727,N_17728,N_17729,N_17730,N_17731,N_17732,N_17733,N_17734,N_17735,N_17736,N_17737,N_17738,N_17739,N_17740,N_17741,N_17742,N_17743,N_17744,N_17745,N_17746,N_17747,N_17748,N_17749,N_17750,N_17751,N_17752,N_17753,N_17754,N_17755,N_17756,N_17757,N_17758,N_17759,N_17760,N_17761,N_17762,N_17763,N_17764,N_17765,N_17766,N_17767,N_17768,N_17769,N_17770,N_17771,N_17772,N_17773,N_17774,N_17775,N_17776,N_17777,N_17778,N_17779,N_17780,N_17781,N_17782,N_17783,N_17784,N_17785,N_17786,N_17787,N_17788,N_17789,N_17790,N_17791,N_17792,N_17793,N_17794,N_17795,N_17796,N_17797,N_17798,N_17799,N_17800,N_17801,N_17802,N_17803,N_17804,N_17805,N_17806,N_17807,N_17808,N_17809,N_17810,N_17811,N_17812,N_17813,N_17814,N_17815,N_17816,N_17817,N_17818,N_17819,N_17820,N_17821,N_17822,N_17823,N_17824,N_17825,N_17826,N_17827,N_17828,N_17829,N_17830,N_17831,N_17832,N_17833,N_17834,N_17835,N_17836,N_17837,N_17838,N_17839,N_17840,N_17841,N_17842,N_17843,N_17844,N_17845,N_17846,N_17847,N_17848,N_17849,N_17850,N_17851,N_17852,N_17853,N_17854,N_17855,N_17856,N_17857,N_17858,N_17859,N_17860,N_17861,N_17862,N_17863,N_17864,N_17865,N_17866,N_17867,N_17868,N_17869,N_17870,N_17871,N_17872,N_17873,N_17874,N_17875,N_17876,N_17877,N_17878,N_17879,N_17880,N_17881,N_17882,N_17883,N_17884,N_17885,N_17886,N_17887,N_17888,N_17889,N_17890,N_17891,N_17892,N_17893,N_17894,N_17895,N_17896,N_17897,N_17898,N_17899,N_17900,N_17901,N_17902,N_17903,N_17904,N_17905,N_17906,N_17907,N_17908,N_17909,N_17910,N_17911,N_17912,N_17913,N_17914,N_17915,N_17916,N_17917,N_17918,N_17919,N_17920,N_17921,N_17922,N_17923,N_17924,N_17925,N_17926,N_17927,N_17928,N_17929,N_17930,N_17931,N_17932,N_17933,N_17934,N_17935,N_17936,N_17937,N_17938,N_17939,N_17940,N_17941,N_17942,N_17943,N_17944,N_17945,N_17946,N_17947,N_17948,N_17949,N_17950,N_17951,N_17952,N_17953,N_17954,N_17955,N_17956,N_17957,N_17958,N_17959,N_17960,N_17961,N_17962,N_17963,N_17964,N_17965,N_17966,N_17967,N_17968,N_17969,N_17970,N_17971,N_17972,N_17973,N_17974,N_17975,N_17976,N_17977,N_17978,N_17979,N_17980,N_17981,N_17982,N_17983,N_17984,N_17985,N_17986,N_17987,N_17988,N_17989,N_17990,N_17991,N_17992,N_17993,N_17994,N_17995,N_17996,N_17997,N_17998,N_17999,N_18000,N_18001,N_18002,N_18003,N_18004,N_18005,N_18006,N_18007,N_18008,N_18009,N_18010,N_18011,N_18012,N_18013,N_18014,N_18015,N_18016,N_18017,N_18018,N_18019,N_18020,N_18021,N_18022,N_18023,N_18024,N_18025,N_18026,N_18027,N_18028,N_18029,N_18030,N_18031,N_18032,N_18033,N_18034,N_18035,N_18036,N_18037,N_18038,N_18039,N_18040,N_18041,N_18042,N_18043,N_18044,N_18045,N_18046,N_18047,N_18048,N_18049,N_18050,N_18051,N_18052,N_18053,N_18054,N_18055,N_18056,N_18057,N_18058,N_18059,N_18060,N_18061,N_18062,N_18063,N_18064,N_18065,N_18066,N_18067,N_18068,N_18069,N_18070,N_18071,N_18072,N_18073,N_18074,N_18075,N_18076,N_18077,N_18078,N_18079,N_18080,N_18081,N_18082,N_18083,N_18084,N_18085,N_18086,N_18087,N_18088,N_18089,N_18090,N_18091,N_18092,N_18093,N_18094,N_18095,N_18096,N_18097,N_18098,N_18099,N_18100,N_18101,N_18102,N_18103,N_18104,N_18105,N_18106,N_18107,N_18108,N_18109,N_18110,N_18111,N_18112,N_18113,N_18114,N_18115,N_18116,N_18117,N_18118,N_18119,N_18120,N_18121,N_18122,N_18123,N_18124,N_18125,N_18126,N_18127,N_18128,N_18129,N_18130,N_18131,N_18132,N_18133,N_18134,N_18135,N_18136,N_18137,N_18138,N_18139,N_18140,N_18141,N_18142,N_18143,N_18144,N_18145,N_18146,N_18147,N_18148,N_18149,N_18150,N_18151,N_18152,N_18153,N_18154,N_18155,N_18156,N_18157,N_18158,N_18159,N_18160,N_18161,N_18162,N_18163,N_18164,N_18165,N_18166,N_18167,N_18168,N_18169,N_18170,N_18171,N_18172,N_18173,N_18174,N_18175,N_18176,N_18177,N_18178,N_18179,N_18180,N_18181,N_18182,N_18183,N_18184,N_18185,N_18186,N_18187,N_18188,N_18189,N_18190,N_18191,N_18192,N_18193,N_18194,N_18195,N_18196,N_18197,N_18198,N_18199,N_18200,N_18201,N_18202,N_18203,N_18204,N_18205,N_18206,N_18207,N_18208,N_18209,N_18210,N_18211,N_18212,N_18213,N_18214,N_18215,N_18216,N_18217,N_18218,N_18219,N_18220,N_18221,N_18222,N_18223,N_18224,N_18225,N_18226,N_18227,N_18228,N_18229,N_18230,N_18231,N_18232,N_18233,N_18234,N_18235,N_18236,N_18237,N_18238,N_18239,N_18240,N_18241,N_18242,N_18243,N_18244,N_18245,N_18246,N_18247,N_18248,N_18249,N_18250,N_18251,N_18252,N_18253,N_18254,N_18255,N_18256,N_18257,N_18258,N_18259,N_18260,N_18261,N_18262,N_18263,N_18264,N_18265,N_18266,N_18267,N_18268,N_18269,N_18270,N_18271,N_18272,N_18273,N_18274,N_18275,N_18276,N_18277,N_18278,N_18279,N_18280,N_18281,N_18282,N_18283,N_18284,N_18285,N_18286,N_18287,N_18288,N_18289,N_18290,N_18291,N_18292,N_18293,N_18294,N_18295,N_18296,N_18297,N_18298,N_18299,N_18300,N_18301,N_18302,N_18303,N_18304,N_18305,N_18306,N_18307,N_18308,N_18309,N_18310,N_18311,N_18312,N_18313,N_18314,N_18315,N_18316,N_18317,N_18318,N_18319,N_18320,N_18321,N_18322,N_18323,N_18324,N_18325,N_18326,N_18327,N_18328,N_18329,N_18330,N_18331,N_18332,N_18333,N_18334,N_18335,N_18336,N_18337,N_18338,N_18339,N_18340,N_18341,N_18342,N_18343,N_18344,N_18345,N_18346,N_18347,N_18348,N_18349,N_18350,N_18351,N_18352,N_18353,N_18354,N_18355,N_18356,N_18357,N_18358,N_18359,N_18360,N_18361,N_18362,N_18363,N_18364,N_18365,N_18366,N_18367,N_18368,N_18369,N_18370,N_18371,N_18372,N_18373,N_18374,N_18375,N_18376,N_18377,N_18378,N_18379,N_18380,N_18381,N_18382,N_18383,N_18384,N_18385,N_18386,N_18387,N_18388,N_18389,N_18390,N_18391,N_18392,N_18393,N_18394,N_18395,N_18396,N_18397,N_18398,N_18399,N_18400,N_18401,N_18402,N_18403,N_18404,N_18405,N_18406,N_18407,N_18408,N_18409,N_18410,N_18411,N_18412,N_18413,N_18414,N_18415,N_18416,N_18417,N_18418,N_18419,N_18420,N_18421,N_18422,N_18423,N_18424,N_18425,N_18426,N_18427,N_18428,N_18429,N_18430,N_18431,N_18432,N_18433,N_18434,N_18435,N_18436,N_18437,N_18438,N_18439,N_18440,N_18441,N_18442,N_18443,N_18444,N_18445,N_18446,N_18447,N_18448,N_18449,N_18450,N_18451,N_18452,N_18453,N_18454,N_18455,N_18456,N_18457,N_18458,N_18459,N_18460,N_18461,N_18462,N_18463,N_18464,N_18465,N_18466,N_18467,N_18468,N_18469,N_18470,N_18471,N_18472,N_18473,N_18474,N_18475,N_18476,N_18477,N_18478,N_18479,N_18480,N_18481,N_18482,N_18483,N_18484,N_18485,N_18486,N_18487,N_18488,N_18489,N_18490,N_18491,N_18492,N_18493,N_18494,N_18495,N_18496,N_18497,N_18498,N_18499,N_18500,N_18501,N_18502,N_18503,N_18504,N_18505,N_18506,N_18507,N_18508,N_18509,N_18510,N_18511,N_18512,N_18513,N_18514,N_18515,N_18516,N_18517,N_18518,N_18519,N_18520,N_18521,N_18522,N_18523,N_18524,N_18525,N_18526,N_18527,N_18528,N_18529,N_18530,N_18531,N_18532,N_18533,N_18534,N_18535,N_18536,N_18537,N_18538,N_18539,N_18540,N_18541,N_18542,N_18543,N_18544,N_18545,N_18546,N_18547,N_18548,N_18549,N_18550,N_18551,N_18552,N_18553,N_18554,N_18555,N_18556,N_18557,N_18558,N_18559,N_18560,N_18561,N_18562,N_18563,N_18564,N_18565,N_18566,N_18567,N_18568,N_18569,N_18570,N_18571,N_18572,N_18573,N_18574,N_18575,N_18576,N_18577,N_18578,N_18579,N_18580,N_18581,N_18582,N_18583,N_18584,N_18585,N_18586,N_18587,N_18588,N_18589,N_18590,N_18591,N_18592,N_18593,N_18594,N_18595,N_18596,N_18597,N_18598,N_18599,N_18600,N_18601,N_18602,N_18603,N_18604,N_18605,N_18606,N_18607,N_18608,N_18609,N_18610,N_18611,N_18612,N_18613,N_18614,N_18615,N_18616,N_18617,N_18618,N_18619,N_18620,N_18621,N_18622,N_18623,N_18624,N_18625,N_18626,N_18627,N_18628,N_18629,N_18630,N_18631,N_18632,N_18633,N_18634,N_18635,N_18636,N_18637,N_18638,N_18639,N_18640,N_18641,N_18642,N_18643,N_18644,N_18645,N_18646,N_18647,N_18648,N_18649,N_18650,N_18651,N_18652,N_18653,N_18654,N_18655,N_18656,N_18657,N_18658,N_18659,N_18660,N_18661,N_18662,N_18663,N_18664,N_18665,N_18666,N_18667,N_18668,N_18669,N_18670,N_18671,N_18672,N_18673,N_18674,N_18675,N_18676,N_18677,N_18678,N_18679,N_18680,N_18681,N_18682,N_18683,N_18684,N_18685,N_18686,N_18687,N_18688,N_18689,N_18690,N_18691,N_18692,N_18693,N_18694,N_18695,N_18696,N_18697,N_18698,N_18699,N_18700,N_18701,N_18702,N_18703,N_18704,N_18705,N_18706,N_18707,N_18708,N_18709,N_18710,N_18711,N_18712,N_18713,N_18714,N_18715,N_18716,N_18717,N_18718,N_18719,N_18720,N_18721,N_18722,N_18723,N_18724,N_18725,N_18726,N_18727,N_18728,N_18729,N_18730,N_18731,N_18732,N_18733,N_18734,N_18735,N_18736,N_18737,N_18738,N_18739,N_18740,N_18741,N_18742,N_18743,N_18744,N_18745,N_18746,N_18747,N_18748,N_18749,N_18750,N_18751,N_18752,N_18753,N_18754,N_18755,N_18756,N_18757,N_18758,N_18759,N_18760,N_18761,N_18762,N_18763,N_18764,N_18765,N_18766,N_18767,N_18768,N_18769,N_18770,N_18771,N_18772,N_18773,N_18774,N_18775,N_18776,N_18777,N_18778,N_18779,N_18780,N_18781,N_18782,N_18783,N_18784,N_18785,N_18786,N_18787,N_18788,N_18789,N_18790,N_18791,N_18792,N_18793,N_18794,N_18795,N_18796,N_18797,N_18798,N_18799,N_18800,N_18801,N_18802,N_18803,N_18804,N_18805,N_18806,N_18807,N_18808,N_18809,N_18810,N_18811,N_18812,N_18813,N_18814,N_18815,N_18816,N_18817,N_18818,N_18819,N_18820,N_18821,N_18822,N_18823,N_18824,N_18825,N_18826,N_18827,N_18828,N_18829,N_18830,N_18831,N_18832,N_18833,N_18834,N_18835,N_18836,N_18837,N_18838,N_18839,N_18840,N_18841,N_18842,N_18843,N_18844,N_18845,N_18846,N_18847,N_18848,N_18849,N_18850,N_18851,N_18852,N_18853,N_18854,N_18855,N_18856,N_18857,N_18858,N_18859,N_18860,N_18861,N_18862,N_18863,N_18864,N_18865,N_18866,N_18867,N_18868,N_18869,N_18870,N_18871,N_18872,N_18873,N_18874,N_18875,N_18876,N_18877,N_18878,N_18879,N_18880,N_18881,N_18882,N_18883,N_18884,N_18885,N_18886,N_18887,N_18888,N_18889,N_18890,N_18891,N_18892,N_18893,N_18894,N_18895,N_18896,N_18897,N_18898,N_18899,N_18900,N_18901,N_18902,N_18903,N_18904,N_18905,N_18906,N_18907,N_18908,N_18909,N_18910,N_18911,N_18912,N_18913,N_18914,N_18915,N_18916,N_18917,N_18918,N_18919,N_18920,N_18921,N_18922,N_18923,N_18924,N_18925,N_18926,N_18927,N_18928,N_18929,N_18930,N_18931,N_18932,N_18933,N_18934,N_18935,N_18936,N_18937,N_18938,N_18939,N_18940,N_18941,N_18942,N_18943,N_18944,N_18945,N_18946,N_18947,N_18948,N_18949,N_18950,N_18951,N_18952,N_18953,N_18954,N_18955,N_18956,N_18957,N_18958,N_18959,N_18960,N_18961,N_18962,N_18963,N_18964,N_18965,N_18966,N_18967,N_18968,N_18969,N_18970,N_18971,N_18972,N_18973,N_18974,N_18975,N_18976,N_18977,N_18978,N_18979,N_18980,N_18981,N_18982,N_18983,N_18984,N_18985,N_18986,N_18987,N_18988,N_18989,N_18990,N_18991,N_18992,N_18993,N_18994,N_18995,N_18996,N_18997,N_18998,N_18999,N_19000,N_19001,N_19002,N_19003,N_19004,N_19005,N_19006,N_19007,N_19008,N_19009,N_19010,N_19011,N_19012,N_19013,N_19014,N_19015,N_19016,N_19017,N_19018,N_19019,N_19020,N_19021,N_19022,N_19023,N_19024,N_19025,N_19026,N_19027,N_19028,N_19029,N_19030,N_19031,N_19032,N_19033,N_19034,N_19035,N_19036,N_19037,N_19038,N_19039,N_19040,N_19041,N_19042,N_19043,N_19044,N_19045,N_19046,N_19047,N_19048,N_19049,N_19050,N_19051,N_19052,N_19053,N_19054,N_19055,N_19056,N_19057,N_19058,N_19059,N_19060,N_19061,N_19062,N_19063,N_19064,N_19065,N_19066,N_19067,N_19068,N_19069,N_19070,N_19071,N_19072,N_19073,N_19074,N_19075,N_19076,N_19077,N_19078,N_19079,N_19080,N_19081,N_19082,N_19083,N_19084,N_19085,N_19086,N_19087,N_19088,N_19089,N_19090,N_19091,N_19092,N_19093,N_19094,N_19095,N_19096,N_19097,N_19098,N_19099,N_19100,N_19101,N_19102,N_19103,N_19104,N_19105,N_19106,N_19107,N_19108,N_19109,N_19110,N_19111,N_19112,N_19113,N_19114,N_19115,N_19116,N_19117,N_19118,N_19119,N_19120,N_19121,N_19122,N_19123,N_19124,N_19125,N_19126,N_19127,N_19128,N_19129,N_19130,N_19131,N_19132,N_19133,N_19134,N_19135,N_19136,N_19137,N_19138,N_19139,N_19140,N_19141,N_19142,N_19143,N_19144,N_19145,N_19146,N_19147,N_19148,N_19149,N_19150,N_19151,N_19152,N_19153,N_19154,N_19155,N_19156,N_19157,N_19158,N_19159,N_19160,N_19161,N_19162,N_19163,N_19164,N_19165,N_19166,N_19167,N_19168,N_19169,N_19170,N_19171,N_19172,N_19173,N_19174,N_19175,N_19176,N_19177,N_19178,N_19179,N_19180,N_19181,N_19182,N_19183,N_19184,N_19185,N_19186,N_19187,N_19188,N_19189,N_19190,N_19191,N_19192,N_19193,N_19194,N_19195,N_19196,N_19197,N_19198,N_19199,N_19200,N_19201,N_19202,N_19203,N_19204,N_19205,N_19206,N_19207,N_19208,N_19209,N_19210,N_19211,N_19212,N_19213,N_19214,N_19215,N_19216,N_19217,N_19218,N_19219,N_19220,N_19221,N_19222,N_19223,N_19224,N_19225,N_19226,N_19227,N_19228,N_19229,N_19230,N_19231,N_19232,N_19233,N_19234,N_19235,N_19236,N_19237,N_19238,N_19239,N_19240,N_19241,N_19242,N_19243,N_19244,N_19245,N_19246,N_19247,N_19248,N_19249,N_19250,N_19251,N_19252,N_19253,N_19254,N_19255,N_19256,N_19257,N_19258,N_19259,N_19260,N_19261,N_19262,N_19263,N_19264,N_19265,N_19266,N_19267,N_19268,N_19269,N_19270,N_19271,N_19272,N_19273,N_19274,N_19275,N_19276,N_19277,N_19278,N_19279,N_19280,N_19281,N_19282,N_19283,N_19284,N_19285,N_19286,N_19287,N_19288,N_19289,N_19290,N_19291,N_19292,N_19293,N_19294,N_19295,N_19296,N_19297,N_19298,N_19299,N_19300,N_19301,N_19302,N_19303,N_19304,N_19305,N_19306,N_19307,N_19308,N_19309,N_19310,N_19311,N_19312,N_19313,N_19314,N_19315,N_19316,N_19317,N_19318,N_19319,N_19320,N_19321,N_19322,N_19323,N_19324,N_19325,N_19326,N_19327,N_19328,N_19329,N_19330,N_19331,N_19332,N_19333,N_19334,N_19335,N_19336,N_19337,N_19338,N_19339,N_19340,N_19341,N_19342,N_19343,N_19344,N_19345,N_19346,N_19347,N_19348,N_19349,N_19350,N_19351,N_19352,N_19353,N_19354,N_19355,N_19356,N_19357,N_19358,N_19359,N_19360,N_19361,N_19362,N_19363,N_19364,N_19365,N_19366,N_19367,N_19368,N_19369,N_19370,N_19371,N_19372,N_19373,N_19374,N_19375,N_19376,N_19377,N_19378,N_19379,N_19380,N_19381,N_19382,N_19383,N_19384,N_19385,N_19386,N_19387,N_19388,N_19389,N_19390,N_19391,N_19392,N_19393,N_19394,N_19395,N_19396,N_19397,N_19398,N_19399,N_19400,N_19401,N_19402,N_19403,N_19404,N_19405,N_19406,N_19407,N_19408,N_19409,N_19410,N_19411,N_19412,N_19413,N_19414,N_19415,N_19416,N_19417,N_19418,N_19419,N_19420,N_19421,N_19422,N_19423,N_19424,N_19425,N_19426,N_19427,N_19428,N_19429,N_19430,N_19431,N_19432,N_19433,N_19434,N_19435,N_19436,N_19437,N_19438,N_19439,N_19440,N_19441,N_19442,N_19443,N_19444,N_19445,N_19446,N_19447,N_19448,N_19449,N_19450,N_19451,N_19452,N_19453,N_19454,N_19455,N_19456,N_19457,N_19458,N_19459,N_19460,N_19461,N_19462,N_19463,N_19464,N_19465,N_19466,N_19467,N_19468,N_19469,N_19470,N_19471,N_19472,N_19473,N_19474,N_19475,N_19476,N_19477,N_19478,N_19479,N_19480,N_19481,N_19482,N_19483,N_19484,N_19485,N_19486,N_19487,N_19488,N_19489,N_19490,N_19491,N_19492,N_19493,N_19494,N_19495,N_19496,N_19497,N_19498,N_19499,N_19500,N_19501,N_19502,N_19503,N_19504,N_19505,N_19506,N_19507,N_19508,N_19509,N_19510,N_19511,N_19512,N_19513,N_19514,N_19515,N_19516,N_19517,N_19518,N_19519,N_19520,N_19521,N_19522,N_19523,N_19524,N_19525,N_19526,N_19527,N_19528,N_19529,N_19530,N_19531,N_19532,N_19533,N_19534,N_19535,N_19536,N_19537,N_19538,N_19539,N_19540,N_19541,N_19542,N_19543,N_19544,N_19545,N_19546,N_19547,N_19548,N_19549,N_19550,N_19551,N_19552,N_19553,N_19554,N_19555,N_19556,N_19557,N_19558,N_19559,N_19560,N_19561,N_19562,N_19563,N_19564,N_19565,N_19566,N_19567,N_19568,N_19569,N_19570,N_19571,N_19572,N_19573,N_19574,N_19575,N_19576,N_19577,N_19578,N_19579,N_19580,N_19581,N_19582,N_19583,N_19584,N_19585,N_19586,N_19587,N_19588,N_19589,N_19590,N_19591,N_19592,N_19593,N_19594,N_19595,N_19596,N_19597,N_19598,N_19599,N_19600,N_19601,N_19602,N_19603,N_19604,N_19605,N_19606,N_19607,N_19608,N_19609,N_19610,N_19611,N_19612,N_19613,N_19614,N_19615,N_19616,N_19617,N_19618,N_19619,N_19620,N_19621,N_19622,N_19623,N_19624,N_19625,N_19626,N_19627,N_19628,N_19629,N_19630,N_19631,N_19632,N_19633,N_19634,N_19635,N_19636,N_19637,N_19638,N_19639,N_19640,N_19641,N_19642,N_19643,N_19644,N_19645,N_19646,N_19647,N_19648,N_19649,N_19650,N_19651,N_19652,N_19653,N_19654,N_19655,N_19656,N_19657,N_19658,N_19659,N_19660,N_19661,N_19662,N_19663,N_19664,N_19665,N_19666,N_19667,N_19668,N_19669,N_19670,N_19671,N_19672,N_19673,N_19674,N_19675,N_19676,N_19677,N_19678,N_19679,N_19680,N_19681,N_19682,N_19683,N_19684,N_19685,N_19686,N_19687,N_19688,N_19689,N_19690,N_19691,N_19692,N_19693,N_19694,N_19695,N_19696,N_19697,N_19698,N_19699,N_19700,N_19701,N_19702,N_19703,N_19704,N_19705,N_19706,N_19707,N_19708,N_19709,N_19710,N_19711,N_19712,N_19713,N_19714,N_19715,N_19716,N_19717,N_19718,N_19719,N_19720,N_19721,N_19722,N_19723,N_19724,N_19725,N_19726,N_19727,N_19728,N_19729,N_19730,N_19731,N_19732,N_19733,N_19734,N_19735,N_19736,N_19737,N_19738,N_19739,N_19740,N_19741,N_19742,N_19743,N_19744,N_19745,N_19746,N_19747,N_19748,N_19749,N_19750,N_19751,N_19752,N_19753,N_19754,N_19755,N_19756,N_19757,N_19758,N_19759,N_19760,N_19761,N_19762,N_19763,N_19764,N_19765,N_19766,N_19767,N_19768,N_19769,N_19770,N_19771,N_19772,N_19773,N_19774,N_19775,N_19776,N_19777,N_19778,N_19779,N_19780,N_19781,N_19782,N_19783,N_19784,N_19785,N_19786,N_19787,N_19788,N_19789,N_19790,N_19791,N_19792,N_19793,N_19794,N_19795,N_19796,N_19797,N_19798,N_19799,N_19800,N_19801,N_19802,N_19803,N_19804,N_19805,N_19806,N_19807,N_19808,N_19809,N_19810,N_19811,N_19812,N_19813,N_19814,N_19815,N_19816,N_19817,N_19818,N_19819,N_19820,N_19821,N_19822,N_19823,N_19824,N_19825,N_19826,N_19827,N_19828,N_19829,N_19830,N_19831,N_19832,N_19833,N_19834,N_19835,N_19836,N_19837,N_19838,N_19839,N_19840,N_19841,N_19842,N_19843,N_19844,N_19845,N_19846,N_19847,N_19848,N_19849,N_19850,N_19851,N_19852,N_19853,N_19854,N_19855,N_19856,N_19857,N_19858,N_19859,N_19860,N_19861,N_19862,N_19863,N_19864,N_19865,N_19866,N_19867,N_19868,N_19869,N_19870,N_19871,N_19872,N_19873,N_19874,N_19875,N_19876,N_19877,N_19878,N_19879,N_19880,N_19881,N_19882,N_19883,N_19884,N_19885,N_19886,N_19887,N_19888,N_19889,N_19890,N_19891,N_19892,N_19893,N_19894,N_19895,N_19896,N_19897,N_19898,N_19899,N_19900,N_19901,N_19902,N_19903,N_19904,N_19905,N_19906,N_19907,N_19908,N_19909,N_19910,N_19911,N_19912,N_19913,N_19914,N_19915,N_19916,N_19917,N_19918,N_19919,N_19920,N_19921,N_19922,N_19923,N_19924,N_19925,N_19926,N_19927,N_19928,N_19929,N_19930,N_19931,N_19932,N_19933,N_19934,N_19935,N_19936,N_19937,N_19938,N_19939,N_19940,N_19941,N_19942,N_19943,N_19944,N_19945,N_19946,N_19947,N_19948,N_19949,N_19950,N_19951,N_19952,N_19953,N_19954,N_19955,N_19956,N_19957,N_19958,N_19959,N_19960,N_19961,N_19962,N_19963,N_19964,N_19965,N_19966,N_19967,N_19968,N_19969,N_19970,N_19971,N_19972,N_19973,N_19974,N_19975,N_19976,N_19977,N_19978,N_19979,N_19980,N_19981,N_19982,N_19983,N_19984,N_19985,N_19986,N_19987,N_19988,N_19989,N_19990,N_19991,N_19992,N_19993,N_19994,N_19995,N_19996,N_19997,N_19998,N_19999,N_20000,N_20001,N_20002,N_20003,N_20004,N_20005,N_20006,N_20007,N_20008,N_20009,N_20010,N_20011,N_20012,N_20013,N_20014,N_20015,N_20016,N_20017,N_20018,N_20019,N_20020,N_20021,N_20022,N_20023,N_20024,N_20025,N_20026,N_20027,N_20028,N_20029,N_20030,N_20031,N_20032,N_20033,N_20034,N_20035,N_20036,N_20037,N_20038,N_20039,N_20040,N_20041,N_20042,N_20043,N_20044,N_20045,N_20046,N_20047,N_20048,N_20049,N_20050,N_20051,N_20052,N_20053,N_20054,N_20055,N_20056,N_20057,N_20058,N_20059,N_20060,N_20061,N_20062,N_20063,N_20064,N_20065,N_20066,N_20067,N_20068,N_20069,N_20070,N_20071,N_20072,N_20073,N_20074,N_20075,N_20076,N_20077,N_20078,N_20079,N_20080,N_20081,N_20082,N_20083,N_20084,N_20085,N_20086,N_20087,N_20088,N_20089,N_20090,N_20091,N_20092,N_20093,N_20094,N_20095,N_20096,N_20097,N_20098,N_20099,N_20100,N_20101,N_20102,N_20103,N_20104,N_20105,N_20106,N_20107,N_20108,N_20109,N_20110,N_20111,N_20112,N_20113,N_20114,N_20115,N_20116,N_20117,N_20118,N_20119,N_20120,N_20121,N_20122,N_20123,N_20124,N_20125,N_20126,N_20127,N_20128,N_20129,N_20130,N_20131,N_20132,N_20133,N_20134,N_20135,N_20136,N_20137,N_20138,N_20139,N_20140,N_20141,N_20142,N_20143,N_20144,N_20145,N_20146,N_20147,N_20148,N_20149,N_20150,N_20151,N_20152,N_20153,N_20154,N_20155,N_20156,N_20157,N_20158,N_20159,N_20160,N_20161,N_20162,N_20163,N_20164,N_20165,N_20166,N_20167,N_20168,N_20169,N_20170,N_20171,N_20172,N_20173,N_20174,N_20175,N_20176,N_20177,N_20178,N_20179,N_20180,N_20181,N_20182,N_20183,N_20184,N_20185,N_20186,N_20187,N_20188,N_20189,N_20190,N_20191,N_20192,N_20193,N_20194,N_20195,N_20196,N_20197,N_20198,N_20199,N_20200,N_20201,N_20202,N_20203,N_20204,N_20205,N_20206,N_20207,N_20208,N_20209,N_20210,N_20211,N_20212,N_20213,N_20214,N_20215,N_20216,N_20217,N_20218,N_20219,N_20220,N_20221,N_20222,N_20223,N_20224,N_20225,N_20226,N_20227,N_20228,N_20229,N_20230,N_20231,N_20232,N_20233,N_20234,N_20235,N_20236,N_20237,N_20238,N_20239,N_20240,N_20241,N_20242,N_20243,N_20244,N_20245,N_20246,N_20247,N_20248,N_20249,N_20250,N_20251,N_20252,N_20253,N_20254,N_20255,N_20256,N_20257,N_20258,N_20259,N_20260,N_20261,N_20262,N_20263,N_20264,N_20265,N_20266,N_20267,N_20268,N_20269,N_20270,N_20271,N_20272,N_20273,N_20274,N_20275,N_20276,N_20277,N_20278,N_20279,N_20280,N_20281,N_20282,N_20283,N_20284,N_20285,N_20286,N_20287,N_20288,N_20289,N_20290,N_20291,N_20292,N_20293,N_20294,N_20295,N_20296,N_20297,N_20298,N_20299,N_20300,N_20301,N_20302,N_20303,N_20304,N_20305,N_20306,N_20307,N_20308,N_20309,N_20310,N_20311,N_20312,N_20313,N_20314,N_20315,N_20316,N_20317,N_20318,N_20319,N_20320,N_20321,N_20322,N_20323,N_20324,N_20325,N_20326,N_20327,N_20328,N_20329,N_20330,N_20331,N_20332,N_20333,N_20334,N_20335,N_20336,N_20337,N_20338,N_20339,N_20340,N_20341,N_20342,N_20343,N_20344,N_20345,N_20346,N_20347,N_20348,N_20349,N_20350,N_20351,N_20352,N_20353,N_20354,N_20355,N_20356,N_20357,N_20358,N_20359,N_20360,N_20361,N_20362,N_20363,N_20364,N_20365,N_20366,N_20367,N_20368,N_20369,N_20370,N_20371,N_20372,N_20373,N_20374,N_20375,N_20376,N_20377,N_20378,N_20379,N_20380,N_20381,N_20382,N_20383,N_20384,N_20385,N_20386,N_20387,N_20388,N_20389,N_20390,N_20391,N_20392,N_20393,N_20394,N_20395,N_20396,N_20397,N_20398,N_20399,N_20400,N_20401,N_20402,N_20403,N_20404,N_20405,N_20406,N_20407,N_20408,N_20409,N_20410,N_20411,N_20412,N_20413,N_20414,N_20415,N_20416,N_20417,N_20418,N_20419,N_20420,N_20421,N_20422,N_20423,N_20424,N_20425,N_20426,N_20427,N_20428,N_20429,N_20430,N_20431,N_20432,N_20433,N_20434,N_20435,N_20436,N_20437,N_20438,N_20439,N_20440,N_20441,N_20442,N_20443,N_20444,N_20445,N_20446,N_20447,N_20448,N_20449,N_20450,N_20451,N_20452,N_20453,N_20454,N_20455,N_20456,N_20457,N_20458,N_20459,N_20460,N_20461,N_20462,N_20463,N_20464,N_20465,N_20466,N_20467,N_20468,N_20469,N_20470,N_20471,N_20472,N_20473,N_20474,N_20475,N_20476,N_20477,N_20478,N_20479,N_20480,N_20481,N_20482,N_20483,N_20484,N_20485,N_20486,N_20487,N_20488,N_20489,N_20490,N_20491,N_20492,N_20493,N_20494,N_20495,N_20496,N_20497,N_20498,N_20499,N_20500,N_20501,N_20502,N_20503,N_20504,N_20505,N_20506,N_20507,N_20508,N_20509,N_20510,N_20511,N_20512,N_20513,N_20514,N_20515,N_20516,N_20517,N_20518,N_20519,N_20520,N_20521,N_20522,N_20523,N_20524,N_20525,N_20526,N_20527,N_20528,N_20529,N_20530,N_20531,N_20532,N_20533,N_20534,N_20535,N_20536,N_20537,N_20538,N_20539,N_20540,N_20541,N_20542,N_20543,N_20544,N_20545,N_20546,N_20547,N_20548,N_20549,N_20550,N_20551,N_20552,N_20553,N_20554,N_20555,N_20556,N_20557,N_20558,N_20559,N_20560,N_20561,N_20562,N_20563,N_20564,N_20565,N_20566,N_20567,N_20568,N_20569,N_20570,N_20571,N_20572,N_20573,N_20574,N_20575,N_20576,N_20577,N_20578,N_20579,N_20580,N_20581,N_20582,N_20583,N_20584,N_20585,N_20586,N_20587,N_20588,N_20589,N_20590,N_20591,N_20592,N_20593,N_20594,N_20595,N_20596,N_20597,N_20598,N_20599,N_20600,N_20601,N_20602,N_20603,N_20604,N_20605,N_20606,N_20607,N_20608,N_20609,N_20610,N_20611,N_20612,N_20613,N_20614,N_20615,N_20616,N_20617,N_20618,N_20619,N_20620,N_20621,N_20622,N_20623,N_20624,N_20625,N_20626,N_20627,N_20628,N_20629,N_20630,N_20631,N_20632,N_20633,N_20634,N_20635,N_20636,N_20637,N_20638,N_20639,N_20640,N_20641,N_20642,N_20643,N_20644,N_20645,N_20646,N_20647,N_20648,N_20649,N_20650,N_20651,N_20652,N_20653,N_20654,N_20655,N_20656,N_20657,N_20658,N_20659,N_20660,N_20661,N_20662,N_20663,N_20664,N_20665,N_20666,N_20667,N_20668,N_20669,N_20670,N_20671,N_20672,N_20673,N_20674,N_20675,N_20676,N_20677,N_20678,N_20679,N_20680,N_20681,N_20682,N_20683,N_20684,N_20685,N_20686,N_20687,N_20688,N_20689,N_20690,N_20691,N_20692,N_20693,N_20694,N_20695,N_20696,N_20697,N_20698,N_20699,N_20700,N_20701,N_20702,N_20703,N_20704,N_20705,N_20706,N_20707,N_20708,N_20709,N_20710,N_20711,N_20712,N_20713,N_20714,N_20715,N_20716,N_20717,N_20718,N_20719,N_20720,N_20721,N_20722,N_20723,N_20724,N_20725,N_20726,N_20727,N_20728,N_20729,N_20730,N_20731,N_20732,N_20733,N_20734,N_20735,N_20736,N_20737,N_20738,N_20739,N_20740,N_20741,N_20742,N_20743,N_20744,N_20745,N_20746,N_20747,N_20748,N_20749,N_20750,N_20751,N_20752,N_20753,N_20754,N_20755,N_20756,N_20757,N_20758,N_20759,N_20760,N_20761,N_20762,N_20763,N_20764,N_20765,N_20766,N_20767,N_20768,N_20769,N_20770,N_20771,N_20772,N_20773,N_20774,N_20775,N_20776,N_20777,N_20778,N_20779,N_20780,N_20781,N_20782,N_20783,N_20784,N_20785,N_20786,N_20787,N_20788,N_20789,N_20790,N_20791,N_20792,N_20793,N_20794,N_20795,N_20796,N_20797,N_20798,N_20799,N_20800,N_20801,N_20802,N_20803,N_20804,N_20805,N_20806,N_20807,N_20808,N_20809,N_20810,N_20811,N_20812,N_20813,N_20814,N_20815,N_20816,N_20817,N_20818,N_20819,N_20820,N_20821,N_20822,N_20823,N_20824,N_20825,N_20826,N_20827,N_20828,N_20829,N_20830,N_20831,N_20832,N_20833,N_20834,N_20835,N_20836,N_20837,N_20838,N_20839,N_20840,N_20841,N_20842,N_20843,N_20844,N_20845,N_20846,N_20847,N_20848,N_20849,N_20850,N_20851,N_20852,N_20853,N_20854,N_20855,N_20856,N_20857,N_20858,N_20859,N_20860,N_20861,N_20862,N_20863,N_20864,N_20865,N_20866,N_20867,N_20868,N_20869,N_20870,N_20871,N_20872,N_20873,N_20874,N_20875,N_20876,N_20877,N_20878,N_20879,N_20880,N_20881,N_20882,N_20883,N_20884,N_20885,N_20886,N_20887,N_20888,N_20889,N_20890,N_20891,N_20892,N_20893,N_20894,N_20895,N_20896,N_20897,N_20898,N_20899,N_20900,N_20901,N_20902,N_20903,N_20904,N_20905,N_20906,N_20907,N_20908,N_20909,N_20910,N_20911,N_20912,N_20913,N_20914,N_20915,N_20916,N_20917,N_20918,N_20919,N_20920,N_20921,N_20922,N_20923,N_20924,N_20925,N_20926,N_20927,N_20928,N_20929,N_20930,N_20931,N_20932,N_20933,N_20934,N_20935,N_20936,N_20937,N_20938,N_20939,N_20940,N_20941,N_20942,N_20943,N_20944,N_20945,N_20946,N_20947,N_20948,N_20949,N_20950,N_20951,N_20952,N_20953,N_20954,N_20955,N_20956,N_20957,N_20958,N_20959,N_20960,N_20961,N_20962,N_20963,N_20964,N_20965,N_20966,N_20967,N_20968,N_20969,N_20970,N_20971,N_20972,N_20973,N_20974,N_20975,N_20976,N_20977,N_20978,N_20979,N_20980,N_20981,N_20982,N_20983,N_20984,N_20985,N_20986,N_20987,N_20988,N_20989,N_20990,N_20991,N_20992,N_20993,N_20994,N_20995,N_20996,N_20997,N_20998,N_20999,N_21000,N_21001,N_21002,N_21003,N_21004,N_21005,N_21006,N_21007,N_21008,N_21009,N_21010,N_21011,N_21012,N_21013,N_21014,N_21015,N_21016,N_21017,N_21018,N_21019,N_21020,N_21021,N_21022,N_21023,N_21024,N_21025,N_21026,N_21027,N_21028,N_21029,N_21030,N_21031,N_21032,N_21033,N_21034,N_21035,N_21036,N_21037,N_21038,N_21039,N_21040,N_21041,N_21042,N_21043,N_21044,N_21045,N_21046,N_21047,N_21048,N_21049,N_21050,N_21051,N_21052,N_21053,N_21054,N_21055,N_21056,N_21057,N_21058,N_21059,N_21060,N_21061,N_21062,N_21063,N_21064,N_21065,N_21066,N_21067,N_21068,N_21069,N_21070,N_21071,N_21072,N_21073,N_21074,N_21075,N_21076,N_21077,N_21078,N_21079,N_21080,N_21081,N_21082,N_21083,N_21084,N_21085,N_21086,N_21087,N_21088,N_21089,N_21090,N_21091,N_21092,N_21093,N_21094,N_21095,N_21096,N_21097,N_21098,N_21099,N_21100,N_21101,N_21102,N_21103,N_21104,N_21105,N_21106,N_21107,N_21108,N_21109,N_21110,N_21111,N_21112,N_21113,N_21114,N_21115,N_21116,N_21117,N_21118,N_21119,N_21120,N_21121,N_21122,N_21123,N_21124,N_21125,N_21126,N_21127,N_21128,N_21129,N_21130,N_21131,N_21132,N_21133,N_21134,N_21135,N_21136,N_21137,N_21138,N_21139,N_21140,N_21141,N_21142,N_21143,N_21144,N_21145,N_21146,N_21147,N_21148,N_21149,N_21150,N_21151,N_21152,N_21153,N_21154,N_21155,N_21156,N_21157,N_21158,N_21159,N_21160,N_21161,N_21162,N_21163,N_21164,N_21165,N_21166,N_21167,N_21168,N_21169,N_21170,N_21171,N_21172,N_21173,N_21174,N_21175,N_21176,N_21177,N_21178,N_21179,N_21180,N_21181,N_21182,N_21183,N_21184,N_21185,N_21186,N_21187,N_21188,N_21189,N_21190,N_21191,N_21192,N_21193,N_21194,N_21195,N_21196,N_21197,N_21198,N_21199,N_21200,N_21201,N_21202,N_21203,N_21204,N_21205,N_21206,N_21207,N_21208,N_21209,N_21210,N_21211,N_21212,N_21213,N_21214,N_21215,N_21216,N_21217,N_21218,N_21219,N_21220,N_21221,N_21222,N_21223,N_21224,N_21225,N_21226,N_21227,N_21228,N_21229,N_21230,N_21231,N_21232,N_21233,N_21234,N_21235,N_21236,N_21237,N_21238,N_21239,N_21240,N_21241,N_21242,N_21243,N_21244,N_21245,N_21246,N_21247,N_21248,N_21249,N_21250,N_21251,N_21252,N_21253,N_21254,N_21255,N_21256,N_21257,N_21258,N_21259,N_21260,N_21261,N_21262,N_21263,N_21264,N_21265,N_21266,N_21267,N_21268,N_21269,N_21270,N_21271,N_21272,N_21273,N_21274,N_21275,N_21276,N_21277,N_21278,N_21279,N_21280,N_21281,N_21282,N_21283,N_21284,N_21285,N_21286,N_21287,N_21288,N_21289,N_21290,N_21291,N_21292,N_21293,N_21294,N_21295,N_21296,N_21297,N_21298,N_21299,N_21300,N_21301,N_21302,N_21303,N_21304,N_21305,N_21306,N_21307,N_21308,N_21309,N_21310,N_21311,N_21312,N_21313,N_21314,N_21315,N_21316,N_21317,N_21318,N_21319,N_21320,N_21321,N_21322,N_21323,N_21324,N_21325,N_21326,N_21327,N_21328,N_21329,N_21330,N_21331,N_21332,N_21333,N_21334,N_21335,N_21336,N_21337,N_21338,N_21339,N_21340,N_21341,N_21342,N_21343,N_21344,N_21345,N_21346,N_21347,N_21348,N_21349,N_21350,N_21351,N_21352,N_21353,N_21354,N_21355,N_21356,N_21357,N_21358,N_21359,N_21360,N_21361,N_21362,N_21363,N_21364,N_21365,N_21366,N_21367,N_21368,N_21369,N_21370,N_21371,N_21372,N_21373,N_21374,N_21375,N_21376,N_21377,N_21378,N_21379,N_21380,N_21381,N_21382,N_21383,N_21384,N_21385,N_21386,N_21387,N_21388,N_21389,N_21390,N_21391,N_21392,N_21393,N_21394,N_21395,N_21396,N_21397,N_21398,N_21399,N_21400,N_21401,N_21402,N_21403,N_21404,N_21405,N_21406,N_21407,N_21408,N_21409,N_21410,N_21411,N_21412,N_21413,N_21414,N_21415,N_21416,N_21417,N_21418,N_21419,N_21420,N_21421,N_21422,N_21423,N_21424,N_21425,N_21426,N_21427,N_21428,N_21429,N_21430,N_21431,N_21432,N_21433,N_21434,N_21435,N_21436,N_21437,N_21438,N_21439,N_21440,N_21441,N_21442,N_21443,N_21444,N_21445,N_21446,N_21447,N_21448,N_21449,N_21450,N_21451,N_21452,N_21453,N_21454,N_21455,N_21456,N_21457,N_21458,N_21459,N_21460,N_21461,N_21462,N_21463,N_21464,N_21465,N_21466,N_21467,N_21468,N_21469,N_21470,N_21471,N_21472,N_21473,N_21474,N_21475,N_21476,N_21477,N_21478,N_21479,N_21480,N_21481,N_21482,N_21483,N_21484,N_21485,N_21486,N_21487,N_21488,N_21489,N_21490,N_21491,N_21492,N_21493,N_21494,N_21495,N_21496,N_21497,N_21498,N_21499,N_21500,N_21501,N_21502,N_21503,N_21504,N_21505,N_21506,N_21507,N_21508,N_21509,N_21510,N_21511,N_21512,N_21513,N_21514,N_21515,N_21516,N_21517,N_21518,N_21519,N_21520,N_21521,N_21522,N_21523,N_21524,N_21525,N_21526,N_21527,N_21528,N_21529,N_21530,N_21531,N_21532,N_21533,N_21534,N_21535,N_21536,N_21537,N_21538,N_21539,N_21540,N_21541,N_21542,N_21543,N_21544,N_21545,N_21546,N_21547,N_21548,N_21549,N_21550,N_21551,N_21552,N_21553,N_21554,N_21555,N_21556,N_21557,N_21558,N_21559,N_21560,N_21561,N_21562,N_21563,N_21564,N_21565,N_21566,N_21567,N_21568,N_21569,N_21570,N_21571,N_21572,N_21573,N_21574,N_21575,N_21576,N_21577,N_21578,N_21579,N_21580,N_21581,N_21582,N_21583,N_21584,N_21585,N_21586,N_21587,N_21588,N_21589,N_21590,N_21591,N_21592,N_21593,N_21594,N_21595,N_21596,N_21597,N_21598,N_21599,N_21600,N_21601,N_21602,N_21603,N_21604,N_21605,N_21606,N_21607,N_21608,N_21609,N_21610,N_21611,N_21612,N_21613,N_21614,N_21615,N_21616,N_21617,N_21618,N_21619,N_21620,N_21621,N_21622,N_21623,N_21624,N_21625,N_21626,N_21627,N_21628,N_21629,N_21630,N_21631,N_21632,N_21633,N_21634,N_21635,N_21636,N_21637,N_21638,N_21639,N_21640,N_21641,N_21642,N_21643,N_21644,N_21645,N_21646,N_21647,N_21648,N_21649,N_21650,N_21651,N_21652,N_21653,N_21654,N_21655,N_21656,N_21657,N_21658,N_21659,N_21660,N_21661,N_21662,N_21663,N_21664,N_21665,N_21666,N_21667,N_21668,N_21669,N_21670,N_21671,N_21672,N_21673,N_21674,N_21675,N_21676,N_21677,N_21678,N_21679,N_21680,N_21681,N_21682,N_21683,N_21684,N_21685,N_21686,N_21687,N_21688,N_21689,N_21690,N_21691,N_21692,N_21693,N_21694,N_21695,N_21696,N_21697,N_21698,N_21699,N_21700,N_21701,N_21702,N_21703,N_21704,N_21705,N_21706,N_21707,N_21708,N_21709,N_21710,N_21711,N_21712,N_21713,N_21714,N_21715,N_21716,N_21717,N_21718,N_21719,N_21720,N_21721,N_21722,N_21723,N_21724,N_21725,N_21726,N_21727,N_21728,N_21729,N_21730,N_21731,N_21732,N_21733,N_21734,N_21735,N_21736,N_21737,N_21738,N_21739,N_21740,N_21741,N_21742,N_21743,N_21744,N_21745,N_21746,N_21747,N_21748,N_21749,N_21750,N_21751,N_21752,N_21753,N_21754,N_21755,N_21756,N_21757,N_21758,N_21759,N_21760,N_21761,N_21762,N_21763,N_21764,N_21765,N_21766,N_21767,N_21768,N_21769,N_21770,N_21771,N_21772,N_21773,N_21774,N_21775,N_21776,N_21777,N_21778,N_21779,N_21780,N_21781,N_21782,N_21783,N_21784,N_21785,N_21786,N_21787,N_21788,N_21789,N_21790,N_21791,N_21792,N_21793,N_21794,N_21795,N_21796,N_21797,N_21798,N_21799,N_21800,N_21801,N_21802,N_21803,N_21804,N_21805,N_21806,N_21807,N_21808,N_21809,N_21810,N_21811,N_21812,N_21813,N_21814,N_21815,N_21816,N_21817,N_21818,N_21819,N_21820,N_21821,N_21822,N_21823,N_21824,N_21825,N_21826,N_21827,N_21828,N_21829,N_21830,N_21831,N_21832,N_21833,N_21834,N_21835,N_21836,N_21837,N_21838,N_21839,N_21840,N_21841,N_21842,N_21843,N_21844,N_21845,N_21846,N_21847,N_21848,N_21849,N_21850,N_21851,N_21852,N_21853,N_21854,N_21855,N_21856,N_21857,N_21858,N_21859,N_21860,N_21861,N_21862,N_21863,N_21864,N_21865,N_21866,N_21867,N_21868,N_21869,N_21870,N_21871,N_21872,N_21873,N_21874,N_21875,N_21876,N_21877,N_21878,N_21879,N_21880,N_21881,N_21882,N_21883,N_21884,N_21885,N_21886,N_21887,N_21888,N_21889,N_21890,N_21891,N_21892,N_21893,N_21894,N_21895,N_21896,N_21897,N_21898,N_21899,N_21900,N_21901,N_21902,N_21903,N_21904,N_21905,N_21906,N_21907,N_21908,N_21909,N_21910,N_21911,N_21912,N_21913,N_21914,N_21915,N_21916,N_21917,N_21918,N_21919,N_21920,N_21921,N_21922,N_21923,N_21924,N_21925,N_21926,N_21927,N_21928,N_21929,N_21930,N_21931,N_21932,N_21933,N_21934,N_21935,N_21936,N_21937,N_21938,N_21939,N_21940,N_21941,N_21942,N_21943,N_21944,N_21945,N_21946,N_21947,N_21948,N_21949,N_21950,N_21951,N_21952,N_21953,N_21954,N_21955,N_21956,N_21957,N_21958,N_21959,N_21960,N_21961,N_21962,N_21963,N_21964,N_21965,N_21966,N_21967,N_21968,N_21969,N_21970,N_21971,N_21972,N_21973,N_21974,N_21975,N_21976,N_21977,N_21978,N_21979,N_21980,N_21981,N_21982,N_21983,N_21984,N_21985,N_21986,N_21987,N_21988,N_21989,N_21990,N_21991,N_21992,N_21993,N_21994,N_21995,N_21996,N_21997,N_21998,N_21999,N_22000,N_22001,N_22002,N_22003,N_22004,N_22005,N_22006,N_22007,N_22008,N_22009,N_22010,N_22011,N_22012,N_22013,N_22014,N_22015,N_22016,N_22017,N_22018,N_22019,N_22020,N_22021,N_22022,N_22023,N_22024,N_22025,N_22026,N_22027,N_22028,N_22029,N_22030,N_22031,N_22032,N_22033,N_22034,N_22035,N_22036,N_22037,N_22038,N_22039,N_22040,N_22041,N_22042,N_22043,N_22044,N_22045,N_22046,N_22047,N_22048,N_22049,N_22050,N_22051,N_22052,N_22053,N_22054,N_22055,N_22056,N_22057,N_22058,N_22059,N_22060,N_22061,N_22062,N_22063,N_22064,N_22065,N_22066,N_22067,N_22068,N_22069,N_22070,N_22071,N_22072,N_22073,N_22074,N_22075,N_22076,N_22077,N_22078,N_22079,N_22080,N_22081,N_22082,N_22083,N_22084,N_22085,N_22086,N_22087,N_22088,N_22089,N_22090,N_22091,N_22092,N_22093,N_22094,N_22095,N_22096,N_22097,N_22098,N_22099,N_22100,N_22101,N_22102,N_22103,N_22104,N_22105,N_22106,N_22107,N_22108,N_22109,N_22110,N_22111,N_22112,N_22113,N_22114,N_22115,N_22116,N_22117,N_22118,N_22119,N_22120,N_22121,N_22122,N_22123,N_22124,N_22125,N_22126,N_22127,N_22128,N_22129,N_22130,N_22131,N_22132,N_22133,N_22134,N_22135,N_22136,N_22137,N_22138,N_22139,N_22140,N_22141,N_22142,N_22143,N_22144,N_22145,N_22146,N_22147,N_22148,N_22149,N_22150,N_22151,N_22152,N_22153,N_22154,N_22155,N_22156,N_22157,N_22158,N_22159,N_22160,N_22161,N_22162,N_22163,N_22164,N_22165,N_22166,N_22167,N_22168,N_22169,N_22170,N_22171,N_22172,N_22173,N_22174,N_22175,N_22176,N_22177,N_22178,N_22179,N_22180,N_22181,N_22182,N_22183,N_22184,N_22185,N_22186,N_22187,N_22188,N_22189,N_22190,N_22191,N_22192,N_22193,N_22194,N_22195,N_22196,N_22197,N_22198,N_22199,N_22200,N_22201,N_22202,N_22203,N_22204,N_22205,N_22206,N_22207,N_22208,N_22209,N_22210,N_22211,N_22212,N_22213,N_22214,N_22215,N_22216,N_22217,N_22218,N_22219,N_22220,N_22221,N_22222,N_22223,N_22224,N_22225,N_22226,N_22227,N_22228,N_22229,N_22230,N_22231,N_22232,N_22233,N_22234,N_22235,N_22236,N_22237,N_22238,N_22239,N_22240,N_22241,N_22242,N_22243,N_22244,N_22245,N_22246,N_22247,N_22248,N_22249,N_22250,N_22251,N_22252,N_22253,N_22254,N_22255,N_22256,N_22257,N_22258,N_22259,N_22260,N_22261,N_22262,N_22263,N_22264,N_22265,N_22266,N_22267,N_22268,N_22269,N_22270,N_22271,N_22272,N_22273,N_22274,N_22275,N_22276,N_22277,N_22278,N_22279,N_22280,N_22281,N_22282,N_22283,N_22284,N_22285,N_22286,N_22287,N_22288,N_22289,N_22290,N_22291,N_22292,N_22293,N_22294,N_22295,N_22296,N_22297,N_22298,N_22299,N_22300,N_22301,N_22302,N_22303,N_22304,N_22305,N_22306,N_22307,N_22308,N_22309,N_22310,N_22311,N_22312,N_22313,N_22314,N_22315,N_22316,N_22317,N_22318,N_22319,N_22320,N_22321,N_22322,N_22323,N_22324,N_22325,N_22326,N_22327,N_22328,N_22329,N_22330,N_22331,N_22332,N_22333,N_22334,N_22335,N_22336,N_22337,N_22338,N_22339,N_22340,N_22341,N_22342,N_22343,N_22344,N_22345,N_22346,N_22347,N_22348,N_22349,N_22350,N_22351,N_22352,N_22353,N_22354,N_22355,N_22356,N_22357,N_22358,N_22359,N_22360,N_22361,N_22362,N_22363,N_22364,N_22365,N_22366,N_22367,N_22368,N_22369,N_22370,N_22371,N_22372,N_22373,N_22374,N_22375,N_22376,N_22377,N_22378,N_22379,N_22380,N_22381,N_22382,N_22383,N_22384,N_22385,N_22386,N_22387,N_22388,N_22389,N_22390,N_22391,N_22392,N_22393,N_22394,N_22395,N_22396,N_22397,N_22398,N_22399,N_22400,N_22401,N_22402,N_22403,N_22404,N_22405,N_22406,N_22407,N_22408,N_22409,N_22410,N_22411,N_22412,N_22413,N_22414,N_22415,N_22416,N_22417,N_22418,N_22419,N_22420,N_22421,N_22422,N_22423,N_22424,N_22425,N_22426,N_22427,N_22428,N_22429,N_22430,N_22431,N_22432,N_22433,N_22434,N_22435,N_22436,N_22437,N_22438,N_22439,N_22440,N_22441,N_22442,N_22443,N_22444,N_22445,N_22446,N_22447,N_22448,N_22449,N_22450,N_22451,N_22452,N_22453,N_22454,N_22455,N_22456,N_22457,N_22458,N_22459,N_22460,N_22461,N_22462,N_22463,N_22464,N_22465,N_22466,N_22467,N_22468,N_22469,N_22470,N_22471,N_22472,N_22473,N_22474,N_22475,N_22476,N_22477,N_22478,N_22479,N_22480,N_22481,N_22482,N_22483,N_22484,N_22485,N_22486,N_22487,N_22488,N_22489,N_22490,N_22491,N_22492,N_22493,N_22494,N_22495,N_22496,N_22497,N_22498,N_22499,N_22500,N_22501,N_22502,N_22503,N_22504,N_22505,N_22506,N_22507,N_22508,N_22509,N_22510,N_22511,N_22512,N_22513,N_22514,N_22515,N_22516,N_22517,N_22518,N_22519,N_22520,N_22521,N_22522,N_22523,N_22524,N_22525,N_22526,N_22527,N_22528,N_22529,N_22530,N_22531,N_22532,N_22533,N_22534,N_22535,N_22536,N_22537,N_22538,N_22539,N_22540,N_22541,N_22542,N_22543,N_22544,N_22545,N_22546,N_22547,N_22548,N_22549,N_22550,N_22551,N_22552,N_22553,N_22554,N_22555,N_22556,N_22557,N_22558,N_22559,N_22560,N_22561,N_22562,N_22563,N_22564,N_22565,N_22566,N_22567,N_22568,N_22569,N_22570,N_22571,N_22572,N_22573,N_22574,N_22575,N_22576,N_22577,N_22578,N_22579,N_22580,N_22581,N_22582,N_22583,N_22584,N_22585,N_22586,N_22587,N_22588,N_22589,N_22590,N_22591,N_22592,N_22593,N_22594,N_22595,N_22596,N_22597,N_22598,N_22599,N_22600,N_22601,N_22602,N_22603,N_22604,N_22605,N_22606,N_22607,N_22608,N_22609,N_22610,N_22611,N_22612,N_22613,N_22614,N_22615,N_22616,N_22617,N_22618,N_22619,N_22620,N_22621,N_22622,N_22623,N_22624,N_22625,N_22626,N_22627,N_22628,N_22629,N_22630,N_22631,N_22632,N_22633,N_22634,N_22635,N_22636,N_22637,N_22638,N_22639,N_22640,N_22641,N_22642,N_22643,N_22644,N_22645,N_22646,N_22647,N_22648,N_22649,N_22650,N_22651,N_22652,N_22653,N_22654,N_22655,N_22656,N_22657,N_22658,N_22659,N_22660,N_22661,N_22662,N_22663,N_22664,N_22665,N_22666,N_22667,N_22668,N_22669,N_22670,N_22671,N_22672,N_22673,N_22674,N_22675,N_22676,N_22677,N_22678,N_22679,N_22680,N_22681,N_22682,N_22683,N_22684,N_22685,N_22686,N_22687,N_22688,N_22689,N_22690,N_22691,N_22692,N_22693,N_22694,N_22695,N_22696,N_22697,N_22698,N_22699,N_22700,N_22701,N_22702,N_22703,N_22704,N_22705,N_22706,N_22707,N_22708,N_22709,N_22710,N_22711,N_22712,N_22713,N_22714,N_22715,N_22716,N_22717,N_22718,N_22719,N_22720,N_22721,N_22722,N_22723,N_22724,N_22725,N_22726,N_22727,N_22728,N_22729,N_22730,N_22731,N_22732,N_22733,N_22734,N_22735,N_22736,N_22737,N_22738,N_22739,N_22740,N_22741,N_22742,N_22743,N_22744,N_22745,N_22746,N_22747,N_22748,N_22749,N_22750,N_22751,N_22752,N_22753,N_22754,N_22755,N_22756,N_22757,N_22758,N_22759,N_22760,N_22761,N_22762,N_22763,N_22764,N_22765,N_22766,N_22767,N_22768,N_22769,N_22770,N_22771,N_22772,N_22773,N_22774,N_22775,N_22776,N_22777,N_22778,N_22779,N_22780,N_22781,N_22782,N_22783,N_22784,N_22785,N_22786,N_22787,N_22788,N_22789,N_22790,N_22791,N_22792,N_22793,N_22794,N_22795,N_22796,N_22797,N_22798,N_22799,N_22800,N_22801,N_22802,N_22803,N_22804,N_22805,N_22806,N_22807,N_22808,N_22809,N_22810,N_22811,N_22812,N_22813,N_22814,N_22815,N_22816,N_22817,N_22818,N_22819,N_22820,N_22821,N_22822,N_22823,N_22824,N_22825,N_22826,N_22827,N_22828,N_22829,N_22830,N_22831,N_22832,N_22833,N_22834,N_22835,N_22836,N_22837,N_22838,N_22839,N_22840,N_22841,N_22842,N_22843,N_22844,N_22845,N_22846,N_22847,N_22848,N_22849,N_22850,N_22851,N_22852,N_22853,N_22854,N_22855,N_22856,N_22857,N_22858,N_22859,N_22860,N_22861,N_22862,N_22863,N_22864,N_22865,N_22866,N_22867,N_22868,N_22869,N_22870,N_22871,N_22872,N_22873,N_22874,N_22875,N_22876,N_22877,N_22878,N_22879,N_22880,N_22881,N_22882,N_22883,N_22884,N_22885,N_22886,N_22887,N_22888,N_22889,N_22890,N_22891,N_22892,N_22893,N_22894,N_22895,N_22896,N_22897,N_22898,N_22899,N_22900,N_22901,N_22902,N_22903,N_22904,N_22905,N_22906,N_22907,N_22908,N_22909,N_22910,N_22911,N_22912,N_22913,N_22914,N_22915,N_22916,N_22917,N_22918,N_22919,N_22920,N_22921,N_22922,N_22923,N_22924,N_22925,N_22926,N_22927,N_22928,N_22929,N_22930,N_22931,N_22932,N_22933,N_22934,N_22935,N_22936,N_22937,N_22938,N_22939,N_22940,N_22941,N_22942,N_22943,N_22944,N_22945,N_22946,N_22947,N_22948,N_22949,N_22950,N_22951,N_22952,N_22953,N_22954,N_22955,N_22956,N_22957,N_22958,N_22959,N_22960,N_22961,N_22962,N_22963,N_22964,N_22965,N_22966,N_22967,N_22968,N_22969,N_22970,N_22971,N_22972,N_22973,N_22974,N_22975,N_22976,N_22977,N_22978,N_22979,N_22980,N_22981,N_22982,N_22983,N_22984,N_22985,N_22986,N_22987,N_22988,N_22989,N_22990,N_22991,N_22992,N_22993,N_22994,N_22995,N_22996,N_22997,N_22998,N_22999,N_23000,N_23001,N_23002,N_23003,N_23004,N_23005,N_23006,N_23007,N_23008,N_23009,N_23010,N_23011,N_23012,N_23013,N_23014,N_23015,N_23016,N_23017,N_23018,N_23019,N_23020,N_23021,N_23022,N_23023,N_23024,N_23025,N_23026,N_23027,N_23028,N_23029,N_23030,N_23031,N_23032,N_23033,N_23034,N_23035,N_23036,N_23037,N_23038,N_23039,N_23040,N_23041,N_23042,N_23043,N_23044,N_23045,N_23046,N_23047,N_23048,N_23049,N_23050,N_23051,N_23052,N_23053,N_23054,N_23055,N_23056,N_23057,N_23058,N_23059,N_23060,N_23061,N_23062,N_23063,N_23064,N_23065,N_23066,N_23067,N_23068,N_23069,N_23070,N_23071,N_23072,N_23073,N_23074,N_23075,N_23076,N_23077,N_23078,N_23079,N_23080,N_23081,N_23082,N_23083,N_23084,N_23085,N_23086,N_23087,N_23088,N_23089,N_23090,N_23091,N_23092,N_23093,N_23094,N_23095,N_23096,N_23097,N_23098,N_23099,N_23100,N_23101,N_23102,N_23103,N_23104,N_23105,N_23106,N_23107,N_23108,N_23109,N_23110,N_23111,N_23112,N_23113,N_23114,N_23115,N_23116,N_23117,N_23118,N_23119,N_23120,N_23121,N_23122,N_23123,N_23124,N_23125,N_23126,N_23127,N_23128,N_23129,N_23130,N_23131,N_23132,N_23133,N_23134,N_23135,N_23136,N_23137,N_23138,N_23139,N_23140,N_23141,N_23142,N_23143,N_23144,N_23145,N_23146,N_23147,N_23148,N_23149,N_23150,N_23151,N_23152,N_23153,N_23154,N_23155,N_23156,N_23157,N_23158,N_23159,N_23160,N_23161,N_23162,N_23163,N_23164,N_23165,N_23166,N_23167,N_23168,N_23169,N_23170,N_23171,N_23172,N_23173,N_23174,N_23175,N_23176,N_23177,N_23178,N_23179,N_23180,N_23181,N_23182,N_23183,N_23184,N_23185,N_23186,N_23187,N_23188,N_23189,N_23190,N_23191,N_23192,N_23193,N_23194,N_23195,N_23196,N_23197,N_23198,N_23199,N_23200,N_23201,N_23202,N_23203,N_23204,N_23205,N_23206,N_23207,N_23208,N_23209,N_23210,N_23211,N_23212,N_23213,N_23214,N_23215,N_23216,N_23217,N_23218,N_23219,N_23220,N_23221,N_23222,N_23223,N_23224,N_23225,N_23226,N_23227,N_23228,N_23229,N_23230,N_23231,N_23232,N_23233,N_23234,N_23235,N_23236,N_23237,N_23238,N_23239,N_23240,N_23241,N_23242,N_23243,N_23244,N_23245,N_23246,N_23247,N_23248,N_23249,N_23250,N_23251,N_23252,N_23253,N_23254,N_23255,N_23256,N_23257,N_23258,N_23259,N_23260,N_23261,N_23262,N_23263,N_23264,N_23265,N_23266,N_23267,N_23268,N_23269,N_23270,N_23271,N_23272,N_23273,N_23274,N_23275,N_23276,N_23277,N_23278,N_23279,N_23280,N_23281,N_23282,N_23283,N_23284,N_23285,N_23286,N_23287,N_23288,N_23289,N_23290,N_23291,N_23292,N_23293,N_23294,N_23295,N_23296,N_23297,N_23298,N_23299,N_23300,N_23301,N_23302,N_23303,N_23304,N_23305,N_23306,N_23307,N_23308,N_23309,N_23310,N_23311,N_23312,N_23313,N_23314,N_23315,N_23316,N_23317,N_23318,N_23319,N_23320,N_23321,N_23322,N_23323,N_23324,N_23325,N_23326,N_23327,N_23328,N_23329,N_23330,N_23331,N_23332,N_23333,N_23334,N_23335,N_23336,N_23337,N_23338,N_23339,N_23340,N_23341,N_23342,N_23343,N_23344,N_23345,N_23346,N_23347,N_23348,N_23349,N_23350,N_23351,N_23352,N_23353,N_23354,N_23355,N_23356,N_23357,N_23358,N_23359,N_23360,N_23361,N_23362,N_23363,N_23364,N_23365,N_23366,N_23367,N_23368,N_23369,N_23370,N_23371,N_23372,N_23373,N_23374,N_23375,N_23376,N_23377,N_23378,N_23379,N_23380,N_23381,N_23382,N_23383,N_23384,N_23385,N_23386,N_23387,N_23388,N_23389,N_23390,N_23391,N_23392,N_23393,N_23394,N_23395,N_23396,N_23397,N_23398,N_23399,N_23400,N_23401,N_23402,N_23403,N_23404,N_23405,N_23406,N_23407,N_23408,N_23409,N_23410,N_23411,N_23412,N_23413,N_23414,N_23415,N_23416,N_23417,N_23418,N_23419,N_23420,N_23421,N_23422,N_23423,N_23424,N_23425,N_23426,N_23427,N_23428,N_23429,N_23430,N_23431,N_23432,N_23433,N_23434,N_23435,N_23436,N_23437,N_23438,N_23439,N_23440,N_23441,N_23442,N_23443,N_23444,N_23445,N_23446,N_23447,N_23448,N_23449,N_23450,N_23451,N_23452,N_23453,N_23454,N_23455,N_23456,N_23457,N_23458,N_23459,N_23460,N_23461,N_23462,N_23463,N_23464,N_23465,N_23466,N_23467,N_23468,N_23469,N_23470,N_23471,N_23472,N_23473,N_23474,N_23475,N_23476,N_23477,N_23478,N_23479,N_23480,N_23481,N_23482,N_23483,N_23484,N_23485,N_23486,N_23487,N_23488,N_23489,N_23490,N_23491,N_23492,N_23493,N_23494,N_23495,N_23496,N_23497,N_23498,N_23499,N_23500,N_23501,N_23502,N_23503,N_23504,N_23505,N_23506,N_23507,N_23508,N_23509,N_23510,N_23511,N_23512,N_23513,N_23514,N_23515,N_23516,N_23517,N_23518,N_23519,N_23520,N_23521,N_23522,N_23523,N_23524,N_23525,N_23526,N_23527,N_23528,N_23529,N_23530,N_23531,N_23532,N_23533,N_23534,N_23535,N_23536,N_23537,N_23538,N_23539,N_23540,N_23541,N_23542,N_23543,N_23544,N_23545,N_23546,N_23547,N_23548,N_23549,N_23550,N_23551,N_23552,N_23553,N_23554,N_23555,N_23556,N_23557,N_23558,N_23559,N_23560,N_23561,N_23562,N_23563,N_23564,N_23565,N_23566,N_23567,N_23568,N_23569,N_23570,N_23571,N_23572,N_23573,N_23574,N_23575,N_23576,N_23577,N_23578,N_23579,N_23580,N_23581,N_23582,N_23583,N_23584,N_23585,N_23586,N_23587,N_23588,N_23589,N_23590,N_23591,N_23592,N_23593,N_23594,N_23595,N_23596,N_23597,N_23598,N_23599,N_23600,N_23601,N_23602,N_23603,N_23604,N_23605,N_23606,N_23607,N_23608,N_23609,N_23610,N_23611,N_23612,N_23613,N_23614,N_23615,N_23616,N_23617,N_23618,N_23619,N_23620,N_23621,N_23622,N_23623,N_23624,N_23625,N_23626,N_23627,N_23628,N_23629,N_23630,N_23631,N_23632,N_23633,N_23634,N_23635,N_23636,N_23637,N_23638,N_23639,N_23640,N_23641,N_23642,N_23643,N_23644,N_23645,N_23646,N_23647,N_23648,N_23649,N_23650,N_23651,N_23652,N_23653,N_23654,N_23655,N_23656,N_23657,N_23658,N_23659,N_23660,N_23661,N_23662,N_23663,N_23664,N_23665,N_23666,N_23667,N_23668,N_23669,N_23670,N_23671,N_23672,N_23673,N_23674,N_23675,N_23676,N_23677,N_23678,N_23679,N_23680,N_23681,N_23682,N_23683,N_23684,N_23685,N_23686,N_23687,N_23688,N_23689,N_23690,N_23691,N_23692,N_23693,N_23694,N_23695,N_23696,N_23697,N_23698,N_23699,N_23700,N_23701,N_23702,N_23703,N_23704,N_23705,N_23706,N_23707,N_23708,N_23709,N_23710,N_23711,N_23712,N_23713,N_23714,N_23715,N_23716,N_23717,N_23718,N_23719,N_23720,N_23721,N_23722,N_23723,N_23724,N_23725,N_23726,N_23727,N_23728,N_23729,N_23730,N_23731,N_23732,N_23733,N_23734,N_23735,N_23736,N_23737,N_23738,N_23739,N_23740,N_23741,N_23742,N_23743,N_23744,N_23745,N_23746,N_23747,N_23748,N_23749,N_23750,N_23751,N_23752,N_23753,N_23754,N_23755,N_23756,N_23757,N_23758,N_23759,N_23760,N_23761,N_23762,N_23763,N_23764,N_23765,N_23766,N_23767,N_23768,N_23769,N_23770,N_23771,N_23772,N_23773,N_23774,N_23775,N_23776,N_23777,N_23778,N_23779,N_23780,N_23781,N_23782,N_23783,N_23784,N_23785,N_23786,N_23787,N_23788,N_23789,N_23790,N_23791,N_23792,N_23793,N_23794,N_23795,N_23796,N_23797,N_23798,N_23799,N_23800,N_23801,N_23802,N_23803,N_23804,N_23805,N_23806,N_23807,N_23808,N_23809,N_23810,N_23811,N_23812,N_23813,N_23814,N_23815,N_23816,N_23817,N_23818,N_23819,N_23820,N_23821,N_23822,N_23823,N_23824,N_23825,N_23826,N_23827,N_23828,N_23829,N_23830,N_23831,N_23832,N_23833,N_23834,N_23835,N_23836,N_23837,N_23838,N_23839,N_23840,N_23841,N_23842,N_23843,N_23844,N_23845,N_23846,N_23847,N_23848,N_23849,N_23850,N_23851,N_23852,N_23853,N_23854,N_23855,N_23856,N_23857,N_23858,N_23859,N_23860,N_23861,N_23862,N_23863,N_23864,N_23865,N_23866,N_23867,N_23868,N_23869,N_23870,N_23871,N_23872,N_23873,N_23874,N_23875,N_23876,N_23877,N_23878,N_23879,N_23880,N_23881,N_23882,N_23883,N_23884,N_23885,N_23886,N_23887,N_23888,N_23889,N_23890,N_23891,N_23892,N_23893,N_23894,N_23895,N_23896,N_23897,N_23898,N_23899,N_23900,N_23901,N_23902,N_23903,N_23904,N_23905,N_23906,N_23907,N_23908,N_23909,N_23910,N_23911,N_23912,N_23913,N_23914,N_23915,N_23916,N_23917,N_23918,N_23919,N_23920,N_23921,N_23922,N_23923,N_23924,N_23925,N_23926,N_23927,N_23928,N_23929,N_23930,N_23931,N_23932,N_23933,N_23934,N_23935,N_23936,N_23937,N_23938,N_23939,N_23940,N_23941,N_23942,N_23943,N_23944,N_23945,N_23946,N_23947,N_23948,N_23949,N_23950,N_23951,N_23952,N_23953,N_23954,N_23955,N_23956,N_23957,N_23958,N_23959,N_23960,N_23961,N_23962,N_23963,N_23964,N_23965,N_23966,N_23967,N_23968,N_23969,N_23970,N_23971,N_23972,N_23973,N_23974,N_23975,N_23976,N_23977,N_23978,N_23979,N_23980,N_23981,N_23982,N_23983,N_23984,N_23985,N_23986,N_23987,N_23988,N_23989,N_23990,N_23991,N_23992,N_23993,N_23994,N_23995,N_23996,N_23997,N_23998,N_23999,N_24000,N_24001,N_24002,N_24003,N_24004,N_24005,N_24006,N_24007,N_24008,N_24009,N_24010,N_24011,N_24012,N_24013,N_24014,N_24015,N_24016,N_24017,N_24018,N_24019,N_24020,N_24021,N_24022,N_24023,N_24024,N_24025,N_24026,N_24027,N_24028,N_24029,N_24030,N_24031,N_24032,N_24033,N_24034,N_24035,N_24036,N_24037,N_24038,N_24039,N_24040,N_24041,N_24042,N_24043,N_24044,N_24045,N_24046,N_24047,N_24048,N_24049,N_24050,N_24051,N_24052,N_24053,N_24054,N_24055,N_24056,N_24057,N_24058,N_24059,N_24060,N_24061,N_24062,N_24063,N_24064,N_24065,N_24066,N_24067,N_24068,N_24069,N_24070,N_24071,N_24072,N_24073,N_24074,N_24075,N_24076,N_24077,N_24078,N_24079,N_24080,N_24081,N_24082,N_24083,N_24084,N_24085,N_24086,N_24087,N_24088,N_24089,N_24090,N_24091,N_24092,N_24093,N_24094,N_24095,N_24096,N_24097,N_24098,N_24099,N_24100,N_24101,N_24102,N_24103,N_24104,N_24105,N_24106,N_24107,N_24108,N_24109,N_24110,N_24111,N_24112,N_24113,N_24114,N_24115,N_24116,N_24117,N_24118,N_24119,N_24120,N_24121,N_24122,N_24123,N_24124,N_24125,N_24126,N_24127,N_24128,N_24129,N_24130,N_24131,N_24132,N_24133,N_24134,N_24135,N_24136,N_24137,N_24138,N_24139,N_24140,N_24141,N_24142,N_24143,N_24144,N_24145,N_24146,N_24147,N_24148,N_24149,N_24150,N_24151,N_24152,N_24153,N_24154,N_24155,N_24156,N_24157,N_24158,N_24159,N_24160,N_24161,N_24162,N_24163,N_24164,N_24165,N_24166,N_24167,N_24168,N_24169,N_24170,N_24171,N_24172,N_24173,N_24174,N_24175,N_24176,N_24177,N_24178,N_24179,N_24180,N_24181,N_24182,N_24183,N_24184,N_24185,N_24186,N_24187,N_24188,N_24189,N_24190,N_24191,N_24192,N_24193,N_24194,N_24195,N_24196,N_24197,N_24198,N_24199,N_24200,N_24201,N_24202,N_24203,N_24204,N_24205,N_24206,N_24207,N_24208,N_24209,N_24210,N_24211,N_24212,N_24213,N_24214,N_24215,N_24216,N_24217,N_24218,N_24219,N_24220,N_24221,N_24222,N_24223,N_24224,N_24225,N_24226,N_24227,N_24228,N_24229,N_24230,N_24231,N_24232,N_24233,N_24234,N_24235,N_24236,N_24237,N_24238,N_24239,N_24240,N_24241,N_24242,N_24243,N_24244,N_24245,N_24246,N_24247,N_24248,N_24249,N_24250,N_24251,N_24252,N_24253,N_24254,N_24255,N_24256,N_24257,N_24258,N_24259,N_24260,N_24261,N_24262,N_24263,N_24264,N_24265,N_24266,N_24267,N_24268,N_24269,N_24270,N_24271,N_24272,N_24273,N_24274,N_24275,N_24276,N_24277,N_24278,N_24279,N_24280,N_24281,N_24282,N_24283,N_24284,N_24285,N_24286,N_24287,N_24288,N_24289,N_24290,N_24291,N_24292,N_24293,N_24294,N_24295,N_24296,N_24297,N_24298,N_24299,N_24300,N_24301,N_24302,N_24303,N_24304,N_24305,N_24306,N_24307,N_24308,N_24309,N_24310,N_24311,N_24312,N_24313,N_24314,N_24315,N_24316,N_24317,N_24318,N_24319,N_24320,N_24321,N_24322,N_24323,N_24324,N_24325,N_24326,N_24327,N_24328,N_24329,N_24330,N_24331,N_24332,N_24333,N_24334,N_24335,N_24336,N_24337,N_24338,N_24339,N_24340,N_24341,N_24342,N_24343,N_24344,N_24345,N_24346,N_24347,N_24348,N_24349,N_24350,N_24351,N_24352,N_24353,N_24354,N_24355,N_24356,N_24357,N_24358,N_24359,N_24360,N_24361,N_24362,N_24363,N_24364,N_24365,N_24366,N_24367,N_24368,N_24369,N_24370,N_24371,N_24372,N_24373,N_24374,N_24375,N_24376,N_24377,N_24378,N_24379,N_24380,N_24381,N_24382,N_24383,N_24384,N_24385,N_24386,N_24387,N_24388,N_24389,N_24390,N_24391,N_24392,N_24393,N_24394,N_24395,N_24396,N_24397,N_24398,N_24399,N_24400,N_24401,N_24402,N_24403,N_24404,N_24405,N_24406,N_24407,N_24408,N_24409,N_24410,N_24411,N_24412,N_24413,N_24414,N_24415,N_24416,N_24417,N_24418,N_24419,N_24420,N_24421,N_24422,N_24423,N_24424,N_24425,N_24426,N_24427,N_24428,N_24429,N_24430,N_24431,N_24432,N_24433,N_24434,N_24435,N_24436,N_24437,N_24438,N_24439,N_24440,N_24441,N_24442,N_24443,N_24444,N_24445,N_24446,N_24447,N_24448,N_24449,N_24450,N_24451,N_24452,N_24453,N_24454,N_24455,N_24456,N_24457,N_24458,N_24459,N_24460,N_24461,N_24462,N_24463,N_24464,N_24465,N_24466,N_24467,N_24468,N_24469,N_24470,N_24471,N_24472,N_24473,N_24474,N_24475,N_24476,N_24477,N_24478,N_24479,N_24480,N_24481,N_24482,N_24483,N_24484,N_24485,N_24486,N_24487,N_24488,N_24489,N_24490,N_24491,N_24492,N_24493,N_24494,N_24495,N_24496,N_24497,N_24498,N_24499,N_24500,N_24501,N_24502,N_24503,N_24504,N_24505,N_24506,N_24507,N_24508,N_24509,N_24510,N_24511,N_24512,N_24513,N_24514,N_24515,N_24516,N_24517,N_24518,N_24519,N_24520,N_24521,N_24522,N_24523,N_24524,N_24525,N_24526,N_24527,N_24528,N_24529,N_24530,N_24531,N_24532,N_24533,N_24534,N_24535,N_24536,N_24537,N_24538,N_24539,N_24540,N_24541,N_24542,N_24543,N_24544,N_24545,N_24546,N_24547,N_24548,N_24549,N_24550,N_24551,N_24552,N_24553,N_24554,N_24555,N_24556,N_24557,N_24558,N_24559,N_24560,N_24561,N_24562,N_24563,N_24564,N_24565,N_24566,N_24567,N_24568,N_24569,N_24570,N_24571,N_24572,N_24573,N_24574,N_24575,N_24576,N_24577,N_24578,N_24579,N_24580,N_24581,N_24582,N_24583,N_24584,N_24585,N_24586,N_24587,N_24588,N_24589,N_24590,N_24591,N_24592,N_24593,N_24594,N_24595,N_24596,N_24597,N_24598,N_24599,N_24600,N_24601,N_24602,N_24603,N_24604,N_24605,N_24606,N_24607,N_24608,N_24609,N_24610,N_24611,N_24612,N_24613,N_24614,N_24615,N_24616,N_24617,N_24618,N_24619,N_24620,N_24621,N_24622,N_24623,N_24624,N_24625,N_24626,N_24627,N_24628,N_24629,N_24630,N_24631,N_24632,N_24633,N_24634,N_24635,N_24636,N_24637,N_24638,N_24639,N_24640,N_24641,N_24642,N_24643,N_24644,N_24645,N_24646,N_24647,N_24648,N_24649,N_24650,N_24651,N_24652,N_24653,N_24654,N_24655,N_24656,N_24657,N_24658,N_24659,N_24660,N_24661,N_24662,N_24663,N_24664,N_24665,N_24666,N_24667,N_24668,N_24669,N_24670,N_24671,N_24672,N_24673,N_24674,N_24675,N_24676,N_24677,N_24678,N_24679,N_24680,N_24681,N_24682,N_24683,N_24684,N_24685,N_24686,N_24687,N_24688,N_24689,N_24690,N_24691,N_24692,N_24693,N_24694,N_24695,N_24696,N_24697,N_24698,N_24699,N_24700,N_24701,N_24702,N_24703,N_24704,N_24705,N_24706,N_24707,N_24708,N_24709,N_24710,N_24711,N_24712,N_24713,N_24714,N_24715,N_24716,N_24717,N_24718,N_24719,N_24720,N_24721,N_24722,N_24723,N_24724,N_24725,N_24726,N_24727,N_24728,N_24729,N_24730,N_24731,N_24732,N_24733,N_24734,N_24735,N_24736,N_24737,N_24738,N_24739,N_24740,N_24741,N_24742,N_24743,N_24744,N_24745,N_24746,N_24747,N_24748,N_24749,N_24750,N_24751,N_24752,N_24753,N_24754,N_24755,N_24756,N_24757,N_24758,N_24759,N_24760,N_24761,N_24762,N_24763,N_24764,N_24765,N_24766,N_24767,N_24768,N_24769,N_24770,N_24771,N_24772,N_24773,N_24774,N_24775,N_24776,N_24777,N_24778,N_24779,N_24780,N_24781,N_24782,N_24783,N_24784,N_24785,N_24786,N_24787,N_24788,N_24789,N_24790,N_24791,N_24792,N_24793,N_24794,N_24795,N_24796,N_24797,N_24798,N_24799,N_24800,N_24801,N_24802,N_24803,N_24804,N_24805,N_24806,N_24807,N_24808,N_24809,N_24810,N_24811,N_24812,N_24813,N_24814,N_24815,N_24816,N_24817,N_24818,N_24819,N_24820,N_24821,N_24822,N_24823,N_24824,N_24825,N_24826,N_24827,N_24828,N_24829,N_24830,N_24831,N_24832,N_24833,N_24834,N_24835,N_24836,N_24837,N_24838,N_24839,N_24840,N_24841,N_24842,N_24843,N_24844,N_24845,N_24846,N_24847,N_24848,N_24849,N_24850,N_24851,N_24852,N_24853,N_24854,N_24855,N_24856,N_24857,N_24858,N_24859,N_24860,N_24861,N_24862,N_24863,N_24864,N_24865,N_24866,N_24867,N_24868,N_24869,N_24870,N_24871,N_24872,N_24873,N_24874,N_24875,N_24876,N_24877,N_24878,N_24879,N_24880,N_24881,N_24882,N_24883,N_24884,N_24885,N_24886,N_24887,N_24888,N_24889,N_24890,N_24891,N_24892,N_24893,N_24894,N_24895,N_24896,N_24897,N_24898,N_24899,N_24900,N_24901,N_24902,N_24903,N_24904,N_24905,N_24906,N_24907,N_24908,N_24909,N_24910,N_24911,N_24912,N_24913,N_24914,N_24915,N_24916,N_24917,N_24918,N_24919,N_24920,N_24921,N_24922,N_24923,N_24924,N_24925,N_24926,N_24927,N_24928,N_24929,N_24930,N_24931,N_24932,N_24933,N_24934,N_24935,N_24936,N_24937,N_24938,N_24939,N_24940,N_24941,N_24942,N_24943,N_24944,N_24945,N_24946,N_24947,N_24948,N_24949,N_24950,N_24951,N_24952,N_24953,N_24954,N_24955,N_24956,N_24957,N_24958,N_24959,N_24960,N_24961,N_24962,N_24963,N_24964,N_24965,N_24966,N_24967,N_24968,N_24969,N_24970,N_24971,N_24972,N_24973,N_24974,N_24975,N_24976,N_24977,N_24978,N_24979,N_24980,N_24981,N_24982,N_24983,N_24984,N_24985,N_24986,N_24987,N_24988,N_24989,N_24990,N_24991,N_24992,N_24993,N_24994,N_24995,N_24996,N_24997,N_24998,N_24999;
nor U0 (N_0,In_1777,In_1593);
nand U1 (N_1,In_1720,In_94);
nor U2 (N_2,In_1027,In_1922);
and U3 (N_3,In_1278,In_846);
or U4 (N_4,In_1877,In_2193);
or U5 (N_5,In_737,In_175);
and U6 (N_6,In_300,In_2389);
nand U7 (N_7,In_930,In_1501);
nor U8 (N_8,In_1186,In_901);
or U9 (N_9,In_2354,In_1938);
nor U10 (N_10,In_1604,In_2299);
nand U11 (N_11,In_1512,In_933);
xnor U12 (N_12,In_637,In_1851);
or U13 (N_13,In_2163,In_550);
or U14 (N_14,In_2238,In_2105);
nand U15 (N_15,In_1330,In_1273);
or U16 (N_16,In_345,In_2149);
and U17 (N_17,In_1509,In_1201);
nand U18 (N_18,In_1312,In_993);
nor U19 (N_19,In_1507,In_314);
and U20 (N_20,In_877,In_327);
nor U21 (N_21,In_1136,In_412);
nand U22 (N_22,In_1216,In_114);
nand U23 (N_23,In_1913,In_2378);
nand U24 (N_24,In_1220,In_1022);
and U25 (N_25,In_822,In_889);
and U26 (N_26,In_1716,In_2349);
nor U27 (N_27,In_1609,In_368);
nand U28 (N_28,In_156,In_1556);
nor U29 (N_29,In_376,In_1217);
or U30 (N_30,In_2229,In_2146);
or U31 (N_31,In_1314,In_1385);
and U32 (N_32,In_613,In_1908);
xor U33 (N_33,In_2,In_1031);
nor U34 (N_34,In_2119,In_1516);
or U35 (N_35,In_1171,In_138);
xor U36 (N_36,In_1260,In_633);
xnor U37 (N_37,In_2458,In_639);
or U38 (N_38,In_2380,In_554);
or U39 (N_39,In_1207,In_1652);
or U40 (N_40,In_1193,In_679);
xnor U41 (N_41,In_939,In_869);
nand U42 (N_42,In_1649,In_2322);
xnor U43 (N_43,In_511,In_2414);
and U44 (N_44,In_2196,In_2495);
or U45 (N_45,In_289,In_955);
or U46 (N_46,In_392,In_572);
nand U47 (N_47,In_2474,In_1533);
nor U48 (N_48,In_235,In_2231);
or U49 (N_49,In_951,In_1748);
and U50 (N_50,In_1384,In_2100);
nor U51 (N_51,In_2009,In_1395);
nand U52 (N_52,In_475,In_99);
xor U53 (N_53,In_2168,In_2485);
nand U54 (N_54,In_780,In_1990);
or U55 (N_55,In_1059,In_8);
nor U56 (N_56,In_1676,In_1537);
nand U57 (N_57,In_204,In_984);
and U58 (N_58,In_2092,In_383);
nand U59 (N_59,In_2399,In_2260);
or U60 (N_60,In_1425,In_1788);
or U61 (N_61,In_2138,In_353);
and U62 (N_62,In_295,In_2139);
or U63 (N_63,In_708,In_1576);
nor U64 (N_64,In_784,In_973);
xnor U65 (N_65,In_1398,In_2239);
or U66 (N_66,In_1830,In_233);
or U67 (N_67,In_1873,In_1888);
or U68 (N_68,In_753,In_277);
and U69 (N_69,In_1852,In_723);
xnor U70 (N_70,In_1636,In_1603);
nand U71 (N_71,In_1587,In_1161);
nand U72 (N_72,In_1903,In_570);
nand U73 (N_73,In_1536,In_1165);
and U74 (N_74,In_636,In_2186);
nor U75 (N_75,In_947,In_2407);
nor U76 (N_76,In_1090,In_1051);
nor U77 (N_77,In_1656,In_131);
and U78 (N_78,In_541,In_979);
and U79 (N_79,In_934,In_1701);
and U80 (N_80,In_504,In_1167);
nand U81 (N_81,In_986,In_2262);
nor U82 (N_82,In_1194,In_663);
nor U83 (N_83,In_789,In_528);
or U84 (N_84,In_2377,In_150);
nor U85 (N_85,In_589,In_1381);
nand U86 (N_86,In_1028,In_472);
and U87 (N_87,In_1807,In_688);
nor U88 (N_88,In_583,In_269);
nand U89 (N_89,In_2003,In_2111);
xnor U90 (N_90,In_924,In_2263);
and U91 (N_91,In_555,In_683);
nand U92 (N_92,In_704,In_2405);
nor U93 (N_93,In_749,In_462);
and U94 (N_94,In_196,In_530);
or U95 (N_95,In_1895,In_378);
and U96 (N_96,In_229,In_1783);
nor U97 (N_97,In_1280,In_638);
xnor U98 (N_98,In_518,In_801);
nand U99 (N_99,In_1155,In_140);
nand U100 (N_100,In_744,In_74);
nand U101 (N_101,In_84,In_1885);
nand U102 (N_102,In_592,In_1372);
nand U103 (N_103,In_425,In_1680);
and U104 (N_104,In_1192,In_2490);
and U105 (N_105,In_1729,In_1421);
and U106 (N_106,In_1778,In_1791);
or U107 (N_107,In_1428,In_1099);
or U108 (N_108,In_265,In_574);
nor U109 (N_109,In_241,In_982);
nor U110 (N_110,In_1154,In_1447);
nor U111 (N_111,In_2288,In_426);
and U112 (N_112,In_1756,In_1141);
and U113 (N_113,In_456,In_699);
and U114 (N_114,In_2167,In_398);
or U115 (N_115,In_2128,In_1858);
nor U116 (N_116,In_891,In_1739);
nand U117 (N_117,In_2312,In_1996);
or U118 (N_118,In_367,In_1145);
and U119 (N_119,In_2079,In_2282);
nor U120 (N_120,In_1911,In_1841);
and U121 (N_121,In_1319,In_143);
nand U122 (N_122,In_2123,In_2051);
or U123 (N_123,In_1763,In_1357);
nor U124 (N_124,In_1891,In_498);
or U125 (N_125,In_1005,In_513);
xor U126 (N_126,In_1714,In_1894);
nor U127 (N_127,In_1519,In_1667);
nor U128 (N_128,In_706,In_1724);
or U129 (N_129,In_1003,In_1061);
and U130 (N_130,In_1478,In_2086);
or U131 (N_131,In_1910,In_2426);
and U132 (N_132,In_1387,In_407);
nand U133 (N_133,In_1475,In_1334);
nor U134 (N_134,In_819,In_245);
xor U135 (N_135,In_689,In_51);
and U136 (N_136,In_1488,In_191);
nand U137 (N_137,In_427,In_2004);
nand U138 (N_138,In_2144,In_2434);
nand U139 (N_139,In_1982,In_1538);
xor U140 (N_140,In_348,In_97);
or U141 (N_141,In_2304,In_1709);
nor U142 (N_142,In_595,In_1147);
nand U143 (N_143,In_2291,In_1964);
nor U144 (N_144,In_1310,In_1403);
nand U145 (N_145,In_1534,In_1723);
and U146 (N_146,In_1801,In_1786);
and U147 (N_147,In_1465,In_1438);
nand U148 (N_148,In_57,In_1793);
and U149 (N_149,In_2406,In_1019);
or U150 (N_150,In_2457,In_1721);
nor U151 (N_151,In_1430,In_66);
nor U152 (N_152,In_1076,In_2439);
or U153 (N_153,In_1139,In_2362);
or U154 (N_154,In_1437,In_2479);
and U155 (N_155,In_2258,In_811);
and U156 (N_156,In_1499,In_1074);
and U157 (N_157,In_1320,In_514);
nor U158 (N_158,In_2428,In_1906);
and U159 (N_159,In_697,In_1782);
nor U160 (N_160,In_1711,In_1215);
or U161 (N_161,In_2121,In_1826);
and U162 (N_162,In_1442,In_1287);
and U163 (N_163,In_32,In_2058);
and U164 (N_164,In_1555,In_2190);
xnor U165 (N_165,In_1079,In_296);
or U166 (N_166,In_2171,In_2348);
nand U167 (N_167,In_1566,In_185);
or U168 (N_168,In_2192,In_52);
or U169 (N_169,In_418,In_1175);
or U170 (N_170,In_2256,In_187);
nor U171 (N_171,In_466,In_2325);
or U172 (N_172,In_162,In_2070);
nor U173 (N_173,In_855,In_1941);
or U174 (N_174,In_414,In_611);
or U175 (N_175,In_420,In_1040);
xor U176 (N_176,In_793,In_1408);
nor U177 (N_177,In_2272,In_2037);
nor U178 (N_178,In_112,In_1283);
or U179 (N_179,In_2015,In_506);
nor U180 (N_180,In_146,In_1484);
and U181 (N_181,In_1670,In_573);
nand U182 (N_182,In_1934,In_1106);
nor U183 (N_183,In_2126,In_2316);
or U184 (N_184,In_1869,In_715);
and U185 (N_185,In_1502,In_1993);
nand U186 (N_186,In_206,In_139);
or U187 (N_187,In_109,In_1704);
nor U188 (N_188,In_1084,In_67);
and U189 (N_189,In_642,In_1168);
nor U190 (N_190,In_2363,In_2477);
nand U191 (N_191,In_2131,In_257);
or U192 (N_192,In_728,In_916);
nand U193 (N_193,In_4,In_1285);
or U194 (N_194,In_2129,In_615);
nand U195 (N_195,In_1418,In_1776);
and U196 (N_196,In_929,In_2243);
nor U197 (N_197,In_807,In_534);
nand U198 (N_198,In_2438,In_2374);
nor U199 (N_199,In_1205,In_2041);
nor U200 (N_200,In_2040,In_1848);
nand U201 (N_201,In_2266,In_137);
and U202 (N_202,In_525,In_2227);
nand U203 (N_203,In_1404,In_1020);
nand U204 (N_204,In_803,In_2404);
xnor U205 (N_205,In_135,In_1731);
nand U206 (N_206,In_2077,In_1780);
nand U207 (N_207,In_1270,In_134);
and U208 (N_208,In_1343,In_2455);
xor U209 (N_209,In_765,In_542);
and U210 (N_210,In_1023,In_409);
nor U211 (N_211,In_1586,In_160);
and U212 (N_212,In_658,In_334);
nand U213 (N_213,In_1160,In_813);
nand U214 (N_214,In_856,In_2435);
nor U215 (N_215,In_2491,In_482);
nor U216 (N_216,In_2246,In_1325);
nor U217 (N_217,In_510,In_2027);
or U218 (N_218,In_1230,In_1500);
nor U219 (N_219,In_1151,In_1364);
or U220 (N_220,In_1617,In_323);
and U221 (N_221,In_1640,In_987);
nor U222 (N_222,In_2225,In_2307);
or U223 (N_223,In_339,In_1299);
and U224 (N_224,In_1561,In_1092);
nand U225 (N_225,In_832,In_2463);
or U226 (N_226,In_2493,In_875);
nor U227 (N_227,In_2364,In_349);
or U228 (N_228,In_1865,In_261);
nand U229 (N_229,In_1683,In_1679);
nand U230 (N_230,In_484,In_1541);
nand U231 (N_231,In_577,In_2460);
xnor U232 (N_232,In_2257,In_2013);
nand U233 (N_233,In_870,In_1738);
nor U234 (N_234,In_1011,In_2099);
nand U235 (N_235,In_2392,In_2475);
nor U236 (N_236,In_1091,In_821);
and U237 (N_237,In_2102,In_1305);
nor U238 (N_238,In_1149,In_288);
and U239 (N_239,In_1846,In_707);
nand U240 (N_240,In_106,In_201);
or U241 (N_241,In_606,In_2470);
or U242 (N_242,In_1184,In_1034);
nor U243 (N_243,In_10,In_214);
nor U244 (N_244,In_1813,In_590);
and U245 (N_245,In_2461,In_2413);
or U246 (N_246,In_2076,In_1489);
nor U247 (N_247,In_2172,In_786);
and U248 (N_248,In_851,In_1132);
and U249 (N_249,In_2344,In_2337);
nor U250 (N_250,In_631,In_58);
and U251 (N_251,In_634,In_1871);
nor U252 (N_252,In_491,In_2039);
nand U253 (N_253,In_1613,In_2203);
nor U254 (N_254,In_1815,In_29);
nor U255 (N_255,In_1014,In_2326);
and U256 (N_256,In_2385,In_122);
nor U257 (N_257,In_1915,In_1472);
and U258 (N_258,In_12,In_325);
and U259 (N_259,In_1390,In_1853);
nor U260 (N_260,In_1864,In_1053);
nor U261 (N_261,In_2187,In_655);
nor U262 (N_262,In_792,In_309);
nand U263 (N_263,In_258,In_2133);
or U264 (N_264,In_1703,In_2006);
xnor U265 (N_265,In_665,In_1562);
nand U266 (N_266,In_1420,In_359);
or U267 (N_267,In_1886,In_2499);
or U268 (N_268,In_343,In_2433);
nor U269 (N_269,In_1176,In_2384);
and U270 (N_270,In_698,In_1767);
nand U271 (N_271,In_157,In_1191);
nor U272 (N_272,In_503,In_1834);
or U273 (N_273,In_1570,In_917);
xor U274 (N_274,In_1306,In_649);
nor U275 (N_275,In_1641,In_620);
and U276 (N_276,In_402,In_0);
nand U277 (N_277,In_1542,In_549);
nand U278 (N_278,In_2035,In_1050);
xor U279 (N_279,In_508,In_1309);
nand U280 (N_280,In_810,In_927);
and U281 (N_281,In_531,In_47);
nor U282 (N_282,In_1758,In_213);
or U283 (N_283,In_1263,In_2248);
nand U284 (N_284,In_1203,In_2114);
nor U285 (N_285,In_1648,In_783);
or U286 (N_286,In_2284,In_331);
nand U287 (N_287,In_1629,In_1557);
nor U288 (N_288,In_28,In_886);
and U289 (N_289,In_1219,In_2369);
nand U290 (N_290,In_2062,In_1238);
and U291 (N_291,In_338,In_711);
and U292 (N_292,In_1423,In_918);
nand U293 (N_293,In_820,In_1304);
or U294 (N_294,In_763,In_1083);
or U295 (N_295,In_2209,In_69);
and U296 (N_296,In_2065,In_975);
nor U297 (N_297,In_643,In_2347);
and U298 (N_298,In_238,In_769);
nand U299 (N_299,In_1233,In_1845);
nand U300 (N_300,In_88,In_1605);
or U301 (N_301,In_2210,In_1214);
and U302 (N_302,In_862,In_2289);
or U303 (N_303,In_2101,In_272);
xnor U304 (N_304,In_1735,In_1268);
and U305 (N_305,In_2333,In_1180);
and U306 (N_306,In_564,In_1284);
or U307 (N_307,In_2387,In_226);
nand U308 (N_308,In_833,In_1972);
or U309 (N_309,In_2021,In_2080);
xor U310 (N_310,In_165,In_712);
xor U311 (N_311,In_2498,In_1487);
xor U312 (N_312,In_1409,In_1948);
nand U313 (N_313,In_1627,In_1611);
or U314 (N_314,In_798,In_546);
or U315 (N_315,In_1123,In_1321);
or U316 (N_316,In_120,In_1039);
or U317 (N_317,In_2419,In_533);
nor U318 (N_318,In_785,In_1410);
xnor U319 (N_319,In_2421,In_678);
or U320 (N_320,In_2340,In_1925);
nand U321 (N_321,In_1503,In_2444);
nand U322 (N_322,In_2223,In_1751);
nor U323 (N_323,In_1292,In_2394);
or U324 (N_324,In_492,In_464);
or U325 (N_325,In_1431,In_1980);
and U326 (N_326,In_1955,In_391);
nor U327 (N_327,In_836,In_1961);
or U328 (N_328,In_1497,In_1339);
or U329 (N_329,In_1317,In_2294);
or U330 (N_330,In_687,In_75);
nand U331 (N_331,In_444,In_664);
and U332 (N_332,In_544,In_1986);
xor U333 (N_333,In_1341,In_1921);
nor U334 (N_334,In_2218,In_1101);
nor U335 (N_335,In_455,In_881);
and U336 (N_336,In_867,In_1222);
nand U337 (N_337,In_1875,In_14);
nor U338 (N_338,In_164,In_2306);
or U339 (N_339,In_1819,In_119);
and U340 (N_340,In_1456,In_1480);
nand U341 (N_341,In_2200,In_365);
and U342 (N_342,In_505,In_404);
nor U343 (N_343,In_1063,In_1206);
nand U344 (N_344,In_770,In_1769);
or U345 (N_345,In_1665,In_597);
and U346 (N_346,In_2224,In_1188);
nor U347 (N_347,In_1983,In_1975);
nor U348 (N_348,In_935,In_2450);
nor U349 (N_349,In_92,In_920);
and U350 (N_350,In_1930,In_1042);
nand U351 (N_351,In_1413,In_1804);
nand U352 (N_352,In_796,In_748);
nor U353 (N_353,In_1087,In_1916);
or U354 (N_354,In_1674,In_1415);
or U355 (N_355,In_1086,In_2481);
or U356 (N_356,In_1144,In_250);
nand U357 (N_357,In_2423,In_9);
or U358 (N_358,In_2127,In_2360);
xor U359 (N_359,In_1114,In_1150);
or U360 (N_360,In_2169,In_337);
nor U361 (N_361,In_1368,In_262);
or U362 (N_362,In_757,In_1999);
nor U363 (N_363,In_1594,In_2467);
xnor U364 (N_364,In_2182,In_1839);
and U365 (N_365,In_253,In_270);
nand U366 (N_366,In_1699,In_2356);
and U367 (N_367,In_1505,In_1137);
and U368 (N_368,In_1109,In_805);
nand U369 (N_369,In_188,In_1997);
or U370 (N_370,In_1047,In_61);
and U371 (N_371,In_2270,In_537);
and U372 (N_372,In_2339,In_415);
nand U373 (N_373,In_1717,In_1377);
or U374 (N_374,In_254,In_76);
nand U375 (N_375,In_2221,In_1812);
or U376 (N_376,In_2030,In_690);
nand U377 (N_377,In_411,In_2269);
or U378 (N_378,In_2252,In_1785);
nand U379 (N_379,In_1279,In_701);
or U380 (N_380,In_1863,In_1029);
nor U381 (N_381,In_2352,In_318);
nor U382 (N_382,In_2233,In_63);
or U383 (N_383,In_2409,In_2032);
or U384 (N_384,In_602,In_450);
nor U385 (N_385,In_2343,In_1159);
nand U386 (N_386,In_2478,In_216);
nor U387 (N_387,In_2287,In_1977);
nand U388 (N_388,In_1077,In_1827);
nor U389 (N_389,In_745,In_1467);
and U390 (N_390,In_104,In_676);
nand U391 (N_391,In_950,In_1770);
or U392 (N_392,In_941,In_2247);
nand U393 (N_393,In_1646,In_1295);
xor U394 (N_394,In_1527,In_93);
nor U395 (N_395,In_1244,In_2104);
and U396 (N_396,In_275,In_1590);
nor U397 (N_397,In_1198,In_2156);
or U398 (N_398,In_1379,In_2427);
or U399 (N_399,In_148,In_1790);
and U400 (N_400,In_2267,In_2154);
or U401 (N_401,In_1104,In_995);
nand U402 (N_402,In_860,In_1252);
nand U403 (N_403,In_1441,In_2273);
nor U404 (N_404,In_895,In_1671);
nand U405 (N_405,In_2096,In_2420);
nand U406 (N_406,In_787,In_834);
or U407 (N_407,In_1904,In_40);
nand U408 (N_408,In_46,In_2026);
nor U409 (N_409,In_2120,In_659);
nor U410 (N_410,In_535,In_2355);
nor U411 (N_411,In_2277,In_1985);
xnor U412 (N_412,In_1917,In_1340);
or U413 (N_413,In_2370,In_424);
nor U414 (N_414,In_307,In_2234);
and U415 (N_415,In_536,In_922);
nand U416 (N_416,In_1406,In_149);
nand U417 (N_417,In_1631,In_848);
and U418 (N_418,In_1811,In_1954);
nand U419 (N_419,In_919,In_560);
xnor U420 (N_420,In_661,In_904);
or U421 (N_421,In_685,In_2057);
nor U422 (N_422,In_1752,In_1070);
xnor U423 (N_423,In_1393,In_1315);
and U424 (N_424,In_1152,In_1949);
or U425 (N_425,In_2497,In_2358);
or U426 (N_426,In_893,In_931);
nor U427 (N_427,In_400,In_2314);
or U428 (N_428,In_1522,In_1234);
and U429 (N_429,In_2353,In_2327);
and U430 (N_430,In_2431,In_1157);
or U431 (N_431,In_1197,In_1033);
nand U432 (N_432,In_623,In_1121);
xnor U433 (N_433,In_1380,In_1081);
or U434 (N_434,In_2417,In_1481);
and U435 (N_435,In_111,In_2335);
xnor U436 (N_436,In_1496,In_1932);
nor U437 (N_437,In_561,In_992);
or U438 (N_438,In_2140,In_2432);
and U439 (N_439,In_2046,In_1890);
or U440 (N_440,In_779,In_1324);
and U441 (N_441,In_286,In_872);
nand U442 (N_442,In_1666,In_1902);
and U443 (N_443,In_333,In_2185);
nor U444 (N_444,In_750,In_33);
xor U445 (N_445,In_1066,In_2278);
and U446 (N_446,In_1789,In_865);
and U447 (N_447,In_1318,In_1936);
nand U448 (N_448,In_1598,In_271);
nand U449 (N_449,In_1745,In_815);
or U450 (N_450,In_1470,In_36);
xor U451 (N_451,In_305,In_842);
nand U452 (N_452,In_1589,In_1759);
xor U453 (N_453,In_1392,In_2195);
and U454 (N_454,In_1582,In_167);
and U455 (N_455,In_2328,In_500);
and U456 (N_456,In_2141,In_923);
or U457 (N_457,In_1988,In_2125);
nand U458 (N_458,In_1477,In_1226);
nand U459 (N_459,In_2476,In_2085);
or U460 (N_460,In_1945,In_1432);
and U461 (N_461,In_2115,In_489);
nor U462 (N_462,In_87,In_1148);
nor U463 (N_463,In_2219,In_600);
nand U464 (N_464,In_791,In_2152);
or U465 (N_465,In_512,In_1898);
or U466 (N_466,In_304,In_16);
nand U467 (N_467,In_878,In_351);
and U468 (N_468,In_1417,In_1950);
or U469 (N_469,In_2158,In_1253);
nand U470 (N_470,In_218,In_1134);
nand U471 (N_471,In_553,In_1411);
nor U472 (N_472,In_2401,In_1082);
and U473 (N_473,In_1612,In_961);
nand U474 (N_474,In_645,In_417);
xnor U475 (N_475,In_1600,In_2279);
nand U476 (N_476,In_1228,In_1107);
nand U477 (N_477,In_1588,In_1914);
nor U478 (N_478,In_1998,In_231);
nor U479 (N_479,In_326,In_1227);
or U480 (N_480,In_1897,In_53);
nor U481 (N_481,In_2334,In_1041);
and U482 (N_482,In_2164,In_2285);
and U483 (N_483,In_652,In_1884);
nand U484 (N_484,In_2212,In_1223);
nor U485 (N_485,In_1422,In_189);
or U486 (N_486,In_680,In_746);
nor U487 (N_487,In_2107,In_1169);
nand U488 (N_488,In_1504,In_2173);
and U489 (N_489,In_1013,In_2073);
xnor U490 (N_490,In_2297,In_340);
or U491 (N_491,In_1374,In_255);
nor U492 (N_492,In_999,In_1730);
nand U493 (N_493,In_396,In_1307);
or U494 (N_494,In_1928,In_1221);
nand U495 (N_495,In_567,In_1211);
nand U496 (N_496,In_190,In_1583);
xor U497 (N_497,In_59,In_976);
xnor U498 (N_498,In_2177,In_2117);
or U499 (N_499,In_1337,In_329);
or U500 (N_500,In_50,In_2056);
nor U501 (N_501,In_1524,In_1185);
nor U502 (N_502,In_221,In_390);
and U503 (N_503,In_1981,In_1568);
nor U504 (N_504,In_437,In_863);
nor U505 (N_505,In_1803,In_1784);
xor U506 (N_506,In_171,In_1828);
or U507 (N_507,In_710,In_163);
nor U508 (N_508,In_1199,In_2063);
nand U509 (N_509,In_408,In_1298);
and U510 (N_510,In_911,In_1135);
and U511 (N_511,In_1657,In_1539);
and U512 (N_512,In_2459,In_1049);
and U513 (N_513,In_1030,In_2245);
nand U514 (N_514,In_228,In_1024);
or U515 (N_515,In_960,In_2228);
or U516 (N_516,In_1755,In_1893);
nor U517 (N_517,In_177,In_1016);
nand U518 (N_518,In_476,In_725);
or U519 (N_519,In_648,In_726);
xnor U520 (N_520,In_2010,In_1262);
nor U521 (N_521,In_2388,In_1558);
xor U522 (N_522,In_1650,In_1951);
nor U523 (N_523,In_885,In_985);
or U524 (N_524,In_515,In_635);
and U525 (N_525,In_1847,In_1446);
nand U526 (N_526,In_375,In_1857);
nand U527 (N_527,In_2110,In_670);
or U528 (N_528,In_1599,In_2087);
nand U529 (N_529,In_496,In_465);
nand U530 (N_530,In_152,In_2162);
xor U531 (N_531,In_1045,In_1878);
and U532 (N_532,In_584,In_1057);
nand U533 (N_533,In_155,In_1741);
nor U534 (N_534,In_1844,In_2078);
or U535 (N_535,In_2205,In_1506);
or U536 (N_536,In_804,In_2264);
or U537 (N_537,In_2019,In_1732);
nand U538 (N_538,In_2466,In_308);
or U539 (N_539,In_2148,In_1126);
nor U540 (N_540,In_95,In_1580);
nand U541 (N_541,In_1391,In_1426);
nor U542 (N_542,In_1573,In_98);
or U543 (N_543,In_1495,In_126);
or U544 (N_544,In_847,In_1009);
nor U545 (N_545,In_2329,In_586);
or U546 (N_546,In_2201,In_1743);
nor U547 (N_547,In_656,In_1718);
nand U548 (N_548,In_1771,In_45);
nor U549 (N_549,In_1688,In_2303);
or U550 (N_550,In_1213,In_945);
nand U551 (N_551,In_1055,In_1054);
and U552 (N_552,In_662,In_458);
nand U553 (N_553,In_2254,In_151);
and U554 (N_554,In_1131,In_641);
nand U555 (N_555,In_1529,In_234);
or U556 (N_556,In_2007,In_1697);
nand U557 (N_557,In_2093,In_259);
and U558 (N_558,In_2211,In_1457);
nand U559 (N_559,In_2456,In_1749);
nand U560 (N_560,In_1901,In_1231);
xnor U561 (N_561,In_1461,In_1471);
or U562 (N_562,In_1080,In_762);
or U563 (N_563,In_1143,In_1610);
nor U564 (N_564,In_692,In_207);
or U565 (N_565,In_2235,In_557);
xnor U566 (N_566,In_741,In_994);
xor U567 (N_567,In_37,In_1378);
or U568 (N_568,In_251,In_86);
and U569 (N_569,In_2346,In_1113);
nor U570 (N_570,In_1440,In_71);
or U571 (N_571,In_956,In_1158);
nor U572 (N_572,In_1282,In_943);
xor U573 (N_573,In_423,In_2082);
and U574 (N_574,In_2043,In_363);
xnor U575 (N_575,In_2000,In_284);
xnor U576 (N_576,In_1064,In_1900);
nand U577 (N_577,In_1254,In_1879);
nor U578 (N_578,In_829,In_478);
nor U579 (N_579,In_1336,In_2008);
nand U580 (N_580,In_481,In_2072);
or U581 (N_581,In_603,In_242);
xor U582 (N_582,In_1272,In_1700);
or U583 (N_583,In_1719,In_1968);
nor U584 (N_584,In_1464,In_2098);
and U585 (N_585,In_2445,In_1919);
nor U586 (N_586,In_1351,In_754);
nor U587 (N_587,In_369,In_2342);
nor U588 (N_588,In_115,In_1726);
nor U589 (N_589,In_1311,In_118);
nor U590 (N_590,In_1255,In_520);
nand U591 (N_591,In_1535,In_2020);
nor U592 (N_592,In_1493,In_1127);
nand U593 (N_593,In_1346,In_1363);
xor U594 (N_594,In_2351,In_1822);
nor U595 (N_595,In_1382,In_1693);
or U596 (N_596,In_773,In_1397);
nor U597 (N_597,In_2055,In_282);
nor U598 (N_598,In_806,In_1036);
nor U599 (N_599,In_694,In_1659);
or U600 (N_600,In_1286,In_1814);
and U601 (N_601,In_490,In_2292);
nor U602 (N_602,In_1043,In_1737);
and U603 (N_603,In_2276,In_446);
and U604 (N_604,In_964,In_1883);
and U605 (N_605,In_1643,In_6);
nand U606 (N_606,In_1069,In_2261);
nor U607 (N_607,In_1825,In_2068);
or U608 (N_608,In_113,In_1491);
and U609 (N_609,In_1817,In_103);
nor U610 (N_610,In_225,In_346);
nand U611 (N_611,In_1479,In_1483);
xnor U612 (N_612,In_2017,In_1689);
nor U613 (N_613,In_2044,In_1823);
nand U614 (N_614,In_558,In_970);
xnor U615 (N_615,In_2022,In_581);
nand U616 (N_616,In_1367,In_2298);
nor U617 (N_617,In_1808,In_967);
nand U618 (N_618,In_1725,In_2451);
nand U619 (N_619,In_24,In_882);
nand U620 (N_620,In_907,In_483);
nor U621 (N_621,In_301,In_1232);
or U622 (N_622,In_1551,In_2372);
and U623 (N_623,In_1002,In_438);
and U624 (N_624,In_230,In_1008);
or U625 (N_625,In_1130,In_946);
nor U626 (N_626,In_1035,In_2053);
or U627 (N_627,In_1933,In_2023);
nand U628 (N_628,In_516,In_321);
or U629 (N_629,In_903,In_2415);
and U630 (N_630,In_1052,In_624);
and U631 (N_631,In_208,In_64);
nor U632 (N_632,In_1574,In_601);
nor U633 (N_633,In_1521,In_1246);
or U634 (N_634,In_540,In_1125);
and U635 (N_635,In_1492,In_1929);
or U636 (N_636,In_1655,In_980);
xnor U637 (N_637,In_782,In_1806);
or U638 (N_638,In_666,In_341);
nand U639 (N_639,In_1829,In_480);
and U640 (N_640,In_2265,In_448);
or U641 (N_641,In_2014,In_2308);
nand U642 (N_642,In_125,In_1436);
or U643 (N_643,In_2489,In_2400);
nor U644 (N_644,In_2130,In_1510);
and U645 (N_645,In_607,In_852);
xnor U646 (N_646,In_1638,In_2472);
or U647 (N_647,In_2207,In_2183);
and U648 (N_648,In_729,In_279);
nand U649 (N_649,In_2170,In_1098);
nor U650 (N_650,In_358,In_1623);
nand U651 (N_651,In_145,In_921);
or U652 (N_652,In_866,In_2052);
and U653 (N_653,In_1448,In_1530);
or U654 (N_654,In_2331,In_1335);
or U655 (N_655,In_361,In_1563);
nor U656 (N_656,In_1698,In_1443);
and U657 (N_657,In_890,In_2050);
xnor U658 (N_658,In_335,In_2382);
nand U659 (N_659,In_1235,In_1577);
nor U660 (N_660,In_72,In_1249);
nand U661 (N_661,In_580,In_1660);
xor U662 (N_662,In_2398,In_182);
and U663 (N_663,In_2106,In_2134);
nand U664 (N_664,In_320,In_62);
and U665 (N_665,In_1918,In_1018);
nand U666 (N_666,In_605,In_2402);
nand U667 (N_667,In_669,In_1178);
nand U668 (N_668,In_174,In_826);
or U669 (N_669,In_445,In_7);
and U670 (N_670,In_25,In_110);
or U671 (N_671,In_610,In_897);
and U672 (N_672,In_355,In_2109);
and U673 (N_673,In_102,In_366);
or U674 (N_674,In_521,In_1969);
xnor U675 (N_675,In_1606,In_1559);
and U676 (N_676,In_1707,In_1747);
nand U677 (N_677,In_827,In_1662);
nand U678 (N_678,In_1552,In_1722);
or U679 (N_679,In_1687,In_1181);
nor U680 (N_680,In_1354,In_733);
or U681 (N_681,In_1237,In_1820);
and U682 (N_682,In_101,In_200);
xor U683 (N_683,In_2159,In_681);
nand U684 (N_684,In_2330,In_399);
xnor U685 (N_685,In_2112,In_2029);
xnor U686 (N_686,In_925,In_117);
nand U687 (N_687,In_2301,In_302);
nor U688 (N_688,In_562,In_1518);
or U689 (N_689,In_1241,In_2259);
nand U690 (N_690,In_760,In_1275);
or U691 (N_691,In_2249,In_566);
nor U692 (N_692,In_35,In_1172);
or U693 (N_693,In_1245,In_1469);
and U694 (N_694,In_1153,In_1289);
nor U695 (N_695,In_705,In_1460);
nand U696 (N_696,In_565,In_654);
or U697 (N_697,In_432,In_332);
or U698 (N_698,In_1764,In_1912);
or U699 (N_699,In_790,In_2084);
nand U700 (N_700,In_374,In_1026);
nand U701 (N_701,In_2274,In_1366);
or U702 (N_702,In_2160,In_1694);
and U703 (N_703,In_2180,In_388);
nor U704 (N_704,In_617,In_342);
xor U705 (N_705,In_1994,In_2375);
nand U706 (N_706,In_1463,In_39);
nand U707 (N_707,In_2145,In_227);
and U708 (N_708,In_285,In_1957);
nand U709 (N_709,In_387,In_1797);
or U710 (N_710,In_1360,In_1291);
nand U711 (N_711,In_1445,In_381);
xnor U712 (N_712,In_1971,In_2066);
or U713 (N_713,In_91,In_1177);
nor U714 (N_714,In_1250,In_463);
nor U715 (N_715,In_273,In_2064);
nand U716 (N_716,In_884,In_1297);
xnor U717 (N_717,In_290,In_1001);
nand U718 (N_718,In_1264,In_1596);
or U719 (N_719,In_1359,In_60);
xor U720 (N_720,In_203,In_718);
and U721 (N_721,In_2373,In_1862);
nor U722 (N_722,In_1787,In_1007);
and U723 (N_723,In_2309,In_1427);
nand U724 (N_724,In_1708,In_1710);
nor U725 (N_725,In_1316,In_2324);
and U726 (N_726,In_291,In_618);
and U727 (N_727,In_1338,In_209);
nor U728 (N_728,In_479,In_1628);
nor U729 (N_729,In_1062,In_1622);
nand U730 (N_730,In_1164,In_1058);
nor U731 (N_731,In_1247,In_828);
nor U732 (N_732,In_394,In_2396);
or U733 (N_733,In_1474,In_2336);
nor U734 (N_734,In_599,In_1096);
or U735 (N_735,In_575,In_859);
nor U736 (N_736,In_2403,In_168);
nand U737 (N_737,In_1774,In_494);
or U738 (N_738,In_2202,In_236);
or U739 (N_739,In_263,In_319);
nand U740 (N_740,In_1116,In_2090);
nor U741 (N_741,In_1508,In_1124);
and U742 (N_742,In_702,In_2395);
xor U743 (N_743,In_2213,In_2113);
or U744 (N_744,In_1386,In_2317);
xnor U745 (N_745,In_2188,In_991);
or U746 (N_746,In_2184,In_1239);
nand U747 (N_747,In_1927,In_2208);
nor U748 (N_748,In_667,In_1088);
xor U749 (N_749,In_1965,In_766);
xnor U750 (N_750,In_2089,In_914);
and U751 (N_751,In_1672,In_401);
nand U752 (N_752,In_1344,In_2416);
nand U753 (N_753,In_1429,In_141);
or U754 (N_754,In_596,In_1715);
nor U755 (N_755,In_1021,In_1290);
nand U756 (N_756,In_2341,In_195);
nor U757 (N_757,In_1943,In_1620);
or U758 (N_758,In_1585,In_1740);
nand U759 (N_759,In_632,In_1696);
nor U760 (N_760,In_347,In_988);
nor U761 (N_761,In_2280,In_2199);
nor U762 (N_762,In_912,In_854);
nand U763 (N_763,In_626,In_684);
xor U764 (N_764,In_1766,In_868);
or U765 (N_765,In_79,In_127);
or U766 (N_766,In_1685,In_1944);
nand U767 (N_767,In_1094,In_193);
nand U768 (N_768,In_280,In_178);
xnor U769 (N_769,In_240,In_640);
xnor U770 (N_770,In_344,In_2147);
or U771 (N_771,In_2217,In_1251);
or U772 (N_772,In_1532,In_1303);
and U773 (N_773,In_845,In_1615);
nand U774 (N_774,In_199,In_1753);
nand U775 (N_775,In_2124,In_952);
or U776 (N_776,In_1112,In_313);
or U777 (N_777,In_501,In_77);
nand U778 (N_778,In_1103,In_880);
nor U779 (N_779,In_1525,In_978);
or U780 (N_780,In_31,In_1405);
nand U781 (N_781,In_2033,In_817);
xnor U782 (N_782,In_244,In_389);
nand U783 (N_783,In_153,In_1179);
nor U784 (N_784,In_591,In_1433);
or U785 (N_785,In_159,In_1402);
or U786 (N_786,In_926,In_421);
or U787 (N_787,In_1905,In_2425);
and U788 (N_788,In_972,In_2095);
or U789 (N_789,In_874,In_630);
or U790 (N_790,In_2045,In_1772);
or U791 (N_791,In_2338,In_1089);
nor U792 (N_792,In_1742,In_2320);
or U793 (N_793,In_2230,In_808);
nand U794 (N_794,In_1695,In_1449);
nor U795 (N_795,In_350,In_1809);
or U796 (N_796,In_416,In_915);
or U797 (N_797,In_1810,In_700);
or U798 (N_798,In_747,In_2059);
nand U799 (N_799,In_2002,In_354);
or U800 (N_800,In_823,In_2462);
or U801 (N_801,In_1342,In_1399);
or U802 (N_802,In_2366,In_2094);
or U803 (N_803,In_2103,In_2232);
nor U804 (N_804,In_2465,In_551);
or U805 (N_805,In_453,In_322);
and U806 (N_806,In_49,In_1816);
or U807 (N_807,In_772,In_981);
and U808 (N_808,In_2253,In_1240);
nor U809 (N_809,In_1383,In_2244);
nand U810 (N_810,In_1775,In_1097);
nand U811 (N_811,In_41,In_1085);
and U812 (N_812,In_1601,In_1684);
nand U813 (N_813,In_2155,In_1434);
and U814 (N_814,In_799,In_1133);
and U815 (N_815,In_2204,In_1195);
or U816 (N_816,In_1108,In_1242);
nor U817 (N_817,In_1453,In_1872);
or U818 (N_818,In_1924,In_1373);
and U819 (N_819,In_1625,In_756);
or U820 (N_820,In_1760,In_1117);
or U821 (N_821,In_297,In_2430);
or U822 (N_822,In_406,In_357);
xnor U823 (N_823,In_1750,In_651);
and U824 (N_824,In_1000,In_1881);
nor U825 (N_825,In_166,In_205);
and U826 (N_826,In_2386,In_2024);
nor U827 (N_827,In_1713,In_128);
and U828 (N_828,In_1956,In_1328);
nand U829 (N_829,In_65,In_13);
nor U830 (N_830,In_1992,In_1329);
or U831 (N_831,In_30,In_2468);
nor U832 (N_832,In_1553,In_1974);
nor U833 (N_833,In_1302,In_1435);
nor U834 (N_834,In_898,In_2496);
and U835 (N_835,In_2393,In_385);
nand U836 (N_836,In_1332,In_1880);
nor U837 (N_837,In_543,In_2486);
and U838 (N_838,In_627,In_502);
nor U839 (N_839,In_614,In_998);
nand U840 (N_840,In_547,In_1038);
nand U841 (N_841,In_1543,In_1182);
nand U842 (N_842,In_22,In_136);
or U843 (N_843,In_2220,In_751);
or U844 (N_844,In_1935,In_1651);
xnor U845 (N_845,In_714,In_966);
and U846 (N_846,In_2137,In_1591);
and U847 (N_847,In_317,In_644);
or U848 (N_848,In_1746,In_1229);
and U849 (N_849,In_15,In_397);
nand U850 (N_850,In_243,In_1068);
or U851 (N_851,In_1269,In_1854);
nand U852 (N_852,In_430,In_1668);
and U853 (N_853,In_1485,In_835);
nor U854 (N_854,In_2319,In_1850);
and U855 (N_855,In_936,In_671);
and U856 (N_856,In_1,In_2189);
nor U857 (N_857,In_2367,In_585);
nor U858 (N_858,In_814,In_858);
or U859 (N_859,In_183,In_371);
nand U860 (N_860,In_2226,In_1396);
or U861 (N_861,In_1736,In_2166);
xnor U862 (N_862,In_686,In_899);
nor U863 (N_863,In_2390,In_433);
and U864 (N_864,In_1976,In_675);
and U865 (N_865,In_169,In_695);
nand U866 (N_866,In_2067,In_1632);
nand U867 (N_867,In_278,In_260);
nand U868 (N_868,In_224,In_2240);
nor U869 (N_869,In_1773,In_2005);
nand U870 (N_870,In_186,In_1189);
xor U871 (N_871,In_1248,In_1937);
xnor U872 (N_872,In_871,In_730);
xnor U873 (N_873,In_21,In_1838);
nor U874 (N_874,In_1712,In_2452);
xnor U875 (N_875,In_1190,In_850);
or U876 (N_876,In_1560,In_1056);
and U877 (N_877,In_778,In_2376);
nand U878 (N_878,In_1006,In_1032);
and U879 (N_879,In_2464,In_682);
nor U880 (N_880,In_460,In_1313);
nor U881 (N_881,In_1037,In_1115);
nand U882 (N_882,In_1486,In_1407);
and U883 (N_883,In_2482,In_857);
or U884 (N_884,In_548,In_1208);
xor U885 (N_885,In_1547,In_55);
xnor U886 (N_886,In_957,In_11);
or U887 (N_887,In_1892,In_1909);
xor U888 (N_888,In_2454,In_443);
and U889 (N_889,In_552,In_816);
nand U890 (N_890,In_1523,In_194);
and U891 (N_891,In_287,In_902);
or U892 (N_892,In_2441,In_1138);
and U893 (N_893,In_2178,In_252);
nor U894 (N_894,In_1682,In_1110);
nor U895 (N_895,In_2488,In_1958);
nor U896 (N_896,In_198,In_1567);
nor U897 (N_897,In_1170,In_1323);
nor U898 (N_898,In_1276,In_1705);
and U899 (N_899,In_497,In_1633);
nor U900 (N_900,In_764,In_26);
and U901 (N_901,In_468,In_556);
nand U902 (N_902,In_1920,In_1706);
nor U903 (N_903,In_219,In_905);
or U904 (N_904,In_1597,In_2150);
nor U905 (N_905,In_1414,In_2332);
xor U906 (N_906,In_619,In_360);
nor U907 (N_907,In_2449,In_974);
nor U908 (N_908,In_2097,In_410);
and U909 (N_909,In_1690,In_1837);
xor U910 (N_910,In_161,In_1616);
nor U911 (N_911,In_1754,In_173);
or U912 (N_912,In_1867,In_1779);
nand U913 (N_913,In_1122,In_900);
nor U914 (N_914,In_202,In_1637);
nor U915 (N_915,In_713,In_1579);
xor U916 (N_916,In_657,In_267);
nor U917 (N_917,In_1048,In_2061);
and U918 (N_918,In_906,In_256);
nand U919 (N_919,In_2484,In_1960);
or U920 (N_920,In_691,In_1347);
and U921 (N_921,In_303,In_1842);
nor U922 (N_922,In_1855,In_539);
or U923 (N_923,In_1288,In_330);
and U924 (N_924,In_1129,In_246);
nand U925 (N_925,In_1451,In_887);
nand U926 (N_926,In_1658,In_1102);
nand U927 (N_927,In_133,In_80);
and U928 (N_928,In_1762,In_2321);
nand U929 (N_929,In_1162,In_2318);
or U930 (N_930,In_1119,In_954);
nor U931 (N_931,In_429,In_740);
nor U932 (N_932,In_2012,In_1991);
or U933 (N_933,In_440,In_1571);
xor U934 (N_934,In_2161,In_721);
nor U935 (N_935,In_292,In_1365);
or U936 (N_936,In_616,In_434);
or U937 (N_937,In_2311,In_2060);
xnor U938 (N_938,In_576,In_170);
nand U939 (N_939,In_940,In_2036);
nor U940 (N_940,In_1966,In_1513);
nor U941 (N_941,In_1095,In_1870);
nor U942 (N_942,In_2295,In_2487);
nand U943 (N_943,In_2088,In_2191);
nand U944 (N_944,In_1293,In_2241);
or U945 (N_945,In_1326,In_364);
nor U946 (N_946,In_1962,In_1602);
xnor U947 (N_947,In_2174,In_1528);
or U948 (N_948,In_738,In_538);
nor U949 (N_949,In_1899,In_1261);
xnor U950 (N_950,In_1271,In_1868);
xor U951 (N_951,In_1946,In_1836);
nand U952 (N_952,In_1459,In_1120);
or U953 (N_953,In_1979,In_477);
or U954 (N_954,In_393,In_27);
and U955 (N_955,In_1970,In_1482);
nand U956 (N_956,In_2176,In_248);
and U957 (N_957,In_68,In_428);
or U958 (N_958,In_1210,In_743);
or U959 (N_959,In_176,In_217);
or U960 (N_960,In_522,In_264);
and U961 (N_961,In_1452,In_2165);
nand U962 (N_962,In_767,In_1277);
and U963 (N_963,In_1661,In_578);
nor U964 (N_964,In_732,In_442);
nand U965 (N_965,In_294,In_910);
or U966 (N_966,In_469,In_2296);
or U967 (N_967,In_647,In_1923);
nand U968 (N_968,In_2492,In_1677);
or U969 (N_969,In_1196,In_315);
nor U970 (N_970,In_1624,In_1256);
and U971 (N_971,In_519,In_1224);
nand U972 (N_972,In_1835,In_274);
nand U973 (N_973,In_1926,In_2038);
and U974 (N_974,In_1554,In_1727);
and U975 (N_975,In_1569,In_281);
nand U976 (N_976,In_384,In_1266);
or U977 (N_977,In_395,In_673);
nand U978 (N_978,In_1744,In_1520);
nor U979 (N_979,In_268,In_1067);
xnor U980 (N_980,In_569,In_959);
or U981 (N_981,In_849,In_2275);
nand U982 (N_982,In_800,In_100);
nor U983 (N_983,In_1371,In_1202);
or U984 (N_984,In_2047,In_18);
nor U985 (N_985,In_2028,In_1963);
and U986 (N_986,In_1673,In_1078);
nor U987 (N_987,In_1866,In_1375);
or U988 (N_988,In_2091,In_44);
nand U989 (N_989,In_660,In_1345);
nand U990 (N_990,In_2365,In_1889);
nor U991 (N_991,In_2081,In_837);
nor U992 (N_992,In_2071,In_1781);
and U993 (N_993,In_629,In_2300);
or U994 (N_994,In_953,In_2323);
nand U995 (N_995,In_298,In_422);
nor U996 (N_996,In_2132,In_1140);
and U997 (N_997,In_1947,In_894);
or U998 (N_998,In_742,In_132);
nand U999 (N_999,In_2151,In_646);
and U1000 (N_1000,In_1859,In_124);
nand U1001 (N_1001,In_1768,In_2175);
nor U1002 (N_1002,In_1012,In_1301);
xor U1003 (N_1003,In_1355,In_1073);
nor U1004 (N_1004,In_938,In_2237);
and U1005 (N_1005,In_1973,In_2075);
or U1006 (N_1006,In_2251,In_2424);
or U1007 (N_1007,In_1548,In_379);
nand U1008 (N_1008,In_154,In_19);
or U1009 (N_1009,In_788,In_838);
nand U1010 (N_1010,In_1653,In_276);
nand U1011 (N_1011,In_1333,In_853);
or U1012 (N_1012,In_2042,In_720);
and U1013 (N_1013,In_1515,In_2083);
nand U1014 (N_1014,In_17,In_768);
or U1015 (N_1015,In_212,In_668);
nor U1016 (N_1016,In_755,In_759);
and U1017 (N_1017,In_1896,In_2198);
nand U1018 (N_1018,In_831,In_781);
nand U1019 (N_1019,In_2293,In_1296);
nor U1020 (N_1020,In_1308,In_1348);
or U1021 (N_1021,In_677,In_123);
or U1022 (N_1022,In_794,In_1907);
nor U1023 (N_1023,In_693,In_2397);
or U1024 (N_1024,In_1204,In_1540);
and U1025 (N_1025,In_942,In_722);
nor U1026 (N_1026,In_948,In_1821);
xor U1027 (N_1027,In_735,In_211);
or U1028 (N_1028,In_1531,In_386);
or U1029 (N_1029,In_2422,In_604);
and U1030 (N_1030,In_1876,In_1394);
or U1031 (N_1031,In_1128,In_2436);
and U1032 (N_1032,In_559,In_1544);
nor U1033 (N_1033,In_493,In_454);
or U1034 (N_1034,In_777,In_2448);
nand U1035 (N_1035,In_1614,In_1225);
nand U1036 (N_1036,In_1840,In_517);
xor U1037 (N_1037,In_1630,In_523);
nand U1038 (N_1038,In_73,In_179);
or U1039 (N_1039,In_526,In_840);
xnor U1040 (N_1040,In_2383,In_650);
nand U1041 (N_1041,In_2412,In_474);
nor U1042 (N_1042,In_824,In_937);
and U1043 (N_1043,In_529,In_266);
and U1044 (N_1044,In_239,In_2215);
xor U1045 (N_1045,In_172,In_1369);
nor U1046 (N_1046,In_2480,In_1065);
or U1047 (N_1047,In_372,In_830);
nor U1048 (N_1048,In_989,In_215);
and U1049 (N_1049,In_1118,In_1546);
nor U1050 (N_1050,In_1856,In_1952);
nor U1051 (N_1051,In_587,In_996);
nand U1052 (N_1052,In_1644,In_2286);
or U1053 (N_1053,In_293,In_144);
nor U1054 (N_1054,In_1831,In_1978);
or U1055 (N_1055,In_2206,In_1075);
nor U1056 (N_1056,In_2381,In_622);
or U1057 (N_1057,In_844,In_2418);
nor U1058 (N_1058,In_1794,In_1327);
nor U1059 (N_1059,In_311,In_594);
xor U1060 (N_1060,In_1578,In_2122);
nor U1061 (N_1061,In_1468,In_1322);
or U1062 (N_1062,In_724,In_1362);
nor U1063 (N_1063,In_545,In_983);
and U1064 (N_1064,In_247,In_1798);
xnor U1065 (N_1065,In_2411,In_2034);
nor U1066 (N_1066,In_461,In_1691);
nand U1067 (N_1067,In_1494,In_965);
nor U1068 (N_1068,In_38,In_2408);
and U1069 (N_1069,In_1654,In_81);
or U1070 (N_1070,In_2074,In_1412);
nand U1071 (N_1071,In_1874,In_1581);
and U1072 (N_1072,In_23,In_1669);
xor U1073 (N_1073,In_405,In_795);
and U1074 (N_1074,In_2368,In_696);
nand U1075 (N_1075,In_83,In_1142);
nand U1076 (N_1076,In_876,In_734);
nor U1077 (N_1077,In_1458,In_752);
xor U1078 (N_1078,In_719,In_1281);
nand U1079 (N_1079,In_608,In_181);
nand U1080 (N_1080,In_377,In_413);
nand U1081 (N_1081,In_1156,In_1401);
nand U1082 (N_1082,In_2310,In_1639);
xnor U1083 (N_1083,In_2216,In_373);
and U1084 (N_1084,In_2157,In_362);
or U1085 (N_1085,In_1200,In_403);
nand U1086 (N_1086,In_2357,In_452);
or U1087 (N_1087,In_1607,In_1989);
nand U1088 (N_1088,In_1795,In_1111);
or U1089 (N_1089,In_1439,In_2494);
and U1090 (N_1090,In_237,In_89);
or U1091 (N_1091,In_1565,In_1664);
nor U1092 (N_1092,In_593,In_1100);
nand U1093 (N_1093,In_1642,In_1675);
xnor U1094 (N_1094,In_1681,In_2153);
and U1095 (N_1095,In_249,In_2443);
nor U1096 (N_1096,In_43,In_571);
xnor U1097 (N_1097,In_324,In_873);
nand U1098 (N_1098,In_130,In_1584);
xor U1099 (N_1099,In_563,In_879);
xor U1100 (N_1100,In_96,In_1358);
nor U1101 (N_1101,In_1173,In_1361);
nor U1102 (N_1102,In_971,In_1843);
xor U1103 (N_1103,In_439,In_5);
nand U1104 (N_1104,In_1824,In_451);
or U1105 (N_1105,In_1267,In_158);
and U1106 (N_1106,In_2001,In_306);
and U1107 (N_1107,In_1564,In_2345);
nand U1108 (N_1108,In_776,In_1647);
nor U1109 (N_1109,In_2197,In_105);
nor U1110 (N_1110,In_486,In_192);
nand U1111 (N_1111,In_968,In_1450);
or U1112 (N_1112,In_312,In_436);
nand U1113 (N_1113,In_449,In_1490);
and U1114 (N_1114,In_1595,In_2446);
and U1115 (N_1115,In_1645,In_283);
or U1116 (N_1116,In_1931,In_1887);
nand U1117 (N_1117,In_568,In_499);
nor U1118 (N_1118,In_1550,In_1959);
and U1119 (N_1119,In_1350,In_818);
and U1120 (N_1120,In_2118,In_1400);
or U1121 (N_1121,In_1734,In_370);
nor U1122 (N_1122,In_2442,In_2222);
xnor U1123 (N_1123,In_2410,In_441);
xnor U1124 (N_1124,In_147,In_1163);
or U1125 (N_1125,In_1987,In_310);
or U1126 (N_1126,In_316,In_129);
nand U1127 (N_1127,In_1618,In_485);
nand U1128 (N_1128,In_1511,In_1004);
xor U1129 (N_1129,In_2361,In_108);
nor U1130 (N_1130,In_1060,In_2236);
nor U1131 (N_1131,In_1765,In_457);
or U1132 (N_1132,In_797,In_928);
nor U1133 (N_1133,In_1995,In_2049);
or U1134 (N_1134,In_1984,In_2069);
or U1135 (N_1135,In_1849,In_716);
or U1136 (N_1136,In_2135,In_1545);
or U1137 (N_1137,In_579,In_2268);
nor U1138 (N_1138,In_771,In_609);
nand U1139 (N_1139,In_932,In_1462);
nor U1140 (N_1140,In_2447,In_2359);
xnor U1141 (N_1141,In_1592,In_1967);
and U1142 (N_1142,In_2108,In_588);
nor U1143 (N_1143,In_621,In_1455);
and U1144 (N_1144,In_1236,In_527);
nor U1145 (N_1145,In_1071,In_1174);
nor U1146 (N_1146,In_82,In_1860);
or U1147 (N_1147,In_625,In_1800);
nand U1148 (N_1148,In_809,In_2283);
nand U1149 (N_1149,In_1796,In_1444);
nor U1150 (N_1150,In_2179,In_598);
nor U1151 (N_1151,In_222,In_864);
and U1152 (N_1152,In_495,In_184);
or U1153 (N_1153,In_892,In_736);
xor U1154 (N_1154,In_2290,In_524);
nor U1155 (N_1155,In_220,In_1072);
nor U1156 (N_1156,In_85,In_356);
nand U1157 (N_1157,In_2143,In_487);
xor U1158 (N_1158,In_1093,In_2469);
nand U1159 (N_1159,In_703,In_672);
nand U1160 (N_1160,In_825,In_1212);
nor U1161 (N_1161,In_419,In_1692);
nor U1162 (N_1162,In_380,In_1243);
nor U1163 (N_1163,In_913,In_509);
nor U1164 (N_1164,In_2483,In_78);
and U1165 (N_1165,In_2194,In_2371);
nand U1166 (N_1166,In_507,In_299);
or U1167 (N_1167,In_1733,In_2453);
xnor U1168 (N_1168,In_1818,In_1044);
nor U1169 (N_1169,In_1939,In_1833);
or U1170 (N_1170,In_1025,In_1861);
xor U1171 (N_1171,In_944,In_990);
and U1172 (N_1172,In_1300,In_431);
or U1173 (N_1173,In_532,In_1218);
nand U1174 (N_1174,In_223,In_116);
or U1175 (N_1175,In_1608,In_1942);
nor U1176 (N_1176,In_1832,In_2136);
nor U1177 (N_1177,In_997,In_1046);
nor U1178 (N_1178,In_90,In_1792);
nor U1179 (N_1179,In_1353,In_2429);
nor U1180 (N_1180,In_1376,In_473);
and U1181 (N_1181,In_352,In_1526);
nand U1182 (N_1182,In_2214,In_1686);
nand U1183 (N_1183,In_962,In_2181);
nand U1184 (N_1184,In_2391,In_2011);
or U1185 (N_1185,In_2440,In_2281);
and U1186 (N_1186,In_739,In_54);
nor U1187 (N_1187,In_775,In_142);
or U1188 (N_1188,In_3,In_1294);
or U1189 (N_1189,In_1757,In_2379);
nand U1190 (N_1190,In_328,In_1498);
nand U1191 (N_1191,In_1265,In_1621);
or U1192 (N_1192,In_197,In_70);
or U1193 (N_1193,In_1466,In_582);
and U1194 (N_1194,In_2473,In_470);
and U1195 (N_1195,In_467,In_977);
and U1196 (N_1196,In_1370,In_1209);
and U1197 (N_1197,In_843,In_2250);
or U1198 (N_1198,In_1634,In_2271);
or U1199 (N_1199,In_2350,In_727);
and U1200 (N_1200,In_435,In_1331);
nand U1201 (N_1201,In_841,In_674);
xor U1202 (N_1202,In_861,In_1728);
and U1203 (N_1203,In_471,In_1017);
nand U1204 (N_1204,In_382,In_1799);
or U1205 (N_1205,In_1805,In_1146);
nand U1206 (N_1206,In_2016,In_1619);
nor U1207 (N_1207,In_34,In_949);
nor U1208 (N_1208,In_1259,In_1575);
or U1209 (N_1209,In_1702,In_1882);
xnor U1210 (N_1210,In_612,In_839);
nand U1211 (N_1211,In_20,In_774);
nor U1212 (N_1212,In_232,In_459);
nand U1213 (N_1213,In_908,In_1352);
nor U1214 (N_1214,In_2048,In_56);
nor U1215 (N_1215,In_447,In_336);
xnor U1216 (N_1216,In_1257,In_2018);
xor U1217 (N_1217,In_2305,In_488);
or U1218 (N_1218,In_2471,In_1802);
and U1219 (N_1219,In_1388,In_709);
nand U1220 (N_1220,In_107,In_1473);
or U1221 (N_1221,In_812,In_48);
nand U1222 (N_1222,In_1419,In_1940);
or U1223 (N_1223,In_1454,In_1274);
nand U1224 (N_1224,In_1476,In_731);
nor U1225 (N_1225,In_1010,In_2302);
nor U1226 (N_1226,In_1356,In_802);
nand U1227 (N_1227,In_2313,In_2315);
nor U1228 (N_1228,In_1678,In_896);
or U1229 (N_1229,In_1635,In_2031);
xnor U1230 (N_1230,In_717,In_1187);
and U1231 (N_1231,In_42,In_1572);
nor U1232 (N_1232,In_1258,In_963);
nor U1233 (N_1233,In_1166,In_888);
and U1234 (N_1234,In_1183,In_2054);
or U1235 (N_1235,In_2437,In_1424);
and U1236 (N_1236,In_1015,In_180);
or U1237 (N_1237,In_969,In_1626);
or U1238 (N_1238,In_883,In_1761);
nor U1239 (N_1239,In_1517,In_1349);
nor U1240 (N_1240,In_1514,In_210);
nand U1241 (N_1241,In_758,In_2025);
or U1242 (N_1242,In_2142,In_1953);
xor U1243 (N_1243,In_121,In_909);
nor U1244 (N_1244,In_761,In_1549);
nand U1245 (N_1245,In_1105,In_1389);
or U1246 (N_1246,In_1663,In_2242);
nor U1247 (N_1247,In_628,In_2116);
and U1248 (N_1248,In_2255,In_1416);
or U1249 (N_1249,In_958,In_653);
and U1250 (N_1250,In_2289,In_2331);
xor U1251 (N_1251,In_1207,In_2025);
or U1252 (N_1252,In_1706,In_26);
nor U1253 (N_1253,In_217,In_1051);
nand U1254 (N_1254,In_1469,In_921);
nor U1255 (N_1255,In_2034,In_2046);
nand U1256 (N_1256,In_338,In_1791);
or U1257 (N_1257,In_1766,In_1930);
and U1258 (N_1258,In_1254,In_277);
and U1259 (N_1259,In_1622,In_1965);
and U1260 (N_1260,In_2009,In_1295);
and U1261 (N_1261,In_1604,In_1103);
or U1262 (N_1262,In_244,In_676);
or U1263 (N_1263,In_2449,In_210);
and U1264 (N_1264,In_528,In_852);
nand U1265 (N_1265,In_451,In_576);
nor U1266 (N_1266,In_845,In_2020);
and U1267 (N_1267,In_2240,In_1712);
and U1268 (N_1268,In_1617,In_1857);
xor U1269 (N_1269,In_174,In_624);
or U1270 (N_1270,In_1648,In_1409);
nand U1271 (N_1271,In_946,In_1194);
or U1272 (N_1272,In_2112,In_1612);
and U1273 (N_1273,In_773,In_1122);
or U1274 (N_1274,In_2238,In_690);
nor U1275 (N_1275,In_497,In_2200);
and U1276 (N_1276,In_1321,In_2094);
xor U1277 (N_1277,In_2468,In_1571);
xor U1278 (N_1278,In_412,In_126);
nand U1279 (N_1279,In_1110,In_1611);
or U1280 (N_1280,In_745,In_1729);
nand U1281 (N_1281,In_1924,In_982);
or U1282 (N_1282,In_1252,In_372);
and U1283 (N_1283,In_2208,In_797);
xnor U1284 (N_1284,In_476,In_1376);
nor U1285 (N_1285,In_2427,In_527);
nand U1286 (N_1286,In_1354,In_1379);
or U1287 (N_1287,In_2348,In_1954);
nand U1288 (N_1288,In_1282,In_177);
and U1289 (N_1289,In_441,In_2281);
and U1290 (N_1290,In_2068,In_2172);
or U1291 (N_1291,In_124,In_1649);
or U1292 (N_1292,In_2092,In_56);
and U1293 (N_1293,In_772,In_1628);
nand U1294 (N_1294,In_1612,In_1383);
or U1295 (N_1295,In_2213,In_1933);
or U1296 (N_1296,In_1793,In_718);
xnor U1297 (N_1297,In_2312,In_1936);
or U1298 (N_1298,In_1897,In_1479);
and U1299 (N_1299,In_1191,In_1406);
nor U1300 (N_1300,In_1388,In_1030);
nand U1301 (N_1301,In_1661,In_1922);
or U1302 (N_1302,In_383,In_2293);
or U1303 (N_1303,In_12,In_1672);
nor U1304 (N_1304,In_1655,In_1552);
xor U1305 (N_1305,In_103,In_0);
and U1306 (N_1306,In_1667,In_1923);
nor U1307 (N_1307,In_394,In_250);
nor U1308 (N_1308,In_2497,In_939);
or U1309 (N_1309,In_880,In_240);
nor U1310 (N_1310,In_1659,In_939);
nand U1311 (N_1311,In_477,In_2096);
nand U1312 (N_1312,In_2476,In_127);
nor U1313 (N_1313,In_612,In_466);
and U1314 (N_1314,In_267,In_93);
and U1315 (N_1315,In_261,In_355);
or U1316 (N_1316,In_1292,In_1945);
and U1317 (N_1317,In_482,In_1812);
or U1318 (N_1318,In_1908,In_956);
xor U1319 (N_1319,In_1087,In_134);
or U1320 (N_1320,In_1699,In_1730);
nand U1321 (N_1321,In_1131,In_1550);
nor U1322 (N_1322,In_1085,In_224);
or U1323 (N_1323,In_1789,In_1712);
nor U1324 (N_1324,In_420,In_406);
nor U1325 (N_1325,In_1441,In_831);
nand U1326 (N_1326,In_544,In_1539);
or U1327 (N_1327,In_1549,In_1342);
and U1328 (N_1328,In_1981,In_1548);
and U1329 (N_1329,In_1973,In_2390);
nand U1330 (N_1330,In_1960,In_2469);
or U1331 (N_1331,In_432,In_1978);
nand U1332 (N_1332,In_743,In_1640);
or U1333 (N_1333,In_241,In_1515);
nor U1334 (N_1334,In_1376,In_215);
or U1335 (N_1335,In_2308,In_2312);
nor U1336 (N_1336,In_1825,In_1547);
nand U1337 (N_1337,In_1637,In_2184);
nand U1338 (N_1338,In_1870,In_2173);
xnor U1339 (N_1339,In_2223,In_762);
xnor U1340 (N_1340,In_1893,In_1507);
nor U1341 (N_1341,In_1071,In_1769);
or U1342 (N_1342,In_2151,In_2432);
nor U1343 (N_1343,In_254,In_2087);
and U1344 (N_1344,In_2312,In_310);
nor U1345 (N_1345,In_2053,In_1569);
or U1346 (N_1346,In_1453,In_1426);
and U1347 (N_1347,In_1655,In_376);
nand U1348 (N_1348,In_132,In_2457);
xnor U1349 (N_1349,In_1966,In_1546);
and U1350 (N_1350,In_1175,In_1917);
and U1351 (N_1351,In_2451,In_364);
or U1352 (N_1352,In_2440,In_1983);
nand U1353 (N_1353,In_1425,In_1210);
nand U1354 (N_1354,In_167,In_663);
or U1355 (N_1355,In_1929,In_343);
and U1356 (N_1356,In_1063,In_893);
nand U1357 (N_1357,In_1961,In_31);
and U1358 (N_1358,In_1991,In_2324);
or U1359 (N_1359,In_1769,In_2377);
nor U1360 (N_1360,In_2023,In_623);
and U1361 (N_1361,In_2305,In_1030);
nor U1362 (N_1362,In_2261,In_278);
and U1363 (N_1363,In_1923,In_1241);
xor U1364 (N_1364,In_45,In_2490);
nand U1365 (N_1365,In_2276,In_189);
or U1366 (N_1366,In_674,In_416);
and U1367 (N_1367,In_463,In_1082);
and U1368 (N_1368,In_740,In_2097);
nor U1369 (N_1369,In_1591,In_1164);
xnor U1370 (N_1370,In_36,In_446);
nand U1371 (N_1371,In_580,In_3);
nand U1372 (N_1372,In_1028,In_2218);
nor U1373 (N_1373,In_2460,In_1135);
or U1374 (N_1374,In_1885,In_1215);
xnor U1375 (N_1375,In_2092,In_1324);
nand U1376 (N_1376,In_468,In_146);
and U1377 (N_1377,In_1997,In_144);
nand U1378 (N_1378,In_814,In_221);
and U1379 (N_1379,In_1276,In_89);
xor U1380 (N_1380,In_2181,In_1595);
nand U1381 (N_1381,In_1632,In_467);
xor U1382 (N_1382,In_1361,In_565);
nand U1383 (N_1383,In_650,In_2119);
nor U1384 (N_1384,In_758,In_1143);
or U1385 (N_1385,In_1724,In_883);
nand U1386 (N_1386,In_1450,In_521);
or U1387 (N_1387,In_2310,In_1628);
xnor U1388 (N_1388,In_418,In_1721);
and U1389 (N_1389,In_2037,In_2085);
and U1390 (N_1390,In_134,In_939);
nor U1391 (N_1391,In_638,In_942);
and U1392 (N_1392,In_2329,In_387);
nand U1393 (N_1393,In_1668,In_1796);
or U1394 (N_1394,In_2084,In_873);
nor U1395 (N_1395,In_1336,In_1453);
nand U1396 (N_1396,In_166,In_1236);
xor U1397 (N_1397,In_1793,In_513);
nand U1398 (N_1398,In_509,In_2279);
and U1399 (N_1399,In_2070,In_1667);
or U1400 (N_1400,In_1498,In_283);
nand U1401 (N_1401,In_1710,In_1711);
nand U1402 (N_1402,In_356,In_1566);
or U1403 (N_1403,In_913,In_200);
nor U1404 (N_1404,In_667,In_150);
nand U1405 (N_1405,In_212,In_1293);
or U1406 (N_1406,In_2196,In_323);
and U1407 (N_1407,In_316,In_2419);
or U1408 (N_1408,In_830,In_643);
or U1409 (N_1409,In_120,In_2290);
nor U1410 (N_1410,In_1284,In_1154);
xor U1411 (N_1411,In_1080,In_2183);
nand U1412 (N_1412,In_196,In_843);
nor U1413 (N_1413,In_1066,In_344);
nor U1414 (N_1414,In_1904,In_385);
nor U1415 (N_1415,In_1723,In_2022);
and U1416 (N_1416,In_1896,In_1956);
nand U1417 (N_1417,In_1816,In_1406);
nor U1418 (N_1418,In_1728,In_622);
or U1419 (N_1419,In_283,In_1050);
nand U1420 (N_1420,In_2289,In_945);
or U1421 (N_1421,In_2355,In_1171);
nor U1422 (N_1422,In_325,In_202);
nand U1423 (N_1423,In_2310,In_1423);
or U1424 (N_1424,In_192,In_1330);
nand U1425 (N_1425,In_2352,In_708);
nor U1426 (N_1426,In_367,In_1916);
nor U1427 (N_1427,In_107,In_711);
nor U1428 (N_1428,In_2101,In_316);
and U1429 (N_1429,In_1405,In_2429);
and U1430 (N_1430,In_789,In_2249);
and U1431 (N_1431,In_325,In_1901);
nor U1432 (N_1432,In_1977,In_1322);
xnor U1433 (N_1433,In_2280,In_1291);
and U1434 (N_1434,In_2399,In_712);
or U1435 (N_1435,In_866,In_1623);
or U1436 (N_1436,In_444,In_1238);
and U1437 (N_1437,In_643,In_1831);
xnor U1438 (N_1438,In_801,In_1890);
nor U1439 (N_1439,In_531,In_1212);
nor U1440 (N_1440,In_415,In_1700);
nor U1441 (N_1441,In_1178,In_2223);
and U1442 (N_1442,In_532,In_1123);
nor U1443 (N_1443,In_58,In_1263);
nor U1444 (N_1444,In_697,In_624);
nor U1445 (N_1445,In_872,In_389);
xor U1446 (N_1446,In_780,In_2443);
and U1447 (N_1447,In_704,In_1368);
nand U1448 (N_1448,In_1315,In_369);
nand U1449 (N_1449,In_194,In_1916);
xnor U1450 (N_1450,In_2343,In_1909);
or U1451 (N_1451,In_6,In_930);
or U1452 (N_1452,In_184,In_1232);
or U1453 (N_1453,In_761,In_1169);
and U1454 (N_1454,In_1908,In_1364);
and U1455 (N_1455,In_1642,In_2499);
nor U1456 (N_1456,In_1969,In_1453);
and U1457 (N_1457,In_1557,In_1324);
nor U1458 (N_1458,In_79,In_1940);
and U1459 (N_1459,In_2167,In_869);
nor U1460 (N_1460,In_1898,In_2158);
and U1461 (N_1461,In_1674,In_2357);
xor U1462 (N_1462,In_1665,In_577);
and U1463 (N_1463,In_969,In_1387);
nor U1464 (N_1464,In_499,In_1113);
xor U1465 (N_1465,In_503,In_2310);
nand U1466 (N_1466,In_1374,In_525);
nor U1467 (N_1467,In_2430,In_984);
or U1468 (N_1468,In_2068,In_2299);
nor U1469 (N_1469,In_2345,In_229);
or U1470 (N_1470,In_465,In_239);
nor U1471 (N_1471,In_262,In_1575);
nor U1472 (N_1472,In_558,In_2445);
nor U1473 (N_1473,In_2073,In_788);
xor U1474 (N_1474,In_1816,In_2351);
xnor U1475 (N_1475,In_1645,In_2130);
xnor U1476 (N_1476,In_2,In_2370);
or U1477 (N_1477,In_844,In_578);
nor U1478 (N_1478,In_2197,In_419);
nand U1479 (N_1479,In_69,In_2139);
or U1480 (N_1480,In_839,In_1935);
or U1481 (N_1481,In_1538,In_716);
nand U1482 (N_1482,In_1299,In_2318);
nor U1483 (N_1483,In_166,In_326);
or U1484 (N_1484,In_2056,In_450);
and U1485 (N_1485,In_223,In_134);
and U1486 (N_1486,In_442,In_974);
and U1487 (N_1487,In_2046,In_1176);
nand U1488 (N_1488,In_2264,In_2051);
and U1489 (N_1489,In_499,In_142);
nand U1490 (N_1490,In_2186,In_2192);
nor U1491 (N_1491,In_2185,In_2333);
and U1492 (N_1492,In_1423,In_2166);
or U1493 (N_1493,In_2316,In_1739);
and U1494 (N_1494,In_997,In_450);
nor U1495 (N_1495,In_1144,In_627);
nor U1496 (N_1496,In_1482,In_219);
and U1497 (N_1497,In_2442,In_2050);
xor U1498 (N_1498,In_557,In_881);
nand U1499 (N_1499,In_848,In_1232);
or U1500 (N_1500,In_1666,In_108);
nand U1501 (N_1501,In_2134,In_1986);
nand U1502 (N_1502,In_104,In_73);
or U1503 (N_1503,In_943,In_2342);
nor U1504 (N_1504,In_176,In_1175);
nor U1505 (N_1505,In_70,In_1448);
nand U1506 (N_1506,In_2354,In_1015);
and U1507 (N_1507,In_1271,In_324);
nor U1508 (N_1508,In_2246,In_1732);
xor U1509 (N_1509,In_2227,In_2149);
nand U1510 (N_1510,In_2345,In_1783);
or U1511 (N_1511,In_490,In_863);
and U1512 (N_1512,In_2401,In_1127);
xnor U1513 (N_1513,In_623,In_1398);
xnor U1514 (N_1514,In_1372,In_877);
nor U1515 (N_1515,In_413,In_472);
nor U1516 (N_1516,In_419,In_873);
nor U1517 (N_1517,In_206,In_1234);
xor U1518 (N_1518,In_2179,In_1875);
nor U1519 (N_1519,In_931,In_157);
nor U1520 (N_1520,In_750,In_1848);
or U1521 (N_1521,In_1428,In_1630);
nand U1522 (N_1522,In_1385,In_1899);
and U1523 (N_1523,In_1969,In_1637);
and U1524 (N_1524,In_2100,In_1011);
nor U1525 (N_1525,In_1586,In_952);
nand U1526 (N_1526,In_1826,In_1092);
and U1527 (N_1527,In_1796,In_1794);
nand U1528 (N_1528,In_395,In_1023);
and U1529 (N_1529,In_1494,In_2330);
nor U1530 (N_1530,In_2220,In_1421);
nor U1531 (N_1531,In_632,In_703);
and U1532 (N_1532,In_193,In_65);
and U1533 (N_1533,In_2400,In_365);
and U1534 (N_1534,In_435,In_502);
nor U1535 (N_1535,In_975,In_1250);
nor U1536 (N_1536,In_2270,In_1311);
or U1537 (N_1537,In_499,In_2016);
and U1538 (N_1538,In_1824,In_369);
or U1539 (N_1539,In_767,In_956);
nor U1540 (N_1540,In_2040,In_1305);
and U1541 (N_1541,In_2409,In_701);
or U1542 (N_1542,In_1043,In_1126);
nand U1543 (N_1543,In_729,In_1131);
and U1544 (N_1544,In_1446,In_1917);
nor U1545 (N_1545,In_717,In_2213);
nor U1546 (N_1546,In_2008,In_1620);
and U1547 (N_1547,In_1224,In_1927);
or U1548 (N_1548,In_898,In_1873);
nand U1549 (N_1549,In_1387,In_1659);
and U1550 (N_1550,In_119,In_1531);
nand U1551 (N_1551,In_711,In_1434);
nand U1552 (N_1552,In_41,In_27);
nor U1553 (N_1553,In_1849,In_1728);
and U1554 (N_1554,In_1456,In_1123);
or U1555 (N_1555,In_2233,In_681);
or U1556 (N_1556,In_2013,In_1728);
or U1557 (N_1557,In_559,In_1622);
and U1558 (N_1558,In_1879,In_50);
or U1559 (N_1559,In_33,In_2184);
nor U1560 (N_1560,In_1392,In_293);
nand U1561 (N_1561,In_642,In_1248);
xnor U1562 (N_1562,In_1609,In_1580);
nor U1563 (N_1563,In_291,In_1067);
nand U1564 (N_1564,In_549,In_194);
and U1565 (N_1565,In_1887,In_2290);
or U1566 (N_1566,In_411,In_1909);
and U1567 (N_1567,In_1665,In_1322);
or U1568 (N_1568,In_167,In_972);
and U1569 (N_1569,In_931,In_1705);
or U1570 (N_1570,In_1241,In_1340);
nor U1571 (N_1571,In_1003,In_364);
nor U1572 (N_1572,In_673,In_2119);
nor U1573 (N_1573,In_838,In_1021);
nor U1574 (N_1574,In_56,In_1175);
or U1575 (N_1575,In_864,In_295);
or U1576 (N_1576,In_905,In_2201);
nor U1577 (N_1577,In_1273,In_2370);
nand U1578 (N_1578,In_488,In_2420);
nand U1579 (N_1579,In_0,In_1355);
and U1580 (N_1580,In_250,In_72);
and U1581 (N_1581,In_530,In_1465);
nand U1582 (N_1582,In_302,In_243);
and U1583 (N_1583,In_310,In_2166);
nor U1584 (N_1584,In_1406,In_1456);
nand U1585 (N_1585,In_2020,In_1319);
nor U1586 (N_1586,In_17,In_1393);
nor U1587 (N_1587,In_390,In_1279);
and U1588 (N_1588,In_76,In_2327);
and U1589 (N_1589,In_1980,In_1547);
nand U1590 (N_1590,In_1248,In_1798);
nand U1591 (N_1591,In_196,In_2221);
and U1592 (N_1592,In_34,In_2045);
nand U1593 (N_1593,In_1751,In_1634);
nand U1594 (N_1594,In_231,In_315);
and U1595 (N_1595,In_1991,In_927);
and U1596 (N_1596,In_2491,In_1625);
or U1597 (N_1597,In_1721,In_527);
and U1598 (N_1598,In_1750,In_645);
nand U1599 (N_1599,In_410,In_1666);
or U1600 (N_1600,In_1414,In_2103);
and U1601 (N_1601,In_970,In_2188);
xor U1602 (N_1602,In_1477,In_220);
nor U1603 (N_1603,In_2321,In_320);
or U1604 (N_1604,In_1908,In_379);
nor U1605 (N_1605,In_564,In_576);
and U1606 (N_1606,In_1507,In_1610);
and U1607 (N_1607,In_2399,In_342);
nand U1608 (N_1608,In_228,In_939);
or U1609 (N_1609,In_502,In_1859);
or U1610 (N_1610,In_1311,In_158);
xnor U1611 (N_1611,In_1606,In_1161);
or U1612 (N_1612,In_1784,In_1001);
nor U1613 (N_1613,In_2407,In_1662);
or U1614 (N_1614,In_864,In_980);
nand U1615 (N_1615,In_314,In_1590);
and U1616 (N_1616,In_1495,In_2268);
nand U1617 (N_1617,In_2345,In_965);
xnor U1618 (N_1618,In_816,In_1502);
xnor U1619 (N_1619,In_423,In_2419);
or U1620 (N_1620,In_2256,In_2461);
nor U1621 (N_1621,In_281,In_1329);
or U1622 (N_1622,In_1975,In_1021);
and U1623 (N_1623,In_1114,In_2219);
nor U1624 (N_1624,In_190,In_708);
nor U1625 (N_1625,In_1820,In_2436);
nand U1626 (N_1626,In_1842,In_1856);
nand U1627 (N_1627,In_911,In_2132);
xor U1628 (N_1628,In_525,In_1160);
and U1629 (N_1629,In_582,In_1864);
xnor U1630 (N_1630,In_304,In_230);
nor U1631 (N_1631,In_203,In_1882);
or U1632 (N_1632,In_951,In_755);
nor U1633 (N_1633,In_1388,In_780);
and U1634 (N_1634,In_927,In_1973);
xnor U1635 (N_1635,In_1785,In_1890);
or U1636 (N_1636,In_903,In_454);
and U1637 (N_1637,In_2196,In_482);
or U1638 (N_1638,In_1690,In_2229);
xnor U1639 (N_1639,In_871,In_864);
and U1640 (N_1640,In_1504,In_2065);
or U1641 (N_1641,In_148,In_2226);
xor U1642 (N_1642,In_242,In_406);
nor U1643 (N_1643,In_1406,In_2484);
or U1644 (N_1644,In_1182,In_257);
and U1645 (N_1645,In_913,In_2177);
or U1646 (N_1646,In_1479,In_1528);
nor U1647 (N_1647,In_1541,In_580);
nand U1648 (N_1648,In_1813,In_828);
xor U1649 (N_1649,In_603,In_1115);
and U1650 (N_1650,In_1632,In_1548);
nand U1651 (N_1651,In_35,In_2049);
and U1652 (N_1652,In_1109,In_1954);
nor U1653 (N_1653,In_1716,In_2328);
nand U1654 (N_1654,In_1457,In_2);
or U1655 (N_1655,In_136,In_913);
nor U1656 (N_1656,In_51,In_1615);
xor U1657 (N_1657,In_508,In_1217);
nand U1658 (N_1658,In_2119,In_2299);
or U1659 (N_1659,In_1080,In_793);
and U1660 (N_1660,In_588,In_1777);
nor U1661 (N_1661,In_91,In_1282);
xnor U1662 (N_1662,In_1648,In_1774);
or U1663 (N_1663,In_2243,In_2115);
nand U1664 (N_1664,In_1797,In_746);
nor U1665 (N_1665,In_601,In_1979);
or U1666 (N_1666,In_1124,In_2378);
xnor U1667 (N_1667,In_640,In_233);
or U1668 (N_1668,In_373,In_1109);
xnor U1669 (N_1669,In_973,In_1665);
or U1670 (N_1670,In_2121,In_1117);
and U1671 (N_1671,In_1914,In_2469);
or U1672 (N_1672,In_2403,In_2282);
nand U1673 (N_1673,In_2389,In_1792);
xnor U1674 (N_1674,In_203,In_1070);
and U1675 (N_1675,In_2329,In_2456);
nor U1676 (N_1676,In_419,In_740);
xor U1677 (N_1677,In_1256,In_530);
nand U1678 (N_1678,In_661,In_589);
xor U1679 (N_1679,In_2495,In_859);
and U1680 (N_1680,In_1898,In_1053);
xor U1681 (N_1681,In_1793,In_473);
or U1682 (N_1682,In_2245,In_1098);
and U1683 (N_1683,In_511,In_1343);
and U1684 (N_1684,In_1222,In_1823);
nand U1685 (N_1685,In_157,In_476);
nor U1686 (N_1686,In_2000,In_1735);
xnor U1687 (N_1687,In_1391,In_1916);
nor U1688 (N_1688,In_179,In_645);
nor U1689 (N_1689,In_2141,In_67);
nand U1690 (N_1690,In_186,In_2193);
xnor U1691 (N_1691,In_542,In_999);
or U1692 (N_1692,In_1398,In_650);
and U1693 (N_1693,In_266,In_507);
and U1694 (N_1694,In_1670,In_338);
and U1695 (N_1695,In_2005,In_1899);
and U1696 (N_1696,In_2272,In_313);
nand U1697 (N_1697,In_2450,In_657);
xor U1698 (N_1698,In_1167,In_1969);
nand U1699 (N_1699,In_665,In_658);
and U1700 (N_1700,In_1288,In_134);
and U1701 (N_1701,In_1711,In_1896);
and U1702 (N_1702,In_350,In_1084);
nand U1703 (N_1703,In_565,In_845);
nor U1704 (N_1704,In_1132,In_2187);
nand U1705 (N_1705,In_975,In_1784);
and U1706 (N_1706,In_30,In_2417);
xor U1707 (N_1707,In_717,In_1574);
nand U1708 (N_1708,In_586,In_1279);
xnor U1709 (N_1709,In_1233,In_2069);
and U1710 (N_1710,In_2498,In_582);
nor U1711 (N_1711,In_7,In_347);
and U1712 (N_1712,In_693,In_541);
and U1713 (N_1713,In_2236,In_1809);
nand U1714 (N_1714,In_70,In_1372);
and U1715 (N_1715,In_819,In_449);
nand U1716 (N_1716,In_328,In_976);
nand U1717 (N_1717,In_2326,In_1766);
nor U1718 (N_1718,In_1815,In_2289);
nand U1719 (N_1719,In_757,In_1791);
nand U1720 (N_1720,In_471,In_1413);
or U1721 (N_1721,In_1331,In_1382);
and U1722 (N_1722,In_2454,In_188);
nor U1723 (N_1723,In_607,In_1595);
nand U1724 (N_1724,In_2102,In_2239);
and U1725 (N_1725,In_1720,In_824);
nor U1726 (N_1726,In_2443,In_241);
nor U1727 (N_1727,In_171,In_2375);
and U1728 (N_1728,In_2147,In_1913);
xor U1729 (N_1729,In_276,In_2);
or U1730 (N_1730,In_726,In_147);
nor U1731 (N_1731,In_1425,In_2367);
nor U1732 (N_1732,In_2267,In_922);
nand U1733 (N_1733,In_2381,In_1931);
or U1734 (N_1734,In_2407,In_1882);
nand U1735 (N_1735,In_2173,In_1990);
or U1736 (N_1736,In_2146,In_2329);
nor U1737 (N_1737,In_1257,In_571);
nand U1738 (N_1738,In_2413,In_3);
xor U1739 (N_1739,In_510,In_901);
or U1740 (N_1740,In_452,In_1374);
and U1741 (N_1741,In_1788,In_1785);
nor U1742 (N_1742,In_1659,In_1398);
xor U1743 (N_1743,In_432,In_39);
or U1744 (N_1744,In_395,In_1017);
nand U1745 (N_1745,In_9,In_732);
or U1746 (N_1746,In_189,In_1982);
nand U1747 (N_1747,In_1385,In_495);
xnor U1748 (N_1748,In_1349,In_1274);
nand U1749 (N_1749,In_2462,In_1362);
nand U1750 (N_1750,In_644,In_2303);
and U1751 (N_1751,In_336,In_473);
nor U1752 (N_1752,In_2351,In_2210);
or U1753 (N_1753,In_1070,In_1914);
nor U1754 (N_1754,In_2485,In_1736);
nor U1755 (N_1755,In_1475,In_1592);
and U1756 (N_1756,In_2146,In_412);
nor U1757 (N_1757,In_1918,In_1932);
nor U1758 (N_1758,In_32,In_262);
nand U1759 (N_1759,In_1224,In_1960);
xor U1760 (N_1760,In_1430,In_360);
and U1761 (N_1761,In_2027,In_1004);
xnor U1762 (N_1762,In_449,In_995);
nand U1763 (N_1763,In_237,In_443);
nor U1764 (N_1764,In_872,In_2320);
or U1765 (N_1765,In_1872,In_1963);
or U1766 (N_1766,In_1620,In_87);
or U1767 (N_1767,In_728,In_1400);
or U1768 (N_1768,In_324,In_430);
nor U1769 (N_1769,In_2258,In_1963);
nor U1770 (N_1770,In_2435,In_416);
nor U1771 (N_1771,In_1774,In_764);
and U1772 (N_1772,In_767,In_1122);
nand U1773 (N_1773,In_581,In_1131);
and U1774 (N_1774,In_1439,In_1788);
or U1775 (N_1775,In_47,In_372);
xor U1776 (N_1776,In_1933,In_973);
nor U1777 (N_1777,In_1698,In_2387);
xor U1778 (N_1778,In_300,In_1562);
xnor U1779 (N_1779,In_343,In_1781);
or U1780 (N_1780,In_912,In_224);
or U1781 (N_1781,In_1043,In_388);
nand U1782 (N_1782,In_1809,In_1060);
nor U1783 (N_1783,In_987,In_518);
or U1784 (N_1784,In_801,In_334);
nor U1785 (N_1785,In_1624,In_2167);
and U1786 (N_1786,In_1913,In_2276);
nor U1787 (N_1787,In_540,In_2130);
and U1788 (N_1788,In_1938,In_2497);
and U1789 (N_1789,In_1347,In_1556);
or U1790 (N_1790,In_1668,In_652);
nand U1791 (N_1791,In_2368,In_1062);
nand U1792 (N_1792,In_1790,In_2492);
xor U1793 (N_1793,In_2168,In_2274);
nor U1794 (N_1794,In_2369,In_223);
nand U1795 (N_1795,In_659,In_1963);
nand U1796 (N_1796,In_465,In_1369);
or U1797 (N_1797,In_395,In_98);
and U1798 (N_1798,In_1293,In_173);
and U1799 (N_1799,In_1882,In_1593);
or U1800 (N_1800,In_345,In_2053);
or U1801 (N_1801,In_2251,In_974);
and U1802 (N_1802,In_61,In_953);
nand U1803 (N_1803,In_2402,In_1056);
xnor U1804 (N_1804,In_1702,In_2429);
nor U1805 (N_1805,In_1866,In_2293);
or U1806 (N_1806,In_2284,In_1686);
and U1807 (N_1807,In_667,In_665);
nand U1808 (N_1808,In_708,In_2239);
and U1809 (N_1809,In_2054,In_37);
and U1810 (N_1810,In_1080,In_131);
nand U1811 (N_1811,In_426,In_34);
or U1812 (N_1812,In_876,In_1245);
and U1813 (N_1813,In_962,In_37);
and U1814 (N_1814,In_1124,In_2045);
and U1815 (N_1815,In_2024,In_874);
or U1816 (N_1816,In_91,In_11);
or U1817 (N_1817,In_1271,In_1363);
nand U1818 (N_1818,In_449,In_740);
nor U1819 (N_1819,In_76,In_2310);
nand U1820 (N_1820,In_1429,In_675);
or U1821 (N_1821,In_998,In_1388);
or U1822 (N_1822,In_239,In_2381);
and U1823 (N_1823,In_1501,In_2302);
or U1824 (N_1824,In_12,In_805);
and U1825 (N_1825,In_723,In_2377);
nor U1826 (N_1826,In_1364,In_1570);
or U1827 (N_1827,In_1974,In_178);
nor U1828 (N_1828,In_1000,In_661);
nand U1829 (N_1829,In_300,In_671);
and U1830 (N_1830,In_2103,In_29);
nor U1831 (N_1831,In_1540,In_1947);
nand U1832 (N_1832,In_1167,In_2333);
nor U1833 (N_1833,In_1227,In_508);
or U1834 (N_1834,In_2285,In_439);
and U1835 (N_1835,In_1284,In_453);
and U1836 (N_1836,In_177,In_1179);
and U1837 (N_1837,In_1194,In_807);
nand U1838 (N_1838,In_729,In_85);
or U1839 (N_1839,In_1314,In_1141);
nand U1840 (N_1840,In_332,In_2091);
nor U1841 (N_1841,In_1902,In_2170);
and U1842 (N_1842,In_476,In_2434);
nand U1843 (N_1843,In_398,In_72);
or U1844 (N_1844,In_1149,In_570);
or U1845 (N_1845,In_1889,In_860);
and U1846 (N_1846,In_1815,In_286);
nand U1847 (N_1847,In_2006,In_764);
nor U1848 (N_1848,In_1379,In_547);
and U1849 (N_1849,In_1306,In_2357);
nor U1850 (N_1850,In_1995,In_938);
nor U1851 (N_1851,In_394,In_393);
or U1852 (N_1852,In_1829,In_92);
and U1853 (N_1853,In_27,In_2221);
and U1854 (N_1854,In_90,In_103);
or U1855 (N_1855,In_91,In_1356);
and U1856 (N_1856,In_1994,In_1145);
and U1857 (N_1857,In_543,In_2262);
and U1858 (N_1858,In_525,In_96);
nor U1859 (N_1859,In_306,In_172);
and U1860 (N_1860,In_1400,In_2246);
and U1861 (N_1861,In_613,In_1410);
nand U1862 (N_1862,In_1619,In_1779);
nor U1863 (N_1863,In_95,In_1845);
and U1864 (N_1864,In_1580,In_442);
and U1865 (N_1865,In_1107,In_1425);
nand U1866 (N_1866,In_858,In_2157);
xnor U1867 (N_1867,In_1713,In_1679);
nor U1868 (N_1868,In_1692,In_2454);
nor U1869 (N_1869,In_342,In_1043);
and U1870 (N_1870,In_1839,In_1371);
nand U1871 (N_1871,In_1946,In_752);
and U1872 (N_1872,In_2025,In_1008);
and U1873 (N_1873,In_2130,In_1099);
or U1874 (N_1874,In_914,In_357);
or U1875 (N_1875,In_545,In_2191);
nor U1876 (N_1876,In_767,In_2208);
and U1877 (N_1877,In_1584,In_1399);
or U1878 (N_1878,In_1131,In_1129);
or U1879 (N_1879,In_1053,In_1740);
or U1880 (N_1880,In_2235,In_192);
xnor U1881 (N_1881,In_1615,In_934);
or U1882 (N_1882,In_1601,In_2440);
nand U1883 (N_1883,In_438,In_837);
nand U1884 (N_1884,In_536,In_1663);
nor U1885 (N_1885,In_237,In_1616);
or U1886 (N_1886,In_1206,In_393);
nor U1887 (N_1887,In_892,In_531);
nor U1888 (N_1888,In_1635,In_981);
or U1889 (N_1889,In_857,In_1155);
and U1890 (N_1890,In_911,In_1021);
nand U1891 (N_1891,In_346,In_1421);
nand U1892 (N_1892,In_819,In_1607);
nor U1893 (N_1893,In_156,In_53);
and U1894 (N_1894,In_894,In_1242);
and U1895 (N_1895,In_1421,In_769);
xnor U1896 (N_1896,In_305,In_2293);
and U1897 (N_1897,In_2241,In_2351);
or U1898 (N_1898,In_441,In_1355);
and U1899 (N_1899,In_904,In_2119);
and U1900 (N_1900,In_357,In_1123);
or U1901 (N_1901,In_1364,In_373);
xor U1902 (N_1902,In_925,In_1951);
and U1903 (N_1903,In_268,In_66);
nor U1904 (N_1904,In_1013,In_2395);
xor U1905 (N_1905,In_1317,In_1525);
and U1906 (N_1906,In_131,In_904);
nor U1907 (N_1907,In_1094,In_1173);
or U1908 (N_1908,In_868,In_2158);
and U1909 (N_1909,In_703,In_675);
nor U1910 (N_1910,In_1378,In_372);
or U1911 (N_1911,In_1581,In_1057);
nand U1912 (N_1912,In_2333,In_1233);
nand U1913 (N_1913,In_2012,In_2033);
or U1914 (N_1914,In_6,In_2215);
nor U1915 (N_1915,In_1374,In_57);
xor U1916 (N_1916,In_1090,In_38);
or U1917 (N_1917,In_1447,In_2334);
or U1918 (N_1918,In_254,In_1916);
nor U1919 (N_1919,In_1959,In_762);
xor U1920 (N_1920,In_1075,In_852);
and U1921 (N_1921,In_2358,In_1672);
nand U1922 (N_1922,In_1888,In_766);
xnor U1923 (N_1923,In_2377,In_1103);
or U1924 (N_1924,In_2311,In_1434);
nor U1925 (N_1925,In_1185,In_2057);
xnor U1926 (N_1926,In_336,In_144);
or U1927 (N_1927,In_1633,In_275);
nand U1928 (N_1928,In_174,In_1872);
or U1929 (N_1929,In_1269,In_1423);
or U1930 (N_1930,In_1398,In_189);
and U1931 (N_1931,In_2248,In_295);
nand U1932 (N_1932,In_1354,In_708);
and U1933 (N_1933,In_2318,In_1191);
and U1934 (N_1934,In_2081,In_425);
or U1935 (N_1935,In_2119,In_2098);
nor U1936 (N_1936,In_1680,In_1616);
and U1937 (N_1937,In_2038,In_1907);
and U1938 (N_1938,In_1387,In_968);
nand U1939 (N_1939,In_479,In_1410);
nand U1940 (N_1940,In_2264,In_1937);
nor U1941 (N_1941,In_2333,In_1936);
xnor U1942 (N_1942,In_1717,In_2417);
and U1943 (N_1943,In_2032,In_207);
nand U1944 (N_1944,In_349,In_616);
or U1945 (N_1945,In_899,In_1148);
or U1946 (N_1946,In_65,In_316);
and U1947 (N_1947,In_154,In_533);
nand U1948 (N_1948,In_996,In_1407);
and U1949 (N_1949,In_2030,In_753);
nor U1950 (N_1950,In_1778,In_1556);
and U1951 (N_1951,In_1746,In_2309);
and U1952 (N_1952,In_2024,In_662);
or U1953 (N_1953,In_1198,In_1782);
nor U1954 (N_1954,In_2192,In_38);
xnor U1955 (N_1955,In_697,In_1688);
nand U1956 (N_1956,In_390,In_239);
or U1957 (N_1957,In_2201,In_47);
nor U1958 (N_1958,In_687,In_1818);
and U1959 (N_1959,In_59,In_1767);
or U1960 (N_1960,In_1104,In_806);
and U1961 (N_1961,In_560,In_2494);
or U1962 (N_1962,In_1193,In_70);
nand U1963 (N_1963,In_376,In_2);
xnor U1964 (N_1964,In_1000,In_1095);
nand U1965 (N_1965,In_2155,In_2048);
xor U1966 (N_1966,In_1632,In_1649);
or U1967 (N_1967,In_1914,In_560);
and U1968 (N_1968,In_2003,In_1238);
nor U1969 (N_1969,In_1312,In_1377);
nand U1970 (N_1970,In_807,In_325);
nand U1971 (N_1971,In_2456,In_1973);
nor U1972 (N_1972,In_273,In_870);
and U1973 (N_1973,In_2475,In_1188);
or U1974 (N_1974,In_383,In_412);
nand U1975 (N_1975,In_69,In_1700);
nor U1976 (N_1976,In_2112,In_501);
or U1977 (N_1977,In_1486,In_762);
or U1978 (N_1978,In_1238,In_2192);
nor U1979 (N_1979,In_346,In_1610);
or U1980 (N_1980,In_1616,In_660);
nor U1981 (N_1981,In_2361,In_486);
nand U1982 (N_1982,In_1455,In_198);
nor U1983 (N_1983,In_1381,In_1235);
or U1984 (N_1984,In_956,In_774);
or U1985 (N_1985,In_2252,In_1796);
or U1986 (N_1986,In_2008,In_1297);
or U1987 (N_1987,In_1860,In_2117);
and U1988 (N_1988,In_518,In_1263);
nand U1989 (N_1989,In_1427,In_2002);
nor U1990 (N_1990,In_282,In_1197);
nor U1991 (N_1991,In_3,In_2157);
or U1992 (N_1992,In_1437,In_922);
nand U1993 (N_1993,In_185,In_873);
nand U1994 (N_1994,In_1931,In_578);
nand U1995 (N_1995,In_1242,In_513);
or U1996 (N_1996,In_1257,In_316);
nor U1997 (N_1997,In_1549,In_121);
nor U1998 (N_1998,In_578,In_1000);
nor U1999 (N_1999,In_1563,In_1878);
nor U2000 (N_2000,In_465,In_1834);
nor U2001 (N_2001,In_734,In_44);
or U2002 (N_2002,In_1316,In_2212);
and U2003 (N_2003,In_396,In_1279);
nor U2004 (N_2004,In_692,In_1513);
xor U2005 (N_2005,In_9,In_1684);
and U2006 (N_2006,In_2267,In_353);
or U2007 (N_2007,In_654,In_7);
and U2008 (N_2008,In_1368,In_1385);
nor U2009 (N_2009,In_1161,In_537);
nand U2010 (N_2010,In_1373,In_2049);
nor U2011 (N_2011,In_2449,In_863);
nand U2012 (N_2012,In_223,In_20);
and U2013 (N_2013,In_2430,In_2086);
or U2014 (N_2014,In_1606,In_1277);
nor U2015 (N_2015,In_1630,In_1672);
and U2016 (N_2016,In_1466,In_144);
and U2017 (N_2017,In_2087,In_2129);
nor U2018 (N_2018,In_503,In_499);
nor U2019 (N_2019,In_998,In_1376);
or U2020 (N_2020,In_971,In_130);
and U2021 (N_2021,In_126,In_1396);
nor U2022 (N_2022,In_1525,In_325);
xor U2023 (N_2023,In_2262,In_1868);
and U2024 (N_2024,In_982,In_482);
and U2025 (N_2025,In_1043,In_2424);
and U2026 (N_2026,In_2309,In_2122);
nor U2027 (N_2027,In_995,In_1896);
nor U2028 (N_2028,In_1796,In_432);
nor U2029 (N_2029,In_499,In_1987);
and U2030 (N_2030,In_645,In_1098);
nand U2031 (N_2031,In_1929,In_375);
and U2032 (N_2032,In_634,In_762);
and U2033 (N_2033,In_698,In_1282);
nand U2034 (N_2034,In_2411,In_500);
nor U2035 (N_2035,In_1239,In_1575);
nand U2036 (N_2036,In_2113,In_2161);
and U2037 (N_2037,In_583,In_66);
xnor U2038 (N_2038,In_148,In_1748);
and U2039 (N_2039,In_2413,In_941);
or U2040 (N_2040,In_1435,In_440);
xor U2041 (N_2041,In_1454,In_2420);
or U2042 (N_2042,In_1544,In_1960);
nand U2043 (N_2043,In_1162,In_1701);
and U2044 (N_2044,In_923,In_147);
nor U2045 (N_2045,In_2274,In_2019);
nor U2046 (N_2046,In_736,In_1586);
nor U2047 (N_2047,In_428,In_789);
nand U2048 (N_2048,In_531,In_1912);
nor U2049 (N_2049,In_2180,In_402);
or U2050 (N_2050,In_531,In_169);
and U2051 (N_2051,In_647,In_2126);
xnor U2052 (N_2052,In_956,In_313);
nor U2053 (N_2053,In_1366,In_2273);
and U2054 (N_2054,In_761,In_243);
or U2055 (N_2055,In_1953,In_2457);
nor U2056 (N_2056,In_1470,In_288);
nor U2057 (N_2057,In_67,In_108);
nand U2058 (N_2058,In_1045,In_506);
xor U2059 (N_2059,In_1507,In_736);
xor U2060 (N_2060,In_305,In_2419);
nor U2061 (N_2061,In_2459,In_2045);
or U2062 (N_2062,In_2365,In_1909);
or U2063 (N_2063,In_1576,In_2236);
nor U2064 (N_2064,In_669,In_21);
xor U2065 (N_2065,In_282,In_1221);
nand U2066 (N_2066,In_83,In_993);
nor U2067 (N_2067,In_91,In_1655);
and U2068 (N_2068,In_443,In_515);
nor U2069 (N_2069,In_2014,In_766);
or U2070 (N_2070,In_71,In_1764);
nor U2071 (N_2071,In_2258,In_542);
nand U2072 (N_2072,In_239,In_2463);
and U2073 (N_2073,In_2387,In_206);
nor U2074 (N_2074,In_672,In_955);
nor U2075 (N_2075,In_1732,In_512);
nor U2076 (N_2076,In_568,In_2373);
nand U2077 (N_2077,In_1918,In_796);
nand U2078 (N_2078,In_2042,In_1742);
or U2079 (N_2079,In_1295,In_1967);
nand U2080 (N_2080,In_1503,In_1010);
nor U2081 (N_2081,In_1429,In_2382);
nand U2082 (N_2082,In_1983,In_1254);
or U2083 (N_2083,In_1491,In_456);
nand U2084 (N_2084,In_1092,In_1039);
and U2085 (N_2085,In_938,In_2137);
nor U2086 (N_2086,In_230,In_2296);
and U2087 (N_2087,In_150,In_1177);
or U2088 (N_2088,In_2307,In_920);
nor U2089 (N_2089,In_1185,In_1553);
or U2090 (N_2090,In_1865,In_1246);
and U2091 (N_2091,In_1528,In_1121);
nor U2092 (N_2092,In_1062,In_445);
nand U2093 (N_2093,In_1007,In_309);
nand U2094 (N_2094,In_57,In_150);
and U2095 (N_2095,In_999,In_329);
nand U2096 (N_2096,In_1928,In_2417);
nand U2097 (N_2097,In_1727,In_397);
and U2098 (N_2098,In_1119,In_1259);
or U2099 (N_2099,In_1298,In_232);
and U2100 (N_2100,In_2018,In_887);
nand U2101 (N_2101,In_892,In_1267);
or U2102 (N_2102,In_2036,In_1525);
and U2103 (N_2103,In_873,In_620);
and U2104 (N_2104,In_82,In_1090);
nor U2105 (N_2105,In_991,In_476);
nor U2106 (N_2106,In_1282,In_922);
nand U2107 (N_2107,In_2329,In_1121);
nand U2108 (N_2108,In_2278,In_1787);
nor U2109 (N_2109,In_1440,In_743);
and U2110 (N_2110,In_2167,In_2373);
nand U2111 (N_2111,In_1213,In_651);
nor U2112 (N_2112,In_2311,In_1067);
or U2113 (N_2113,In_929,In_1634);
or U2114 (N_2114,In_214,In_2001);
and U2115 (N_2115,In_442,In_765);
xor U2116 (N_2116,In_2406,In_2062);
nand U2117 (N_2117,In_749,In_1002);
nor U2118 (N_2118,In_1815,In_764);
or U2119 (N_2119,In_337,In_1176);
and U2120 (N_2120,In_1022,In_725);
nor U2121 (N_2121,In_1365,In_1036);
nand U2122 (N_2122,In_421,In_2241);
nand U2123 (N_2123,In_1525,In_1152);
or U2124 (N_2124,In_751,In_20);
and U2125 (N_2125,In_2403,In_1520);
nor U2126 (N_2126,In_106,In_757);
nor U2127 (N_2127,In_1522,In_2157);
and U2128 (N_2128,In_2169,In_1533);
or U2129 (N_2129,In_1078,In_1704);
xnor U2130 (N_2130,In_485,In_188);
nand U2131 (N_2131,In_1581,In_2416);
and U2132 (N_2132,In_841,In_2410);
and U2133 (N_2133,In_1304,In_2442);
nor U2134 (N_2134,In_2270,In_2400);
and U2135 (N_2135,In_1616,In_1634);
or U2136 (N_2136,In_8,In_1692);
or U2137 (N_2137,In_1679,In_1467);
nor U2138 (N_2138,In_2250,In_228);
xnor U2139 (N_2139,In_505,In_498);
nand U2140 (N_2140,In_645,In_310);
nor U2141 (N_2141,In_306,In_977);
nand U2142 (N_2142,In_767,In_198);
nand U2143 (N_2143,In_429,In_1404);
nor U2144 (N_2144,In_1988,In_411);
xnor U2145 (N_2145,In_1186,In_1793);
and U2146 (N_2146,In_1522,In_2496);
nand U2147 (N_2147,In_2138,In_743);
and U2148 (N_2148,In_573,In_2393);
or U2149 (N_2149,In_1256,In_16);
nor U2150 (N_2150,In_1720,In_1773);
nand U2151 (N_2151,In_1147,In_1564);
nor U2152 (N_2152,In_1854,In_696);
nor U2153 (N_2153,In_269,In_1483);
nor U2154 (N_2154,In_1650,In_200);
and U2155 (N_2155,In_218,In_2349);
nand U2156 (N_2156,In_1379,In_471);
or U2157 (N_2157,In_2151,In_832);
nand U2158 (N_2158,In_2374,In_1719);
xnor U2159 (N_2159,In_716,In_1238);
nor U2160 (N_2160,In_1158,In_2121);
nor U2161 (N_2161,In_1552,In_2424);
or U2162 (N_2162,In_2203,In_58);
nor U2163 (N_2163,In_1271,In_2281);
nor U2164 (N_2164,In_2189,In_2201);
nand U2165 (N_2165,In_1860,In_1289);
nand U2166 (N_2166,In_1584,In_852);
nand U2167 (N_2167,In_1201,In_643);
nor U2168 (N_2168,In_1557,In_2057);
nor U2169 (N_2169,In_243,In_682);
xor U2170 (N_2170,In_1926,In_2098);
nand U2171 (N_2171,In_335,In_238);
or U2172 (N_2172,In_1182,In_1802);
and U2173 (N_2173,In_128,In_1676);
xor U2174 (N_2174,In_2484,In_1844);
nor U2175 (N_2175,In_1540,In_172);
nor U2176 (N_2176,In_1640,In_1098);
nor U2177 (N_2177,In_243,In_1746);
or U2178 (N_2178,In_822,In_1951);
or U2179 (N_2179,In_2127,In_2224);
and U2180 (N_2180,In_2359,In_783);
and U2181 (N_2181,In_1411,In_1165);
nand U2182 (N_2182,In_188,In_935);
xnor U2183 (N_2183,In_987,In_694);
or U2184 (N_2184,In_1317,In_1709);
nand U2185 (N_2185,In_2231,In_662);
or U2186 (N_2186,In_548,In_1330);
nand U2187 (N_2187,In_609,In_682);
or U2188 (N_2188,In_691,In_2289);
or U2189 (N_2189,In_2036,In_1538);
nor U2190 (N_2190,In_2139,In_744);
nand U2191 (N_2191,In_862,In_315);
nand U2192 (N_2192,In_1817,In_1776);
nor U2193 (N_2193,In_1743,In_1660);
nand U2194 (N_2194,In_717,In_1477);
and U2195 (N_2195,In_1993,In_1721);
nor U2196 (N_2196,In_1744,In_125);
nor U2197 (N_2197,In_2142,In_1125);
nand U2198 (N_2198,In_595,In_1881);
nor U2199 (N_2199,In_1180,In_146);
nand U2200 (N_2200,In_622,In_1415);
nand U2201 (N_2201,In_1716,In_1529);
or U2202 (N_2202,In_1478,In_2028);
nand U2203 (N_2203,In_73,In_920);
and U2204 (N_2204,In_2437,In_1956);
nor U2205 (N_2205,In_435,In_242);
nor U2206 (N_2206,In_1038,In_2099);
nand U2207 (N_2207,In_248,In_908);
nand U2208 (N_2208,In_1235,In_457);
or U2209 (N_2209,In_841,In_791);
or U2210 (N_2210,In_364,In_695);
xnor U2211 (N_2211,In_95,In_1217);
nor U2212 (N_2212,In_1357,In_417);
nand U2213 (N_2213,In_519,In_1596);
and U2214 (N_2214,In_139,In_2192);
and U2215 (N_2215,In_2078,In_1692);
or U2216 (N_2216,In_1137,In_1361);
nor U2217 (N_2217,In_147,In_777);
nor U2218 (N_2218,In_1860,In_1692);
and U2219 (N_2219,In_1779,In_371);
or U2220 (N_2220,In_1301,In_476);
and U2221 (N_2221,In_2391,In_139);
nand U2222 (N_2222,In_1784,In_2026);
and U2223 (N_2223,In_1781,In_348);
and U2224 (N_2224,In_2221,In_2352);
or U2225 (N_2225,In_729,In_740);
xnor U2226 (N_2226,In_722,In_1397);
xnor U2227 (N_2227,In_610,In_531);
nor U2228 (N_2228,In_552,In_976);
xor U2229 (N_2229,In_1721,In_1801);
xnor U2230 (N_2230,In_959,In_986);
nand U2231 (N_2231,In_1827,In_206);
nand U2232 (N_2232,In_2486,In_1302);
or U2233 (N_2233,In_2454,In_965);
nor U2234 (N_2234,In_2140,In_2149);
nor U2235 (N_2235,In_1588,In_1684);
or U2236 (N_2236,In_12,In_1169);
and U2237 (N_2237,In_1245,In_1976);
nor U2238 (N_2238,In_1807,In_1739);
or U2239 (N_2239,In_1565,In_1552);
and U2240 (N_2240,In_1486,In_176);
or U2241 (N_2241,In_1723,In_1773);
xnor U2242 (N_2242,In_1335,In_980);
nor U2243 (N_2243,In_848,In_1437);
nor U2244 (N_2244,In_1502,In_2219);
or U2245 (N_2245,In_858,In_1540);
and U2246 (N_2246,In_1482,In_1619);
or U2247 (N_2247,In_1412,In_1536);
nand U2248 (N_2248,In_1027,In_598);
and U2249 (N_2249,In_331,In_394);
nor U2250 (N_2250,In_2204,In_290);
nor U2251 (N_2251,In_47,In_1430);
or U2252 (N_2252,In_969,In_434);
nor U2253 (N_2253,In_1624,In_1032);
nand U2254 (N_2254,In_2378,In_2031);
or U2255 (N_2255,In_1533,In_2401);
nand U2256 (N_2256,In_881,In_889);
or U2257 (N_2257,In_1824,In_736);
nor U2258 (N_2258,In_1675,In_2190);
nand U2259 (N_2259,In_2483,In_1026);
nand U2260 (N_2260,In_1537,In_2190);
nand U2261 (N_2261,In_2149,In_418);
and U2262 (N_2262,In_1024,In_157);
xnor U2263 (N_2263,In_632,In_1263);
nand U2264 (N_2264,In_621,In_154);
nor U2265 (N_2265,In_1397,In_946);
or U2266 (N_2266,In_1096,In_2355);
and U2267 (N_2267,In_1598,In_1082);
nand U2268 (N_2268,In_562,In_947);
nand U2269 (N_2269,In_2449,In_1106);
nand U2270 (N_2270,In_261,In_1577);
or U2271 (N_2271,In_2118,In_1);
xor U2272 (N_2272,In_87,In_1224);
and U2273 (N_2273,In_1607,In_1155);
and U2274 (N_2274,In_1529,In_2071);
nand U2275 (N_2275,In_581,In_834);
and U2276 (N_2276,In_1466,In_1084);
and U2277 (N_2277,In_1511,In_2446);
or U2278 (N_2278,In_632,In_2331);
nand U2279 (N_2279,In_1944,In_2);
and U2280 (N_2280,In_2066,In_1278);
nor U2281 (N_2281,In_102,In_2279);
and U2282 (N_2282,In_766,In_994);
nor U2283 (N_2283,In_1886,In_1316);
nand U2284 (N_2284,In_700,In_2205);
nand U2285 (N_2285,In_2276,In_1553);
and U2286 (N_2286,In_1532,In_1850);
nor U2287 (N_2287,In_1000,In_861);
nor U2288 (N_2288,In_1921,In_1174);
nand U2289 (N_2289,In_2152,In_580);
and U2290 (N_2290,In_1877,In_167);
xnor U2291 (N_2291,In_881,In_2473);
and U2292 (N_2292,In_1866,In_1399);
and U2293 (N_2293,In_673,In_1701);
nor U2294 (N_2294,In_1007,In_1274);
nor U2295 (N_2295,In_1695,In_1055);
nor U2296 (N_2296,In_1702,In_448);
nand U2297 (N_2297,In_302,In_1967);
and U2298 (N_2298,In_1685,In_832);
nor U2299 (N_2299,In_848,In_205);
and U2300 (N_2300,In_2139,In_1193);
or U2301 (N_2301,In_613,In_354);
or U2302 (N_2302,In_981,In_1836);
and U2303 (N_2303,In_509,In_1442);
nor U2304 (N_2304,In_1039,In_367);
nor U2305 (N_2305,In_638,In_1029);
and U2306 (N_2306,In_412,In_158);
or U2307 (N_2307,In_1575,In_1102);
nand U2308 (N_2308,In_462,In_1893);
xor U2309 (N_2309,In_1690,In_2185);
nand U2310 (N_2310,In_822,In_263);
or U2311 (N_2311,In_2168,In_2328);
nor U2312 (N_2312,In_1820,In_1993);
and U2313 (N_2313,In_315,In_2487);
or U2314 (N_2314,In_1161,In_390);
or U2315 (N_2315,In_1801,In_1573);
nand U2316 (N_2316,In_2362,In_1416);
or U2317 (N_2317,In_129,In_71);
nor U2318 (N_2318,In_251,In_1290);
nand U2319 (N_2319,In_765,In_1282);
or U2320 (N_2320,In_1809,In_1292);
nand U2321 (N_2321,In_919,In_1269);
or U2322 (N_2322,In_1632,In_2476);
or U2323 (N_2323,In_293,In_1718);
nor U2324 (N_2324,In_2212,In_2176);
nor U2325 (N_2325,In_1958,In_384);
nor U2326 (N_2326,In_2225,In_2137);
nand U2327 (N_2327,In_1824,In_2168);
or U2328 (N_2328,In_1748,In_2166);
nor U2329 (N_2329,In_2108,In_349);
nand U2330 (N_2330,In_1736,In_393);
nor U2331 (N_2331,In_2276,In_27);
nor U2332 (N_2332,In_434,In_2018);
nor U2333 (N_2333,In_130,In_425);
nand U2334 (N_2334,In_315,In_155);
nor U2335 (N_2335,In_904,In_1679);
nand U2336 (N_2336,In_2090,In_144);
nand U2337 (N_2337,In_1886,In_166);
or U2338 (N_2338,In_2319,In_1878);
and U2339 (N_2339,In_542,In_1786);
and U2340 (N_2340,In_967,In_1222);
or U2341 (N_2341,In_1989,In_2028);
nand U2342 (N_2342,In_186,In_953);
nand U2343 (N_2343,In_834,In_1540);
nand U2344 (N_2344,In_1722,In_1274);
and U2345 (N_2345,In_2222,In_604);
nor U2346 (N_2346,In_457,In_738);
or U2347 (N_2347,In_183,In_2357);
xor U2348 (N_2348,In_58,In_2150);
nand U2349 (N_2349,In_403,In_2121);
nand U2350 (N_2350,In_114,In_231);
and U2351 (N_2351,In_1423,In_1319);
nand U2352 (N_2352,In_2287,In_2250);
and U2353 (N_2353,In_1620,In_486);
and U2354 (N_2354,In_662,In_707);
and U2355 (N_2355,In_224,In_154);
nor U2356 (N_2356,In_270,In_1662);
xor U2357 (N_2357,In_2191,In_565);
nand U2358 (N_2358,In_606,In_833);
or U2359 (N_2359,In_2076,In_1368);
and U2360 (N_2360,In_1632,In_1245);
nor U2361 (N_2361,In_1347,In_2347);
and U2362 (N_2362,In_39,In_265);
xnor U2363 (N_2363,In_850,In_1157);
and U2364 (N_2364,In_572,In_759);
or U2365 (N_2365,In_54,In_2394);
and U2366 (N_2366,In_540,In_2486);
and U2367 (N_2367,In_2466,In_1191);
or U2368 (N_2368,In_1816,In_1446);
or U2369 (N_2369,In_286,In_1969);
or U2370 (N_2370,In_6,In_1697);
or U2371 (N_2371,In_1801,In_914);
nand U2372 (N_2372,In_2093,In_2336);
nand U2373 (N_2373,In_528,In_1036);
or U2374 (N_2374,In_239,In_1848);
or U2375 (N_2375,In_1959,In_2160);
and U2376 (N_2376,In_2479,In_81);
and U2377 (N_2377,In_1073,In_1723);
nand U2378 (N_2378,In_894,In_62);
and U2379 (N_2379,In_808,In_211);
and U2380 (N_2380,In_344,In_1097);
nor U2381 (N_2381,In_703,In_2438);
nor U2382 (N_2382,In_768,In_1236);
or U2383 (N_2383,In_2018,In_2369);
or U2384 (N_2384,In_1406,In_2435);
or U2385 (N_2385,In_1482,In_1187);
nor U2386 (N_2386,In_1827,In_1385);
xor U2387 (N_2387,In_60,In_1253);
and U2388 (N_2388,In_1089,In_2264);
and U2389 (N_2389,In_1345,In_2409);
nor U2390 (N_2390,In_2296,In_2470);
and U2391 (N_2391,In_354,In_1176);
and U2392 (N_2392,In_278,In_1737);
nand U2393 (N_2393,In_865,In_1526);
or U2394 (N_2394,In_1124,In_1221);
nor U2395 (N_2395,In_65,In_733);
and U2396 (N_2396,In_271,In_2206);
nand U2397 (N_2397,In_221,In_1134);
or U2398 (N_2398,In_1520,In_349);
nand U2399 (N_2399,In_1617,In_1799);
nand U2400 (N_2400,In_885,In_547);
or U2401 (N_2401,In_640,In_720);
or U2402 (N_2402,In_1500,In_2137);
xor U2403 (N_2403,In_676,In_1558);
or U2404 (N_2404,In_1497,In_200);
and U2405 (N_2405,In_301,In_468);
nand U2406 (N_2406,In_521,In_1082);
xnor U2407 (N_2407,In_191,In_593);
and U2408 (N_2408,In_1756,In_429);
nand U2409 (N_2409,In_2337,In_1830);
and U2410 (N_2410,In_1778,In_1633);
or U2411 (N_2411,In_603,In_2308);
nand U2412 (N_2412,In_1291,In_1607);
xnor U2413 (N_2413,In_268,In_1540);
and U2414 (N_2414,In_2173,In_909);
nor U2415 (N_2415,In_2163,In_1134);
or U2416 (N_2416,In_1118,In_1479);
nand U2417 (N_2417,In_2455,In_724);
nand U2418 (N_2418,In_1153,In_1225);
xor U2419 (N_2419,In_1473,In_1584);
or U2420 (N_2420,In_1185,In_2373);
nand U2421 (N_2421,In_1603,In_1258);
xnor U2422 (N_2422,In_1668,In_2217);
and U2423 (N_2423,In_149,In_2363);
and U2424 (N_2424,In_1657,In_2106);
or U2425 (N_2425,In_1336,In_1955);
nand U2426 (N_2426,In_558,In_1603);
nor U2427 (N_2427,In_2496,In_2008);
and U2428 (N_2428,In_371,In_2006);
nor U2429 (N_2429,In_1899,In_729);
xnor U2430 (N_2430,In_742,In_351);
and U2431 (N_2431,In_51,In_1317);
or U2432 (N_2432,In_1278,In_89);
or U2433 (N_2433,In_1682,In_680);
nor U2434 (N_2434,In_989,In_772);
nand U2435 (N_2435,In_552,In_1757);
and U2436 (N_2436,In_1562,In_1284);
xnor U2437 (N_2437,In_2395,In_891);
and U2438 (N_2438,In_1071,In_2076);
nor U2439 (N_2439,In_1936,In_955);
xor U2440 (N_2440,In_1682,In_212);
and U2441 (N_2441,In_1015,In_935);
and U2442 (N_2442,In_1397,In_1538);
and U2443 (N_2443,In_806,In_1677);
and U2444 (N_2444,In_2308,In_856);
nor U2445 (N_2445,In_856,In_98);
or U2446 (N_2446,In_555,In_1568);
or U2447 (N_2447,In_587,In_1004);
nor U2448 (N_2448,In_2254,In_1403);
and U2449 (N_2449,In_887,In_1467);
and U2450 (N_2450,In_507,In_2183);
nor U2451 (N_2451,In_2450,In_536);
and U2452 (N_2452,In_1492,In_31);
nand U2453 (N_2453,In_590,In_880);
nor U2454 (N_2454,In_370,In_1584);
or U2455 (N_2455,In_2475,In_2097);
nand U2456 (N_2456,In_2043,In_1344);
and U2457 (N_2457,In_1181,In_1375);
nor U2458 (N_2458,In_660,In_338);
and U2459 (N_2459,In_1667,In_356);
nand U2460 (N_2460,In_1450,In_232);
and U2461 (N_2461,In_2068,In_1864);
nand U2462 (N_2462,In_1672,In_2425);
nor U2463 (N_2463,In_740,In_1251);
nand U2464 (N_2464,In_1660,In_933);
nand U2465 (N_2465,In_1179,In_679);
nand U2466 (N_2466,In_16,In_385);
and U2467 (N_2467,In_304,In_205);
or U2468 (N_2468,In_1109,In_762);
nand U2469 (N_2469,In_557,In_1216);
or U2470 (N_2470,In_2217,In_1937);
and U2471 (N_2471,In_124,In_307);
nand U2472 (N_2472,In_502,In_546);
or U2473 (N_2473,In_1202,In_2463);
nor U2474 (N_2474,In_768,In_633);
and U2475 (N_2475,In_1049,In_1196);
or U2476 (N_2476,In_576,In_1619);
xor U2477 (N_2477,In_1590,In_2269);
or U2478 (N_2478,In_1099,In_2434);
and U2479 (N_2479,In_114,In_449);
nand U2480 (N_2480,In_1299,In_1250);
and U2481 (N_2481,In_611,In_882);
nor U2482 (N_2482,In_1016,In_1601);
or U2483 (N_2483,In_1431,In_2112);
or U2484 (N_2484,In_2119,In_2019);
nand U2485 (N_2485,In_571,In_1580);
and U2486 (N_2486,In_567,In_227);
or U2487 (N_2487,In_1988,In_1853);
and U2488 (N_2488,In_1882,In_516);
nand U2489 (N_2489,In_1778,In_1106);
nand U2490 (N_2490,In_1675,In_302);
or U2491 (N_2491,In_182,In_2226);
nor U2492 (N_2492,In_1101,In_759);
nand U2493 (N_2493,In_485,In_576);
nand U2494 (N_2494,In_1206,In_355);
and U2495 (N_2495,In_2063,In_1417);
or U2496 (N_2496,In_209,In_1063);
nor U2497 (N_2497,In_734,In_338);
and U2498 (N_2498,In_1117,In_196);
nor U2499 (N_2499,In_1494,In_221);
nand U2500 (N_2500,In_1079,In_2426);
nand U2501 (N_2501,In_1199,In_2177);
and U2502 (N_2502,In_163,In_1176);
or U2503 (N_2503,In_1654,In_728);
nand U2504 (N_2504,In_201,In_140);
or U2505 (N_2505,In_2366,In_1904);
nand U2506 (N_2506,In_752,In_557);
or U2507 (N_2507,In_2327,In_587);
nor U2508 (N_2508,In_1520,In_2476);
and U2509 (N_2509,In_1370,In_44);
nand U2510 (N_2510,In_840,In_2454);
or U2511 (N_2511,In_1241,In_366);
and U2512 (N_2512,In_1020,In_113);
nor U2513 (N_2513,In_137,In_261);
nand U2514 (N_2514,In_1517,In_434);
nand U2515 (N_2515,In_1173,In_2028);
nor U2516 (N_2516,In_132,In_970);
nand U2517 (N_2517,In_2301,In_3);
or U2518 (N_2518,In_1743,In_2398);
or U2519 (N_2519,In_912,In_1133);
nor U2520 (N_2520,In_390,In_921);
and U2521 (N_2521,In_1383,In_1789);
or U2522 (N_2522,In_1783,In_600);
nand U2523 (N_2523,In_1433,In_2179);
or U2524 (N_2524,In_373,In_1248);
and U2525 (N_2525,In_198,In_1339);
nor U2526 (N_2526,In_2419,In_1255);
and U2527 (N_2527,In_620,In_151);
and U2528 (N_2528,In_89,In_1532);
and U2529 (N_2529,In_1925,In_30);
xnor U2530 (N_2530,In_884,In_1324);
or U2531 (N_2531,In_1109,In_504);
nor U2532 (N_2532,In_1968,In_861);
xnor U2533 (N_2533,In_202,In_1132);
nand U2534 (N_2534,In_438,In_1890);
or U2535 (N_2535,In_405,In_391);
nand U2536 (N_2536,In_1569,In_627);
or U2537 (N_2537,In_211,In_1739);
nor U2538 (N_2538,In_1122,In_596);
or U2539 (N_2539,In_930,In_2356);
nor U2540 (N_2540,In_2046,In_92);
xor U2541 (N_2541,In_98,In_1071);
nand U2542 (N_2542,In_1233,In_2353);
nand U2543 (N_2543,In_768,In_1378);
nand U2544 (N_2544,In_76,In_1910);
nor U2545 (N_2545,In_2434,In_2283);
nor U2546 (N_2546,In_2459,In_1674);
nand U2547 (N_2547,In_963,In_1965);
nand U2548 (N_2548,In_424,In_861);
or U2549 (N_2549,In_1814,In_1657);
nand U2550 (N_2550,In_1397,In_1889);
xor U2551 (N_2551,In_237,In_578);
or U2552 (N_2552,In_2374,In_2430);
nor U2553 (N_2553,In_2145,In_1706);
nand U2554 (N_2554,In_2348,In_1917);
nand U2555 (N_2555,In_587,In_1516);
nand U2556 (N_2556,In_789,In_2205);
and U2557 (N_2557,In_760,In_1406);
or U2558 (N_2558,In_1109,In_369);
nand U2559 (N_2559,In_1199,In_887);
xor U2560 (N_2560,In_1378,In_2031);
xnor U2561 (N_2561,In_1267,In_68);
nand U2562 (N_2562,In_1057,In_149);
nand U2563 (N_2563,In_407,In_1100);
nor U2564 (N_2564,In_779,In_1999);
or U2565 (N_2565,In_433,In_2416);
and U2566 (N_2566,In_1300,In_2452);
and U2567 (N_2567,In_1764,In_2081);
and U2568 (N_2568,In_1786,In_2281);
or U2569 (N_2569,In_2446,In_332);
nor U2570 (N_2570,In_968,In_1230);
nand U2571 (N_2571,In_36,In_189);
nor U2572 (N_2572,In_891,In_1951);
xor U2573 (N_2573,In_353,In_272);
nor U2574 (N_2574,In_1873,In_1755);
nand U2575 (N_2575,In_1764,In_1744);
and U2576 (N_2576,In_680,In_1933);
nand U2577 (N_2577,In_93,In_1862);
and U2578 (N_2578,In_1781,In_1430);
or U2579 (N_2579,In_31,In_2268);
and U2580 (N_2580,In_1595,In_986);
nor U2581 (N_2581,In_965,In_292);
or U2582 (N_2582,In_1615,In_2248);
or U2583 (N_2583,In_1850,In_971);
and U2584 (N_2584,In_2459,In_2356);
or U2585 (N_2585,In_160,In_189);
nand U2586 (N_2586,In_1855,In_2040);
nand U2587 (N_2587,In_1973,In_1556);
and U2588 (N_2588,In_1406,In_795);
nor U2589 (N_2589,In_1727,In_2182);
and U2590 (N_2590,In_1469,In_1516);
and U2591 (N_2591,In_2263,In_1983);
xor U2592 (N_2592,In_2182,In_1774);
nor U2593 (N_2593,In_334,In_911);
and U2594 (N_2594,In_1126,In_2026);
or U2595 (N_2595,In_1151,In_2075);
nand U2596 (N_2596,In_1850,In_1810);
xnor U2597 (N_2597,In_259,In_1860);
and U2598 (N_2598,In_1505,In_822);
or U2599 (N_2599,In_62,In_2326);
or U2600 (N_2600,In_24,In_239);
or U2601 (N_2601,In_1773,In_173);
nand U2602 (N_2602,In_824,In_799);
xnor U2603 (N_2603,In_561,In_1014);
and U2604 (N_2604,In_1153,In_724);
nand U2605 (N_2605,In_1020,In_282);
nor U2606 (N_2606,In_1024,In_1847);
xnor U2607 (N_2607,In_2025,In_1199);
or U2608 (N_2608,In_1129,In_564);
xor U2609 (N_2609,In_453,In_467);
or U2610 (N_2610,In_1066,In_2470);
nor U2611 (N_2611,In_2392,In_12);
and U2612 (N_2612,In_899,In_644);
and U2613 (N_2613,In_980,In_2110);
xor U2614 (N_2614,In_1041,In_2284);
and U2615 (N_2615,In_1765,In_682);
or U2616 (N_2616,In_916,In_1049);
nand U2617 (N_2617,In_336,In_54);
or U2618 (N_2618,In_1181,In_1439);
and U2619 (N_2619,In_158,In_1926);
nor U2620 (N_2620,In_540,In_2208);
or U2621 (N_2621,In_1709,In_1353);
and U2622 (N_2622,In_2053,In_2339);
nand U2623 (N_2623,In_211,In_2100);
or U2624 (N_2624,In_1405,In_2328);
nor U2625 (N_2625,In_1010,In_1696);
nand U2626 (N_2626,In_2263,In_1950);
nand U2627 (N_2627,In_2488,In_1893);
xor U2628 (N_2628,In_2109,In_1466);
nand U2629 (N_2629,In_1120,In_771);
nand U2630 (N_2630,In_556,In_2098);
xor U2631 (N_2631,In_1019,In_1223);
or U2632 (N_2632,In_660,In_468);
and U2633 (N_2633,In_1044,In_1063);
nor U2634 (N_2634,In_1931,In_1671);
nand U2635 (N_2635,In_635,In_1656);
xnor U2636 (N_2636,In_1737,In_83);
nor U2637 (N_2637,In_1585,In_1204);
and U2638 (N_2638,In_2001,In_2015);
or U2639 (N_2639,In_572,In_481);
and U2640 (N_2640,In_1631,In_1329);
nor U2641 (N_2641,In_787,In_1133);
and U2642 (N_2642,In_1935,In_36);
nor U2643 (N_2643,In_996,In_619);
nor U2644 (N_2644,In_1693,In_348);
or U2645 (N_2645,In_1778,In_2451);
nand U2646 (N_2646,In_862,In_2111);
and U2647 (N_2647,In_1289,In_2194);
and U2648 (N_2648,In_2185,In_2499);
nor U2649 (N_2649,In_1922,In_1183);
or U2650 (N_2650,In_492,In_1731);
xor U2651 (N_2651,In_2364,In_653);
nor U2652 (N_2652,In_1061,In_589);
nand U2653 (N_2653,In_1269,In_1070);
and U2654 (N_2654,In_2321,In_1291);
and U2655 (N_2655,In_2196,In_1169);
nor U2656 (N_2656,In_187,In_2118);
nand U2657 (N_2657,In_242,In_2188);
and U2658 (N_2658,In_318,In_987);
and U2659 (N_2659,In_389,In_1045);
nor U2660 (N_2660,In_1437,In_1708);
nand U2661 (N_2661,In_301,In_286);
and U2662 (N_2662,In_2372,In_1466);
nand U2663 (N_2663,In_1716,In_169);
nor U2664 (N_2664,In_1836,In_2062);
nand U2665 (N_2665,In_1631,In_2348);
and U2666 (N_2666,In_1230,In_2114);
nor U2667 (N_2667,In_2349,In_2322);
and U2668 (N_2668,In_133,In_1758);
and U2669 (N_2669,In_1918,In_1268);
nor U2670 (N_2670,In_191,In_1678);
or U2671 (N_2671,In_2464,In_1315);
or U2672 (N_2672,In_2005,In_395);
nand U2673 (N_2673,In_1191,In_1438);
or U2674 (N_2674,In_550,In_742);
nor U2675 (N_2675,In_917,In_1185);
nor U2676 (N_2676,In_1180,In_375);
and U2677 (N_2677,In_2042,In_274);
nand U2678 (N_2678,In_1194,In_336);
or U2679 (N_2679,In_2,In_2373);
or U2680 (N_2680,In_446,In_22);
xnor U2681 (N_2681,In_1116,In_667);
nand U2682 (N_2682,In_245,In_538);
nor U2683 (N_2683,In_2150,In_2489);
nor U2684 (N_2684,In_1458,In_1849);
or U2685 (N_2685,In_662,In_129);
nor U2686 (N_2686,In_313,In_1339);
nand U2687 (N_2687,In_2281,In_275);
xnor U2688 (N_2688,In_2172,In_2075);
or U2689 (N_2689,In_429,In_2275);
or U2690 (N_2690,In_1966,In_2386);
or U2691 (N_2691,In_156,In_1940);
nand U2692 (N_2692,In_209,In_1304);
nand U2693 (N_2693,In_801,In_957);
nand U2694 (N_2694,In_138,In_646);
nor U2695 (N_2695,In_1483,In_306);
and U2696 (N_2696,In_1842,In_2468);
or U2697 (N_2697,In_2252,In_733);
nor U2698 (N_2698,In_1609,In_1800);
or U2699 (N_2699,In_26,In_986);
and U2700 (N_2700,In_1213,In_307);
xnor U2701 (N_2701,In_2012,In_2122);
or U2702 (N_2702,In_2306,In_1638);
and U2703 (N_2703,In_1508,In_1234);
nand U2704 (N_2704,In_1184,In_1823);
and U2705 (N_2705,In_2339,In_713);
nand U2706 (N_2706,In_1913,In_101);
and U2707 (N_2707,In_1791,In_474);
nor U2708 (N_2708,In_231,In_723);
or U2709 (N_2709,In_1294,In_1330);
and U2710 (N_2710,In_1052,In_30);
or U2711 (N_2711,In_369,In_45);
or U2712 (N_2712,In_549,In_976);
and U2713 (N_2713,In_2085,In_990);
nand U2714 (N_2714,In_223,In_776);
or U2715 (N_2715,In_2161,In_258);
and U2716 (N_2716,In_2273,In_2274);
nor U2717 (N_2717,In_1869,In_1930);
or U2718 (N_2718,In_1089,In_872);
nand U2719 (N_2719,In_987,In_2187);
xnor U2720 (N_2720,In_1853,In_608);
or U2721 (N_2721,In_649,In_2459);
nand U2722 (N_2722,In_1304,In_1136);
and U2723 (N_2723,In_1209,In_360);
nor U2724 (N_2724,In_174,In_2415);
nor U2725 (N_2725,In_2492,In_410);
nor U2726 (N_2726,In_1246,In_499);
nor U2727 (N_2727,In_1881,In_312);
and U2728 (N_2728,In_2150,In_1586);
or U2729 (N_2729,In_1923,In_308);
or U2730 (N_2730,In_1419,In_1288);
or U2731 (N_2731,In_870,In_1216);
xor U2732 (N_2732,In_1725,In_2322);
nand U2733 (N_2733,In_545,In_2013);
nand U2734 (N_2734,In_663,In_2445);
nor U2735 (N_2735,In_1365,In_2321);
nor U2736 (N_2736,In_399,In_1291);
nor U2737 (N_2737,In_1871,In_470);
or U2738 (N_2738,In_2015,In_2044);
nor U2739 (N_2739,In_1941,In_479);
and U2740 (N_2740,In_1004,In_1651);
or U2741 (N_2741,In_2232,In_890);
and U2742 (N_2742,In_495,In_2449);
or U2743 (N_2743,In_2179,In_885);
or U2744 (N_2744,In_1248,In_1262);
xor U2745 (N_2745,In_856,In_185);
nand U2746 (N_2746,In_1889,In_930);
or U2747 (N_2747,In_613,In_1078);
and U2748 (N_2748,In_382,In_1816);
xor U2749 (N_2749,In_1187,In_981);
or U2750 (N_2750,In_1438,In_224);
and U2751 (N_2751,In_12,In_2128);
and U2752 (N_2752,In_2300,In_2351);
or U2753 (N_2753,In_524,In_188);
or U2754 (N_2754,In_1794,In_1183);
nor U2755 (N_2755,In_1731,In_757);
nand U2756 (N_2756,In_1164,In_1691);
nor U2757 (N_2757,In_520,In_932);
nor U2758 (N_2758,In_847,In_1277);
xnor U2759 (N_2759,In_2005,In_759);
nand U2760 (N_2760,In_1817,In_1221);
or U2761 (N_2761,In_1851,In_227);
and U2762 (N_2762,In_1206,In_1368);
nor U2763 (N_2763,In_455,In_2339);
and U2764 (N_2764,In_2496,In_1295);
nand U2765 (N_2765,In_1603,In_458);
nor U2766 (N_2766,In_1675,In_1678);
nand U2767 (N_2767,In_180,In_1273);
and U2768 (N_2768,In_596,In_2399);
nand U2769 (N_2769,In_534,In_244);
and U2770 (N_2770,In_1871,In_641);
nor U2771 (N_2771,In_1408,In_81);
nor U2772 (N_2772,In_1262,In_2085);
and U2773 (N_2773,In_2118,In_1341);
xor U2774 (N_2774,In_2424,In_1988);
or U2775 (N_2775,In_1411,In_2301);
and U2776 (N_2776,In_823,In_348);
nor U2777 (N_2777,In_1941,In_952);
nor U2778 (N_2778,In_139,In_806);
xnor U2779 (N_2779,In_196,In_1543);
nand U2780 (N_2780,In_1604,In_564);
nand U2781 (N_2781,In_281,In_2143);
or U2782 (N_2782,In_971,In_683);
or U2783 (N_2783,In_2319,In_302);
or U2784 (N_2784,In_991,In_68);
nand U2785 (N_2785,In_59,In_1703);
nand U2786 (N_2786,In_2121,In_442);
or U2787 (N_2787,In_2172,In_102);
and U2788 (N_2788,In_382,In_671);
nand U2789 (N_2789,In_1916,In_755);
nor U2790 (N_2790,In_1214,In_1944);
xnor U2791 (N_2791,In_642,In_2099);
nand U2792 (N_2792,In_2267,In_12);
or U2793 (N_2793,In_997,In_874);
or U2794 (N_2794,In_1211,In_869);
and U2795 (N_2795,In_1136,In_216);
and U2796 (N_2796,In_924,In_1213);
or U2797 (N_2797,In_206,In_378);
and U2798 (N_2798,In_111,In_2115);
and U2799 (N_2799,In_1720,In_2420);
nor U2800 (N_2800,In_2214,In_1861);
and U2801 (N_2801,In_87,In_1935);
nor U2802 (N_2802,In_218,In_132);
nand U2803 (N_2803,In_819,In_2463);
xor U2804 (N_2804,In_1798,In_1875);
and U2805 (N_2805,In_1873,In_1212);
nand U2806 (N_2806,In_438,In_334);
and U2807 (N_2807,In_1860,In_672);
or U2808 (N_2808,In_229,In_1349);
and U2809 (N_2809,In_2257,In_1171);
xnor U2810 (N_2810,In_1327,In_958);
xor U2811 (N_2811,In_1674,In_401);
or U2812 (N_2812,In_2132,In_1458);
and U2813 (N_2813,In_1395,In_2056);
xnor U2814 (N_2814,In_2036,In_1721);
nor U2815 (N_2815,In_1563,In_794);
and U2816 (N_2816,In_159,In_932);
and U2817 (N_2817,In_2251,In_1793);
and U2818 (N_2818,In_1964,In_343);
and U2819 (N_2819,In_1604,In_513);
and U2820 (N_2820,In_2313,In_2033);
nand U2821 (N_2821,In_1327,In_263);
xnor U2822 (N_2822,In_907,In_2404);
nor U2823 (N_2823,In_2294,In_1945);
and U2824 (N_2824,In_1634,In_173);
nor U2825 (N_2825,In_568,In_1834);
or U2826 (N_2826,In_172,In_177);
nor U2827 (N_2827,In_1796,In_485);
and U2828 (N_2828,In_404,In_1763);
and U2829 (N_2829,In_809,In_1170);
and U2830 (N_2830,In_2348,In_998);
or U2831 (N_2831,In_1739,In_1694);
and U2832 (N_2832,In_2436,In_2399);
xnor U2833 (N_2833,In_335,In_470);
nor U2834 (N_2834,In_647,In_2268);
or U2835 (N_2835,In_2059,In_546);
and U2836 (N_2836,In_1533,In_644);
or U2837 (N_2837,In_1394,In_2472);
xnor U2838 (N_2838,In_559,In_1261);
and U2839 (N_2839,In_1009,In_147);
and U2840 (N_2840,In_1231,In_1427);
xor U2841 (N_2841,In_233,In_1957);
nand U2842 (N_2842,In_1780,In_1437);
and U2843 (N_2843,In_39,In_1653);
nor U2844 (N_2844,In_411,In_1535);
nor U2845 (N_2845,In_1178,In_403);
and U2846 (N_2846,In_930,In_1820);
nor U2847 (N_2847,In_445,In_1307);
nand U2848 (N_2848,In_741,In_864);
and U2849 (N_2849,In_115,In_1933);
nand U2850 (N_2850,In_1517,In_1536);
or U2851 (N_2851,In_2051,In_246);
and U2852 (N_2852,In_1087,In_1196);
nand U2853 (N_2853,In_445,In_97);
and U2854 (N_2854,In_1179,In_1430);
nor U2855 (N_2855,In_386,In_997);
and U2856 (N_2856,In_771,In_1253);
nor U2857 (N_2857,In_1748,In_1652);
nand U2858 (N_2858,In_1272,In_2285);
or U2859 (N_2859,In_2357,In_1161);
nand U2860 (N_2860,In_2347,In_2139);
and U2861 (N_2861,In_1270,In_998);
and U2862 (N_2862,In_1865,In_1058);
nor U2863 (N_2863,In_36,In_1433);
nand U2864 (N_2864,In_1284,In_1488);
or U2865 (N_2865,In_605,In_1567);
nand U2866 (N_2866,In_1156,In_1950);
or U2867 (N_2867,In_1836,In_1674);
nand U2868 (N_2868,In_1369,In_414);
or U2869 (N_2869,In_1540,In_1712);
or U2870 (N_2870,In_1380,In_953);
nor U2871 (N_2871,In_1009,In_1686);
nor U2872 (N_2872,In_2111,In_1828);
nand U2873 (N_2873,In_514,In_1891);
nand U2874 (N_2874,In_1763,In_1454);
xor U2875 (N_2875,In_1627,In_1785);
xnor U2876 (N_2876,In_2105,In_136);
xor U2877 (N_2877,In_63,In_1570);
nor U2878 (N_2878,In_498,In_69);
or U2879 (N_2879,In_2218,In_422);
and U2880 (N_2880,In_1183,In_535);
and U2881 (N_2881,In_1384,In_2);
xnor U2882 (N_2882,In_2213,In_1914);
or U2883 (N_2883,In_694,In_949);
xor U2884 (N_2884,In_2051,In_2223);
nand U2885 (N_2885,In_1936,In_2126);
and U2886 (N_2886,In_80,In_2462);
and U2887 (N_2887,In_482,In_2319);
nand U2888 (N_2888,In_1400,In_437);
or U2889 (N_2889,In_2200,In_1245);
nor U2890 (N_2890,In_2247,In_2000);
nand U2891 (N_2891,In_2364,In_1209);
nand U2892 (N_2892,In_4,In_2176);
nand U2893 (N_2893,In_2256,In_918);
or U2894 (N_2894,In_2349,In_294);
and U2895 (N_2895,In_1912,In_660);
and U2896 (N_2896,In_1193,In_571);
nor U2897 (N_2897,In_578,In_837);
nor U2898 (N_2898,In_113,In_1383);
nor U2899 (N_2899,In_898,In_35);
nor U2900 (N_2900,In_135,In_1758);
or U2901 (N_2901,In_1528,In_1145);
nand U2902 (N_2902,In_1389,In_2011);
and U2903 (N_2903,In_477,In_1455);
nand U2904 (N_2904,In_1675,In_64);
nand U2905 (N_2905,In_95,In_791);
nor U2906 (N_2906,In_2039,In_1185);
or U2907 (N_2907,In_233,In_1088);
and U2908 (N_2908,In_1534,In_154);
nand U2909 (N_2909,In_1998,In_2451);
xor U2910 (N_2910,In_2145,In_1222);
nand U2911 (N_2911,In_573,In_2306);
nand U2912 (N_2912,In_1790,In_1155);
and U2913 (N_2913,In_221,In_2497);
nor U2914 (N_2914,In_2059,In_1806);
and U2915 (N_2915,In_1724,In_1653);
nor U2916 (N_2916,In_810,In_2195);
or U2917 (N_2917,In_48,In_989);
or U2918 (N_2918,In_774,In_1335);
nor U2919 (N_2919,In_745,In_268);
nor U2920 (N_2920,In_1171,In_1859);
nor U2921 (N_2921,In_2476,In_1987);
nor U2922 (N_2922,In_474,In_1157);
nor U2923 (N_2923,In_1949,In_396);
or U2924 (N_2924,In_1199,In_1209);
nand U2925 (N_2925,In_1398,In_175);
nor U2926 (N_2926,In_2093,In_728);
nor U2927 (N_2927,In_2167,In_2090);
and U2928 (N_2928,In_937,In_927);
nand U2929 (N_2929,In_400,In_658);
and U2930 (N_2930,In_1914,In_1199);
nand U2931 (N_2931,In_2317,In_557);
and U2932 (N_2932,In_342,In_64);
or U2933 (N_2933,In_1596,In_67);
or U2934 (N_2934,In_578,In_634);
or U2935 (N_2935,In_1701,In_2423);
nor U2936 (N_2936,In_1369,In_1816);
or U2937 (N_2937,In_1957,In_1421);
xnor U2938 (N_2938,In_1533,In_442);
or U2939 (N_2939,In_1187,In_1196);
or U2940 (N_2940,In_1156,In_1070);
nand U2941 (N_2941,In_864,In_661);
and U2942 (N_2942,In_1751,In_2183);
and U2943 (N_2943,In_627,In_1863);
nand U2944 (N_2944,In_1707,In_1017);
nor U2945 (N_2945,In_2393,In_539);
or U2946 (N_2946,In_1524,In_2284);
nor U2947 (N_2947,In_160,In_1195);
nand U2948 (N_2948,In_519,In_216);
nor U2949 (N_2949,In_2146,In_1403);
and U2950 (N_2950,In_588,In_1193);
nor U2951 (N_2951,In_1731,In_776);
nor U2952 (N_2952,In_2109,In_1935);
or U2953 (N_2953,In_1467,In_2318);
xor U2954 (N_2954,In_2325,In_632);
nand U2955 (N_2955,In_894,In_2405);
nand U2956 (N_2956,In_29,In_1878);
xor U2957 (N_2957,In_500,In_596);
nor U2958 (N_2958,In_1092,In_1109);
or U2959 (N_2959,In_880,In_288);
nor U2960 (N_2960,In_495,In_198);
and U2961 (N_2961,In_1961,In_671);
xor U2962 (N_2962,In_1461,In_2353);
or U2963 (N_2963,In_300,In_369);
and U2964 (N_2964,In_150,In_94);
or U2965 (N_2965,In_643,In_386);
or U2966 (N_2966,In_174,In_1930);
nand U2967 (N_2967,In_768,In_2468);
or U2968 (N_2968,In_107,In_1979);
xnor U2969 (N_2969,In_612,In_2025);
and U2970 (N_2970,In_1282,In_1005);
xnor U2971 (N_2971,In_929,In_237);
or U2972 (N_2972,In_838,In_2173);
nand U2973 (N_2973,In_2081,In_2254);
nand U2974 (N_2974,In_843,In_1277);
xor U2975 (N_2975,In_13,In_395);
or U2976 (N_2976,In_855,In_1107);
and U2977 (N_2977,In_2446,In_1912);
nand U2978 (N_2978,In_1209,In_1226);
nand U2979 (N_2979,In_2428,In_39);
xnor U2980 (N_2980,In_749,In_2365);
nor U2981 (N_2981,In_1228,In_1520);
nand U2982 (N_2982,In_1236,In_164);
and U2983 (N_2983,In_1219,In_2);
or U2984 (N_2984,In_780,In_771);
xnor U2985 (N_2985,In_1242,In_1722);
and U2986 (N_2986,In_2258,In_1221);
xnor U2987 (N_2987,In_1041,In_1258);
and U2988 (N_2988,In_772,In_1513);
nor U2989 (N_2989,In_948,In_820);
and U2990 (N_2990,In_1636,In_16);
nor U2991 (N_2991,In_95,In_1475);
nand U2992 (N_2992,In_1909,In_1303);
nor U2993 (N_2993,In_967,In_2081);
or U2994 (N_2994,In_2020,In_1738);
nor U2995 (N_2995,In_913,In_1045);
and U2996 (N_2996,In_680,In_1038);
xor U2997 (N_2997,In_1560,In_474);
xor U2998 (N_2998,In_806,In_2484);
and U2999 (N_2999,In_218,In_1527);
or U3000 (N_3000,In_282,In_1315);
nor U3001 (N_3001,In_1358,In_1708);
or U3002 (N_3002,In_696,In_1613);
xor U3003 (N_3003,In_1547,In_616);
xor U3004 (N_3004,In_2421,In_2263);
xor U3005 (N_3005,In_1380,In_922);
and U3006 (N_3006,In_1117,In_2190);
or U3007 (N_3007,In_841,In_2382);
nor U3008 (N_3008,In_1939,In_1141);
or U3009 (N_3009,In_2465,In_1050);
and U3010 (N_3010,In_606,In_18);
or U3011 (N_3011,In_1975,In_1916);
or U3012 (N_3012,In_1650,In_1163);
nor U3013 (N_3013,In_530,In_1683);
and U3014 (N_3014,In_38,In_989);
and U3015 (N_3015,In_980,In_1178);
or U3016 (N_3016,In_124,In_1347);
nand U3017 (N_3017,In_2459,In_528);
nor U3018 (N_3018,In_1557,In_157);
or U3019 (N_3019,In_935,In_2366);
nor U3020 (N_3020,In_2172,In_2111);
and U3021 (N_3021,In_1743,In_1498);
and U3022 (N_3022,In_901,In_2101);
nand U3023 (N_3023,In_1129,In_504);
nor U3024 (N_3024,In_538,In_2474);
nand U3025 (N_3025,In_629,In_1667);
nand U3026 (N_3026,In_2222,In_1863);
or U3027 (N_3027,In_2372,In_1991);
nor U3028 (N_3028,In_2216,In_983);
nor U3029 (N_3029,In_804,In_703);
nand U3030 (N_3030,In_1459,In_760);
nand U3031 (N_3031,In_1997,In_2189);
or U3032 (N_3032,In_2191,In_959);
nand U3033 (N_3033,In_1433,In_1678);
nand U3034 (N_3034,In_53,In_1724);
or U3035 (N_3035,In_2077,In_1332);
or U3036 (N_3036,In_761,In_1701);
nor U3037 (N_3037,In_1109,In_1130);
nor U3038 (N_3038,In_619,In_2249);
or U3039 (N_3039,In_553,In_1113);
nand U3040 (N_3040,In_924,In_1088);
nand U3041 (N_3041,In_189,In_780);
or U3042 (N_3042,In_2338,In_154);
or U3043 (N_3043,In_1128,In_1152);
nand U3044 (N_3044,In_718,In_1217);
xor U3045 (N_3045,In_2322,In_1899);
xnor U3046 (N_3046,In_596,In_127);
nand U3047 (N_3047,In_165,In_959);
or U3048 (N_3048,In_1750,In_341);
and U3049 (N_3049,In_1223,In_852);
nor U3050 (N_3050,In_1793,In_1421);
or U3051 (N_3051,In_324,In_593);
or U3052 (N_3052,In_1887,In_105);
nand U3053 (N_3053,In_679,In_1442);
nand U3054 (N_3054,In_680,In_7);
xor U3055 (N_3055,In_877,In_2162);
nand U3056 (N_3056,In_526,In_1032);
and U3057 (N_3057,In_735,In_2432);
or U3058 (N_3058,In_2252,In_142);
nor U3059 (N_3059,In_1982,In_2291);
nand U3060 (N_3060,In_141,In_579);
xor U3061 (N_3061,In_438,In_2246);
and U3062 (N_3062,In_754,In_1585);
nand U3063 (N_3063,In_1792,In_2059);
or U3064 (N_3064,In_1436,In_1474);
or U3065 (N_3065,In_750,In_416);
xor U3066 (N_3066,In_1998,In_106);
nand U3067 (N_3067,In_2055,In_2202);
nand U3068 (N_3068,In_2250,In_584);
nand U3069 (N_3069,In_1051,In_2445);
xnor U3070 (N_3070,In_2388,In_2079);
or U3071 (N_3071,In_1572,In_746);
nor U3072 (N_3072,In_2197,In_481);
and U3073 (N_3073,In_2070,In_1478);
or U3074 (N_3074,In_1811,In_2392);
or U3075 (N_3075,In_1284,In_304);
nor U3076 (N_3076,In_125,In_1829);
and U3077 (N_3077,In_577,In_838);
nand U3078 (N_3078,In_1489,In_1877);
and U3079 (N_3079,In_1738,In_2074);
nor U3080 (N_3080,In_1001,In_1587);
nand U3081 (N_3081,In_2329,In_553);
and U3082 (N_3082,In_338,In_1541);
or U3083 (N_3083,In_2276,In_500);
or U3084 (N_3084,In_1465,In_524);
nand U3085 (N_3085,In_2232,In_1929);
or U3086 (N_3086,In_1106,In_1229);
nor U3087 (N_3087,In_1983,In_874);
nand U3088 (N_3088,In_191,In_1054);
nand U3089 (N_3089,In_2480,In_1194);
nor U3090 (N_3090,In_1464,In_45);
nor U3091 (N_3091,In_464,In_579);
nand U3092 (N_3092,In_2003,In_2404);
nor U3093 (N_3093,In_1097,In_2412);
nor U3094 (N_3094,In_1153,In_2493);
nor U3095 (N_3095,In_35,In_867);
nor U3096 (N_3096,In_1502,In_2193);
xor U3097 (N_3097,In_1321,In_409);
nand U3098 (N_3098,In_1320,In_331);
nor U3099 (N_3099,In_1754,In_2159);
and U3100 (N_3100,In_1147,In_1418);
and U3101 (N_3101,In_1390,In_1015);
or U3102 (N_3102,In_2474,In_419);
nor U3103 (N_3103,In_518,In_2198);
nor U3104 (N_3104,In_19,In_1052);
nor U3105 (N_3105,In_1693,In_2442);
and U3106 (N_3106,In_1736,In_616);
xnor U3107 (N_3107,In_383,In_2244);
nand U3108 (N_3108,In_1924,In_1975);
nor U3109 (N_3109,In_1146,In_790);
or U3110 (N_3110,In_770,In_1001);
nor U3111 (N_3111,In_659,In_1329);
nor U3112 (N_3112,In_955,In_0);
nand U3113 (N_3113,In_962,In_950);
nand U3114 (N_3114,In_2209,In_1885);
and U3115 (N_3115,In_288,In_1389);
nand U3116 (N_3116,In_458,In_1385);
nand U3117 (N_3117,In_1003,In_134);
nand U3118 (N_3118,In_2126,In_618);
nor U3119 (N_3119,In_1124,In_2498);
or U3120 (N_3120,In_1806,In_2080);
nand U3121 (N_3121,In_1626,In_1637);
nand U3122 (N_3122,In_445,In_1654);
nor U3123 (N_3123,In_1893,In_2298);
nor U3124 (N_3124,In_934,In_1222);
xor U3125 (N_3125,N_1905,N_672);
nand U3126 (N_3126,N_1387,N_2549);
or U3127 (N_3127,N_767,N_1457);
or U3128 (N_3128,N_999,N_1100);
nand U3129 (N_3129,N_2292,N_2783);
nand U3130 (N_3130,N_1941,N_3031);
xor U3131 (N_3131,N_833,N_1324);
nor U3132 (N_3132,N_1462,N_2958);
or U3133 (N_3133,N_627,N_639);
xor U3134 (N_3134,N_2085,N_549);
xnor U3135 (N_3135,N_2172,N_1302);
and U3136 (N_3136,N_470,N_37);
nor U3137 (N_3137,N_682,N_1276);
nand U3138 (N_3138,N_2686,N_2241);
xnor U3139 (N_3139,N_468,N_2423);
nor U3140 (N_3140,N_2496,N_1374);
nand U3141 (N_3141,N_530,N_460);
and U3142 (N_3142,N_1014,N_663);
nor U3143 (N_3143,N_1416,N_2111);
xnor U3144 (N_3144,N_343,N_2823);
nor U3145 (N_3145,N_2690,N_1062);
nand U3146 (N_3146,N_567,N_818);
nand U3147 (N_3147,N_2953,N_2448);
and U3148 (N_3148,N_2112,N_730);
nand U3149 (N_3149,N_798,N_638);
nor U3150 (N_3150,N_2136,N_2158);
or U3151 (N_3151,N_2539,N_2135);
nand U3152 (N_3152,N_1344,N_1343);
nor U3153 (N_3153,N_1694,N_946);
and U3154 (N_3154,N_1898,N_1563);
and U3155 (N_3155,N_1669,N_2190);
and U3156 (N_3156,N_2796,N_1951);
nor U3157 (N_3157,N_2835,N_1974);
and U3158 (N_3158,N_1006,N_1066);
nor U3159 (N_3159,N_2705,N_1723);
or U3160 (N_3160,N_834,N_2692);
xor U3161 (N_3161,N_2729,N_1867);
xor U3162 (N_3162,N_2821,N_843);
nand U3163 (N_3163,N_413,N_1753);
nor U3164 (N_3164,N_386,N_1980);
and U3165 (N_3165,N_1902,N_1573);
nor U3166 (N_3166,N_2401,N_1703);
and U3167 (N_3167,N_1923,N_93);
nor U3168 (N_3168,N_1238,N_2664);
nand U3169 (N_3169,N_1284,N_1636);
nand U3170 (N_3170,N_254,N_2441);
and U3171 (N_3171,N_2340,N_2788);
and U3172 (N_3172,N_1068,N_1015);
nand U3173 (N_3173,N_3103,N_921);
nor U3174 (N_3174,N_2892,N_1056);
nand U3175 (N_3175,N_2765,N_2442);
and U3176 (N_3176,N_2063,N_1945);
nor U3177 (N_3177,N_1317,N_2597);
and U3178 (N_3178,N_1977,N_1787);
and U3179 (N_3179,N_891,N_1791);
and U3180 (N_3180,N_2894,N_744);
nor U3181 (N_3181,N_2504,N_2088);
nor U3182 (N_3182,N_2403,N_2255);
or U3183 (N_3183,N_2616,N_2097);
or U3184 (N_3184,N_2305,N_216);
or U3185 (N_3185,N_56,N_2507);
nor U3186 (N_3186,N_621,N_712);
nor U3187 (N_3187,N_2219,N_931);
nor U3188 (N_3188,N_560,N_1048);
and U3189 (N_3189,N_2643,N_2168);
or U3190 (N_3190,N_2907,N_3061);
and U3191 (N_3191,N_864,N_2060);
nor U3192 (N_3192,N_2931,N_2672);
nand U3193 (N_3193,N_1871,N_511);
nand U3194 (N_3194,N_2175,N_2527);
xnor U3195 (N_3195,N_1175,N_2189);
nand U3196 (N_3196,N_1551,N_561);
nor U3197 (N_3197,N_1866,N_2499);
nor U3198 (N_3198,N_1187,N_1390);
nor U3199 (N_3199,N_2809,N_581);
xor U3200 (N_3200,N_2472,N_570);
xor U3201 (N_3201,N_1389,N_1382);
nor U3202 (N_3202,N_3066,N_2843);
nor U3203 (N_3203,N_1385,N_708);
nand U3204 (N_3204,N_158,N_2486);
or U3205 (N_3205,N_134,N_2421);
nand U3206 (N_3206,N_1067,N_1953);
xnor U3207 (N_3207,N_1598,N_2460);
nand U3208 (N_3208,N_3123,N_1307);
or U3209 (N_3209,N_205,N_2346);
nor U3210 (N_3210,N_2438,N_3016);
or U3211 (N_3211,N_1111,N_1314);
or U3212 (N_3212,N_1201,N_1522);
xnor U3213 (N_3213,N_365,N_1113);
nor U3214 (N_3214,N_2627,N_1635);
and U3215 (N_3215,N_913,N_251);
nand U3216 (N_3216,N_1024,N_1439);
or U3217 (N_3217,N_2864,N_3018);
nor U3218 (N_3218,N_1252,N_2262);
nor U3219 (N_3219,N_2431,N_1400);
nand U3220 (N_3220,N_1095,N_2008);
nor U3221 (N_3221,N_903,N_2997);
xnor U3222 (N_3222,N_152,N_33);
or U3223 (N_3223,N_1286,N_2533);
and U3224 (N_3224,N_958,N_3118);
nand U3225 (N_3225,N_476,N_1486);
nor U3226 (N_3226,N_1948,N_1991);
nor U3227 (N_3227,N_2230,N_303);
or U3228 (N_3228,N_1641,N_1215);
and U3229 (N_3229,N_1299,N_139);
nor U3230 (N_3230,N_2167,N_2480);
nor U3231 (N_3231,N_574,N_2573);
nor U3232 (N_3232,N_2933,N_1608);
xnor U3233 (N_3233,N_424,N_1047);
nor U3234 (N_3234,N_25,N_778);
nand U3235 (N_3235,N_2681,N_284);
nand U3236 (N_3236,N_195,N_2270);
nand U3237 (N_3237,N_421,N_1291);
xor U3238 (N_3238,N_1101,N_1073);
and U3239 (N_3239,N_43,N_28);
xor U3240 (N_3240,N_1103,N_2444);
nand U3241 (N_3241,N_358,N_318);
or U3242 (N_3242,N_1338,N_1607);
nand U3243 (N_3243,N_1294,N_2591);
and U3244 (N_3244,N_990,N_836);
and U3245 (N_3245,N_2372,N_2861);
nand U3246 (N_3246,N_2583,N_1290);
and U3247 (N_3247,N_896,N_121);
nor U3248 (N_3248,N_670,N_746);
or U3249 (N_3249,N_2212,N_2083);
nor U3250 (N_3250,N_1449,N_2887);
or U3251 (N_3251,N_2736,N_1209);
and U3252 (N_3252,N_2826,N_2320);
nor U3253 (N_3253,N_1182,N_211);
xnor U3254 (N_3254,N_376,N_2016);
nand U3255 (N_3255,N_847,N_2091);
or U3256 (N_3256,N_1535,N_740);
and U3257 (N_3257,N_2181,N_1967);
or U3258 (N_3258,N_204,N_3027);
nor U3259 (N_3259,N_630,N_1473);
and U3260 (N_3260,N_1492,N_242);
nand U3261 (N_3261,N_1041,N_1506);
nand U3262 (N_3262,N_1196,N_1153);
or U3263 (N_3263,N_475,N_2704);
or U3264 (N_3264,N_2268,N_2081);
and U3265 (N_3265,N_1216,N_1203);
or U3266 (N_3266,N_295,N_1633);
or U3267 (N_3267,N_2179,N_2793);
or U3268 (N_3268,N_698,N_1002);
nor U3269 (N_3269,N_2165,N_2808);
nand U3270 (N_3270,N_846,N_2984);
or U3271 (N_3271,N_1807,N_1230);
nor U3272 (N_3272,N_2250,N_430);
nor U3273 (N_3273,N_1279,N_1982);
or U3274 (N_3274,N_2155,N_2059);
and U3275 (N_3275,N_917,N_1058);
nand U3276 (N_3276,N_1013,N_499);
nor U3277 (N_3277,N_1806,N_1225);
nand U3278 (N_3278,N_2824,N_2131);
nor U3279 (N_3279,N_2501,N_1192);
or U3280 (N_3280,N_2508,N_2767);
nor U3281 (N_3281,N_2598,N_354);
nor U3282 (N_3282,N_416,N_2866);
nand U3283 (N_3283,N_2578,N_861);
nor U3284 (N_3284,N_217,N_1186);
or U3285 (N_3285,N_2934,N_1969);
nand U3286 (N_3286,N_42,N_1232);
nand U3287 (N_3287,N_2411,N_1033);
nor U3288 (N_3288,N_918,N_2891);
nor U3289 (N_3289,N_2668,N_531);
or U3290 (N_3290,N_1701,N_2568);
or U3291 (N_3291,N_1968,N_940);
nand U3292 (N_3292,N_426,N_3072);
nand U3293 (N_3293,N_973,N_1571);
nor U3294 (N_3294,N_617,N_144);
or U3295 (N_3295,N_1149,N_200);
or U3296 (N_3296,N_3013,N_775);
xor U3297 (N_3297,N_369,N_1759);
and U3298 (N_3298,N_1285,N_327);
or U3299 (N_3299,N_856,N_2337);
or U3300 (N_3300,N_1763,N_2080);
or U3301 (N_3301,N_515,N_306);
or U3302 (N_3302,N_1964,N_1802);
nand U3303 (N_3303,N_232,N_206);
nor U3304 (N_3304,N_1083,N_540);
and U3305 (N_3305,N_664,N_1361);
nand U3306 (N_3306,N_502,N_1913);
and U3307 (N_3307,N_1767,N_736);
and U3308 (N_3308,N_768,N_881);
and U3309 (N_3309,N_1016,N_82);
nand U3310 (N_3310,N_6,N_3006);
or U3311 (N_3311,N_2939,N_2723);
or U3312 (N_3312,N_260,N_3001);
or U3313 (N_3313,N_427,N_745);
nor U3314 (N_3314,N_985,N_162);
nor U3315 (N_3315,N_113,N_2656);
and U3316 (N_3316,N_494,N_2970);
nor U3317 (N_3317,N_1538,N_1962);
nand U3318 (N_3318,N_1081,N_2755);
nand U3319 (N_3319,N_1444,N_874);
xnor U3320 (N_3320,N_399,N_2043);
or U3321 (N_3321,N_1834,N_1123);
xnor U3322 (N_3322,N_637,N_1638);
nand U3323 (N_3323,N_2127,N_3008);
nor U3324 (N_3324,N_2886,N_1292);
nand U3325 (N_3325,N_3068,N_2717);
xnor U3326 (N_3326,N_1342,N_2046);
nand U3327 (N_3327,N_2806,N_1243);
nand U3328 (N_3328,N_2235,N_2816);
or U3329 (N_3329,N_1340,N_1096);
or U3330 (N_3330,N_1861,N_693);
nand U3331 (N_3331,N_1679,N_2065);
and U3332 (N_3332,N_484,N_145);
or U3333 (N_3333,N_2464,N_207);
nor U3334 (N_3334,N_509,N_2074);
or U3335 (N_3335,N_1405,N_2474);
xor U3336 (N_3336,N_2555,N_474);
nand U3337 (N_3337,N_3025,N_583);
nor U3338 (N_3338,N_976,N_2126);
and U3339 (N_3339,N_347,N_904);
nor U3340 (N_3340,N_3073,N_220);
nand U3341 (N_3341,N_292,N_2195);
nand U3342 (N_3342,N_535,N_457);
or U3343 (N_3343,N_3036,N_2895);
xor U3344 (N_3344,N_1725,N_450);
or U3345 (N_3345,N_1553,N_1503);
nand U3346 (N_3346,N_3105,N_1424);
and U3347 (N_3347,N_2357,N_719);
nand U3348 (N_3348,N_2638,N_1370);
nand U3349 (N_3349,N_669,N_1729);
nand U3350 (N_3350,N_2014,N_2893);
or U3351 (N_3351,N_3117,N_2351);
or U3352 (N_3352,N_3059,N_490);
nor U3353 (N_3353,N_1334,N_2554);
or U3354 (N_3354,N_1689,N_3055);
nand U3355 (N_3355,N_1911,N_1784);
and U3356 (N_3356,N_289,N_1327);
or U3357 (N_3357,N_2106,N_3096);
nor U3358 (N_3358,N_3104,N_877);
nand U3359 (N_3359,N_704,N_2880);
xnor U3360 (N_3360,N_529,N_871);
and U3361 (N_3361,N_290,N_1137);
or U3362 (N_3362,N_594,N_2992);
and U3363 (N_3363,N_3044,N_1921);
nand U3364 (N_3364,N_1748,N_2450);
xnor U3365 (N_3365,N_1773,N_1580);
xor U3366 (N_3366,N_2951,N_1171);
and U3367 (N_3367,N_954,N_1337);
nor U3368 (N_3368,N_364,N_1749);
or U3369 (N_3369,N_1899,N_485);
or U3370 (N_3370,N_2682,N_1667);
or U3371 (N_3371,N_2354,N_1539);
nor U3372 (N_3372,N_2968,N_715);
nand U3373 (N_3373,N_1322,N_1975);
nor U3374 (N_3374,N_1960,N_71);
and U3375 (N_3375,N_2979,N_1581);
nor U3376 (N_3376,N_87,N_701);
nor U3377 (N_3377,N_462,N_451);
nor U3378 (N_3378,N_2304,N_2227);
and U3379 (N_3379,N_3020,N_374);
or U3380 (N_3380,N_47,N_3034);
nand U3381 (N_3381,N_2815,N_1534);
nor U3382 (N_3382,N_414,N_1010);
or U3383 (N_3383,N_1797,N_2698);
nand U3384 (N_3384,N_156,N_507);
nand U3385 (N_3385,N_1819,N_525);
nor U3386 (N_3386,N_1330,N_2244);
or U3387 (N_3387,N_3005,N_2528);
nor U3388 (N_3388,N_2201,N_1349);
xor U3389 (N_3389,N_2814,N_2021);
nor U3390 (N_3390,N_2999,N_1464);
nand U3391 (N_3391,N_1345,N_264);
or U3392 (N_3392,N_105,N_1606);
or U3393 (N_3393,N_2829,N_2276);
or U3394 (N_3394,N_900,N_588);
nand U3395 (N_3395,N_930,N_1843);
xnor U3396 (N_3396,N_2,N_130);
nor U3397 (N_3397,N_805,N_202);
nor U3398 (N_3398,N_679,N_2204);
nor U3399 (N_3399,N_1484,N_1611);
nand U3400 (N_3400,N_2224,N_2649);
nand U3401 (N_3401,N_756,N_1125);
nor U3402 (N_3402,N_2852,N_1386);
and U3403 (N_3403,N_458,N_2948);
nor U3404 (N_3404,N_1256,N_2322);
or U3405 (N_3405,N_294,N_366);
and U3406 (N_3406,N_991,N_1208);
and U3407 (N_3407,N_1637,N_645);
nor U3408 (N_3408,N_791,N_684);
or U3409 (N_3409,N_1161,N_2713);
and U3410 (N_3410,N_0,N_2130);
or U3411 (N_3411,N_677,N_2856);
and U3412 (N_3412,N_442,N_74);
or U3413 (N_3413,N_610,N_2696);
or U3414 (N_3414,N_1379,N_892);
and U3415 (N_3415,N_944,N_1779);
nor U3416 (N_3416,N_1297,N_1803);
xor U3417 (N_3417,N_1304,N_1001);
nand U3418 (N_3418,N_2994,N_982);
or U3419 (N_3419,N_2524,N_2567);
or U3420 (N_3420,N_67,N_398);
or U3421 (N_3421,N_1839,N_1778);
or U3422 (N_3422,N_1687,N_691);
xnor U3423 (N_3423,N_100,N_1102);
nand U3424 (N_3424,N_909,N_1875);
and U3425 (N_3425,N_852,N_1076);
or U3426 (N_3426,N_151,N_2150);
nand U3427 (N_3427,N_2327,N_1339);
and U3428 (N_3428,N_854,N_1454);
and U3429 (N_3429,N_397,N_1207);
nand U3430 (N_3430,N_2239,N_981);
and U3431 (N_3431,N_2885,N_497);
or U3432 (N_3432,N_1533,N_411);
or U3433 (N_3433,N_1904,N_2369);
xor U3434 (N_3434,N_2274,N_616);
nand U3435 (N_3435,N_920,N_2557);
or U3436 (N_3436,N_977,N_1954);
nor U3437 (N_3437,N_1670,N_1713);
nand U3438 (N_3438,N_456,N_2355);
nand U3439 (N_3439,N_1718,N_1381);
xnor U3440 (N_3440,N_826,N_3076);
and U3441 (N_3441,N_2537,N_3039);
nor U3442 (N_3442,N_1659,N_668);
nand U3443 (N_3443,N_2799,N_132);
xor U3444 (N_3444,N_59,N_1895);
and U3445 (N_3445,N_723,N_1907);
nand U3446 (N_3446,N_1318,N_1560);
or U3447 (N_3447,N_1532,N_3115);
or U3448 (N_3448,N_1512,N_1692);
nand U3449 (N_3449,N_2810,N_77);
nand U3450 (N_3450,N_2918,N_935);
or U3451 (N_3451,N_1764,N_1456);
nor U3452 (N_3452,N_1796,N_832);
or U3453 (N_3453,N_1654,N_964);
nand U3454 (N_3454,N_2173,N_2608);
nand U3455 (N_3455,N_1828,N_2670);
or U3456 (N_3456,N_76,N_2650);
or U3457 (N_3457,N_2912,N_461);
xor U3458 (N_3458,N_1422,N_573);
xor U3459 (N_3459,N_2641,N_705);
nand U3460 (N_3460,N_2914,N_875);
and U3461 (N_3461,N_131,N_1280);
or U3462 (N_3462,N_1399,N_2716);
nor U3463 (N_3463,N_248,N_2804);
and U3464 (N_3464,N_116,N_128);
nor U3465 (N_3465,N_2099,N_1086);
nor U3466 (N_3466,N_111,N_1568);
nand U3467 (N_3467,N_3060,N_3112);
nand U3468 (N_3468,N_3097,N_159);
nor U3469 (N_3469,N_1212,N_972);
and U3470 (N_3470,N_1179,N_2640);
xnor U3471 (N_3471,N_7,N_2881);
nand U3472 (N_3472,N_1917,N_766);
or U3473 (N_3473,N_1321,N_2915);
and U3474 (N_3474,N_2440,N_177);
nand U3475 (N_3475,N_1181,N_1910);
or U3476 (N_3476,N_2153,N_186);
or U3477 (N_3477,N_4,N_2802);
xnor U3478 (N_3478,N_1210,N_2217);
nor U3479 (N_3479,N_1946,N_1319);
nor U3480 (N_3480,N_1425,N_1218);
nand U3481 (N_3481,N_824,N_941);
or U3482 (N_3482,N_2922,N_2618);
or U3483 (N_3483,N_1929,N_269);
or U3484 (N_3484,N_929,N_422);
or U3485 (N_3485,N_1554,N_1599);
and U3486 (N_3486,N_1846,N_2837);
and U3487 (N_3487,N_2560,N_1265);
nor U3488 (N_3488,N_1621,N_1516);
or U3489 (N_3489,N_2581,N_2515);
xor U3490 (N_3490,N_2410,N_2770);
or U3491 (N_3491,N_356,N_368);
nor U3492 (N_3492,N_2620,N_2936);
or U3493 (N_3493,N_1524,N_1150);
and U3494 (N_3494,N_1949,N_2663);
and U3495 (N_3495,N_2742,N_2741);
nor U3496 (N_3496,N_3070,N_1341);
nor U3497 (N_3497,N_1720,N_2138);
or U3498 (N_3498,N_1766,N_2040);
nor U3499 (N_3499,N_2003,N_1859);
nand U3500 (N_3500,N_2781,N_974);
nor U3501 (N_3501,N_169,N_1305);
or U3502 (N_3502,N_2259,N_2558);
nand U3503 (N_3503,N_1359,N_2120);
nor U3504 (N_3504,N_170,N_245);
xnor U3505 (N_3505,N_2842,N_2542);
nor U3506 (N_3506,N_1590,N_1008);
and U3507 (N_3507,N_555,N_681);
and U3508 (N_3508,N_2456,N_819);
nor U3509 (N_3509,N_2971,N_1079);
nand U3510 (N_3510,N_2148,N_415);
nand U3511 (N_3511,N_1412,N_2418);
or U3512 (N_3512,N_2252,N_2865);
and U3513 (N_3513,N_1777,N_2694);
or U3514 (N_3514,N_2405,N_2812);
and U3515 (N_3515,N_1116,N_897);
or U3516 (N_3516,N_2853,N_2391);
or U3517 (N_3517,N_1675,N_3028);
nand U3518 (N_3518,N_2913,N_820);
and U3519 (N_3519,N_118,N_51);
and U3520 (N_3520,N_2037,N_815);
nand U3521 (N_3521,N_2392,N_1475);
nor U3522 (N_3522,N_3049,N_784);
or U3523 (N_3523,N_1589,N_2163);
nor U3524 (N_3524,N_781,N_1523);
or U3525 (N_3525,N_1393,N_2703);
or U3526 (N_3526,N_867,N_2169);
nor U3527 (N_3527,N_1690,N_890);
or U3528 (N_3528,N_3122,N_2813);
nor U3529 (N_3529,N_2273,N_198);
or U3530 (N_3530,N_2414,N_774);
nand U3531 (N_3531,N_1956,N_2595);
nor U3532 (N_3532,N_2209,N_432);
nand U3533 (N_3533,N_1624,N_94);
xnor U3534 (N_3534,N_1431,N_870);
or U3535 (N_3535,N_2141,N_2399);
nor U3536 (N_3536,N_2010,N_1548);
or U3537 (N_3537,N_2445,N_3109);
and U3538 (N_3538,N_439,N_138);
nor U3539 (N_3539,N_648,N_1817);
xor U3540 (N_3540,N_2094,N_1901);
nor U3541 (N_3541,N_2902,N_1021);
and U3542 (N_3542,N_2147,N_2950);
nor U3543 (N_3543,N_2345,N_2651);
xnor U3544 (N_3544,N_661,N_279);
nor U3545 (N_3545,N_1601,N_2774);
nor U3546 (N_3546,N_2429,N_1053);
nor U3547 (N_3547,N_665,N_271);
nor U3548 (N_3548,N_1430,N_3056);
and U3549 (N_3549,N_2706,N_1751);
xor U3550 (N_3550,N_2561,N_2031);
nand U3551 (N_3551,N_629,N_1813);
nand U3552 (N_3552,N_547,N_2188);
nand U3553 (N_3553,N_405,N_1501);
nor U3554 (N_3554,N_243,N_420);
nor U3555 (N_3555,N_1356,N_2875);
or U3556 (N_3556,N_1029,N_122);
nor U3557 (N_3557,N_2693,N_2437);
and U3558 (N_3558,N_2619,N_1529);
and U3559 (N_3559,N_1657,N_1891);
or U3560 (N_3560,N_1195,N_1678);
nor U3561 (N_3561,N_1268,N_2408);
or U3562 (N_3562,N_3009,N_1780);
nand U3563 (N_3563,N_1856,N_1310);
nand U3564 (N_3564,N_2100,N_1709);
nand U3565 (N_3565,N_987,N_607);
nor U3566 (N_3566,N_1760,N_687);
and U3567 (N_3567,N_2870,N_2174);
or U3568 (N_3568,N_700,N_2069);
nand U3569 (N_3569,N_1206,N_2500);
nor U3570 (N_3570,N_1189,N_579);
nor U3571 (N_3571,N_855,N_2301);
and U3572 (N_3572,N_2538,N_1556);
or U3573 (N_3573,N_1615,N_686);
nand U3574 (N_3574,N_208,N_1199);
nand U3575 (N_3575,N_656,N_3051);
nand U3576 (N_3576,N_319,N_526);
and U3577 (N_3577,N_2574,N_2653);
nand U3578 (N_3578,N_2458,N_2792);
or U3579 (N_3579,N_1362,N_384);
xnor U3580 (N_3580,N_2336,N_2628);
nor U3581 (N_3581,N_2848,N_1197);
nand U3582 (N_3582,N_2286,N_2535);
and U3583 (N_3583,N_1061,N_556);
nor U3584 (N_3584,N_647,N_1827);
xnor U3585 (N_3585,N_2733,N_886);
nor U3586 (N_3586,N_335,N_1744);
and U3587 (N_3587,N_1831,N_1401);
and U3588 (N_3588,N_680,N_2314);
and U3589 (N_3589,N_1629,N_2284);
or U3590 (N_3590,N_48,N_1887);
and U3591 (N_3591,N_2413,N_780);
and U3592 (N_3592,N_919,N_472);
or U3593 (N_3593,N_1620,N_1298);
xor U3594 (N_3594,N_235,N_57);
and U3595 (N_3595,N_1335,N_1578);
or U3596 (N_3596,N_2800,N_1998);
nor U3597 (N_3597,N_1158,N_1848);
or U3598 (N_3598,N_1639,N_2660);
nand U3599 (N_3599,N_2621,N_92);
and U3600 (N_3600,N_1747,N_240);
nand U3601 (N_3601,N_2859,N_1128);
or U3602 (N_3602,N_446,N_1202);
nand U3603 (N_3603,N_3,N_3022);
or U3604 (N_3604,N_2326,N_1732);
nand U3605 (N_3605,N_2047,N_2030);
or U3606 (N_3606,N_835,N_960);
nand U3607 (N_3607,N_710,N_965);
or U3608 (N_3608,N_651,N_1733);
and U3609 (N_3609,N_3000,N_626);
nand U3610 (N_3610,N_2778,N_258);
nor U3611 (N_3611,N_3041,N_2087);
and U3612 (N_3612,N_2009,N_1055);
nor U3613 (N_3613,N_695,N_1497);
xor U3614 (N_3614,N_2543,N_2226);
xnor U3615 (N_3615,N_589,N_2983);
nand U3616 (N_3616,N_38,N_1190);
xnor U3617 (N_3617,N_823,N_844);
nor U3618 (N_3618,N_699,N_1559);
nor U3619 (N_3619,N_595,N_1513);
nand U3620 (N_3620,N_1889,N_2697);
and U3621 (N_3621,N_326,N_2362);
nand U3622 (N_3622,N_2571,N_1287);
nor U3623 (N_3623,N_1549,N_389);
and U3624 (N_3624,N_157,N_21);
or U3625 (N_3625,N_2211,N_283);
nor U3626 (N_3626,N_1712,N_728);
or U3627 (N_3627,N_1377,N_1973);
or U3628 (N_3628,N_2991,N_148);
nor U3629 (N_3629,N_2665,N_2454);
and U3630 (N_3630,N_2750,N_436);
nor U3631 (N_3631,N_1163,N_716);
or U3632 (N_3632,N_2143,N_2465);
or U3633 (N_3633,N_2688,N_2605);
and U3634 (N_3634,N_2176,N_2722);
xor U3635 (N_3635,N_166,N_83);
nor U3636 (N_3636,N_1269,N_1574);
nor U3637 (N_3637,N_2109,N_1000);
and U3638 (N_3638,N_1826,N_239);
or U3639 (N_3639,N_532,N_392);
xor U3640 (N_3640,N_739,N_2115);
nor U3641 (N_3641,N_1541,N_2559);
and U3642 (N_3642,N_49,N_1936);
nand U3643 (N_3643,N_1035,N_905);
and U3644 (N_3644,N_720,N_2844);
or U3645 (N_3645,N_1445,N_1988);
xor U3646 (N_3646,N_2358,N_2961);
and U3647 (N_3647,N_1688,N_199);
nor U3648 (N_3648,N_1371,N_3082);
or U3649 (N_3649,N_1699,N_950);
nor U3650 (N_3650,N_73,N_1653);
nand U3651 (N_3651,N_2678,N_40);
or U3652 (N_3652,N_265,N_1728);
or U3653 (N_3653,N_1427,N_296);
nand U3654 (N_3654,N_2376,N_1138);
and U3655 (N_3655,N_582,N_14);
nor U3656 (N_3656,N_1063,N_278);
nand U3657 (N_3657,N_1612,N_816);
nor U3658 (N_3658,N_2280,N_1112);
nor U3659 (N_3659,N_2636,N_1972);
and U3660 (N_3660,N_809,N_2116);
nor U3661 (N_3661,N_1333,N_53);
nand U3662 (N_3662,N_1239,N_792);
nand U3663 (N_3663,N_1115,N_68);
nand U3664 (N_3664,N_2363,N_236);
nand U3665 (N_3665,N_2182,N_483);
and U3666 (N_3666,N_1418,N_2609);
nor U3667 (N_3667,N_2064,N_962);
and U3668 (N_3668,N_1562,N_1172);
or U3669 (N_3669,N_323,N_1697);
and U3670 (N_3670,N_2378,N_2124);
or U3671 (N_3671,N_2022,N_282);
xnor U3672 (N_3672,N_696,N_280);
nand U3673 (N_3673,N_2811,N_160);
nand U3674 (N_3674,N_1488,N_1680);
nand U3675 (N_3675,N_2348,N_1993);
nand U3676 (N_3676,N_123,N_3095);
xnor U3677 (N_3677,N_901,N_879);
or U3678 (N_3678,N_3040,N_2632);
or U3679 (N_3679,N_1658,N_2530);
xor U3680 (N_3680,N_2828,N_1525);
and U3681 (N_3681,N_153,N_653);
nand U3682 (N_3682,N_2954,N_759);
xor U3683 (N_3683,N_850,N_2002);
nor U3684 (N_3684,N_106,N_1261);
or U3685 (N_3685,N_657,N_2242);
nand U3686 (N_3686,N_1643,N_1544);
and U3687 (N_3687,N_1104,N_1300);
and U3688 (N_3688,N_60,N_523);
or U3689 (N_3689,N_2753,N_2884);
nand U3690 (N_3690,N_1278,N_787);
and U3691 (N_3691,N_109,N_1586);
nor U3692 (N_3692,N_2727,N_2714);
xor U3693 (N_3693,N_2025,N_1582);
and U3694 (N_3694,N_266,N_2385);
and U3695 (N_3695,N_2724,N_2617);
nand U3696 (N_3696,N_1626,N_142);
and U3697 (N_3697,N_2684,N_1419);
nand U3698 (N_3698,N_1110,N_1645);
and U3699 (N_3699,N_1518,N_110);
nor U3700 (N_3700,N_1815,N_1649);
or U3701 (N_3701,N_55,N_1080);
or U3702 (N_3702,N_1900,N_2596);
or U3703 (N_3703,N_1227,N_2001);
nand U3704 (N_3704,N_2566,N_1625);
nor U3705 (N_3705,N_98,N_3021);
nand U3706 (N_3706,N_2850,N_1436);
nor U3707 (N_3707,N_2956,N_2086);
xor U3708 (N_3708,N_26,N_622);
or U3709 (N_3709,N_1369,N_2927);
xnor U3710 (N_3710,N_328,N_2779);
xnor U3711 (N_3711,N_1691,N_1821);
nand U3712 (N_3712,N_2263,N_2290);
and U3713 (N_3713,N_1970,N_2726);
nand U3714 (N_3714,N_1027,N_2117);
nor U3715 (N_3715,N_625,N_2243);
nand U3716 (N_3716,N_259,N_602);
nor U3717 (N_3717,N_1622,N_2762);
or U3718 (N_3718,N_659,N_2387);
or U3719 (N_3719,N_2383,N_2349);
nand U3720 (N_3720,N_312,N_311);
nand U3721 (N_3721,N_1470,N_2103);
nand U3722 (N_3722,N_821,N_789);
nor U3723 (N_3723,N_1628,N_300);
nor U3724 (N_3724,N_1698,N_1438);
and U3725 (N_3725,N_1223,N_2073);
xnor U3726 (N_3726,N_3081,N_2334);
nor U3727 (N_3727,N_1485,N_1987);
and U3728 (N_3728,N_2271,N_1376);
and U3729 (N_3729,N_336,N_2093);
nor U3730 (N_3730,N_1451,N_1075);
or U3731 (N_3731,N_2154,N_1696);
or U3732 (N_3732,N_2166,N_1452);
nor U3733 (N_3733,N_3077,N_924);
xnor U3734 (N_3734,N_1157,N_1046);
nor U3735 (N_3735,N_1947,N_277);
nor U3736 (N_3736,N_1229,N_2308);
nor U3737 (N_3737,N_2098,N_183);
and U3738 (N_3738,N_2461,N_2180);
and U3739 (N_3739,N_1860,N_2398);
nand U3740 (N_3740,N_2102,N_1566);
nand U3741 (N_3741,N_2585,N_609);
nand U3742 (N_3742,N_2937,N_273);
nor U3743 (N_3743,N_3017,N_2592);
nand U3744 (N_3744,N_808,N_1458);
nor U3745 (N_3745,N_2580,N_2862);
nand U3746 (N_3746,N_3012,N_718);
and U3747 (N_3747,N_2514,N_888);
and U3748 (N_3748,N_1352,N_765);
nand U3749 (N_3749,N_1476,N_2552);
or U3750 (N_3750,N_752,N_1880);
or U3751 (N_3751,N_1648,N_760);
xnor U3752 (N_3752,N_1221,N_500);
nor U3753 (N_3753,N_2962,N_2790);
xor U3754 (N_3754,N_1833,N_1782);
nor U3755 (N_3755,N_2945,N_949);
nor U3756 (N_3756,N_2976,N_1937);
or U3757 (N_3757,N_1737,N_2677);
nor U3758 (N_3758,N_2921,N_2151);
or U3759 (N_3759,N_2562,N_914);
xnor U3760 (N_3760,N_2987,N_2447);
and U3761 (N_3761,N_911,N_2452);
nor U3762 (N_3762,N_321,N_2613);
or U3763 (N_3763,N_52,N_1521);
and U3764 (N_3764,N_1736,N_2860);
and U3765 (N_3765,N_2773,N_112);
nand U3766 (N_3766,N_3069,N_1668);
nor U3767 (N_3767,N_1384,N_732);
or U3768 (N_3768,N_2789,N_1986);
nand U3769 (N_3769,N_633,N_1990);
xnor U3770 (N_3770,N_2488,N_448);
or U3771 (N_3771,N_1237,N_1939);
xnor U3772 (N_3772,N_1303,N_1976);
nor U3773 (N_3773,N_224,N_810);
nor U3774 (N_3774,N_1402,N_741);
xor U3775 (N_3775,N_2134,N_2898);
nand U3776 (N_3776,N_2610,N_1994);
nor U3777 (N_3777,N_2475,N_2654);
and U3778 (N_3778,N_257,N_263);
and U3779 (N_3779,N_2161,N_674);
nand U3780 (N_3780,N_2746,N_1519);
xor U3781 (N_3781,N_333,N_3007);
nand U3782 (N_3782,N_1739,N_1312);
nor U3783 (N_3783,N_1672,N_382);
or U3784 (N_3784,N_2307,N_2666);
nand U3785 (N_3785,N_2359,N_937);
and U3786 (N_3786,N_2419,N_1919);
and U3787 (N_3787,N_883,N_2646);
or U3788 (N_3788,N_1037,N_943);
nor U3789 (N_3789,N_2377,N_261);
nand U3790 (N_3790,N_1575,N_2614);
nor U3791 (N_3791,N_2687,N_1801);
and U3792 (N_3792,N_2302,N_1007);
and U3793 (N_3793,N_58,N_2353);
nand U3794 (N_3794,N_2457,N_1442);
nand U3795 (N_3795,N_2890,N_599);
and U3796 (N_3796,N_2079,N_2089);
xor U3797 (N_3797,N_514,N_2960);
nor U3798 (N_3798,N_2295,N_334);
nor U3799 (N_3799,N_1489,N_1685);
nor U3800 (N_3800,N_898,N_683);
or U3801 (N_3801,N_1930,N_1034);
nand U3802 (N_3802,N_308,N_520);
nor U3803 (N_3803,N_2974,N_2162);
nor U3804 (N_3804,N_2647,N_2170);
and U3805 (N_3805,N_187,N_666);
nand U3806 (N_3806,N_769,N_992);
or U3807 (N_3807,N_959,N_1603);
nand U3808 (N_3808,N_2849,N_428);
or U3809 (N_3809,N_3083,N_3093);
nor U3810 (N_3810,N_1865,N_2888);
nor U3811 (N_3811,N_2751,N_2851);
nor U3812 (N_3812,N_2825,N_1557);
nand U3813 (N_3813,N_2026,N_1288);
nor U3814 (N_3814,N_41,N_2625);
and U3815 (N_3815,N_2076,N_471);
nand U3816 (N_3816,N_1446,N_611);
xnor U3817 (N_3817,N_390,N_3075);
or U3818 (N_3818,N_1478,N_1673);
nor U3819 (N_3819,N_803,N_2207);
xor U3820 (N_3820,N_2932,N_801);
nor U3821 (N_3821,N_2070,N_1325);
nand U3822 (N_3822,N_2801,N_2246);
nand U3823 (N_3823,N_1886,N_1135);
or U3824 (N_3824,N_1121,N_1091);
nor U3825 (N_3825,N_2240,N_673);
or U3826 (N_3826,N_1,N_1686);
nand U3827 (N_3827,N_1348,N_2525);
or U3828 (N_3828,N_2743,N_314);
or U3829 (N_3829,N_2468,N_1329);
and U3830 (N_3830,N_1864,N_1616);
nor U3831 (N_3831,N_1862,N_2487);
or U3832 (N_3832,N_2381,N_136);
nor U3833 (N_3833,N_1731,N_3004);
nor U3834 (N_3834,N_997,N_2142);
or U3835 (N_3835,N_449,N_868);
nor U3836 (N_3836,N_2764,N_619);
or U3837 (N_3837,N_1025,N_355);
xnor U3838 (N_3838,N_1248,N_2900);
and U3839 (N_3839,N_1408,N_750);
or U3840 (N_3840,N_2119,N_578);
nand U3841 (N_3841,N_2702,N_2210);
nor U3842 (N_3842,N_493,N_3085);
or U3843 (N_3843,N_800,N_1585);
and U3844 (N_3844,N_2634,N_2463);
and U3845 (N_3845,N_1714,N_1765);
and U3846 (N_3846,N_1719,N_1366);
or U3847 (N_3847,N_3078,N_1716);
nor U3848 (N_3848,N_2637,N_1162);
xnor U3849 (N_3849,N_85,N_2213);
nand U3850 (N_3850,N_1961,N_2310);
nand U3851 (N_3851,N_771,N_1108);
nand U3852 (N_3852,N_23,N_2061);
xnor U3853 (N_3853,N_988,N_2642);
and U3854 (N_3854,N_178,N_1674);
nor U3855 (N_3855,N_2629,N_3032);
xnor U3856 (N_3856,N_2004,N_1543);
nor U3857 (N_3857,N_1272,N_443);
and U3858 (N_3858,N_2333,N_827);
xnor U3859 (N_3859,N_1072,N_17);
nor U3860 (N_3860,N_614,N_1213);
nor U3861 (N_3861,N_894,N_1868);
or U3862 (N_3862,N_3033,N_851);
nor U3863 (N_3863,N_270,N_2516);
or U3864 (N_3864,N_2869,N_2685);
and U3865 (N_3865,N_1406,N_604);
or U3866 (N_3866,N_1498,N_412);
or U3867 (N_3867,N_2606,N_1051);
nand U3868 (N_3868,N_893,N_508);
xor U3869 (N_3869,N_858,N_214);
and U3870 (N_3870,N_2425,N_1705);
nand U3871 (N_3871,N_2989,N_1928);
nor U3872 (N_3872,N_2156,N_1769);
xnor U3873 (N_3873,N_880,N_887);
nor U3874 (N_3874,N_2267,N_1373);
nor U3875 (N_3875,N_2655,N_1005);
nand U3876 (N_3876,N_2517,N_1482);
nand U3877 (N_3877,N_1360,N_2101);
or U3878 (N_3878,N_302,N_124);
nand U3879 (N_3879,N_711,N_1060);
or U3880 (N_3880,N_2492,N_1109);
nand U3881 (N_3881,N_84,N_2144);
or U3882 (N_3882,N_101,N_304);
and U3883 (N_3883,N_2082,N_1480);
and U3884 (N_3884,N_2721,N_2066);
xor U3885 (N_3885,N_88,N_2588);
or U3886 (N_3886,N_3100,N_545);
and U3887 (N_3887,N_454,N_662);
and U3888 (N_3888,N_2459,N_2312);
nand U3889 (N_3889,N_1623,N_1959);
nor U3890 (N_3890,N_1935,N_753);
nor U3891 (N_3891,N_706,N_2745);
nand U3892 (N_3892,N_1942,N_2712);
or U3893 (N_3893,N_2797,N_378);
or U3894 (N_3894,N_1065,N_1440);
nor U3895 (N_3895,N_536,N_1089);
nand U3896 (N_3896,N_2965,N_2546);
and U3897 (N_3897,N_3101,N_348);
and U3898 (N_3898,N_1289,N_181);
and U3899 (N_3899,N_3099,N_1695);
nand U3900 (N_3900,N_1106,N_2897);
nor U3901 (N_3901,N_2365,N_1465);
and U3902 (N_3902,N_36,N_2433);
or U3903 (N_3903,N_2453,N_1471);
or U3904 (N_3904,N_1794,N_1903);
nand U3905 (N_3905,N_1433,N_510);
nor U3906 (N_3906,N_2041,N_876);
xnor U3907 (N_3907,N_2541,N_2187);
nor U3908 (N_3908,N_978,N_1052);
xor U3909 (N_3909,N_1879,N_2756);
or U3910 (N_3910,N_2318,N_2247);
and U3911 (N_3911,N_2957,N_1914);
nand U3912 (N_3912,N_30,N_936);
nor U3913 (N_3913,N_2878,N_1421);
nand U3914 (N_3914,N_2981,N_2324);
or U3915 (N_3915,N_603,N_2584);
and U3916 (N_3916,N_1447,N_1932);
nand U3917 (N_3917,N_1320,N_2128);
and U3918 (N_3918,N_218,N_1235);
nand U3919 (N_3919,N_1761,N_1650);
nand U3920 (N_3920,N_2123,N_1854);
xor U3921 (N_3921,N_623,N_1613);
nor U3922 (N_3922,N_301,N_2489);
or U3923 (N_3923,N_797,N_938);
nand U3924 (N_3924,N_63,N_1164);
or U3925 (N_3925,N_632,N_1681);
nand U3926 (N_3926,N_2969,N_1461);
xnor U3927 (N_3927,N_1789,N_297);
and U3928 (N_3928,N_409,N_2389);
nand U3929 (N_3929,N_994,N_505);
and U3930 (N_3930,N_2872,N_963);
nor U3931 (N_3931,N_1874,N_822);
and U3932 (N_3932,N_1129,N_857);
and U3933 (N_3933,N_2035,N_783);
or U3934 (N_3934,N_807,N_1140);
nor U3935 (N_3935,N_926,N_2281);
and U3936 (N_3936,N_2200,N_1792);
nand U3937 (N_3937,N_675,N_2840);
nor U3938 (N_3938,N_3003,N_1323);
or U3939 (N_3939,N_3089,N_165);
nor U3940 (N_3940,N_115,N_2012);
nand U3941 (N_3941,N_1336,N_91);
nor U3942 (N_3942,N_2502,N_1222);
nand U3943 (N_3943,N_2661,N_2577);
or U3944 (N_3944,N_908,N_1564);
nand U3945 (N_3945,N_1814,N_2737);
nor U3946 (N_3946,N_2972,N_2422);
nor U3947 (N_3947,N_1798,N_1592);
nand U3948 (N_3948,N_1200,N_975);
and U3949 (N_3949,N_188,N_506);
nand U3950 (N_3950,N_1144,N_2771);
xor U3951 (N_3951,N_2140,N_1277);
nor U3952 (N_3952,N_2332,N_1133);
nand U3953 (N_3953,N_1398,N_853);
or U3954 (N_3954,N_2803,N_431);
xor U3955 (N_3955,N_2473,N_2973);
and U3956 (N_3956,N_2947,N_213);
and U3957 (N_3957,N_1550,N_1240);
nand U3958 (N_3958,N_2739,N_814);
xor U3959 (N_3959,N_1511,N_717);
nor U3960 (N_3960,N_1985,N_2044);
and U3961 (N_3961,N_2402,N_606);
or U3962 (N_3962,N_1165,N_1070);
nor U3963 (N_3963,N_1676,N_313);
or U3964 (N_3964,N_518,N_1453);
and U3965 (N_3965,N_3079,N_1250);
nand U3966 (N_3966,N_2747,N_2145);
nor U3967 (N_3967,N_2446,N_1849);
and U3968 (N_3968,N_2191,N_2734);
xnor U3969 (N_3969,N_1594,N_1166);
and U3970 (N_3970,N_2725,N_189);
or U3971 (N_3971,N_272,N_425);
nor U3972 (N_3972,N_230,N_3014);
or U3973 (N_3973,N_2034,N_2194);
nor U3974 (N_3974,N_2356,N_848);
and U3975 (N_3975,N_2294,N_2768);
or U3976 (N_3976,N_1479,N_2786);
nor U3977 (N_3977,N_1122,N_2769);
or U3978 (N_3978,N_1394,N_2223);
or U3979 (N_3979,N_554,N_1126);
or U3980 (N_3980,N_2586,N_1906);
xnor U3981 (N_3981,N_1472,N_624);
nor U3982 (N_3982,N_1403,N_396);
or U3983 (N_3983,N_2260,N_2415);
and U3984 (N_3984,N_1118,N_1282);
and U3985 (N_3985,N_2700,N_1825);
nand U3986 (N_3986,N_1829,N_1087);
nand U3987 (N_3987,N_1364,N_168);
nand U3988 (N_3988,N_2096,N_496);
nor U3989 (N_3989,N_176,N_869);
and U3990 (N_3990,N_2171,N_380);
nor U3991 (N_3991,N_1558,N_50);
nand U3992 (N_3992,N_782,N_2715);
xor U3993 (N_3993,N_1742,N_1308);
nor U3994 (N_3994,N_2510,N_175);
nand U3995 (N_3995,N_2285,N_65);
nand U3996 (N_3996,N_2277,N_2113);
nor U3997 (N_3997,N_482,N_3050);
or U3998 (N_3998,N_2491,N_226);
or U3999 (N_3999,N_542,N_2794);
nor U4000 (N_4000,N_66,N_276);
and U4001 (N_4001,N_2234,N_947);
or U4002 (N_4002,N_1940,N_2784);
nor U4003 (N_4003,N_2582,N_480);
and U4004 (N_4004,N_2400,N_2090);
nor U4005 (N_4005,N_192,N_299);
xnor U4006 (N_4006,N_1170,N_146);
xnor U4007 (N_4007,N_1855,N_546);
nor U4008 (N_4008,N_360,N_2671);
or U4009 (N_4009,N_370,N_3023);
or U4010 (N_4010,N_2820,N_1781);
nand U4011 (N_4011,N_2478,N_2795);
or U4012 (N_4012,N_1735,N_2523);
and U4013 (N_4013,N_2269,N_1042);
nand U4014 (N_4014,N_114,N_2048);
nor U4015 (N_4015,N_1642,N_1786);
or U4016 (N_4016,N_631,N_2328);
nand U4017 (N_4017,N_1411,N_2910);
nor U4018 (N_4018,N_2760,N_1840);
and U4019 (N_4019,N_1837,N_2321);
nand U4020 (N_4020,N_13,N_605);
and U4021 (N_4021,N_634,N_2785);
nor U4022 (N_4022,N_2020,N_2291);
xor U4023 (N_4023,N_307,N_481);
or U4024 (N_4024,N_400,N_285);
nor U4025 (N_4025,N_2303,N_126);
xnor U4026 (N_4026,N_2718,N_394);
nand U4027 (N_4027,N_11,N_80);
nand U4028 (N_4028,N_2652,N_2225);
nor U4029 (N_4029,N_3067,N_2758);
nor U4030 (N_4030,N_1741,N_2908);
nand U4031 (N_4031,N_488,N_1178);
nor U4032 (N_4032,N_863,N_2575);
or U4033 (N_4033,N_469,N_512);
nand U4034 (N_4034,N_2522,N_1809);
nand U4035 (N_4035,N_1893,N_1916);
nand U4036 (N_4036,N_367,N_1293);
and U4037 (N_4037,N_1605,N_1414);
nand U4038 (N_4038,N_423,N_1168);
nand U4039 (N_4039,N_381,N_1727);
nand U4040 (N_4040,N_2709,N_1365);
and U4041 (N_4041,N_1395,N_2635);
nor U4042 (N_4042,N_828,N_517);
nor U4043 (N_4043,N_2874,N_1019);
nor U4044 (N_4044,N_129,N_1684);
and U4045 (N_4045,N_2680,N_3080);
and U4046 (N_4046,N_957,N_346);
nand U4047 (N_4047,N_1857,N_2338);
and U4048 (N_4048,N_2384,N_1026);
nand U4049 (N_4049,N_2645,N_2838);
and U4050 (N_4050,N_983,N_2108);
or U4051 (N_4051,N_246,N_2467);
and U4052 (N_4052,N_1838,N_2896);
or U4053 (N_4053,N_1306,N_1528);
and U4054 (N_4054,N_1254,N_221);
nand U4055 (N_4055,N_1413,N_534);
or U4056 (N_4056,N_137,N_1872);
nand U4057 (N_4057,N_572,N_330);
and U4058 (N_4058,N_1296,N_383);
nor U4059 (N_4059,N_54,N_2393);
nand U4060 (N_4060,N_902,N_1758);
nand U4061 (N_4061,N_1579,N_78);
or U4062 (N_4062,N_1824,N_179);
or U4063 (N_4063,N_2350,N_1094);
xnor U4064 (N_4064,N_979,N_906);
nor U4065 (N_4065,N_1788,N_417);
and U4066 (N_4066,N_2374,N_1388);
or U4067 (N_4067,N_252,N_3106);
or U4068 (N_4068,N_2479,N_799);
or U4069 (N_4069,N_3110,N_2599);
and U4070 (N_4070,N_2509,N_440);
or U4071 (N_4071,N_2352,N_1925);
or U4072 (N_4072,N_1708,N_2245);
and U4073 (N_4073,N_107,N_2624);
xor U4074 (N_4074,N_1820,N_3024);
nor U4075 (N_4075,N_1823,N_702);
and U4076 (N_4076,N_184,N_751);
nor U4077 (N_4077,N_377,N_1432);
and U4078 (N_4078,N_2287,N_418);
or U4079 (N_4079,N_338,N_2503);
nand U4080 (N_4080,N_349,N_2611);
nor U4081 (N_4081,N_1927,N_1743);
nand U4082 (N_4082,N_2323,N_120);
and U4083 (N_4083,N_1818,N_1666);
or U4084 (N_4084,N_1555,N_62);
or U4085 (N_4085,N_2042,N_628);
nand U4086 (N_4086,N_654,N_2300);
or U4087 (N_4087,N_197,N_402);
and U4088 (N_4088,N_845,N_3116);
or U4089 (N_4089,N_1469,N_2521);
and U4090 (N_4090,N_3102,N_1570);
or U4091 (N_4091,N_2231,N_363);
and U4092 (N_4092,N_250,N_2899);
xor U4093 (N_4093,N_2926,N_453);
nand U4094 (N_4094,N_817,N_1090);
or U4095 (N_4095,N_1944,N_2253);
and U4096 (N_4096,N_690,N_794);
nand U4097 (N_4097,N_1346,N_2133);
and U4098 (N_4098,N_433,N_1591);
nor U4099 (N_4099,N_215,N_2317);
xnor U4100 (N_4100,N_2434,N_247);
and U4101 (N_4101,N_2550,N_3038);
nand U4102 (N_4102,N_636,N_2335);
nor U4103 (N_4103,N_2995,N_2763);
nand U4104 (N_4104,N_234,N_1214);
nand U4105 (N_4105,N_2553,N_1883);
nand U4106 (N_4106,N_2289,N_644);
nand U4107 (N_4107,N_2867,N_2924);
xnor U4108 (N_4108,N_344,N_3062);
xnor U4109 (N_4109,N_1631,N_1409);
nand U4110 (N_4110,N_2053,N_1313);
xor U4111 (N_4111,N_371,N_967);
or U4112 (N_4112,N_655,N_1311);
or U4113 (N_4113,N_615,N_1142);
and U4114 (N_4114,N_1152,N_46);
and U4115 (N_4115,N_2279,N_44);
nand U4116 (N_4116,N_1030,N_2299);
or U4117 (N_4117,N_1380,N_445);
nand U4118 (N_4118,N_2761,N_2551);
xnor U4119 (N_4119,N_785,N_2701);
nand U4120 (N_4120,N_2033,N_489);
and U4121 (N_4121,N_1757,N_2909);
and U4122 (N_4122,N_1176,N_180);
nand U4123 (N_4123,N_1147,N_2249);
nand U4124 (N_4124,N_20,N_18);
nor U4125 (N_4125,N_22,N_1738);
nor U4126 (N_4126,N_196,N_2205);
nand U4127 (N_4127,N_1074,N_1315);
nand U4128 (N_4128,N_652,N_2361);
xnor U4129 (N_4129,N_1092,N_2316);
and U4130 (N_4130,N_640,N_1234);
and U4131 (N_4131,N_1527,N_1466);
nor U4132 (N_4132,N_737,N_1114);
nor U4133 (N_4133,N_1193,N_558);
and U4134 (N_4134,N_1491,N_2451);
and U4135 (N_4135,N_642,N_293);
and U4136 (N_4136,N_1177,N_1131);
and U4137 (N_4137,N_2938,N_2529);
xnor U4138 (N_4138,N_1915,N_1448);
nand U4139 (N_4139,N_3092,N_2506);
nor U4140 (N_4140,N_1540,N_726);
and U4141 (N_4141,N_571,N_61);
nor U4142 (N_4142,N_993,N_928);
or U4143 (N_4143,N_1264,N_587);
xnor U4144 (N_4144,N_1044,N_2237);
xnor U4145 (N_4145,N_1266,N_968);
nand U4146 (N_4146,N_2738,N_1220);
and U4147 (N_4147,N_2710,N_1211);
nand U4148 (N_4148,N_2942,N_2719);
xor U4149 (N_4149,N_3048,N_2772);
nand U4150 (N_4150,N_1542,N_5);
xnor U4151 (N_4151,N_2007,N_2594);
or U4152 (N_4152,N_2548,N_1355);
or U4153 (N_4153,N_1926,N_694);
or U4154 (N_4154,N_125,N_274);
nand U4155 (N_4155,N_1159,N_566);
and U4156 (N_4156,N_1064,N_1136);
nor U4157 (N_4157,N_667,N_1124);
nor U4158 (N_4158,N_1517,N_2845);
and U4159 (N_4159,N_2490,N_1955);
nand U4160 (N_4160,N_1271,N_3029);
nor U4161 (N_4161,N_1878,N_2056);
nor U4162 (N_4162,N_1351,N_231);
and U4163 (N_4163,N_2185,N_2282);
or U4164 (N_4164,N_2214,N_2373);
or U4165 (N_4165,N_34,N_3084);
nor U4166 (N_4166,N_434,N_1146);
nand U4167 (N_4167,N_329,N_291);
nor U4168 (N_4168,N_1995,N_459);
nand U4169 (N_4169,N_763,N_2390);
xnor U4170 (N_4170,N_676,N_2905);
or U4171 (N_4171,N_1281,N_2977);
nor U4172 (N_4172,N_2417,N_403);
and U4173 (N_4173,N_2344,N_393);
and U4174 (N_4174,N_2184,N_406);
or U4175 (N_4175,N_770,N_1774);
xor U4176 (N_4176,N_1258,N_1888);
or U4177 (N_4177,N_734,N_2602);
nand U4178 (N_4178,N_1184,N_559);
or U4179 (N_4179,N_1255,N_1347);
nor U4180 (N_4180,N_1706,N_1226);
nor U4181 (N_4181,N_2364,N_1107);
and U4182 (N_4182,N_16,N_703);
nand U4183 (N_4183,N_298,N_544);
xnor U4184 (N_4184,N_167,N_2615);
and U4185 (N_4185,N_150,N_2857);
and U4186 (N_4186,N_1530,N_724);
nand U4187 (N_4187,N_473,N_1850);
nand U4188 (N_4188,N_89,N_1017);
nand U4189 (N_4189,N_1350,N_1309);
or U4190 (N_4190,N_539,N_1704);
nor U4191 (N_4191,N_1429,N_952);
nand U4192 (N_4192,N_1804,N_455);
nand U4193 (N_4193,N_463,N_2325);
nand U4194 (N_4194,N_1617,N_2946);
or U4195 (N_4195,N_1963,N_1500);
or U4196 (N_4196,N_2683,N_600);
and U4197 (N_4197,N_2218,N_2832);
or U4198 (N_4198,N_2375,N_2028);
nor U4199 (N_4199,N_796,N_649);
or U4200 (N_4200,N_2511,N_2505);
nor U4201 (N_4201,N_2107,N_2980);
and U4202 (N_4202,N_149,N_1671);
or U4203 (N_4203,N_825,N_161);
and U4204 (N_4204,N_2265,N_320);
nand U4205 (N_4205,N_2493,N_689);
nand U4206 (N_4206,N_1151,N_2360);
nand U4207 (N_4207,N_580,N_8);
nor U4208 (N_4208,N_1577,N_1597);
and U4209 (N_4209,N_2068,N_2426);
nor U4210 (N_4210,N_268,N_477);
and U4211 (N_4211,N_2476,N_491);
and U4212 (N_4212,N_504,N_980);
xor U4213 (N_4213,N_2626,N_872);
nand U4214 (N_4214,N_793,N_961);
nand U4215 (N_4215,N_743,N_2222);
xor U4216 (N_4216,N_2339,N_2943);
nor U4217 (N_4217,N_340,N_64);
nand U4218 (N_4218,N_1423,N_806);
and U4219 (N_4219,N_3088,N_2644);
and U4220 (N_4220,N_650,N_2062);
nor U4221 (N_4221,N_1032,N_2371);
nand U4222 (N_4222,N_533,N_2532);
nor U4223 (N_4223,N_1331,N_2871);
nand U4224 (N_4224,N_1145,N_1841);
nor U4225 (N_4225,N_2545,N_884);
and U4226 (N_4226,N_951,N_2331);
xnor U4227 (N_4227,N_1020,N_2579);
or U4228 (N_4228,N_1918,N_2967);
nor U4229 (N_4229,N_447,N_345);
nor U4230 (N_4230,N_10,N_564);
nor U4231 (N_4231,N_1664,N_2673);
and U4232 (N_4232,N_286,N_2963);
xor U4233 (N_4233,N_1853,N_1922);
or U4234 (N_4234,N_970,N_209);
nand U4235 (N_4235,N_212,N_316);
or U4236 (N_4236,N_692,N_2587);
nand U4237 (N_4237,N_1397,N_2855);
nor U4238 (N_4238,N_788,N_2600);
nor U4239 (N_4239,N_590,N_839);
nand U4240 (N_4240,N_524,N_1455);
nor U4241 (N_4241,N_1830,N_3043);
xnor U4242 (N_4242,N_305,N_1909);
and U4243 (N_4243,N_1652,N_795);
nor U4244 (N_4244,N_373,N_671);
xnor U4245 (N_4245,N_410,N_2978);
nand U4246 (N_4246,N_2822,N_2038);
nand U4247 (N_4247,N_1367,N_2341);
nand U4248 (N_4248,N_2203,N_1054);
or U4249 (N_4249,N_1627,N_1651);
nand U4250 (N_4250,N_2298,N_1217);
nor U4251 (N_4251,N_408,N_2482);
or U4252 (N_4252,N_1614,N_467);
or U4253 (N_4253,N_2833,N_361);
or U4254 (N_4254,N_2313,N_2854);
or U4255 (N_4255,N_1410,N_2216);
nand U4256 (N_4256,N_777,N_1526);
and U4257 (N_4257,N_1800,N_966);
or U4258 (N_4258,N_1567,N_1082);
nor U4259 (N_4259,N_915,N_1039);
or U4260 (N_4260,N_1383,N_1180);
nor U4261 (N_4261,N_1022,N_1957);
or U4262 (N_4262,N_1632,N_2911);
nor U4263 (N_4263,N_729,N_81);
nor U4264 (N_4264,N_838,N_754);
nor U4265 (N_4265,N_2254,N_1700);
and U4266 (N_4266,N_1934,N_1011);
nor U4267 (N_4267,N_1565,N_738);
xnor U4268 (N_4268,N_1481,N_2759);
nand U4269 (N_4269,N_709,N_194);
and U4270 (N_4270,N_164,N_1085);
nand U4271 (N_4271,N_721,N_2805);
xnor U4272 (N_4272,N_3011,N_932);
and U4273 (N_4273,N_1069,N_1253);
nor U4274 (N_4274,N_776,N_1609);
nor U4275 (N_4275,N_1630,N_108);
and U4276 (N_4276,N_2232,N_1012);
and U4277 (N_4277,N_102,N_238);
nor U4278 (N_4278,N_747,N_1505);
or U4279 (N_4279,N_315,N_437);
or U4280 (N_4280,N_2757,N_538);
nand U4281 (N_4281,N_3052,N_1656);
and U4282 (N_4282,N_643,N_563);
and U4283 (N_4283,N_3064,N_2847);
xor U4284 (N_4284,N_2569,N_141);
and U4285 (N_4285,N_2197,N_228);
xnor U4286 (N_4286,N_2024,N_748);
and U4287 (N_4287,N_2982,N_591);
or U4288 (N_4288,N_1604,N_1191);
nand U4289 (N_4289,N_1795,N_466);
and U4290 (N_4290,N_2306,N_1257);
nand U4291 (N_4291,N_2483,N_757);
nor U4292 (N_4292,N_2777,N_1785);
and U4293 (N_4293,N_2157,N_550);
and U4294 (N_4294,N_2975,N_163);
nand U4295 (N_4295,N_2728,N_395);
nand U4296 (N_4296,N_3037,N_733);
and U4297 (N_4297,N_288,N_2397);
nand U4298 (N_4298,N_1241,N_948);
or U4299 (N_4299,N_1882,N_1971);
or U4300 (N_4300,N_3010,N_1045);
nor U4301 (N_4301,N_2818,N_912);
nand U4302 (N_4302,N_764,N_1682);
nand U4303 (N_4303,N_12,N_2831);
nor U4304 (N_4304,N_2368,N_1508);
and U4305 (N_4305,N_1105,N_1148);
and U4306 (N_4306,N_1663,N_3107);
or U4307 (N_4307,N_1835,N_2966);
and U4308 (N_4308,N_1375,N_2988);
and U4309 (N_4309,N_934,N_501);
or U4310 (N_4310,N_2283,N_1894);
nand U4311 (N_4311,N_1845,N_790);
nor U4312 (N_4312,N_2699,N_2462);
nor U4313 (N_4313,N_2744,N_2986);
or U4314 (N_4314,N_2051,N_618);
or U4315 (N_4315,N_1487,N_2477);
or U4316 (N_4316,N_2072,N_1897);
and U4317 (N_4317,N_29,N_3111);
or U4318 (N_4318,N_387,N_1117);
and U4319 (N_4319,N_1808,N_241);
or U4320 (N_4320,N_1173,N_2612);
nor U4321 (N_4321,N_953,N_557);
or U4322 (N_4322,N_2882,N_1477);
nor U4323 (N_4323,N_3046,N_1520);
or U4324 (N_4324,N_804,N_70);
or U4325 (N_4325,N_2045,N_1873);
and U4326 (N_4326,N_2215,N_2730);
nand U4327 (N_4327,N_1301,N_2556);
or U4328 (N_4328,N_331,N_1434);
and U4329 (N_4329,N_3054,N_2689);
nand U4330 (N_4330,N_731,N_2104);
xnor U4331 (N_4331,N_1920,N_1536);
nand U4332 (N_4332,N_2432,N_2424);
or U4333 (N_4333,N_1965,N_2928);
nand U4334 (N_4334,N_2749,N_24);
nand U4335 (N_4335,N_2122,N_1665);
and U4336 (N_4336,N_758,N_1130);
or U4337 (N_4337,N_762,N_2466);
or U4338 (N_4338,N_1584,N_2382);
nor U4339 (N_4339,N_1463,N_2676);
nor U4340 (N_4340,N_2817,N_841);
or U4341 (N_4341,N_2780,N_2208);
nand U4342 (N_4342,N_1099,N_147);
nand U4343 (N_4343,N_2075,N_830);
nor U4344 (N_4344,N_1372,N_31);
nor U4345 (N_4345,N_1499,N_3035);
nor U4346 (N_4346,N_3042,N_19);
nor U4347 (N_4347,N_2563,N_2748);
xor U4348 (N_4348,N_375,N_1141);
xor U4349 (N_4349,N_1246,N_3094);
or U4350 (N_4350,N_749,N_1999);
and U4351 (N_4351,N_2540,N_2311);
or U4352 (N_4352,N_1793,N_522);
nor U4353 (N_4353,N_813,N_281);
or U4354 (N_4354,N_487,N_1618);
and U4355 (N_4355,N_2050,N_79);
or U4356 (N_4356,N_3108,N_2152);
nor U4357 (N_4357,N_2006,N_1474);
or U4358 (N_4358,N_1494,N_849);
nor U4359 (N_4359,N_956,N_593);
or U4360 (N_4360,N_3124,N_2416);
or U4361 (N_4361,N_1468,N_2428);
xnor U4362 (N_4362,N_255,N_2873);
nor U4363 (N_4363,N_256,N_1049);
and U4364 (N_4364,N_2435,N_2386);
xnor U4365 (N_4365,N_1710,N_2409);
nor U4366 (N_4366,N_1989,N_1154);
nor U4367 (N_4367,N_75,N_2343);
xnor U4368 (N_4368,N_317,N_2940);
nand U4369 (N_4369,N_2054,N_1852);
nor U4370 (N_4370,N_1693,N_1028);
nand U4371 (N_4371,N_2512,N_543);
xnor U4372 (N_4372,N_1707,N_2039);
and U4373 (N_4373,N_154,N_1031);
xnor U4374 (N_4374,N_899,N_2930);
nand U4375 (N_4375,N_608,N_492);
or U4376 (N_4376,N_1702,N_310);
xor U4377 (N_4377,N_2648,N_1260);
xor U4378 (N_4378,N_1870,N_2593);
or U4379 (N_4379,N_597,N_2766);
and U4380 (N_4380,N_2484,N_2278);
nor U4381 (N_4381,N_2055,N_1391);
nor U4382 (N_4382,N_219,N_773);
and U4383 (N_4383,N_1504,N_1952);
nor U4384 (N_4384,N_2667,N_2944);
and U4385 (N_4385,N_3091,N_1205);
and U4386 (N_4386,N_287,N_1043);
nor U4387 (N_4387,N_1332,N_3002);
or U4388 (N_4388,N_513,N_562);
nor U4389 (N_4389,N_2836,N_586);
nor U4390 (N_4390,N_2164,N_2220);
nor U4391 (N_4391,N_2221,N_925);
or U4392 (N_4392,N_32,N_1224);
and U4393 (N_4393,N_2105,N_601);
or U4394 (N_4394,N_859,N_1851);
nand U4395 (N_4395,N_97,N_986);
and U4396 (N_4396,N_1502,N_90);
nor U4397 (N_4397,N_193,N_1139);
or U4398 (N_4398,N_516,N_1933);
or U4399 (N_4399,N_2005,N_1495);
nand U4400 (N_4400,N_984,N_2330);
and U4401 (N_4401,N_707,N_45);
and U4402 (N_4402,N_1437,N_2659);
nor U4403 (N_4403,N_351,N_1537);
and U4404 (N_4404,N_1392,N_401);
nand U4405 (N_4405,N_2993,N_727);
or U4406 (N_4406,N_2883,N_2903);
xor U4407 (N_4407,N_1596,N_249);
nand U4408 (N_4408,N_103,N_2146);
nor U4409 (N_4409,N_2470,N_2266);
nand U4410 (N_4410,N_1435,N_761);
or U4411 (N_4411,N_2901,N_1247);
nand U4412 (N_4412,N_2544,N_2439);
nor U4413 (N_4413,N_140,N_565);
xnor U4414 (N_4414,N_3121,N_1745);
and U4415 (N_4415,N_1228,N_2394);
nand U4416 (N_4416,N_568,N_171);
or U4417 (N_4417,N_1812,N_1004);
nor U4418 (N_4418,N_3063,N_2572);
nand U4419 (N_4419,N_464,N_2819);
or U4420 (N_4420,N_407,N_1531);
and U4421 (N_4421,N_1884,N_860);
nor U4422 (N_4422,N_385,N_2919);
or U4423 (N_4423,N_873,N_2296);
or U4424 (N_4424,N_86,N_1924);
nand U4425 (N_4425,N_2469,N_227);
and U4426 (N_4426,N_862,N_127);
xnor U4427 (N_4427,N_2633,N_971);
nor U4428 (N_4428,N_2846,N_2084);
nand U4429 (N_4429,N_1003,N_2834);
and U4430 (N_4430,N_478,N_528);
nand U4431 (N_4431,N_3087,N_1450);
and U4432 (N_4432,N_3114,N_725);
nand U4433 (N_4433,N_2202,N_922);
nor U4434 (N_4434,N_1634,N_2827);
or U4435 (N_4435,N_1490,N_1167);
xnor U4436 (N_4436,N_2430,N_1507);
or U4437 (N_4437,N_1711,N_866);
or U4438 (N_4438,N_1583,N_1983);
and U4439 (N_4439,N_2679,N_2121);
nand U4440 (N_4440,N_9,N_2513);
nand U4441 (N_4441,N_945,N_1244);
nor U4442 (N_4442,N_2078,N_104);
or U4443 (N_4443,N_840,N_1885);
xor U4444 (N_4444,N_135,N_592);
or U4445 (N_4445,N_223,N_2455);
nand U4446 (N_4446,N_527,N_2708);
nor U4447 (N_4447,N_379,N_1077);
and U4448 (N_4448,N_2603,N_2256);
or U4449 (N_4449,N_1127,N_253);
nor U4450 (N_4450,N_1847,N_1561);
nor U4451 (N_4451,N_541,N_35);
or U4452 (N_4452,N_1647,N_2029);
or U4453 (N_4453,N_2192,N_596);
or U4454 (N_4454,N_1892,N_1134);
nor U4455 (N_4455,N_2139,N_2735);
nor U4456 (N_4456,N_2998,N_2449);
and U4457 (N_4457,N_1510,N_1771);
nor U4458 (N_4458,N_1943,N_3090);
xnor U4459 (N_4459,N_1776,N_2067);
or U4460 (N_4460,N_1805,N_998);
or U4461 (N_4461,N_1890,N_325);
or U4462 (N_4462,N_2395,N_2720);
nand U4463 (N_4463,N_1552,N_2436);
xor U4464 (N_4464,N_2347,N_2023);
nand U4465 (N_4465,N_620,N_1183);
nand U4466 (N_4466,N_2160,N_1515);
or U4467 (N_4467,N_1236,N_2916);
nand U4468 (N_4468,N_2071,N_1251);
nand U4469 (N_4469,N_713,N_2052);
nor U4470 (N_4470,N_812,N_1071);
nand U4471 (N_4471,N_742,N_2206);
nand U4472 (N_4472,N_1259,N_2495);
nand U4473 (N_4473,N_1770,N_3045);
and U4474 (N_4474,N_1378,N_1646);
or U4475 (N_4475,N_2879,N_2707);
xor U4476 (N_4476,N_2531,N_117);
and U4477 (N_4477,N_2791,N_2519);
or U4478 (N_4478,N_2196,N_1156);
or U4479 (N_4479,N_2732,N_2787);
and U4480 (N_4480,N_1231,N_2018);
xnor U4481 (N_4481,N_786,N_1772);
nand U4482 (N_4482,N_1775,N_1018);
or U4483 (N_4483,N_2536,N_2198);
or U4484 (N_4484,N_2639,N_1368);
or U4485 (N_4485,N_2342,N_2258);
or U4486 (N_4486,N_2379,N_2711);
nand U4487 (N_4487,N_811,N_1755);
nor U4488 (N_4488,N_1040,N_2607);
nand U4489 (N_4489,N_2118,N_99);
nand U4490 (N_4490,N_3053,N_404);
nor U4491 (N_4491,N_1655,N_895);
and U4492 (N_4492,N_2858,N_1160);
or U4493 (N_4493,N_444,N_910);
xnor U4494 (N_4494,N_2238,N_837);
nand U4495 (N_4495,N_1023,N_2674);
or U4496 (N_4496,N_1602,N_1404);
and U4497 (N_4497,N_2917,N_1545);
nor U4498 (N_4498,N_722,N_685);
xnor U4499 (N_4499,N_2830,N_203);
nor U4500 (N_4500,N_1966,N_2443);
nand U4501 (N_4501,N_1715,N_955);
nand U4502 (N_4502,N_1569,N_1950);
and U4503 (N_4503,N_2534,N_1120);
and U4504 (N_4504,N_1263,N_1858);
or U4505 (N_4505,N_521,N_2754);
nor U4506 (N_4506,N_182,N_324);
and U4507 (N_4507,N_1644,N_889);
or U4508 (N_4508,N_2015,N_429);
nand U4509 (N_4509,N_688,N_1799);
and U4510 (N_4510,N_1415,N_585);
or U4511 (N_4511,N_2923,N_2114);
and U4512 (N_4512,N_2996,N_2485);
nor U4513 (N_4513,N_1661,N_2494);
or U4514 (N_4514,N_2839,N_3026);
nand U4515 (N_4515,N_2964,N_1842);
or U4516 (N_4516,N_1816,N_2798);
nor U4517 (N_4517,N_225,N_2057);
or U4518 (N_4518,N_1358,N_337);
nor U4519 (N_4519,N_995,N_1363);
or U4520 (N_4520,N_569,N_1460);
and U4521 (N_4521,N_1316,N_1619);
and U4522 (N_4522,N_635,N_2985);
or U4523 (N_4523,N_452,N_1036);
or U4524 (N_4524,N_2199,N_2027);
nand U4525 (N_4525,N_1881,N_1084);
nor U4526 (N_4526,N_2370,N_939);
and U4527 (N_4527,N_3086,N_3119);
nand U4528 (N_4528,N_486,N_2740);
nor U4529 (N_4529,N_1595,N_1869);
or U4530 (N_4530,N_2293,N_2272);
nor U4531 (N_4531,N_1877,N_552);
or U4532 (N_4532,N_438,N_2949);
nor U4533 (N_4533,N_362,N_1912);
or U4534 (N_4534,N_357,N_2229);
and U4535 (N_4535,N_1931,N_3057);
nand U4536 (N_4536,N_1009,N_1810);
nand U4537 (N_4537,N_927,N_1908);
nor U4538 (N_4538,N_2019,N_1059);
or U4539 (N_4539,N_1832,N_1185);
nand U4540 (N_4540,N_2178,N_2427);
xor U4541 (N_4541,N_1204,N_1295);
and U4542 (N_4542,N_772,N_1496);
nor U4543 (N_4543,N_2658,N_2013);
nand U4544 (N_4544,N_2959,N_2863);
and U4545 (N_4545,N_2367,N_1509);
and U4546 (N_4546,N_15,N_2925);
and U4547 (N_4547,N_1600,N_2319);
and U4548 (N_4548,N_885,N_441);
nand U4549 (N_4549,N_1588,N_2990);
xnor U4550 (N_4550,N_2481,N_1979);
nand U4551 (N_4551,N_1093,N_244);
and U4552 (N_4552,N_3019,N_1420);
or U4553 (N_4553,N_210,N_2518);
nand U4554 (N_4554,N_339,N_2236);
nand U4555 (N_4555,N_714,N_2631);
nand U4556 (N_4556,N_678,N_1188);
nand U4557 (N_4557,N_1198,N_2941);
or U4558 (N_4558,N_267,N_1143);
xnor U4559 (N_4559,N_1593,N_1417);
and U4560 (N_4560,N_882,N_2388);
nor U4561 (N_4561,N_1249,N_275);
xor U4562 (N_4562,N_2776,N_1283);
nand U4563 (N_4563,N_2183,N_435);
nand U4564 (N_4564,N_1790,N_1811);
nor U4565 (N_4565,N_1467,N_1483);
nand U4566 (N_4566,N_2412,N_372);
nand U4567 (N_4567,N_2251,N_465);
nand U4568 (N_4568,N_1273,N_2309);
nor U4569 (N_4569,N_1098,N_2132);
nor U4570 (N_4570,N_1328,N_537);
or U4571 (N_4571,N_865,N_916);
nor U4572 (N_4572,N_612,N_1267);
nor U4573 (N_4573,N_1997,N_2497);
nor U4574 (N_4574,N_1441,N_1958);
and U4575 (N_4575,N_1547,N_2904);
and U4576 (N_4576,N_613,N_341);
or U4577 (N_4577,N_1783,N_69);
nor U4578 (N_4578,N_1844,N_350);
xnor U4579 (N_4579,N_2315,N_172);
nor U4580 (N_4580,N_598,N_1754);
nand U4581 (N_4581,N_1938,N_185);
nand U4582 (N_4582,N_2775,N_2526);
xor U4583 (N_4583,N_1057,N_1717);
or U4584 (N_4584,N_1587,N_2011);
and U4585 (N_4585,N_1836,N_2929);
nor U4586 (N_4586,N_1896,N_1822);
nor U4587 (N_4587,N_1640,N_2159);
nand U4588 (N_4588,N_1981,N_1233);
nand U4589 (N_4589,N_133,N_3120);
xnor U4590 (N_4590,N_3113,N_923);
or U4591 (N_4591,N_519,N_1610);
or U4592 (N_4592,N_1984,N_2275);
nor U4593 (N_4593,N_174,N_1262);
xor U4594 (N_4594,N_3015,N_229);
or U4595 (N_4595,N_201,N_190);
nor U4596 (N_4596,N_1978,N_2193);
nand U4597 (N_4597,N_173,N_2889);
or U4598 (N_4598,N_2876,N_222);
xnor U4599 (N_4599,N_878,N_2077);
nand U4600 (N_4600,N_342,N_1174);
nand U4601 (N_4601,N_1275,N_1357);
or U4602 (N_4602,N_2955,N_72);
nor U4603 (N_4603,N_697,N_2396);
and U4604 (N_4604,N_2589,N_1724);
or U4605 (N_4605,N_1326,N_1050);
and U4606 (N_4606,N_503,N_2877);
nor U4607 (N_4607,N_3065,N_388);
nor U4608 (N_4608,N_1407,N_1119);
and U4609 (N_4609,N_1683,N_1576);
nand U4610 (N_4610,N_2297,N_3074);
and U4611 (N_4611,N_1354,N_2233);
nand U4612 (N_4612,N_1730,N_802);
nor U4613 (N_4613,N_2731,N_1245);
xor U4614 (N_4614,N_1428,N_2420);
nand U4615 (N_4615,N_2935,N_2058);
nor U4616 (N_4616,N_1353,N_1274);
and U4617 (N_4617,N_1514,N_735);
or U4618 (N_4618,N_27,N_1746);
or U4619 (N_4619,N_1677,N_2380);
nand U4620 (N_4620,N_2017,N_2366);
or U4621 (N_4621,N_143,N_2868);
and U4622 (N_4622,N_2906,N_829);
and U4623 (N_4623,N_2952,N_2590);
nand U4624 (N_4624,N_95,N_391);
and U4625 (N_4625,N_2137,N_1996);
nand U4626 (N_4626,N_2691,N_575);
or U4627 (N_4627,N_1740,N_96);
or U4628 (N_4628,N_641,N_2471);
and U4629 (N_4629,N_1219,N_2675);
or U4630 (N_4630,N_2329,N_2604);
xor U4631 (N_4631,N_2564,N_359);
nand U4632 (N_4632,N_1493,N_419);
nand U4633 (N_4633,N_933,N_2000);
nand U4634 (N_4634,N_2807,N_1876);
or U4635 (N_4635,N_842,N_2752);
or U4636 (N_4636,N_2406,N_233);
nand U4637 (N_4637,N_1660,N_1242);
or U4638 (N_4638,N_576,N_2257);
nand U4639 (N_4639,N_2669,N_2288);
nand U4640 (N_4640,N_1992,N_2110);
nand U4641 (N_4641,N_479,N_309);
nor U4642 (N_4642,N_1426,N_352);
nor U4643 (N_4643,N_660,N_989);
xnor U4644 (N_4644,N_2248,N_2630);
nor U4645 (N_4645,N_2576,N_577);
nand U4646 (N_4646,N_2570,N_2782);
nor U4647 (N_4647,N_779,N_646);
nand U4648 (N_4648,N_1396,N_322);
or U4649 (N_4649,N_2032,N_2404);
nand U4650 (N_4650,N_2622,N_2498);
nand U4651 (N_4651,N_2601,N_2092);
nand U4652 (N_4652,N_1132,N_2095);
xnor U4653 (N_4653,N_2125,N_332);
xor U4654 (N_4654,N_1270,N_658);
xnor U4655 (N_4655,N_2049,N_262);
or U4656 (N_4656,N_1756,N_942);
and U4657 (N_4657,N_2920,N_1078);
or U4658 (N_4658,N_2149,N_119);
or U4659 (N_4659,N_1169,N_353);
and U4660 (N_4660,N_1750,N_1572);
and U4661 (N_4661,N_1194,N_498);
nor U4662 (N_4662,N_1768,N_584);
nand U4663 (N_4663,N_495,N_907);
or U4664 (N_4664,N_548,N_2186);
or U4665 (N_4665,N_191,N_996);
xnor U4666 (N_4666,N_1155,N_1726);
xor U4667 (N_4667,N_2547,N_1097);
and U4668 (N_4668,N_2662,N_1863);
nor U4669 (N_4669,N_3098,N_1038);
and U4670 (N_4670,N_1443,N_2228);
nor U4671 (N_4671,N_1662,N_3058);
xor U4672 (N_4672,N_755,N_1734);
and U4673 (N_4673,N_2407,N_2623);
and U4674 (N_4674,N_3071,N_3030);
or U4675 (N_4675,N_1721,N_831);
nand U4676 (N_4676,N_2695,N_2520);
and U4677 (N_4677,N_3047,N_969);
nand U4678 (N_4678,N_2264,N_551);
nand U4679 (N_4679,N_2657,N_553);
or U4680 (N_4680,N_1546,N_2036);
or U4681 (N_4681,N_2565,N_1722);
and U4682 (N_4682,N_2261,N_39);
nor U4683 (N_4683,N_1088,N_2841);
and U4684 (N_4684,N_237,N_2177);
nor U4685 (N_4685,N_2129,N_155);
nand U4686 (N_4686,N_1762,N_1752);
and U4687 (N_4687,N_1459,N_2269);
and U4688 (N_4688,N_2003,N_2001);
or U4689 (N_4689,N_1285,N_1479);
or U4690 (N_4690,N_779,N_94);
nand U4691 (N_4691,N_432,N_1896);
nor U4692 (N_4692,N_408,N_362);
nor U4693 (N_4693,N_288,N_2665);
and U4694 (N_4694,N_1882,N_1626);
nor U4695 (N_4695,N_2838,N_2682);
and U4696 (N_4696,N_1106,N_1168);
nand U4697 (N_4697,N_45,N_2600);
and U4698 (N_4698,N_3003,N_2219);
or U4699 (N_4699,N_1025,N_1827);
and U4700 (N_4700,N_405,N_188);
nor U4701 (N_4701,N_2578,N_2067);
nor U4702 (N_4702,N_597,N_2282);
nor U4703 (N_4703,N_112,N_255);
or U4704 (N_4704,N_2023,N_2853);
nor U4705 (N_4705,N_1589,N_127);
and U4706 (N_4706,N_2454,N_2594);
xor U4707 (N_4707,N_2690,N_1226);
xnor U4708 (N_4708,N_664,N_128);
and U4709 (N_4709,N_812,N_1676);
nand U4710 (N_4710,N_373,N_1366);
nor U4711 (N_4711,N_1824,N_650);
or U4712 (N_4712,N_913,N_1704);
or U4713 (N_4713,N_1149,N_802);
or U4714 (N_4714,N_2136,N_146);
and U4715 (N_4715,N_166,N_620);
nand U4716 (N_4716,N_1947,N_1812);
and U4717 (N_4717,N_546,N_1069);
nor U4718 (N_4718,N_2768,N_155);
xnor U4719 (N_4719,N_637,N_2314);
nand U4720 (N_4720,N_2157,N_459);
xnor U4721 (N_4721,N_1896,N_468);
nand U4722 (N_4722,N_238,N_505);
and U4723 (N_4723,N_2168,N_2429);
and U4724 (N_4724,N_64,N_1093);
and U4725 (N_4725,N_782,N_2491);
nor U4726 (N_4726,N_1265,N_2779);
or U4727 (N_4727,N_931,N_2384);
and U4728 (N_4728,N_121,N_551);
or U4729 (N_4729,N_815,N_1638);
and U4730 (N_4730,N_1013,N_2595);
xnor U4731 (N_4731,N_2482,N_2352);
nor U4732 (N_4732,N_1460,N_2104);
or U4733 (N_4733,N_682,N_1320);
or U4734 (N_4734,N_810,N_985);
nand U4735 (N_4735,N_1729,N_1716);
nor U4736 (N_4736,N_50,N_1351);
nand U4737 (N_4737,N_2833,N_2644);
nor U4738 (N_4738,N_2342,N_1681);
or U4739 (N_4739,N_82,N_1824);
nand U4740 (N_4740,N_1663,N_629);
nand U4741 (N_4741,N_2388,N_56);
nand U4742 (N_4742,N_1066,N_2900);
nand U4743 (N_4743,N_2578,N_1367);
and U4744 (N_4744,N_1338,N_2606);
nor U4745 (N_4745,N_2552,N_2846);
nand U4746 (N_4746,N_2184,N_410);
and U4747 (N_4747,N_1273,N_171);
nand U4748 (N_4748,N_1934,N_1875);
xnor U4749 (N_4749,N_1066,N_2922);
nor U4750 (N_4750,N_2311,N_2872);
and U4751 (N_4751,N_1015,N_2434);
nand U4752 (N_4752,N_408,N_2618);
and U4753 (N_4753,N_2077,N_48);
or U4754 (N_4754,N_1438,N_2784);
nand U4755 (N_4755,N_2450,N_1188);
nor U4756 (N_4756,N_2429,N_458);
and U4757 (N_4757,N_2130,N_2771);
nor U4758 (N_4758,N_1806,N_918);
xnor U4759 (N_4759,N_428,N_2484);
xor U4760 (N_4760,N_1819,N_2341);
and U4761 (N_4761,N_1049,N_1913);
nand U4762 (N_4762,N_330,N_1794);
xor U4763 (N_4763,N_2737,N_301);
and U4764 (N_4764,N_1144,N_2756);
or U4765 (N_4765,N_1403,N_1610);
or U4766 (N_4766,N_1760,N_2016);
nor U4767 (N_4767,N_242,N_682);
and U4768 (N_4768,N_1925,N_2495);
nand U4769 (N_4769,N_1287,N_1138);
xnor U4770 (N_4770,N_2416,N_2938);
and U4771 (N_4771,N_1381,N_1609);
and U4772 (N_4772,N_2127,N_2807);
xnor U4773 (N_4773,N_95,N_202);
and U4774 (N_4774,N_333,N_1265);
or U4775 (N_4775,N_412,N_2836);
and U4776 (N_4776,N_573,N_267);
or U4777 (N_4777,N_1863,N_2598);
and U4778 (N_4778,N_508,N_2193);
nand U4779 (N_4779,N_2175,N_351);
and U4780 (N_4780,N_1582,N_1566);
nand U4781 (N_4781,N_179,N_1232);
and U4782 (N_4782,N_2043,N_817);
nand U4783 (N_4783,N_2863,N_1444);
nand U4784 (N_4784,N_2807,N_1358);
or U4785 (N_4785,N_1519,N_3055);
nand U4786 (N_4786,N_286,N_1444);
and U4787 (N_4787,N_1995,N_1743);
and U4788 (N_4788,N_1771,N_2462);
nor U4789 (N_4789,N_1881,N_2975);
nand U4790 (N_4790,N_492,N_2831);
nor U4791 (N_4791,N_2359,N_1329);
nand U4792 (N_4792,N_1358,N_477);
and U4793 (N_4793,N_2243,N_1062);
nand U4794 (N_4794,N_2587,N_184);
nor U4795 (N_4795,N_232,N_344);
nor U4796 (N_4796,N_196,N_1117);
or U4797 (N_4797,N_97,N_1102);
nor U4798 (N_4798,N_1915,N_2808);
or U4799 (N_4799,N_2360,N_1546);
and U4800 (N_4800,N_215,N_2569);
nand U4801 (N_4801,N_449,N_2348);
xor U4802 (N_4802,N_908,N_637);
nor U4803 (N_4803,N_377,N_1871);
xnor U4804 (N_4804,N_378,N_441);
or U4805 (N_4805,N_1135,N_2844);
and U4806 (N_4806,N_311,N_345);
or U4807 (N_4807,N_2426,N_969);
and U4808 (N_4808,N_2505,N_1286);
xor U4809 (N_4809,N_428,N_1550);
or U4810 (N_4810,N_2002,N_1551);
nand U4811 (N_4811,N_1979,N_1497);
or U4812 (N_4812,N_1989,N_317);
and U4813 (N_4813,N_402,N_1476);
or U4814 (N_4814,N_193,N_2263);
nor U4815 (N_4815,N_2646,N_2412);
or U4816 (N_4816,N_2699,N_1252);
or U4817 (N_4817,N_383,N_339);
and U4818 (N_4818,N_65,N_3124);
nor U4819 (N_4819,N_2290,N_2476);
and U4820 (N_4820,N_2725,N_2072);
nor U4821 (N_4821,N_2826,N_596);
or U4822 (N_4822,N_2320,N_321);
xor U4823 (N_4823,N_1907,N_863);
or U4824 (N_4824,N_2596,N_1851);
xor U4825 (N_4825,N_1205,N_1451);
or U4826 (N_4826,N_1964,N_2396);
and U4827 (N_4827,N_1015,N_240);
nand U4828 (N_4828,N_1437,N_2528);
nor U4829 (N_4829,N_1943,N_904);
nand U4830 (N_4830,N_2574,N_2253);
nor U4831 (N_4831,N_1866,N_859);
or U4832 (N_4832,N_2161,N_1378);
nor U4833 (N_4833,N_1580,N_812);
or U4834 (N_4834,N_2036,N_719);
and U4835 (N_4835,N_361,N_742);
nand U4836 (N_4836,N_328,N_2792);
or U4837 (N_4837,N_500,N_562);
nand U4838 (N_4838,N_1255,N_2341);
xnor U4839 (N_4839,N_1365,N_3053);
nand U4840 (N_4840,N_1619,N_2060);
and U4841 (N_4841,N_1641,N_2328);
or U4842 (N_4842,N_155,N_2884);
nand U4843 (N_4843,N_2993,N_2079);
or U4844 (N_4844,N_914,N_2375);
or U4845 (N_4845,N_2283,N_2808);
nand U4846 (N_4846,N_2478,N_1159);
nor U4847 (N_4847,N_1069,N_1117);
xnor U4848 (N_4848,N_2824,N_21);
nand U4849 (N_4849,N_2331,N_1709);
or U4850 (N_4850,N_2521,N_1437);
or U4851 (N_4851,N_2905,N_105);
and U4852 (N_4852,N_3009,N_602);
nand U4853 (N_4853,N_384,N_942);
nor U4854 (N_4854,N_1735,N_2934);
nand U4855 (N_4855,N_2399,N_13);
nand U4856 (N_4856,N_1799,N_485);
nand U4857 (N_4857,N_2900,N_2459);
xor U4858 (N_4858,N_504,N_527);
nor U4859 (N_4859,N_459,N_3102);
or U4860 (N_4860,N_448,N_216);
nand U4861 (N_4861,N_2803,N_1318);
nand U4862 (N_4862,N_1326,N_2470);
nor U4863 (N_4863,N_1989,N_109);
and U4864 (N_4864,N_1357,N_2612);
and U4865 (N_4865,N_2218,N_933);
or U4866 (N_4866,N_2970,N_351);
nand U4867 (N_4867,N_2611,N_401);
nand U4868 (N_4868,N_52,N_663);
or U4869 (N_4869,N_1974,N_2257);
or U4870 (N_4870,N_583,N_2739);
xnor U4871 (N_4871,N_1421,N_2098);
or U4872 (N_4872,N_79,N_1532);
and U4873 (N_4873,N_1155,N_2640);
xnor U4874 (N_4874,N_276,N_2966);
nand U4875 (N_4875,N_829,N_2963);
nand U4876 (N_4876,N_391,N_2314);
nor U4877 (N_4877,N_2843,N_2397);
nand U4878 (N_4878,N_2454,N_1615);
nand U4879 (N_4879,N_1157,N_2294);
or U4880 (N_4880,N_167,N_1610);
and U4881 (N_4881,N_1516,N_2837);
or U4882 (N_4882,N_1911,N_1116);
and U4883 (N_4883,N_138,N_2185);
and U4884 (N_4884,N_2674,N_499);
xnor U4885 (N_4885,N_1176,N_2815);
or U4886 (N_4886,N_2698,N_1541);
nand U4887 (N_4887,N_386,N_78);
nor U4888 (N_4888,N_2550,N_641);
or U4889 (N_4889,N_2882,N_1905);
and U4890 (N_4890,N_161,N_11);
nor U4891 (N_4891,N_1456,N_2152);
nor U4892 (N_4892,N_1785,N_1867);
and U4893 (N_4893,N_2064,N_2605);
xnor U4894 (N_4894,N_1768,N_2912);
or U4895 (N_4895,N_18,N_996);
xnor U4896 (N_4896,N_180,N_2036);
and U4897 (N_4897,N_283,N_378);
and U4898 (N_4898,N_2471,N_2673);
or U4899 (N_4899,N_333,N_2861);
xor U4900 (N_4900,N_2337,N_288);
nor U4901 (N_4901,N_1608,N_2627);
nand U4902 (N_4902,N_699,N_3020);
nor U4903 (N_4903,N_2007,N_2084);
nor U4904 (N_4904,N_455,N_465);
or U4905 (N_4905,N_910,N_530);
nor U4906 (N_4906,N_1803,N_19);
nor U4907 (N_4907,N_1487,N_1311);
and U4908 (N_4908,N_2054,N_1905);
nor U4909 (N_4909,N_658,N_2479);
nor U4910 (N_4910,N_1656,N_1889);
xor U4911 (N_4911,N_1134,N_282);
nor U4912 (N_4912,N_3040,N_2733);
and U4913 (N_4913,N_2003,N_2137);
xnor U4914 (N_4914,N_2147,N_1623);
and U4915 (N_4915,N_2175,N_957);
or U4916 (N_4916,N_205,N_1006);
or U4917 (N_4917,N_1997,N_822);
nor U4918 (N_4918,N_3052,N_2727);
or U4919 (N_4919,N_2611,N_2320);
nand U4920 (N_4920,N_3122,N_251);
xnor U4921 (N_4921,N_56,N_1407);
nand U4922 (N_4922,N_1135,N_1017);
xnor U4923 (N_4923,N_1012,N_446);
nand U4924 (N_4924,N_2949,N_1335);
and U4925 (N_4925,N_69,N_2304);
and U4926 (N_4926,N_2370,N_960);
or U4927 (N_4927,N_2439,N_2621);
xnor U4928 (N_4928,N_1979,N_1130);
or U4929 (N_4929,N_4,N_302);
or U4930 (N_4930,N_420,N_2680);
nor U4931 (N_4931,N_2382,N_1593);
and U4932 (N_4932,N_1904,N_1260);
and U4933 (N_4933,N_2056,N_1950);
and U4934 (N_4934,N_2667,N_2254);
nor U4935 (N_4935,N_1958,N_2080);
or U4936 (N_4936,N_825,N_1276);
and U4937 (N_4937,N_965,N_156);
nor U4938 (N_4938,N_955,N_2232);
or U4939 (N_4939,N_964,N_1844);
nor U4940 (N_4940,N_1739,N_654);
nand U4941 (N_4941,N_1672,N_193);
nand U4942 (N_4942,N_614,N_1805);
nand U4943 (N_4943,N_597,N_711);
nand U4944 (N_4944,N_1507,N_804);
and U4945 (N_4945,N_2421,N_1931);
nand U4946 (N_4946,N_510,N_122);
nor U4947 (N_4947,N_95,N_1117);
or U4948 (N_4948,N_3106,N_1904);
xnor U4949 (N_4949,N_246,N_1068);
or U4950 (N_4950,N_2034,N_2454);
and U4951 (N_4951,N_1482,N_1079);
and U4952 (N_4952,N_1203,N_1804);
or U4953 (N_4953,N_1942,N_2321);
nor U4954 (N_4954,N_1614,N_1885);
nor U4955 (N_4955,N_2961,N_2043);
nand U4956 (N_4956,N_519,N_598);
xnor U4957 (N_4957,N_1671,N_147);
and U4958 (N_4958,N_1105,N_2476);
or U4959 (N_4959,N_641,N_2031);
nor U4960 (N_4960,N_3012,N_2143);
and U4961 (N_4961,N_2035,N_2786);
nor U4962 (N_4962,N_331,N_74);
xnor U4963 (N_4963,N_984,N_2617);
nand U4964 (N_4964,N_1977,N_1373);
nand U4965 (N_4965,N_2465,N_481);
and U4966 (N_4966,N_1453,N_309);
nor U4967 (N_4967,N_127,N_1618);
xnor U4968 (N_4968,N_1910,N_2012);
and U4969 (N_4969,N_484,N_2093);
and U4970 (N_4970,N_1960,N_1876);
and U4971 (N_4971,N_1235,N_2794);
xor U4972 (N_4972,N_2796,N_2295);
nor U4973 (N_4973,N_227,N_1640);
and U4974 (N_4974,N_83,N_326);
and U4975 (N_4975,N_740,N_2425);
nor U4976 (N_4976,N_2977,N_2399);
nand U4977 (N_4977,N_742,N_977);
nor U4978 (N_4978,N_3006,N_579);
and U4979 (N_4979,N_159,N_1782);
nor U4980 (N_4980,N_2483,N_2723);
and U4981 (N_4981,N_2768,N_2227);
xor U4982 (N_4982,N_924,N_1031);
nand U4983 (N_4983,N_128,N_2929);
or U4984 (N_4984,N_1245,N_3104);
nor U4985 (N_4985,N_908,N_424);
xnor U4986 (N_4986,N_160,N_2134);
or U4987 (N_4987,N_1133,N_919);
and U4988 (N_4988,N_2465,N_111);
or U4989 (N_4989,N_379,N_316);
xor U4990 (N_4990,N_1082,N_403);
xnor U4991 (N_4991,N_241,N_2747);
and U4992 (N_4992,N_2738,N_1627);
nor U4993 (N_4993,N_3101,N_839);
nand U4994 (N_4994,N_1099,N_2101);
nand U4995 (N_4995,N_77,N_2615);
or U4996 (N_4996,N_2244,N_596);
or U4997 (N_4997,N_616,N_636);
or U4998 (N_4998,N_2293,N_2071);
nor U4999 (N_4999,N_1152,N_2293);
and U5000 (N_5000,N_1326,N_122);
nand U5001 (N_5001,N_576,N_3011);
and U5002 (N_5002,N_1253,N_1390);
nand U5003 (N_5003,N_551,N_1877);
and U5004 (N_5004,N_465,N_56);
or U5005 (N_5005,N_1491,N_870);
and U5006 (N_5006,N_2665,N_1479);
or U5007 (N_5007,N_1290,N_850);
nor U5008 (N_5008,N_2066,N_241);
nor U5009 (N_5009,N_1704,N_2813);
nor U5010 (N_5010,N_2443,N_2870);
or U5011 (N_5011,N_2005,N_1241);
nand U5012 (N_5012,N_252,N_1679);
nand U5013 (N_5013,N_2676,N_1717);
and U5014 (N_5014,N_2575,N_621);
or U5015 (N_5015,N_2291,N_1938);
and U5016 (N_5016,N_598,N_2881);
nand U5017 (N_5017,N_1359,N_1632);
nor U5018 (N_5018,N_605,N_1086);
and U5019 (N_5019,N_120,N_1185);
xnor U5020 (N_5020,N_1700,N_720);
and U5021 (N_5021,N_1535,N_563);
nor U5022 (N_5022,N_753,N_1321);
and U5023 (N_5023,N_889,N_2035);
or U5024 (N_5024,N_257,N_1457);
and U5025 (N_5025,N_81,N_1415);
and U5026 (N_5026,N_952,N_2667);
nand U5027 (N_5027,N_1697,N_2895);
or U5028 (N_5028,N_832,N_1035);
or U5029 (N_5029,N_2330,N_1745);
nand U5030 (N_5030,N_1581,N_756);
nor U5031 (N_5031,N_648,N_520);
nand U5032 (N_5032,N_2282,N_598);
nor U5033 (N_5033,N_2272,N_159);
or U5034 (N_5034,N_1999,N_1889);
or U5035 (N_5035,N_1674,N_547);
and U5036 (N_5036,N_1704,N_1669);
or U5037 (N_5037,N_1007,N_1309);
nand U5038 (N_5038,N_810,N_157);
nor U5039 (N_5039,N_3009,N_2287);
nor U5040 (N_5040,N_1995,N_2715);
nor U5041 (N_5041,N_1008,N_1738);
xnor U5042 (N_5042,N_766,N_2719);
or U5043 (N_5043,N_1969,N_1362);
nor U5044 (N_5044,N_445,N_1972);
and U5045 (N_5045,N_413,N_1466);
and U5046 (N_5046,N_970,N_1410);
nor U5047 (N_5047,N_2344,N_307);
or U5048 (N_5048,N_37,N_2191);
or U5049 (N_5049,N_2600,N_961);
or U5050 (N_5050,N_1291,N_2816);
nand U5051 (N_5051,N_1752,N_493);
nor U5052 (N_5052,N_1350,N_733);
or U5053 (N_5053,N_2071,N_228);
nand U5054 (N_5054,N_1478,N_247);
and U5055 (N_5055,N_2394,N_531);
xnor U5056 (N_5056,N_1343,N_1396);
nor U5057 (N_5057,N_701,N_1311);
nand U5058 (N_5058,N_827,N_1736);
and U5059 (N_5059,N_1321,N_883);
and U5060 (N_5060,N_2635,N_2310);
and U5061 (N_5061,N_1037,N_2830);
xor U5062 (N_5062,N_2046,N_2039);
and U5063 (N_5063,N_1066,N_456);
and U5064 (N_5064,N_59,N_2617);
xnor U5065 (N_5065,N_1711,N_3097);
nor U5066 (N_5066,N_2428,N_1070);
or U5067 (N_5067,N_1809,N_1171);
or U5068 (N_5068,N_2526,N_1915);
nand U5069 (N_5069,N_2913,N_2489);
nor U5070 (N_5070,N_2241,N_1917);
nand U5071 (N_5071,N_1290,N_2538);
or U5072 (N_5072,N_2872,N_2377);
nor U5073 (N_5073,N_2379,N_2437);
nand U5074 (N_5074,N_2547,N_2265);
or U5075 (N_5075,N_999,N_2104);
xor U5076 (N_5076,N_2961,N_2937);
xnor U5077 (N_5077,N_2116,N_3085);
or U5078 (N_5078,N_414,N_2647);
or U5079 (N_5079,N_1036,N_1926);
nand U5080 (N_5080,N_2841,N_1291);
or U5081 (N_5081,N_1225,N_82);
or U5082 (N_5082,N_1072,N_1378);
and U5083 (N_5083,N_2759,N_1553);
or U5084 (N_5084,N_304,N_1760);
and U5085 (N_5085,N_1812,N_77);
and U5086 (N_5086,N_111,N_1138);
and U5087 (N_5087,N_868,N_100);
nor U5088 (N_5088,N_225,N_1914);
nand U5089 (N_5089,N_3046,N_505);
nor U5090 (N_5090,N_1842,N_1798);
and U5091 (N_5091,N_205,N_71);
nand U5092 (N_5092,N_770,N_382);
or U5093 (N_5093,N_2064,N_1379);
or U5094 (N_5094,N_1061,N_2852);
and U5095 (N_5095,N_506,N_1795);
nand U5096 (N_5096,N_1108,N_1963);
and U5097 (N_5097,N_2565,N_487);
nand U5098 (N_5098,N_592,N_1578);
and U5099 (N_5099,N_1762,N_78);
or U5100 (N_5100,N_135,N_810);
or U5101 (N_5101,N_2705,N_2779);
xnor U5102 (N_5102,N_2122,N_3086);
nand U5103 (N_5103,N_652,N_908);
nor U5104 (N_5104,N_1863,N_1132);
nand U5105 (N_5105,N_2805,N_579);
nor U5106 (N_5106,N_146,N_2513);
nand U5107 (N_5107,N_2662,N_2270);
and U5108 (N_5108,N_59,N_759);
nor U5109 (N_5109,N_1335,N_1588);
or U5110 (N_5110,N_2541,N_1143);
nand U5111 (N_5111,N_2504,N_2879);
xor U5112 (N_5112,N_2925,N_2993);
nor U5113 (N_5113,N_28,N_2712);
or U5114 (N_5114,N_2675,N_844);
nand U5115 (N_5115,N_1780,N_730);
or U5116 (N_5116,N_2319,N_2876);
nand U5117 (N_5117,N_477,N_1857);
or U5118 (N_5118,N_291,N_2623);
nand U5119 (N_5119,N_2013,N_1293);
xnor U5120 (N_5120,N_411,N_1126);
nand U5121 (N_5121,N_623,N_27);
nor U5122 (N_5122,N_573,N_477);
xnor U5123 (N_5123,N_2954,N_318);
and U5124 (N_5124,N_1916,N_1985);
nor U5125 (N_5125,N_2678,N_2811);
and U5126 (N_5126,N_83,N_2634);
nor U5127 (N_5127,N_1842,N_2832);
or U5128 (N_5128,N_2857,N_2977);
or U5129 (N_5129,N_3029,N_1748);
nand U5130 (N_5130,N_313,N_1014);
nand U5131 (N_5131,N_1440,N_2608);
or U5132 (N_5132,N_580,N_2317);
nor U5133 (N_5133,N_645,N_2942);
nor U5134 (N_5134,N_581,N_129);
nor U5135 (N_5135,N_899,N_2059);
and U5136 (N_5136,N_741,N_2288);
nand U5137 (N_5137,N_1547,N_3003);
nand U5138 (N_5138,N_823,N_318);
nor U5139 (N_5139,N_2385,N_2114);
or U5140 (N_5140,N_562,N_2137);
or U5141 (N_5141,N_2510,N_2426);
nand U5142 (N_5142,N_1623,N_2129);
nor U5143 (N_5143,N_2321,N_68);
and U5144 (N_5144,N_1739,N_2363);
and U5145 (N_5145,N_1872,N_1216);
or U5146 (N_5146,N_1076,N_2308);
nor U5147 (N_5147,N_605,N_2349);
xnor U5148 (N_5148,N_2908,N_2395);
xnor U5149 (N_5149,N_1685,N_3014);
nor U5150 (N_5150,N_2371,N_636);
nor U5151 (N_5151,N_995,N_1056);
nor U5152 (N_5152,N_699,N_2822);
xnor U5153 (N_5153,N_3121,N_801);
nand U5154 (N_5154,N_382,N_2045);
nor U5155 (N_5155,N_2711,N_2317);
or U5156 (N_5156,N_2813,N_555);
and U5157 (N_5157,N_2537,N_336);
or U5158 (N_5158,N_500,N_1258);
and U5159 (N_5159,N_1172,N_452);
nand U5160 (N_5160,N_2209,N_1574);
and U5161 (N_5161,N_201,N_834);
xnor U5162 (N_5162,N_1484,N_1483);
nand U5163 (N_5163,N_2416,N_629);
and U5164 (N_5164,N_1904,N_2376);
or U5165 (N_5165,N_1387,N_1967);
and U5166 (N_5166,N_1842,N_2968);
and U5167 (N_5167,N_1581,N_508);
and U5168 (N_5168,N_2141,N_540);
or U5169 (N_5169,N_813,N_2388);
and U5170 (N_5170,N_1884,N_2483);
nand U5171 (N_5171,N_1757,N_2737);
or U5172 (N_5172,N_1341,N_1442);
nor U5173 (N_5173,N_1998,N_1444);
nand U5174 (N_5174,N_2224,N_2467);
nor U5175 (N_5175,N_698,N_931);
nor U5176 (N_5176,N_1522,N_1435);
or U5177 (N_5177,N_2953,N_46);
nand U5178 (N_5178,N_746,N_659);
and U5179 (N_5179,N_1725,N_2152);
or U5180 (N_5180,N_1872,N_184);
nor U5181 (N_5181,N_709,N_702);
nand U5182 (N_5182,N_1727,N_1438);
nor U5183 (N_5183,N_1385,N_623);
or U5184 (N_5184,N_1150,N_145);
and U5185 (N_5185,N_119,N_1405);
and U5186 (N_5186,N_452,N_2589);
or U5187 (N_5187,N_458,N_1532);
or U5188 (N_5188,N_864,N_1228);
and U5189 (N_5189,N_1290,N_125);
nand U5190 (N_5190,N_1522,N_2656);
nand U5191 (N_5191,N_190,N_2758);
and U5192 (N_5192,N_142,N_208);
and U5193 (N_5193,N_2012,N_664);
and U5194 (N_5194,N_2284,N_2340);
nor U5195 (N_5195,N_989,N_3042);
or U5196 (N_5196,N_1267,N_3118);
and U5197 (N_5197,N_669,N_611);
xnor U5198 (N_5198,N_1520,N_2033);
xnor U5199 (N_5199,N_304,N_1434);
nor U5200 (N_5200,N_1868,N_226);
xnor U5201 (N_5201,N_1692,N_577);
nor U5202 (N_5202,N_2910,N_2172);
nor U5203 (N_5203,N_2622,N_1003);
nor U5204 (N_5204,N_2846,N_328);
and U5205 (N_5205,N_684,N_2732);
nor U5206 (N_5206,N_3068,N_1018);
nand U5207 (N_5207,N_1504,N_68);
nand U5208 (N_5208,N_2781,N_2505);
nand U5209 (N_5209,N_841,N_1132);
xnor U5210 (N_5210,N_2051,N_1822);
or U5211 (N_5211,N_657,N_2894);
nor U5212 (N_5212,N_2560,N_1011);
xor U5213 (N_5213,N_2926,N_2780);
nor U5214 (N_5214,N_1293,N_2532);
nor U5215 (N_5215,N_505,N_1506);
nand U5216 (N_5216,N_1527,N_1665);
nand U5217 (N_5217,N_2289,N_733);
nand U5218 (N_5218,N_2051,N_2053);
or U5219 (N_5219,N_138,N_2416);
or U5220 (N_5220,N_2812,N_1599);
nor U5221 (N_5221,N_975,N_1443);
nand U5222 (N_5222,N_645,N_2711);
and U5223 (N_5223,N_2957,N_2919);
nor U5224 (N_5224,N_899,N_1513);
and U5225 (N_5225,N_2350,N_1729);
nor U5226 (N_5226,N_1931,N_1530);
and U5227 (N_5227,N_2032,N_1728);
or U5228 (N_5228,N_172,N_2817);
nor U5229 (N_5229,N_989,N_2820);
xnor U5230 (N_5230,N_718,N_1676);
nor U5231 (N_5231,N_13,N_593);
or U5232 (N_5232,N_1659,N_1552);
and U5233 (N_5233,N_2377,N_192);
or U5234 (N_5234,N_105,N_25);
and U5235 (N_5235,N_2429,N_752);
xnor U5236 (N_5236,N_1314,N_2759);
nor U5237 (N_5237,N_1116,N_2634);
and U5238 (N_5238,N_3081,N_2743);
or U5239 (N_5239,N_1611,N_320);
nand U5240 (N_5240,N_170,N_1869);
nand U5241 (N_5241,N_2190,N_2116);
nor U5242 (N_5242,N_1764,N_939);
and U5243 (N_5243,N_402,N_1146);
nand U5244 (N_5244,N_2294,N_2461);
or U5245 (N_5245,N_1180,N_545);
xor U5246 (N_5246,N_1280,N_731);
and U5247 (N_5247,N_2399,N_1429);
xnor U5248 (N_5248,N_1319,N_1792);
nand U5249 (N_5249,N_2831,N_1834);
xor U5250 (N_5250,N_2748,N_1478);
nor U5251 (N_5251,N_1936,N_1518);
nor U5252 (N_5252,N_2532,N_1823);
and U5253 (N_5253,N_223,N_1557);
or U5254 (N_5254,N_2671,N_1511);
and U5255 (N_5255,N_2448,N_290);
nor U5256 (N_5256,N_1854,N_1141);
and U5257 (N_5257,N_303,N_1966);
nor U5258 (N_5258,N_990,N_1226);
or U5259 (N_5259,N_481,N_2758);
nand U5260 (N_5260,N_1437,N_1930);
nand U5261 (N_5261,N_3108,N_3092);
nand U5262 (N_5262,N_307,N_2775);
nor U5263 (N_5263,N_1529,N_329);
or U5264 (N_5264,N_1708,N_2838);
nor U5265 (N_5265,N_2729,N_1661);
nor U5266 (N_5266,N_2684,N_88);
nand U5267 (N_5267,N_2804,N_2652);
and U5268 (N_5268,N_1928,N_59);
xnor U5269 (N_5269,N_1770,N_2607);
and U5270 (N_5270,N_1365,N_181);
nor U5271 (N_5271,N_252,N_835);
nand U5272 (N_5272,N_2056,N_85);
nand U5273 (N_5273,N_1515,N_291);
and U5274 (N_5274,N_489,N_1632);
and U5275 (N_5275,N_2450,N_810);
nand U5276 (N_5276,N_2109,N_3048);
and U5277 (N_5277,N_687,N_2798);
and U5278 (N_5278,N_3054,N_2871);
xnor U5279 (N_5279,N_1193,N_278);
or U5280 (N_5280,N_2198,N_265);
nor U5281 (N_5281,N_8,N_2556);
or U5282 (N_5282,N_636,N_344);
nor U5283 (N_5283,N_2307,N_2522);
nor U5284 (N_5284,N_1352,N_1998);
and U5285 (N_5285,N_81,N_2563);
xnor U5286 (N_5286,N_746,N_619);
xnor U5287 (N_5287,N_2452,N_1056);
nor U5288 (N_5288,N_1006,N_592);
or U5289 (N_5289,N_1489,N_759);
or U5290 (N_5290,N_2819,N_856);
nor U5291 (N_5291,N_2458,N_1281);
nand U5292 (N_5292,N_2274,N_296);
and U5293 (N_5293,N_156,N_3021);
nand U5294 (N_5294,N_1568,N_2202);
nand U5295 (N_5295,N_205,N_1399);
and U5296 (N_5296,N_1362,N_2103);
nor U5297 (N_5297,N_628,N_48);
nand U5298 (N_5298,N_2403,N_1998);
nor U5299 (N_5299,N_1276,N_1053);
or U5300 (N_5300,N_2854,N_1769);
nand U5301 (N_5301,N_2451,N_1285);
or U5302 (N_5302,N_923,N_2793);
nand U5303 (N_5303,N_2040,N_527);
nor U5304 (N_5304,N_1571,N_2905);
and U5305 (N_5305,N_258,N_1340);
nand U5306 (N_5306,N_962,N_2973);
nor U5307 (N_5307,N_2519,N_1775);
xor U5308 (N_5308,N_2715,N_2390);
nand U5309 (N_5309,N_1991,N_2053);
nor U5310 (N_5310,N_1785,N_333);
or U5311 (N_5311,N_982,N_1103);
nand U5312 (N_5312,N_2274,N_2124);
nor U5313 (N_5313,N_691,N_1239);
nand U5314 (N_5314,N_2544,N_1548);
and U5315 (N_5315,N_4,N_2967);
or U5316 (N_5316,N_927,N_1145);
xor U5317 (N_5317,N_713,N_1670);
xnor U5318 (N_5318,N_783,N_2949);
nor U5319 (N_5319,N_1267,N_87);
and U5320 (N_5320,N_2590,N_2409);
and U5321 (N_5321,N_850,N_18);
nor U5322 (N_5322,N_2450,N_1157);
or U5323 (N_5323,N_1005,N_707);
nor U5324 (N_5324,N_314,N_2093);
nor U5325 (N_5325,N_1031,N_2334);
nand U5326 (N_5326,N_1207,N_2900);
and U5327 (N_5327,N_2358,N_173);
nor U5328 (N_5328,N_3047,N_1242);
and U5329 (N_5329,N_2260,N_2893);
nor U5330 (N_5330,N_3062,N_590);
xor U5331 (N_5331,N_1983,N_2261);
xnor U5332 (N_5332,N_1254,N_1576);
and U5333 (N_5333,N_462,N_2823);
or U5334 (N_5334,N_1093,N_2871);
and U5335 (N_5335,N_831,N_1516);
nand U5336 (N_5336,N_395,N_858);
nand U5337 (N_5337,N_259,N_1983);
and U5338 (N_5338,N_459,N_555);
nor U5339 (N_5339,N_916,N_671);
nor U5340 (N_5340,N_746,N_1754);
or U5341 (N_5341,N_1380,N_2590);
nor U5342 (N_5342,N_269,N_1234);
nand U5343 (N_5343,N_1931,N_238);
nor U5344 (N_5344,N_1000,N_3120);
nor U5345 (N_5345,N_2100,N_3080);
nor U5346 (N_5346,N_1860,N_2784);
and U5347 (N_5347,N_2012,N_2359);
xor U5348 (N_5348,N_2835,N_197);
xnor U5349 (N_5349,N_1025,N_282);
and U5350 (N_5350,N_1477,N_2635);
and U5351 (N_5351,N_1156,N_2192);
or U5352 (N_5352,N_1632,N_2726);
and U5353 (N_5353,N_675,N_1393);
nand U5354 (N_5354,N_3104,N_1115);
and U5355 (N_5355,N_1966,N_1216);
nor U5356 (N_5356,N_2115,N_2310);
nor U5357 (N_5357,N_1820,N_2465);
and U5358 (N_5358,N_1701,N_1989);
or U5359 (N_5359,N_1874,N_1120);
or U5360 (N_5360,N_1267,N_2004);
or U5361 (N_5361,N_2469,N_217);
nor U5362 (N_5362,N_2969,N_746);
nor U5363 (N_5363,N_2300,N_1598);
nor U5364 (N_5364,N_643,N_1391);
and U5365 (N_5365,N_443,N_911);
and U5366 (N_5366,N_467,N_2783);
nand U5367 (N_5367,N_69,N_329);
nand U5368 (N_5368,N_1256,N_1251);
nand U5369 (N_5369,N_1201,N_837);
and U5370 (N_5370,N_2585,N_2992);
and U5371 (N_5371,N_1555,N_971);
nor U5372 (N_5372,N_2263,N_2985);
xnor U5373 (N_5373,N_2895,N_681);
or U5374 (N_5374,N_2410,N_517);
or U5375 (N_5375,N_2385,N_2216);
xor U5376 (N_5376,N_1097,N_3006);
or U5377 (N_5377,N_111,N_33);
xor U5378 (N_5378,N_2903,N_1440);
nand U5379 (N_5379,N_313,N_1609);
or U5380 (N_5380,N_2120,N_823);
or U5381 (N_5381,N_741,N_2142);
and U5382 (N_5382,N_1746,N_1455);
nor U5383 (N_5383,N_2740,N_1028);
nand U5384 (N_5384,N_381,N_124);
nand U5385 (N_5385,N_2858,N_2027);
nand U5386 (N_5386,N_1225,N_2398);
nor U5387 (N_5387,N_677,N_1163);
and U5388 (N_5388,N_57,N_2327);
nor U5389 (N_5389,N_1768,N_2776);
nor U5390 (N_5390,N_2193,N_339);
or U5391 (N_5391,N_1255,N_2826);
nand U5392 (N_5392,N_1913,N_754);
or U5393 (N_5393,N_689,N_1985);
or U5394 (N_5394,N_2615,N_1025);
nand U5395 (N_5395,N_1532,N_93);
nand U5396 (N_5396,N_2672,N_1500);
nor U5397 (N_5397,N_1078,N_2770);
nand U5398 (N_5398,N_1011,N_815);
nand U5399 (N_5399,N_359,N_413);
or U5400 (N_5400,N_135,N_1194);
nand U5401 (N_5401,N_879,N_90);
and U5402 (N_5402,N_1698,N_593);
nand U5403 (N_5403,N_1422,N_1652);
nor U5404 (N_5404,N_1698,N_2044);
or U5405 (N_5405,N_479,N_908);
and U5406 (N_5406,N_2958,N_520);
or U5407 (N_5407,N_1821,N_1047);
and U5408 (N_5408,N_255,N_1366);
and U5409 (N_5409,N_2246,N_2573);
nand U5410 (N_5410,N_2989,N_207);
nor U5411 (N_5411,N_1926,N_2182);
and U5412 (N_5412,N_1725,N_2854);
nor U5413 (N_5413,N_428,N_179);
nor U5414 (N_5414,N_1360,N_159);
or U5415 (N_5415,N_632,N_460);
or U5416 (N_5416,N_866,N_1800);
and U5417 (N_5417,N_1504,N_103);
nand U5418 (N_5418,N_2103,N_1803);
or U5419 (N_5419,N_2329,N_1415);
or U5420 (N_5420,N_2129,N_1124);
and U5421 (N_5421,N_2514,N_2711);
nand U5422 (N_5422,N_1151,N_1632);
nand U5423 (N_5423,N_814,N_2645);
nand U5424 (N_5424,N_633,N_1033);
and U5425 (N_5425,N_2588,N_1302);
and U5426 (N_5426,N_2809,N_2439);
nand U5427 (N_5427,N_1347,N_3055);
nand U5428 (N_5428,N_420,N_148);
nand U5429 (N_5429,N_3032,N_2867);
nand U5430 (N_5430,N_2171,N_2215);
and U5431 (N_5431,N_1068,N_2169);
nor U5432 (N_5432,N_1785,N_2857);
nand U5433 (N_5433,N_912,N_2356);
nor U5434 (N_5434,N_1449,N_2564);
and U5435 (N_5435,N_1591,N_98);
xnor U5436 (N_5436,N_1032,N_1844);
and U5437 (N_5437,N_853,N_1716);
nand U5438 (N_5438,N_682,N_1468);
or U5439 (N_5439,N_1240,N_2453);
or U5440 (N_5440,N_1443,N_1117);
xor U5441 (N_5441,N_1336,N_2912);
nand U5442 (N_5442,N_3059,N_1525);
or U5443 (N_5443,N_2568,N_1287);
nor U5444 (N_5444,N_674,N_1861);
or U5445 (N_5445,N_2974,N_2105);
nor U5446 (N_5446,N_410,N_289);
nor U5447 (N_5447,N_2443,N_2101);
and U5448 (N_5448,N_2927,N_2406);
xnor U5449 (N_5449,N_720,N_127);
nor U5450 (N_5450,N_448,N_2535);
and U5451 (N_5451,N_361,N_736);
or U5452 (N_5452,N_157,N_1585);
nor U5453 (N_5453,N_2702,N_176);
or U5454 (N_5454,N_1500,N_1015);
and U5455 (N_5455,N_434,N_4);
nand U5456 (N_5456,N_1581,N_2665);
or U5457 (N_5457,N_1195,N_220);
or U5458 (N_5458,N_464,N_208);
nand U5459 (N_5459,N_1405,N_171);
or U5460 (N_5460,N_2263,N_3045);
nor U5461 (N_5461,N_2404,N_1292);
and U5462 (N_5462,N_2896,N_502);
and U5463 (N_5463,N_1633,N_797);
or U5464 (N_5464,N_126,N_2208);
or U5465 (N_5465,N_2737,N_532);
xnor U5466 (N_5466,N_2413,N_2509);
and U5467 (N_5467,N_2544,N_1469);
or U5468 (N_5468,N_2354,N_1081);
or U5469 (N_5469,N_1477,N_1633);
nand U5470 (N_5470,N_921,N_2793);
or U5471 (N_5471,N_1298,N_2260);
and U5472 (N_5472,N_549,N_1016);
nor U5473 (N_5473,N_2592,N_3123);
nand U5474 (N_5474,N_644,N_2714);
or U5475 (N_5475,N_3055,N_1459);
nand U5476 (N_5476,N_2894,N_702);
and U5477 (N_5477,N_651,N_2307);
nor U5478 (N_5478,N_2224,N_576);
or U5479 (N_5479,N_2230,N_256);
or U5480 (N_5480,N_746,N_2007);
xor U5481 (N_5481,N_111,N_1809);
nand U5482 (N_5482,N_1585,N_2486);
and U5483 (N_5483,N_374,N_2);
and U5484 (N_5484,N_2635,N_2327);
or U5485 (N_5485,N_1976,N_1348);
nand U5486 (N_5486,N_1760,N_2220);
nor U5487 (N_5487,N_899,N_636);
nand U5488 (N_5488,N_288,N_2720);
and U5489 (N_5489,N_1325,N_3003);
nand U5490 (N_5490,N_189,N_1637);
or U5491 (N_5491,N_2304,N_2198);
and U5492 (N_5492,N_135,N_869);
and U5493 (N_5493,N_450,N_1061);
and U5494 (N_5494,N_250,N_2921);
xnor U5495 (N_5495,N_846,N_1588);
nor U5496 (N_5496,N_1773,N_2269);
or U5497 (N_5497,N_2620,N_946);
nand U5498 (N_5498,N_1158,N_2180);
nor U5499 (N_5499,N_856,N_2253);
or U5500 (N_5500,N_113,N_2546);
nor U5501 (N_5501,N_1850,N_2798);
or U5502 (N_5502,N_2067,N_839);
or U5503 (N_5503,N_959,N_803);
nand U5504 (N_5504,N_666,N_1902);
xnor U5505 (N_5505,N_2311,N_1563);
and U5506 (N_5506,N_1694,N_2025);
nor U5507 (N_5507,N_1730,N_2257);
and U5508 (N_5508,N_546,N_2685);
or U5509 (N_5509,N_1477,N_2324);
nor U5510 (N_5510,N_212,N_2650);
nand U5511 (N_5511,N_2222,N_2621);
and U5512 (N_5512,N_2616,N_2761);
nor U5513 (N_5513,N_1423,N_1521);
nor U5514 (N_5514,N_1112,N_1691);
nor U5515 (N_5515,N_2509,N_1505);
nand U5516 (N_5516,N_2080,N_1361);
and U5517 (N_5517,N_2721,N_671);
and U5518 (N_5518,N_2487,N_1765);
nand U5519 (N_5519,N_465,N_299);
or U5520 (N_5520,N_2122,N_1543);
nor U5521 (N_5521,N_689,N_1545);
nor U5522 (N_5522,N_1850,N_213);
or U5523 (N_5523,N_1474,N_649);
nand U5524 (N_5524,N_1578,N_2644);
nand U5525 (N_5525,N_1189,N_2162);
and U5526 (N_5526,N_1055,N_198);
xnor U5527 (N_5527,N_693,N_352);
xor U5528 (N_5528,N_304,N_898);
nor U5529 (N_5529,N_2611,N_2336);
nand U5530 (N_5530,N_3069,N_2417);
or U5531 (N_5531,N_2693,N_1297);
or U5532 (N_5532,N_594,N_158);
nand U5533 (N_5533,N_2407,N_1817);
nor U5534 (N_5534,N_1799,N_1670);
or U5535 (N_5535,N_1087,N_2972);
and U5536 (N_5536,N_8,N_2616);
and U5537 (N_5537,N_1497,N_3094);
nand U5538 (N_5538,N_3078,N_1341);
nand U5539 (N_5539,N_560,N_2183);
nand U5540 (N_5540,N_905,N_215);
xor U5541 (N_5541,N_2158,N_1264);
or U5542 (N_5542,N_796,N_2931);
or U5543 (N_5543,N_500,N_171);
nand U5544 (N_5544,N_3008,N_104);
nand U5545 (N_5545,N_1339,N_2208);
or U5546 (N_5546,N_2638,N_1362);
nand U5547 (N_5547,N_2300,N_2883);
nand U5548 (N_5548,N_2869,N_620);
and U5549 (N_5549,N_2113,N_672);
nand U5550 (N_5550,N_2938,N_1191);
nand U5551 (N_5551,N_248,N_2074);
nand U5552 (N_5552,N_533,N_1437);
nor U5553 (N_5553,N_1853,N_1168);
and U5554 (N_5554,N_419,N_54);
xnor U5555 (N_5555,N_2339,N_2535);
or U5556 (N_5556,N_1751,N_58);
nor U5557 (N_5557,N_2141,N_225);
nor U5558 (N_5558,N_1326,N_518);
nand U5559 (N_5559,N_2429,N_1722);
nand U5560 (N_5560,N_2945,N_372);
nand U5561 (N_5561,N_1292,N_1350);
xor U5562 (N_5562,N_55,N_1819);
and U5563 (N_5563,N_731,N_2514);
nand U5564 (N_5564,N_1872,N_1349);
and U5565 (N_5565,N_626,N_2238);
and U5566 (N_5566,N_449,N_2395);
or U5567 (N_5567,N_1910,N_3067);
and U5568 (N_5568,N_542,N_334);
or U5569 (N_5569,N_1676,N_666);
or U5570 (N_5570,N_72,N_1856);
and U5571 (N_5571,N_3019,N_3066);
nor U5572 (N_5572,N_1899,N_2011);
xnor U5573 (N_5573,N_2253,N_114);
and U5574 (N_5574,N_62,N_836);
nor U5575 (N_5575,N_2776,N_2433);
and U5576 (N_5576,N_3010,N_2672);
or U5577 (N_5577,N_1281,N_1373);
or U5578 (N_5578,N_470,N_2308);
and U5579 (N_5579,N_891,N_1264);
and U5580 (N_5580,N_1835,N_698);
and U5581 (N_5581,N_2186,N_746);
or U5582 (N_5582,N_1909,N_2247);
nor U5583 (N_5583,N_1516,N_159);
nand U5584 (N_5584,N_1061,N_1828);
xor U5585 (N_5585,N_3124,N_2173);
nor U5586 (N_5586,N_768,N_1110);
nand U5587 (N_5587,N_2317,N_3116);
xnor U5588 (N_5588,N_1656,N_230);
or U5589 (N_5589,N_994,N_1999);
and U5590 (N_5590,N_1977,N_545);
nor U5591 (N_5591,N_1403,N_2273);
nor U5592 (N_5592,N_1121,N_2344);
or U5593 (N_5593,N_2224,N_1731);
nor U5594 (N_5594,N_2979,N_1469);
or U5595 (N_5595,N_1035,N_1560);
nand U5596 (N_5596,N_230,N_1151);
and U5597 (N_5597,N_2229,N_550);
and U5598 (N_5598,N_472,N_39);
nor U5599 (N_5599,N_791,N_646);
and U5600 (N_5600,N_2614,N_2010);
nand U5601 (N_5601,N_1009,N_2887);
nor U5602 (N_5602,N_2456,N_522);
nor U5603 (N_5603,N_2943,N_2703);
and U5604 (N_5604,N_2803,N_1165);
or U5605 (N_5605,N_599,N_1587);
nand U5606 (N_5606,N_1328,N_340);
and U5607 (N_5607,N_2119,N_1243);
nand U5608 (N_5608,N_1291,N_2264);
nand U5609 (N_5609,N_2373,N_1722);
nand U5610 (N_5610,N_1633,N_1163);
nand U5611 (N_5611,N_1462,N_3001);
nor U5612 (N_5612,N_2739,N_775);
nor U5613 (N_5613,N_776,N_2596);
and U5614 (N_5614,N_604,N_2405);
xor U5615 (N_5615,N_2448,N_2125);
and U5616 (N_5616,N_2330,N_1459);
or U5617 (N_5617,N_785,N_1086);
nor U5618 (N_5618,N_1189,N_2629);
and U5619 (N_5619,N_2411,N_1034);
nand U5620 (N_5620,N_1576,N_2445);
or U5621 (N_5621,N_320,N_722);
nor U5622 (N_5622,N_2150,N_628);
nor U5623 (N_5623,N_1252,N_1318);
xor U5624 (N_5624,N_1497,N_1971);
and U5625 (N_5625,N_321,N_1332);
nand U5626 (N_5626,N_497,N_363);
xor U5627 (N_5627,N_1606,N_277);
xnor U5628 (N_5628,N_253,N_540);
and U5629 (N_5629,N_2969,N_2613);
and U5630 (N_5630,N_1075,N_2790);
nor U5631 (N_5631,N_1597,N_1853);
nor U5632 (N_5632,N_1999,N_2381);
nand U5633 (N_5633,N_446,N_483);
or U5634 (N_5634,N_2377,N_1367);
or U5635 (N_5635,N_607,N_474);
or U5636 (N_5636,N_1622,N_2694);
or U5637 (N_5637,N_360,N_1000);
nand U5638 (N_5638,N_2281,N_1325);
or U5639 (N_5639,N_961,N_2206);
nand U5640 (N_5640,N_1825,N_1625);
nand U5641 (N_5641,N_397,N_1502);
nand U5642 (N_5642,N_2607,N_1130);
nand U5643 (N_5643,N_2234,N_2525);
nand U5644 (N_5644,N_2764,N_2854);
nand U5645 (N_5645,N_725,N_2527);
nand U5646 (N_5646,N_1889,N_2958);
and U5647 (N_5647,N_1332,N_1145);
and U5648 (N_5648,N_1769,N_2924);
nand U5649 (N_5649,N_1618,N_459);
and U5650 (N_5650,N_1838,N_2374);
nor U5651 (N_5651,N_640,N_2281);
or U5652 (N_5652,N_2829,N_2526);
nor U5653 (N_5653,N_439,N_2630);
and U5654 (N_5654,N_1238,N_13);
nand U5655 (N_5655,N_1119,N_522);
nor U5656 (N_5656,N_299,N_2362);
nand U5657 (N_5657,N_250,N_903);
nand U5658 (N_5658,N_2129,N_1830);
nor U5659 (N_5659,N_2755,N_1447);
or U5660 (N_5660,N_2600,N_2227);
or U5661 (N_5661,N_1133,N_928);
nand U5662 (N_5662,N_3069,N_2743);
nand U5663 (N_5663,N_2356,N_1553);
and U5664 (N_5664,N_2650,N_82);
nand U5665 (N_5665,N_652,N_2653);
or U5666 (N_5666,N_325,N_2900);
and U5667 (N_5667,N_1411,N_758);
and U5668 (N_5668,N_1925,N_1579);
and U5669 (N_5669,N_2594,N_2373);
nand U5670 (N_5670,N_1871,N_1295);
or U5671 (N_5671,N_2789,N_352);
or U5672 (N_5672,N_2605,N_252);
or U5673 (N_5673,N_2992,N_1613);
nor U5674 (N_5674,N_2623,N_1913);
and U5675 (N_5675,N_405,N_2965);
nor U5676 (N_5676,N_535,N_1885);
and U5677 (N_5677,N_1233,N_2017);
and U5678 (N_5678,N_3001,N_1880);
nand U5679 (N_5679,N_68,N_2300);
xnor U5680 (N_5680,N_1410,N_552);
or U5681 (N_5681,N_2383,N_1199);
and U5682 (N_5682,N_333,N_2845);
and U5683 (N_5683,N_3022,N_445);
and U5684 (N_5684,N_2901,N_2518);
and U5685 (N_5685,N_2612,N_2882);
and U5686 (N_5686,N_1338,N_786);
nand U5687 (N_5687,N_1907,N_519);
or U5688 (N_5688,N_1300,N_628);
or U5689 (N_5689,N_1883,N_2917);
nor U5690 (N_5690,N_2302,N_2370);
and U5691 (N_5691,N_247,N_2332);
nand U5692 (N_5692,N_2725,N_1168);
nor U5693 (N_5693,N_1372,N_310);
nand U5694 (N_5694,N_1924,N_1743);
or U5695 (N_5695,N_2625,N_2485);
nor U5696 (N_5696,N_1268,N_2896);
nor U5697 (N_5697,N_854,N_2274);
nor U5698 (N_5698,N_1879,N_2897);
xor U5699 (N_5699,N_1352,N_2201);
or U5700 (N_5700,N_1109,N_2094);
or U5701 (N_5701,N_1505,N_1329);
and U5702 (N_5702,N_1809,N_169);
and U5703 (N_5703,N_2120,N_1033);
nand U5704 (N_5704,N_2119,N_792);
and U5705 (N_5705,N_292,N_3062);
and U5706 (N_5706,N_1259,N_2325);
nor U5707 (N_5707,N_1654,N_2210);
or U5708 (N_5708,N_1722,N_447);
or U5709 (N_5709,N_1099,N_2074);
or U5710 (N_5710,N_2448,N_1672);
nand U5711 (N_5711,N_1712,N_3076);
or U5712 (N_5712,N_141,N_2527);
nand U5713 (N_5713,N_2230,N_430);
nor U5714 (N_5714,N_2535,N_2106);
and U5715 (N_5715,N_331,N_2878);
and U5716 (N_5716,N_1803,N_2705);
nor U5717 (N_5717,N_1145,N_348);
nor U5718 (N_5718,N_1492,N_62);
or U5719 (N_5719,N_2617,N_1875);
and U5720 (N_5720,N_2583,N_2655);
xor U5721 (N_5721,N_1765,N_1619);
xor U5722 (N_5722,N_2743,N_1051);
xor U5723 (N_5723,N_3093,N_241);
xor U5724 (N_5724,N_739,N_665);
or U5725 (N_5725,N_2627,N_80);
and U5726 (N_5726,N_1487,N_1268);
and U5727 (N_5727,N_2722,N_2024);
xnor U5728 (N_5728,N_1072,N_617);
nand U5729 (N_5729,N_1817,N_371);
and U5730 (N_5730,N_1561,N_1286);
or U5731 (N_5731,N_1676,N_1413);
nor U5732 (N_5732,N_2785,N_2241);
or U5733 (N_5733,N_627,N_2121);
xnor U5734 (N_5734,N_2370,N_209);
nor U5735 (N_5735,N_182,N_1526);
or U5736 (N_5736,N_2473,N_2142);
nor U5737 (N_5737,N_1294,N_1136);
and U5738 (N_5738,N_1100,N_904);
and U5739 (N_5739,N_276,N_2135);
nor U5740 (N_5740,N_80,N_1679);
nand U5741 (N_5741,N_170,N_2684);
and U5742 (N_5742,N_609,N_1825);
or U5743 (N_5743,N_2806,N_1376);
nor U5744 (N_5744,N_456,N_352);
or U5745 (N_5745,N_271,N_345);
nand U5746 (N_5746,N_1377,N_2725);
nor U5747 (N_5747,N_1961,N_2320);
and U5748 (N_5748,N_240,N_1283);
nor U5749 (N_5749,N_2,N_1183);
nor U5750 (N_5750,N_3094,N_1112);
or U5751 (N_5751,N_1784,N_2653);
nor U5752 (N_5752,N_2195,N_1865);
or U5753 (N_5753,N_2805,N_2811);
and U5754 (N_5754,N_2781,N_2152);
and U5755 (N_5755,N_1289,N_1259);
and U5756 (N_5756,N_1611,N_961);
nor U5757 (N_5757,N_1503,N_1531);
xnor U5758 (N_5758,N_279,N_1663);
and U5759 (N_5759,N_2746,N_1671);
nand U5760 (N_5760,N_1906,N_252);
xnor U5761 (N_5761,N_472,N_325);
and U5762 (N_5762,N_2989,N_311);
or U5763 (N_5763,N_458,N_1783);
and U5764 (N_5764,N_341,N_171);
nor U5765 (N_5765,N_2162,N_1352);
or U5766 (N_5766,N_1193,N_2739);
xor U5767 (N_5767,N_3114,N_2644);
nand U5768 (N_5768,N_2042,N_2779);
and U5769 (N_5769,N_2162,N_2455);
nor U5770 (N_5770,N_2232,N_1931);
or U5771 (N_5771,N_2512,N_3008);
nand U5772 (N_5772,N_214,N_425);
or U5773 (N_5773,N_49,N_542);
xnor U5774 (N_5774,N_111,N_715);
and U5775 (N_5775,N_1052,N_3028);
nand U5776 (N_5776,N_937,N_1870);
xor U5777 (N_5777,N_1953,N_1810);
and U5778 (N_5778,N_155,N_674);
and U5779 (N_5779,N_1450,N_2307);
nor U5780 (N_5780,N_2105,N_2598);
or U5781 (N_5781,N_2653,N_1381);
nor U5782 (N_5782,N_2610,N_127);
and U5783 (N_5783,N_918,N_870);
or U5784 (N_5784,N_217,N_1046);
and U5785 (N_5785,N_1689,N_1223);
xor U5786 (N_5786,N_2689,N_1488);
nor U5787 (N_5787,N_1383,N_1281);
or U5788 (N_5788,N_83,N_285);
and U5789 (N_5789,N_1378,N_2406);
or U5790 (N_5790,N_569,N_628);
and U5791 (N_5791,N_2099,N_2755);
nand U5792 (N_5792,N_2329,N_95);
or U5793 (N_5793,N_454,N_1351);
nand U5794 (N_5794,N_2901,N_90);
or U5795 (N_5795,N_2858,N_1865);
nor U5796 (N_5796,N_2134,N_3037);
xnor U5797 (N_5797,N_937,N_1710);
and U5798 (N_5798,N_2952,N_1845);
nor U5799 (N_5799,N_2758,N_2478);
nand U5800 (N_5800,N_1105,N_2432);
nor U5801 (N_5801,N_2979,N_2670);
and U5802 (N_5802,N_1007,N_753);
nor U5803 (N_5803,N_2130,N_2968);
nor U5804 (N_5804,N_2720,N_1211);
nor U5805 (N_5805,N_1318,N_3113);
nor U5806 (N_5806,N_80,N_2960);
nor U5807 (N_5807,N_2786,N_1073);
or U5808 (N_5808,N_2837,N_2988);
nor U5809 (N_5809,N_1119,N_1856);
or U5810 (N_5810,N_780,N_359);
nand U5811 (N_5811,N_2278,N_2019);
or U5812 (N_5812,N_695,N_1);
nor U5813 (N_5813,N_950,N_111);
and U5814 (N_5814,N_1962,N_1475);
nor U5815 (N_5815,N_1281,N_1748);
xor U5816 (N_5816,N_1599,N_2607);
or U5817 (N_5817,N_737,N_2083);
or U5818 (N_5818,N_2870,N_673);
xor U5819 (N_5819,N_2899,N_1368);
and U5820 (N_5820,N_2534,N_1169);
nand U5821 (N_5821,N_373,N_3074);
and U5822 (N_5822,N_594,N_1885);
or U5823 (N_5823,N_715,N_1582);
nor U5824 (N_5824,N_1749,N_1319);
and U5825 (N_5825,N_2804,N_398);
nand U5826 (N_5826,N_2945,N_1563);
nand U5827 (N_5827,N_36,N_82);
and U5828 (N_5828,N_3100,N_2334);
or U5829 (N_5829,N_1101,N_2488);
nor U5830 (N_5830,N_2752,N_372);
nor U5831 (N_5831,N_809,N_2933);
nand U5832 (N_5832,N_401,N_2696);
and U5833 (N_5833,N_178,N_1734);
and U5834 (N_5834,N_2363,N_2785);
or U5835 (N_5835,N_1385,N_2786);
nand U5836 (N_5836,N_2666,N_2076);
and U5837 (N_5837,N_2676,N_1532);
xor U5838 (N_5838,N_714,N_1149);
and U5839 (N_5839,N_1039,N_1316);
xor U5840 (N_5840,N_194,N_1735);
nand U5841 (N_5841,N_2564,N_59);
nor U5842 (N_5842,N_72,N_2540);
or U5843 (N_5843,N_207,N_797);
and U5844 (N_5844,N_960,N_2294);
or U5845 (N_5845,N_2357,N_212);
or U5846 (N_5846,N_190,N_1260);
or U5847 (N_5847,N_1378,N_1038);
or U5848 (N_5848,N_1919,N_1475);
and U5849 (N_5849,N_601,N_1423);
or U5850 (N_5850,N_868,N_1027);
nand U5851 (N_5851,N_1698,N_232);
and U5852 (N_5852,N_1531,N_1414);
and U5853 (N_5853,N_247,N_2676);
nor U5854 (N_5854,N_2641,N_1036);
and U5855 (N_5855,N_1369,N_1663);
and U5856 (N_5856,N_112,N_462);
and U5857 (N_5857,N_1054,N_2468);
nand U5858 (N_5858,N_2835,N_1554);
xor U5859 (N_5859,N_2298,N_726);
or U5860 (N_5860,N_321,N_792);
and U5861 (N_5861,N_1140,N_1103);
nor U5862 (N_5862,N_143,N_938);
nor U5863 (N_5863,N_267,N_922);
nand U5864 (N_5864,N_2744,N_2886);
xnor U5865 (N_5865,N_1828,N_1060);
and U5866 (N_5866,N_2371,N_2760);
nand U5867 (N_5867,N_1056,N_1782);
and U5868 (N_5868,N_1072,N_2632);
nand U5869 (N_5869,N_759,N_1577);
nand U5870 (N_5870,N_1699,N_2580);
nand U5871 (N_5871,N_1373,N_1471);
nand U5872 (N_5872,N_1220,N_272);
nand U5873 (N_5873,N_3079,N_760);
nor U5874 (N_5874,N_1367,N_1472);
or U5875 (N_5875,N_2985,N_712);
nor U5876 (N_5876,N_1673,N_3064);
nor U5877 (N_5877,N_1724,N_628);
nand U5878 (N_5878,N_413,N_2172);
nor U5879 (N_5879,N_1974,N_2546);
nand U5880 (N_5880,N_2832,N_669);
nand U5881 (N_5881,N_2019,N_676);
nor U5882 (N_5882,N_172,N_2341);
or U5883 (N_5883,N_2746,N_1788);
nor U5884 (N_5884,N_1081,N_970);
nor U5885 (N_5885,N_955,N_2877);
and U5886 (N_5886,N_1579,N_2527);
nand U5887 (N_5887,N_1875,N_2322);
xor U5888 (N_5888,N_1222,N_2096);
or U5889 (N_5889,N_1068,N_552);
and U5890 (N_5890,N_1602,N_1540);
or U5891 (N_5891,N_397,N_2162);
or U5892 (N_5892,N_2126,N_1274);
and U5893 (N_5893,N_2217,N_1036);
nor U5894 (N_5894,N_1979,N_840);
nand U5895 (N_5895,N_413,N_2001);
nor U5896 (N_5896,N_1801,N_414);
or U5897 (N_5897,N_1159,N_495);
nand U5898 (N_5898,N_2156,N_2187);
or U5899 (N_5899,N_494,N_924);
nand U5900 (N_5900,N_2881,N_112);
and U5901 (N_5901,N_1150,N_1686);
xor U5902 (N_5902,N_308,N_2191);
and U5903 (N_5903,N_2701,N_1269);
nand U5904 (N_5904,N_752,N_2059);
or U5905 (N_5905,N_783,N_1223);
and U5906 (N_5906,N_896,N_3105);
or U5907 (N_5907,N_1324,N_1224);
nor U5908 (N_5908,N_2688,N_2394);
or U5909 (N_5909,N_1474,N_777);
nand U5910 (N_5910,N_1454,N_1260);
or U5911 (N_5911,N_813,N_622);
nor U5912 (N_5912,N_158,N_1669);
and U5913 (N_5913,N_180,N_1953);
nor U5914 (N_5914,N_2480,N_2163);
and U5915 (N_5915,N_275,N_3065);
xnor U5916 (N_5916,N_353,N_508);
xnor U5917 (N_5917,N_574,N_941);
nor U5918 (N_5918,N_928,N_2975);
and U5919 (N_5919,N_2571,N_2317);
nor U5920 (N_5920,N_123,N_2119);
and U5921 (N_5921,N_2281,N_2921);
or U5922 (N_5922,N_1824,N_931);
xnor U5923 (N_5923,N_1477,N_543);
and U5924 (N_5924,N_445,N_14);
nor U5925 (N_5925,N_2473,N_2799);
or U5926 (N_5926,N_466,N_1947);
and U5927 (N_5927,N_799,N_103);
nor U5928 (N_5928,N_2975,N_1519);
or U5929 (N_5929,N_2395,N_2486);
nor U5930 (N_5930,N_1798,N_46);
nor U5931 (N_5931,N_223,N_891);
or U5932 (N_5932,N_3088,N_2611);
or U5933 (N_5933,N_2511,N_2432);
xnor U5934 (N_5934,N_863,N_2209);
nand U5935 (N_5935,N_1803,N_3004);
or U5936 (N_5936,N_1450,N_403);
nand U5937 (N_5937,N_296,N_837);
nand U5938 (N_5938,N_1438,N_1740);
nand U5939 (N_5939,N_1025,N_2273);
xor U5940 (N_5940,N_1537,N_2085);
nor U5941 (N_5941,N_1014,N_40);
nor U5942 (N_5942,N_2161,N_2615);
or U5943 (N_5943,N_1353,N_992);
xnor U5944 (N_5944,N_2480,N_2697);
xnor U5945 (N_5945,N_1226,N_1267);
xor U5946 (N_5946,N_801,N_2488);
nor U5947 (N_5947,N_889,N_3107);
or U5948 (N_5948,N_674,N_1544);
xnor U5949 (N_5949,N_645,N_2483);
or U5950 (N_5950,N_2280,N_1206);
nand U5951 (N_5951,N_1266,N_2586);
nor U5952 (N_5952,N_1424,N_3104);
nand U5953 (N_5953,N_1400,N_2755);
xor U5954 (N_5954,N_2321,N_7);
and U5955 (N_5955,N_602,N_1044);
or U5956 (N_5956,N_883,N_1671);
or U5957 (N_5957,N_664,N_1142);
and U5958 (N_5958,N_2572,N_2570);
nand U5959 (N_5959,N_2135,N_534);
nand U5960 (N_5960,N_474,N_176);
nor U5961 (N_5961,N_3007,N_2352);
and U5962 (N_5962,N_1336,N_980);
nand U5963 (N_5963,N_973,N_2364);
or U5964 (N_5964,N_2844,N_2409);
or U5965 (N_5965,N_1021,N_1638);
nand U5966 (N_5966,N_2484,N_261);
nand U5967 (N_5967,N_2546,N_1125);
nand U5968 (N_5968,N_2557,N_782);
nand U5969 (N_5969,N_2084,N_2493);
and U5970 (N_5970,N_2046,N_2761);
or U5971 (N_5971,N_646,N_868);
or U5972 (N_5972,N_1809,N_527);
nand U5973 (N_5973,N_2382,N_2792);
nand U5974 (N_5974,N_2436,N_642);
or U5975 (N_5975,N_2189,N_519);
nor U5976 (N_5976,N_2119,N_2327);
nand U5977 (N_5977,N_361,N_2255);
xnor U5978 (N_5978,N_1977,N_783);
or U5979 (N_5979,N_361,N_1126);
and U5980 (N_5980,N_1521,N_3098);
nor U5981 (N_5981,N_2852,N_1653);
or U5982 (N_5982,N_1647,N_1766);
and U5983 (N_5983,N_2969,N_838);
or U5984 (N_5984,N_512,N_1318);
nor U5985 (N_5985,N_1763,N_2992);
and U5986 (N_5986,N_1847,N_1093);
nor U5987 (N_5987,N_493,N_220);
nor U5988 (N_5988,N_1758,N_452);
or U5989 (N_5989,N_591,N_3072);
and U5990 (N_5990,N_2932,N_1055);
nand U5991 (N_5991,N_1220,N_1703);
nor U5992 (N_5992,N_429,N_837);
nand U5993 (N_5993,N_545,N_2456);
nor U5994 (N_5994,N_2369,N_2191);
and U5995 (N_5995,N_979,N_2080);
xnor U5996 (N_5996,N_3098,N_1407);
or U5997 (N_5997,N_2019,N_313);
and U5998 (N_5998,N_50,N_456);
or U5999 (N_5999,N_181,N_1780);
xor U6000 (N_6000,N_3004,N_1647);
or U6001 (N_6001,N_2538,N_1961);
nor U6002 (N_6002,N_2982,N_3062);
or U6003 (N_6003,N_1806,N_506);
or U6004 (N_6004,N_487,N_2193);
nor U6005 (N_6005,N_2860,N_863);
nor U6006 (N_6006,N_135,N_2929);
or U6007 (N_6007,N_2322,N_1231);
nor U6008 (N_6008,N_1540,N_3100);
nor U6009 (N_6009,N_2734,N_2858);
nand U6010 (N_6010,N_2938,N_63);
xor U6011 (N_6011,N_1126,N_741);
and U6012 (N_6012,N_1086,N_2128);
nor U6013 (N_6013,N_700,N_871);
and U6014 (N_6014,N_65,N_176);
nand U6015 (N_6015,N_2990,N_2060);
nor U6016 (N_6016,N_2443,N_2905);
nand U6017 (N_6017,N_200,N_1312);
nor U6018 (N_6018,N_470,N_1667);
or U6019 (N_6019,N_3051,N_1997);
and U6020 (N_6020,N_642,N_2565);
and U6021 (N_6021,N_867,N_1432);
or U6022 (N_6022,N_2104,N_229);
or U6023 (N_6023,N_454,N_178);
xor U6024 (N_6024,N_134,N_2145);
and U6025 (N_6025,N_930,N_950);
nor U6026 (N_6026,N_853,N_2167);
nor U6027 (N_6027,N_1973,N_2079);
and U6028 (N_6028,N_1938,N_2388);
nor U6029 (N_6029,N_1875,N_943);
and U6030 (N_6030,N_3069,N_2578);
nor U6031 (N_6031,N_296,N_2371);
and U6032 (N_6032,N_1791,N_220);
nor U6033 (N_6033,N_709,N_2631);
nand U6034 (N_6034,N_1046,N_839);
or U6035 (N_6035,N_267,N_842);
and U6036 (N_6036,N_786,N_915);
nand U6037 (N_6037,N_1614,N_2671);
nand U6038 (N_6038,N_2624,N_2716);
or U6039 (N_6039,N_1015,N_1033);
and U6040 (N_6040,N_2409,N_2063);
and U6041 (N_6041,N_144,N_1489);
and U6042 (N_6042,N_3027,N_1438);
and U6043 (N_6043,N_1569,N_18);
or U6044 (N_6044,N_2037,N_2691);
or U6045 (N_6045,N_2482,N_1653);
and U6046 (N_6046,N_1779,N_698);
nand U6047 (N_6047,N_1206,N_1735);
nand U6048 (N_6048,N_2269,N_1692);
or U6049 (N_6049,N_2614,N_2163);
nand U6050 (N_6050,N_2775,N_1365);
or U6051 (N_6051,N_1329,N_1263);
xnor U6052 (N_6052,N_606,N_785);
nor U6053 (N_6053,N_1734,N_1305);
nand U6054 (N_6054,N_2657,N_709);
and U6055 (N_6055,N_2029,N_1282);
xor U6056 (N_6056,N_1366,N_909);
or U6057 (N_6057,N_2549,N_765);
nor U6058 (N_6058,N_996,N_420);
nand U6059 (N_6059,N_333,N_247);
and U6060 (N_6060,N_1464,N_2773);
and U6061 (N_6061,N_244,N_81);
and U6062 (N_6062,N_2982,N_3054);
nand U6063 (N_6063,N_37,N_3033);
xnor U6064 (N_6064,N_676,N_52);
nand U6065 (N_6065,N_2459,N_2071);
nand U6066 (N_6066,N_1773,N_1033);
or U6067 (N_6067,N_701,N_1539);
nand U6068 (N_6068,N_2484,N_1930);
nor U6069 (N_6069,N_1594,N_1444);
nand U6070 (N_6070,N_1030,N_1444);
or U6071 (N_6071,N_2195,N_1261);
nor U6072 (N_6072,N_1662,N_19);
or U6073 (N_6073,N_1430,N_2200);
or U6074 (N_6074,N_1253,N_135);
and U6075 (N_6075,N_67,N_421);
or U6076 (N_6076,N_1139,N_3090);
nand U6077 (N_6077,N_828,N_614);
xnor U6078 (N_6078,N_958,N_2174);
and U6079 (N_6079,N_1500,N_1654);
and U6080 (N_6080,N_22,N_1940);
xor U6081 (N_6081,N_1971,N_1414);
nand U6082 (N_6082,N_568,N_495);
and U6083 (N_6083,N_1504,N_1720);
xor U6084 (N_6084,N_1348,N_271);
xnor U6085 (N_6085,N_2186,N_1178);
nand U6086 (N_6086,N_1692,N_1965);
or U6087 (N_6087,N_2871,N_1259);
nor U6088 (N_6088,N_783,N_1009);
and U6089 (N_6089,N_2632,N_593);
xnor U6090 (N_6090,N_1977,N_2037);
xor U6091 (N_6091,N_3077,N_603);
nor U6092 (N_6092,N_2811,N_132);
and U6093 (N_6093,N_2779,N_2244);
nor U6094 (N_6094,N_1631,N_253);
and U6095 (N_6095,N_1250,N_1727);
nor U6096 (N_6096,N_2404,N_993);
and U6097 (N_6097,N_2652,N_1551);
nor U6098 (N_6098,N_597,N_2422);
and U6099 (N_6099,N_1216,N_25);
xnor U6100 (N_6100,N_1030,N_2407);
and U6101 (N_6101,N_2504,N_1744);
and U6102 (N_6102,N_1388,N_2084);
and U6103 (N_6103,N_1470,N_2160);
and U6104 (N_6104,N_999,N_2597);
and U6105 (N_6105,N_1943,N_248);
nand U6106 (N_6106,N_1866,N_389);
or U6107 (N_6107,N_2806,N_338);
nand U6108 (N_6108,N_2637,N_55);
or U6109 (N_6109,N_2709,N_906);
or U6110 (N_6110,N_78,N_910);
nand U6111 (N_6111,N_2605,N_1172);
or U6112 (N_6112,N_1115,N_1181);
and U6113 (N_6113,N_1198,N_1952);
nor U6114 (N_6114,N_2074,N_2729);
and U6115 (N_6115,N_1307,N_189);
nand U6116 (N_6116,N_483,N_1787);
nor U6117 (N_6117,N_1945,N_1519);
and U6118 (N_6118,N_31,N_2640);
and U6119 (N_6119,N_2751,N_1894);
nor U6120 (N_6120,N_396,N_719);
or U6121 (N_6121,N_386,N_879);
nor U6122 (N_6122,N_2381,N_635);
nand U6123 (N_6123,N_2191,N_2789);
xor U6124 (N_6124,N_1999,N_1126);
nor U6125 (N_6125,N_1685,N_2289);
or U6126 (N_6126,N_1121,N_924);
nor U6127 (N_6127,N_2485,N_1359);
nor U6128 (N_6128,N_2994,N_424);
nor U6129 (N_6129,N_2238,N_1126);
xor U6130 (N_6130,N_127,N_2359);
nor U6131 (N_6131,N_821,N_606);
nor U6132 (N_6132,N_1168,N_3055);
nand U6133 (N_6133,N_2349,N_2497);
and U6134 (N_6134,N_3068,N_182);
xor U6135 (N_6135,N_944,N_1046);
xnor U6136 (N_6136,N_1516,N_532);
and U6137 (N_6137,N_21,N_364);
or U6138 (N_6138,N_1708,N_2362);
or U6139 (N_6139,N_2459,N_2268);
or U6140 (N_6140,N_1096,N_2082);
xor U6141 (N_6141,N_2869,N_1214);
xnor U6142 (N_6142,N_1135,N_1869);
and U6143 (N_6143,N_1811,N_991);
nand U6144 (N_6144,N_2448,N_778);
or U6145 (N_6145,N_2173,N_378);
and U6146 (N_6146,N_876,N_921);
or U6147 (N_6147,N_372,N_2861);
or U6148 (N_6148,N_648,N_2045);
xor U6149 (N_6149,N_1078,N_2158);
xnor U6150 (N_6150,N_2820,N_1347);
xor U6151 (N_6151,N_3088,N_2163);
nand U6152 (N_6152,N_1305,N_1561);
and U6153 (N_6153,N_2069,N_2029);
nor U6154 (N_6154,N_2206,N_938);
nand U6155 (N_6155,N_1302,N_2493);
or U6156 (N_6156,N_2095,N_187);
and U6157 (N_6157,N_1931,N_458);
xor U6158 (N_6158,N_391,N_2481);
nand U6159 (N_6159,N_1140,N_2189);
nor U6160 (N_6160,N_511,N_606);
xnor U6161 (N_6161,N_86,N_2920);
nor U6162 (N_6162,N_2526,N_953);
or U6163 (N_6163,N_1977,N_580);
or U6164 (N_6164,N_2485,N_1147);
or U6165 (N_6165,N_1130,N_1003);
nand U6166 (N_6166,N_2105,N_48);
xor U6167 (N_6167,N_2770,N_1487);
and U6168 (N_6168,N_1016,N_862);
nor U6169 (N_6169,N_1943,N_817);
or U6170 (N_6170,N_1820,N_168);
or U6171 (N_6171,N_2554,N_2602);
and U6172 (N_6172,N_3001,N_485);
nand U6173 (N_6173,N_519,N_2270);
nor U6174 (N_6174,N_2593,N_1015);
or U6175 (N_6175,N_3014,N_414);
nand U6176 (N_6176,N_2058,N_132);
nand U6177 (N_6177,N_882,N_1770);
nand U6178 (N_6178,N_199,N_2984);
or U6179 (N_6179,N_2095,N_1469);
and U6180 (N_6180,N_2501,N_2371);
nor U6181 (N_6181,N_2598,N_2401);
and U6182 (N_6182,N_2410,N_957);
or U6183 (N_6183,N_2580,N_2641);
or U6184 (N_6184,N_2250,N_2177);
nand U6185 (N_6185,N_2429,N_2068);
and U6186 (N_6186,N_2621,N_175);
nand U6187 (N_6187,N_2702,N_755);
nand U6188 (N_6188,N_2660,N_2815);
or U6189 (N_6189,N_1698,N_1661);
nor U6190 (N_6190,N_2147,N_1503);
and U6191 (N_6191,N_2341,N_1438);
nand U6192 (N_6192,N_1811,N_1169);
or U6193 (N_6193,N_1136,N_3117);
nor U6194 (N_6194,N_303,N_1345);
nand U6195 (N_6195,N_200,N_1091);
nor U6196 (N_6196,N_2642,N_2463);
nand U6197 (N_6197,N_475,N_486);
and U6198 (N_6198,N_1138,N_1388);
or U6199 (N_6199,N_2019,N_2491);
nor U6200 (N_6200,N_757,N_631);
nor U6201 (N_6201,N_2963,N_778);
or U6202 (N_6202,N_2105,N_2050);
or U6203 (N_6203,N_1573,N_426);
nor U6204 (N_6204,N_3094,N_1494);
xor U6205 (N_6205,N_668,N_1749);
and U6206 (N_6206,N_1563,N_1187);
or U6207 (N_6207,N_1820,N_1306);
nand U6208 (N_6208,N_1381,N_1890);
nor U6209 (N_6209,N_256,N_571);
nand U6210 (N_6210,N_2130,N_1900);
or U6211 (N_6211,N_2539,N_2507);
xnor U6212 (N_6212,N_3024,N_398);
nand U6213 (N_6213,N_2075,N_2951);
nand U6214 (N_6214,N_1422,N_587);
or U6215 (N_6215,N_2886,N_2354);
or U6216 (N_6216,N_2469,N_1370);
and U6217 (N_6217,N_225,N_1460);
nand U6218 (N_6218,N_1326,N_1863);
nor U6219 (N_6219,N_815,N_428);
xor U6220 (N_6220,N_2777,N_2062);
and U6221 (N_6221,N_2862,N_57);
and U6222 (N_6222,N_463,N_2988);
or U6223 (N_6223,N_1383,N_90);
nor U6224 (N_6224,N_70,N_2689);
or U6225 (N_6225,N_588,N_92);
xnor U6226 (N_6226,N_1383,N_971);
nand U6227 (N_6227,N_2590,N_218);
or U6228 (N_6228,N_218,N_2101);
nand U6229 (N_6229,N_3010,N_946);
nor U6230 (N_6230,N_1220,N_1177);
or U6231 (N_6231,N_1403,N_2143);
and U6232 (N_6232,N_1149,N_611);
nor U6233 (N_6233,N_949,N_2004);
nand U6234 (N_6234,N_2207,N_2857);
and U6235 (N_6235,N_2367,N_2724);
nor U6236 (N_6236,N_605,N_909);
nand U6237 (N_6237,N_3025,N_1922);
and U6238 (N_6238,N_786,N_1327);
or U6239 (N_6239,N_1757,N_2256);
nor U6240 (N_6240,N_2387,N_268);
xnor U6241 (N_6241,N_1300,N_1413);
or U6242 (N_6242,N_1055,N_1920);
xor U6243 (N_6243,N_1645,N_39);
and U6244 (N_6244,N_854,N_2760);
or U6245 (N_6245,N_1579,N_194);
nand U6246 (N_6246,N_775,N_1842);
and U6247 (N_6247,N_2673,N_2294);
and U6248 (N_6248,N_3097,N_202);
nor U6249 (N_6249,N_2299,N_1374);
or U6250 (N_6250,N_4995,N_3526);
or U6251 (N_6251,N_4989,N_5648);
or U6252 (N_6252,N_6195,N_5448);
or U6253 (N_6253,N_5328,N_5036);
and U6254 (N_6254,N_4045,N_3170);
nor U6255 (N_6255,N_6113,N_5654);
and U6256 (N_6256,N_3731,N_3367);
nor U6257 (N_6257,N_5830,N_4486);
or U6258 (N_6258,N_4612,N_3685);
nand U6259 (N_6259,N_5649,N_6078);
or U6260 (N_6260,N_5238,N_4571);
xnor U6261 (N_6261,N_5864,N_5829);
xnor U6262 (N_6262,N_5529,N_6147);
or U6263 (N_6263,N_5401,N_4850);
nor U6264 (N_6264,N_5091,N_5753);
nor U6265 (N_6265,N_3648,N_4716);
nor U6266 (N_6266,N_3505,N_4117);
nand U6267 (N_6267,N_6213,N_3424);
nor U6268 (N_6268,N_4355,N_5996);
and U6269 (N_6269,N_4519,N_3907);
or U6270 (N_6270,N_3352,N_5471);
or U6271 (N_6271,N_3711,N_6132);
nor U6272 (N_6272,N_3329,N_4199);
xor U6273 (N_6273,N_6084,N_5418);
xnor U6274 (N_6274,N_6107,N_6098);
and U6275 (N_6275,N_3607,N_6206);
nand U6276 (N_6276,N_4491,N_4668);
nor U6277 (N_6277,N_5114,N_3641);
or U6278 (N_6278,N_5916,N_3373);
nor U6279 (N_6279,N_6119,N_5509);
and U6280 (N_6280,N_3843,N_3776);
and U6281 (N_6281,N_3457,N_5889);
or U6282 (N_6282,N_4891,N_5852);
and U6283 (N_6283,N_5749,N_3873);
nand U6284 (N_6284,N_4903,N_5031);
and U6285 (N_6285,N_5914,N_6096);
and U6286 (N_6286,N_3328,N_5717);
nor U6287 (N_6287,N_5267,N_3800);
and U6288 (N_6288,N_3276,N_5050);
nand U6289 (N_6289,N_3626,N_5912);
xor U6290 (N_6290,N_4312,N_4569);
and U6291 (N_6291,N_3871,N_4804);
nor U6292 (N_6292,N_5883,N_3551);
and U6293 (N_6293,N_4391,N_4530);
or U6294 (N_6294,N_6011,N_3959);
or U6295 (N_6295,N_3847,N_5986);
or U6296 (N_6296,N_5508,N_5432);
nor U6297 (N_6297,N_3693,N_5604);
or U6298 (N_6298,N_3490,N_5952);
nor U6299 (N_6299,N_4548,N_3649);
nand U6300 (N_6300,N_4135,N_6022);
and U6301 (N_6301,N_4930,N_4229);
nor U6302 (N_6302,N_6235,N_3438);
and U6303 (N_6303,N_3804,N_4696);
or U6304 (N_6304,N_4921,N_4998);
and U6305 (N_6305,N_5246,N_5705);
nand U6306 (N_6306,N_4556,N_4823);
or U6307 (N_6307,N_3202,N_3310);
xnor U6308 (N_6308,N_3579,N_5668);
nor U6309 (N_6309,N_5940,N_4647);
nand U6310 (N_6310,N_3340,N_3857);
and U6311 (N_6311,N_3706,N_5278);
nand U6312 (N_6312,N_5924,N_4197);
and U6313 (N_6313,N_5728,N_4186);
or U6314 (N_6314,N_3998,N_4070);
or U6315 (N_6315,N_5547,N_6155);
nand U6316 (N_6316,N_4038,N_3391);
and U6317 (N_6317,N_3760,N_3627);
or U6318 (N_6318,N_5151,N_5707);
and U6319 (N_6319,N_3259,N_4590);
nor U6320 (N_6320,N_5299,N_4351);
nor U6321 (N_6321,N_5398,N_5186);
nor U6322 (N_6322,N_5195,N_4061);
nand U6323 (N_6323,N_4093,N_5569);
nand U6324 (N_6324,N_3159,N_5853);
or U6325 (N_6325,N_3495,N_4940);
or U6326 (N_6326,N_4410,N_3503);
xor U6327 (N_6327,N_6158,N_5546);
nor U6328 (N_6328,N_5202,N_4790);
nor U6329 (N_6329,N_5810,N_4177);
nor U6330 (N_6330,N_3617,N_3605);
nor U6331 (N_6331,N_3958,N_6072);
and U6332 (N_6332,N_4183,N_4568);
nor U6333 (N_6333,N_4015,N_5295);
nand U6334 (N_6334,N_5363,N_5866);
nor U6335 (N_6335,N_5500,N_4616);
xor U6336 (N_6336,N_4709,N_4623);
nand U6337 (N_6337,N_5727,N_4000);
and U6338 (N_6338,N_5170,N_3318);
or U6339 (N_6339,N_4832,N_5575);
nor U6340 (N_6340,N_3355,N_5780);
and U6341 (N_6341,N_6171,N_5785);
and U6342 (N_6342,N_3929,N_3566);
nor U6343 (N_6343,N_3307,N_4213);
xor U6344 (N_6344,N_6198,N_4599);
or U6345 (N_6345,N_3976,N_5906);
or U6346 (N_6346,N_4083,N_4439);
or U6347 (N_6347,N_4253,N_3395);
nand U6348 (N_6348,N_5157,N_4359);
nor U6349 (N_6349,N_5832,N_4985);
nor U6350 (N_6350,N_4110,N_5543);
or U6351 (N_6351,N_5870,N_4602);
nor U6352 (N_6352,N_4649,N_5112);
nor U6353 (N_6353,N_6057,N_6238);
nand U6354 (N_6354,N_6202,N_6153);
and U6355 (N_6355,N_3910,N_5488);
nand U6356 (N_6356,N_5739,N_4467);
or U6357 (N_6357,N_4248,N_3175);
nand U6358 (N_6358,N_5570,N_3813);
nand U6359 (N_6359,N_5066,N_5819);
nand U6360 (N_6360,N_4218,N_4763);
nand U6361 (N_6361,N_3981,N_4841);
nand U6362 (N_6362,N_5439,N_6149);
or U6363 (N_6363,N_4222,N_4095);
and U6364 (N_6364,N_6073,N_4446);
or U6365 (N_6365,N_4682,N_5937);
nand U6366 (N_6366,N_3768,N_4689);
nor U6367 (N_6367,N_5571,N_5352);
nor U6368 (N_6368,N_4484,N_4140);
and U6369 (N_6369,N_3619,N_3214);
nor U6370 (N_6370,N_5791,N_5153);
nand U6371 (N_6371,N_3348,N_5628);
nand U6372 (N_6372,N_4471,N_3745);
or U6373 (N_6373,N_4944,N_5752);
or U6374 (N_6374,N_4494,N_4040);
and U6375 (N_6375,N_4799,N_4288);
or U6376 (N_6376,N_5284,N_3577);
or U6377 (N_6377,N_5614,N_5100);
or U6378 (N_6378,N_4300,N_4963);
and U6379 (N_6379,N_4788,N_5169);
nor U6380 (N_6380,N_5121,N_4955);
nor U6381 (N_6381,N_3718,N_6001);
nand U6382 (N_6382,N_4969,N_3903);
and U6383 (N_6383,N_5213,N_3185);
nor U6384 (N_6384,N_5436,N_5927);
xor U6385 (N_6385,N_4711,N_3836);
xnor U6386 (N_6386,N_5068,N_4984);
and U6387 (N_6387,N_5878,N_3812);
nand U6388 (N_6388,N_3676,N_4683);
nand U6389 (N_6389,N_4736,N_5840);
nand U6390 (N_6390,N_4988,N_3927);
or U6391 (N_6391,N_5577,N_3137);
or U6392 (N_6392,N_3674,N_5960);
or U6393 (N_6393,N_3212,N_4806);
and U6394 (N_6394,N_3508,N_4585);
xor U6395 (N_6395,N_5959,N_3742);
nand U6396 (N_6396,N_3798,N_4113);
or U6397 (N_6397,N_4124,N_4746);
or U6398 (N_6398,N_3472,N_5079);
and U6399 (N_6399,N_3828,N_3824);
or U6400 (N_6400,N_5150,N_3523);
or U6401 (N_6401,N_5836,N_6112);
nand U6402 (N_6402,N_3858,N_4870);
nand U6403 (N_6403,N_5998,N_3967);
nor U6404 (N_6404,N_5722,N_4332);
and U6405 (N_6405,N_5601,N_5737);
nand U6406 (N_6406,N_4700,N_5913);
nand U6407 (N_6407,N_4348,N_4155);
nor U6408 (N_6408,N_3247,N_4094);
nor U6409 (N_6409,N_4295,N_5143);
and U6410 (N_6410,N_3404,N_3942);
xor U6411 (N_6411,N_3970,N_5592);
and U6412 (N_6412,N_3293,N_4800);
xor U6413 (N_6413,N_4915,N_5107);
xnor U6414 (N_6414,N_4503,N_5655);
or U6415 (N_6415,N_3298,N_3938);
or U6416 (N_6416,N_5474,N_5264);
and U6417 (N_6417,N_5414,N_6070);
nand U6418 (N_6418,N_5108,N_4693);
and U6419 (N_6419,N_4398,N_3385);
and U6420 (N_6420,N_4992,N_5220);
nand U6421 (N_6421,N_5227,N_4490);
nor U6422 (N_6422,N_3270,N_5392);
nand U6423 (N_6423,N_4150,N_5076);
and U6424 (N_6424,N_3721,N_4570);
and U6425 (N_6425,N_5233,N_4810);
and U6426 (N_6426,N_4836,N_3698);
and U6427 (N_6427,N_4239,N_4485);
or U6428 (N_6428,N_3628,N_5035);
and U6429 (N_6429,N_5751,N_3525);
xor U6430 (N_6430,N_4852,N_3468);
nand U6431 (N_6431,N_6244,N_5452);
nand U6432 (N_6432,N_3415,N_4655);
or U6433 (N_6433,N_5052,N_6047);
and U6434 (N_6434,N_4873,N_5973);
nor U6435 (N_6435,N_4115,N_4301);
nand U6436 (N_6436,N_5026,N_5833);
and U6437 (N_6437,N_5189,N_6225);
nand U6438 (N_6438,N_6043,N_3380);
or U6439 (N_6439,N_4376,N_5311);
or U6440 (N_6440,N_3941,N_3463);
nand U6441 (N_6441,N_5764,N_4077);
and U6442 (N_6442,N_4950,N_5908);
nor U6443 (N_6443,N_3728,N_3635);
or U6444 (N_6444,N_3912,N_3799);
nor U6445 (N_6445,N_3530,N_4691);
xnor U6446 (N_6446,N_3750,N_3849);
and U6447 (N_6447,N_5119,N_3889);
or U6448 (N_6448,N_4887,N_3286);
and U6449 (N_6449,N_5417,N_4851);
nor U6450 (N_6450,N_4418,N_4436);
and U6451 (N_6451,N_3229,N_5435);
nor U6452 (N_6452,N_5265,N_5967);
or U6453 (N_6453,N_3713,N_4378);
nor U6454 (N_6454,N_3216,N_5879);
and U6455 (N_6455,N_3834,N_4047);
or U6456 (N_6456,N_5095,N_3371);
nor U6457 (N_6457,N_4215,N_5535);
nand U6458 (N_6458,N_3213,N_5191);
nand U6459 (N_6459,N_5564,N_4712);
or U6460 (N_6460,N_5607,N_4803);
nand U6461 (N_6461,N_5097,N_5443);
nor U6462 (N_6462,N_4444,N_4920);
nor U6463 (N_6463,N_4327,N_6178);
and U6464 (N_6464,N_5362,N_4085);
nand U6465 (N_6465,N_4505,N_5963);
nand U6466 (N_6466,N_5083,N_5183);
nor U6467 (N_6467,N_3146,N_5797);
and U6468 (N_6468,N_5355,N_3336);
xnor U6469 (N_6469,N_3892,N_3994);
nor U6470 (N_6470,N_3547,N_3545);
xor U6471 (N_6471,N_4193,N_3261);
or U6472 (N_6472,N_6229,N_5877);
and U6473 (N_6473,N_3414,N_4660);
or U6474 (N_6474,N_3369,N_6191);
or U6475 (N_6475,N_6227,N_3399);
xnor U6476 (N_6476,N_3322,N_4564);
nor U6477 (N_6477,N_3955,N_5680);
and U6478 (N_6478,N_5816,N_4922);
xor U6479 (N_6479,N_4425,N_5742);
and U6480 (N_6480,N_5656,N_3152);
nor U6481 (N_6481,N_4194,N_5968);
nor U6482 (N_6482,N_3816,N_4086);
nor U6483 (N_6483,N_3471,N_3956);
nor U6484 (N_6484,N_4825,N_4837);
nand U6485 (N_6485,N_4948,N_5621);
nand U6486 (N_6486,N_5925,N_4914);
nand U6487 (N_6487,N_4573,N_4879);
and U6488 (N_6488,N_3499,N_3954);
and U6489 (N_6489,N_5622,N_3808);
or U6490 (N_6490,N_3492,N_4156);
and U6491 (N_6491,N_5433,N_3602);
or U6492 (N_6492,N_5402,N_4518);
xnor U6493 (N_6493,N_6049,N_4692);
and U6494 (N_6494,N_4235,N_4760);
or U6495 (N_6495,N_4596,N_6033);
nor U6496 (N_6496,N_5792,N_5982);
and U6497 (N_6497,N_3363,N_6060);
or U6498 (N_6498,N_4274,N_5812);
nor U6499 (N_6499,N_3507,N_3469);
or U6500 (N_6500,N_5702,N_3802);
or U6501 (N_6501,N_6136,N_3567);
and U6502 (N_6502,N_3256,N_3376);
xnor U6503 (N_6503,N_5568,N_4357);
nor U6504 (N_6504,N_4118,N_4091);
and U6505 (N_6505,N_4553,N_5905);
nand U6506 (N_6506,N_5451,N_6247);
or U6507 (N_6507,N_5788,N_5980);
or U6508 (N_6508,N_4328,N_5391);
nor U6509 (N_6509,N_4284,N_5673);
nand U6510 (N_6510,N_5958,N_5353);
nand U6511 (N_6511,N_4601,N_5842);
xor U6512 (N_6512,N_5007,N_5152);
nand U6513 (N_6513,N_3983,N_4149);
nand U6514 (N_6514,N_4438,N_5125);
nor U6515 (N_6515,N_5023,N_4924);
or U6516 (N_6516,N_5351,N_5505);
nand U6517 (N_6517,N_6005,N_5281);
nand U6518 (N_6518,N_3700,N_5336);
nand U6519 (N_6519,N_3925,N_5799);
xnor U6520 (N_6520,N_5693,N_6192);
nor U6521 (N_6521,N_3278,N_4014);
nor U6522 (N_6522,N_5422,N_5455);
and U6523 (N_6523,N_4515,N_4429);
nand U6524 (N_6524,N_5521,N_3444);
nand U6525 (N_6525,N_4326,N_4740);
and U6526 (N_6526,N_3207,N_3630);
and U6527 (N_6527,N_3921,N_5424);
nor U6528 (N_6528,N_4111,N_3274);
and U6529 (N_6529,N_5857,N_3156);
or U6530 (N_6530,N_3279,N_4058);
and U6531 (N_6531,N_6087,N_6125);
or U6532 (N_6532,N_5754,N_3429);
and U6533 (N_6533,N_3255,N_4982);
or U6534 (N_6534,N_3366,N_5054);
xnor U6535 (N_6535,N_6030,N_4893);
or U6536 (N_6536,N_3896,N_3143);
nor U6537 (N_6537,N_4258,N_4533);
nor U6538 (N_6538,N_3901,N_4659);
nand U6539 (N_6539,N_3829,N_3940);
or U6540 (N_6540,N_4853,N_4074);
xnor U6541 (N_6541,N_5969,N_4360);
and U6542 (N_6542,N_3634,N_5827);
or U6543 (N_6543,N_4170,N_4742);
nand U6544 (N_6544,N_5472,N_3754);
or U6545 (N_6545,N_4190,N_3879);
and U6546 (N_6546,N_5240,N_3263);
xor U6547 (N_6547,N_4002,N_3999);
nor U6548 (N_6548,N_4353,N_3647);
or U6549 (N_6549,N_6196,N_4007);
nor U6550 (N_6550,N_3194,N_3859);
xnor U6551 (N_6551,N_4771,N_3953);
nand U6552 (N_6552,N_6199,N_5122);
or U6553 (N_6553,N_6146,N_4130);
or U6554 (N_6554,N_4237,N_3864);
and U6555 (N_6555,N_5061,N_5863);
nor U6556 (N_6556,N_3260,N_5469);
and U6557 (N_6557,N_4703,N_4653);
nor U6558 (N_6558,N_5658,N_6120);
or U6559 (N_6559,N_3656,N_3947);
nor U6560 (N_6560,N_5588,N_4175);
nand U6561 (N_6561,N_3625,N_3632);
and U6562 (N_6562,N_4182,N_5217);
nand U6563 (N_6563,N_3769,N_5408);
nor U6564 (N_6564,N_3313,N_5104);
xnor U6565 (N_6565,N_4880,N_4428);
nor U6566 (N_6566,N_5364,N_3467);
nand U6567 (N_6567,N_5201,N_5550);
nor U6568 (N_6568,N_4377,N_5949);
nor U6569 (N_6569,N_5179,N_4939);
and U6570 (N_6570,N_3381,N_5389);
nor U6571 (N_6571,N_4902,N_5804);
nor U6572 (N_6572,N_6134,N_3362);
nor U6573 (N_6573,N_3480,N_3250);
nand U6574 (N_6574,N_3677,N_6215);
nand U6575 (N_6575,N_4534,N_3482);
xor U6576 (N_6576,N_4981,N_3494);
nand U6577 (N_6577,N_5706,N_4871);
and U6578 (N_6578,N_4666,N_3411);
and U6579 (N_6579,N_5997,N_5222);
or U6580 (N_6580,N_6089,N_5513);
and U6581 (N_6581,N_6203,N_5667);
or U6582 (N_6582,N_4004,N_4168);
and U6583 (N_6583,N_4911,N_3778);
nor U6584 (N_6584,N_5709,N_3218);
nand U6585 (N_6585,N_4042,N_3190);
nand U6586 (N_6586,N_3624,N_4162);
and U6587 (N_6587,N_5345,N_5897);
or U6588 (N_6588,N_5549,N_5946);
and U6589 (N_6589,N_5659,N_4999);
nor U6590 (N_6590,N_3756,N_3510);
nand U6591 (N_6591,N_3680,N_4480);
nand U6592 (N_6592,N_3631,N_4610);
or U6593 (N_6593,N_4629,N_5890);
nand U6594 (N_6594,N_5845,N_4122);
and U6595 (N_6595,N_5617,N_3403);
and U6596 (N_6596,N_5985,N_3845);
nor U6597 (N_6597,N_3794,N_3564);
or U6598 (N_6598,N_3345,N_4751);
xnor U6599 (N_6599,N_3868,N_3957);
or U6600 (N_6600,N_4392,N_4492);
and U6601 (N_6601,N_4977,N_4416);
or U6602 (N_6602,N_4039,N_3637);
or U6603 (N_6603,N_5479,N_4424);
or U6604 (N_6604,N_3127,N_6014);
nand U6605 (N_6605,N_5524,N_6248);
nand U6606 (N_6606,N_5239,N_5361);
or U6607 (N_6607,N_3219,N_4005);
xnor U6608 (N_6608,N_5590,N_4625);
nor U6609 (N_6609,N_4497,N_6038);
and U6610 (N_6610,N_4638,N_4673);
and U6611 (N_6611,N_3265,N_5721);
nor U6612 (N_6612,N_5263,N_4909);
nor U6613 (N_6613,N_5411,N_3930);
nand U6614 (N_6614,N_4611,N_6108);
nand U6615 (N_6615,N_4769,N_4159);
or U6616 (N_6616,N_3665,N_4698);
nor U6617 (N_6617,N_4013,N_4049);
nor U6618 (N_6618,N_6103,N_5768);
or U6619 (N_6619,N_4308,N_4952);
or U6620 (N_6620,N_4139,N_3126);
and U6621 (N_6621,N_4905,N_4757);
or U6622 (N_6622,N_3147,N_4056);
nor U6623 (N_6623,N_4230,N_5350);
or U6624 (N_6624,N_4964,N_5964);
and U6625 (N_6625,N_3611,N_4405);
nand U6626 (N_6626,N_3243,N_5493);
nor U6627 (N_6627,N_4630,N_5939);
nand U6628 (N_6628,N_4830,N_5403);
nor U6629 (N_6629,N_5140,N_5113);
nand U6630 (N_6630,N_4198,N_4634);
nand U6631 (N_6631,N_3923,N_5898);
xnor U6632 (N_6632,N_4859,N_4334);
or U6633 (N_6633,N_5538,N_4942);
nand U6634 (N_6634,N_4502,N_5972);
nor U6635 (N_6635,N_3161,N_5921);
or U6636 (N_6636,N_3600,N_4646);
nand U6637 (N_6637,N_4145,N_3984);
nand U6638 (N_6638,N_5974,N_4310);
and U6639 (N_6639,N_5697,N_3866);
nand U6640 (N_6640,N_3246,N_5789);
or U6641 (N_6641,N_4100,N_3620);
and U6642 (N_6642,N_3242,N_4926);
nor U6643 (N_6643,N_6150,N_3818);
nor U6644 (N_6644,N_5394,N_5209);
nand U6645 (N_6645,N_3236,N_5626);
and U6646 (N_6646,N_5450,N_3304);
nor U6647 (N_6647,N_5808,N_3945);
nor U6648 (N_6648,N_5970,N_3296);
xor U6649 (N_6649,N_6045,N_3454);
nor U6650 (N_6650,N_3477,N_4172);
or U6651 (N_6651,N_4275,N_6181);
nand U6652 (N_6652,N_4267,N_3643);
nor U6653 (N_6653,N_3785,N_6000);
xor U6654 (N_6654,N_3158,N_5650);
or U6655 (N_6655,N_5623,N_4731);
nor U6656 (N_6656,N_5087,N_4913);
and U6657 (N_6657,N_3153,N_5642);
nand U6658 (N_6658,N_5047,N_3460);
or U6659 (N_6659,N_6032,N_3675);
xor U6660 (N_6660,N_5466,N_3389);
nor U6661 (N_6661,N_4741,N_4456);
nor U6662 (N_6662,N_4245,N_3556);
nor U6663 (N_6663,N_5670,N_3715);
or U6664 (N_6664,N_4090,N_5040);
xnor U6665 (N_6665,N_5307,N_5449);
nand U6666 (N_6666,N_4477,N_4527);
nand U6667 (N_6667,N_3406,N_6218);
and U6668 (N_6668,N_4531,N_3448);
nor U6669 (N_6669,N_3163,N_4550);
and U6670 (N_6670,N_3944,N_4675);
nand U6671 (N_6671,N_4037,N_3330);
nor U6672 (N_6672,N_4448,N_4369);
xor U6673 (N_6673,N_3826,N_5676);
nor U6674 (N_6674,N_5126,N_4028);
nand U6675 (N_6675,N_4744,N_3610);
and U6676 (N_6676,N_5532,N_5343);
and U6677 (N_6677,N_3478,N_5732);
and U6678 (N_6678,N_6077,N_5716);
xnor U6679 (N_6679,N_4032,N_5894);
nand U6680 (N_6680,N_4104,N_4030);
nor U6681 (N_6681,N_3601,N_4558);
nand U6682 (N_6682,N_5269,N_4350);
nand U6683 (N_6683,N_5303,N_3405);
xnor U6684 (N_6684,N_3401,N_3384);
nor U6685 (N_6685,N_4762,N_4725);
or U6686 (N_6686,N_5206,N_4877);
or U6687 (N_6687,N_5426,N_4787);
or U6688 (N_6688,N_3428,N_5111);
and U6689 (N_6689,N_3209,N_5724);
nand U6690 (N_6690,N_6226,N_3266);
xor U6691 (N_6691,N_3741,N_3306);
nor U6692 (N_6692,N_3734,N_4244);
and U6693 (N_6693,N_5064,N_5270);
nand U6694 (N_6694,N_4076,N_4994);
nor U6695 (N_6695,N_3379,N_5086);
nand U6696 (N_6696,N_3689,N_4478);
nor U6697 (N_6697,N_5211,N_3682);
or U6698 (N_6698,N_4665,N_3814);
nor U6699 (N_6699,N_3583,N_5520);
nand U6700 (N_6700,N_5275,N_3425);
nor U6701 (N_6701,N_5933,N_6129);
xor U6702 (N_6702,N_5161,N_5357);
nor U6703 (N_6703,N_4344,N_4609);
and U6704 (N_6704,N_5678,N_3419);
and U6705 (N_6705,N_3426,N_4413);
or U6706 (N_6706,N_4817,N_4900);
nor U6707 (N_6707,N_5483,N_6207);
nor U6708 (N_6708,N_4525,N_5643);
or U6709 (N_6709,N_5823,N_4191);
nand U6710 (N_6710,N_4722,N_5682);
xnor U6711 (N_6711,N_3702,N_4204);
nor U6712 (N_6712,N_5283,N_6062);
nand U6713 (N_6713,N_3420,N_3188);
nor U6714 (N_6714,N_4081,N_4956);
nand U6715 (N_6715,N_5156,N_3561);
nand U6716 (N_6716,N_5164,N_6019);
nand U6717 (N_6717,N_4708,N_5254);
or U6718 (N_6718,N_3179,N_3596);
and U6719 (N_6719,N_5349,N_3732);
or U6720 (N_6720,N_4027,N_3897);
and U6721 (N_6721,N_5429,N_5598);
or U6722 (N_6722,N_5955,N_3996);
or U6723 (N_6723,N_3320,N_4819);
xor U6724 (N_6724,N_4943,N_4098);
nor U6725 (N_6725,N_3408,N_4765);
or U6726 (N_6726,N_3144,N_3821);
nand U6727 (N_6727,N_4577,N_5486);
nor U6728 (N_6728,N_5942,N_3807);
or U6729 (N_6729,N_4580,N_3797);
and U6730 (N_6730,N_4057,N_6074);
nand U6731 (N_6731,N_4381,N_3134);
nor U6732 (N_6732,N_6243,N_3877);
xor U6733 (N_6733,N_5367,N_3453);
and U6734 (N_6734,N_4846,N_4962);
and U6735 (N_6735,N_5399,N_3479);
or U6736 (N_6736,N_4506,N_5105);
and U6737 (N_6737,N_4624,N_6105);
or U6738 (N_6738,N_3346,N_5242);
nor U6739 (N_6739,N_3882,N_5463);
and U6740 (N_6740,N_5175,N_4896);
or U6741 (N_6741,N_3975,N_5374);
nor U6742 (N_6742,N_5306,N_5454);
xor U6743 (N_6743,N_5860,N_5699);
or U6744 (N_6744,N_4496,N_5244);
nor U6745 (N_6745,N_4532,N_5821);
or U6746 (N_6746,N_5608,N_5226);
xnor U6747 (N_6747,N_5517,N_3578);
nor U6748 (N_6748,N_4633,N_5779);
xor U6749 (N_6749,N_4205,N_6180);
nand U6750 (N_6750,N_5178,N_4663);
or U6751 (N_6751,N_4294,N_3173);
nor U6752 (N_6752,N_4521,N_5625);
and U6753 (N_6753,N_5177,N_5024);
and U6754 (N_6754,N_3299,N_3904);
and U6755 (N_6755,N_3888,N_3377);
xor U6756 (N_6756,N_5322,N_5205);
nand U6757 (N_6757,N_3705,N_5188);
or U6758 (N_6758,N_5218,N_3842);
or U6759 (N_6759,N_4802,N_4544);
and U6760 (N_6760,N_6128,N_3770);
or U6761 (N_6761,N_5118,N_5669);
or U6762 (N_6762,N_6131,N_5712);
or U6763 (N_6763,N_3445,N_6015);
nor U6764 (N_6764,N_3652,N_3613);
xor U6765 (N_6765,N_5021,N_3129);
and U6766 (N_6766,N_3961,N_3555);
or U6767 (N_6767,N_6086,N_4559);
and U6768 (N_6768,N_5379,N_4246);
nand U6769 (N_6769,N_6233,N_3511);
xnor U6770 (N_6770,N_3844,N_4415);
or U6771 (N_6771,N_5708,N_3527);
or U6772 (N_6772,N_5534,N_5761);
and U6773 (N_6773,N_4023,N_4881);
and U6774 (N_6774,N_4127,N_5839);
and U6775 (N_6775,N_6106,N_5675);
and U6776 (N_6776,N_5018,N_3982);
nor U6777 (N_6777,N_3370,N_5376);
and U6778 (N_6778,N_3990,N_4174);
or U6779 (N_6779,N_6154,N_4766);
and U6780 (N_6780,N_4273,N_3972);
and U6781 (N_6781,N_4396,N_5070);
or U6782 (N_6782,N_6140,N_3980);
and U6783 (N_6783,N_5372,N_4228);
or U6784 (N_6784,N_3149,N_5638);
and U6785 (N_6785,N_3598,N_5581);
or U6786 (N_6786,N_5567,N_3271);
nor U6787 (N_6787,N_4287,N_4789);
nand U6788 (N_6788,N_4243,N_5231);
or U6789 (N_6789,N_5044,N_6221);
and U6790 (N_6790,N_4866,N_5308);
or U6791 (N_6791,N_5323,N_4791);
nand U6792 (N_6792,N_6048,N_3730);
nand U6793 (N_6793,N_4073,N_5920);
or U6794 (N_6794,N_4974,N_4466);
nand U6795 (N_6795,N_3751,N_6122);
nand U6796 (N_6796,N_4109,N_3582);
nor U6797 (N_6797,N_3431,N_5232);
nand U6798 (N_6798,N_3323,N_3333);
or U6799 (N_6799,N_6182,N_5045);
nor U6800 (N_6800,N_4935,N_5146);
nand U6801 (N_6801,N_5525,N_3334);
nor U6802 (N_6802,N_5874,N_3154);
nor U6803 (N_6803,N_4838,N_3563);
or U6804 (N_6804,N_4656,N_3180);
nand U6805 (N_6805,N_5497,N_4821);
and U6806 (N_6806,N_3885,N_5022);
nor U6807 (N_6807,N_4538,N_5533);
or U6808 (N_6808,N_5034,N_6246);
nand U6809 (N_6809,N_6219,N_4221);
nor U6810 (N_6810,N_4454,N_5548);
or U6811 (N_6811,N_4200,N_3253);
nand U6812 (N_6812,N_4260,N_5129);
and U6813 (N_6813,N_6026,N_5165);
and U6814 (N_6814,N_3833,N_5356);
nand U6815 (N_6815,N_4508,N_5947);
or U6816 (N_6816,N_4726,N_4707);
nor U6817 (N_6817,N_6017,N_6174);
nor U6818 (N_6818,N_3817,N_4869);
or U6819 (N_6819,N_3659,N_3189);
nor U6820 (N_6820,N_5092,N_5116);
or U6821 (N_6821,N_5666,N_6138);
or U6822 (N_6822,N_3252,N_3660);
nand U6823 (N_6823,N_3764,N_4210);
and U6824 (N_6824,N_5679,N_3865);
and U6825 (N_6825,N_5983,N_3164);
or U6826 (N_6826,N_5762,N_4212);
nor U6827 (N_6827,N_3558,N_5695);
nor U6828 (N_6828,N_5008,N_3402);
nand U6829 (N_6829,N_6160,N_5934);
nand U6830 (N_6830,N_3827,N_4959);
and U6831 (N_6831,N_5542,N_5338);
nand U6832 (N_6832,N_3781,N_3560);
or U6833 (N_6833,N_6222,N_4727);
nor U6834 (N_6834,N_3321,N_5221);
and U6835 (N_6835,N_3187,N_4071);
or U6836 (N_6836,N_5807,N_5730);
nor U6837 (N_6837,N_5750,N_4142);
or U6838 (N_6838,N_5080,N_3772);
nor U6839 (N_6839,N_4279,N_3926);
and U6840 (N_6840,N_3233,N_4730);
and U6841 (N_6841,N_3568,N_3695);
nor U6842 (N_6842,N_4263,N_5854);
and U6843 (N_6843,N_5719,N_5616);
nand U6844 (N_6844,N_6184,N_4890);
nor U6845 (N_6845,N_4364,N_5478);
or U6846 (N_6846,N_3172,N_4238);
and U6847 (N_6847,N_3540,N_5591);
or U6848 (N_6848,N_4844,N_6130);
and U6849 (N_6849,N_6241,N_4811);
and U6850 (N_6850,N_4276,N_4101);
nand U6851 (N_6851,N_5348,N_3417);
xnor U6852 (N_6852,N_5440,N_4933);
xor U6853 (N_6853,N_3554,N_3230);
nor U6854 (N_6854,N_3432,N_5711);
nand U6855 (N_6855,N_5358,N_4997);
and U6856 (N_6856,N_4878,N_4192);
xnor U6857 (N_6857,N_4857,N_5174);
xor U6858 (N_6858,N_3142,N_5917);
nand U6859 (N_6859,N_6109,N_3969);
nor U6860 (N_6860,N_4349,N_3709);
nand U6861 (N_6861,N_4719,N_5181);
or U6862 (N_6862,N_4163,N_5258);
xnor U6863 (N_6863,N_3839,N_4099);
and U6864 (N_6864,N_5948,N_4055);
or U6865 (N_6865,N_5740,N_6245);
nand U6866 (N_6866,N_4917,N_6002);
nand U6867 (N_6867,N_3733,N_6080);
nand U6868 (N_6868,N_4667,N_5539);
nand U6869 (N_6869,N_6053,N_4361);
and U6870 (N_6870,N_3132,N_4925);
or U6871 (N_6871,N_4148,N_5039);
nor U6872 (N_6872,N_4586,N_3400);
and U6873 (N_6873,N_3290,N_4388);
nand U6874 (N_6874,N_5745,N_5133);
nand U6875 (N_6875,N_5207,N_5847);
nand U6876 (N_6876,N_5991,N_5900);
nor U6877 (N_6877,N_4211,N_4219);
and U6878 (N_6878,N_3777,N_5359);
nor U6879 (N_6879,N_5470,N_4437);
and U6880 (N_6880,N_5510,N_4044);
nand U6881 (N_6881,N_6110,N_5834);
and U6882 (N_6882,N_3918,N_6175);
nor U6883 (N_6883,N_5545,N_4591);
nand U6884 (N_6884,N_5896,N_5406);
xor U6885 (N_6885,N_3151,N_5115);
or U6886 (N_6886,N_3518,N_4339);
and U6887 (N_6887,N_3268,N_3716);
xor U6888 (N_6888,N_5051,N_5371);
nand U6889 (N_6889,N_4702,N_4835);
nand U6890 (N_6890,N_3475,N_3763);
and U6891 (N_6891,N_4445,N_3489);
nor U6892 (N_6892,N_4291,N_4723);
or U6893 (N_6893,N_5926,N_4654);
and U6894 (N_6894,N_5868,N_4220);
nand U6895 (N_6895,N_4152,N_5720);
nor U6896 (N_6896,N_5009,N_3962);
or U6897 (N_6897,N_3287,N_4059);
and U6898 (N_6898,N_5117,N_3894);
nand U6899 (N_6899,N_3522,N_6051);
or U6900 (N_6900,N_5554,N_3316);
or U6901 (N_6901,N_5130,N_5431);
and U6902 (N_6902,N_4587,N_3739);
nor U6903 (N_6903,N_3491,N_4608);
and U6904 (N_6904,N_4322,N_3344);
and U6905 (N_6905,N_3735,N_6056);
nor U6906 (N_6906,N_5314,N_5415);
nand U6907 (N_6907,N_3876,N_3282);
nor U6908 (N_6908,N_4898,N_3240);
and U6909 (N_6909,N_4207,N_3589);
nor U6910 (N_6910,N_5794,N_3992);
nor U6911 (N_6911,N_3786,N_5773);
or U6912 (N_6912,N_4314,N_4426);
nand U6913 (N_6913,N_4010,N_5337);
nor U6914 (N_6914,N_4286,N_4578);
nor U6915 (N_6915,N_4468,N_5067);
nor U6916 (N_6916,N_5690,N_4252);
or U6917 (N_6917,N_4845,N_6230);
and U6918 (N_6918,N_3811,N_4764);
nor U6919 (N_6919,N_5817,N_4195);
xor U6920 (N_6920,N_3315,N_5046);
xnor U6921 (N_6921,N_4600,N_4927);
nand U6922 (N_6922,N_4885,N_5778);
nor U6923 (N_6923,N_3683,N_3758);
xnor U6924 (N_6924,N_4143,N_5468);
nor U6925 (N_6925,N_5128,N_6216);
and U6926 (N_6926,N_3646,N_5541);
and U6927 (N_6927,N_5918,N_4807);
nand U6928 (N_6928,N_3791,N_3753);
nor U6929 (N_6929,N_3803,N_4138);
and U6930 (N_6930,N_4345,N_5462);
nand U6931 (N_6931,N_5019,N_3446);
or U6932 (N_6932,N_4597,N_6115);
and U6933 (N_6933,N_4366,N_3837);
or U6934 (N_6934,N_5503,N_5298);
nor U6935 (N_6935,N_5776,N_3916);
nor U6936 (N_6936,N_5060,N_5634);
and U6937 (N_6937,N_3182,N_4639);
or U6938 (N_6938,N_5312,N_5378);
nor U6939 (N_6939,N_4697,N_4967);
nand U6940 (N_6940,N_4618,N_5726);
or U6941 (N_6941,N_5010,N_4065);
and U6942 (N_6942,N_3409,N_6090);
nand U6943 (N_6943,N_5282,N_4661);
nand U6944 (N_6944,N_4316,N_5645);
or U6945 (N_6945,N_5966,N_4779);
or U6946 (N_6946,N_5253,N_4588);
or U6947 (N_6947,N_3297,N_5257);
or U6948 (N_6948,N_4451,N_4884);
nor U6949 (N_6949,N_6009,N_4442);
and U6950 (N_6950,N_5249,N_5210);
or U6951 (N_6951,N_3269,N_4021);
and U6952 (N_6952,N_3436,N_3145);
nor U6953 (N_6953,N_5006,N_3225);
or U6954 (N_6954,N_5587,N_4465);
nor U6955 (N_6955,N_4129,N_3870);
and U6956 (N_6956,N_4979,N_5346);
and U6957 (N_6957,N_3933,N_3277);
nor U6958 (N_6958,N_3875,N_4006);
and U6959 (N_6959,N_5419,N_4333);
nand U6960 (N_6960,N_5200,N_4302);
nand U6961 (N_6961,N_4681,N_5928);
or U6962 (N_6962,N_3997,N_3456);
and U6963 (N_6963,N_5261,N_5280);
and U6964 (N_6964,N_4387,N_6228);
nand U6965 (N_6965,N_5951,N_3413);
nor U6966 (N_6966,N_4256,N_5806);
and U6967 (N_6967,N_4912,N_5409);
nand U6968 (N_6968,N_3539,N_4566);
nand U6969 (N_6969,N_4102,N_3538);
nand U6970 (N_6970,N_5197,N_3559);
and U6971 (N_6971,N_3548,N_5340);
xnor U6972 (N_6972,N_3337,N_3943);
nor U6973 (N_6973,N_4458,N_4923);
nor U6974 (N_6974,N_6081,N_6020);
or U6975 (N_6975,N_3639,N_5093);
and U6976 (N_6976,N_3746,N_4747);
or U6977 (N_6977,N_3884,N_4217);
nor U6978 (N_6978,N_3410,N_5689);
nor U6979 (N_6979,N_5134,N_3993);
or U6980 (N_6980,N_4343,N_4463);
or U6981 (N_6981,N_4144,N_5015);
nand U6982 (N_6982,N_3973,N_5573);
nor U6983 (N_6983,N_4918,N_3465);
xnor U6984 (N_6984,N_5137,N_5757);
nand U6985 (N_6985,N_4582,N_5001);
xor U6986 (N_6986,N_3343,N_4319);
nand U6987 (N_6987,N_4907,N_4450);
nand U6988 (N_6988,N_4272,N_4372);
nor U6989 (N_6989,N_6220,N_3549);
or U6990 (N_6990,N_4283,N_4208);
and U6991 (N_6991,N_5743,N_6208);
xor U6992 (N_6992,N_5826,N_5783);
xnor U6993 (N_6993,N_6156,N_4938);
and U6994 (N_6994,N_5744,N_3840);
nor U6995 (N_6995,N_3234,N_5159);
and U6996 (N_6996,N_3931,N_5481);
nor U6997 (N_6997,N_4676,N_3232);
xor U6998 (N_6998,N_5600,N_6099);
xnor U6999 (N_6999,N_5259,N_3815);
and U7000 (N_7000,N_3254,N_3198);
or U7001 (N_7001,N_3932,N_3919);
and U7002 (N_7002,N_4908,N_4321);
nor U7003 (N_7003,N_5241,N_6139);
and U7004 (N_7004,N_4051,N_5393);
or U7005 (N_7005,N_3466,N_6162);
nand U7006 (N_7006,N_6082,N_3393);
or U7007 (N_7007,N_6183,N_5075);
or U7008 (N_7008,N_4814,N_3248);
or U7009 (N_7009,N_3686,N_4572);
xnor U7010 (N_7010,N_4399,N_3536);
nor U7011 (N_7011,N_5496,N_5652);
nor U7012 (N_7012,N_6027,N_5811);
xnor U7013 (N_7013,N_3291,N_5798);
nor U7014 (N_7014,N_5230,N_3908);
and U7015 (N_7015,N_5309,N_4268);
nand U7016 (N_7016,N_3902,N_6239);
nand U7017 (N_7017,N_5506,N_3862);
and U7018 (N_7018,N_3832,N_5574);
nor U7019 (N_7019,N_4628,N_5701);
nor U7020 (N_7020,N_4356,N_5565);
nand U7021 (N_7021,N_5131,N_4562);
xnor U7022 (N_7022,N_3338,N_4820);
nand U7023 (N_7023,N_3327,N_6091);
nand U7024 (N_7024,N_5330,N_4461);
nand U7025 (N_7025,N_5915,N_6037);
or U7026 (N_7026,N_3354,N_3985);
xnor U7027 (N_7027,N_3874,N_4464);
or U7028 (N_7028,N_4367,N_3283);
xnor U7029 (N_7029,N_5793,N_4735);
xor U7030 (N_7030,N_4593,N_3618);
and U7031 (N_7031,N_4643,N_4603);
and U7032 (N_7032,N_3661,N_4713);
xnor U7033 (N_7033,N_4409,N_3220);
and U7034 (N_7034,N_6059,N_6177);
xor U7035 (N_7035,N_3765,N_3178);
nor U7036 (N_7036,N_3169,N_6028);
and U7037 (N_7037,N_5476,N_4983);
and U7038 (N_7038,N_4054,N_4003);
or U7039 (N_7039,N_3339,N_5032);
and U7040 (N_7040,N_5511,N_4986);
xnor U7041 (N_7041,N_4916,N_5321);
xor U7042 (N_7042,N_3780,N_5420);
nand U7043 (N_7043,N_5480,N_5148);
nor U7044 (N_7044,N_4605,N_5090);
xor U7045 (N_7045,N_3697,N_4313);
and U7046 (N_7046,N_4501,N_6104);
nand U7047 (N_7047,N_4685,N_6224);
nand U7048 (N_7048,N_3606,N_6166);
nand U7049 (N_7049,N_4335,N_5229);
and U7050 (N_7050,N_3788,N_4325);
nor U7051 (N_7051,N_3789,N_5305);
and U7052 (N_7052,N_3534,N_3440);
nand U7053 (N_7053,N_5360,N_6012);
and U7054 (N_7054,N_4622,N_5224);
and U7055 (N_7055,N_3964,N_5315);
or U7056 (N_7056,N_4395,N_5846);
or U7057 (N_7057,N_3288,N_5995);
or U7058 (N_7058,N_5957,N_3880);
and U7059 (N_7059,N_5786,N_5016);
nand U7060 (N_7060,N_5180,N_4247);
nand U7061 (N_7061,N_4323,N_4872);
or U7062 (N_7062,N_4020,N_4563);
nor U7063 (N_7063,N_3856,N_5936);
or U7064 (N_7064,N_4154,N_4889);
or U7065 (N_7065,N_5954,N_5333);
or U7066 (N_7066,N_4116,N_5805);
and U7067 (N_7067,N_3719,N_5203);
nand U7068 (N_7068,N_6186,N_5869);
xor U7069 (N_7069,N_4827,N_4473);
xnor U7070 (N_7070,N_6041,N_5672);
or U7071 (N_7071,N_4340,N_6079);
nand U7072 (N_7072,N_6170,N_5425);
nor U7073 (N_7073,N_4670,N_5551);
or U7074 (N_7074,N_3303,N_5589);
nor U7075 (N_7075,N_5560,N_6034);
nand U7076 (N_7076,N_3201,N_5442);
nor U7077 (N_7077,N_4022,N_3636);
nor U7078 (N_7078,N_3574,N_5632);
and U7079 (N_7079,N_3434,N_3524);
xnor U7080 (N_7080,N_5494,N_4842);
nor U7081 (N_7081,N_4389,N_5759);
and U7082 (N_7082,N_3383,N_4309);
nand U7083 (N_7083,N_3612,N_4862);
xor U7084 (N_7084,N_4785,N_5850);
nand U7085 (N_7085,N_3591,N_3581);
or U7086 (N_7086,N_4557,N_5310);
and U7087 (N_7087,N_5585,N_3965);
nand U7088 (N_7088,N_5456,N_5266);
nor U7089 (N_7089,N_6249,N_4227);
nand U7090 (N_7090,N_4421,N_4402);
or U7091 (N_7091,N_3285,N_3552);
or U7092 (N_7092,N_5013,N_5501);
and U7093 (N_7093,N_4718,N_3917);
nor U7094 (N_7094,N_3519,N_5731);
xnor U7095 (N_7095,N_4112,N_5074);
nor U7096 (N_7096,N_5553,N_5445);
nand U7097 (N_7097,N_3437,N_5631);
and U7098 (N_7098,N_3590,N_5859);
and U7099 (N_7099,N_3311,N_4107);
xor U7100 (N_7100,N_6067,N_5272);
nand U7101 (N_7101,N_4018,N_5944);
or U7102 (N_7102,N_4576,N_5048);
nand U7103 (N_7103,N_3521,N_3914);
or U7104 (N_7104,N_3160,N_4695);
and U7105 (N_7105,N_5110,N_6240);
xor U7106 (N_7106,N_5313,N_3621);
and U7107 (N_7107,N_5005,N_5460);
nor U7108 (N_7108,N_4160,N_4931);
and U7109 (N_7109,N_6121,N_3615);
nand U7110 (N_7110,N_4688,N_4855);
and U7111 (N_7111,N_6021,N_6164);
or U7112 (N_7112,N_4504,N_4812);
nor U7113 (N_7113,N_6165,N_5423);
and U7114 (N_7114,N_3708,N_5698);
nor U7115 (N_7115,N_5902,N_3165);
nor U7116 (N_7116,N_3520,N_5292);
nor U7117 (N_7117,N_5089,N_4520);
nor U7118 (N_7118,N_5563,N_5147);
and U7119 (N_7119,N_5862,N_4831);
nor U7120 (N_7120,N_5612,N_4883);
and U7121 (N_7121,N_3841,N_5527);
nand U7122 (N_7122,N_4250,N_4216);
nor U7123 (N_7123,N_6205,N_4242);
or U7124 (N_7124,N_4180,N_5085);
nand U7125 (N_7125,N_4318,N_5302);
and U7126 (N_7126,N_4946,N_5848);
nand U7127 (N_7127,N_3737,N_4662);
or U7128 (N_7128,N_4011,N_4937);
nor U7129 (N_7129,N_5756,N_4386);
nor U7130 (N_7130,N_5279,N_4380);
and U7131 (N_7131,N_4848,N_4374);
nand U7132 (N_7132,N_4960,N_4875);
xor U7133 (N_7133,N_4342,N_3125);
nand U7134 (N_7134,N_5383,N_4176);
or U7135 (N_7135,N_3638,N_4336);
or U7136 (N_7136,N_5787,N_3543);
or U7137 (N_7137,N_4016,N_5559);
nor U7138 (N_7138,N_6050,N_4223);
nand U7139 (N_7139,N_4080,N_4828);
and U7140 (N_7140,N_4271,N_5236);
nor U7141 (N_7141,N_5903,N_4337);
xnor U7142 (N_7142,N_5965,N_4784);
nand U7143 (N_7143,N_6194,N_3439);
and U7144 (N_7144,N_5605,N_4128);
nand U7145 (N_7145,N_3386,N_3805);
or U7146 (N_7146,N_5580,N_5518);
nand U7147 (N_7147,N_4516,N_4513);
nand U7148 (N_7148,N_4971,N_5922);
or U7149 (N_7149,N_3644,N_5030);
or U7150 (N_7150,N_5646,N_3474);
nand U7151 (N_7151,N_4774,N_4996);
and U7152 (N_7152,N_4126,N_4499);
or U7153 (N_7153,N_5892,N_3669);
and U7154 (N_7154,N_5931,N_6023);
and U7155 (N_7155,N_5370,N_4134);
and U7156 (N_7156,N_3810,N_3378);
nor U7157 (N_7157,N_3459,N_4854);
and U7158 (N_7158,N_4748,N_5684);
and U7159 (N_7159,N_4236,N_4365);
nand U7160 (N_7160,N_5871,N_4452);
nand U7161 (N_7161,N_4285,N_5000);
and U7162 (N_7162,N_3139,N_3820);
nor U7163 (N_7163,N_5291,N_4184);
nand U7164 (N_7164,N_6169,N_5741);
or U7165 (N_7165,N_4690,N_5331);
xor U7166 (N_7166,N_4901,N_4441);
xor U7167 (N_7167,N_3915,N_5677);
nand U7168 (N_7168,N_3496,N_3128);
xor U7169 (N_7169,N_4745,N_3963);
nor U7170 (N_7170,N_4581,N_5556);
or U7171 (N_7171,N_5685,N_4867);
or U7172 (N_7172,N_4621,N_5162);
or U7173 (N_7173,N_3934,N_3629);
nor U7174 (N_7174,N_3663,N_4928);
nor U7175 (N_7175,N_5099,N_4072);
nand U7176 (N_7176,N_4783,N_5136);
and U7177 (N_7177,N_5286,N_4957);
xnor U7178 (N_7178,N_3863,N_5572);
and U7179 (N_7179,N_3640,N_4255);
xor U7180 (N_7180,N_6111,N_3712);
nor U7181 (N_7181,N_4575,N_4460);
nand U7182 (N_7182,N_4103,N_4607);
or U7183 (N_7183,N_5938,N_5132);
or U7184 (N_7184,N_5977,N_3135);
or U7185 (N_7185,N_3515,N_4778);
or U7186 (N_7186,N_5994,N_5341);
or U7187 (N_7187,N_6142,N_5499);
and U7188 (N_7188,N_5397,N_5327);
and U7189 (N_7189,N_4249,N_4026);
and U7190 (N_7190,N_3319,N_4632);
and U7191 (N_7191,N_4861,N_4796);
or U7192 (N_7192,N_5464,N_4839);
nand U7193 (N_7193,N_3883,N_3869);
xnor U7194 (N_7194,N_5733,N_6161);
and U7195 (N_7195,N_3570,N_4650);
nor U7196 (N_7196,N_5519,N_3407);
nor U7197 (N_7197,N_3727,N_3544);
nand U7198 (N_7198,N_3427,N_4407);
nor U7199 (N_7199,N_4598,N_5407);
nand U7200 (N_7200,N_3767,N_4082);
or U7201 (N_7201,N_4843,N_6172);
nand U7202 (N_7202,N_5725,N_4978);
nand U7203 (N_7203,N_3238,N_3174);
or U7204 (N_7204,N_3262,N_5444);
nor U7205 (N_7205,N_4834,N_3208);
nand U7206 (N_7206,N_4232,N_5155);
and U7207 (N_7207,N_3657,N_5058);
nand U7208 (N_7208,N_5713,N_4459);
nor U7209 (N_7209,N_4173,N_5057);
and U7210 (N_7210,N_5714,N_5929);
nor U7211 (N_7211,N_4620,N_5971);
or U7212 (N_7212,N_6016,N_4953);
and U7213 (N_7213,N_5071,N_5017);
xnor U7214 (N_7214,N_4715,N_3483);
nand U7215 (N_7215,N_5584,N_5760);
nor U7216 (N_7216,N_3517,N_5184);
and U7217 (N_7217,N_4910,N_4987);
nand U7218 (N_7218,N_3891,N_4234);
nand U7219 (N_7219,N_4231,N_5289);
and U7220 (N_7220,N_6193,N_4589);
nor U7221 (N_7221,N_5620,N_3694);
nand U7222 (N_7222,N_4767,N_5260);
or U7223 (N_7223,N_4482,N_4805);
nor U7224 (N_7224,N_3196,N_5381);
and U7225 (N_7225,N_3357,N_3920);
nor U7226 (N_7226,N_3599,N_5557);
nand U7227 (N_7227,N_3237,N_6061);
and U7228 (N_7228,N_4801,N_5802);
nor U7229 (N_7229,N_3387,N_5907);
and U7230 (N_7230,N_4958,N_6058);
or U7231 (N_7231,N_4761,N_5077);
or U7232 (N_7232,N_5990,N_3418);
nand U7233 (N_7233,N_3476,N_3793);
nor U7234 (N_7234,N_4346,N_4541);
and U7235 (N_7235,N_5029,N_4768);
nor U7236 (N_7236,N_3701,N_4594);
or U7237 (N_7237,N_4067,N_3761);
nand U7238 (N_7238,N_5098,N_4529);
nor U7239 (N_7239,N_3542,N_4961);
nand U7240 (N_7240,N_6188,N_5273);
nor U7241 (N_7241,N_5094,N_5641);
and U7242 (N_7242,N_5653,N_3922);
nand U7243 (N_7243,N_5182,N_3795);
and U7244 (N_7244,N_5168,N_5251);
nor U7245 (N_7245,N_4536,N_5380);
nor U7246 (N_7246,N_3977,N_5686);
nor U7247 (N_7247,N_3911,N_4411);
nand U7248 (N_7248,N_3672,N_5630);
or U7249 (N_7249,N_4419,N_4296);
and U7250 (N_7250,N_5204,N_5828);
or U7251 (N_7251,N_5274,N_3295);
nand U7252 (N_7252,N_3633,N_4546);
nor U7253 (N_7253,N_6013,N_5300);
and U7254 (N_7254,N_3743,N_5139);
nor U7255 (N_7255,N_4137,N_3995);
and U7256 (N_7256,N_3595,N_5326);
and U7257 (N_7257,N_5490,N_4679);
and U7258 (N_7258,N_3819,N_4254);
and U7259 (N_7259,N_3688,N_6126);
and U7260 (N_7260,N_3806,N_5056);
or U7261 (N_7261,N_5796,N_3155);
nor U7262 (N_7262,N_3244,N_4752);
or U7263 (N_7263,N_4031,N_4737);
nor U7264 (N_7264,N_5615,N_5199);
nand U7265 (N_7265,N_4008,N_4431);
and U7266 (N_7266,N_5710,N_3852);
and U7267 (N_7267,N_4824,N_5491);
xnor U7268 (N_7268,N_3860,N_4808);
or U7269 (N_7269,N_4009,N_5109);
or U7270 (N_7270,N_4717,N_3571);
nor U7271 (N_7271,N_4430,N_3575);
and U7272 (N_7272,N_3308,N_4976);
nand U7273 (N_7273,N_5096,N_3205);
xnor U7274 (N_7274,N_4792,N_4084);
or U7275 (N_7275,N_4592,N_3493);
nand U7276 (N_7276,N_3140,N_4829);
nand U7277 (N_7277,N_4060,N_6052);
nand U7278 (N_7278,N_4382,N_3325);
nand U7279 (N_7279,N_4899,N_3667);
nand U7280 (N_7280,N_4729,N_5683);
and U7281 (N_7281,N_3740,N_3779);
nand U7282 (N_7282,N_4375,N_6088);
nand U7283 (N_7283,N_5377,N_4487);
nor U7284 (N_7284,N_3231,N_5910);
nor U7285 (N_7285,N_4579,N_6044);
nand U7286 (N_7286,N_4069,N_3239);
or U7287 (N_7287,N_4780,N_3662);
nand U7288 (N_7288,N_4390,N_5961);
nor U7289 (N_7289,N_3349,N_3394);
or U7290 (N_7290,N_5578,N_3890);
and U7291 (N_7291,N_5294,N_3141);
or U7292 (N_7292,N_5194,N_4171);
and U7293 (N_7293,N_3485,N_5586);
or U7294 (N_7294,N_5664,N_5962);
nand U7295 (N_7295,N_4196,N_4427);
and U7296 (N_7296,N_4226,N_4657);
nand U7297 (N_7297,N_3898,N_3861);
nand U7298 (N_7298,N_3309,N_4535);
and U7299 (N_7299,N_4640,N_3846);
nor U7300 (N_7300,N_5458,N_5055);
nor U7301 (N_7301,N_3441,N_5627);
and U7302 (N_7302,N_5694,N_6083);
or U7303 (N_7303,N_5765,N_4560);
or U7304 (N_7304,N_5867,N_4106);
nand U7305 (N_7305,N_3498,N_4063);
and U7306 (N_7306,N_3312,N_5042);
and U7307 (N_7307,N_4919,N_4293);
or U7308 (N_7308,N_5212,N_4932);
nor U7309 (N_7309,N_6092,N_3531);
nor U7310 (N_7310,N_4315,N_3284);
nand U7311 (N_7311,N_5662,N_4626);
nand U7312 (N_7312,N_3831,N_5809);
and U7313 (N_7313,N_5784,N_3704);
or U7314 (N_7314,N_5271,N_4251);
nor U7315 (N_7315,N_5651,N_3184);
nor U7316 (N_7316,N_4179,N_5438);
or U7317 (N_7317,N_3830,N_5457);
or U7318 (N_7318,N_5288,N_6071);
and U7319 (N_7319,N_3430,N_3867);
nand U7320 (N_7320,N_3736,N_3801);
or U7321 (N_7321,N_4096,N_6007);
nand U7322 (N_7322,N_4141,N_5801);
nand U7323 (N_7323,N_5225,N_5629);
and U7324 (N_7324,N_5858,N_3787);
or U7325 (N_7325,N_4187,N_5606);
or U7326 (N_7326,N_3241,N_4941);
nor U7327 (N_7327,N_5734,N_5909);
or U7328 (N_7328,N_4338,N_5437);
nor U7329 (N_7329,N_6031,N_3614);
nand U7330 (N_7330,N_4029,N_4017);
nand U7331 (N_7331,N_3335,N_3854);
and U7332 (N_7332,N_5540,N_5876);
nor U7333 (N_7333,N_3668,N_6076);
nor U7334 (N_7334,N_3528,N_3452);
xnor U7335 (N_7335,N_6065,N_5396);
nand U7336 (N_7336,N_3257,N_5999);
nand U7337 (N_7337,N_4470,N_3300);
or U7338 (N_7338,N_5103,N_5003);
or U7339 (N_7339,N_4358,N_3960);
nand U7340 (N_7340,N_5561,N_6054);
or U7341 (N_7341,N_4847,N_3809);
nor U7342 (N_7342,N_4157,N_4542);
and U7343 (N_7343,N_4495,N_4617);
xnor U7344 (N_7344,N_6025,N_5884);
xor U7345 (N_7345,N_4161,N_4833);
and U7346 (N_7346,N_3372,N_6036);
and U7347 (N_7347,N_4423,N_3684);
and U7348 (N_7348,N_3162,N_6004);
nor U7349 (N_7349,N_5771,N_4097);
nor U7350 (N_7350,N_4209,N_4151);
or U7351 (N_7351,N_4121,N_5335);
nor U7352 (N_7352,N_3587,N_5700);
nand U7353 (N_7353,N_3724,N_4476);
xor U7354 (N_7354,N_4403,N_4614);
nor U7355 (N_7355,N_5639,N_5893);
nor U7356 (N_7356,N_3171,N_5102);
or U7357 (N_7357,N_4201,N_4972);
or U7358 (N_7358,N_5214,N_5888);
nand U7359 (N_7359,N_4108,N_3604);
or U7360 (N_7360,N_3473,N_5536);
nand U7361 (N_7361,N_3783,N_4202);
and U7362 (N_7362,N_6117,N_4401);
and U7363 (N_7363,N_4324,N_5755);
nand U7364 (N_7364,N_5611,N_5256);
nand U7365 (N_7365,N_6159,N_3398);
xnor U7366 (N_7366,N_5404,N_3991);
nor U7367 (N_7367,N_3899,N_3966);
xor U7368 (N_7368,N_5989,N_4329);
nor U7369 (N_7369,N_4773,N_3203);
and U7370 (N_7370,N_5465,N_5012);
nor U7371 (N_7371,N_3365,N_6152);
nand U7372 (N_7372,N_5738,N_3138);
or U7373 (N_7373,N_3666,N_3585);
nand U7374 (N_7374,N_6127,N_4053);
nand U7375 (N_7375,N_4131,N_4120);
or U7376 (N_7376,N_3989,N_3341);
nand U7377 (N_7377,N_3872,N_4756);
nand U7378 (N_7378,N_3514,N_5453);
nor U7379 (N_7379,N_5703,N_3314);
nor U7380 (N_7380,N_3717,N_4320);
nor U7381 (N_7381,N_4024,N_5681);
nand U7382 (N_7382,N_5166,N_4370);
or U7383 (N_7383,N_3691,N_4658);
xnor U7384 (N_7384,N_6237,N_5566);
nand U7385 (N_7385,N_3562,N_6046);
nand U7386 (N_7386,N_3375,N_5339);
or U7387 (N_7387,N_5487,N_5234);
nor U7388 (N_7388,N_5160,N_3580);
and U7389 (N_7389,N_4876,N_3851);
nor U7390 (N_7390,N_4781,N_4945);
and U7391 (N_7391,N_5772,N_5502);
nand U7392 (N_7392,N_6069,N_5385);
nor U7393 (N_7393,N_5223,N_5430);
or U7394 (N_7394,N_4584,N_6040);
xnor U7395 (N_7395,N_3324,N_4408);
nand U7396 (N_7396,N_5319,N_3774);
or U7397 (N_7397,N_3771,N_5555);
nand U7398 (N_7398,N_4904,N_3651);
or U7399 (N_7399,N_5824,N_5981);
nand U7400 (N_7400,N_3673,N_4816);
nor U7401 (N_7401,N_4305,N_5163);
nand U7402 (N_7402,N_5069,N_5498);
and U7403 (N_7403,N_3699,N_4509);
nor U7404 (N_7404,N_5636,N_6236);
or U7405 (N_7405,N_4687,N_5081);
or U7406 (N_7406,N_4936,N_5187);
xnor U7407 (N_7407,N_4164,N_5062);
nand U7408 (N_7408,N_5841,N_3210);
nor U7409 (N_7409,N_6210,N_3449);
or U7410 (N_7410,N_5950,N_4443);
nand U7411 (N_7411,N_3565,N_4136);
xor U7412 (N_7412,N_4606,N_4543);
or U7413 (N_7413,N_5317,N_3825);
or U7414 (N_7414,N_4772,N_5800);
nor U7415 (N_7415,N_4782,N_4259);
and U7416 (N_7416,N_6075,N_5663);
or U7417 (N_7417,N_6024,N_5386);
or U7418 (N_7418,N_6118,N_3762);
and U7419 (N_7419,N_3167,N_4311);
nand U7420 (N_7420,N_5988,N_4720);
and U7421 (N_7421,N_4089,N_3168);
and U7422 (N_7422,N_4728,N_5523);
nand U7423 (N_7423,N_4524,N_5123);
and U7424 (N_7424,N_6189,N_3616);
xnor U7425 (N_7425,N_4297,N_3359);
nand U7426 (N_7426,N_4354,N_5746);
nand U7427 (N_7427,N_5945,N_3221);
nor U7428 (N_7428,N_5172,N_5923);
or U7429 (N_7429,N_3512,N_5171);
nor U7430 (N_7430,N_4793,N_4475);
nand U7431 (N_7431,N_5758,N_3245);
xor U7432 (N_7432,N_3416,N_5904);
and U7433 (N_7433,N_5149,N_4035);
nand U7434 (N_7434,N_4732,N_4241);
and U7435 (N_7435,N_3356,N_5373);
xor U7436 (N_7436,N_4511,N_6163);
or U7437 (N_7437,N_3195,N_4734);
nand U7438 (N_7438,N_3458,N_5384);
or U7439 (N_7439,N_3553,N_5885);
nor U7440 (N_7440,N_5775,N_5382);
nand U7441 (N_7441,N_5537,N_5135);
nand U7442 (N_7442,N_6145,N_5935);
xnor U7443 (N_7443,N_5582,N_3374);
nor U7444 (N_7444,N_5011,N_5579);
nor U7445 (N_7445,N_6209,N_5691);
nand U7446 (N_7446,N_3486,N_4934);
and U7447 (N_7447,N_5530,N_3131);
nor U7448 (N_7448,N_4677,N_3749);
and U7449 (N_7449,N_3532,N_4379);
nand U7450 (N_7450,N_5843,N_4672);
xor U7451 (N_7451,N_4888,N_5992);
nor U7452 (N_7452,N_4303,N_3222);
and U7453 (N_7453,N_5886,N_3258);
nor U7454 (N_7454,N_3950,N_3752);
or U7455 (N_7455,N_3396,N_5790);
xor U7456 (N_7456,N_4394,N_5004);
nor U7457 (N_7457,N_5268,N_5594);
or U7458 (N_7458,N_4257,N_4758);
nor U7459 (N_7459,N_4025,N_4119);
nand U7460 (N_7460,N_5647,N_3726);
and U7461 (N_7461,N_3550,N_6214);
and U7462 (N_7462,N_3949,N_3347);
nand U7463 (N_7463,N_4507,N_3443);
nor U7464 (N_7464,N_4906,N_3557);
and U7465 (N_7465,N_5979,N_4412);
or U7466 (N_7466,N_4214,N_4331);
nor U7467 (N_7467,N_4483,N_6102);
or U7468 (N_7468,N_3597,N_5072);
or U7469 (N_7469,N_4706,N_5173);
nand U7470 (N_7470,N_3573,N_3148);
xnor U7471 (N_7471,N_4203,N_3584);
or U7472 (N_7472,N_5434,N_3784);
nor U7473 (N_7473,N_3506,N_3759);
and U7474 (N_7474,N_4269,N_4397);
nand U7475 (N_7475,N_3952,N_4278);
nor U7476 (N_7476,N_3192,N_3166);
nand U7477 (N_7477,N_4341,N_4488);
or U7478 (N_7478,N_4738,N_5596);
nand U7479 (N_7479,N_4863,N_4627);
nand U7480 (N_7480,N_3157,N_5671);
and U7481 (N_7481,N_5368,N_6097);
or U7482 (N_7482,N_3855,N_4079);
or U7483 (N_7483,N_5106,N_4786);
nand U7484 (N_7484,N_4500,N_3650);
nor U7485 (N_7485,N_6187,N_4514);
nor U7486 (N_7486,N_3586,N_3305);
nor U7487 (N_7487,N_5285,N_4481);
or U7488 (N_7488,N_5911,N_4864);
or U7489 (N_7489,N_4277,N_5041);
nor U7490 (N_7490,N_4545,N_6114);
nand U7491 (N_7491,N_6116,N_3537);
or U7492 (N_7492,N_5489,N_5332);
and U7493 (N_7493,N_3609,N_5250);
or U7494 (N_7494,N_5369,N_4078);
or U7495 (N_7495,N_4261,N_4561);
nor U7496 (N_7496,N_3447,N_3516);
nand U7497 (N_7497,N_5400,N_3878);
and U7498 (N_7498,N_5459,N_4019);
or U7499 (N_7499,N_5899,N_3541);
nor U7500 (N_7500,N_4895,N_6035);
or U7501 (N_7501,N_5814,N_5516);
nand U7502 (N_7502,N_4292,N_4547);
nand U7503 (N_7503,N_4555,N_5053);
or U7504 (N_7504,N_4970,N_4433);
and U7505 (N_7505,N_4860,N_5049);
or U7506 (N_7506,N_4166,N_4775);
nor U7507 (N_7507,N_5825,N_4306);
xor U7508 (N_7508,N_5851,N_3968);
nand U7509 (N_7509,N_6063,N_5583);
nand U7510 (N_7510,N_4363,N_5901);
or U7511 (N_7511,N_5033,N_4114);
nor U7512 (N_7512,N_5696,N_5296);
or U7513 (N_7513,N_4701,N_3588);
and U7514 (N_7514,N_3464,N_6124);
nor U7515 (N_7515,N_5593,N_5522);
nand U7516 (N_7516,N_6157,N_4479);
xnor U7517 (N_7517,N_4794,N_3687);
nand U7518 (N_7518,N_4822,N_4147);
or U7519 (N_7519,N_6066,N_5795);
or U7520 (N_7520,N_5735,N_5815);
nor U7521 (N_7521,N_6018,N_3191);
nand U7522 (N_7522,N_4894,N_3714);
nor U7523 (N_7523,N_3267,N_6010);
and U7524 (N_7524,N_5120,N_3678);
nand U7525 (N_7525,N_5637,N_3681);
nor U7526 (N_7526,N_5073,N_4798);
nand U7527 (N_7527,N_3513,N_5803);
or U7528 (N_7528,N_4636,N_4674);
or U7529 (N_7529,N_4635,N_4462);
or U7530 (N_7530,N_5277,N_6234);
and U7531 (N_7531,N_3294,N_5838);
and U7532 (N_7532,N_5492,N_3368);
and U7533 (N_7533,N_3593,N_4167);
nor U7534 (N_7534,N_3302,N_3744);
and U7535 (N_7535,N_4897,N_4537);
or U7536 (N_7536,N_4991,N_5262);
nor U7537 (N_7537,N_4280,N_5599);
or U7538 (N_7538,N_5930,N_5252);
xor U7539 (N_7539,N_5993,N_5065);
or U7540 (N_7540,N_3461,N_5427);
and U7541 (N_7541,N_5603,N_6003);
xnor U7542 (N_7542,N_3200,N_4680);
nor U7543 (N_7543,N_3703,N_5657);
or U7544 (N_7544,N_4755,N_5101);
or U7545 (N_7545,N_4856,N_4453);
and U7546 (N_7546,N_3360,N_5609);
nor U7547 (N_7547,N_5882,N_5953);
or U7548 (N_7548,N_4240,N_4264);
xor U7549 (N_7549,N_4615,N_4489);
and U7550 (N_7550,N_4750,N_4165);
nor U7551 (N_7551,N_3433,N_4400);
nand U7552 (N_7552,N_6167,N_4565);
nand U7553 (N_7553,N_5818,N_3747);
or U7554 (N_7554,N_3249,N_6144);
nor U7555 (N_7555,N_3848,N_6179);
or U7556 (N_7556,N_3193,N_4385);
and U7557 (N_7557,N_3150,N_3390);
nor U7558 (N_7558,N_4317,N_6232);
xor U7559 (N_7559,N_4743,N_3500);
nand U7560 (N_7560,N_3136,N_3273);
nand U7561 (N_7561,N_4724,N_3442);
nor U7562 (N_7562,N_4549,N_3792);
xor U7563 (N_7563,N_3351,N_5835);
nand U7564 (N_7564,N_4265,N_5865);
nor U7565 (N_7565,N_3773,N_3738);
nor U7566 (N_7566,N_6197,N_3881);
nand U7567 (N_7567,N_5660,N_5082);
or U7568 (N_7568,N_4645,N_5255);
nand U7569 (N_7569,N_5334,N_4282);
nor U7570 (N_7570,N_3204,N_3909);
nand U7571 (N_7571,N_5624,N_3217);
nor U7572 (N_7572,N_3264,N_5142);
nand U7573 (N_7573,N_6176,N_3301);
nand U7574 (N_7574,N_4092,N_6148);
or U7575 (N_7575,N_3358,N_3670);
nand U7576 (N_7576,N_3462,N_3664);
nand U7577 (N_7577,N_5774,N_4414);
and U7578 (N_7578,N_5467,N_4699);
or U7579 (N_7579,N_4526,N_5344);
nand U7580 (N_7580,N_4973,N_5873);
or U7581 (N_7581,N_5661,N_4980);
and U7582 (N_7582,N_5141,N_4968);
nand U7583 (N_7583,N_4352,N_3723);
nand U7584 (N_7584,N_4493,N_4554);
or U7585 (N_7585,N_4498,N_3572);
nor U7586 (N_7586,N_3757,N_5576);
xor U7587 (N_7587,N_3422,N_4678);
xnor U7588 (N_7588,N_4849,N_4714);
xor U7589 (N_7589,N_4189,N_5196);
or U7590 (N_7590,N_5297,N_4759);
nand U7591 (N_7591,N_3133,N_5932);
nand U7592 (N_7592,N_3481,N_3487);
nand U7593 (N_7593,N_5856,N_4733);
xnor U7594 (N_7594,N_4474,N_5597);
and U7595 (N_7595,N_5635,N_3317);
or U7596 (N_7596,N_4383,N_3215);
nor U7597 (N_7597,N_4062,N_4664);
and U7598 (N_7598,N_3979,N_4225);
or U7599 (N_7599,N_4123,N_3533);
or U7600 (N_7600,N_3822,N_3353);
and U7601 (N_7601,N_5688,N_4754);
or U7602 (N_7602,N_4469,N_5514);
and U7603 (N_7603,N_3710,N_5844);
nand U7604 (N_7604,N_5084,N_5887);
nor U7605 (N_7605,N_5304,N_4088);
or U7606 (N_7606,N_3186,N_5248);
and U7607 (N_7607,N_5613,N_5831);
or U7608 (N_7608,N_5880,N_4826);
nand U7609 (N_7609,N_4512,N_4583);
nand U7610 (N_7610,N_5190,N_3350);
nand U7611 (N_7611,N_4637,N_6231);
nand U7612 (N_7612,N_6211,N_5602);
nor U7613 (N_7613,N_4146,N_5777);
nor U7614 (N_7614,N_4947,N_4132);
and U7615 (N_7615,N_5822,N_6173);
and U7616 (N_7616,N_5329,N_5037);
or U7617 (N_7617,N_4739,N_4648);
and U7618 (N_7618,N_4705,N_4631);
or U7619 (N_7619,N_4125,N_4133);
nor U7620 (N_7620,N_3978,N_4432);
nor U7621 (N_7621,N_4954,N_5154);
nand U7622 (N_7622,N_5562,N_5477);
or U7623 (N_7623,N_6135,N_3223);
xnor U7624 (N_7624,N_4813,N_4420);
nor U7625 (N_7625,N_3835,N_3235);
and U7626 (N_7626,N_5595,N_6093);
nand U7627 (N_7627,N_5941,N_4868);
or U7628 (N_7628,N_4052,N_4012);
nand U7629 (N_7629,N_3272,N_3451);
nand U7630 (N_7630,N_5316,N_5059);
and U7631 (N_7631,N_5674,N_5318);
nor U7632 (N_7632,N_3900,N_4281);
nor U7633 (N_7633,N_5144,N_5837);
nand U7634 (N_7634,N_4510,N_6123);
nor U7635 (N_7635,N_3206,N_5020);
nor U7636 (N_7636,N_4262,N_3275);
nor U7637 (N_7637,N_3642,N_3895);
nand U7638 (N_7638,N_3893,N_3987);
and U7639 (N_7639,N_5495,N_4455);
or U7640 (N_7640,N_5552,N_3576);
nand U7641 (N_7641,N_5167,N_4169);
xnor U7642 (N_7642,N_5813,N_5124);
and U7643 (N_7643,N_4041,N_5028);
xor U7644 (N_7644,N_4540,N_5644);
nor U7645 (N_7645,N_3361,N_5881);
and U7646 (N_7646,N_5390,N_3509);
and U7647 (N_7647,N_4641,N_5038);
or U7648 (N_7648,N_3951,N_3211);
and U7649 (N_7649,N_3696,N_5484);
nor U7650 (N_7650,N_4158,N_4036);
nand U7651 (N_7651,N_3782,N_4362);
nor U7652 (N_7652,N_5461,N_4882);
and U7653 (N_7653,N_5528,N_4671);
nand U7654 (N_7654,N_5891,N_4770);
or U7655 (N_7655,N_5687,N_3364);
or U7656 (N_7656,N_3450,N_3488);
nand U7657 (N_7657,N_3936,N_3280);
nor U7658 (N_7658,N_4075,N_6133);
nand U7659 (N_7659,N_5320,N_5447);
or U7660 (N_7660,N_3382,N_4528);
nor U7661 (N_7661,N_4449,N_4068);
xnor U7662 (N_7662,N_5287,N_3748);
nand U7663 (N_7663,N_3470,N_5192);
xnor U7664 (N_7664,N_4033,N_4181);
and U7665 (N_7665,N_4299,N_6137);
or U7666 (N_7666,N_4371,N_5365);
or U7667 (N_7667,N_3608,N_3502);
xnor U7668 (N_7668,N_3653,N_6204);
nand U7669 (N_7669,N_4749,N_5872);
nor U7670 (N_7670,N_4753,N_3974);
xnor U7671 (N_7671,N_5193,N_5388);
nand U7672 (N_7672,N_6100,N_4066);
and U7673 (N_7673,N_4087,N_4347);
and U7674 (N_7674,N_4417,N_4686);
or U7675 (N_7675,N_3720,N_4373);
nand U7676 (N_7676,N_5078,N_4050);
and U7677 (N_7677,N_4304,N_4435);
nor U7678 (N_7678,N_4178,N_5976);
or U7679 (N_7679,N_5619,N_6212);
and U7680 (N_7680,N_5441,N_5145);
and U7681 (N_7681,N_6143,N_4567);
xor U7682 (N_7682,N_5943,N_6029);
nand U7683 (N_7683,N_4523,N_4892);
nor U7684 (N_7684,N_4552,N_3397);
or U7685 (N_7685,N_3227,N_5387);
or U7686 (N_7686,N_3435,N_4595);
xnor U7687 (N_7687,N_5002,N_6151);
nor U7688 (N_7688,N_3905,N_4457);
nand U7689 (N_7689,N_3725,N_5428);
or U7690 (N_7690,N_4815,N_5770);
or U7691 (N_7691,N_5919,N_5198);
nand U7692 (N_7692,N_5747,N_5748);
xnor U7693 (N_7693,N_5014,N_5043);
nor U7694 (N_7694,N_3504,N_5413);
or U7695 (N_7695,N_4684,N_5715);
or U7696 (N_7696,N_4551,N_3392);
nand U7697 (N_7697,N_5704,N_6190);
or U7698 (N_7698,N_6141,N_4694);
or U7699 (N_7699,N_5176,N_3887);
nor U7700 (N_7700,N_6217,N_4289);
xor U7701 (N_7701,N_5324,N_4406);
nor U7702 (N_7702,N_5158,N_3130);
nand U7703 (N_7703,N_4048,N_5618);
or U7704 (N_7704,N_5342,N_4652);
and U7705 (N_7705,N_5729,N_5558);
nor U7706 (N_7706,N_3850,N_4307);
and U7707 (N_7707,N_5975,N_6185);
nor U7708 (N_7708,N_5228,N_6200);
xnor U7709 (N_7709,N_5416,N_5978);
nand U7710 (N_7710,N_6223,N_5633);
nand U7711 (N_7711,N_3388,N_5526);
or U7712 (N_7712,N_4266,N_5512);
or U7713 (N_7713,N_5290,N_3766);
or U7714 (N_7714,N_5395,N_5185);
or U7715 (N_7715,N_3412,N_3948);
nand U7716 (N_7716,N_4795,N_4886);
or U7717 (N_7717,N_5723,N_5354);
or U7718 (N_7718,N_5504,N_3455);
and U7719 (N_7719,N_3937,N_5138);
and U7720 (N_7720,N_4865,N_4797);
and U7721 (N_7721,N_4858,N_5473);
or U7722 (N_7722,N_5247,N_4949);
nand U7723 (N_7723,N_4669,N_3592);
nand U7724 (N_7724,N_6095,N_3181);
nor U7725 (N_7725,N_3928,N_4298);
and U7726 (N_7726,N_5820,N_6168);
or U7727 (N_7727,N_5610,N_5956);
nand U7728 (N_7728,N_3183,N_3988);
xnor U7729 (N_7729,N_4404,N_5782);
and U7730 (N_7730,N_4619,N_5446);
or U7731 (N_7731,N_5410,N_3421);
nor U7732 (N_7732,N_6101,N_4965);
and U7733 (N_7733,N_5216,N_5243);
or U7734 (N_7734,N_3658,N_5088);
nor U7735 (N_7735,N_5665,N_5245);
nor U7736 (N_7736,N_4368,N_5421);
nor U7737 (N_7737,N_3484,N_3707);
xnor U7738 (N_7738,N_5781,N_4153);
or U7739 (N_7739,N_6242,N_4185);
or U7740 (N_7740,N_4522,N_4704);
nand U7741 (N_7741,N_3906,N_3594);
and U7742 (N_7742,N_3331,N_3603);
nor U7743 (N_7743,N_4840,N_3913);
xor U7744 (N_7744,N_4651,N_4434);
nor U7745 (N_7745,N_3671,N_3790);
or U7746 (N_7746,N_5482,N_3654);
and U7747 (N_7747,N_5063,N_4105);
or U7748 (N_7748,N_6085,N_5276);
nor U7749 (N_7749,N_3281,N_3946);
and U7750 (N_7750,N_5531,N_3823);
and U7751 (N_7751,N_5763,N_3535);
or U7752 (N_7752,N_5640,N_4043);
nand U7753 (N_7753,N_3886,N_4472);
and U7754 (N_7754,N_3775,N_4393);
nor U7755 (N_7755,N_3292,N_3986);
nor U7756 (N_7756,N_3497,N_3853);
or U7757 (N_7757,N_4517,N_5219);
and U7758 (N_7758,N_6039,N_5855);
and U7759 (N_7759,N_4034,N_4233);
xor U7760 (N_7760,N_5215,N_4604);
nor U7761 (N_7761,N_4990,N_5767);
nand U7762 (N_7762,N_5485,N_3228);
nor U7763 (N_7763,N_4966,N_4224);
nor U7764 (N_7764,N_3939,N_5301);
or U7765 (N_7765,N_4440,N_6064);
nor U7766 (N_7766,N_3729,N_4613);
nand U7767 (N_7767,N_6068,N_3289);
nor U7768 (N_7768,N_5237,N_5027);
and U7769 (N_7769,N_4188,N_4818);
and U7770 (N_7770,N_4929,N_5347);
nor U7771 (N_7771,N_3197,N_3569);
xnor U7772 (N_7772,N_5127,N_5208);
nor U7773 (N_7773,N_5736,N_4270);
xor U7774 (N_7774,N_3971,N_3722);
nor U7775 (N_7775,N_4777,N_5766);
nor U7776 (N_7776,N_4447,N_5987);
nor U7777 (N_7777,N_4574,N_4330);
nor U7778 (N_7778,N_3176,N_4874);
or U7779 (N_7779,N_5507,N_4064);
or U7780 (N_7780,N_5861,N_4644);
nand U7781 (N_7781,N_3623,N_6201);
or U7782 (N_7782,N_3226,N_3546);
nand U7783 (N_7783,N_5984,N_4710);
or U7784 (N_7784,N_4539,N_3679);
nor U7785 (N_7785,N_3177,N_3755);
nand U7786 (N_7786,N_3622,N_3326);
nand U7787 (N_7787,N_5849,N_3796);
nor U7788 (N_7788,N_5235,N_4046);
nand U7789 (N_7789,N_5412,N_4001);
nand U7790 (N_7790,N_6094,N_3645);
nor U7791 (N_7791,N_4422,N_5405);
nand U7792 (N_7792,N_5025,N_4993);
or U7793 (N_7793,N_5692,N_4776);
nand U7794 (N_7794,N_5375,N_4809);
xnor U7795 (N_7795,N_5769,N_3501);
xor U7796 (N_7796,N_3251,N_4951);
nand U7797 (N_7797,N_5544,N_6055);
and U7798 (N_7798,N_3224,N_6006);
and U7799 (N_7799,N_3332,N_5515);
and U7800 (N_7800,N_4975,N_3692);
nand U7801 (N_7801,N_3199,N_3529);
and U7802 (N_7802,N_5325,N_4642);
nor U7803 (N_7803,N_4384,N_5895);
nor U7804 (N_7804,N_3423,N_5293);
and U7805 (N_7805,N_6008,N_3838);
nor U7806 (N_7806,N_3924,N_6042);
or U7807 (N_7807,N_5718,N_3342);
nand U7808 (N_7808,N_3655,N_4206);
or U7809 (N_7809,N_4721,N_3690);
or U7810 (N_7810,N_5366,N_3935);
or U7811 (N_7811,N_5475,N_5875);
nand U7812 (N_7812,N_4290,N_5163);
and U7813 (N_7813,N_5402,N_4118);
and U7814 (N_7814,N_4646,N_5848);
nor U7815 (N_7815,N_5250,N_4591);
nand U7816 (N_7816,N_5807,N_4073);
nand U7817 (N_7817,N_4552,N_5986);
nand U7818 (N_7818,N_3224,N_4247);
nor U7819 (N_7819,N_4635,N_6216);
and U7820 (N_7820,N_3861,N_4353);
and U7821 (N_7821,N_3836,N_4834);
and U7822 (N_7822,N_4532,N_4427);
or U7823 (N_7823,N_5724,N_4805);
nand U7824 (N_7824,N_6246,N_5504);
nor U7825 (N_7825,N_5213,N_5751);
nand U7826 (N_7826,N_6133,N_5337);
nand U7827 (N_7827,N_4242,N_3266);
xor U7828 (N_7828,N_4422,N_3538);
and U7829 (N_7829,N_3885,N_3886);
and U7830 (N_7830,N_5100,N_5446);
or U7831 (N_7831,N_3747,N_5984);
nor U7832 (N_7832,N_4681,N_4238);
nand U7833 (N_7833,N_5797,N_3960);
and U7834 (N_7834,N_3510,N_5498);
nor U7835 (N_7835,N_4903,N_3687);
nand U7836 (N_7836,N_4200,N_5639);
and U7837 (N_7837,N_4457,N_5269);
nand U7838 (N_7838,N_4077,N_5696);
or U7839 (N_7839,N_5499,N_4344);
nor U7840 (N_7840,N_4927,N_5150);
or U7841 (N_7841,N_3801,N_5649);
or U7842 (N_7842,N_4994,N_3527);
or U7843 (N_7843,N_4835,N_5425);
or U7844 (N_7844,N_3972,N_3544);
nor U7845 (N_7845,N_3632,N_3379);
and U7846 (N_7846,N_3154,N_3437);
or U7847 (N_7847,N_6082,N_4741);
nand U7848 (N_7848,N_4496,N_4852);
xor U7849 (N_7849,N_5526,N_4088);
nand U7850 (N_7850,N_4114,N_3254);
and U7851 (N_7851,N_6188,N_3415);
or U7852 (N_7852,N_4203,N_3263);
nand U7853 (N_7853,N_6172,N_3713);
and U7854 (N_7854,N_5090,N_3133);
and U7855 (N_7855,N_3736,N_3467);
nand U7856 (N_7856,N_4398,N_3528);
xor U7857 (N_7857,N_4688,N_5550);
nor U7858 (N_7858,N_6167,N_4767);
or U7859 (N_7859,N_4315,N_4216);
nor U7860 (N_7860,N_5363,N_5486);
and U7861 (N_7861,N_4031,N_6221);
nand U7862 (N_7862,N_5561,N_4367);
nor U7863 (N_7863,N_5232,N_4709);
nor U7864 (N_7864,N_5003,N_3639);
or U7865 (N_7865,N_4073,N_3349);
or U7866 (N_7866,N_5004,N_3732);
nor U7867 (N_7867,N_3128,N_5372);
xor U7868 (N_7868,N_4780,N_5342);
nor U7869 (N_7869,N_5544,N_5047);
nand U7870 (N_7870,N_4256,N_6074);
and U7871 (N_7871,N_3439,N_4659);
or U7872 (N_7872,N_5645,N_3257);
and U7873 (N_7873,N_5360,N_3838);
and U7874 (N_7874,N_4648,N_4519);
nand U7875 (N_7875,N_4080,N_3356);
nand U7876 (N_7876,N_3540,N_3740);
and U7877 (N_7877,N_4878,N_4367);
or U7878 (N_7878,N_3294,N_4311);
or U7879 (N_7879,N_4137,N_4121);
nand U7880 (N_7880,N_3548,N_5618);
or U7881 (N_7881,N_5007,N_3408);
or U7882 (N_7882,N_4497,N_5701);
nor U7883 (N_7883,N_4814,N_6116);
or U7884 (N_7884,N_5796,N_5334);
nand U7885 (N_7885,N_3907,N_5231);
or U7886 (N_7886,N_4423,N_4717);
nand U7887 (N_7887,N_5781,N_5048);
nand U7888 (N_7888,N_4317,N_5550);
nor U7889 (N_7889,N_3258,N_3806);
and U7890 (N_7890,N_4730,N_4930);
and U7891 (N_7891,N_4641,N_3722);
or U7892 (N_7892,N_5983,N_4585);
and U7893 (N_7893,N_4358,N_4846);
xnor U7894 (N_7894,N_5094,N_3320);
and U7895 (N_7895,N_5342,N_4608);
nor U7896 (N_7896,N_3475,N_3248);
or U7897 (N_7897,N_3819,N_6063);
nand U7898 (N_7898,N_3223,N_3681);
or U7899 (N_7899,N_5326,N_3549);
xor U7900 (N_7900,N_5946,N_3756);
nand U7901 (N_7901,N_5419,N_3635);
nor U7902 (N_7902,N_4879,N_3272);
or U7903 (N_7903,N_5523,N_4587);
nand U7904 (N_7904,N_5308,N_4355);
and U7905 (N_7905,N_4669,N_5045);
nor U7906 (N_7906,N_6224,N_4572);
nand U7907 (N_7907,N_5462,N_5208);
or U7908 (N_7908,N_4561,N_4289);
nand U7909 (N_7909,N_5851,N_3561);
xnor U7910 (N_7910,N_3893,N_3333);
and U7911 (N_7911,N_4569,N_3352);
or U7912 (N_7912,N_4028,N_4944);
and U7913 (N_7913,N_3865,N_4638);
nor U7914 (N_7914,N_4636,N_3683);
nor U7915 (N_7915,N_5884,N_3645);
or U7916 (N_7916,N_5543,N_3848);
nand U7917 (N_7917,N_5977,N_3773);
xnor U7918 (N_7918,N_5825,N_3649);
nor U7919 (N_7919,N_5674,N_4538);
nor U7920 (N_7920,N_3516,N_3409);
nor U7921 (N_7921,N_4725,N_3408);
nand U7922 (N_7922,N_3486,N_4656);
or U7923 (N_7923,N_5886,N_3779);
nand U7924 (N_7924,N_5195,N_3612);
or U7925 (N_7925,N_4599,N_5927);
nor U7926 (N_7926,N_3985,N_3974);
and U7927 (N_7927,N_5329,N_3395);
xor U7928 (N_7928,N_5221,N_3686);
xor U7929 (N_7929,N_4141,N_3299);
xor U7930 (N_7930,N_5275,N_5321);
and U7931 (N_7931,N_5011,N_3126);
nor U7932 (N_7932,N_5358,N_5101);
or U7933 (N_7933,N_6071,N_5618);
or U7934 (N_7934,N_5502,N_4067);
or U7935 (N_7935,N_3920,N_5771);
xnor U7936 (N_7936,N_5384,N_5121);
nor U7937 (N_7937,N_3962,N_3748);
nor U7938 (N_7938,N_4584,N_4317);
xor U7939 (N_7939,N_5145,N_3439);
nand U7940 (N_7940,N_3705,N_3972);
nor U7941 (N_7941,N_5971,N_5548);
or U7942 (N_7942,N_4580,N_3219);
or U7943 (N_7943,N_4525,N_5120);
and U7944 (N_7944,N_6043,N_6161);
or U7945 (N_7945,N_5650,N_4706);
nand U7946 (N_7946,N_4408,N_5872);
nor U7947 (N_7947,N_6171,N_3707);
and U7948 (N_7948,N_5103,N_6068);
nand U7949 (N_7949,N_4422,N_4902);
nand U7950 (N_7950,N_3285,N_5158);
nor U7951 (N_7951,N_5931,N_6001);
nand U7952 (N_7952,N_5666,N_5158);
nor U7953 (N_7953,N_4919,N_3227);
nand U7954 (N_7954,N_5899,N_4982);
and U7955 (N_7955,N_5282,N_5129);
or U7956 (N_7956,N_5952,N_5808);
nand U7957 (N_7957,N_4030,N_3861);
nand U7958 (N_7958,N_6160,N_4378);
nand U7959 (N_7959,N_5560,N_6024);
nor U7960 (N_7960,N_5944,N_4949);
nor U7961 (N_7961,N_3678,N_4007);
xor U7962 (N_7962,N_4499,N_3224);
or U7963 (N_7963,N_3452,N_6096);
nor U7964 (N_7964,N_4458,N_4407);
or U7965 (N_7965,N_5009,N_4453);
xnor U7966 (N_7966,N_4360,N_5905);
nor U7967 (N_7967,N_5920,N_3422);
and U7968 (N_7968,N_4533,N_4173);
and U7969 (N_7969,N_5730,N_3951);
nand U7970 (N_7970,N_4823,N_6218);
and U7971 (N_7971,N_3633,N_4138);
or U7972 (N_7972,N_4752,N_4700);
and U7973 (N_7973,N_3206,N_5476);
and U7974 (N_7974,N_5965,N_4483);
xor U7975 (N_7975,N_5033,N_3306);
nand U7976 (N_7976,N_4368,N_4031);
nor U7977 (N_7977,N_5220,N_5382);
and U7978 (N_7978,N_3232,N_3254);
and U7979 (N_7979,N_5878,N_5505);
and U7980 (N_7980,N_5689,N_4547);
nand U7981 (N_7981,N_5699,N_3211);
and U7982 (N_7982,N_4001,N_4383);
xnor U7983 (N_7983,N_4593,N_3314);
nand U7984 (N_7984,N_4503,N_3525);
nor U7985 (N_7985,N_5876,N_6094);
xor U7986 (N_7986,N_3427,N_5792);
nand U7987 (N_7987,N_5716,N_3625);
or U7988 (N_7988,N_4468,N_4312);
and U7989 (N_7989,N_3696,N_6228);
or U7990 (N_7990,N_5913,N_5709);
and U7991 (N_7991,N_3125,N_3789);
nand U7992 (N_7992,N_4672,N_4671);
nand U7993 (N_7993,N_3668,N_5527);
or U7994 (N_7994,N_4644,N_5611);
or U7995 (N_7995,N_5520,N_5100);
and U7996 (N_7996,N_5647,N_3941);
nor U7997 (N_7997,N_3736,N_5252);
and U7998 (N_7998,N_4321,N_4071);
nor U7999 (N_7999,N_5380,N_5112);
nor U8000 (N_8000,N_4230,N_5876);
or U8001 (N_8001,N_4325,N_5778);
nor U8002 (N_8002,N_4712,N_4387);
and U8003 (N_8003,N_3324,N_6014);
nand U8004 (N_8004,N_3501,N_5336);
xor U8005 (N_8005,N_3967,N_5073);
xor U8006 (N_8006,N_4504,N_5926);
nor U8007 (N_8007,N_3886,N_3844);
and U8008 (N_8008,N_3988,N_3758);
nand U8009 (N_8009,N_5153,N_4202);
or U8010 (N_8010,N_5087,N_5736);
xnor U8011 (N_8011,N_3395,N_4002);
nor U8012 (N_8012,N_4067,N_4388);
nor U8013 (N_8013,N_4374,N_3707);
or U8014 (N_8014,N_5507,N_4809);
xor U8015 (N_8015,N_4152,N_5029);
or U8016 (N_8016,N_4776,N_5702);
xnor U8017 (N_8017,N_4315,N_4946);
or U8018 (N_8018,N_5981,N_4710);
or U8019 (N_8019,N_3125,N_3703);
nand U8020 (N_8020,N_3956,N_3777);
xnor U8021 (N_8021,N_4403,N_6178);
nor U8022 (N_8022,N_5240,N_4951);
nor U8023 (N_8023,N_3547,N_5057);
nor U8024 (N_8024,N_5455,N_3576);
nor U8025 (N_8025,N_6149,N_4591);
xor U8026 (N_8026,N_3772,N_4792);
nand U8027 (N_8027,N_3627,N_3174);
xnor U8028 (N_8028,N_3659,N_4365);
or U8029 (N_8029,N_6233,N_5111);
nor U8030 (N_8030,N_4204,N_5127);
and U8031 (N_8031,N_3246,N_5804);
nand U8032 (N_8032,N_3673,N_4866);
nand U8033 (N_8033,N_3411,N_4724);
nor U8034 (N_8034,N_3868,N_5385);
nand U8035 (N_8035,N_6116,N_5501);
nor U8036 (N_8036,N_5909,N_3218);
nand U8037 (N_8037,N_4531,N_5457);
or U8038 (N_8038,N_3289,N_3932);
and U8039 (N_8039,N_4264,N_5228);
or U8040 (N_8040,N_3455,N_5201);
xor U8041 (N_8041,N_4294,N_6085);
nor U8042 (N_8042,N_4690,N_6090);
nor U8043 (N_8043,N_4817,N_4040);
and U8044 (N_8044,N_4257,N_4658);
or U8045 (N_8045,N_5149,N_5253);
or U8046 (N_8046,N_3249,N_5431);
or U8047 (N_8047,N_6181,N_4263);
and U8048 (N_8048,N_3849,N_3442);
or U8049 (N_8049,N_5868,N_3709);
or U8050 (N_8050,N_3630,N_5824);
and U8051 (N_8051,N_5291,N_4656);
or U8052 (N_8052,N_6202,N_5353);
nand U8053 (N_8053,N_4091,N_5762);
and U8054 (N_8054,N_4913,N_3970);
xor U8055 (N_8055,N_5959,N_3146);
or U8056 (N_8056,N_6234,N_3225);
or U8057 (N_8057,N_5495,N_3179);
xor U8058 (N_8058,N_5515,N_4021);
or U8059 (N_8059,N_3938,N_3192);
xor U8060 (N_8060,N_4824,N_3644);
nor U8061 (N_8061,N_5698,N_5220);
or U8062 (N_8062,N_3581,N_3865);
or U8063 (N_8063,N_5008,N_5774);
nor U8064 (N_8064,N_4126,N_4002);
nor U8065 (N_8065,N_4121,N_4048);
nand U8066 (N_8066,N_5568,N_3306);
or U8067 (N_8067,N_4441,N_4413);
and U8068 (N_8068,N_3249,N_4090);
nand U8069 (N_8069,N_5376,N_5805);
nor U8070 (N_8070,N_5452,N_3402);
nand U8071 (N_8071,N_5037,N_5999);
nand U8072 (N_8072,N_4438,N_5760);
nand U8073 (N_8073,N_5407,N_4673);
nand U8074 (N_8074,N_3821,N_3987);
nand U8075 (N_8075,N_5583,N_4493);
and U8076 (N_8076,N_5859,N_3548);
nand U8077 (N_8077,N_3215,N_4749);
nand U8078 (N_8078,N_5492,N_6057);
nor U8079 (N_8079,N_4386,N_4957);
nand U8080 (N_8080,N_5428,N_3527);
nor U8081 (N_8081,N_5450,N_6041);
and U8082 (N_8082,N_5457,N_3992);
nor U8083 (N_8083,N_4220,N_3416);
xnor U8084 (N_8084,N_5731,N_5226);
and U8085 (N_8085,N_5397,N_5737);
nor U8086 (N_8086,N_5638,N_5938);
or U8087 (N_8087,N_4714,N_3347);
and U8088 (N_8088,N_4351,N_3150);
and U8089 (N_8089,N_3533,N_3806);
xnor U8090 (N_8090,N_3300,N_4824);
or U8091 (N_8091,N_4320,N_5363);
and U8092 (N_8092,N_5083,N_4724);
or U8093 (N_8093,N_4828,N_4280);
and U8094 (N_8094,N_4997,N_4361);
nor U8095 (N_8095,N_4291,N_3444);
nand U8096 (N_8096,N_4256,N_4628);
nand U8097 (N_8097,N_4616,N_5184);
nand U8098 (N_8098,N_4580,N_4480);
nand U8099 (N_8099,N_4429,N_4983);
xnor U8100 (N_8100,N_5318,N_3888);
or U8101 (N_8101,N_6041,N_4799);
nand U8102 (N_8102,N_4848,N_5450);
and U8103 (N_8103,N_4225,N_6122);
nand U8104 (N_8104,N_3612,N_6131);
and U8105 (N_8105,N_3598,N_4201);
and U8106 (N_8106,N_3286,N_5729);
nor U8107 (N_8107,N_5721,N_5782);
nor U8108 (N_8108,N_3713,N_5805);
nor U8109 (N_8109,N_3133,N_4082);
nand U8110 (N_8110,N_3996,N_3740);
nand U8111 (N_8111,N_4050,N_5118);
xor U8112 (N_8112,N_4216,N_4579);
nand U8113 (N_8113,N_4857,N_3404);
nor U8114 (N_8114,N_5364,N_3727);
and U8115 (N_8115,N_4087,N_3229);
nor U8116 (N_8116,N_5309,N_5393);
nor U8117 (N_8117,N_5704,N_5706);
and U8118 (N_8118,N_6236,N_5647);
nand U8119 (N_8119,N_4593,N_5617);
nand U8120 (N_8120,N_3936,N_5218);
and U8121 (N_8121,N_4019,N_5873);
nor U8122 (N_8122,N_6143,N_4472);
and U8123 (N_8123,N_5097,N_3992);
nand U8124 (N_8124,N_4962,N_4228);
nor U8125 (N_8125,N_4596,N_4521);
nand U8126 (N_8126,N_3154,N_5957);
or U8127 (N_8127,N_4774,N_5257);
nor U8128 (N_8128,N_5189,N_4472);
nand U8129 (N_8129,N_6022,N_6079);
xor U8130 (N_8130,N_6006,N_3760);
or U8131 (N_8131,N_4951,N_3248);
and U8132 (N_8132,N_5548,N_3709);
nor U8133 (N_8133,N_5243,N_4735);
nand U8134 (N_8134,N_3404,N_3745);
or U8135 (N_8135,N_6041,N_5401);
nand U8136 (N_8136,N_5456,N_4333);
nor U8137 (N_8137,N_4190,N_5363);
and U8138 (N_8138,N_5843,N_4238);
nor U8139 (N_8139,N_5477,N_5222);
or U8140 (N_8140,N_5819,N_4597);
nor U8141 (N_8141,N_3472,N_3915);
or U8142 (N_8142,N_4217,N_4299);
or U8143 (N_8143,N_6147,N_4221);
and U8144 (N_8144,N_3229,N_5302);
or U8145 (N_8145,N_5084,N_3812);
xor U8146 (N_8146,N_5665,N_5916);
nand U8147 (N_8147,N_4328,N_5058);
and U8148 (N_8148,N_4527,N_4348);
xnor U8149 (N_8149,N_6016,N_4758);
and U8150 (N_8150,N_4014,N_4026);
nand U8151 (N_8151,N_4941,N_5716);
nand U8152 (N_8152,N_6006,N_3326);
nor U8153 (N_8153,N_6231,N_3892);
nor U8154 (N_8154,N_5061,N_4363);
and U8155 (N_8155,N_5695,N_4879);
nor U8156 (N_8156,N_4419,N_3607);
xnor U8157 (N_8157,N_4487,N_5744);
nand U8158 (N_8158,N_4588,N_5584);
or U8159 (N_8159,N_6045,N_4366);
or U8160 (N_8160,N_5094,N_4131);
or U8161 (N_8161,N_3794,N_3716);
or U8162 (N_8162,N_3957,N_3288);
nor U8163 (N_8163,N_4295,N_3552);
nor U8164 (N_8164,N_5865,N_5891);
nor U8165 (N_8165,N_6098,N_3305);
nand U8166 (N_8166,N_4194,N_4445);
nand U8167 (N_8167,N_3607,N_4274);
nand U8168 (N_8168,N_3267,N_4801);
nand U8169 (N_8169,N_4935,N_4104);
nand U8170 (N_8170,N_5643,N_4818);
and U8171 (N_8171,N_5111,N_5870);
nand U8172 (N_8172,N_6230,N_5925);
and U8173 (N_8173,N_5423,N_5582);
nand U8174 (N_8174,N_5664,N_5590);
nor U8175 (N_8175,N_3716,N_5361);
nand U8176 (N_8176,N_5699,N_3765);
or U8177 (N_8177,N_4328,N_5779);
or U8178 (N_8178,N_5472,N_3920);
nand U8179 (N_8179,N_4433,N_3288);
and U8180 (N_8180,N_5089,N_5478);
nor U8181 (N_8181,N_4560,N_3443);
xor U8182 (N_8182,N_4038,N_5565);
or U8183 (N_8183,N_3716,N_5353);
nand U8184 (N_8184,N_4314,N_6168);
nand U8185 (N_8185,N_4516,N_4490);
nor U8186 (N_8186,N_3903,N_5487);
nor U8187 (N_8187,N_5706,N_5106);
or U8188 (N_8188,N_3353,N_4797);
nor U8189 (N_8189,N_5473,N_3497);
or U8190 (N_8190,N_5660,N_3143);
xor U8191 (N_8191,N_5716,N_5198);
and U8192 (N_8192,N_5932,N_5002);
nor U8193 (N_8193,N_3741,N_5882);
xor U8194 (N_8194,N_6029,N_5004);
and U8195 (N_8195,N_4367,N_4435);
nand U8196 (N_8196,N_4301,N_3553);
nand U8197 (N_8197,N_5757,N_6046);
or U8198 (N_8198,N_5651,N_4024);
and U8199 (N_8199,N_3623,N_5204);
nor U8200 (N_8200,N_4526,N_5781);
nor U8201 (N_8201,N_3272,N_4752);
xor U8202 (N_8202,N_4994,N_5630);
nor U8203 (N_8203,N_5181,N_3619);
nor U8204 (N_8204,N_4440,N_5446);
or U8205 (N_8205,N_4325,N_5958);
nand U8206 (N_8206,N_3904,N_5248);
nand U8207 (N_8207,N_3470,N_6127);
nor U8208 (N_8208,N_3486,N_6186);
and U8209 (N_8209,N_5679,N_5932);
and U8210 (N_8210,N_3648,N_4705);
or U8211 (N_8211,N_5392,N_5881);
nand U8212 (N_8212,N_4512,N_5894);
nand U8213 (N_8213,N_4409,N_4898);
nand U8214 (N_8214,N_4689,N_5106);
nor U8215 (N_8215,N_3534,N_3400);
nand U8216 (N_8216,N_5680,N_4087);
or U8217 (N_8217,N_5285,N_5397);
or U8218 (N_8218,N_5885,N_3350);
or U8219 (N_8219,N_5837,N_4805);
nor U8220 (N_8220,N_3657,N_6021);
nand U8221 (N_8221,N_5522,N_3440);
nor U8222 (N_8222,N_4675,N_5344);
and U8223 (N_8223,N_5227,N_6029);
xor U8224 (N_8224,N_5167,N_4661);
or U8225 (N_8225,N_3584,N_5759);
xor U8226 (N_8226,N_5343,N_5913);
nand U8227 (N_8227,N_3287,N_3633);
or U8228 (N_8228,N_4646,N_4142);
or U8229 (N_8229,N_4153,N_6144);
and U8230 (N_8230,N_4647,N_4778);
and U8231 (N_8231,N_4627,N_3673);
and U8232 (N_8232,N_5365,N_3793);
nor U8233 (N_8233,N_4837,N_4946);
nand U8234 (N_8234,N_6079,N_6092);
nand U8235 (N_8235,N_4994,N_3611);
nand U8236 (N_8236,N_3988,N_4969);
or U8237 (N_8237,N_5696,N_5419);
nand U8238 (N_8238,N_3734,N_3260);
nand U8239 (N_8239,N_5769,N_6213);
and U8240 (N_8240,N_4409,N_3630);
or U8241 (N_8241,N_4613,N_6060);
nand U8242 (N_8242,N_3914,N_5722);
xnor U8243 (N_8243,N_6218,N_4721);
or U8244 (N_8244,N_4566,N_4955);
nand U8245 (N_8245,N_4222,N_4932);
and U8246 (N_8246,N_4654,N_3867);
nor U8247 (N_8247,N_5787,N_5840);
nand U8248 (N_8248,N_4789,N_3797);
nor U8249 (N_8249,N_4227,N_5764);
and U8250 (N_8250,N_3596,N_3523);
and U8251 (N_8251,N_4361,N_4647);
or U8252 (N_8252,N_3229,N_4691);
and U8253 (N_8253,N_4899,N_5395);
nand U8254 (N_8254,N_3186,N_3865);
or U8255 (N_8255,N_3324,N_3207);
xnor U8256 (N_8256,N_5897,N_3858);
and U8257 (N_8257,N_4976,N_5016);
or U8258 (N_8258,N_6241,N_3719);
nor U8259 (N_8259,N_3438,N_6119);
xnor U8260 (N_8260,N_3696,N_3777);
nor U8261 (N_8261,N_3296,N_5164);
or U8262 (N_8262,N_6208,N_6170);
nand U8263 (N_8263,N_5712,N_5685);
and U8264 (N_8264,N_4415,N_5354);
or U8265 (N_8265,N_4944,N_3139);
and U8266 (N_8266,N_4319,N_4788);
xnor U8267 (N_8267,N_4605,N_6043);
nand U8268 (N_8268,N_5265,N_4820);
nand U8269 (N_8269,N_5227,N_4865);
nor U8270 (N_8270,N_3627,N_5926);
and U8271 (N_8271,N_4787,N_5303);
or U8272 (N_8272,N_6223,N_5802);
nor U8273 (N_8273,N_3845,N_5525);
nor U8274 (N_8274,N_6119,N_3213);
or U8275 (N_8275,N_3871,N_4942);
nand U8276 (N_8276,N_3867,N_5139);
nand U8277 (N_8277,N_4513,N_3264);
xor U8278 (N_8278,N_5637,N_5499);
xnor U8279 (N_8279,N_5987,N_5043);
nand U8280 (N_8280,N_6174,N_4097);
and U8281 (N_8281,N_4033,N_5348);
nand U8282 (N_8282,N_5606,N_4095);
xnor U8283 (N_8283,N_4316,N_3969);
and U8284 (N_8284,N_4344,N_4769);
nor U8285 (N_8285,N_3494,N_5111);
nand U8286 (N_8286,N_4731,N_6055);
nor U8287 (N_8287,N_6110,N_6204);
nand U8288 (N_8288,N_5472,N_3902);
nand U8289 (N_8289,N_5193,N_5781);
nand U8290 (N_8290,N_6080,N_5418);
or U8291 (N_8291,N_4090,N_4804);
xnor U8292 (N_8292,N_4313,N_6229);
and U8293 (N_8293,N_5128,N_3576);
nand U8294 (N_8294,N_4612,N_5368);
nor U8295 (N_8295,N_3348,N_5411);
xor U8296 (N_8296,N_4731,N_5637);
or U8297 (N_8297,N_3927,N_6033);
xnor U8298 (N_8298,N_6047,N_6125);
and U8299 (N_8299,N_5577,N_3831);
nor U8300 (N_8300,N_6219,N_5590);
nand U8301 (N_8301,N_3375,N_5460);
or U8302 (N_8302,N_3780,N_5318);
and U8303 (N_8303,N_6163,N_5213);
xor U8304 (N_8304,N_5224,N_5137);
nand U8305 (N_8305,N_5244,N_3152);
nor U8306 (N_8306,N_3332,N_3966);
nor U8307 (N_8307,N_4907,N_3515);
or U8308 (N_8308,N_3525,N_5701);
nor U8309 (N_8309,N_4228,N_3766);
xor U8310 (N_8310,N_4916,N_4968);
nor U8311 (N_8311,N_3158,N_6208);
and U8312 (N_8312,N_5132,N_4510);
nand U8313 (N_8313,N_5416,N_4758);
nand U8314 (N_8314,N_5103,N_3898);
and U8315 (N_8315,N_3538,N_4219);
and U8316 (N_8316,N_3666,N_3702);
nand U8317 (N_8317,N_5194,N_4232);
and U8318 (N_8318,N_3829,N_3566);
nand U8319 (N_8319,N_4435,N_5321);
xnor U8320 (N_8320,N_6181,N_3616);
xnor U8321 (N_8321,N_5137,N_5954);
xor U8322 (N_8322,N_3814,N_4338);
nor U8323 (N_8323,N_6180,N_3647);
nand U8324 (N_8324,N_3889,N_3547);
or U8325 (N_8325,N_5882,N_5702);
nor U8326 (N_8326,N_3884,N_5148);
nor U8327 (N_8327,N_3167,N_3555);
nor U8328 (N_8328,N_4608,N_4974);
nor U8329 (N_8329,N_5684,N_5691);
nand U8330 (N_8330,N_5586,N_3790);
xnor U8331 (N_8331,N_5353,N_5433);
nor U8332 (N_8332,N_3984,N_4500);
nand U8333 (N_8333,N_5487,N_4544);
and U8334 (N_8334,N_4369,N_4660);
xnor U8335 (N_8335,N_3896,N_3934);
or U8336 (N_8336,N_3575,N_4616);
and U8337 (N_8337,N_4428,N_3225);
nor U8338 (N_8338,N_3508,N_3286);
or U8339 (N_8339,N_4588,N_3250);
and U8340 (N_8340,N_6030,N_3308);
and U8341 (N_8341,N_4873,N_5978);
nor U8342 (N_8342,N_3946,N_3475);
or U8343 (N_8343,N_3700,N_4501);
nand U8344 (N_8344,N_3918,N_5848);
nand U8345 (N_8345,N_3912,N_4815);
nor U8346 (N_8346,N_4643,N_5235);
or U8347 (N_8347,N_5692,N_3917);
xor U8348 (N_8348,N_4868,N_6006);
nor U8349 (N_8349,N_4600,N_3653);
nor U8350 (N_8350,N_3591,N_3946);
nand U8351 (N_8351,N_3650,N_3896);
or U8352 (N_8352,N_3133,N_3782);
or U8353 (N_8353,N_5697,N_5066);
nand U8354 (N_8354,N_6091,N_3553);
nand U8355 (N_8355,N_5486,N_5224);
xnor U8356 (N_8356,N_3129,N_3706);
and U8357 (N_8357,N_5680,N_4691);
or U8358 (N_8358,N_4959,N_5253);
and U8359 (N_8359,N_3933,N_3920);
nand U8360 (N_8360,N_5020,N_3731);
or U8361 (N_8361,N_4403,N_3513);
and U8362 (N_8362,N_5924,N_3335);
nor U8363 (N_8363,N_6122,N_5958);
and U8364 (N_8364,N_6215,N_6232);
nand U8365 (N_8365,N_5435,N_3215);
nand U8366 (N_8366,N_4250,N_4499);
nor U8367 (N_8367,N_5370,N_4133);
and U8368 (N_8368,N_3158,N_3922);
nor U8369 (N_8369,N_3594,N_3189);
nor U8370 (N_8370,N_5371,N_3231);
or U8371 (N_8371,N_3239,N_3741);
nand U8372 (N_8372,N_5895,N_5640);
or U8373 (N_8373,N_4368,N_5704);
or U8374 (N_8374,N_6159,N_6201);
xor U8375 (N_8375,N_6107,N_6091);
nor U8376 (N_8376,N_5464,N_4430);
or U8377 (N_8377,N_5681,N_5956);
or U8378 (N_8378,N_5829,N_3950);
and U8379 (N_8379,N_5825,N_5947);
xnor U8380 (N_8380,N_5020,N_5894);
or U8381 (N_8381,N_5601,N_3771);
and U8382 (N_8382,N_4602,N_5321);
or U8383 (N_8383,N_5533,N_5716);
or U8384 (N_8384,N_4018,N_5571);
nor U8385 (N_8385,N_5428,N_5919);
or U8386 (N_8386,N_4300,N_4097);
xnor U8387 (N_8387,N_3643,N_4207);
nor U8388 (N_8388,N_6120,N_3440);
nor U8389 (N_8389,N_4695,N_4118);
nor U8390 (N_8390,N_3542,N_3200);
or U8391 (N_8391,N_5865,N_5336);
nor U8392 (N_8392,N_3548,N_5424);
and U8393 (N_8393,N_3663,N_5273);
or U8394 (N_8394,N_4795,N_5196);
or U8395 (N_8395,N_3337,N_6177);
nor U8396 (N_8396,N_4265,N_5859);
or U8397 (N_8397,N_3692,N_4444);
or U8398 (N_8398,N_4738,N_4488);
nor U8399 (N_8399,N_3739,N_3895);
or U8400 (N_8400,N_5355,N_4267);
or U8401 (N_8401,N_4600,N_4295);
nor U8402 (N_8402,N_5581,N_5876);
xnor U8403 (N_8403,N_5294,N_3334);
xor U8404 (N_8404,N_4358,N_3449);
and U8405 (N_8405,N_3812,N_3891);
or U8406 (N_8406,N_5827,N_3232);
nor U8407 (N_8407,N_3693,N_6244);
nor U8408 (N_8408,N_3266,N_4308);
nor U8409 (N_8409,N_6069,N_4924);
nor U8410 (N_8410,N_3218,N_3762);
nand U8411 (N_8411,N_4562,N_3228);
and U8412 (N_8412,N_5879,N_4972);
xor U8413 (N_8413,N_3177,N_4056);
nand U8414 (N_8414,N_3326,N_5497);
and U8415 (N_8415,N_5983,N_3759);
and U8416 (N_8416,N_4937,N_4671);
or U8417 (N_8417,N_4734,N_5022);
nand U8418 (N_8418,N_5507,N_4879);
xnor U8419 (N_8419,N_4735,N_4374);
or U8420 (N_8420,N_4346,N_4323);
and U8421 (N_8421,N_3647,N_4902);
nor U8422 (N_8422,N_3515,N_5924);
or U8423 (N_8423,N_4986,N_5070);
xnor U8424 (N_8424,N_5094,N_4651);
nor U8425 (N_8425,N_5573,N_5721);
nand U8426 (N_8426,N_5216,N_6079);
nand U8427 (N_8427,N_3780,N_3596);
or U8428 (N_8428,N_5869,N_6128);
nor U8429 (N_8429,N_5170,N_5275);
and U8430 (N_8430,N_4415,N_4795);
nor U8431 (N_8431,N_5316,N_3952);
and U8432 (N_8432,N_5529,N_4783);
nand U8433 (N_8433,N_4104,N_3939);
nor U8434 (N_8434,N_6065,N_3992);
or U8435 (N_8435,N_4892,N_6012);
and U8436 (N_8436,N_3981,N_5681);
xnor U8437 (N_8437,N_4652,N_3940);
and U8438 (N_8438,N_6127,N_4724);
or U8439 (N_8439,N_4490,N_3177);
xnor U8440 (N_8440,N_5654,N_5392);
or U8441 (N_8441,N_6239,N_5154);
or U8442 (N_8442,N_3471,N_3775);
nor U8443 (N_8443,N_4016,N_3425);
and U8444 (N_8444,N_3388,N_3250);
nor U8445 (N_8445,N_5212,N_3498);
and U8446 (N_8446,N_3747,N_5355);
and U8447 (N_8447,N_3627,N_5695);
or U8448 (N_8448,N_5897,N_4258);
nand U8449 (N_8449,N_5481,N_3859);
nand U8450 (N_8450,N_3389,N_5380);
nand U8451 (N_8451,N_5533,N_3253);
xor U8452 (N_8452,N_4033,N_5073);
nand U8453 (N_8453,N_3385,N_5744);
nor U8454 (N_8454,N_4059,N_3308);
and U8455 (N_8455,N_4569,N_5604);
xor U8456 (N_8456,N_4242,N_4365);
nand U8457 (N_8457,N_5212,N_5201);
xor U8458 (N_8458,N_5646,N_5406);
or U8459 (N_8459,N_3536,N_3714);
nor U8460 (N_8460,N_5629,N_3747);
nor U8461 (N_8461,N_3949,N_4156);
nor U8462 (N_8462,N_5716,N_4471);
xor U8463 (N_8463,N_4749,N_5913);
and U8464 (N_8464,N_4306,N_3967);
nand U8465 (N_8465,N_4924,N_4478);
xor U8466 (N_8466,N_6109,N_5667);
nand U8467 (N_8467,N_3904,N_3262);
or U8468 (N_8468,N_3840,N_4610);
xor U8469 (N_8469,N_4187,N_3916);
nor U8470 (N_8470,N_4531,N_4896);
nor U8471 (N_8471,N_4077,N_6199);
nand U8472 (N_8472,N_3866,N_5228);
nor U8473 (N_8473,N_3244,N_5375);
and U8474 (N_8474,N_4756,N_3844);
or U8475 (N_8475,N_5080,N_5201);
and U8476 (N_8476,N_6057,N_4457);
nand U8477 (N_8477,N_5427,N_3474);
nand U8478 (N_8478,N_4515,N_5529);
and U8479 (N_8479,N_3390,N_3649);
xor U8480 (N_8480,N_4236,N_3179);
nor U8481 (N_8481,N_4133,N_3308);
and U8482 (N_8482,N_3674,N_3514);
and U8483 (N_8483,N_4586,N_4865);
xnor U8484 (N_8484,N_3165,N_3676);
and U8485 (N_8485,N_4696,N_3970);
and U8486 (N_8486,N_5318,N_5012);
nand U8487 (N_8487,N_4498,N_4330);
xor U8488 (N_8488,N_3154,N_5690);
nand U8489 (N_8489,N_5991,N_3450);
or U8490 (N_8490,N_5478,N_5506);
xor U8491 (N_8491,N_4601,N_5173);
nor U8492 (N_8492,N_4199,N_3384);
or U8493 (N_8493,N_4771,N_5443);
or U8494 (N_8494,N_4040,N_4077);
nor U8495 (N_8495,N_5496,N_6052);
xnor U8496 (N_8496,N_3809,N_5516);
nand U8497 (N_8497,N_5721,N_3456);
nand U8498 (N_8498,N_4248,N_3147);
and U8499 (N_8499,N_3988,N_3768);
nor U8500 (N_8500,N_3350,N_6143);
and U8501 (N_8501,N_3152,N_3125);
and U8502 (N_8502,N_5553,N_4512);
and U8503 (N_8503,N_6019,N_5309);
or U8504 (N_8504,N_4576,N_5895);
and U8505 (N_8505,N_3582,N_5791);
nand U8506 (N_8506,N_4665,N_3308);
nand U8507 (N_8507,N_3771,N_5674);
nor U8508 (N_8508,N_4038,N_4371);
nand U8509 (N_8509,N_3463,N_4835);
and U8510 (N_8510,N_4144,N_4784);
or U8511 (N_8511,N_4077,N_5473);
or U8512 (N_8512,N_5283,N_3558);
or U8513 (N_8513,N_5790,N_5576);
and U8514 (N_8514,N_4992,N_5167);
or U8515 (N_8515,N_3286,N_5194);
nand U8516 (N_8516,N_5730,N_4176);
nor U8517 (N_8517,N_4411,N_3189);
nand U8518 (N_8518,N_3438,N_3439);
nand U8519 (N_8519,N_3616,N_6168);
and U8520 (N_8520,N_3449,N_3841);
or U8521 (N_8521,N_4147,N_4837);
or U8522 (N_8522,N_4119,N_5593);
nor U8523 (N_8523,N_5867,N_3440);
nand U8524 (N_8524,N_4913,N_4644);
nand U8525 (N_8525,N_5334,N_4792);
or U8526 (N_8526,N_3475,N_6018);
and U8527 (N_8527,N_5675,N_4366);
or U8528 (N_8528,N_6079,N_4838);
and U8529 (N_8529,N_5778,N_5032);
nand U8530 (N_8530,N_5695,N_5585);
nor U8531 (N_8531,N_5291,N_4414);
nor U8532 (N_8532,N_5331,N_3784);
nor U8533 (N_8533,N_5127,N_4832);
or U8534 (N_8534,N_4855,N_4489);
nor U8535 (N_8535,N_4013,N_4607);
nand U8536 (N_8536,N_3500,N_3237);
nor U8537 (N_8537,N_3135,N_5948);
or U8538 (N_8538,N_5220,N_4530);
and U8539 (N_8539,N_6134,N_4457);
nor U8540 (N_8540,N_5692,N_4390);
or U8541 (N_8541,N_3184,N_6034);
nand U8542 (N_8542,N_3323,N_3926);
nand U8543 (N_8543,N_4917,N_5924);
and U8544 (N_8544,N_6238,N_5399);
nor U8545 (N_8545,N_3232,N_3152);
and U8546 (N_8546,N_3860,N_3283);
nand U8547 (N_8547,N_5022,N_5629);
and U8548 (N_8548,N_5150,N_5086);
xor U8549 (N_8549,N_5988,N_4812);
nor U8550 (N_8550,N_3834,N_3608);
and U8551 (N_8551,N_5469,N_4765);
xnor U8552 (N_8552,N_5647,N_4388);
and U8553 (N_8553,N_5368,N_5105);
or U8554 (N_8554,N_5508,N_4721);
and U8555 (N_8555,N_5317,N_5907);
nand U8556 (N_8556,N_5946,N_6074);
nor U8557 (N_8557,N_4015,N_5928);
or U8558 (N_8558,N_3609,N_4634);
nand U8559 (N_8559,N_5736,N_5109);
or U8560 (N_8560,N_3315,N_4195);
or U8561 (N_8561,N_5323,N_3827);
nand U8562 (N_8562,N_4801,N_3266);
or U8563 (N_8563,N_5684,N_5666);
nor U8564 (N_8564,N_5663,N_5856);
and U8565 (N_8565,N_5380,N_3182);
nor U8566 (N_8566,N_4509,N_6159);
nand U8567 (N_8567,N_4148,N_5364);
xor U8568 (N_8568,N_3923,N_4308);
nand U8569 (N_8569,N_4175,N_3913);
nand U8570 (N_8570,N_4198,N_5019);
and U8571 (N_8571,N_5155,N_5265);
nor U8572 (N_8572,N_5891,N_3876);
nand U8573 (N_8573,N_4846,N_5410);
nand U8574 (N_8574,N_6059,N_3795);
nor U8575 (N_8575,N_4479,N_4246);
and U8576 (N_8576,N_5874,N_6180);
nand U8577 (N_8577,N_3631,N_4104);
nor U8578 (N_8578,N_4320,N_5166);
or U8579 (N_8579,N_3438,N_4026);
or U8580 (N_8580,N_4306,N_3268);
nand U8581 (N_8581,N_5128,N_4253);
xor U8582 (N_8582,N_3994,N_4479);
or U8583 (N_8583,N_3663,N_5390);
nor U8584 (N_8584,N_4078,N_4418);
nand U8585 (N_8585,N_3445,N_4486);
and U8586 (N_8586,N_4192,N_3809);
nand U8587 (N_8587,N_5793,N_4694);
or U8588 (N_8588,N_5894,N_5437);
nor U8589 (N_8589,N_4441,N_5290);
nand U8590 (N_8590,N_4242,N_4376);
nor U8591 (N_8591,N_5752,N_4370);
nor U8592 (N_8592,N_5846,N_4993);
nor U8593 (N_8593,N_3565,N_4516);
or U8594 (N_8594,N_4699,N_4261);
or U8595 (N_8595,N_4280,N_3128);
nand U8596 (N_8596,N_3501,N_4505);
or U8597 (N_8597,N_3834,N_4040);
nor U8598 (N_8598,N_3457,N_5943);
xnor U8599 (N_8599,N_5071,N_3718);
nor U8600 (N_8600,N_3199,N_3685);
or U8601 (N_8601,N_5264,N_5258);
and U8602 (N_8602,N_5322,N_3356);
nor U8603 (N_8603,N_3436,N_5046);
and U8604 (N_8604,N_5679,N_6225);
nand U8605 (N_8605,N_3171,N_3401);
xor U8606 (N_8606,N_6147,N_6185);
nand U8607 (N_8607,N_3578,N_4581);
nor U8608 (N_8608,N_5322,N_4376);
nor U8609 (N_8609,N_5638,N_6055);
nor U8610 (N_8610,N_5593,N_3168);
nor U8611 (N_8611,N_3870,N_3716);
or U8612 (N_8612,N_6235,N_5435);
nand U8613 (N_8613,N_3521,N_3431);
and U8614 (N_8614,N_5833,N_4570);
nor U8615 (N_8615,N_4865,N_3286);
or U8616 (N_8616,N_5974,N_3696);
nor U8617 (N_8617,N_3324,N_5240);
nand U8618 (N_8618,N_5318,N_5409);
and U8619 (N_8619,N_3479,N_6006);
nor U8620 (N_8620,N_4517,N_4785);
or U8621 (N_8621,N_5648,N_5273);
or U8622 (N_8622,N_3356,N_5885);
nor U8623 (N_8623,N_3737,N_4311);
nand U8624 (N_8624,N_3362,N_4445);
nor U8625 (N_8625,N_5124,N_3885);
nand U8626 (N_8626,N_4381,N_3744);
xnor U8627 (N_8627,N_5706,N_3735);
or U8628 (N_8628,N_4712,N_5534);
nand U8629 (N_8629,N_5216,N_4256);
nand U8630 (N_8630,N_4317,N_3297);
nor U8631 (N_8631,N_5076,N_5310);
and U8632 (N_8632,N_5160,N_4988);
nand U8633 (N_8633,N_4769,N_4257);
nand U8634 (N_8634,N_6025,N_5058);
or U8635 (N_8635,N_6001,N_4930);
or U8636 (N_8636,N_5043,N_5819);
nor U8637 (N_8637,N_4504,N_3474);
xor U8638 (N_8638,N_4056,N_5176);
and U8639 (N_8639,N_4016,N_5594);
and U8640 (N_8640,N_4808,N_5258);
nand U8641 (N_8641,N_4589,N_3610);
or U8642 (N_8642,N_5630,N_5666);
and U8643 (N_8643,N_4394,N_4243);
nor U8644 (N_8644,N_3312,N_4558);
and U8645 (N_8645,N_3295,N_4998);
and U8646 (N_8646,N_4848,N_5288);
nor U8647 (N_8647,N_3313,N_4990);
xor U8648 (N_8648,N_5378,N_3678);
nand U8649 (N_8649,N_5311,N_4097);
and U8650 (N_8650,N_4045,N_3658);
and U8651 (N_8651,N_3823,N_4187);
nor U8652 (N_8652,N_5661,N_3424);
nand U8653 (N_8653,N_4487,N_5664);
and U8654 (N_8654,N_5083,N_4031);
nand U8655 (N_8655,N_3200,N_3487);
xor U8656 (N_8656,N_5672,N_4729);
nand U8657 (N_8657,N_5415,N_5587);
nand U8658 (N_8658,N_3817,N_3390);
and U8659 (N_8659,N_3329,N_5647);
nand U8660 (N_8660,N_3496,N_4481);
or U8661 (N_8661,N_5534,N_4708);
or U8662 (N_8662,N_4231,N_3220);
nand U8663 (N_8663,N_4009,N_6210);
xnor U8664 (N_8664,N_5750,N_3406);
nand U8665 (N_8665,N_5983,N_5086);
nor U8666 (N_8666,N_4636,N_5501);
or U8667 (N_8667,N_4464,N_6205);
nor U8668 (N_8668,N_3376,N_5768);
nand U8669 (N_8669,N_3631,N_3246);
xnor U8670 (N_8670,N_4679,N_4733);
or U8671 (N_8671,N_3174,N_3185);
nand U8672 (N_8672,N_5169,N_5624);
or U8673 (N_8673,N_3613,N_4328);
nor U8674 (N_8674,N_3624,N_5558);
nand U8675 (N_8675,N_3990,N_6237);
or U8676 (N_8676,N_3630,N_5884);
nand U8677 (N_8677,N_3526,N_5105);
nor U8678 (N_8678,N_5369,N_6215);
nor U8679 (N_8679,N_5458,N_3319);
and U8680 (N_8680,N_3766,N_3337);
nor U8681 (N_8681,N_4699,N_4600);
or U8682 (N_8682,N_3530,N_6172);
and U8683 (N_8683,N_4086,N_4577);
nand U8684 (N_8684,N_3574,N_4981);
nor U8685 (N_8685,N_3980,N_4937);
xnor U8686 (N_8686,N_4066,N_5773);
xor U8687 (N_8687,N_3839,N_4192);
xnor U8688 (N_8688,N_4380,N_5619);
nor U8689 (N_8689,N_3336,N_5309);
or U8690 (N_8690,N_4693,N_5591);
nand U8691 (N_8691,N_3135,N_4472);
and U8692 (N_8692,N_3899,N_4893);
and U8693 (N_8693,N_5300,N_4080);
or U8694 (N_8694,N_4517,N_5839);
nor U8695 (N_8695,N_5474,N_4675);
or U8696 (N_8696,N_3560,N_5546);
or U8697 (N_8697,N_6025,N_5597);
nand U8698 (N_8698,N_4165,N_5928);
and U8699 (N_8699,N_5509,N_3891);
nand U8700 (N_8700,N_5888,N_4858);
and U8701 (N_8701,N_5250,N_4553);
xnor U8702 (N_8702,N_4230,N_5424);
and U8703 (N_8703,N_6138,N_5868);
or U8704 (N_8704,N_3907,N_3221);
and U8705 (N_8705,N_3774,N_3446);
xor U8706 (N_8706,N_5809,N_3736);
and U8707 (N_8707,N_3413,N_5464);
nor U8708 (N_8708,N_6063,N_3381);
nor U8709 (N_8709,N_3231,N_5767);
or U8710 (N_8710,N_3692,N_3388);
or U8711 (N_8711,N_5240,N_3233);
nor U8712 (N_8712,N_4730,N_3547);
nor U8713 (N_8713,N_3440,N_5938);
or U8714 (N_8714,N_3804,N_3648);
nand U8715 (N_8715,N_4686,N_6229);
or U8716 (N_8716,N_4912,N_5754);
nor U8717 (N_8717,N_4811,N_4832);
nand U8718 (N_8718,N_4579,N_6226);
and U8719 (N_8719,N_5162,N_3358);
nor U8720 (N_8720,N_5470,N_5156);
or U8721 (N_8721,N_6173,N_6216);
and U8722 (N_8722,N_5734,N_5419);
and U8723 (N_8723,N_3144,N_4740);
xnor U8724 (N_8724,N_4997,N_3737);
nor U8725 (N_8725,N_4828,N_5504);
or U8726 (N_8726,N_4104,N_6129);
nand U8727 (N_8727,N_3939,N_3647);
or U8728 (N_8728,N_4522,N_3603);
xnor U8729 (N_8729,N_3617,N_3956);
and U8730 (N_8730,N_5862,N_4888);
and U8731 (N_8731,N_3368,N_3164);
and U8732 (N_8732,N_5839,N_3145);
and U8733 (N_8733,N_4001,N_5403);
xor U8734 (N_8734,N_6215,N_4556);
nor U8735 (N_8735,N_3566,N_4734);
and U8736 (N_8736,N_3885,N_5166);
xor U8737 (N_8737,N_4245,N_5686);
xnor U8738 (N_8738,N_5765,N_5713);
nand U8739 (N_8739,N_3959,N_5072);
nor U8740 (N_8740,N_6086,N_4598);
and U8741 (N_8741,N_5760,N_6039);
nor U8742 (N_8742,N_3749,N_4285);
or U8743 (N_8743,N_3261,N_6148);
or U8744 (N_8744,N_3950,N_3349);
or U8745 (N_8745,N_5964,N_5180);
and U8746 (N_8746,N_3703,N_4884);
or U8747 (N_8747,N_3498,N_4902);
nor U8748 (N_8748,N_3500,N_3972);
and U8749 (N_8749,N_4370,N_3931);
and U8750 (N_8750,N_3578,N_3733);
nor U8751 (N_8751,N_4469,N_5082);
nand U8752 (N_8752,N_4069,N_4936);
or U8753 (N_8753,N_3366,N_3679);
and U8754 (N_8754,N_4566,N_5227);
or U8755 (N_8755,N_5481,N_4841);
or U8756 (N_8756,N_5815,N_3330);
nor U8757 (N_8757,N_3298,N_6068);
nor U8758 (N_8758,N_5384,N_6009);
nor U8759 (N_8759,N_3386,N_3261);
or U8760 (N_8760,N_3665,N_4999);
or U8761 (N_8761,N_6118,N_3629);
nor U8762 (N_8762,N_6233,N_3688);
xor U8763 (N_8763,N_5705,N_5215);
or U8764 (N_8764,N_3928,N_5890);
or U8765 (N_8765,N_3334,N_3605);
or U8766 (N_8766,N_4315,N_4037);
or U8767 (N_8767,N_3301,N_4561);
and U8768 (N_8768,N_5185,N_4221);
or U8769 (N_8769,N_3524,N_3499);
xnor U8770 (N_8770,N_3831,N_4913);
nor U8771 (N_8771,N_4490,N_4270);
xnor U8772 (N_8772,N_5691,N_6051);
or U8773 (N_8773,N_3685,N_4141);
nor U8774 (N_8774,N_5176,N_3785);
or U8775 (N_8775,N_5037,N_5785);
nand U8776 (N_8776,N_5483,N_4520);
nor U8777 (N_8777,N_5538,N_4380);
nor U8778 (N_8778,N_4585,N_4006);
and U8779 (N_8779,N_5183,N_6002);
and U8780 (N_8780,N_5069,N_3853);
nand U8781 (N_8781,N_5702,N_3964);
nand U8782 (N_8782,N_3444,N_5269);
xnor U8783 (N_8783,N_4368,N_5400);
nand U8784 (N_8784,N_6161,N_5899);
or U8785 (N_8785,N_5759,N_5184);
nor U8786 (N_8786,N_4219,N_3393);
xnor U8787 (N_8787,N_5119,N_5826);
and U8788 (N_8788,N_4441,N_3885);
and U8789 (N_8789,N_3269,N_3927);
or U8790 (N_8790,N_3702,N_6010);
nand U8791 (N_8791,N_4861,N_3741);
nand U8792 (N_8792,N_3125,N_3339);
and U8793 (N_8793,N_5017,N_6029);
nor U8794 (N_8794,N_4689,N_3583);
nor U8795 (N_8795,N_5738,N_6109);
and U8796 (N_8796,N_5422,N_5486);
nand U8797 (N_8797,N_5281,N_3452);
and U8798 (N_8798,N_6088,N_5087);
and U8799 (N_8799,N_6156,N_5533);
nor U8800 (N_8800,N_4484,N_4678);
nand U8801 (N_8801,N_3191,N_6063);
nand U8802 (N_8802,N_4610,N_5313);
or U8803 (N_8803,N_3159,N_5835);
nand U8804 (N_8804,N_4847,N_3286);
or U8805 (N_8805,N_5270,N_5581);
nor U8806 (N_8806,N_6202,N_4417);
nand U8807 (N_8807,N_4411,N_5700);
or U8808 (N_8808,N_3481,N_4826);
nor U8809 (N_8809,N_4074,N_3723);
nand U8810 (N_8810,N_3598,N_5567);
or U8811 (N_8811,N_5289,N_6183);
or U8812 (N_8812,N_3129,N_4905);
nand U8813 (N_8813,N_3310,N_4126);
nand U8814 (N_8814,N_5495,N_5644);
or U8815 (N_8815,N_3214,N_4186);
nand U8816 (N_8816,N_3673,N_4588);
nand U8817 (N_8817,N_3806,N_3783);
nor U8818 (N_8818,N_3644,N_6218);
nand U8819 (N_8819,N_3252,N_5053);
and U8820 (N_8820,N_3990,N_5562);
or U8821 (N_8821,N_4269,N_3916);
or U8822 (N_8822,N_4778,N_3662);
or U8823 (N_8823,N_5026,N_4546);
and U8824 (N_8824,N_4527,N_5559);
nand U8825 (N_8825,N_5134,N_5825);
nand U8826 (N_8826,N_5128,N_5087);
nor U8827 (N_8827,N_3343,N_4787);
and U8828 (N_8828,N_4075,N_4290);
nand U8829 (N_8829,N_3217,N_5777);
or U8830 (N_8830,N_4330,N_3559);
nand U8831 (N_8831,N_3639,N_3741);
xor U8832 (N_8832,N_5603,N_3142);
nor U8833 (N_8833,N_4771,N_4730);
xnor U8834 (N_8834,N_3855,N_5377);
and U8835 (N_8835,N_5331,N_4887);
and U8836 (N_8836,N_3479,N_3709);
nand U8837 (N_8837,N_5263,N_4437);
or U8838 (N_8838,N_4693,N_5581);
and U8839 (N_8839,N_5057,N_4700);
xor U8840 (N_8840,N_4880,N_4887);
nor U8841 (N_8841,N_5087,N_3878);
nand U8842 (N_8842,N_5007,N_4334);
and U8843 (N_8843,N_3581,N_5679);
nor U8844 (N_8844,N_3449,N_5268);
and U8845 (N_8845,N_5815,N_5482);
or U8846 (N_8846,N_4279,N_5322);
nor U8847 (N_8847,N_4709,N_4081);
nor U8848 (N_8848,N_6208,N_5274);
nor U8849 (N_8849,N_3307,N_5173);
or U8850 (N_8850,N_3665,N_4161);
and U8851 (N_8851,N_6048,N_4654);
and U8852 (N_8852,N_5197,N_3514);
or U8853 (N_8853,N_3971,N_3283);
and U8854 (N_8854,N_5252,N_5820);
or U8855 (N_8855,N_5374,N_3661);
and U8856 (N_8856,N_4233,N_4087);
xor U8857 (N_8857,N_4505,N_5325);
nand U8858 (N_8858,N_5390,N_3622);
nand U8859 (N_8859,N_4045,N_5245);
or U8860 (N_8860,N_5900,N_5333);
and U8861 (N_8861,N_4514,N_4468);
nand U8862 (N_8862,N_4606,N_4030);
nor U8863 (N_8863,N_4470,N_4152);
or U8864 (N_8864,N_4155,N_3959);
and U8865 (N_8865,N_3954,N_6182);
and U8866 (N_8866,N_4685,N_6075);
nor U8867 (N_8867,N_5472,N_3935);
nor U8868 (N_8868,N_4853,N_3990);
and U8869 (N_8869,N_4538,N_5326);
or U8870 (N_8870,N_5558,N_5373);
xor U8871 (N_8871,N_4684,N_5098);
nand U8872 (N_8872,N_5666,N_3966);
or U8873 (N_8873,N_5335,N_4019);
or U8874 (N_8874,N_5101,N_4387);
or U8875 (N_8875,N_5153,N_4985);
or U8876 (N_8876,N_5537,N_5070);
and U8877 (N_8877,N_5394,N_5680);
nand U8878 (N_8878,N_3282,N_4135);
or U8879 (N_8879,N_4435,N_3294);
nand U8880 (N_8880,N_3843,N_6199);
nand U8881 (N_8881,N_5357,N_6025);
nand U8882 (N_8882,N_5101,N_4367);
nor U8883 (N_8883,N_3488,N_4085);
nand U8884 (N_8884,N_4025,N_6112);
nor U8885 (N_8885,N_5339,N_3587);
nand U8886 (N_8886,N_4631,N_3364);
or U8887 (N_8887,N_4729,N_3507);
nand U8888 (N_8888,N_3322,N_5872);
nand U8889 (N_8889,N_3793,N_3721);
xor U8890 (N_8890,N_3542,N_3533);
xor U8891 (N_8891,N_4099,N_4807);
or U8892 (N_8892,N_3404,N_4004);
or U8893 (N_8893,N_4892,N_3405);
xor U8894 (N_8894,N_4111,N_6144);
nand U8895 (N_8895,N_3876,N_6180);
nand U8896 (N_8896,N_5797,N_3484);
or U8897 (N_8897,N_3826,N_4424);
nor U8898 (N_8898,N_4745,N_5372);
nand U8899 (N_8899,N_5516,N_3423);
or U8900 (N_8900,N_4083,N_5803);
and U8901 (N_8901,N_5161,N_3738);
nor U8902 (N_8902,N_5823,N_6116);
or U8903 (N_8903,N_4819,N_4140);
nand U8904 (N_8904,N_5377,N_4848);
nand U8905 (N_8905,N_5798,N_4695);
nand U8906 (N_8906,N_5109,N_3264);
or U8907 (N_8907,N_3510,N_5168);
or U8908 (N_8908,N_4240,N_5892);
or U8909 (N_8909,N_3691,N_5612);
and U8910 (N_8910,N_5115,N_5793);
or U8911 (N_8911,N_3797,N_3480);
xor U8912 (N_8912,N_5530,N_5008);
nand U8913 (N_8913,N_3341,N_5816);
nand U8914 (N_8914,N_5925,N_5611);
and U8915 (N_8915,N_3668,N_3416);
or U8916 (N_8916,N_3646,N_3212);
nor U8917 (N_8917,N_5022,N_4062);
or U8918 (N_8918,N_4783,N_4349);
and U8919 (N_8919,N_4886,N_6092);
nand U8920 (N_8920,N_5760,N_3652);
nand U8921 (N_8921,N_5970,N_4946);
or U8922 (N_8922,N_3481,N_5736);
nand U8923 (N_8923,N_3430,N_4222);
and U8924 (N_8924,N_4226,N_5686);
and U8925 (N_8925,N_3422,N_5910);
nand U8926 (N_8926,N_5774,N_4996);
or U8927 (N_8927,N_3996,N_3603);
and U8928 (N_8928,N_3425,N_6013);
xor U8929 (N_8929,N_4198,N_5555);
xnor U8930 (N_8930,N_4737,N_5181);
or U8931 (N_8931,N_4302,N_5972);
and U8932 (N_8932,N_3815,N_3133);
nor U8933 (N_8933,N_3709,N_5336);
and U8934 (N_8934,N_5075,N_3349);
nand U8935 (N_8935,N_4804,N_5267);
nand U8936 (N_8936,N_5648,N_4803);
nand U8937 (N_8937,N_4583,N_4295);
nor U8938 (N_8938,N_5502,N_4057);
nor U8939 (N_8939,N_5677,N_4863);
nand U8940 (N_8940,N_5377,N_3533);
nand U8941 (N_8941,N_4172,N_5941);
nor U8942 (N_8942,N_4889,N_3287);
or U8943 (N_8943,N_5933,N_4048);
and U8944 (N_8944,N_5771,N_4123);
nor U8945 (N_8945,N_6032,N_6199);
or U8946 (N_8946,N_4136,N_4882);
xnor U8947 (N_8947,N_4075,N_6152);
xnor U8948 (N_8948,N_4849,N_3154);
nand U8949 (N_8949,N_6222,N_5871);
xnor U8950 (N_8950,N_4243,N_5887);
xnor U8951 (N_8951,N_5599,N_5075);
nor U8952 (N_8952,N_5919,N_3305);
nor U8953 (N_8953,N_4049,N_3354);
xnor U8954 (N_8954,N_3281,N_4295);
and U8955 (N_8955,N_3702,N_5718);
nor U8956 (N_8956,N_5046,N_3772);
nor U8957 (N_8957,N_5568,N_6163);
or U8958 (N_8958,N_5164,N_4400);
nor U8959 (N_8959,N_5345,N_5129);
nor U8960 (N_8960,N_4394,N_5097);
or U8961 (N_8961,N_5245,N_6055);
and U8962 (N_8962,N_6001,N_4106);
and U8963 (N_8963,N_3796,N_5957);
or U8964 (N_8964,N_3237,N_4095);
or U8965 (N_8965,N_5629,N_5642);
and U8966 (N_8966,N_4796,N_3510);
nand U8967 (N_8967,N_6061,N_5016);
nor U8968 (N_8968,N_6037,N_3766);
nand U8969 (N_8969,N_4688,N_5308);
nand U8970 (N_8970,N_4819,N_5175);
nand U8971 (N_8971,N_5606,N_4274);
and U8972 (N_8972,N_4153,N_5896);
nor U8973 (N_8973,N_5494,N_4835);
and U8974 (N_8974,N_3126,N_5769);
nor U8975 (N_8975,N_3808,N_5025);
xor U8976 (N_8976,N_4215,N_4193);
and U8977 (N_8977,N_5091,N_4595);
nor U8978 (N_8978,N_5596,N_4213);
nor U8979 (N_8979,N_4672,N_5159);
nand U8980 (N_8980,N_3325,N_5677);
and U8981 (N_8981,N_5408,N_3974);
and U8982 (N_8982,N_4139,N_5424);
nor U8983 (N_8983,N_5551,N_5438);
nor U8984 (N_8984,N_5551,N_3826);
and U8985 (N_8985,N_4914,N_5295);
nor U8986 (N_8986,N_6209,N_4603);
or U8987 (N_8987,N_5392,N_5531);
and U8988 (N_8988,N_6151,N_5162);
nor U8989 (N_8989,N_4959,N_3349);
and U8990 (N_8990,N_3859,N_3700);
nor U8991 (N_8991,N_5491,N_5381);
or U8992 (N_8992,N_3218,N_4641);
or U8993 (N_8993,N_3249,N_5194);
nand U8994 (N_8994,N_6018,N_5834);
nor U8995 (N_8995,N_4894,N_5891);
and U8996 (N_8996,N_5445,N_3909);
nor U8997 (N_8997,N_4708,N_5922);
nor U8998 (N_8998,N_3312,N_5620);
and U8999 (N_8999,N_5793,N_4178);
xor U9000 (N_9000,N_4942,N_3506);
nand U9001 (N_9001,N_4454,N_3907);
or U9002 (N_9002,N_5555,N_5925);
xnor U9003 (N_9003,N_3384,N_5676);
nor U9004 (N_9004,N_4874,N_3776);
nand U9005 (N_9005,N_4959,N_3296);
or U9006 (N_9006,N_6005,N_4439);
or U9007 (N_9007,N_6026,N_4960);
nor U9008 (N_9008,N_5929,N_4754);
and U9009 (N_9009,N_5306,N_5834);
nand U9010 (N_9010,N_4971,N_4309);
nor U9011 (N_9011,N_5840,N_3938);
nand U9012 (N_9012,N_4282,N_4026);
xnor U9013 (N_9013,N_4128,N_5852);
nor U9014 (N_9014,N_5219,N_6229);
nor U9015 (N_9015,N_3503,N_4906);
or U9016 (N_9016,N_4415,N_3325);
xor U9017 (N_9017,N_4027,N_5446);
and U9018 (N_9018,N_3131,N_5844);
nor U9019 (N_9019,N_3436,N_6008);
and U9020 (N_9020,N_3248,N_5001);
nand U9021 (N_9021,N_5127,N_5253);
nor U9022 (N_9022,N_5321,N_4883);
or U9023 (N_9023,N_4283,N_3495);
or U9024 (N_9024,N_3265,N_4735);
or U9025 (N_9025,N_4702,N_5714);
or U9026 (N_9026,N_3595,N_4994);
and U9027 (N_9027,N_4678,N_3723);
or U9028 (N_9028,N_4671,N_5202);
or U9029 (N_9029,N_4273,N_4132);
nor U9030 (N_9030,N_5753,N_5999);
or U9031 (N_9031,N_3421,N_3991);
xnor U9032 (N_9032,N_5678,N_3501);
or U9033 (N_9033,N_5331,N_4037);
xor U9034 (N_9034,N_4893,N_5705);
xnor U9035 (N_9035,N_3894,N_5080);
nor U9036 (N_9036,N_5512,N_4655);
nand U9037 (N_9037,N_4877,N_4961);
nand U9038 (N_9038,N_4175,N_4862);
and U9039 (N_9039,N_4888,N_5016);
or U9040 (N_9040,N_4149,N_6027);
or U9041 (N_9041,N_6160,N_5754);
or U9042 (N_9042,N_5700,N_3126);
or U9043 (N_9043,N_5321,N_4150);
nor U9044 (N_9044,N_3598,N_4894);
or U9045 (N_9045,N_3646,N_5109);
or U9046 (N_9046,N_5512,N_5092);
xnor U9047 (N_9047,N_5022,N_4404);
nor U9048 (N_9048,N_3813,N_3169);
or U9049 (N_9049,N_4061,N_4709);
xor U9050 (N_9050,N_5679,N_5620);
or U9051 (N_9051,N_4870,N_5407);
nand U9052 (N_9052,N_5937,N_4955);
xnor U9053 (N_9053,N_5465,N_5521);
and U9054 (N_9054,N_3474,N_5331);
and U9055 (N_9055,N_5888,N_4306);
nor U9056 (N_9056,N_4025,N_4526);
nand U9057 (N_9057,N_4510,N_5178);
and U9058 (N_9058,N_4622,N_5864);
or U9059 (N_9059,N_3178,N_4992);
nand U9060 (N_9060,N_6028,N_4212);
and U9061 (N_9061,N_3583,N_4806);
nand U9062 (N_9062,N_5290,N_3863);
nand U9063 (N_9063,N_5156,N_5738);
and U9064 (N_9064,N_4089,N_6182);
xor U9065 (N_9065,N_5489,N_3667);
and U9066 (N_9066,N_5747,N_4695);
nor U9067 (N_9067,N_3893,N_3777);
nor U9068 (N_9068,N_5611,N_4446);
nand U9069 (N_9069,N_4075,N_5069);
and U9070 (N_9070,N_4874,N_3989);
nand U9071 (N_9071,N_3987,N_3664);
nor U9072 (N_9072,N_3484,N_4051);
or U9073 (N_9073,N_5716,N_5750);
nor U9074 (N_9074,N_3786,N_4017);
and U9075 (N_9075,N_5040,N_4071);
nor U9076 (N_9076,N_5421,N_3550);
or U9077 (N_9077,N_5905,N_5752);
nand U9078 (N_9078,N_3639,N_3373);
or U9079 (N_9079,N_5938,N_4114);
or U9080 (N_9080,N_4453,N_5873);
nor U9081 (N_9081,N_3136,N_3205);
xor U9082 (N_9082,N_5491,N_4461);
and U9083 (N_9083,N_3125,N_5993);
or U9084 (N_9084,N_3614,N_4810);
nand U9085 (N_9085,N_3346,N_4859);
or U9086 (N_9086,N_4150,N_4499);
and U9087 (N_9087,N_4650,N_4557);
nand U9088 (N_9088,N_5270,N_3493);
nand U9089 (N_9089,N_5164,N_4407);
and U9090 (N_9090,N_5333,N_5787);
and U9091 (N_9091,N_4469,N_4264);
nand U9092 (N_9092,N_5424,N_3449);
and U9093 (N_9093,N_3486,N_4575);
or U9094 (N_9094,N_4166,N_6093);
nand U9095 (N_9095,N_5767,N_4317);
and U9096 (N_9096,N_5317,N_5606);
and U9097 (N_9097,N_3280,N_4868);
xor U9098 (N_9098,N_3668,N_6185);
or U9099 (N_9099,N_5260,N_3130);
or U9100 (N_9100,N_5187,N_3792);
nor U9101 (N_9101,N_3340,N_5566);
or U9102 (N_9102,N_5087,N_5454);
xor U9103 (N_9103,N_5862,N_5424);
xnor U9104 (N_9104,N_5369,N_4246);
or U9105 (N_9105,N_5374,N_6220);
nand U9106 (N_9106,N_4249,N_3516);
or U9107 (N_9107,N_4349,N_4971);
nor U9108 (N_9108,N_5578,N_4783);
nor U9109 (N_9109,N_4165,N_3259);
nand U9110 (N_9110,N_3340,N_5784);
or U9111 (N_9111,N_4611,N_3789);
nor U9112 (N_9112,N_4388,N_4178);
or U9113 (N_9113,N_4587,N_4060);
and U9114 (N_9114,N_4180,N_5005);
nor U9115 (N_9115,N_6177,N_5950);
or U9116 (N_9116,N_6122,N_5795);
nand U9117 (N_9117,N_5791,N_3787);
and U9118 (N_9118,N_5758,N_4389);
nand U9119 (N_9119,N_5353,N_6147);
nor U9120 (N_9120,N_5537,N_3153);
nand U9121 (N_9121,N_4978,N_4001);
xor U9122 (N_9122,N_5650,N_3805);
and U9123 (N_9123,N_5926,N_4020);
and U9124 (N_9124,N_5809,N_6162);
and U9125 (N_9125,N_4966,N_5939);
or U9126 (N_9126,N_5384,N_5451);
or U9127 (N_9127,N_3732,N_5620);
nor U9128 (N_9128,N_5718,N_5737);
and U9129 (N_9129,N_5492,N_5601);
nor U9130 (N_9130,N_5050,N_3293);
and U9131 (N_9131,N_3717,N_4306);
or U9132 (N_9132,N_4780,N_4272);
nand U9133 (N_9133,N_4121,N_3199);
and U9134 (N_9134,N_5636,N_5205);
or U9135 (N_9135,N_4487,N_3724);
nor U9136 (N_9136,N_3345,N_5843);
nand U9137 (N_9137,N_5374,N_5673);
nor U9138 (N_9138,N_3254,N_4975);
and U9139 (N_9139,N_3582,N_3386);
or U9140 (N_9140,N_5450,N_3764);
nand U9141 (N_9141,N_4922,N_4450);
nor U9142 (N_9142,N_5133,N_4747);
and U9143 (N_9143,N_5121,N_4254);
or U9144 (N_9144,N_4579,N_5464);
nor U9145 (N_9145,N_5362,N_4680);
and U9146 (N_9146,N_5089,N_4717);
and U9147 (N_9147,N_4981,N_4474);
and U9148 (N_9148,N_5652,N_3495);
nor U9149 (N_9149,N_3558,N_3429);
or U9150 (N_9150,N_4722,N_5804);
and U9151 (N_9151,N_3255,N_5395);
xnor U9152 (N_9152,N_4079,N_5877);
nand U9153 (N_9153,N_3310,N_4639);
nand U9154 (N_9154,N_4601,N_5468);
and U9155 (N_9155,N_3949,N_3377);
nand U9156 (N_9156,N_4780,N_4935);
xor U9157 (N_9157,N_4943,N_4986);
or U9158 (N_9158,N_5725,N_5042);
and U9159 (N_9159,N_5435,N_3486);
nor U9160 (N_9160,N_3676,N_3881);
nand U9161 (N_9161,N_4077,N_3350);
and U9162 (N_9162,N_4362,N_6142);
nor U9163 (N_9163,N_4680,N_5368);
and U9164 (N_9164,N_3714,N_4519);
nand U9165 (N_9165,N_3244,N_4628);
nor U9166 (N_9166,N_6238,N_3744);
nor U9167 (N_9167,N_5821,N_5703);
nor U9168 (N_9168,N_4490,N_3340);
xor U9169 (N_9169,N_4626,N_4962);
or U9170 (N_9170,N_3311,N_5194);
nor U9171 (N_9171,N_4663,N_4574);
nor U9172 (N_9172,N_4659,N_6079);
nor U9173 (N_9173,N_5852,N_5558);
and U9174 (N_9174,N_5530,N_6068);
and U9175 (N_9175,N_4400,N_5708);
nand U9176 (N_9176,N_3565,N_4979);
nor U9177 (N_9177,N_3432,N_3217);
or U9178 (N_9178,N_6040,N_4706);
xor U9179 (N_9179,N_3887,N_3759);
nand U9180 (N_9180,N_3736,N_4274);
nor U9181 (N_9181,N_5421,N_3619);
nor U9182 (N_9182,N_4536,N_3427);
and U9183 (N_9183,N_3881,N_3208);
nand U9184 (N_9184,N_6183,N_4050);
or U9185 (N_9185,N_4441,N_4028);
nand U9186 (N_9186,N_5053,N_5964);
nand U9187 (N_9187,N_4574,N_3566);
or U9188 (N_9188,N_3495,N_5943);
or U9189 (N_9189,N_4145,N_4199);
xor U9190 (N_9190,N_6212,N_5561);
nand U9191 (N_9191,N_3213,N_3732);
nor U9192 (N_9192,N_3793,N_6202);
or U9193 (N_9193,N_5117,N_5587);
nor U9194 (N_9194,N_5113,N_4156);
or U9195 (N_9195,N_3379,N_5998);
and U9196 (N_9196,N_4426,N_3687);
or U9197 (N_9197,N_3376,N_5297);
and U9198 (N_9198,N_4189,N_5917);
nor U9199 (N_9199,N_3825,N_3495);
or U9200 (N_9200,N_5536,N_3525);
and U9201 (N_9201,N_4177,N_5819);
nor U9202 (N_9202,N_6031,N_5203);
nor U9203 (N_9203,N_4828,N_6107);
and U9204 (N_9204,N_4544,N_5877);
nand U9205 (N_9205,N_5038,N_4751);
or U9206 (N_9206,N_5560,N_5208);
nand U9207 (N_9207,N_4813,N_4359);
nand U9208 (N_9208,N_4877,N_3812);
nor U9209 (N_9209,N_5970,N_4236);
and U9210 (N_9210,N_4167,N_3336);
or U9211 (N_9211,N_5157,N_3259);
nor U9212 (N_9212,N_5249,N_4131);
nor U9213 (N_9213,N_3566,N_3320);
xor U9214 (N_9214,N_5839,N_5617);
and U9215 (N_9215,N_4027,N_5283);
and U9216 (N_9216,N_4617,N_4640);
nand U9217 (N_9217,N_4651,N_5944);
or U9218 (N_9218,N_4104,N_3356);
or U9219 (N_9219,N_3674,N_5505);
nor U9220 (N_9220,N_5624,N_5606);
and U9221 (N_9221,N_6153,N_3544);
nand U9222 (N_9222,N_5819,N_4984);
nor U9223 (N_9223,N_4845,N_3920);
and U9224 (N_9224,N_6096,N_5352);
xnor U9225 (N_9225,N_4806,N_4086);
nand U9226 (N_9226,N_5337,N_5979);
nor U9227 (N_9227,N_3804,N_5019);
and U9228 (N_9228,N_3639,N_5152);
or U9229 (N_9229,N_3994,N_5354);
and U9230 (N_9230,N_6150,N_4092);
or U9231 (N_9231,N_5843,N_3288);
nor U9232 (N_9232,N_4358,N_4178);
nor U9233 (N_9233,N_3512,N_5134);
and U9234 (N_9234,N_4278,N_5044);
nor U9235 (N_9235,N_3762,N_4744);
xnor U9236 (N_9236,N_5304,N_5718);
nor U9237 (N_9237,N_4587,N_5905);
and U9238 (N_9238,N_4305,N_3477);
nand U9239 (N_9239,N_3271,N_3874);
or U9240 (N_9240,N_5881,N_4815);
xnor U9241 (N_9241,N_3628,N_5209);
xor U9242 (N_9242,N_4254,N_4839);
or U9243 (N_9243,N_4681,N_5577);
or U9244 (N_9244,N_4029,N_3763);
nand U9245 (N_9245,N_3156,N_3787);
and U9246 (N_9246,N_5417,N_5332);
or U9247 (N_9247,N_5307,N_5046);
nor U9248 (N_9248,N_3807,N_3877);
or U9249 (N_9249,N_5957,N_3932);
and U9250 (N_9250,N_5078,N_4845);
xor U9251 (N_9251,N_5966,N_5164);
or U9252 (N_9252,N_4031,N_4320);
or U9253 (N_9253,N_3562,N_6113);
or U9254 (N_9254,N_5516,N_3297);
and U9255 (N_9255,N_3487,N_4994);
or U9256 (N_9256,N_5095,N_4605);
nand U9257 (N_9257,N_4025,N_5701);
and U9258 (N_9258,N_4714,N_3595);
nand U9259 (N_9259,N_3304,N_5681);
nor U9260 (N_9260,N_6096,N_5912);
nor U9261 (N_9261,N_3574,N_4780);
and U9262 (N_9262,N_3232,N_5285);
nor U9263 (N_9263,N_6062,N_4432);
or U9264 (N_9264,N_5603,N_5233);
or U9265 (N_9265,N_4035,N_4879);
or U9266 (N_9266,N_4796,N_3429);
or U9267 (N_9267,N_3400,N_6137);
xor U9268 (N_9268,N_3213,N_3623);
xor U9269 (N_9269,N_6123,N_3243);
or U9270 (N_9270,N_3772,N_3938);
or U9271 (N_9271,N_6170,N_5987);
or U9272 (N_9272,N_4368,N_4168);
and U9273 (N_9273,N_5592,N_3285);
and U9274 (N_9274,N_4558,N_4555);
nor U9275 (N_9275,N_5472,N_4118);
nor U9276 (N_9276,N_5563,N_3498);
or U9277 (N_9277,N_6240,N_3761);
nand U9278 (N_9278,N_5358,N_5572);
and U9279 (N_9279,N_4786,N_6053);
nor U9280 (N_9280,N_5733,N_5517);
nand U9281 (N_9281,N_3733,N_5804);
nand U9282 (N_9282,N_5898,N_5863);
nand U9283 (N_9283,N_5320,N_3500);
xnor U9284 (N_9284,N_3628,N_5820);
xor U9285 (N_9285,N_4276,N_5177);
nor U9286 (N_9286,N_4294,N_5491);
nor U9287 (N_9287,N_4982,N_6057);
nor U9288 (N_9288,N_4842,N_3833);
nor U9289 (N_9289,N_5645,N_5016);
or U9290 (N_9290,N_5608,N_6166);
nand U9291 (N_9291,N_3831,N_3760);
xnor U9292 (N_9292,N_4515,N_4390);
nand U9293 (N_9293,N_5501,N_6058);
or U9294 (N_9294,N_6093,N_4989);
or U9295 (N_9295,N_6152,N_4790);
nand U9296 (N_9296,N_3937,N_3855);
nand U9297 (N_9297,N_6067,N_6153);
xnor U9298 (N_9298,N_4358,N_3786);
nand U9299 (N_9299,N_5811,N_4858);
or U9300 (N_9300,N_4083,N_5746);
and U9301 (N_9301,N_3806,N_4630);
nor U9302 (N_9302,N_4549,N_5051);
and U9303 (N_9303,N_5852,N_4763);
xor U9304 (N_9304,N_4524,N_5789);
or U9305 (N_9305,N_3865,N_3408);
nand U9306 (N_9306,N_3781,N_5561);
or U9307 (N_9307,N_4789,N_3569);
nand U9308 (N_9308,N_3997,N_4385);
xnor U9309 (N_9309,N_5436,N_3613);
nor U9310 (N_9310,N_4946,N_3913);
nand U9311 (N_9311,N_3591,N_6084);
nand U9312 (N_9312,N_5629,N_3689);
nor U9313 (N_9313,N_4530,N_6198);
and U9314 (N_9314,N_3204,N_5477);
and U9315 (N_9315,N_4470,N_3275);
and U9316 (N_9316,N_3772,N_6166);
and U9317 (N_9317,N_4697,N_5268);
and U9318 (N_9318,N_3164,N_6201);
nor U9319 (N_9319,N_3151,N_3456);
nand U9320 (N_9320,N_3806,N_5862);
and U9321 (N_9321,N_4673,N_3273);
xor U9322 (N_9322,N_4965,N_3632);
nand U9323 (N_9323,N_3282,N_3472);
or U9324 (N_9324,N_4214,N_5100);
and U9325 (N_9325,N_6203,N_5380);
xnor U9326 (N_9326,N_4040,N_3385);
nor U9327 (N_9327,N_4562,N_3265);
nand U9328 (N_9328,N_3802,N_3524);
or U9329 (N_9329,N_5139,N_3953);
or U9330 (N_9330,N_5353,N_5598);
nand U9331 (N_9331,N_5166,N_4694);
nor U9332 (N_9332,N_5621,N_3238);
and U9333 (N_9333,N_6093,N_5444);
or U9334 (N_9334,N_4321,N_4092);
and U9335 (N_9335,N_5288,N_5254);
and U9336 (N_9336,N_5868,N_4834);
or U9337 (N_9337,N_6220,N_4533);
and U9338 (N_9338,N_5519,N_3224);
nand U9339 (N_9339,N_3970,N_5127);
or U9340 (N_9340,N_3685,N_4398);
and U9341 (N_9341,N_3718,N_4770);
nor U9342 (N_9342,N_3604,N_3204);
nor U9343 (N_9343,N_3814,N_4442);
nor U9344 (N_9344,N_3579,N_3212);
or U9345 (N_9345,N_4018,N_4900);
nand U9346 (N_9346,N_4192,N_5771);
nand U9347 (N_9347,N_3913,N_6047);
and U9348 (N_9348,N_3750,N_5827);
and U9349 (N_9349,N_3726,N_3807);
nand U9350 (N_9350,N_4355,N_4748);
or U9351 (N_9351,N_5328,N_4153);
or U9352 (N_9352,N_6243,N_5593);
nand U9353 (N_9353,N_4045,N_6158);
xor U9354 (N_9354,N_5223,N_4740);
nor U9355 (N_9355,N_5370,N_4402);
and U9356 (N_9356,N_3251,N_5263);
and U9357 (N_9357,N_5020,N_3266);
nor U9358 (N_9358,N_4348,N_3671);
or U9359 (N_9359,N_5219,N_3513);
nor U9360 (N_9360,N_4114,N_3732);
and U9361 (N_9361,N_5047,N_5730);
or U9362 (N_9362,N_5974,N_4947);
or U9363 (N_9363,N_4328,N_3747);
nor U9364 (N_9364,N_5873,N_5564);
or U9365 (N_9365,N_5992,N_4380);
and U9366 (N_9366,N_5834,N_5960);
and U9367 (N_9367,N_3495,N_4321);
nand U9368 (N_9368,N_3892,N_4427);
or U9369 (N_9369,N_4505,N_5311);
or U9370 (N_9370,N_4733,N_4588);
nand U9371 (N_9371,N_6237,N_5970);
or U9372 (N_9372,N_5882,N_4671);
or U9373 (N_9373,N_4007,N_4904);
nand U9374 (N_9374,N_6188,N_6119);
nor U9375 (N_9375,N_7042,N_7465);
nand U9376 (N_9376,N_7723,N_7611);
and U9377 (N_9377,N_7250,N_6579);
and U9378 (N_9378,N_7526,N_9182);
or U9379 (N_9379,N_8368,N_6362);
xor U9380 (N_9380,N_7629,N_8364);
and U9381 (N_9381,N_8761,N_9064);
and U9382 (N_9382,N_6940,N_7527);
nand U9383 (N_9383,N_8358,N_6492);
and U9384 (N_9384,N_9018,N_8956);
or U9385 (N_9385,N_7531,N_7539);
xor U9386 (N_9386,N_7325,N_6517);
or U9387 (N_9387,N_8806,N_7862);
nor U9388 (N_9388,N_8402,N_9042);
xnor U9389 (N_9389,N_9045,N_6439);
nor U9390 (N_9390,N_8188,N_8271);
and U9391 (N_9391,N_7841,N_6381);
or U9392 (N_9392,N_6534,N_8598);
or U9393 (N_9393,N_8937,N_8419);
and U9394 (N_9394,N_7508,N_8820);
or U9395 (N_9395,N_8818,N_9370);
and U9396 (N_9396,N_7823,N_7356);
nor U9397 (N_9397,N_6435,N_6327);
nand U9398 (N_9398,N_7968,N_8879);
or U9399 (N_9399,N_8672,N_6460);
xnor U9400 (N_9400,N_6514,N_8446);
or U9401 (N_9401,N_6309,N_9242);
nor U9402 (N_9402,N_8864,N_8670);
nor U9403 (N_9403,N_7678,N_8757);
nor U9404 (N_9404,N_7159,N_8284);
and U9405 (N_9405,N_8273,N_8390);
nand U9406 (N_9406,N_8912,N_6795);
nand U9407 (N_9407,N_8294,N_8308);
nor U9408 (N_9408,N_8160,N_7446);
nor U9409 (N_9409,N_6403,N_8902);
or U9410 (N_9410,N_6556,N_7610);
nor U9411 (N_9411,N_6464,N_8771);
nor U9412 (N_9412,N_6284,N_8023);
nand U9413 (N_9413,N_7075,N_6837);
nor U9414 (N_9414,N_8449,N_8957);
nor U9415 (N_9415,N_7914,N_7309);
nor U9416 (N_9416,N_8240,N_7009);
and U9417 (N_9417,N_8664,N_6920);
nand U9418 (N_9418,N_6694,N_6800);
nand U9419 (N_9419,N_7580,N_7085);
or U9420 (N_9420,N_6443,N_6322);
nand U9421 (N_9421,N_7155,N_9146);
nor U9422 (N_9422,N_8319,N_6640);
or U9423 (N_9423,N_6862,N_9207);
nor U9424 (N_9424,N_7944,N_6298);
or U9425 (N_9425,N_9154,N_6393);
xor U9426 (N_9426,N_7530,N_6814);
or U9427 (N_9427,N_6392,N_8648);
or U9428 (N_9428,N_9253,N_7910);
or U9429 (N_9429,N_7813,N_6421);
nor U9430 (N_9430,N_6723,N_8790);
and U9431 (N_9431,N_8517,N_6567);
nor U9432 (N_9432,N_9195,N_6949);
or U9433 (N_9433,N_8293,N_8016);
xor U9434 (N_9434,N_8650,N_9280);
or U9435 (N_9435,N_8069,N_7570);
nor U9436 (N_9436,N_7206,N_7463);
or U9437 (N_9437,N_6356,N_7421);
or U9438 (N_9438,N_7341,N_8719);
xor U9439 (N_9439,N_7403,N_8167);
nor U9440 (N_9440,N_8909,N_6951);
xnor U9441 (N_9441,N_7943,N_8387);
and U9442 (N_9442,N_7670,N_7899);
and U9443 (N_9443,N_8625,N_7761);
nor U9444 (N_9444,N_9362,N_6319);
nand U9445 (N_9445,N_6876,N_7495);
or U9446 (N_9446,N_8888,N_7077);
nor U9447 (N_9447,N_7415,N_7783);
nand U9448 (N_9448,N_9212,N_6527);
nand U9449 (N_9449,N_8137,N_8938);
or U9450 (N_9450,N_8378,N_9032);
nand U9451 (N_9451,N_7193,N_6990);
nand U9452 (N_9452,N_8635,N_7971);
and U9453 (N_9453,N_9368,N_6830);
or U9454 (N_9454,N_6373,N_8191);
and U9455 (N_9455,N_6615,N_9299);
and U9456 (N_9456,N_8179,N_8389);
nor U9457 (N_9457,N_8032,N_8923);
or U9458 (N_9458,N_7828,N_7467);
nor U9459 (N_9459,N_7171,N_7079);
and U9460 (N_9460,N_8096,N_6497);
xnor U9461 (N_9461,N_7080,N_9246);
xor U9462 (N_9462,N_9293,N_9098);
nand U9463 (N_9463,N_8576,N_8758);
or U9464 (N_9464,N_7811,N_8425);
xor U9465 (N_9465,N_7252,N_6646);
and U9466 (N_9466,N_8241,N_7720);
or U9467 (N_9467,N_7787,N_6467);
or U9468 (N_9468,N_9282,N_7614);
or U9469 (N_9469,N_7868,N_7220);
nor U9470 (N_9470,N_9174,N_8507);
and U9471 (N_9471,N_6960,N_8537);
nand U9472 (N_9472,N_8285,N_9155);
nor U9473 (N_9473,N_8875,N_6654);
and U9474 (N_9474,N_8570,N_7615);
nand U9475 (N_9475,N_7988,N_6890);
and U9476 (N_9476,N_7638,N_8014);
nand U9477 (N_9477,N_8680,N_7168);
nor U9478 (N_9478,N_7843,N_9294);
or U9479 (N_9479,N_9164,N_9276);
or U9480 (N_9480,N_8310,N_6907);
nand U9481 (N_9481,N_7222,N_7386);
or U9482 (N_9482,N_6746,N_7151);
and U9483 (N_9483,N_9260,N_8227);
nand U9484 (N_9484,N_6906,N_7141);
and U9485 (N_9485,N_7507,N_7484);
nor U9486 (N_9486,N_7546,N_7249);
xor U9487 (N_9487,N_9076,N_8990);
nor U9488 (N_9488,N_8590,N_7837);
xnor U9489 (N_9489,N_7535,N_8185);
and U9490 (N_9490,N_7086,N_6379);
or U9491 (N_9491,N_6871,N_8954);
nand U9492 (N_9492,N_7722,N_7390);
or U9493 (N_9493,N_7644,N_7095);
or U9494 (N_9494,N_8184,N_7959);
nor U9495 (N_9495,N_7822,N_8560);
or U9496 (N_9496,N_6698,N_8112);
or U9497 (N_9497,N_7800,N_6586);
and U9498 (N_9498,N_6677,N_7450);
xnor U9499 (N_9499,N_6748,N_7596);
and U9500 (N_9500,N_6589,N_8101);
nand U9501 (N_9501,N_8165,N_6751);
nand U9502 (N_9502,N_6543,N_8600);
nand U9503 (N_9503,N_8058,N_7618);
or U9504 (N_9504,N_9129,N_6399);
nor U9505 (N_9505,N_6669,N_8151);
and U9506 (N_9506,N_6338,N_7270);
nor U9507 (N_9507,N_7634,N_8838);
and U9508 (N_9508,N_8350,N_8495);
and U9509 (N_9509,N_9215,N_7917);
nor U9510 (N_9510,N_6518,N_8655);
nor U9511 (N_9511,N_9308,N_6811);
nor U9512 (N_9512,N_8638,N_7461);
nor U9513 (N_9513,N_8244,N_7926);
nand U9514 (N_9514,N_6550,N_7727);
and U9515 (N_9515,N_9204,N_6537);
and U9516 (N_9516,N_7370,N_9340);
or U9517 (N_9517,N_6482,N_6509);
nor U9518 (N_9518,N_7902,N_7040);
and U9519 (N_9519,N_7200,N_8707);
nand U9520 (N_9520,N_6846,N_7778);
nand U9521 (N_9521,N_6584,N_9249);
xor U9522 (N_9522,N_7442,N_8235);
and U9523 (N_9523,N_8824,N_8252);
nand U9524 (N_9524,N_9345,N_8012);
xnor U9525 (N_9525,N_6348,N_8817);
or U9526 (N_9526,N_6899,N_8815);
or U9527 (N_9527,N_7651,N_9237);
nor U9528 (N_9528,N_7806,N_6858);
nand U9529 (N_9529,N_6511,N_8287);
or U9530 (N_9530,N_6821,N_7675);
nor U9531 (N_9531,N_8970,N_6981);
nand U9532 (N_9532,N_8582,N_8504);
nand U9533 (N_9533,N_7032,N_8836);
and U9534 (N_9534,N_6732,N_6630);
or U9535 (N_9535,N_6786,N_7205);
xor U9536 (N_9536,N_6258,N_8437);
and U9537 (N_9537,N_6631,N_6813);
or U9538 (N_9538,N_7276,N_7329);
nor U9539 (N_9539,N_7107,N_7848);
and U9540 (N_9540,N_8343,N_9248);
xnor U9541 (N_9541,N_8667,N_8053);
nand U9542 (N_9542,N_9097,N_7704);
nand U9543 (N_9543,N_7184,N_8456);
nand U9544 (N_9544,N_8626,N_9144);
nor U9545 (N_9545,N_6402,N_9319);
nand U9546 (N_9546,N_6715,N_7517);
nand U9547 (N_9547,N_8086,N_7267);
xor U9548 (N_9548,N_8210,N_9329);
or U9549 (N_9549,N_6962,N_8386);
or U9550 (N_9550,N_6691,N_7133);
and U9551 (N_9551,N_9092,N_6977);
nand U9552 (N_9552,N_6323,N_7850);
nor U9553 (N_9553,N_8519,N_7440);
nand U9554 (N_9554,N_6726,N_7647);
nor U9555 (N_9555,N_8653,N_7524);
nand U9556 (N_9556,N_7795,N_9017);
xnor U9557 (N_9557,N_7585,N_8445);
xor U9558 (N_9558,N_8769,N_6620);
nand U9559 (N_9559,N_7738,N_6762);
and U9560 (N_9560,N_7594,N_7542);
and U9561 (N_9561,N_6538,N_6848);
and U9562 (N_9562,N_6847,N_7877);
and U9563 (N_9563,N_7802,N_6626);
nand U9564 (N_9564,N_6883,N_7472);
or U9565 (N_9565,N_6891,N_6695);
or U9566 (N_9566,N_8860,N_8300);
nand U9567 (N_9567,N_9219,N_7181);
or U9568 (N_9568,N_8286,N_8298);
and U9569 (N_9569,N_7924,N_7096);
and U9570 (N_9570,N_6581,N_8347);
nor U9571 (N_9571,N_8391,N_9348);
xor U9572 (N_9572,N_7545,N_6855);
nor U9573 (N_9573,N_7895,N_8931);
and U9574 (N_9574,N_7257,N_8475);
or U9575 (N_9575,N_9229,N_8780);
nand U9576 (N_9576,N_8070,N_8976);
or U9577 (N_9577,N_6599,N_7069);
nor U9578 (N_9578,N_9022,N_7555);
nor U9579 (N_9579,N_6875,N_6828);
or U9580 (N_9580,N_7058,N_6588);
and U9581 (N_9581,N_8968,N_6461);
nand U9582 (N_9582,N_7713,N_7881);
and U9583 (N_9583,N_9305,N_9016);
or U9584 (N_9584,N_9354,N_7093);
and U9585 (N_9585,N_7127,N_8066);
nand U9586 (N_9586,N_7488,N_8479);
and U9587 (N_9587,N_7278,N_7012);
nand U9588 (N_9588,N_7046,N_8181);
xor U9589 (N_9589,N_8833,N_6470);
or U9590 (N_9590,N_7504,N_8356);
nor U9591 (N_9591,N_7265,N_9178);
nand U9592 (N_9592,N_6354,N_6820);
or U9593 (N_9593,N_8804,N_8708);
xnor U9594 (N_9594,N_7909,N_7664);
xor U9595 (N_9595,N_8334,N_6713);
xor U9596 (N_9596,N_8321,N_7221);
or U9597 (N_9597,N_7563,N_8313);
and U9598 (N_9598,N_8071,N_7029);
and U9599 (N_9599,N_7103,N_9287);
nand U9600 (N_9600,N_8048,N_8760);
and U9601 (N_9601,N_6709,N_8972);
and U9602 (N_9602,N_7575,N_6616);
or U9603 (N_9603,N_7204,N_8764);
and U9604 (N_9604,N_6682,N_8890);
or U9605 (N_9605,N_8506,N_7589);
nand U9606 (N_9606,N_8718,N_7553);
and U9607 (N_9607,N_7426,N_8794);
or U9608 (N_9608,N_8684,N_8800);
or U9609 (N_9609,N_7853,N_7842);
nor U9610 (N_9610,N_8554,N_7925);
or U9611 (N_9611,N_7211,N_7769);
nand U9612 (N_9612,N_7662,N_8778);
and U9613 (N_9613,N_7225,N_6498);
nand U9614 (N_9614,N_6448,N_7964);
or U9615 (N_9615,N_7581,N_6851);
or U9616 (N_9616,N_8689,N_7289);
nor U9617 (N_9617,N_6295,N_7084);
nand U9618 (N_9618,N_9044,N_7963);
nor U9619 (N_9619,N_7628,N_7339);
nand U9620 (N_9620,N_8835,N_8630);
and U9621 (N_9621,N_8127,N_6635);
and U9622 (N_9622,N_8601,N_8195);
and U9623 (N_9623,N_8589,N_6427);
xor U9624 (N_9624,N_8644,N_8398);
nor U9625 (N_9625,N_7477,N_8340);
nand U9626 (N_9626,N_8255,N_8631);
and U9627 (N_9627,N_7021,N_8197);
nand U9628 (N_9628,N_7398,N_7473);
nor U9629 (N_9629,N_7956,N_8234);
nand U9630 (N_9630,N_7022,N_7226);
nand U9631 (N_9631,N_6844,N_8460);
nor U9632 (N_9632,N_7344,N_7750);
and U9633 (N_9633,N_7153,N_7897);
nand U9634 (N_9634,N_8779,N_7790);
nor U9635 (N_9635,N_7516,N_7346);
or U9636 (N_9636,N_8344,N_9245);
or U9637 (N_9637,N_6803,N_9190);
and U9638 (N_9638,N_7468,N_8455);
nand U9639 (N_9639,N_9366,N_6401);
nor U9640 (N_9640,N_8411,N_7561);
nor U9641 (N_9641,N_7019,N_8503);
and U9642 (N_9642,N_8816,N_8700);
nand U9643 (N_9643,N_8556,N_7500);
or U9644 (N_9644,N_9310,N_6783);
xnor U9645 (N_9645,N_8702,N_6739);
nand U9646 (N_9646,N_6566,N_8588);
or U9647 (N_9647,N_6915,N_7846);
nor U9648 (N_9648,N_9119,N_8772);
nand U9649 (N_9649,N_6604,N_7810);
nand U9650 (N_9650,N_7711,N_8637);
or U9651 (N_9651,N_7100,N_8480);
nor U9652 (N_9652,N_7701,N_8033);
xnor U9653 (N_9653,N_6596,N_7824);
nand U9654 (N_9654,N_9250,N_9373);
or U9655 (N_9655,N_7026,N_6299);
xor U9656 (N_9656,N_7799,N_6359);
nor U9657 (N_9657,N_8567,N_6325);
and U9658 (N_9658,N_6572,N_6312);
or U9659 (N_9659,N_8125,N_8499);
nand U9660 (N_9660,N_8327,N_8073);
nand U9661 (N_9661,N_6539,N_9316);
and U9662 (N_9662,N_8385,N_8049);
and U9663 (N_9663,N_8921,N_7432);
xor U9664 (N_9664,N_8516,N_8855);
and U9665 (N_9665,N_6430,N_8738);
xor U9666 (N_9666,N_6911,N_6655);
or U9667 (N_9667,N_7246,N_6928);
nor U9668 (N_9668,N_8647,N_8302);
or U9669 (N_9669,N_7937,N_6363);
nand U9670 (N_9670,N_8842,N_7751);
or U9671 (N_9671,N_6866,N_7203);
nor U9672 (N_9672,N_7933,N_8652);
or U9673 (N_9673,N_8254,N_6597);
nand U9674 (N_9674,N_7893,N_8064);
nand U9675 (N_9675,N_8010,N_8353);
nor U9676 (N_9676,N_7719,N_7429);
nand U9677 (N_9677,N_7891,N_7401);
nor U9678 (N_9678,N_7603,N_8412);
nand U9679 (N_9679,N_6457,N_8553);
and U9680 (N_9680,N_7187,N_9341);
nand U9681 (N_9681,N_7873,N_7927);
and U9682 (N_9682,N_8436,N_6884);
nor U9683 (N_9683,N_8314,N_9079);
and U9684 (N_9684,N_8427,N_7299);
or U9685 (N_9685,N_8533,N_7152);
nor U9686 (N_9686,N_8654,N_8575);
and U9687 (N_9687,N_6958,N_6303);
and U9688 (N_9688,N_6600,N_6838);
nor U9689 (N_9689,N_9189,N_8805);
or U9690 (N_9690,N_7202,N_8896);
and U9691 (N_9691,N_6510,N_6384);
and U9692 (N_9692,N_7875,N_7852);
nor U9693 (N_9693,N_9109,N_6921);
xnor U9694 (N_9694,N_9241,N_6361);
and U9695 (N_9695,N_9014,N_6488);
nor U9696 (N_9696,N_6781,N_8607);
xor U9697 (N_9697,N_9142,N_8936);
or U9698 (N_9698,N_8062,N_8220);
nor U9699 (N_9699,N_9012,N_6856);
xor U9700 (N_9700,N_8279,N_6693);
or U9701 (N_9701,N_6346,N_8611);
and U9702 (N_9702,N_7113,N_8737);
nand U9703 (N_9703,N_7903,N_6557);
nand U9704 (N_9704,N_6901,N_6852);
or U9705 (N_9705,N_7595,N_8004);
or U9706 (N_9706,N_6975,N_7300);
nor U9707 (N_9707,N_7164,N_7118);
or U9708 (N_9708,N_6668,N_8483);
xnor U9709 (N_9709,N_8682,N_8563);
xnor U9710 (N_9710,N_8116,N_7597);
or U9711 (N_9711,N_6500,N_6993);
and U9712 (N_9712,N_9179,N_6913);
nand U9713 (N_9713,N_6255,N_8376);
nand U9714 (N_9714,N_9027,N_6274);
nand U9715 (N_9715,N_7115,N_6663);
or U9716 (N_9716,N_8548,N_7537);
nor U9717 (N_9717,N_8162,N_7345);
or U9718 (N_9718,N_9001,N_7218);
or U9719 (N_9719,N_9325,N_7502);
or U9720 (N_9720,N_6397,N_7287);
nand U9721 (N_9721,N_8180,N_7682);
and U9722 (N_9722,N_6853,N_7142);
and U9723 (N_9723,N_8852,N_8424);
or U9724 (N_9724,N_6825,N_8819);
and U9725 (N_9725,N_9166,N_8336);
and U9726 (N_9726,N_6903,N_9257);
and U9727 (N_9727,N_8623,N_7143);
or U9728 (N_9728,N_6347,N_6969);
nor U9729 (N_9729,N_8546,N_6914);
or U9730 (N_9730,N_9176,N_8617);
or U9731 (N_9731,N_7528,N_9162);
nand U9732 (N_9732,N_9073,N_7260);
or U9733 (N_9733,N_8793,N_7389);
nor U9734 (N_9734,N_8950,N_7420);
or U9735 (N_9735,N_8155,N_6269);
nor U9736 (N_9736,N_6545,N_6657);
xor U9737 (N_9737,N_6938,N_8782);
or U9738 (N_9738,N_8512,N_7489);
and U9739 (N_9739,N_6744,N_7134);
nand U9740 (N_9740,N_8774,N_6519);
or U9741 (N_9741,N_7938,N_8669);
or U9742 (N_9742,N_6730,N_6313);
nand U9743 (N_9743,N_8742,N_6777);
or U9744 (N_9744,N_8106,N_9095);
or U9745 (N_9745,N_7957,N_8482);
and U9746 (N_9746,N_8551,N_7631);
nor U9747 (N_9747,N_8001,N_6861);
and U9748 (N_9748,N_8018,N_8857);
and U9749 (N_9749,N_7369,N_7241);
or U9750 (N_9750,N_6614,N_7251);
nor U9751 (N_9751,N_6704,N_6967);
nand U9752 (N_9752,N_7213,N_7407);
nand U9753 (N_9753,N_6585,N_6923);
and U9754 (N_9754,N_7612,N_6966);
xnor U9755 (N_9755,N_9202,N_7292);
nor U9756 (N_9756,N_8126,N_8372);
nor U9757 (N_9757,N_7905,N_8943);
xnor U9758 (N_9758,N_7665,N_7397);
nor U9759 (N_9759,N_9235,N_7510);
nand U9760 (N_9760,N_6377,N_8699);
xor U9761 (N_9761,N_6441,N_7471);
nand U9762 (N_9762,N_7636,N_6449);
or U9763 (N_9763,N_7364,N_7742);
and U9764 (N_9764,N_7577,N_9297);
nor U9765 (N_9765,N_9284,N_7781);
nand U9766 (N_9766,N_7695,N_8107);
or U9767 (N_9767,N_6477,N_8691);
xor U9768 (N_9768,N_9364,N_9055);
and U9769 (N_9769,N_7643,N_7734);
nand U9770 (N_9770,N_8170,N_8930);
or U9771 (N_9771,N_7598,N_9254);
or U9772 (N_9772,N_6963,N_7900);
and U9773 (N_9773,N_6289,N_8196);
and U9774 (N_9774,N_6308,N_6973);
or U9775 (N_9775,N_8434,N_8426);
or U9776 (N_9776,N_8830,N_9331);
nor U9777 (N_9777,N_8924,N_8296);
nand U9778 (N_9778,N_7915,N_8122);
and U9779 (N_9779,N_7703,N_8187);
and U9780 (N_9780,N_9118,N_8253);
or U9781 (N_9781,N_7583,N_8612);
nand U9782 (N_9782,N_7316,N_7335);
or U9783 (N_9783,N_8939,N_6957);
nor U9784 (N_9784,N_6612,N_8510);
or U9785 (N_9785,N_7874,N_8881);
and U9786 (N_9786,N_7175,N_8174);
or U9787 (N_9787,N_8593,N_8995);
and U9788 (N_9788,N_7515,N_7074);
and U9789 (N_9789,N_8451,N_9301);
or U9790 (N_9790,N_8734,N_8743);
and U9791 (N_9791,N_8850,N_7499);
and U9792 (N_9792,N_7928,N_7621);
or U9793 (N_9793,N_9181,N_6650);
and U9794 (N_9794,N_6294,N_9085);
nand U9795 (N_9795,N_9337,N_7511);
and U9796 (N_9796,N_7466,N_8132);
or U9797 (N_9797,N_6961,N_6251);
nor U9798 (N_9798,N_7313,N_7448);
xnor U9799 (N_9799,N_7361,N_6782);
nand U9800 (N_9800,N_6512,N_8471);
nand U9801 (N_9801,N_9357,N_8470);
nand U9802 (N_9802,N_9049,N_9127);
nor U9803 (N_9803,N_8662,N_8869);
and U9804 (N_9804,N_7885,N_8666);
or U9805 (N_9805,N_8574,N_6678);
xnor U9806 (N_9806,N_7214,N_6341);
nand U9807 (N_9807,N_6476,N_9264);
xor U9808 (N_9808,N_8932,N_8105);
or U9809 (N_9809,N_9062,N_8231);
and U9810 (N_9810,N_8831,N_7812);
nand U9811 (N_9811,N_8534,N_6651);
nand U9812 (N_9812,N_8044,N_7840);
and U9813 (N_9813,N_8986,N_8604);
nand U9814 (N_9814,N_8728,N_8587);
nand U9815 (N_9815,N_7041,N_8673);
nand U9816 (N_9816,N_6605,N_7002);
nand U9817 (N_9817,N_9028,N_6710);
nand U9818 (N_9818,N_6302,N_7307);
and U9819 (N_9819,N_7973,N_7709);
or U9820 (N_9820,N_9259,N_6578);
and U9821 (N_9821,N_8068,N_6767);
nor U9822 (N_9822,N_7733,N_6475);
nor U9823 (N_9823,N_6653,N_9227);
or U9824 (N_9824,N_7952,N_8169);
nor U9825 (N_9825,N_6328,N_9153);
nor U9826 (N_9826,N_8660,N_6424);
and U9827 (N_9827,N_8404,N_6689);
nor U9828 (N_9828,N_7512,N_7072);
xnor U9829 (N_9829,N_6802,N_7858);
xnor U9830 (N_9830,N_6956,N_8891);
or U9831 (N_9831,N_7375,N_8320);
or U9832 (N_9832,N_7712,N_8549);
and U9833 (N_9833,N_8362,N_6388);
nand U9834 (N_9834,N_7383,N_9123);
xnor U9835 (N_9835,N_8827,N_8003);
nor U9836 (N_9836,N_9191,N_8110);
nor U9837 (N_9837,N_7690,N_8929);
xor U9838 (N_9838,N_8710,N_7784);
and U9839 (N_9839,N_8409,N_6270);
or U9840 (N_9840,N_9161,N_8982);
and U9841 (N_9841,N_7607,N_6897);
or U9842 (N_9842,N_8811,N_9145);
nand U9843 (N_9843,N_8478,N_7653);
and U9844 (N_9844,N_9105,N_8920);
and U9845 (N_9845,N_7691,N_7569);
nor U9846 (N_9846,N_7459,N_6924);
nand U9847 (N_9847,N_9196,N_7136);
nor U9848 (N_9848,N_6877,N_7324);
and U9849 (N_9849,N_8952,N_6547);
nor U9850 (N_9850,N_7892,N_8668);
nand U9851 (N_9851,N_8428,N_6278);
nand U9852 (N_9852,N_9110,N_8877);
and U9853 (N_9853,N_6807,N_7371);
nor U9854 (N_9854,N_9074,N_7384);
nand U9855 (N_9855,N_7441,N_7088);
nor U9856 (N_9856,N_8410,N_8717);
nor U9857 (N_9857,N_6394,N_6314);
or U9858 (N_9858,N_7405,N_7229);
and U9859 (N_9859,N_8215,N_8773);
and U9860 (N_9860,N_8243,N_7068);
nand U9861 (N_9861,N_9054,N_8077);
xnor U9862 (N_9862,N_8616,N_7754);
or U9863 (N_9863,N_8913,N_8304);
and U9864 (N_9864,N_9268,N_6491);
xor U9865 (N_9865,N_7391,N_7408);
nand U9866 (N_9866,N_7060,N_6880);
and U9867 (N_9867,N_8239,N_8258);
and U9868 (N_9868,N_6854,N_7280);
or U9869 (N_9869,N_8971,N_6315);
and U9870 (N_9870,N_7995,N_9283);
xor U9871 (N_9871,N_7839,N_8490);
nand U9872 (N_9872,N_9005,N_7192);
nand U9873 (N_9873,N_8569,N_9006);
nor U9874 (N_9874,N_7201,N_6559);
nor U9875 (N_9875,N_9071,N_7686);
nor U9876 (N_9876,N_8352,N_6434);
nand U9877 (N_9877,N_8887,N_6796);
nor U9878 (N_9878,N_8900,N_7648);
nor U9879 (N_9879,N_7574,N_6808);
nor U9880 (N_9880,N_8550,N_9184);
nor U9881 (N_9881,N_6874,N_9233);
or U9882 (N_9882,N_9157,N_6812);
and U9883 (N_9883,N_6280,N_7025);
nor U9884 (N_9884,N_7496,N_6860);
and U9885 (N_9885,N_8619,N_9117);
nand U9886 (N_9886,N_8401,N_8371);
or U9887 (N_9887,N_7987,N_7481);
and U9888 (N_9888,N_8661,N_8159);
or U9889 (N_9889,N_7290,N_6902);
nor U9890 (N_9890,N_7059,N_6505);
nor U9891 (N_9891,N_8658,N_6842);
nand U9892 (N_9892,N_8872,N_6942);
or U9893 (N_9893,N_8634,N_9034);
or U9894 (N_9894,N_6889,N_8984);
or U9895 (N_9895,N_9024,N_9343);
and U9896 (N_9896,N_9312,N_6624);
xor U9897 (N_9897,N_8297,N_7105);
nor U9898 (N_9898,N_9239,N_9205);
and U9899 (N_9899,N_7011,N_8208);
nor U9900 (N_9900,N_8884,N_6414);
nor U9901 (N_9901,N_8275,N_7234);
nand U9902 (N_9902,N_8380,N_6932);
and U9903 (N_9903,N_7359,N_7522);
or U9904 (N_9904,N_7626,N_7454);
nor U9905 (N_9905,N_6826,N_7692);
nor U9906 (N_9906,N_6964,N_9172);
nand U9907 (N_9907,N_9177,N_9163);
nand U9908 (N_9908,N_6987,N_6592);
xnor U9909 (N_9909,N_7239,N_7972);
xor U9910 (N_9910,N_8289,N_8212);
nand U9911 (N_9911,N_6878,N_7008);
nand U9912 (N_9912,N_8687,N_7745);
xor U9913 (N_9913,N_6641,N_6273);
xnor U9914 (N_9914,N_7036,N_8494);
and U9915 (N_9915,N_8305,N_7970);
and U9916 (N_9916,N_8733,N_8705);
nand U9917 (N_9917,N_8420,N_6420);
and U9918 (N_9918,N_7082,N_7934);
nand U9919 (N_9919,N_7419,N_7182);
xor U9920 (N_9920,N_7919,N_7039);
nor U9921 (N_9921,N_6291,N_6413);
nor U9922 (N_9922,N_7736,N_8663);
or U9923 (N_9923,N_9000,N_8632);
xnor U9924 (N_9924,N_6368,N_6804);
nor U9925 (N_9925,N_8138,N_8505);
nand U9926 (N_9926,N_8057,N_7803);
and U9927 (N_9927,N_7123,N_7102);
or U9928 (N_9928,N_7078,N_7689);
or U9929 (N_9929,N_7590,N_6935);
nand U9930 (N_9930,N_8531,N_7132);
nand U9931 (N_9931,N_8992,N_7976);
nor U9932 (N_9932,N_7993,N_6340);
and U9933 (N_9933,N_9334,N_8866);
nand U9934 (N_9934,N_7797,N_8458);
nand U9935 (N_9935,N_7998,N_6773);
and U9936 (N_9936,N_7360,N_9291);
and U9937 (N_9937,N_6410,N_7275);
nand U9938 (N_9938,N_7043,N_6575);
nand U9939 (N_9939,N_8768,N_8038);
and U9940 (N_9940,N_7668,N_8328);
and U9941 (N_9941,N_8621,N_6540);
and U9942 (N_9942,N_7235,N_7137);
or U9943 (N_9943,N_6743,N_7677);
and U9944 (N_9944,N_9252,N_7376);
nand U9945 (N_9945,N_8889,N_8147);
nand U9946 (N_9946,N_8226,N_6521);
and U9947 (N_9947,N_7263,N_9160);
nand U9948 (N_9948,N_7104,N_6644);
nand U9949 (N_9949,N_6944,N_9351);
and U9950 (N_9950,N_6916,N_8052);
or U9951 (N_9951,N_7989,N_7223);
nand U9952 (N_9952,N_9168,N_7298);
and U9953 (N_9953,N_6714,N_6406);
and U9954 (N_9954,N_9369,N_6623);
xor U9955 (N_9955,N_7438,N_6737);
nor U9956 (N_9956,N_7062,N_9170);
and U9957 (N_9957,N_8539,N_7655);
or U9958 (N_9958,N_9339,N_6771);
nand U9959 (N_9959,N_8676,N_7788);
and U9960 (N_9960,N_7097,N_8853);
nor U9961 (N_9961,N_7573,N_7955);
xnor U9962 (N_9962,N_7417,N_9167);
xnor U9963 (N_9963,N_8770,N_7098);
or U9964 (N_9964,N_6985,N_7253);
and U9965 (N_9965,N_7404,N_7550);
nand U9966 (N_9966,N_9159,N_6317);
nor U9967 (N_9967,N_7264,N_8461);
nor U9968 (N_9968,N_7023,N_7092);
nor U9969 (N_9969,N_8087,N_6790);
nor U9970 (N_9970,N_8342,N_6879);
or U9971 (N_9971,N_7741,N_8466);
nand U9972 (N_9972,N_8194,N_6984);
or U9973 (N_9973,N_8486,N_8154);
or U9974 (N_9974,N_6670,N_7625);
nor U9975 (N_9975,N_7073,N_8910);
nor U9976 (N_9976,N_9020,N_7210);
xor U9977 (N_9977,N_8749,N_9372);
nor U9978 (N_9978,N_8883,N_8514);
or U9979 (N_9979,N_6617,N_7949);
and U9980 (N_9980,N_9272,N_7174);
and U9981 (N_9981,N_8198,N_7470);
or U9982 (N_9982,N_6904,N_8435);
nand U9983 (N_9983,N_9266,N_6632);
or U9984 (N_9984,N_7282,N_8595);
nor U9985 (N_9985,N_6755,N_9061);
nand U9986 (N_9986,N_8586,N_6307);
xor U9987 (N_9987,N_6418,N_8581);
and U9988 (N_9988,N_7633,N_9203);
nand U9989 (N_9989,N_7645,N_7744);
nor U9990 (N_9990,N_7529,N_8933);
or U9991 (N_9991,N_6661,N_7310);
xnor U9992 (N_9992,N_7746,N_9009);
xnor U9993 (N_9993,N_8250,N_6285);
or U9994 (N_9994,N_9296,N_8114);
nand U9995 (N_9995,N_8642,N_8907);
and U9996 (N_9996,N_6671,N_7053);
and U9997 (N_9997,N_7558,N_9234);
or U9998 (N_9998,N_8019,N_7262);
and U9999 (N_9999,N_6367,N_6887);
xor U10000 (N_10000,N_7362,N_6840);
and U10001 (N_10001,N_6472,N_7619);
xor U10002 (N_10002,N_8735,N_6995);
nand U10003 (N_10003,N_8585,N_8246);
nor U10004 (N_10004,N_8885,N_7464);
nand U10005 (N_10005,N_8109,N_7271);
and U10006 (N_10006,N_9147,N_9226);
nand U10007 (N_10007,N_9093,N_8624);
xnor U10008 (N_10008,N_7064,N_8597);
or U10009 (N_10009,N_8843,N_7392);
nand U10010 (N_10010,N_7821,N_7962);
nor U10011 (N_10011,N_7122,N_6440);
nor U10012 (N_10012,N_9043,N_7666);
or U10013 (N_10013,N_7337,N_7560);
nand U10014 (N_10014,N_7992,N_7854);
nand U10015 (N_10015,N_7605,N_8861);
and U10016 (N_10016,N_7863,N_8508);
nor U10017 (N_10017,N_8944,N_8224);
nand U10018 (N_10018,N_9148,N_9288);
and U10019 (N_10019,N_7980,N_8894);
nor U10020 (N_10020,N_8288,N_9231);
or U10021 (N_10021,N_8379,N_7676);
nor U10022 (N_10022,N_9100,N_7879);
or U10023 (N_10023,N_7150,N_6252);
nor U10024 (N_10024,N_8094,N_7487);
nor U10025 (N_10025,N_8899,N_6666);
nor U10026 (N_10026,N_8628,N_7311);
nand U10027 (N_10027,N_6526,N_9030);
and U10028 (N_10028,N_8264,N_7483);
nand U10029 (N_10029,N_6426,N_7439);
or U10030 (N_10030,N_7209,N_8060);
or U10031 (N_10031,N_7534,N_7776);
or U10032 (N_10032,N_6996,N_8645);
and U10033 (N_10033,N_6636,N_7034);
or U10034 (N_10034,N_8878,N_7154);
nor U10035 (N_10035,N_7509,N_6728);
nor U10036 (N_10036,N_8382,N_7394);
nand U10037 (N_10037,N_8736,N_8725);
and U10038 (N_10038,N_8829,N_7749);
nand U10039 (N_10039,N_6642,N_6416);
or U10040 (N_10040,N_7694,N_7377);
nand U10041 (N_10041,N_7326,N_8762);
nand U10042 (N_10042,N_7038,N_7183);
and U10043 (N_10043,N_8211,N_6647);
nand U10044 (N_10044,N_6711,N_8182);
nor U10045 (N_10045,N_8848,N_6324);
nand U10046 (N_10046,N_6685,N_9130);
or U10047 (N_10047,N_8694,N_6515);
nand U10048 (N_10048,N_6465,N_9292);
nand U10049 (N_10049,N_7281,N_8801);
or U10050 (N_10050,N_6369,N_7197);
nand U10051 (N_10051,N_7354,N_9267);
and U10052 (N_10052,N_7565,N_8370);
nor U10053 (N_10053,N_6257,N_8265);
nor U10054 (N_10054,N_9141,N_8791);
nand U10055 (N_10055,N_8825,N_7630);
nor U10056 (N_10056,N_7434,N_7693);
and U10057 (N_10057,N_6652,N_8919);
or U10058 (N_10058,N_6774,N_9371);
nor U10059 (N_10059,N_7052,N_7671);
nor U10060 (N_10060,N_6374,N_8803);
xnor U10061 (N_10061,N_8030,N_7433);
nand U10062 (N_10062,N_7721,N_8397);
and U10063 (N_10063,N_7756,N_7935);
nand U10064 (N_10064,N_8134,N_6703);
and U10065 (N_10065,N_7567,N_9165);
or U10066 (N_10066,N_7170,N_9324);
and U10067 (N_10067,N_7227,N_8839);
nor U10068 (N_10068,N_6979,N_7024);
and U10069 (N_10069,N_8236,N_6506);
or U10070 (N_10070,N_6542,N_6841);
nor U10071 (N_10071,N_7767,N_8205);
nor U10072 (N_10072,N_8695,N_8345);
nand U10073 (N_10073,N_8953,N_7673);
or U10074 (N_10074,N_7007,N_6483);
nor U10075 (N_10075,N_7111,N_8037);
and U10076 (N_10076,N_9361,N_7230);
and U10077 (N_10077,N_7887,N_8629);
and U10078 (N_10078,N_9091,N_8429);
and U10079 (N_10079,N_8452,N_8186);
or U10080 (N_10080,N_7240,N_9180);
nor U10081 (N_10081,N_6283,N_8746);
and U10082 (N_10082,N_6953,N_8100);
or U10083 (N_10083,N_8123,N_6999);
and U10084 (N_10084,N_7536,N_9317);
or U10085 (N_10085,N_8189,N_7188);
nand U10086 (N_10086,N_6532,N_6300);
nand U10087 (N_10087,N_6311,N_7317);
xor U10088 (N_10088,N_7231,N_9213);
nor U10089 (N_10089,N_8121,N_9046);
and U10090 (N_10090,N_9221,N_8416);
nand U10091 (N_10091,N_7932,N_6687);
or U10092 (N_10092,N_6576,N_9086);
nor U10093 (N_10093,N_6574,N_7554);
nand U10094 (N_10094,N_6591,N_7936);
nor U10095 (N_10095,N_8492,N_6446);
nand U10096 (N_10096,N_8139,N_8978);
and U10097 (N_10097,N_6835,N_8974);
and U10098 (N_10098,N_8515,N_8316);
nor U10099 (N_10099,N_9019,N_6989);
nor U10100 (N_10100,N_8025,N_8522);
nor U10101 (N_10101,N_7358,N_6364);
nor U10102 (N_10102,N_7521,N_7768);
and U10103 (N_10103,N_9295,N_8043);
nand U10104 (N_10104,N_7525,N_6272);
or U10105 (N_10105,N_6729,N_9037);
xnor U10106 (N_10106,N_6447,N_8407);
or U10107 (N_10107,N_9112,N_9188);
nor U10108 (N_10108,N_6681,N_7600);
and U10109 (N_10109,N_7349,N_6633);
nand U10110 (N_10110,N_6972,N_7679);
and U10111 (N_10111,N_8767,N_8331);
xnor U10112 (N_10112,N_7945,N_6569);
or U10113 (N_10113,N_7380,N_6458);
nor U10114 (N_10114,N_9303,N_9094);
nor U10115 (N_10115,N_8322,N_6925);
xor U10116 (N_10116,N_7366,N_7451);
nand U10117 (N_10117,N_7958,N_9186);
and U10118 (N_10118,N_8491,N_8729);
or U10119 (N_10119,N_6643,N_7268);
nor U10120 (N_10120,N_8704,N_8050);
or U10121 (N_10121,N_9333,N_6387);
and U10122 (N_10122,N_6965,N_6868);
nand U10123 (N_10123,N_8530,N_6827);
nor U10124 (N_10124,N_7259,N_7876);
nand U10125 (N_10125,N_8097,N_8219);
xor U10126 (N_10126,N_8432,N_8755);
nor U10127 (N_10127,N_8262,N_7923);
or U10128 (N_10128,N_8724,N_7707);
and U10129 (N_10129,N_8979,N_6780);
nor U10130 (N_10130,N_7237,N_8065);
and U10131 (N_10131,N_7888,N_8727);
and U10132 (N_10132,N_6281,N_6727);
nand U10133 (N_10133,N_8608,N_8168);
nor U10134 (N_10134,N_6912,N_8991);
nor U10135 (N_10135,N_6717,N_8745);
xnor U10136 (N_10136,N_8649,N_7172);
nor U10137 (N_10137,N_6353,N_8088);
or U10138 (N_10138,N_9132,N_8488);
xnor U10139 (N_10139,N_8339,N_8166);
or U10140 (N_10140,N_8141,N_6553);
and U10141 (N_10141,N_8274,N_7195);
and U10142 (N_10142,N_8020,N_6770);
or U10143 (N_10143,N_8266,N_6480);
and U10144 (N_10144,N_9136,N_6776);
or U10145 (N_10145,N_8237,N_9125);
or U10146 (N_10146,N_7000,N_6756);
xor U10147 (N_10147,N_6383,N_7301);
or U10148 (N_10148,N_8079,N_6442);
nand U10149 (N_10149,N_8309,N_8242);
nor U10150 (N_10150,N_9330,N_8373);
nor U10151 (N_10151,N_8789,N_6952);
nor U10152 (N_10152,N_8080,N_7423);
and U10153 (N_10153,N_7493,N_6785);
xnor U10154 (N_10154,N_7162,N_8882);
nor U10155 (N_10155,N_6358,N_6371);
nand U10156 (N_10156,N_8459,N_7367);
and U10157 (N_10157,N_6593,N_9356);
or U10158 (N_10158,N_8828,N_8248);
xnor U10159 (N_10159,N_7735,N_6445);
nand U10160 (N_10160,N_6331,N_7385);
or U10161 (N_10161,N_8009,N_6590);
nor U10162 (N_10162,N_8161,N_8959);
nand U10163 (N_10163,N_8200,N_8218);
and U10164 (N_10164,N_7207,N_6991);
and U10165 (N_10165,N_9078,N_9175);
nand U10166 (N_10166,N_7413,N_8024);
and U10167 (N_10167,N_7001,N_7551);
and U10168 (N_10168,N_7990,N_6757);
xor U10169 (N_10169,N_8315,N_7700);
and U10170 (N_10170,N_6336,N_6775);
and U10171 (N_10171,N_6976,N_9270);
or U10172 (N_10172,N_7334,N_8622);
nor U10173 (N_10173,N_9194,N_8821);
nand U10174 (N_10174,N_6885,N_8078);
nor U10175 (N_10175,N_7556,N_8809);
xnor U10176 (N_10176,N_7368,N_7258);
xnor U10177 (N_10177,N_7699,N_9075);
nand U10178 (N_10178,N_7018,N_8787);
nand U10179 (N_10179,N_8703,N_6554);
nor U10180 (N_10180,N_6759,N_8209);
nor U10181 (N_10181,N_9004,N_6917);
nand U10182 (N_10182,N_7743,N_8561);
nor U10183 (N_10183,N_7867,N_8418);
or U10184 (N_10184,N_7130,N_7121);
or U10185 (N_10185,N_8173,N_7149);
nor U10186 (N_10186,N_7942,N_7728);
xor U10187 (N_10187,N_7480,N_7578);
xor U10188 (N_10188,N_6747,N_9116);
or U10189 (N_10189,N_6594,N_7739);
nor U10190 (N_10190,N_7835,N_7786);
nand U10191 (N_10191,N_9143,N_8464);
nand U10192 (N_10192,N_7880,N_7304);
nor U10193 (N_10193,N_8618,N_7110);
nor U10194 (N_10194,N_6888,N_6734);
nand U10195 (N_10195,N_6941,N_7445);
and U10196 (N_10196,N_8841,N_9047);
and U10197 (N_10197,N_7027,N_7663);
or U10198 (N_10198,N_8034,N_7146);
nor U10199 (N_10199,N_6437,N_8812);
and U10200 (N_10200,N_7406,N_6486);
nor U10201 (N_10201,N_8941,N_8477);
and U10202 (N_10202,N_6609,N_7161);
or U10203 (N_10203,N_7114,N_7028);
nand U10204 (N_10204,N_7049,N_7180);
xnor U10205 (N_10205,N_8228,N_9051);
or U10206 (N_10206,N_9021,N_7825);
and U10207 (N_10207,N_8892,N_7513);
nand U10208 (N_10208,N_6560,N_8216);
nand U10209 (N_10209,N_6264,N_8130);
and U10210 (N_10210,N_7091,N_8777);
or U10211 (N_10211,N_8529,N_8665);
nor U10212 (N_10212,N_8047,N_7051);
and U10213 (N_10213,N_6528,N_9133);
nand U10214 (N_10214,N_6980,N_7144);
nor U10215 (N_10215,N_7979,N_8783);
xor U10216 (N_10216,N_6417,N_8964);
nand U10217 (N_10217,N_8263,N_7793);
xor U10218 (N_10218,N_8457,N_7312);
and U10219 (N_10219,N_6824,N_7941);
nand U10220 (N_10220,N_8115,N_7055);
nand U10221 (N_10221,N_6724,N_7568);
xor U10222 (N_10222,N_7277,N_7762);
and U10223 (N_10223,N_8150,N_8511);
nor U10224 (N_10224,N_7494,N_7347);
xor U10225 (N_10225,N_9104,N_6404);
or U10226 (N_10226,N_8400,N_9198);
nor U10227 (N_10227,N_6968,N_7809);
and U10228 (N_10228,N_6524,N_9122);
nand U10229 (N_10229,N_8797,N_7179);
nand U10230 (N_10230,N_6546,N_8826);
nor U10231 (N_10231,N_8131,N_8965);
nor U10232 (N_10232,N_9336,N_7190);
or U10233 (N_10233,N_8084,N_8988);
xor U10234 (N_10234,N_9033,N_7593);
nand U10235 (N_10235,N_8193,N_8657);
nand U10236 (N_10236,N_7238,N_8987);
nor U10237 (N_10237,N_7562,N_6872);
nor U10238 (N_10238,N_8192,N_7991);
or U10239 (N_10239,N_6892,N_8311);
or U10240 (N_10240,N_7763,N_8544);
nand U10241 (N_10241,N_8000,N_6731);
and U10242 (N_10242,N_8914,N_6250);
xnor U10243 (N_10243,N_7138,N_9214);
nand U10244 (N_10244,N_6400,N_9003);
and U10245 (N_10245,N_7948,N_7109);
or U10246 (N_10246,N_7714,N_7045);
and U10247 (N_10247,N_8871,N_8355);
nand U10248 (N_10248,N_9069,N_9304);
nor U10249 (N_10249,N_7336,N_8290);
or U10250 (N_10250,N_8798,N_6881);
nand U10251 (N_10251,N_8813,N_6798);
xor U10252 (N_10252,N_8693,N_6423);
or U10253 (N_10253,N_8027,N_7048);
or U10254 (N_10254,N_7350,N_7747);
or U10255 (N_10255,N_7939,N_8524);
nor U10256 (N_10256,N_7303,N_9306);
nand U10257 (N_10257,N_8834,N_6428);
nor U10258 (N_10258,N_8442,N_7503);
nand U10259 (N_10259,N_8880,N_6271);
xnor U10260 (N_10260,N_7982,N_8688);
or U10261 (N_10261,N_7967,N_6637);
nand U10262 (N_10262,N_8474,N_7004);
nand U10263 (N_10263,N_6351,N_7169);
nand U10264 (N_10264,N_7050,N_9101);
xnor U10265 (N_10265,N_8498,N_8213);
and U10266 (N_10266,N_9355,N_8118);
nand U10267 (N_10267,N_9328,N_6634);
or U10268 (N_10268,N_8751,N_8810);
nand U10269 (N_10269,N_8579,N_8481);
nand U10270 (N_10270,N_6425,N_6660);
nand U10271 (N_10271,N_7332,N_9216);
and U10272 (N_10272,N_7791,N_8363);
nor U10273 (N_10273,N_9039,N_8814);
and U10274 (N_10274,N_8164,N_6789);
xor U10275 (N_10275,N_8859,N_7120);
nand U10276 (N_10276,N_8918,N_7564);
and U10277 (N_10277,N_6555,N_6758);
or U10278 (N_10278,N_6873,N_9192);
nand U10279 (N_10279,N_8858,N_7212);
nand U10280 (N_10280,N_6304,N_8111);
nand U10281 (N_10281,N_6679,N_6548);
and U10282 (N_10282,N_7912,N_8041);
nand U10283 (N_10283,N_7165,N_8225);
or U10284 (N_10284,N_6863,N_7889);
or U10285 (N_10285,N_7906,N_9124);
and U10286 (N_10286,N_9262,N_7255);
and U10287 (N_10287,N_8354,N_6845);
nor U10288 (N_10288,N_9307,N_6343);
xnor U10289 (N_10289,N_9065,N_8753);
nor U10290 (N_10290,N_7894,N_7076);
xor U10291 (N_10291,N_7861,N_7492);
and U10292 (N_10292,N_8002,N_7119);
or U10293 (N_10293,N_8754,N_7145);
nand U10294 (N_10294,N_7708,N_6843);
nor U10295 (N_10295,N_6686,N_6610);
and U10296 (N_10296,N_9251,N_9279);
nand U10297 (N_10297,N_9106,N_7228);
nor U10298 (N_10298,N_8731,N_7860);
or U10299 (N_10299,N_6870,N_7520);
and U10300 (N_10300,N_7117,N_7057);
nor U10301 (N_10301,N_8583,N_8740);
and U10302 (N_10302,N_8444,N_8439);
and U10303 (N_10303,N_9072,N_8750);
nor U10304 (N_10304,N_7245,N_9058);
nand U10305 (N_10305,N_8868,N_9289);
nor U10306 (N_10306,N_7981,N_8348);
or U10307 (N_10307,N_8245,N_8969);
nor U10308 (N_10308,N_7920,N_7482);
nand U10309 (N_10309,N_8083,N_7849);
nand U10310 (N_10310,N_7158,N_6974);
or U10311 (N_10311,N_8431,N_8962);
or U10312 (N_10312,N_8656,N_8463);
nand U10313 (N_10313,N_6375,N_7646);
or U10314 (N_10314,N_6342,N_9238);
and U10315 (N_10315,N_6948,N_6489);
nor U10316 (N_10316,N_9224,N_8799);
xor U10317 (N_10317,N_7997,N_6765);
or U10318 (N_10318,N_8925,N_7950);
and U10319 (N_10319,N_9199,N_8636);
or U10320 (N_10320,N_8949,N_9023);
nand U10321 (N_10321,N_8261,N_9008);
and U10322 (N_10322,N_8641,N_8120);
nand U10323 (N_10323,N_7216,N_8605);
and U10324 (N_10324,N_7705,N_9120);
nand U10325 (N_10325,N_7807,N_8312);
nor U10326 (N_10326,N_6573,N_7497);
nand U10327 (N_10327,N_8365,N_6345);
nor U10328 (N_10328,N_8103,N_6766);
and U10329 (N_10329,N_7116,N_6419);
nand U10330 (N_10330,N_8697,N_7244);
nand U10331 (N_10331,N_7031,N_6267);
nor U10332 (N_10332,N_7017,N_8578);
nor U10333 (N_10333,N_8613,N_8521);
nand U10334 (N_10334,N_8388,N_9126);
and U10335 (N_10335,N_6849,N_6794);
and U10336 (N_10336,N_9139,N_9083);
and U10337 (N_10337,N_7864,N_8552);
and U10338 (N_10338,N_6541,N_7549);
nand U10339 (N_10339,N_9346,N_7777);
nand U10340 (N_10340,N_7816,N_9225);
nand U10341 (N_10341,N_8876,N_7189);
nand U10342 (N_10342,N_6564,N_6919);
xor U10343 (N_10343,N_8329,N_7037);
and U10344 (N_10344,N_7412,N_6411);
or U10345 (N_10345,N_9332,N_7966);
nand U10346 (N_10346,N_7737,N_6718);
or U10347 (N_10347,N_9185,N_7748);
nor U10348 (N_10348,N_6268,N_8602);
xor U10349 (N_10349,N_6301,N_6530);
and U10350 (N_10350,N_6262,N_6265);
or U10351 (N_10351,N_7851,N_7156);
and U10352 (N_10352,N_7160,N_6997);
and U10353 (N_10353,N_8904,N_7819);
and U10354 (N_10354,N_8571,N_7759);
or U10355 (N_10355,N_7946,N_7805);
or U10356 (N_10356,N_7236,N_7306);
nor U10357 (N_10357,N_7030,N_8152);
nand U10358 (N_10358,N_7285,N_6478);
and U10359 (N_10359,N_6683,N_7978);
xor U10360 (N_10360,N_6344,N_6279);
or U10361 (N_10361,N_8098,N_6286);
or U10362 (N_10362,N_8763,N_7327);
nand U10363 (N_10363,N_9128,N_6690);
nand U10364 (N_10364,N_9278,N_9263);
nor U10365 (N_10365,N_7314,N_8863);
nor U10366 (N_10366,N_7176,N_8157);
nand U10367 (N_10367,N_9089,N_7177);
nand U10368 (N_10368,N_7424,N_7224);
nor U10369 (N_10369,N_9273,N_8752);
and U10370 (N_10370,N_7702,N_9025);
or U10371 (N_10371,N_7818,N_6337);
nand U10372 (N_10372,N_9256,N_7641);
nand U10373 (N_10373,N_9031,N_7639);
xor U10374 (N_10374,N_9258,N_6939);
and U10375 (N_10375,N_8846,N_7261);
nor U10376 (N_10376,N_6986,N_7725);
or U10377 (N_10377,N_7951,N_8580);
nor U10378 (N_10378,N_8639,N_8893);
nand U10379 (N_10379,N_6462,N_8485);
and U10380 (N_10380,N_8775,N_8766);
and U10381 (N_10381,N_6474,N_8720);
or U10382 (N_10382,N_8865,N_7033);
nand U10383 (N_10383,N_7185,N_7071);
or U10384 (N_10384,N_6469,N_7295);
nor U10385 (N_10385,N_8465,N_8406);
nand U10386 (N_10386,N_6582,N_7013);
nand U10387 (N_10387,N_6716,N_6568);
nor U10388 (N_10388,N_7273,N_7400);
nor U10389 (N_10389,N_7425,N_9015);
and U10390 (N_10390,N_9041,N_6396);
nand U10391 (N_10391,N_9321,N_8946);
nand U10392 (N_10392,N_8067,N_8403);
and U10393 (N_10393,N_6950,N_8092);
xor U10394 (N_10394,N_8538,N_6436);
or U10395 (N_10395,N_9099,N_7469);
nor U10396 (N_10396,N_6750,N_8698);
and U10397 (N_10397,N_8129,N_8292);
nor U10398 (N_10398,N_6372,N_8562);
nor U10399 (N_10399,N_8558,N_9002);
nand U10400 (N_10400,N_9201,N_8721);
nor U10401 (N_10401,N_7857,N_8399);
or U10402 (N_10402,N_9149,N_8395);
and U10403 (N_10403,N_7579,N_9210);
nor U10404 (N_10404,N_8202,N_8295);
nor U10405 (N_10405,N_6433,N_7576);
xor U10406 (N_10406,N_8183,N_9365);
xor U10407 (N_10407,N_6333,N_9029);
or U10408 (N_10408,N_8862,N_9320);
or U10409 (N_10409,N_8926,N_6900);
nor U10410 (N_10410,N_8359,N_8895);
nor U10411 (N_10411,N_7294,N_8566);
nand U10412 (N_10412,N_9350,N_7833);
nor U10413 (N_10413,N_7163,N_6772);
nand U10414 (N_10414,N_7242,N_6378);
and U10415 (N_10415,N_8547,N_6955);
nand U10416 (N_10416,N_6988,N_6619);
and U10417 (N_10417,N_6390,N_8501);
xor U10418 (N_10418,N_8467,N_8396);
nand U10419 (N_10419,N_7775,N_8886);
or U10420 (N_10420,N_9088,N_8659);
xnor U10421 (N_10421,N_8958,N_8917);
or U10422 (N_10422,N_7302,N_7872);
or U10423 (N_10423,N_7352,N_6741);
nor U10424 (N_10424,N_9050,N_8915);
nand U10425 (N_10425,N_6625,N_6882);
and U10426 (N_10426,N_8844,N_7687);
or U10427 (N_10427,N_7969,N_6688);
nand U10428 (N_10428,N_9090,N_6992);
xnor U10429 (N_10429,N_8135,N_7908);
nor U10430 (N_10430,N_8542,N_7755);
nand U10431 (N_10431,N_6494,N_6551);
or U10432 (N_10432,N_6673,N_9261);
and U10433 (N_10433,N_7540,N_6908);
and U10434 (N_10434,N_8375,N_7771);
nand U10435 (N_10435,N_7353,N_6595);
nand U10436 (N_10436,N_7789,N_7315);
xnor U10437 (N_10437,N_6806,N_7986);
or U10438 (N_10438,N_7283,N_6805);
nor U10439 (N_10439,N_8807,N_8765);
nor U10440 (N_10440,N_6598,N_8201);
and U10441 (N_10441,N_8493,N_8633);
xor U10442 (N_10442,N_7514,N_8942);
nor U10443 (N_10443,N_8796,N_8678);
or U10444 (N_10444,N_7566,N_8433);
nand U10445 (N_10445,N_8394,N_9187);
or U10446 (N_10446,N_6495,N_8911);
and U10447 (N_10447,N_6649,N_7486);
and U10448 (N_10448,N_6719,N_8408);
nand U10449 (N_10449,N_7274,N_7476);
xnor U10450 (N_10450,N_9113,N_6405);
nand U10451 (N_10451,N_6662,N_8854);
nand U10452 (N_10452,N_6503,N_6725);
nand U10453 (N_10453,N_8781,N_7617);
nor U10454 (N_10454,N_8747,N_6699);
or U10455 (N_10455,N_8916,N_9137);
or U10456 (N_10456,N_6602,N_9115);
nand U10457 (N_10457,N_7297,N_7571);
and U10458 (N_10458,N_9318,N_9218);
nor U10459 (N_10459,N_7616,N_8153);
or U10460 (N_10460,N_6459,N_9363);
and U10461 (N_10461,N_8421,N_8996);
nand U10462 (N_10462,N_6608,N_8093);
nand U10463 (N_10463,N_7054,N_6360);
nor U10464 (N_10464,N_7918,N_7559);
or U10465 (N_10465,N_9048,N_7661);
nor U10466 (N_10466,N_7961,N_6496);
xor U10467 (N_10467,N_8383,N_9359);
or U10468 (N_10468,N_7485,N_8430);
nor U10469 (N_10469,N_7323,N_6937);
nor U10470 (N_10470,N_7624,N_6513);
or U10471 (N_10471,N_8545,N_7284);
and U10472 (N_10472,N_7217,N_9140);
or U10473 (N_10473,N_8983,N_7930);
and U10474 (N_10474,N_6930,N_7794);
or U10475 (N_10475,N_8454,N_7447);
and U10476 (N_10476,N_6927,N_7977);
nor U10477 (N_10477,N_8960,N_7428);
nand U10478 (N_10478,N_7319,N_7649);
and U10479 (N_10479,N_8994,N_7208);
or U10480 (N_10480,N_8646,N_6697);
nor U10481 (N_10481,N_6791,N_7680);
nand U10482 (N_10482,N_7372,N_9067);
or U10483 (N_10483,N_8620,N_9070);
nand U10484 (N_10484,N_8948,N_9068);
and U10485 (N_10485,N_8785,N_8091);
nand U10486 (N_10486,N_6466,N_7010);
xnor U10487 (N_10487,N_9243,N_8072);
and U10488 (N_10488,N_6395,N_8832);
xor U10489 (N_10489,N_7591,N_7416);
and U10490 (N_10490,N_8377,N_6839);
nand U10491 (N_10491,N_7318,N_7538);
and U10492 (N_10492,N_8317,N_7804);
nor U10493 (N_10493,N_6571,N_9035);
or U10494 (N_10494,N_7826,N_8591);
and U10495 (N_10495,N_7065,N_6810);
nand U10496 (N_10496,N_8055,N_8716);
nor U10497 (N_10497,N_8823,N_6665);
nand U10498 (N_10498,N_7770,N_8028);
and U10499 (N_10499,N_9286,N_8935);
or U10500 (N_10500,N_7965,N_6493);
or U10501 (N_10501,N_7654,N_6306);
and U10502 (N_10502,N_6745,N_6701);
xor U10503 (N_10503,N_7219,N_9158);
nor U10504 (N_10504,N_7198,N_8171);
or U10505 (N_10505,N_9314,N_8045);
nand U10506 (N_10506,N_7443,N_8759);
nor U10507 (N_10507,N_6754,N_7462);
nand U10508 (N_10508,N_7698,N_7457);
and U10509 (N_10509,N_6797,N_8318);
nand U10510 (N_10510,N_8690,N_7393);
and U10511 (N_10511,N_6580,N_8374);
nand U10512 (N_10512,N_8963,N_7572);
or U10513 (N_10513,N_8269,N_7994);
xnor U10514 (N_10514,N_8222,N_8627);
or U10515 (N_10515,N_7139,N_7409);
or U10516 (N_10516,N_7399,N_8232);
nand U10517 (N_10517,N_7491,N_8175);
nor U10518 (N_10518,N_6983,N_9374);
xor U10519 (N_10519,N_9230,N_8543);
nand U10520 (N_10520,N_6894,N_6994);
nor U10521 (N_10521,N_6680,N_7288);
nand U10522 (N_10522,N_7015,N_8238);
nor U10523 (N_10523,N_7656,N_7764);
or U10524 (N_10524,N_7178,N_8908);
and U10525 (N_10525,N_8675,N_8035);
and U10526 (N_10526,N_8686,N_6415);
or U10527 (N_10527,N_8448,N_7904);
xnor U10528 (N_10528,N_7829,N_7620);
and U10529 (N_10529,N_6629,N_8874);
xnor U10530 (N_10530,N_7757,N_8177);
and U10531 (N_10531,N_8528,N_6659);
nand U10532 (N_10532,N_8325,N_6857);
nor U10533 (N_10533,N_6451,N_6529);
or U10534 (N_10534,N_7166,N_7272);
and U10535 (N_10535,N_9323,N_8472);
xnor U10536 (N_10536,N_6339,N_6409);
nand U10537 (N_10537,N_8301,N_6708);
nor U10538 (N_10538,N_7518,N_6705);
nand U10539 (N_10539,N_7801,N_8870);
or U10540 (N_10540,N_9290,N_6752);
and U10541 (N_10541,N_7760,N_6606);
xor U10542 (N_10542,N_9300,N_7135);
and U10543 (N_10543,N_8999,N_7411);
and U10544 (N_10544,N_6293,N_8788);
and U10545 (N_10545,N_6763,N_6829);
and U10546 (N_10546,N_6261,N_7147);
nor U10547 (N_10547,N_8381,N_6639);
nor U10548 (N_10548,N_8140,N_8029);
nor U10549 (N_10549,N_7911,N_8095);
and U10550 (N_10550,N_7541,N_7817);
and U10551 (N_10551,N_8163,N_8609);
nor U10552 (N_10552,N_8980,N_8808);
and U10553 (N_10553,N_9077,N_6738);
and U10554 (N_10554,N_7020,N_8178);
or U10555 (N_10555,N_8172,N_6276);
and U10556 (N_10556,N_6332,N_7836);
and U10557 (N_10557,N_7293,N_7333);
nand U10558 (N_10558,N_7449,N_8090);
nor U10559 (N_10559,N_6787,N_9084);
nand U10560 (N_10560,N_6429,N_7131);
nand U10561 (N_10561,N_7328,N_6277);
or U10562 (N_10562,N_7431,N_7148);
nor U10563 (N_10563,N_8577,N_9285);
or U10564 (N_10564,N_9135,N_7544);
xor U10565 (N_10565,N_7286,N_7627);
nand U10566 (N_10566,N_7608,N_9134);
and U10567 (N_10567,N_8257,N_7381);
nand U10568 (N_10568,N_9026,N_7808);
or U10569 (N_10569,N_7552,N_6656);
or U10570 (N_10570,N_6531,N_6809);
and U10571 (N_10571,N_6929,N_6864);
or U10572 (N_10572,N_6702,N_8903);
nand U10573 (N_10573,N_9010,N_7254);
xnor U10574 (N_10574,N_8786,N_8489);
nand U10575 (N_10575,N_7232,N_8555);
nand U10576 (N_10576,N_9150,N_6382);
nor U10577 (N_10577,N_8509,N_9335);
nand U10578 (N_10578,N_7601,N_9066);
and U10579 (N_10579,N_7774,N_7730);
or U10580 (N_10580,N_9255,N_6454);
xor U10581 (N_10581,N_8744,N_7669);
or U10582 (N_10582,N_7427,N_7716);
nor U10583 (N_10583,N_7436,N_6674);
xor U10584 (N_10584,N_7586,N_8099);
nor U10585 (N_10585,N_7779,N_6833);
xor U10586 (N_10586,N_7931,N_6784);
and U10587 (N_10587,N_6318,N_6453);
nand U10588 (N_10588,N_7519,N_7753);
or U10589 (N_10589,N_7523,N_9131);
nor U10590 (N_10590,N_8535,N_6648);
or U10591 (N_10591,N_9038,N_7338);
nand U10592 (N_10592,N_7815,N_7063);
or U10593 (N_10593,N_7896,N_7191);
nor U10594 (N_10594,N_6818,N_7090);
nor U10595 (N_10595,N_9096,N_6385);
or U10596 (N_10596,N_8527,N_6970);
nor U10597 (N_10597,N_8156,N_7732);
nand U10598 (N_10598,N_6733,N_8873);
or U10599 (N_10599,N_8414,N_7321);
or U10600 (N_10600,N_7547,N_6706);
or U10601 (N_10601,N_8026,N_6801);
nand U10602 (N_10602,N_8945,N_9367);
and U10603 (N_10603,N_7898,N_8701);
and U10604 (N_10604,N_8573,N_6523);
or U10605 (N_10605,N_7683,N_8784);
and U10606 (N_10606,N_7604,N_6779);
nor U10607 (N_10607,N_8715,N_6507);
or U10608 (N_10608,N_7320,N_6934);
nand U10609 (N_10609,N_6607,N_8203);
and U10610 (N_10610,N_8967,N_7173);
nor U10611 (N_10611,N_7871,N_6769);
xor U10612 (N_10612,N_6722,N_9007);
or U10613 (N_10613,N_6520,N_8143);
and U10614 (N_10614,N_7724,N_8564);
and U10615 (N_10615,N_8144,N_6945);
nand U10616 (N_10616,N_7061,N_8063);
nand U10617 (N_10617,N_6552,N_8145);
xnor U10618 (N_10618,N_9036,N_7081);
nor U10619 (N_10619,N_8158,N_8723);
and U10620 (N_10620,N_8603,N_7587);
nor U10621 (N_10621,N_7351,N_7623);
nor U10622 (N_10622,N_8393,N_6561);
nand U10623 (N_10623,N_8113,N_6485);
or U10624 (N_10624,N_7954,N_7960);
xor U10625 (N_10625,N_7410,N_6740);
nor U10626 (N_10626,N_8278,N_9108);
nor U10627 (N_10627,N_8007,N_7599);
nor U10628 (N_10628,N_7247,N_8540);
and U10629 (N_10629,N_7688,N_8361);
nand U10630 (N_10630,N_8951,N_6501);
or U10631 (N_10631,N_8119,N_7475);
nor U10632 (N_10632,N_8247,N_9151);
xor U10633 (N_10633,N_9081,N_7355);
nand U10634 (N_10634,N_6365,N_6735);
or U10635 (N_10635,N_8367,N_8392);
nand U10636 (N_10636,N_8513,N_8845);
nor U10637 (N_10637,N_6736,N_8726);
nor U10638 (N_10638,N_8867,N_6587);
xor U10639 (N_10639,N_8102,N_7798);
nor U10640 (N_10640,N_7907,N_6672);
nand U10641 (N_10641,N_8204,N_7430);
or U10642 (N_10642,N_9313,N_8947);
nand U10643 (N_10643,N_8671,N_7388);
and U10644 (N_10644,N_7758,N_7718);
xnor U10645 (N_10645,N_8051,N_7458);
xnor U10646 (N_10646,N_8681,N_6601);
nor U10647 (N_10647,N_8966,N_8961);
or U10648 (N_10648,N_6391,N_8468);
xnor U10649 (N_10649,N_7343,N_9052);
and U10650 (N_10650,N_6412,N_7305);
xor U10651 (N_10651,N_7652,N_9277);
and U10652 (N_10652,N_6931,N_7348);
nand U10653 (N_10653,N_7395,N_7921);
nor U10654 (N_10654,N_9040,N_7548);
and U10655 (N_10655,N_7913,N_9102);
xnor U10656 (N_10656,N_8005,N_8306);
and U10657 (N_10657,N_8713,N_6947);
and U10658 (N_10658,N_7070,N_7418);
or U10659 (N_10659,N_7878,N_6905);
and U10660 (N_10660,N_8709,N_8712);
nand U10661 (N_10661,N_6910,N_8856);
or U10662 (N_10662,N_6712,N_7501);
and U10663 (N_10663,N_8108,N_8384);
xor U10664 (N_10664,N_8341,N_7983);
xor U10665 (N_10665,N_8369,N_7752);
xnor U10666 (N_10666,N_8413,N_8473);
or U10667 (N_10667,N_8977,N_6760);
nand U10668 (N_10668,N_6959,N_8054);
nand U10669 (N_10669,N_8940,N_8074);
nor U10670 (N_10670,N_8332,N_9063);
nand U10671 (N_10671,N_9056,N_9342);
nor U10672 (N_10672,N_7382,N_7901);
xnor U10673 (N_10673,N_9327,N_6350);
or U10674 (N_10674,N_7947,N_6893);
or U10675 (N_10675,N_8450,N_7083);
and U10676 (N_10676,N_6622,N_6692);
and U10677 (N_10677,N_6352,N_9352);
nor U10678 (N_10678,N_6778,N_7112);
and U10679 (N_10679,N_7330,N_7248);
nand U10680 (N_10680,N_7782,N_8502);
or U10681 (N_10681,N_8249,N_6310);
nor U10682 (N_10682,N_6822,N_8851);
or U10683 (N_10683,N_8441,N_6380);
nand U10684 (N_10684,N_9173,N_8706);
and U10685 (N_10685,N_8031,N_8303);
or U10686 (N_10686,N_9265,N_8229);
nor U10687 (N_10687,N_8124,N_7157);
and U10688 (N_10688,N_6452,N_7832);
or U10689 (N_10689,N_9244,N_7582);
nor U10690 (N_10690,N_7291,N_7984);
xnor U10691 (N_10691,N_8415,N_7814);
nand U10692 (N_10692,N_7697,N_7796);
or U10693 (N_10693,N_8973,N_8565);
or U10694 (N_10694,N_6799,N_8059);
nor U10695 (N_10695,N_8523,N_6525);
nand U10696 (N_10696,N_8338,N_7374);
or U10697 (N_10697,N_8606,N_8922);
and U10698 (N_10698,N_8651,N_9220);
nand U10699 (N_10699,N_7108,N_6676);
or U10700 (N_10700,N_7322,N_7437);
xnor U10701 (N_10701,N_7435,N_6468);
nand U10702 (N_10702,N_8281,N_8270);
and U10703 (N_10703,N_9217,N_8142);
nor U10704 (N_10704,N_8283,N_8256);
and U10705 (N_10705,N_7772,N_8267);
or U10706 (N_10706,N_8022,N_7588);
nand U10707 (N_10707,N_6253,N_6898);
nor U10708 (N_10708,N_8849,N_8233);
nand U10709 (N_10709,N_7167,N_8360);
and U10710 (N_10710,N_6922,N_6831);
nor U10711 (N_10711,N_8405,N_7044);
nand U10712 (N_10712,N_8042,N_7452);
and U10713 (N_10713,N_9011,N_6815);
nor U10714 (N_10714,N_6761,N_7215);
nand U10715 (N_10715,N_6613,N_6366);
xor U10716 (N_10716,N_7101,N_8207);
or U10717 (N_10717,N_9360,N_8685);
nand U10718 (N_10718,N_6954,N_6490);
and U10719 (N_10719,N_9271,N_8081);
or U10720 (N_10720,N_7831,N_7847);
nor U10721 (N_10721,N_8674,N_7035);
or U10722 (N_10722,N_8323,N_6479);
nor U10723 (N_10723,N_6816,N_9302);
nand U10724 (N_10724,N_7067,N_7474);
nand U10725 (N_10725,N_7792,N_8259);
and U10726 (N_10726,N_7532,N_8730);
or U10727 (N_10727,N_8993,N_9053);
nor U10728 (N_10728,N_6432,N_6753);
nor U10729 (N_10729,N_6450,N_6936);
nand U10730 (N_10730,N_7922,N_7444);
or U10731 (N_10731,N_9358,N_9197);
and U10732 (N_10732,N_9349,N_7672);
and U10733 (N_10733,N_8997,N_6407);
or U10734 (N_10734,N_6577,N_8462);
nand U10735 (N_10735,N_7194,N_8199);
or U10736 (N_10736,N_6749,N_7866);
xnor U10737 (N_10737,N_8440,N_9236);
or U10738 (N_10738,N_8268,N_6329);
and U10739 (N_10739,N_7613,N_6316);
or U10740 (N_10740,N_8837,N_9315);
nor U10741 (N_10741,N_8559,N_8525);
nor U10742 (N_10742,N_6764,N_7365);
and U10743 (N_10743,N_8075,N_8277);
and U10744 (N_10744,N_7642,N_8928);
or U10745 (N_10745,N_8351,N_6408);
or U10746 (N_10746,N_9309,N_7453);
or U10747 (N_10747,N_7883,N_6533);
and U10748 (N_10748,N_7660,N_8722);
xor U10749 (N_10749,N_6266,N_7196);
xor U10750 (N_10750,N_6370,N_8040);
nor U10751 (N_10751,N_9156,N_8975);
xor U10752 (N_10752,N_9211,N_7650);
xnor U10753 (N_10753,N_7592,N_8223);
nand U10754 (N_10754,N_7066,N_8330);
and U10755 (N_10755,N_8104,N_6508);
nor U10756 (N_10756,N_7890,N_9338);
or U10757 (N_10757,N_9057,N_7685);
and U10758 (N_10758,N_9114,N_9274);
or U10759 (N_10759,N_7780,N_8592);
nor U10760 (N_10760,N_8324,N_6287);
or U10761 (N_10761,N_8148,N_8732);
xor U10762 (N_10762,N_8584,N_7740);
xor U10763 (N_10763,N_7379,N_7606);
nand U10764 (N_10764,N_6275,N_8417);
and U10765 (N_10765,N_8905,N_9269);
and U10766 (N_10766,N_8217,N_6792);
nor U10767 (N_10767,N_7014,N_7602);
xor U10768 (N_10768,N_6334,N_7696);
and U10769 (N_10769,N_8282,N_8897);
xor U10770 (N_10770,N_6290,N_7140);
nor U10771 (N_10771,N_8496,N_7865);
or U10772 (N_10772,N_8272,N_8572);
and U10773 (N_10773,N_9223,N_7296);
or U10774 (N_10774,N_8692,N_7609);
xor U10775 (N_10775,N_7882,N_9171);
or U10776 (N_10776,N_7996,N_6946);
nand U10777 (N_10777,N_9208,N_6487);
and U10778 (N_10778,N_6886,N_8036);
and U10779 (N_10779,N_7456,N_6455);
nand U10780 (N_10780,N_9275,N_7674);
nor U10781 (N_10781,N_7199,N_8739);
or U10782 (N_10782,N_6422,N_9193);
or U10783 (N_10783,N_8423,N_6768);
nor U10784 (N_10784,N_6742,N_7533);
xnor U10785 (N_10785,N_8260,N_7269);
nor U10786 (N_10786,N_6971,N_9080);
nor U10787 (N_10787,N_7681,N_8251);
nand U10788 (N_10788,N_7099,N_6696);
and U10789 (N_10789,N_6867,N_7827);
xnor U10790 (N_10790,N_7667,N_6918);
nand U10791 (N_10791,N_9082,N_7506);
xnor U10792 (N_10792,N_6896,N_8989);
and U10793 (N_10793,N_7785,N_6355);
nand U10794 (N_10794,N_7357,N_8536);
or U10795 (N_10795,N_6628,N_6398);
or U10796 (N_10796,N_6297,N_8021);
nor U10797 (N_10797,N_6335,N_6865);
and U10798 (N_10798,N_6823,N_8008);
nand U10799 (N_10799,N_7363,N_8955);
or U10800 (N_10800,N_7460,N_8748);
nand U10801 (N_10801,N_7490,N_7006);
or U10802 (N_10802,N_6357,N_7396);
and U10803 (N_10803,N_8349,N_7640);
nand U10804 (N_10804,N_6516,N_8015);
nor U10805 (N_10805,N_7884,N_9209);
and U10806 (N_10806,N_6502,N_8333);
nand U10807 (N_10807,N_6263,N_7279);
nand U10808 (N_10808,N_7256,N_8039);
xor U10809 (N_10809,N_8056,N_8679);
or U10810 (N_10810,N_7331,N_7126);
nand U10811 (N_10811,N_7056,N_6320);
or U10812 (N_10812,N_8291,N_6330);
nor U10813 (N_10813,N_7729,N_7543);
nor U10814 (N_10814,N_6481,N_7498);
nor U10815 (N_10815,N_6471,N_7657);
nor U10816 (N_10816,N_6562,N_6535);
nand U10817 (N_10817,N_7974,N_7684);
or U10818 (N_10818,N_6832,N_8568);
nand U10819 (N_10819,N_7340,N_6721);
or U10820 (N_10820,N_6431,N_6536);
or U10821 (N_10821,N_8776,N_7342);
nand U10822 (N_10822,N_6895,N_8357);
or U10823 (N_10823,N_6259,N_9200);
nor U10824 (N_10824,N_7622,N_8795);
nor U10825 (N_10825,N_7637,N_6684);
or U10826 (N_10826,N_7455,N_7706);
or U10827 (N_10827,N_8006,N_7975);
nand U10828 (N_10828,N_8443,N_7635);
xnor U10829 (N_10829,N_6627,N_9138);
nor U10830 (N_10830,N_9087,N_7125);
and U10831 (N_10831,N_8117,N_8133);
or U10832 (N_10832,N_6707,N_8146);
or U10833 (N_10833,N_8447,N_7859);
nor U10834 (N_10834,N_7632,N_7886);
xor U10835 (N_10835,N_9222,N_8176);
or U10836 (N_10836,N_6658,N_6788);
and U10837 (N_10837,N_6700,N_6563);
or U10838 (N_10838,N_6504,N_8985);
nor U10839 (N_10839,N_8594,N_6667);
xnor U10840 (N_10840,N_9206,N_9121);
or U10841 (N_10841,N_6998,N_7855);
nand U10842 (N_10842,N_8335,N_9281);
nand U10843 (N_10843,N_6565,N_6484);
and U10844 (N_10844,N_7243,N_6618);
nor U10845 (N_10845,N_6611,N_7479);
nor U10846 (N_10846,N_7766,N_6817);
or U10847 (N_10847,N_9322,N_6456);
nor U10848 (N_10848,N_6621,N_7870);
or U10849 (N_10849,N_6850,N_7087);
or U10850 (N_10850,N_8714,N_7844);
nand U10851 (N_10851,N_7940,N_8599);
nand U10852 (N_10852,N_6549,N_7999);
or U10853 (N_10853,N_7773,N_8640);
and U10854 (N_10854,N_8927,N_6570);
nor U10855 (N_10855,N_8085,N_7308);
and U10856 (N_10856,N_7414,N_7387);
nor U10857 (N_10857,N_6376,N_8596);
or U10858 (N_10858,N_8046,N_6819);
nor U10859 (N_10859,N_6473,N_7402);
nor U10860 (N_10860,N_8520,N_8013);
and U10861 (N_10861,N_7047,N_8614);
or U10862 (N_10862,N_7422,N_8276);
and U10863 (N_10863,N_7124,N_7266);
xnor U10864 (N_10864,N_8683,N_6675);
or U10865 (N_10865,N_7715,N_6386);
and U10866 (N_10866,N_6499,N_9183);
or U10867 (N_10867,N_8898,N_8076);
or U10868 (N_10868,N_8677,N_8981);
nand U10869 (N_10869,N_8149,N_8082);
nand U10870 (N_10870,N_7869,N_7845);
nand U10871 (N_10871,N_7128,N_8906);
nor U10872 (N_10872,N_8299,N_8847);
nor U10873 (N_10873,N_9013,N_6305);
and U10874 (N_10874,N_8089,N_7233);
nand U10875 (N_10875,N_6943,N_9353);
or U10876 (N_10876,N_8532,N_6389);
nand U10877 (N_10877,N_8557,N_9347);
xor U10878 (N_10878,N_6836,N_7710);
or U10879 (N_10879,N_8230,N_6326);
nor U10880 (N_10880,N_8741,N_9059);
and U10881 (N_10881,N_6444,N_6438);
nor U10882 (N_10882,N_7856,N_9107);
nand U10883 (N_10883,N_9060,N_6558);
nor U10884 (N_10884,N_8221,N_6603);
and U10885 (N_10885,N_7378,N_8206);
nor U10886 (N_10886,N_8998,N_7765);
or U10887 (N_10887,N_8422,N_8643);
and U10888 (N_10888,N_7731,N_8518);
or U10889 (N_10889,N_7953,N_6978);
and U10890 (N_10890,N_6859,N_7985);
or U10891 (N_10891,N_8346,N_6638);
nand U10892 (N_10892,N_7929,N_7003);
or U10893 (N_10893,N_7659,N_8469);
or U10894 (N_10894,N_7505,N_6260);
or U10895 (N_10895,N_8214,N_6793);
or U10896 (N_10896,N_8487,N_6645);
nand U10897 (N_10897,N_7717,N_7005);
nor U10898 (N_10898,N_6349,N_9103);
nor U10899 (N_10899,N_6282,N_7089);
nand U10900 (N_10900,N_6982,N_6664);
and U10901 (N_10901,N_7478,N_7557);
and U10902 (N_10902,N_8500,N_8901);
nor U10903 (N_10903,N_8017,N_8307);
nand U10904 (N_10904,N_9247,N_6834);
nor U10905 (N_10905,N_8497,N_7838);
xnor U10906 (N_10906,N_6933,N_6321);
nand U10907 (N_10907,N_7916,N_8061);
or U10908 (N_10908,N_7129,N_9311);
nand U10909 (N_10909,N_9169,N_8453);
nand U10910 (N_10910,N_8756,N_6909);
nor U10911 (N_10911,N_7094,N_6256);
nor U10912 (N_10912,N_6544,N_8011);
nand U10913 (N_10913,N_8326,N_6583);
nand U10914 (N_10914,N_8526,N_9344);
nand U10915 (N_10915,N_8476,N_7373);
and U10916 (N_10916,N_8840,N_9152);
nor U10917 (N_10917,N_7584,N_7830);
nor U10918 (N_10918,N_8484,N_6254);
and U10919 (N_10919,N_9232,N_8366);
nand U10920 (N_10920,N_6296,N_9111);
nand U10921 (N_10921,N_6292,N_9240);
and U10922 (N_10922,N_8438,N_6288);
or U10923 (N_10923,N_6720,N_8934);
and U10924 (N_10924,N_8280,N_7820);
nor U10925 (N_10925,N_8615,N_6869);
nor U10926 (N_10926,N_6522,N_6926);
nand U10927 (N_10927,N_8190,N_8802);
nor U10928 (N_10928,N_8136,N_8696);
nor U10929 (N_10929,N_9298,N_7186);
nor U10930 (N_10930,N_8610,N_8541);
and U10931 (N_10931,N_8337,N_8822);
nand U10932 (N_10932,N_7658,N_9326);
xor U10933 (N_10933,N_8792,N_7016);
nand U10934 (N_10934,N_8711,N_7726);
and U10935 (N_10935,N_7834,N_8128);
and U10936 (N_10936,N_7106,N_6463);
nand U10937 (N_10937,N_9228,N_7156);
nor U10938 (N_10938,N_8242,N_7058);
nand U10939 (N_10939,N_6730,N_9075);
nand U10940 (N_10940,N_7719,N_8057);
and U10941 (N_10941,N_8490,N_8473);
and U10942 (N_10942,N_8852,N_7481);
or U10943 (N_10943,N_7079,N_7154);
and U10944 (N_10944,N_7268,N_8244);
or U10945 (N_10945,N_8632,N_6430);
or U10946 (N_10946,N_6374,N_9132);
nor U10947 (N_10947,N_6955,N_8441);
nor U10948 (N_10948,N_7312,N_8312);
or U10949 (N_10949,N_7586,N_6803);
xnor U10950 (N_10950,N_8049,N_7661);
nand U10951 (N_10951,N_8007,N_8717);
and U10952 (N_10952,N_7578,N_6491);
and U10953 (N_10953,N_6831,N_9338);
and U10954 (N_10954,N_8100,N_6570);
or U10955 (N_10955,N_9295,N_6479);
or U10956 (N_10956,N_8283,N_8091);
or U10957 (N_10957,N_8517,N_7760);
xor U10958 (N_10958,N_9179,N_7847);
xor U10959 (N_10959,N_8616,N_8124);
and U10960 (N_10960,N_8844,N_6964);
and U10961 (N_10961,N_8197,N_8152);
xnor U10962 (N_10962,N_8954,N_8876);
nand U10963 (N_10963,N_9196,N_6762);
nor U10964 (N_10964,N_8931,N_9116);
nor U10965 (N_10965,N_8722,N_7150);
and U10966 (N_10966,N_7672,N_8053);
nand U10967 (N_10967,N_8749,N_6707);
or U10968 (N_10968,N_6805,N_7125);
xor U10969 (N_10969,N_9255,N_9078);
xnor U10970 (N_10970,N_7234,N_6840);
nand U10971 (N_10971,N_6824,N_8530);
nand U10972 (N_10972,N_7656,N_7884);
and U10973 (N_10973,N_8219,N_8112);
or U10974 (N_10974,N_8441,N_7566);
and U10975 (N_10975,N_7122,N_8001);
xnor U10976 (N_10976,N_7556,N_6697);
or U10977 (N_10977,N_8217,N_6683);
and U10978 (N_10978,N_7313,N_6745);
nor U10979 (N_10979,N_8708,N_6510);
nand U10980 (N_10980,N_7670,N_8768);
or U10981 (N_10981,N_8803,N_6684);
nor U10982 (N_10982,N_6654,N_7178);
xnor U10983 (N_10983,N_7041,N_8882);
nand U10984 (N_10984,N_6814,N_8588);
xor U10985 (N_10985,N_8217,N_7048);
and U10986 (N_10986,N_6753,N_8026);
xor U10987 (N_10987,N_7824,N_9186);
and U10988 (N_10988,N_6648,N_9263);
or U10989 (N_10989,N_8196,N_6364);
nor U10990 (N_10990,N_7074,N_6350);
and U10991 (N_10991,N_6512,N_6750);
or U10992 (N_10992,N_7665,N_6586);
and U10993 (N_10993,N_8551,N_9270);
nor U10994 (N_10994,N_6254,N_7420);
nand U10995 (N_10995,N_7490,N_6535);
or U10996 (N_10996,N_7005,N_7539);
nand U10997 (N_10997,N_9153,N_7311);
or U10998 (N_10998,N_8532,N_8463);
nor U10999 (N_10999,N_7053,N_7974);
nor U11000 (N_11000,N_6452,N_7238);
and U11001 (N_11001,N_9176,N_8711);
xor U11002 (N_11002,N_8901,N_6288);
nand U11003 (N_11003,N_9073,N_8614);
nand U11004 (N_11004,N_6624,N_7421);
nand U11005 (N_11005,N_6778,N_8845);
or U11006 (N_11006,N_9020,N_6643);
nor U11007 (N_11007,N_7889,N_8073);
nand U11008 (N_11008,N_7570,N_6526);
and U11009 (N_11009,N_9215,N_7872);
or U11010 (N_11010,N_7202,N_6581);
xor U11011 (N_11011,N_7707,N_7848);
nand U11012 (N_11012,N_6578,N_6996);
and U11013 (N_11013,N_6864,N_7442);
nor U11014 (N_11014,N_6847,N_7648);
and U11015 (N_11015,N_8181,N_9058);
nand U11016 (N_11016,N_8288,N_7398);
or U11017 (N_11017,N_8739,N_7508);
nor U11018 (N_11018,N_7458,N_8204);
nand U11019 (N_11019,N_8934,N_7025);
nor U11020 (N_11020,N_7627,N_6754);
or U11021 (N_11021,N_7359,N_7210);
nand U11022 (N_11022,N_7346,N_9051);
nand U11023 (N_11023,N_7395,N_8558);
or U11024 (N_11024,N_6644,N_7547);
xnor U11025 (N_11025,N_9172,N_8155);
nor U11026 (N_11026,N_7306,N_6542);
and U11027 (N_11027,N_8443,N_7823);
nor U11028 (N_11028,N_7852,N_8786);
and U11029 (N_11029,N_7202,N_8087);
and U11030 (N_11030,N_8693,N_8326);
and U11031 (N_11031,N_7508,N_7024);
or U11032 (N_11032,N_8797,N_8358);
xnor U11033 (N_11033,N_7655,N_7739);
and U11034 (N_11034,N_9088,N_9348);
or U11035 (N_11035,N_8808,N_7997);
and U11036 (N_11036,N_8097,N_7431);
or U11037 (N_11037,N_7567,N_7703);
xnor U11038 (N_11038,N_7339,N_8404);
and U11039 (N_11039,N_7561,N_8734);
xnor U11040 (N_11040,N_6791,N_6755);
or U11041 (N_11041,N_8115,N_8873);
or U11042 (N_11042,N_8800,N_8851);
nor U11043 (N_11043,N_7675,N_8675);
or U11044 (N_11044,N_9159,N_8420);
or U11045 (N_11045,N_7929,N_8872);
or U11046 (N_11046,N_9310,N_7392);
or U11047 (N_11047,N_8787,N_8236);
or U11048 (N_11048,N_8044,N_6317);
and U11049 (N_11049,N_8552,N_8926);
and U11050 (N_11050,N_7121,N_6836);
or U11051 (N_11051,N_8182,N_7619);
and U11052 (N_11052,N_8818,N_6980);
or U11053 (N_11053,N_9018,N_9011);
and U11054 (N_11054,N_8973,N_8838);
nand U11055 (N_11055,N_9089,N_7229);
xor U11056 (N_11056,N_6872,N_9074);
nand U11057 (N_11057,N_9183,N_8905);
nor U11058 (N_11058,N_7016,N_7785);
nand U11059 (N_11059,N_6912,N_7720);
and U11060 (N_11060,N_7410,N_7287);
or U11061 (N_11061,N_9131,N_7283);
and U11062 (N_11062,N_7882,N_6998);
or U11063 (N_11063,N_7647,N_9103);
or U11064 (N_11064,N_8416,N_7120);
xnor U11065 (N_11065,N_7447,N_9321);
nand U11066 (N_11066,N_7488,N_6919);
and U11067 (N_11067,N_6959,N_8496);
nor U11068 (N_11068,N_9268,N_8317);
or U11069 (N_11069,N_7320,N_6919);
and U11070 (N_11070,N_8409,N_6353);
nand U11071 (N_11071,N_7229,N_9339);
nand U11072 (N_11072,N_7015,N_9328);
or U11073 (N_11073,N_8272,N_6639);
xor U11074 (N_11074,N_8704,N_8929);
nand U11075 (N_11075,N_8148,N_7672);
or U11076 (N_11076,N_7914,N_7656);
xor U11077 (N_11077,N_8799,N_6725);
and U11078 (N_11078,N_7349,N_7438);
nand U11079 (N_11079,N_7864,N_7173);
nor U11080 (N_11080,N_7689,N_7511);
and U11081 (N_11081,N_8878,N_6527);
nor U11082 (N_11082,N_8756,N_8052);
or U11083 (N_11083,N_8961,N_8610);
nor U11084 (N_11084,N_7161,N_6620);
or U11085 (N_11085,N_6969,N_7215);
nand U11086 (N_11086,N_8385,N_8321);
nor U11087 (N_11087,N_7755,N_8634);
or U11088 (N_11088,N_6360,N_8669);
xor U11089 (N_11089,N_6883,N_9003);
nor U11090 (N_11090,N_6701,N_7758);
or U11091 (N_11091,N_9260,N_8774);
or U11092 (N_11092,N_7035,N_7060);
and U11093 (N_11093,N_8244,N_8080);
nor U11094 (N_11094,N_6715,N_8444);
nand U11095 (N_11095,N_7697,N_7156);
or U11096 (N_11096,N_6868,N_8242);
or U11097 (N_11097,N_8062,N_8569);
and U11098 (N_11098,N_6610,N_7515);
xnor U11099 (N_11099,N_6438,N_8919);
or U11100 (N_11100,N_7242,N_8377);
nand U11101 (N_11101,N_7255,N_6487);
nand U11102 (N_11102,N_6519,N_7275);
or U11103 (N_11103,N_6799,N_8025);
nand U11104 (N_11104,N_7685,N_9218);
nand U11105 (N_11105,N_7272,N_8181);
or U11106 (N_11106,N_6827,N_8293);
or U11107 (N_11107,N_7976,N_6903);
or U11108 (N_11108,N_6593,N_8110);
and U11109 (N_11109,N_7769,N_9281);
nand U11110 (N_11110,N_8939,N_7421);
nor U11111 (N_11111,N_6345,N_7473);
or U11112 (N_11112,N_7079,N_6605);
or U11113 (N_11113,N_8053,N_7277);
xnor U11114 (N_11114,N_7573,N_8161);
nor U11115 (N_11115,N_6477,N_7351);
xnor U11116 (N_11116,N_9325,N_9330);
nand U11117 (N_11117,N_6876,N_7301);
nor U11118 (N_11118,N_6404,N_6386);
or U11119 (N_11119,N_6478,N_8217);
or U11120 (N_11120,N_8706,N_8389);
or U11121 (N_11121,N_6495,N_9167);
and U11122 (N_11122,N_6973,N_9102);
nand U11123 (N_11123,N_8406,N_7058);
nor U11124 (N_11124,N_8104,N_9187);
nor U11125 (N_11125,N_7929,N_8642);
nor U11126 (N_11126,N_7289,N_6616);
or U11127 (N_11127,N_8226,N_7556);
or U11128 (N_11128,N_7088,N_6987);
nor U11129 (N_11129,N_8275,N_8519);
nand U11130 (N_11130,N_6740,N_7430);
xnor U11131 (N_11131,N_6821,N_9184);
nor U11132 (N_11132,N_7027,N_7999);
or U11133 (N_11133,N_8142,N_8825);
xnor U11134 (N_11134,N_8089,N_6448);
nand U11135 (N_11135,N_6804,N_7655);
or U11136 (N_11136,N_8324,N_9174);
nor U11137 (N_11137,N_8182,N_6421);
nand U11138 (N_11138,N_7453,N_6587);
nand U11139 (N_11139,N_7440,N_9199);
or U11140 (N_11140,N_7836,N_6428);
nor U11141 (N_11141,N_6876,N_9332);
and U11142 (N_11142,N_7005,N_8732);
nand U11143 (N_11143,N_9051,N_7974);
and U11144 (N_11144,N_8889,N_8739);
or U11145 (N_11145,N_7067,N_6363);
nand U11146 (N_11146,N_7108,N_6447);
and U11147 (N_11147,N_6706,N_7049);
nor U11148 (N_11148,N_6673,N_7902);
nand U11149 (N_11149,N_6475,N_8699);
or U11150 (N_11150,N_8317,N_7188);
xnor U11151 (N_11151,N_7063,N_9283);
nor U11152 (N_11152,N_7637,N_7856);
or U11153 (N_11153,N_6480,N_7168);
or U11154 (N_11154,N_9250,N_6487);
nor U11155 (N_11155,N_9328,N_6254);
or U11156 (N_11156,N_7336,N_8680);
or U11157 (N_11157,N_6746,N_7330);
nand U11158 (N_11158,N_6908,N_7625);
nor U11159 (N_11159,N_7718,N_6575);
nor U11160 (N_11160,N_6491,N_9060);
and U11161 (N_11161,N_8222,N_6606);
nor U11162 (N_11162,N_6602,N_9334);
or U11163 (N_11163,N_7717,N_8471);
or U11164 (N_11164,N_7275,N_8267);
or U11165 (N_11165,N_7627,N_7113);
nand U11166 (N_11166,N_8523,N_8118);
or U11167 (N_11167,N_7428,N_7809);
and U11168 (N_11168,N_9357,N_9137);
nand U11169 (N_11169,N_8873,N_7824);
nand U11170 (N_11170,N_7592,N_7607);
nand U11171 (N_11171,N_8451,N_8534);
nand U11172 (N_11172,N_7587,N_6269);
or U11173 (N_11173,N_7377,N_6534);
xnor U11174 (N_11174,N_7363,N_6953);
and U11175 (N_11175,N_8129,N_8144);
or U11176 (N_11176,N_8683,N_9074);
and U11177 (N_11177,N_9267,N_8756);
and U11178 (N_11178,N_6391,N_6490);
and U11179 (N_11179,N_6412,N_8208);
or U11180 (N_11180,N_7997,N_7489);
and U11181 (N_11181,N_6344,N_8259);
or U11182 (N_11182,N_9167,N_8699);
and U11183 (N_11183,N_7159,N_8005);
and U11184 (N_11184,N_8973,N_6674);
or U11185 (N_11185,N_7562,N_6525);
nand U11186 (N_11186,N_9284,N_6407);
xnor U11187 (N_11187,N_6416,N_7495);
nor U11188 (N_11188,N_8291,N_7183);
and U11189 (N_11189,N_9215,N_6753);
or U11190 (N_11190,N_7430,N_8137);
nor U11191 (N_11191,N_7112,N_8665);
and U11192 (N_11192,N_6784,N_7217);
xnor U11193 (N_11193,N_7779,N_6434);
nand U11194 (N_11194,N_6874,N_9155);
nand U11195 (N_11195,N_7470,N_6935);
nor U11196 (N_11196,N_7761,N_6638);
and U11197 (N_11197,N_6969,N_6287);
or U11198 (N_11198,N_8985,N_8237);
or U11199 (N_11199,N_7275,N_7493);
or U11200 (N_11200,N_8483,N_6730);
or U11201 (N_11201,N_7165,N_8620);
or U11202 (N_11202,N_8513,N_6389);
xnor U11203 (N_11203,N_8837,N_6259);
and U11204 (N_11204,N_8389,N_7213);
xor U11205 (N_11205,N_9232,N_7045);
xnor U11206 (N_11206,N_6728,N_8327);
or U11207 (N_11207,N_7232,N_8206);
nor U11208 (N_11208,N_7526,N_7065);
nand U11209 (N_11209,N_7958,N_6793);
nand U11210 (N_11210,N_6697,N_8230);
or U11211 (N_11211,N_8646,N_9286);
nor U11212 (N_11212,N_6455,N_8786);
and U11213 (N_11213,N_7411,N_8592);
and U11214 (N_11214,N_8705,N_7220);
xnor U11215 (N_11215,N_7560,N_6319);
nor U11216 (N_11216,N_7757,N_7374);
or U11217 (N_11217,N_7539,N_6797);
and U11218 (N_11218,N_8911,N_7585);
nor U11219 (N_11219,N_8155,N_8979);
xor U11220 (N_11220,N_8012,N_6831);
nand U11221 (N_11221,N_8421,N_9244);
nor U11222 (N_11222,N_8396,N_7941);
nand U11223 (N_11223,N_8294,N_7399);
or U11224 (N_11224,N_6274,N_9106);
and U11225 (N_11225,N_7908,N_8236);
or U11226 (N_11226,N_6716,N_6552);
nand U11227 (N_11227,N_6905,N_9097);
and U11228 (N_11228,N_8947,N_8844);
xnor U11229 (N_11229,N_7115,N_8552);
or U11230 (N_11230,N_7678,N_6609);
or U11231 (N_11231,N_9284,N_7816);
and U11232 (N_11232,N_7552,N_8397);
nor U11233 (N_11233,N_8957,N_6521);
nor U11234 (N_11234,N_7254,N_6768);
nor U11235 (N_11235,N_9326,N_8358);
xnor U11236 (N_11236,N_8990,N_6667);
and U11237 (N_11237,N_8316,N_7596);
nor U11238 (N_11238,N_9115,N_8125);
nor U11239 (N_11239,N_6525,N_8754);
or U11240 (N_11240,N_7390,N_8623);
nand U11241 (N_11241,N_8569,N_6581);
nor U11242 (N_11242,N_7342,N_6750);
and U11243 (N_11243,N_6633,N_7583);
nor U11244 (N_11244,N_7422,N_8144);
xor U11245 (N_11245,N_7050,N_6618);
or U11246 (N_11246,N_6834,N_8210);
or U11247 (N_11247,N_7922,N_6291);
nor U11248 (N_11248,N_8118,N_9216);
and U11249 (N_11249,N_6332,N_8560);
nand U11250 (N_11250,N_7226,N_6491);
nand U11251 (N_11251,N_6412,N_6981);
nand U11252 (N_11252,N_8944,N_6636);
and U11253 (N_11253,N_8722,N_7831);
nor U11254 (N_11254,N_8777,N_6424);
or U11255 (N_11255,N_8677,N_6530);
nand U11256 (N_11256,N_6487,N_7655);
nand U11257 (N_11257,N_7620,N_7996);
or U11258 (N_11258,N_7264,N_6875);
or U11259 (N_11259,N_8395,N_8848);
nand U11260 (N_11260,N_8763,N_7518);
xor U11261 (N_11261,N_7147,N_6704);
nand U11262 (N_11262,N_8279,N_7089);
nand U11263 (N_11263,N_7482,N_8260);
and U11264 (N_11264,N_6942,N_7594);
nor U11265 (N_11265,N_7406,N_8554);
or U11266 (N_11266,N_6593,N_8933);
nand U11267 (N_11267,N_6367,N_8785);
and U11268 (N_11268,N_7540,N_6755);
nor U11269 (N_11269,N_6899,N_9054);
and U11270 (N_11270,N_6312,N_7810);
or U11271 (N_11271,N_7194,N_7714);
nor U11272 (N_11272,N_8389,N_6453);
and U11273 (N_11273,N_6778,N_7366);
nor U11274 (N_11274,N_7296,N_8264);
xor U11275 (N_11275,N_7077,N_6608);
and U11276 (N_11276,N_8282,N_7964);
nor U11277 (N_11277,N_8031,N_7324);
or U11278 (N_11278,N_9286,N_7527);
or U11279 (N_11279,N_7002,N_9346);
nand U11280 (N_11280,N_9028,N_8918);
or U11281 (N_11281,N_8832,N_8591);
nand U11282 (N_11282,N_7086,N_8740);
nor U11283 (N_11283,N_8974,N_9014);
and U11284 (N_11284,N_6555,N_7300);
nor U11285 (N_11285,N_7174,N_8583);
nor U11286 (N_11286,N_8941,N_7023);
nand U11287 (N_11287,N_6264,N_6730);
nor U11288 (N_11288,N_9041,N_8773);
nor U11289 (N_11289,N_6734,N_8125);
nor U11290 (N_11290,N_6560,N_7551);
and U11291 (N_11291,N_8520,N_8512);
nand U11292 (N_11292,N_8060,N_7578);
nor U11293 (N_11293,N_7458,N_8476);
and U11294 (N_11294,N_9117,N_7166);
nor U11295 (N_11295,N_8339,N_8012);
nand U11296 (N_11296,N_8854,N_6649);
xor U11297 (N_11297,N_7031,N_7077);
xnor U11298 (N_11298,N_8716,N_8066);
nor U11299 (N_11299,N_8377,N_6763);
nand U11300 (N_11300,N_6296,N_8700);
nand U11301 (N_11301,N_7437,N_8024);
nand U11302 (N_11302,N_9141,N_8070);
xor U11303 (N_11303,N_7729,N_8560);
nand U11304 (N_11304,N_9225,N_7886);
or U11305 (N_11305,N_9334,N_7200);
nand U11306 (N_11306,N_6704,N_6955);
xnor U11307 (N_11307,N_7625,N_8758);
and U11308 (N_11308,N_7207,N_7040);
nor U11309 (N_11309,N_9079,N_6597);
or U11310 (N_11310,N_7908,N_6452);
nand U11311 (N_11311,N_7206,N_8907);
xnor U11312 (N_11312,N_8709,N_8026);
nand U11313 (N_11313,N_6995,N_8224);
nand U11314 (N_11314,N_6408,N_6602);
or U11315 (N_11315,N_7469,N_9047);
or U11316 (N_11316,N_7726,N_7858);
or U11317 (N_11317,N_6324,N_7281);
nand U11318 (N_11318,N_6898,N_7020);
and U11319 (N_11319,N_9212,N_7015);
or U11320 (N_11320,N_9159,N_7293);
nand U11321 (N_11321,N_6396,N_8446);
or U11322 (N_11322,N_6874,N_7224);
and U11323 (N_11323,N_9114,N_7930);
and U11324 (N_11324,N_7632,N_6921);
and U11325 (N_11325,N_7325,N_8382);
nor U11326 (N_11326,N_6617,N_8331);
nor U11327 (N_11327,N_6356,N_8320);
and U11328 (N_11328,N_6734,N_9008);
and U11329 (N_11329,N_7023,N_6894);
nand U11330 (N_11330,N_8424,N_7870);
and U11331 (N_11331,N_8201,N_8840);
or U11332 (N_11332,N_8180,N_9010);
nand U11333 (N_11333,N_6342,N_6863);
or U11334 (N_11334,N_9302,N_8434);
and U11335 (N_11335,N_7155,N_7255);
nor U11336 (N_11336,N_6864,N_7209);
nand U11337 (N_11337,N_6322,N_7368);
nor U11338 (N_11338,N_6687,N_7905);
nand U11339 (N_11339,N_8469,N_7061);
or U11340 (N_11340,N_6989,N_8914);
and U11341 (N_11341,N_8438,N_8972);
nor U11342 (N_11342,N_7102,N_6833);
xor U11343 (N_11343,N_8151,N_6876);
xnor U11344 (N_11344,N_9283,N_8672);
nor U11345 (N_11345,N_8702,N_8567);
nand U11346 (N_11346,N_8332,N_7282);
nor U11347 (N_11347,N_6262,N_6396);
nand U11348 (N_11348,N_7908,N_7000);
xnor U11349 (N_11349,N_6794,N_6734);
nand U11350 (N_11350,N_7236,N_9127);
nor U11351 (N_11351,N_8283,N_6731);
xor U11352 (N_11352,N_8004,N_9209);
or U11353 (N_11353,N_9078,N_6302);
nor U11354 (N_11354,N_7103,N_7207);
nand U11355 (N_11355,N_8740,N_7721);
xor U11356 (N_11356,N_7565,N_9262);
nand U11357 (N_11357,N_8312,N_7164);
and U11358 (N_11358,N_6407,N_9208);
or U11359 (N_11359,N_6343,N_7134);
xor U11360 (N_11360,N_8781,N_6530);
xnor U11361 (N_11361,N_8552,N_7990);
xnor U11362 (N_11362,N_7602,N_7029);
nor U11363 (N_11363,N_8937,N_9317);
nand U11364 (N_11364,N_7714,N_9101);
nor U11365 (N_11365,N_9016,N_6304);
or U11366 (N_11366,N_7824,N_7435);
nand U11367 (N_11367,N_6908,N_7878);
and U11368 (N_11368,N_8539,N_8227);
nand U11369 (N_11369,N_7627,N_7015);
and U11370 (N_11370,N_6551,N_6264);
nand U11371 (N_11371,N_8197,N_7006);
or U11372 (N_11372,N_7668,N_7551);
and U11373 (N_11373,N_8098,N_7998);
nor U11374 (N_11374,N_6587,N_8305);
nor U11375 (N_11375,N_6260,N_9113);
nor U11376 (N_11376,N_6740,N_9040);
xor U11377 (N_11377,N_8534,N_8896);
xor U11378 (N_11378,N_6398,N_8879);
nand U11379 (N_11379,N_8163,N_8088);
and U11380 (N_11380,N_6624,N_7320);
and U11381 (N_11381,N_6930,N_7555);
nand U11382 (N_11382,N_8371,N_8921);
xnor U11383 (N_11383,N_8334,N_6577);
nand U11384 (N_11384,N_7772,N_8807);
xor U11385 (N_11385,N_6461,N_9318);
xnor U11386 (N_11386,N_8775,N_8366);
nand U11387 (N_11387,N_7456,N_7338);
nor U11388 (N_11388,N_7657,N_6397);
and U11389 (N_11389,N_7262,N_8210);
nor U11390 (N_11390,N_6335,N_8367);
nand U11391 (N_11391,N_6372,N_7870);
or U11392 (N_11392,N_8504,N_7819);
nor U11393 (N_11393,N_8139,N_7094);
and U11394 (N_11394,N_7707,N_6645);
nor U11395 (N_11395,N_7598,N_8841);
and U11396 (N_11396,N_8985,N_6741);
xor U11397 (N_11397,N_8997,N_8642);
or U11398 (N_11398,N_9046,N_9295);
and U11399 (N_11399,N_8735,N_7012);
nor U11400 (N_11400,N_7121,N_8348);
nor U11401 (N_11401,N_8936,N_9022);
and U11402 (N_11402,N_8857,N_8561);
or U11403 (N_11403,N_7074,N_6601);
and U11404 (N_11404,N_6328,N_6535);
or U11405 (N_11405,N_6627,N_7941);
nor U11406 (N_11406,N_7817,N_9094);
and U11407 (N_11407,N_6721,N_8778);
or U11408 (N_11408,N_9021,N_9125);
xor U11409 (N_11409,N_8931,N_6567);
nor U11410 (N_11410,N_6449,N_7204);
or U11411 (N_11411,N_8715,N_7895);
and U11412 (N_11412,N_6300,N_7122);
or U11413 (N_11413,N_7270,N_6665);
nand U11414 (N_11414,N_9374,N_7158);
nor U11415 (N_11415,N_8114,N_7063);
xnor U11416 (N_11416,N_8393,N_8045);
nor U11417 (N_11417,N_8410,N_8387);
nand U11418 (N_11418,N_6573,N_9279);
nand U11419 (N_11419,N_6942,N_9182);
and U11420 (N_11420,N_7589,N_8944);
nor U11421 (N_11421,N_7530,N_9129);
nor U11422 (N_11422,N_8837,N_7806);
or U11423 (N_11423,N_8555,N_6284);
and U11424 (N_11424,N_8540,N_8818);
and U11425 (N_11425,N_7143,N_6604);
and U11426 (N_11426,N_8467,N_6851);
nor U11427 (N_11427,N_6486,N_8376);
nor U11428 (N_11428,N_6432,N_7722);
and U11429 (N_11429,N_8280,N_9338);
or U11430 (N_11430,N_6819,N_7930);
or U11431 (N_11431,N_7548,N_8774);
or U11432 (N_11432,N_6903,N_6837);
and U11433 (N_11433,N_9202,N_6322);
nand U11434 (N_11434,N_7848,N_9191);
nor U11435 (N_11435,N_7372,N_8948);
nand U11436 (N_11436,N_7089,N_8082);
nand U11437 (N_11437,N_9321,N_6844);
and U11438 (N_11438,N_7457,N_7501);
nor U11439 (N_11439,N_8835,N_8970);
nand U11440 (N_11440,N_7212,N_9146);
or U11441 (N_11441,N_8327,N_6825);
nand U11442 (N_11442,N_8991,N_6636);
or U11443 (N_11443,N_6549,N_8838);
nor U11444 (N_11444,N_8042,N_7695);
nor U11445 (N_11445,N_6944,N_8525);
nor U11446 (N_11446,N_8969,N_8230);
and U11447 (N_11447,N_6499,N_9047);
and U11448 (N_11448,N_8233,N_6580);
or U11449 (N_11449,N_9066,N_8974);
nand U11450 (N_11450,N_8656,N_6275);
nor U11451 (N_11451,N_7209,N_8161);
nor U11452 (N_11452,N_6659,N_8856);
nor U11453 (N_11453,N_8610,N_6740);
nor U11454 (N_11454,N_7192,N_6574);
nand U11455 (N_11455,N_8153,N_9137);
and U11456 (N_11456,N_6973,N_6816);
and U11457 (N_11457,N_7074,N_7655);
or U11458 (N_11458,N_6685,N_8358);
or U11459 (N_11459,N_8354,N_7014);
and U11460 (N_11460,N_8514,N_7871);
nor U11461 (N_11461,N_8726,N_7697);
xnor U11462 (N_11462,N_7482,N_7265);
or U11463 (N_11463,N_8289,N_6927);
or U11464 (N_11464,N_7564,N_7115);
nand U11465 (N_11465,N_8397,N_8631);
or U11466 (N_11466,N_7028,N_7361);
nor U11467 (N_11467,N_8403,N_9055);
nand U11468 (N_11468,N_7984,N_8203);
or U11469 (N_11469,N_6720,N_8914);
and U11470 (N_11470,N_7846,N_8910);
or U11471 (N_11471,N_7492,N_9232);
xnor U11472 (N_11472,N_8657,N_8484);
nor U11473 (N_11473,N_7723,N_8830);
or U11474 (N_11474,N_8392,N_7558);
and U11475 (N_11475,N_8585,N_8812);
nor U11476 (N_11476,N_8660,N_8386);
and U11477 (N_11477,N_8098,N_8120);
and U11478 (N_11478,N_9078,N_7475);
or U11479 (N_11479,N_6576,N_7818);
and U11480 (N_11480,N_6693,N_7867);
xor U11481 (N_11481,N_6570,N_7069);
nand U11482 (N_11482,N_8667,N_7518);
nand U11483 (N_11483,N_7242,N_7816);
nor U11484 (N_11484,N_8269,N_8839);
or U11485 (N_11485,N_8638,N_8436);
and U11486 (N_11486,N_8253,N_8672);
and U11487 (N_11487,N_7048,N_7572);
nand U11488 (N_11488,N_8425,N_8510);
or U11489 (N_11489,N_8406,N_8056);
nand U11490 (N_11490,N_7484,N_8501);
nor U11491 (N_11491,N_6813,N_9306);
or U11492 (N_11492,N_7610,N_7178);
nor U11493 (N_11493,N_6404,N_8020);
nor U11494 (N_11494,N_6654,N_7374);
or U11495 (N_11495,N_8881,N_7304);
nand U11496 (N_11496,N_7922,N_7196);
xnor U11497 (N_11497,N_7749,N_8245);
nand U11498 (N_11498,N_7442,N_9255);
or U11499 (N_11499,N_8209,N_7100);
and U11500 (N_11500,N_7742,N_7723);
nand U11501 (N_11501,N_6537,N_7035);
nand U11502 (N_11502,N_9359,N_8715);
nand U11503 (N_11503,N_6457,N_7148);
and U11504 (N_11504,N_7273,N_6622);
nand U11505 (N_11505,N_8069,N_7817);
xor U11506 (N_11506,N_6645,N_6635);
or U11507 (N_11507,N_6347,N_7748);
nor U11508 (N_11508,N_6860,N_6730);
nor U11509 (N_11509,N_8803,N_6629);
nor U11510 (N_11510,N_7101,N_7841);
nor U11511 (N_11511,N_8171,N_7711);
or U11512 (N_11512,N_8496,N_6762);
and U11513 (N_11513,N_8803,N_8304);
xnor U11514 (N_11514,N_7662,N_8503);
xor U11515 (N_11515,N_8836,N_9225);
nand U11516 (N_11516,N_6556,N_7983);
xnor U11517 (N_11517,N_8002,N_8196);
nor U11518 (N_11518,N_9152,N_8573);
nor U11519 (N_11519,N_8351,N_7611);
nand U11520 (N_11520,N_7439,N_9169);
nor U11521 (N_11521,N_7178,N_8329);
nand U11522 (N_11522,N_7216,N_7028);
xor U11523 (N_11523,N_8950,N_8439);
and U11524 (N_11524,N_7060,N_8259);
or U11525 (N_11525,N_6955,N_8400);
nor U11526 (N_11526,N_8660,N_6769);
nor U11527 (N_11527,N_8033,N_8066);
nor U11528 (N_11528,N_6707,N_8225);
or U11529 (N_11529,N_6326,N_7828);
or U11530 (N_11530,N_9138,N_7522);
nor U11531 (N_11531,N_7289,N_8181);
nor U11532 (N_11532,N_7279,N_8507);
or U11533 (N_11533,N_7078,N_9140);
or U11534 (N_11534,N_6711,N_8873);
or U11535 (N_11535,N_6879,N_7562);
or U11536 (N_11536,N_8754,N_9350);
or U11537 (N_11537,N_7655,N_8466);
and U11538 (N_11538,N_6759,N_8223);
or U11539 (N_11539,N_8966,N_8037);
nor U11540 (N_11540,N_6369,N_6339);
and U11541 (N_11541,N_7614,N_6472);
nand U11542 (N_11542,N_6745,N_8198);
xnor U11543 (N_11543,N_7093,N_7228);
xnor U11544 (N_11544,N_6934,N_8007);
nand U11545 (N_11545,N_6518,N_6523);
and U11546 (N_11546,N_8053,N_6808);
nor U11547 (N_11547,N_6642,N_9076);
and U11548 (N_11548,N_8955,N_8151);
nand U11549 (N_11549,N_7645,N_8848);
or U11550 (N_11550,N_7673,N_8437);
or U11551 (N_11551,N_6822,N_8421);
or U11552 (N_11552,N_8659,N_8190);
nor U11553 (N_11553,N_7376,N_8438);
xnor U11554 (N_11554,N_6980,N_8398);
xnor U11555 (N_11555,N_7140,N_9117);
or U11556 (N_11556,N_7691,N_7632);
and U11557 (N_11557,N_9132,N_6889);
nand U11558 (N_11558,N_9257,N_8030);
nor U11559 (N_11559,N_8883,N_8019);
xor U11560 (N_11560,N_9128,N_7111);
or U11561 (N_11561,N_7976,N_7140);
or U11562 (N_11562,N_8850,N_7733);
or U11563 (N_11563,N_7212,N_7330);
nor U11564 (N_11564,N_9141,N_8277);
or U11565 (N_11565,N_7518,N_7502);
nand U11566 (N_11566,N_9134,N_6374);
nor U11567 (N_11567,N_8081,N_6862);
or U11568 (N_11568,N_7919,N_6584);
nor U11569 (N_11569,N_7013,N_7973);
or U11570 (N_11570,N_6749,N_7510);
nand U11571 (N_11571,N_8048,N_7727);
and U11572 (N_11572,N_8262,N_8447);
and U11573 (N_11573,N_8566,N_7549);
nand U11574 (N_11574,N_8607,N_9228);
nand U11575 (N_11575,N_9176,N_6321);
and U11576 (N_11576,N_7797,N_7293);
nand U11577 (N_11577,N_8770,N_8734);
nand U11578 (N_11578,N_7308,N_7606);
or U11579 (N_11579,N_7361,N_8005);
xor U11580 (N_11580,N_9110,N_6425);
xor U11581 (N_11581,N_8329,N_8953);
and U11582 (N_11582,N_7015,N_7779);
and U11583 (N_11583,N_7726,N_7406);
or U11584 (N_11584,N_8199,N_8648);
nand U11585 (N_11585,N_7683,N_8381);
or U11586 (N_11586,N_7102,N_7516);
nor U11587 (N_11587,N_8570,N_7512);
or U11588 (N_11588,N_8854,N_9083);
or U11589 (N_11589,N_7898,N_8837);
or U11590 (N_11590,N_7637,N_6622);
and U11591 (N_11591,N_7099,N_6894);
nor U11592 (N_11592,N_9079,N_6799);
or U11593 (N_11593,N_8815,N_8437);
and U11594 (N_11594,N_7682,N_7044);
and U11595 (N_11595,N_8841,N_8534);
or U11596 (N_11596,N_9015,N_8152);
or U11597 (N_11597,N_8008,N_6329);
nand U11598 (N_11598,N_8079,N_8781);
or U11599 (N_11599,N_7479,N_7896);
and U11600 (N_11600,N_6480,N_6429);
nor U11601 (N_11601,N_6294,N_8622);
nand U11602 (N_11602,N_8934,N_8633);
nand U11603 (N_11603,N_7703,N_8939);
and U11604 (N_11604,N_9338,N_9060);
and U11605 (N_11605,N_6783,N_8514);
or U11606 (N_11606,N_7361,N_9179);
or U11607 (N_11607,N_6844,N_8014);
and U11608 (N_11608,N_6778,N_9171);
and U11609 (N_11609,N_8295,N_7338);
and U11610 (N_11610,N_8558,N_7264);
nand U11611 (N_11611,N_7612,N_9293);
nor U11612 (N_11612,N_6913,N_7373);
or U11613 (N_11613,N_7786,N_7340);
and U11614 (N_11614,N_9058,N_8231);
or U11615 (N_11615,N_8701,N_6914);
nand U11616 (N_11616,N_8360,N_7234);
nor U11617 (N_11617,N_6549,N_8295);
and U11618 (N_11618,N_6951,N_6915);
or U11619 (N_11619,N_6585,N_7717);
and U11620 (N_11620,N_8909,N_8996);
nand U11621 (N_11621,N_8622,N_8237);
and U11622 (N_11622,N_8049,N_9219);
nor U11623 (N_11623,N_7770,N_6664);
nor U11624 (N_11624,N_7684,N_6538);
or U11625 (N_11625,N_6303,N_8327);
nor U11626 (N_11626,N_9032,N_9027);
and U11627 (N_11627,N_6897,N_8978);
xnor U11628 (N_11628,N_7162,N_9117);
nand U11629 (N_11629,N_7348,N_6900);
xnor U11630 (N_11630,N_9188,N_9166);
and U11631 (N_11631,N_7785,N_9150);
nor U11632 (N_11632,N_7556,N_7939);
or U11633 (N_11633,N_8947,N_6985);
nand U11634 (N_11634,N_7488,N_6628);
and U11635 (N_11635,N_8522,N_8409);
xnor U11636 (N_11636,N_8995,N_6981);
nor U11637 (N_11637,N_7917,N_6600);
or U11638 (N_11638,N_9101,N_6632);
nand U11639 (N_11639,N_6998,N_6992);
xnor U11640 (N_11640,N_7026,N_7179);
or U11641 (N_11641,N_8432,N_6568);
xor U11642 (N_11642,N_7646,N_8569);
or U11643 (N_11643,N_8324,N_9217);
xnor U11644 (N_11644,N_6762,N_8004);
or U11645 (N_11645,N_6316,N_8761);
and U11646 (N_11646,N_6373,N_8639);
or U11647 (N_11647,N_6689,N_7624);
and U11648 (N_11648,N_7458,N_6793);
or U11649 (N_11649,N_7533,N_7362);
nor U11650 (N_11650,N_7039,N_8461);
nor U11651 (N_11651,N_8123,N_8735);
nor U11652 (N_11652,N_9100,N_8878);
nand U11653 (N_11653,N_6253,N_9342);
nand U11654 (N_11654,N_7081,N_7309);
and U11655 (N_11655,N_6256,N_8147);
and U11656 (N_11656,N_7504,N_6846);
or U11657 (N_11657,N_8251,N_9023);
or U11658 (N_11658,N_8847,N_8773);
or U11659 (N_11659,N_7885,N_7786);
and U11660 (N_11660,N_8973,N_8691);
xnor U11661 (N_11661,N_7931,N_9363);
or U11662 (N_11662,N_8101,N_7051);
nand U11663 (N_11663,N_7518,N_7821);
nand U11664 (N_11664,N_9340,N_8858);
or U11665 (N_11665,N_8679,N_7355);
or U11666 (N_11666,N_8617,N_7155);
xnor U11667 (N_11667,N_8911,N_6372);
or U11668 (N_11668,N_9352,N_7008);
and U11669 (N_11669,N_6428,N_9084);
and U11670 (N_11670,N_6292,N_8011);
or U11671 (N_11671,N_9256,N_9301);
nand U11672 (N_11672,N_8052,N_8739);
and U11673 (N_11673,N_7706,N_7753);
nand U11674 (N_11674,N_7088,N_6702);
or U11675 (N_11675,N_7036,N_7516);
or U11676 (N_11676,N_8199,N_6545);
nor U11677 (N_11677,N_7129,N_7399);
or U11678 (N_11678,N_9168,N_8666);
and U11679 (N_11679,N_7572,N_8668);
nor U11680 (N_11680,N_7204,N_8774);
nand U11681 (N_11681,N_6627,N_7147);
or U11682 (N_11682,N_8833,N_8144);
and U11683 (N_11683,N_8379,N_7233);
or U11684 (N_11684,N_8887,N_9206);
and U11685 (N_11685,N_7448,N_8972);
and U11686 (N_11686,N_6895,N_8821);
or U11687 (N_11687,N_6550,N_8801);
nand U11688 (N_11688,N_6477,N_6484);
xor U11689 (N_11689,N_7762,N_7804);
nor U11690 (N_11690,N_6790,N_8898);
nor U11691 (N_11691,N_8264,N_7424);
nand U11692 (N_11692,N_9114,N_7987);
or U11693 (N_11693,N_8198,N_7800);
nand U11694 (N_11694,N_7339,N_8848);
or U11695 (N_11695,N_7492,N_8673);
and U11696 (N_11696,N_8354,N_6947);
or U11697 (N_11697,N_7884,N_9164);
and U11698 (N_11698,N_7123,N_7650);
and U11699 (N_11699,N_8920,N_6571);
and U11700 (N_11700,N_7505,N_6420);
xor U11701 (N_11701,N_8685,N_9225);
nor U11702 (N_11702,N_7295,N_8868);
and U11703 (N_11703,N_8548,N_9206);
and U11704 (N_11704,N_7264,N_7865);
and U11705 (N_11705,N_8464,N_8400);
and U11706 (N_11706,N_7286,N_8763);
or U11707 (N_11707,N_8077,N_7167);
and U11708 (N_11708,N_8193,N_8968);
and U11709 (N_11709,N_8371,N_7568);
nor U11710 (N_11710,N_6716,N_7316);
nand U11711 (N_11711,N_8042,N_9272);
or U11712 (N_11712,N_7294,N_8257);
nand U11713 (N_11713,N_6411,N_9004);
and U11714 (N_11714,N_7544,N_7790);
nand U11715 (N_11715,N_8551,N_8497);
nor U11716 (N_11716,N_8133,N_9056);
nand U11717 (N_11717,N_8153,N_6443);
or U11718 (N_11718,N_8625,N_7452);
nor U11719 (N_11719,N_9342,N_8163);
and U11720 (N_11720,N_8786,N_7387);
nor U11721 (N_11721,N_8004,N_7987);
and U11722 (N_11722,N_7478,N_7923);
or U11723 (N_11723,N_8407,N_6492);
nor U11724 (N_11724,N_8954,N_7558);
and U11725 (N_11725,N_6998,N_7640);
or U11726 (N_11726,N_7973,N_6833);
xnor U11727 (N_11727,N_8338,N_7596);
nor U11728 (N_11728,N_8906,N_9167);
nor U11729 (N_11729,N_9209,N_8778);
nor U11730 (N_11730,N_6964,N_7483);
and U11731 (N_11731,N_8066,N_7412);
or U11732 (N_11732,N_8755,N_7900);
or U11733 (N_11733,N_6515,N_8023);
and U11734 (N_11734,N_8377,N_7382);
nor U11735 (N_11735,N_8541,N_8861);
and U11736 (N_11736,N_6290,N_8918);
and U11737 (N_11737,N_7333,N_8943);
xnor U11738 (N_11738,N_8188,N_8258);
nand U11739 (N_11739,N_6299,N_8500);
nand U11740 (N_11740,N_9229,N_8346);
nor U11741 (N_11741,N_8752,N_7225);
or U11742 (N_11742,N_7485,N_9349);
or U11743 (N_11743,N_7850,N_8269);
nor U11744 (N_11744,N_8200,N_8073);
nand U11745 (N_11745,N_7208,N_7168);
nand U11746 (N_11746,N_8787,N_8556);
nor U11747 (N_11747,N_6763,N_7523);
and U11748 (N_11748,N_7549,N_8196);
or U11749 (N_11749,N_6288,N_7956);
nand U11750 (N_11750,N_7314,N_7566);
or U11751 (N_11751,N_6989,N_6297);
nor U11752 (N_11752,N_7790,N_9289);
nand U11753 (N_11753,N_8386,N_8204);
xnor U11754 (N_11754,N_7056,N_6829);
nand U11755 (N_11755,N_8310,N_7355);
nand U11756 (N_11756,N_6613,N_6912);
or U11757 (N_11757,N_9038,N_6698);
nand U11758 (N_11758,N_6276,N_8011);
or U11759 (N_11759,N_9266,N_7850);
or U11760 (N_11760,N_8673,N_9102);
nor U11761 (N_11761,N_6675,N_8168);
or U11762 (N_11762,N_6567,N_8578);
nand U11763 (N_11763,N_7476,N_6596);
and U11764 (N_11764,N_7092,N_6367);
and U11765 (N_11765,N_8808,N_8128);
or U11766 (N_11766,N_7736,N_6414);
nor U11767 (N_11767,N_8691,N_6516);
nor U11768 (N_11768,N_6983,N_6788);
nor U11769 (N_11769,N_7087,N_7207);
and U11770 (N_11770,N_9171,N_8628);
nor U11771 (N_11771,N_7160,N_6927);
xnor U11772 (N_11772,N_8390,N_7837);
or U11773 (N_11773,N_7482,N_8314);
nand U11774 (N_11774,N_7254,N_7672);
nor U11775 (N_11775,N_8875,N_8561);
xor U11776 (N_11776,N_8080,N_6750);
nor U11777 (N_11777,N_8574,N_9331);
xnor U11778 (N_11778,N_8036,N_8393);
or U11779 (N_11779,N_7270,N_8823);
or U11780 (N_11780,N_6327,N_8596);
nor U11781 (N_11781,N_6961,N_6845);
nor U11782 (N_11782,N_6946,N_9338);
nor U11783 (N_11783,N_9224,N_6716);
or U11784 (N_11784,N_7665,N_9019);
and U11785 (N_11785,N_7121,N_6390);
nor U11786 (N_11786,N_7601,N_7863);
or U11787 (N_11787,N_8301,N_6279);
nand U11788 (N_11788,N_8887,N_7260);
and U11789 (N_11789,N_8048,N_8037);
or U11790 (N_11790,N_6892,N_8598);
or U11791 (N_11791,N_7735,N_9306);
nor U11792 (N_11792,N_6473,N_8534);
or U11793 (N_11793,N_8395,N_8489);
nor U11794 (N_11794,N_8206,N_8879);
and U11795 (N_11795,N_7593,N_8368);
or U11796 (N_11796,N_6922,N_9307);
or U11797 (N_11797,N_7974,N_6710);
xnor U11798 (N_11798,N_7942,N_8862);
nor U11799 (N_11799,N_7162,N_8975);
nand U11800 (N_11800,N_7808,N_7117);
nand U11801 (N_11801,N_6405,N_7485);
nand U11802 (N_11802,N_7752,N_7245);
nor U11803 (N_11803,N_8478,N_7212);
xnor U11804 (N_11804,N_7283,N_9204);
nor U11805 (N_11805,N_7554,N_8385);
and U11806 (N_11806,N_7581,N_8947);
and U11807 (N_11807,N_8563,N_6887);
and U11808 (N_11808,N_8221,N_7133);
nand U11809 (N_11809,N_8313,N_6258);
xor U11810 (N_11810,N_8801,N_8660);
xor U11811 (N_11811,N_8784,N_7909);
nand U11812 (N_11812,N_6303,N_6952);
nor U11813 (N_11813,N_6766,N_9348);
nor U11814 (N_11814,N_6334,N_8625);
nor U11815 (N_11815,N_6816,N_9078);
and U11816 (N_11816,N_6756,N_8081);
or U11817 (N_11817,N_9261,N_7322);
and U11818 (N_11818,N_7028,N_8926);
nand U11819 (N_11819,N_7703,N_9073);
nand U11820 (N_11820,N_7745,N_8469);
nand U11821 (N_11821,N_7495,N_8585);
xnor U11822 (N_11822,N_6626,N_7856);
or U11823 (N_11823,N_9343,N_8093);
and U11824 (N_11824,N_7727,N_6949);
nand U11825 (N_11825,N_8372,N_8963);
or U11826 (N_11826,N_6470,N_7287);
nor U11827 (N_11827,N_8414,N_8954);
nand U11828 (N_11828,N_6503,N_9290);
xor U11829 (N_11829,N_9143,N_8309);
and U11830 (N_11830,N_8450,N_8983);
nor U11831 (N_11831,N_6374,N_6578);
xnor U11832 (N_11832,N_7240,N_6671);
and U11833 (N_11833,N_8674,N_8377);
xnor U11834 (N_11834,N_7839,N_7321);
and U11835 (N_11835,N_8120,N_8883);
nor U11836 (N_11836,N_7158,N_7146);
nor U11837 (N_11837,N_7836,N_8462);
xor U11838 (N_11838,N_9262,N_8825);
nor U11839 (N_11839,N_6550,N_7268);
and U11840 (N_11840,N_8751,N_7127);
and U11841 (N_11841,N_8681,N_8127);
and U11842 (N_11842,N_9270,N_9036);
or U11843 (N_11843,N_8537,N_7290);
xnor U11844 (N_11844,N_7706,N_6731);
nor U11845 (N_11845,N_8465,N_6731);
xnor U11846 (N_11846,N_7709,N_8936);
or U11847 (N_11847,N_8012,N_7951);
or U11848 (N_11848,N_6463,N_7402);
or U11849 (N_11849,N_6449,N_8884);
and U11850 (N_11850,N_8988,N_6887);
and U11851 (N_11851,N_7062,N_7944);
or U11852 (N_11852,N_8371,N_7818);
nand U11853 (N_11853,N_8585,N_8061);
or U11854 (N_11854,N_8781,N_6470);
nand U11855 (N_11855,N_8604,N_8911);
nand U11856 (N_11856,N_9296,N_9315);
nor U11857 (N_11857,N_7024,N_8689);
and U11858 (N_11858,N_7753,N_6357);
nand U11859 (N_11859,N_8651,N_6802);
or U11860 (N_11860,N_8293,N_7562);
nand U11861 (N_11861,N_6922,N_6680);
nand U11862 (N_11862,N_6461,N_6926);
nand U11863 (N_11863,N_8081,N_6984);
nand U11864 (N_11864,N_8120,N_9137);
or U11865 (N_11865,N_7585,N_8355);
or U11866 (N_11866,N_7800,N_6626);
or U11867 (N_11867,N_7725,N_8774);
nor U11868 (N_11868,N_6567,N_7531);
nor U11869 (N_11869,N_7533,N_7105);
and U11870 (N_11870,N_8302,N_7738);
nor U11871 (N_11871,N_7437,N_9050);
or U11872 (N_11872,N_8962,N_9272);
nand U11873 (N_11873,N_6713,N_7953);
nand U11874 (N_11874,N_6979,N_6425);
or U11875 (N_11875,N_7989,N_7226);
xnor U11876 (N_11876,N_9315,N_8110);
or U11877 (N_11877,N_7180,N_7691);
nand U11878 (N_11878,N_6887,N_8683);
or U11879 (N_11879,N_8852,N_9143);
and U11880 (N_11880,N_6361,N_6355);
nor U11881 (N_11881,N_9059,N_7876);
nor U11882 (N_11882,N_9047,N_9153);
nor U11883 (N_11883,N_9210,N_9131);
nand U11884 (N_11884,N_8411,N_8019);
nor U11885 (N_11885,N_7686,N_9229);
nor U11886 (N_11886,N_7013,N_9309);
nand U11887 (N_11887,N_9006,N_8716);
nand U11888 (N_11888,N_9073,N_8711);
and U11889 (N_11889,N_7579,N_9101);
nand U11890 (N_11890,N_6524,N_7282);
nor U11891 (N_11891,N_7694,N_8784);
or U11892 (N_11892,N_7730,N_7334);
and U11893 (N_11893,N_7500,N_8675);
and U11894 (N_11894,N_8268,N_7975);
nor U11895 (N_11895,N_8597,N_9257);
nor U11896 (N_11896,N_7317,N_6876);
nand U11897 (N_11897,N_7820,N_8557);
xnor U11898 (N_11898,N_8131,N_9115);
nand U11899 (N_11899,N_9374,N_8762);
nor U11900 (N_11900,N_8735,N_6466);
nand U11901 (N_11901,N_6437,N_8006);
and U11902 (N_11902,N_6757,N_6833);
nor U11903 (N_11903,N_7088,N_7104);
nand U11904 (N_11904,N_7781,N_6776);
or U11905 (N_11905,N_8984,N_7151);
xnor U11906 (N_11906,N_7879,N_6772);
nor U11907 (N_11907,N_6439,N_7916);
or U11908 (N_11908,N_6525,N_6600);
nor U11909 (N_11909,N_7017,N_6684);
and U11910 (N_11910,N_6705,N_9162);
and U11911 (N_11911,N_7489,N_8168);
nand U11912 (N_11912,N_7713,N_7699);
nand U11913 (N_11913,N_8217,N_7569);
or U11914 (N_11914,N_8461,N_6391);
nor U11915 (N_11915,N_7957,N_8733);
and U11916 (N_11916,N_8645,N_6717);
and U11917 (N_11917,N_6906,N_7084);
or U11918 (N_11918,N_8530,N_7318);
nand U11919 (N_11919,N_7502,N_8005);
or U11920 (N_11920,N_8225,N_9116);
nor U11921 (N_11921,N_8276,N_7415);
and U11922 (N_11922,N_8514,N_7689);
or U11923 (N_11923,N_8537,N_6994);
and U11924 (N_11924,N_6661,N_9043);
and U11925 (N_11925,N_6448,N_8220);
xor U11926 (N_11926,N_7475,N_8396);
and U11927 (N_11927,N_9025,N_7194);
nor U11928 (N_11928,N_8306,N_6949);
nand U11929 (N_11929,N_7037,N_9276);
nand U11930 (N_11930,N_9351,N_7244);
nand U11931 (N_11931,N_8925,N_8331);
or U11932 (N_11932,N_9291,N_7952);
nor U11933 (N_11933,N_8173,N_8638);
or U11934 (N_11934,N_7335,N_8549);
or U11935 (N_11935,N_7471,N_6298);
nand U11936 (N_11936,N_9061,N_8543);
nor U11937 (N_11937,N_8536,N_6574);
or U11938 (N_11938,N_8455,N_7922);
nor U11939 (N_11939,N_7161,N_8705);
nor U11940 (N_11940,N_8003,N_7571);
and U11941 (N_11941,N_8500,N_7469);
nand U11942 (N_11942,N_7169,N_6864);
and U11943 (N_11943,N_7924,N_7397);
or U11944 (N_11944,N_8639,N_8824);
nand U11945 (N_11945,N_6699,N_7915);
nor U11946 (N_11946,N_6521,N_6558);
or U11947 (N_11947,N_7353,N_8050);
nand U11948 (N_11948,N_7505,N_7776);
or U11949 (N_11949,N_6995,N_7297);
or U11950 (N_11950,N_8888,N_8994);
nand U11951 (N_11951,N_8800,N_6444);
nand U11952 (N_11952,N_8716,N_7528);
xor U11953 (N_11953,N_6768,N_7823);
or U11954 (N_11954,N_6789,N_8464);
or U11955 (N_11955,N_7726,N_6298);
and U11956 (N_11956,N_7638,N_8780);
or U11957 (N_11957,N_8444,N_8960);
xor U11958 (N_11958,N_8279,N_6973);
nor U11959 (N_11959,N_9350,N_7970);
and U11960 (N_11960,N_8300,N_7031);
xnor U11961 (N_11961,N_6696,N_7272);
nand U11962 (N_11962,N_8647,N_7517);
nor U11963 (N_11963,N_9203,N_7207);
nor U11964 (N_11964,N_8613,N_6634);
nor U11965 (N_11965,N_8777,N_7694);
nand U11966 (N_11966,N_7257,N_6635);
xor U11967 (N_11967,N_7322,N_6676);
nand U11968 (N_11968,N_6816,N_9290);
or U11969 (N_11969,N_9078,N_6270);
nor U11970 (N_11970,N_9061,N_8526);
nor U11971 (N_11971,N_8353,N_7695);
and U11972 (N_11972,N_8091,N_7552);
or U11973 (N_11973,N_9267,N_9084);
or U11974 (N_11974,N_7883,N_8429);
or U11975 (N_11975,N_6856,N_8885);
or U11976 (N_11976,N_8998,N_8744);
nor U11977 (N_11977,N_7511,N_8898);
xnor U11978 (N_11978,N_7693,N_9097);
and U11979 (N_11979,N_9146,N_8704);
or U11980 (N_11980,N_8358,N_6951);
or U11981 (N_11981,N_6381,N_9064);
xor U11982 (N_11982,N_7379,N_8751);
nand U11983 (N_11983,N_7615,N_8990);
nand U11984 (N_11984,N_6493,N_7500);
and U11985 (N_11985,N_7465,N_8892);
and U11986 (N_11986,N_7000,N_8288);
nand U11987 (N_11987,N_9010,N_8760);
and U11988 (N_11988,N_7509,N_8541);
nor U11989 (N_11989,N_8175,N_6552);
nor U11990 (N_11990,N_6375,N_8745);
nor U11991 (N_11991,N_8512,N_8005);
xor U11992 (N_11992,N_8480,N_9035);
nand U11993 (N_11993,N_6925,N_7328);
nor U11994 (N_11994,N_6285,N_7915);
or U11995 (N_11995,N_8220,N_6893);
nand U11996 (N_11996,N_9297,N_6279);
xor U11997 (N_11997,N_9047,N_8789);
nor U11998 (N_11998,N_8801,N_7597);
nand U11999 (N_11999,N_8025,N_8562);
and U12000 (N_12000,N_7726,N_7072);
nand U12001 (N_12001,N_9083,N_7434);
nand U12002 (N_12002,N_7817,N_7532);
nor U12003 (N_12003,N_6859,N_9277);
nand U12004 (N_12004,N_7502,N_8734);
nand U12005 (N_12005,N_7010,N_6754);
and U12006 (N_12006,N_7712,N_9033);
nand U12007 (N_12007,N_7854,N_6669);
xor U12008 (N_12008,N_8761,N_8179);
nand U12009 (N_12009,N_8976,N_6846);
nand U12010 (N_12010,N_7142,N_6949);
nor U12011 (N_12011,N_9094,N_6927);
nor U12012 (N_12012,N_7167,N_8573);
or U12013 (N_12013,N_7468,N_7385);
and U12014 (N_12014,N_6972,N_8428);
or U12015 (N_12015,N_8554,N_8865);
and U12016 (N_12016,N_8783,N_7409);
nand U12017 (N_12017,N_7722,N_6479);
xnor U12018 (N_12018,N_7047,N_6445);
xor U12019 (N_12019,N_7819,N_6976);
nand U12020 (N_12020,N_7344,N_8116);
nor U12021 (N_12021,N_6773,N_7289);
and U12022 (N_12022,N_6251,N_7789);
nand U12023 (N_12023,N_7644,N_9260);
nand U12024 (N_12024,N_7763,N_9209);
nor U12025 (N_12025,N_7487,N_8827);
or U12026 (N_12026,N_7503,N_6642);
nand U12027 (N_12027,N_9193,N_9168);
xor U12028 (N_12028,N_6348,N_8628);
nand U12029 (N_12029,N_8381,N_6599);
xnor U12030 (N_12030,N_7363,N_7526);
nand U12031 (N_12031,N_8796,N_6874);
xnor U12032 (N_12032,N_9326,N_7730);
and U12033 (N_12033,N_6651,N_6347);
nand U12034 (N_12034,N_7348,N_9244);
or U12035 (N_12035,N_7171,N_6969);
nand U12036 (N_12036,N_6727,N_6774);
nor U12037 (N_12037,N_8380,N_6701);
nor U12038 (N_12038,N_7525,N_7695);
or U12039 (N_12039,N_7529,N_8172);
or U12040 (N_12040,N_8997,N_8273);
or U12041 (N_12041,N_8301,N_8863);
nand U12042 (N_12042,N_8070,N_8928);
nor U12043 (N_12043,N_7073,N_6765);
and U12044 (N_12044,N_7101,N_7027);
and U12045 (N_12045,N_9063,N_6553);
or U12046 (N_12046,N_6816,N_7555);
nand U12047 (N_12047,N_8579,N_6553);
and U12048 (N_12048,N_7107,N_9177);
and U12049 (N_12049,N_6474,N_6349);
and U12050 (N_12050,N_9014,N_8131);
nor U12051 (N_12051,N_6253,N_6361);
and U12052 (N_12052,N_9170,N_7845);
nand U12053 (N_12053,N_8089,N_7498);
nand U12054 (N_12054,N_8673,N_6853);
and U12055 (N_12055,N_7278,N_8916);
or U12056 (N_12056,N_6261,N_6847);
or U12057 (N_12057,N_8043,N_8821);
and U12058 (N_12058,N_7356,N_9279);
and U12059 (N_12059,N_9007,N_8495);
nor U12060 (N_12060,N_6526,N_7518);
nand U12061 (N_12061,N_7717,N_8405);
nor U12062 (N_12062,N_6733,N_8993);
or U12063 (N_12063,N_6830,N_9016);
and U12064 (N_12064,N_6740,N_9270);
xor U12065 (N_12065,N_6878,N_8047);
and U12066 (N_12066,N_6353,N_8628);
or U12067 (N_12067,N_8383,N_9018);
and U12068 (N_12068,N_9357,N_7365);
nor U12069 (N_12069,N_6889,N_9213);
or U12070 (N_12070,N_7359,N_9184);
or U12071 (N_12071,N_8578,N_8738);
nor U12072 (N_12072,N_7017,N_8302);
nor U12073 (N_12073,N_9354,N_7005);
nor U12074 (N_12074,N_6888,N_7623);
xor U12075 (N_12075,N_9140,N_7397);
or U12076 (N_12076,N_6879,N_6741);
nor U12077 (N_12077,N_7664,N_7017);
nand U12078 (N_12078,N_8285,N_7070);
or U12079 (N_12079,N_7807,N_7372);
nor U12080 (N_12080,N_9120,N_6476);
nand U12081 (N_12081,N_6560,N_8646);
nor U12082 (N_12082,N_9153,N_6759);
and U12083 (N_12083,N_8308,N_8040);
nand U12084 (N_12084,N_8638,N_6833);
nand U12085 (N_12085,N_9318,N_7493);
nand U12086 (N_12086,N_6670,N_6598);
or U12087 (N_12087,N_9349,N_8926);
and U12088 (N_12088,N_8952,N_7073);
nand U12089 (N_12089,N_7553,N_9221);
nor U12090 (N_12090,N_8489,N_8710);
nor U12091 (N_12091,N_7598,N_9241);
nand U12092 (N_12092,N_7087,N_6352);
or U12093 (N_12093,N_7553,N_6663);
nor U12094 (N_12094,N_8796,N_9195);
and U12095 (N_12095,N_7816,N_8632);
xnor U12096 (N_12096,N_8105,N_7773);
nor U12097 (N_12097,N_7719,N_7421);
or U12098 (N_12098,N_8069,N_8553);
and U12099 (N_12099,N_6359,N_6720);
nand U12100 (N_12100,N_6507,N_8553);
nand U12101 (N_12101,N_6746,N_7709);
or U12102 (N_12102,N_8854,N_8722);
and U12103 (N_12103,N_7760,N_7674);
or U12104 (N_12104,N_6723,N_7219);
nor U12105 (N_12105,N_8895,N_6988);
nor U12106 (N_12106,N_8585,N_9239);
or U12107 (N_12107,N_8238,N_8648);
xnor U12108 (N_12108,N_9187,N_9288);
or U12109 (N_12109,N_8770,N_8838);
or U12110 (N_12110,N_7195,N_7440);
or U12111 (N_12111,N_8754,N_7628);
or U12112 (N_12112,N_9256,N_7413);
and U12113 (N_12113,N_9302,N_6363);
xor U12114 (N_12114,N_7065,N_6295);
nand U12115 (N_12115,N_8291,N_7675);
or U12116 (N_12116,N_8871,N_6376);
xnor U12117 (N_12117,N_6706,N_7134);
and U12118 (N_12118,N_7997,N_8416);
or U12119 (N_12119,N_8831,N_6286);
or U12120 (N_12120,N_7057,N_8044);
or U12121 (N_12121,N_7164,N_8855);
nand U12122 (N_12122,N_9061,N_7283);
nand U12123 (N_12123,N_6405,N_8805);
or U12124 (N_12124,N_7120,N_7474);
nor U12125 (N_12125,N_6617,N_6458);
or U12126 (N_12126,N_7046,N_6823);
nor U12127 (N_12127,N_7410,N_6796);
and U12128 (N_12128,N_6339,N_7152);
or U12129 (N_12129,N_8333,N_8453);
xor U12130 (N_12130,N_9331,N_6616);
or U12131 (N_12131,N_8546,N_7810);
and U12132 (N_12132,N_7670,N_7834);
or U12133 (N_12133,N_8701,N_6647);
or U12134 (N_12134,N_8373,N_6387);
nand U12135 (N_12135,N_7095,N_8066);
nor U12136 (N_12136,N_6559,N_7705);
or U12137 (N_12137,N_9267,N_7640);
or U12138 (N_12138,N_8742,N_6794);
nand U12139 (N_12139,N_6546,N_8067);
or U12140 (N_12140,N_7908,N_8935);
nor U12141 (N_12141,N_7727,N_9170);
and U12142 (N_12142,N_8827,N_7255);
or U12143 (N_12143,N_8271,N_7712);
or U12144 (N_12144,N_8766,N_6969);
nor U12145 (N_12145,N_7778,N_7875);
and U12146 (N_12146,N_7824,N_9202);
nor U12147 (N_12147,N_8723,N_6368);
and U12148 (N_12148,N_7867,N_6376);
nor U12149 (N_12149,N_7287,N_8443);
nor U12150 (N_12150,N_7834,N_9011);
nand U12151 (N_12151,N_9085,N_8687);
and U12152 (N_12152,N_7990,N_8316);
nor U12153 (N_12153,N_8498,N_7668);
nor U12154 (N_12154,N_6719,N_8379);
or U12155 (N_12155,N_6276,N_6727);
xnor U12156 (N_12156,N_7645,N_8430);
nand U12157 (N_12157,N_6931,N_9194);
or U12158 (N_12158,N_8258,N_7682);
and U12159 (N_12159,N_8052,N_7198);
nand U12160 (N_12160,N_8115,N_8579);
or U12161 (N_12161,N_8142,N_6918);
or U12162 (N_12162,N_8787,N_9000);
nor U12163 (N_12163,N_8500,N_6764);
nand U12164 (N_12164,N_7264,N_7518);
xor U12165 (N_12165,N_7794,N_8327);
and U12166 (N_12166,N_8263,N_7866);
or U12167 (N_12167,N_6811,N_8264);
nor U12168 (N_12168,N_7580,N_6580);
or U12169 (N_12169,N_6842,N_7256);
or U12170 (N_12170,N_9070,N_9304);
or U12171 (N_12171,N_8002,N_8336);
nor U12172 (N_12172,N_6534,N_9211);
and U12173 (N_12173,N_8334,N_9074);
and U12174 (N_12174,N_6756,N_7499);
nand U12175 (N_12175,N_7748,N_9124);
and U12176 (N_12176,N_8852,N_7430);
or U12177 (N_12177,N_8906,N_7807);
or U12178 (N_12178,N_8565,N_7941);
nand U12179 (N_12179,N_7349,N_9180);
nand U12180 (N_12180,N_7862,N_9156);
or U12181 (N_12181,N_7270,N_7997);
nand U12182 (N_12182,N_8554,N_9020);
nor U12183 (N_12183,N_6707,N_6792);
or U12184 (N_12184,N_6386,N_6596);
or U12185 (N_12185,N_9371,N_8128);
and U12186 (N_12186,N_9327,N_8109);
or U12187 (N_12187,N_8347,N_6885);
nor U12188 (N_12188,N_8450,N_6424);
and U12189 (N_12189,N_9035,N_9267);
and U12190 (N_12190,N_6429,N_7026);
nor U12191 (N_12191,N_6424,N_9122);
or U12192 (N_12192,N_8669,N_8438);
nand U12193 (N_12193,N_8982,N_6646);
nand U12194 (N_12194,N_8943,N_8919);
or U12195 (N_12195,N_8126,N_8296);
nor U12196 (N_12196,N_7756,N_8244);
and U12197 (N_12197,N_8760,N_6365);
nor U12198 (N_12198,N_8447,N_6572);
nor U12199 (N_12199,N_8906,N_9250);
or U12200 (N_12200,N_8805,N_8323);
or U12201 (N_12201,N_8202,N_9361);
or U12202 (N_12202,N_6968,N_9363);
xor U12203 (N_12203,N_8113,N_6724);
and U12204 (N_12204,N_8975,N_8990);
nand U12205 (N_12205,N_7309,N_6777);
or U12206 (N_12206,N_6806,N_7528);
nor U12207 (N_12207,N_8475,N_7370);
nand U12208 (N_12208,N_6622,N_7701);
or U12209 (N_12209,N_8726,N_7067);
nand U12210 (N_12210,N_7329,N_8992);
and U12211 (N_12211,N_8010,N_6531);
nand U12212 (N_12212,N_6626,N_6572);
nand U12213 (N_12213,N_7816,N_8001);
nor U12214 (N_12214,N_6769,N_6890);
and U12215 (N_12215,N_6825,N_8366);
nor U12216 (N_12216,N_7071,N_7731);
or U12217 (N_12217,N_8543,N_7354);
and U12218 (N_12218,N_6566,N_8582);
nand U12219 (N_12219,N_6958,N_8211);
nor U12220 (N_12220,N_8976,N_9234);
nand U12221 (N_12221,N_8131,N_6404);
and U12222 (N_12222,N_7712,N_8187);
or U12223 (N_12223,N_8772,N_7281);
nand U12224 (N_12224,N_8405,N_8433);
and U12225 (N_12225,N_6301,N_7166);
xnor U12226 (N_12226,N_8467,N_6634);
or U12227 (N_12227,N_8840,N_9125);
or U12228 (N_12228,N_8371,N_6653);
and U12229 (N_12229,N_7101,N_6584);
xor U12230 (N_12230,N_8054,N_6384);
and U12231 (N_12231,N_9087,N_6367);
nand U12232 (N_12232,N_9264,N_9238);
and U12233 (N_12233,N_7920,N_7753);
nor U12234 (N_12234,N_6363,N_7547);
or U12235 (N_12235,N_6498,N_8841);
nand U12236 (N_12236,N_7333,N_7202);
and U12237 (N_12237,N_8022,N_6894);
or U12238 (N_12238,N_7345,N_7333);
and U12239 (N_12239,N_9182,N_8644);
and U12240 (N_12240,N_8021,N_9371);
xor U12241 (N_12241,N_7696,N_6826);
nor U12242 (N_12242,N_9328,N_7013);
nor U12243 (N_12243,N_6509,N_7913);
nand U12244 (N_12244,N_7001,N_7689);
nor U12245 (N_12245,N_7091,N_6510);
xnor U12246 (N_12246,N_8349,N_8983);
nor U12247 (N_12247,N_7525,N_8185);
nand U12248 (N_12248,N_8046,N_9263);
nand U12249 (N_12249,N_9141,N_6949);
nand U12250 (N_12250,N_6550,N_6865);
nand U12251 (N_12251,N_8889,N_8295);
nor U12252 (N_12252,N_7778,N_7063);
nand U12253 (N_12253,N_6385,N_9258);
and U12254 (N_12254,N_8541,N_6553);
and U12255 (N_12255,N_9081,N_6412);
nand U12256 (N_12256,N_6495,N_8076);
and U12257 (N_12257,N_8819,N_6650);
or U12258 (N_12258,N_7009,N_7621);
or U12259 (N_12259,N_6472,N_8779);
or U12260 (N_12260,N_7646,N_7410);
nor U12261 (N_12261,N_7684,N_8745);
nor U12262 (N_12262,N_8637,N_9186);
nor U12263 (N_12263,N_9341,N_6423);
nor U12264 (N_12264,N_8704,N_8129);
nor U12265 (N_12265,N_8321,N_7998);
or U12266 (N_12266,N_8446,N_7653);
nor U12267 (N_12267,N_7245,N_8176);
or U12268 (N_12268,N_7977,N_8638);
and U12269 (N_12269,N_7980,N_7344);
and U12270 (N_12270,N_8485,N_8645);
and U12271 (N_12271,N_9207,N_8305);
nand U12272 (N_12272,N_8803,N_6753);
xnor U12273 (N_12273,N_7941,N_7712);
xor U12274 (N_12274,N_8192,N_6855);
nor U12275 (N_12275,N_7892,N_7716);
nand U12276 (N_12276,N_7370,N_6321);
nor U12277 (N_12277,N_9129,N_7062);
and U12278 (N_12278,N_6508,N_6489);
or U12279 (N_12279,N_9114,N_6912);
or U12280 (N_12280,N_6604,N_8289);
nand U12281 (N_12281,N_8504,N_8461);
xnor U12282 (N_12282,N_8801,N_7759);
and U12283 (N_12283,N_8941,N_6666);
and U12284 (N_12284,N_7891,N_7033);
nor U12285 (N_12285,N_9343,N_6472);
and U12286 (N_12286,N_6473,N_8809);
and U12287 (N_12287,N_7577,N_9120);
and U12288 (N_12288,N_7804,N_8628);
xor U12289 (N_12289,N_8111,N_6788);
nor U12290 (N_12290,N_9282,N_6501);
or U12291 (N_12291,N_7031,N_9159);
and U12292 (N_12292,N_7785,N_7961);
and U12293 (N_12293,N_7297,N_8618);
nor U12294 (N_12294,N_6567,N_8202);
or U12295 (N_12295,N_6290,N_6423);
xor U12296 (N_12296,N_8882,N_6789);
or U12297 (N_12297,N_6716,N_8678);
nand U12298 (N_12298,N_8749,N_8386);
and U12299 (N_12299,N_7653,N_8805);
nor U12300 (N_12300,N_7611,N_8448);
or U12301 (N_12301,N_8145,N_6872);
nor U12302 (N_12302,N_8871,N_6588);
nor U12303 (N_12303,N_6600,N_7416);
nor U12304 (N_12304,N_9193,N_7565);
or U12305 (N_12305,N_8377,N_6709);
nand U12306 (N_12306,N_6526,N_8960);
nand U12307 (N_12307,N_8956,N_8376);
nand U12308 (N_12308,N_7325,N_6884);
and U12309 (N_12309,N_6723,N_7615);
and U12310 (N_12310,N_6479,N_9365);
and U12311 (N_12311,N_8813,N_9257);
and U12312 (N_12312,N_9161,N_8677);
and U12313 (N_12313,N_7199,N_9032);
xnor U12314 (N_12314,N_9304,N_8958);
and U12315 (N_12315,N_6593,N_7274);
nor U12316 (N_12316,N_6408,N_7220);
and U12317 (N_12317,N_9357,N_7609);
nor U12318 (N_12318,N_6942,N_6832);
and U12319 (N_12319,N_7324,N_8267);
and U12320 (N_12320,N_7440,N_7115);
and U12321 (N_12321,N_6474,N_8631);
nor U12322 (N_12322,N_7848,N_8235);
and U12323 (N_12323,N_7566,N_6657);
or U12324 (N_12324,N_8945,N_6250);
xor U12325 (N_12325,N_8731,N_7009);
or U12326 (N_12326,N_6914,N_9136);
xor U12327 (N_12327,N_6423,N_7355);
nor U12328 (N_12328,N_8556,N_7479);
nand U12329 (N_12329,N_7606,N_6796);
nor U12330 (N_12330,N_7771,N_9025);
nand U12331 (N_12331,N_8268,N_9237);
nor U12332 (N_12332,N_7635,N_9032);
nand U12333 (N_12333,N_8648,N_6485);
nand U12334 (N_12334,N_8311,N_8194);
nor U12335 (N_12335,N_7706,N_8918);
or U12336 (N_12336,N_7812,N_7937);
nand U12337 (N_12337,N_8101,N_6394);
nand U12338 (N_12338,N_9096,N_7849);
and U12339 (N_12339,N_6917,N_7444);
or U12340 (N_12340,N_7880,N_8801);
nand U12341 (N_12341,N_9002,N_9309);
or U12342 (N_12342,N_6307,N_7183);
xnor U12343 (N_12343,N_8831,N_8346);
nor U12344 (N_12344,N_7454,N_8124);
nor U12345 (N_12345,N_7635,N_7306);
and U12346 (N_12346,N_7042,N_7369);
and U12347 (N_12347,N_7784,N_8720);
nand U12348 (N_12348,N_7021,N_8691);
nand U12349 (N_12349,N_6593,N_8195);
and U12350 (N_12350,N_6459,N_6341);
nand U12351 (N_12351,N_7957,N_7569);
or U12352 (N_12352,N_6676,N_8860);
nor U12353 (N_12353,N_6617,N_7567);
and U12354 (N_12354,N_9344,N_9253);
or U12355 (N_12355,N_7248,N_8322);
or U12356 (N_12356,N_6757,N_6661);
or U12357 (N_12357,N_7297,N_6915);
xnor U12358 (N_12358,N_7450,N_8263);
nand U12359 (N_12359,N_6792,N_7140);
nand U12360 (N_12360,N_8424,N_9234);
or U12361 (N_12361,N_8614,N_7324);
nand U12362 (N_12362,N_9034,N_7652);
or U12363 (N_12363,N_7139,N_8601);
or U12364 (N_12364,N_9133,N_8064);
xor U12365 (N_12365,N_6573,N_8367);
nor U12366 (N_12366,N_8656,N_9041);
nor U12367 (N_12367,N_7362,N_6347);
nand U12368 (N_12368,N_9142,N_8358);
and U12369 (N_12369,N_8741,N_7794);
or U12370 (N_12370,N_7565,N_6965);
nor U12371 (N_12371,N_6505,N_7499);
nand U12372 (N_12372,N_6970,N_8011);
and U12373 (N_12373,N_7660,N_9148);
and U12374 (N_12374,N_6719,N_7882);
and U12375 (N_12375,N_8329,N_8570);
or U12376 (N_12376,N_6424,N_7333);
nand U12377 (N_12377,N_6422,N_8726);
nor U12378 (N_12378,N_6784,N_7411);
nor U12379 (N_12379,N_7489,N_7388);
and U12380 (N_12380,N_7100,N_6504);
or U12381 (N_12381,N_8729,N_7118);
or U12382 (N_12382,N_7010,N_7346);
xor U12383 (N_12383,N_6574,N_7020);
nand U12384 (N_12384,N_8540,N_8218);
nand U12385 (N_12385,N_6414,N_9313);
and U12386 (N_12386,N_6889,N_9206);
and U12387 (N_12387,N_8672,N_7318);
nor U12388 (N_12388,N_6787,N_8108);
nor U12389 (N_12389,N_7908,N_7967);
or U12390 (N_12390,N_8657,N_8487);
nor U12391 (N_12391,N_8529,N_8225);
nand U12392 (N_12392,N_6751,N_9261);
or U12393 (N_12393,N_6942,N_6782);
nor U12394 (N_12394,N_6269,N_6668);
or U12395 (N_12395,N_7209,N_6803);
nor U12396 (N_12396,N_8862,N_6642);
or U12397 (N_12397,N_6465,N_9322);
or U12398 (N_12398,N_7504,N_7578);
or U12399 (N_12399,N_8655,N_7675);
and U12400 (N_12400,N_7457,N_7293);
and U12401 (N_12401,N_8359,N_8411);
and U12402 (N_12402,N_7886,N_6450);
and U12403 (N_12403,N_8922,N_8548);
or U12404 (N_12404,N_8983,N_9162);
nor U12405 (N_12405,N_7361,N_6693);
nand U12406 (N_12406,N_8046,N_9224);
and U12407 (N_12407,N_7663,N_8985);
and U12408 (N_12408,N_8395,N_6697);
and U12409 (N_12409,N_8321,N_8478);
nor U12410 (N_12410,N_7075,N_9043);
xnor U12411 (N_12411,N_8618,N_8975);
nand U12412 (N_12412,N_8029,N_6287);
nor U12413 (N_12413,N_7803,N_7791);
nor U12414 (N_12414,N_8127,N_7270);
nand U12415 (N_12415,N_7597,N_8574);
nand U12416 (N_12416,N_7056,N_7643);
and U12417 (N_12417,N_7758,N_7669);
or U12418 (N_12418,N_6899,N_7388);
nand U12419 (N_12419,N_6587,N_8756);
nor U12420 (N_12420,N_6317,N_8163);
nor U12421 (N_12421,N_8467,N_7863);
and U12422 (N_12422,N_8356,N_6318);
xor U12423 (N_12423,N_7185,N_8661);
or U12424 (N_12424,N_7750,N_7734);
nand U12425 (N_12425,N_6667,N_6252);
nor U12426 (N_12426,N_8616,N_8349);
xnor U12427 (N_12427,N_6448,N_7025);
nand U12428 (N_12428,N_6396,N_8244);
and U12429 (N_12429,N_6753,N_6904);
nand U12430 (N_12430,N_8106,N_8154);
and U12431 (N_12431,N_7085,N_7858);
and U12432 (N_12432,N_8458,N_8694);
nand U12433 (N_12433,N_8167,N_9053);
nand U12434 (N_12434,N_6955,N_8372);
nand U12435 (N_12435,N_6485,N_8602);
nor U12436 (N_12436,N_8615,N_6778);
nand U12437 (N_12437,N_8815,N_8754);
nand U12438 (N_12438,N_7507,N_8589);
or U12439 (N_12439,N_6536,N_8775);
nor U12440 (N_12440,N_8079,N_6316);
or U12441 (N_12441,N_8573,N_8645);
nor U12442 (N_12442,N_7779,N_7039);
or U12443 (N_12443,N_9313,N_6697);
nor U12444 (N_12444,N_6907,N_6888);
nand U12445 (N_12445,N_6631,N_6734);
or U12446 (N_12446,N_8225,N_8004);
xnor U12447 (N_12447,N_6632,N_8883);
and U12448 (N_12448,N_7874,N_6596);
nor U12449 (N_12449,N_9363,N_6729);
xnor U12450 (N_12450,N_7605,N_8750);
or U12451 (N_12451,N_7475,N_8845);
or U12452 (N_12452,N_7060,N_9140);
or U12453 (N_12453,N_7751,N_7749);
xor U12454 (N_12454,N_6921,N_7297);
and U12455 (N_12455,N_6862,N_7324);
or U12456 (N_12456,N_6373,N_7490);
and U12457 (N_12457,N_8149,N_8992);
nand U12458 (N_12458,N_8750,N_7135);
nand U12459 (N_12459,N_9059,N_8870);
and U12460 (N_12460,N_7078,N_7346);
and U12461 (N_12461,N_8217,N_8193);
nand U12462 (N_12462,N_8833,N_8656);
or U12463 (N_12463,N_9044,N_7262);
nor U12464 (N_12464,N_8699,N_7096);
nor U12465 (N_12465,N_7733,N_8134);
and U12466 (N_12466,N_6398,N_6764);
and U12467 (N_12467,N_6558,N_6984);
nand U12468 (N_12468,N_6574,N_8936);
nor U12469 (N_12469,N_6291,N_7232);
or U12470 (N_12470,N_7417,N_7041);
nand U12471 (N_12471,N_7442,N_8925);
xor U12472 (N_12472,N_7283,N_7032);
nor U12473 (N_12473,N_8142,N_8584);
nor U12474 (N_12474,N_8688,N_6994);
nand U12475 (N_12475,N_8901,N_7419);
nor U12476 (N_12476,N_8552,N_6869);
nand U12477 (N_12477,N_6664,N_7511);
nand U12478 (N_12478,N_7098,N_7384);
and U12479 (N_12479,N_6910,N_8224);
or U12480 (N_12480,N_6588,N_7014);
and U12481 (N_12481,N_9016,N_9333);
nor U12482 (N_12482,N_9187,N_8624);
and U12483 (N_12483,N_8770,N_6386);
and U12484 (N_12484,N_7015,N_8260);
nor U12485 (N_12485,N_8780,N_9077);
or U12486 (N_12486,N_6987,N_8606);
and U12487 (N_12487,N_8158,N_7256);
xnor U12488 (N_12488,N_7075,N_6542);
nand U12489 (N_12489,N_9087,N_8025);
xnor U12490 (N_12490,N_7191,N_9150);
nor U12491 (N_12491,N_6475,N_7130);
nor U12492 (N_12492,N_7187,N_9165);
xor U12493 (N_12493,N_7579,N_8053);
xnor U12494 (N_12494,N_6989,N_8655);
xor U12495 (N_12495,N_7273,N_7010);
or U12496 (N_12496,N_8113,N_8203);
xnor U12497 (N_12497,N_8527,N_8062);
nand U12498 (N_12498,N_7782,N_8813);
nor U12499 (N_12499,N_6582,N_8472);
xor U12500 (N_12500,N_11055,N_10610);
nor U12501 (N_12501,N_12232,N_11214);
xor U12502 (N_12502,N_10285,N_11054);
nand U12503 (N_12503,N_11928,N_10094);
nand U12504 (N_12504,N_11243,N_10740);
nand U12505 (N_12505,N_10977,N_10962);
and U12506 (N_12506,N_11517,N_10246);
and U12507 (N_12507,N_9703,N_12416);
or U12508 (N_12508,N_11232,N_11339);
nand U12509 (N_12509,N_10053,N_12068);
nor U12510 (N_12510,N_10098,N_11516);
and U12511 (N_12511,N_12472,N_12222);
nand U12512 (N_12512,N_11707,N_12059);
and U12513 (N_12513,N_9831,N_10140);
xnor U12514 (N_12514,N_10825,N_10444);
nor U12515 (N_12515,N_10580,N_12090);
nor U12516 (N_12516,N_9524,N_10671);
and U12517 (N_12517,N_9784,N_10733);
and U12518 (N_12518,N_10250,N_10472);
nor U12519 (N_12519,N_10205,N_9931);
nand U12520 (N_12520,N_10649,N_10142);
and U12521 (N_12521,N_10223,N_11894);
nand U12522 (N_12522,N_12364,N_9755);
and U12523 (N_12523,N_10373,N_10229);
nand U12524 (N_12524,N_11669,N_11605);
nand U12525 (N_12525,N_10691,N_10305);
nand U12526 (N_12526,N_11804,N_12430);
nor U12527 (N_12527,N_11245,N_9471);
and U12528 (N_12528,N_10522,N_11515);
xnor U12529 (N_12529,N_12259,N_9624);
nand U12530 (N_12530,N_9453,N_9674);
and U12531 (N_12531,N_12077,N_10040);
and U12532 (N_12532,N_9950,N_11814);
nor U12533 (N_12533,N_11832,N_10923);
or U12534 (N_12534,N_10348,N_9615);
and U12535 (N_12535,N_9846,N_10490);
or U12536 (N_12536,N_10982,N_12214);
nor U12537 (N_12537,N_11174,N_9722);
nand U12538 (N_12538,N_10259,N_11029);
or U12539 (N_12539,N_12372,N_10380);
nor U12540 (N_12540,N_11428,N_10203);
nand U12541 (N_12541,N_9810,N_10817);
nor U12542 (N_12542,N_12235,N_11062);
or U12543 (N_12543,N_12443,N_11385);
and U12544 (N_12544,N_9893,N_10949);
nor U12545 (N_12545,N_11848,N_10861);
nor U12546 (N_12546,N_11246,N_12124);
xnor U12547 (N_12547,N_12081,N_10614);
and U12548 (N_12548,N_12027,N_9886);
or U12549 (N_12549,N_10020,N_9751);
nor U12550 (N_12550,N_10720,N_10448);
and U12551 (N_12551,N_10736,N_10811);
nand U12552 (N_12552,N_10968,N_11914);
and U12553 (N_12553,N_12127,N_12265);
xor U12554 (N_12554,N_11336,N_10168);
or U12555 (N_12555,N_10376,N_9616);
or U12556 (N_12556,N_9861,N_9550);
and U12557 (N_12557,N_9654,N_11315);
or U12558 (N_12558,N_11985,N_11125);
and U12559 (N_12559,N_12038,N_9957);
nor U12560 (N_12560,N_10925,N_11744);
and U12561 (N_12561,N_11291,N_12238);
nand U12562 (N_12562,N_9902,N_10676);
or U12563 (N_12563,N_10821,N_10441);
nor U12564 (N_12564,N_10104,N_9948);
or U12565 (N_12565,N_12340,N_9705);
or U12566 (N_12566,N_9862,N_12107);
nor U12567 (N_12567,N_10848,N_12114);
nor U12568 (N_12568,N_12035,N_11788);
nor U12569 (N_12569,N_9586,N_12278);
and U12570 (N_12570,N_9603,N_9549);
nor U12571 (N_12571,N_11687,N_11645);
nand U12572 (N_12572,N_10775,N_10976);
xor U12573 (N_12573,N_9590,N_10129);
or U12574 (N_12574,N_10728,N_12036);
or U12575 (N_12575,N_11564,N_10113);
and U12576 (N_12576,N_12078,N_11553);
xnor U12577 (N_12577,N_9546,N_11791);
nor U12578 (N_12578,N_10661,N_12147);
nor U12579 (N_12579,N_10716,N_11922);
nor U12580 (N_12580,N_9439,N_10729);
or U12581 (N_12581,N_12141,N_10902);
or U12582 (N_12582,N_10268,N_11492);
nand U12583 (N_12583,N_11462,N_10572);
nor U12584 (N_12584,N_12252,N_11453);
nor U12585 (N_12585,N_10605,N_11854);
nand U12586 (N_12586,N_11407,N_12311);
and U12587 (N_12587,N_9564,N_12013);
or U12588 (N_12588,N_11562,N_10946);
and U12589 (N_12589,N_9860,N_10469);
or U12590 (N_12590,N_9462,N_10742);
or U12591 (N_12591,N_11878,N_10571);
nor U12592 (N_12592,N_10018,N_10263);
and U12593 (N_12593,N_11548,N_12272);
nand U12594 (N_12594,N_12125,N_10764);
and U12595 (N_12595,N_10627,N_11745);
and U12596 (N_12596,N_9881,N_11676);
and U12597 (N_12597,N_11499,N_9608);
nor U12598 (N_12598,N_12053,N_12057);
and U12599 (N_12599,N_10478,N_10758);
nand U12600 (N_12600,N_11983,N_11488);
and U12601 (N_12601,N_9850,N_11699);
nor U12602 (N_12602,N_11239,N_12434);
or U12603 (N_12603,N_12387,N_12312);
or U12604 (N_12604,N_10843,N_9528);
nand U12605 (N_12605,N_10032,N_12096);
nor U12606 (N_12606,N_10783,N_10896);
xor U12607 (N_12607,N_11066,N_9620);
nor U12608 (N_12608,N_12220,N_11594);
nand U12609 (N_12609,N_11166,N_11793);
nor U12610 (N_12610,N_10646,N_11325);
xor U12611 (N_12611,N_11240,N_12492);
and U12612 (N_12612,N_12136,N_11244);
and U12613 (N_12613,N_11588,N_11609);
and U12614 (N_12614,N_11004,N_12483);
and U12615 (N_12615,N_11368,N_12155);
nor U12616 (N_12616,N_9712,N_10533);
nor U12617 (N_12617,N_10501,N_9801);
nor U12618 (N_12618,N_11843,N_11184);
xnor U12619 (N_12619,N_11220,N_9949);
nand U12620 (N_12620,N_10678,N_11003);
nor U12621 (N_12621,N_12007,N_12242);
nand U12622 (N_12622,N_11427,N_10143);
and U12623 (N_12623,N_12411,N_12092);
or U12624 (N_12624,N_12052,N_11082);
or U12625 (N_12625,N_9644,N_11680);
nor U12626 (N_12626,N_11992,N_9976);
and U12627 (N_12627,N_11803,N_9568);
nand U12628 (N_12628,N_11432,N_11704);
or U12629 (N_12629,N_10064,N_11312);
nor U12630 (N_12630,N_9899,N_11413);
or U12631 (N_12631,N_9570,N_11394);
nand U12632 (N_12632,N_9464,N_11895);
and U12633 (N_12633,N_9660,N_12054);
nand U12634 (N_12634,N_11995,N_11752);
nand U12635 (N_12635,N_11307,N_11048);
nand U12636 (N_12636,N_9484,N_10643);
nand U12637 (N_12637,N_10264,N_11450);
nand U12638 (N_12638,N_11287,N_9809);
nor U12639 (N_12639,N_10166,N_10051);
xnor U12640 (N_12640,N_10419,N_9786);
nand U12641 (N_12641,N_11087,N_11402);
and U12642 (N_12642,N_11648,N_12412);
xor U12643 (N_12643,N_9687,N_9494);
nand U12644 (N_12644,N_10632,N_11792);
nand U12645 (N_12645,N_11417,N_12117);
nand U12646 (N_12646,N_10206,N_11389);
nand U12647 (N_12647,N_11891,N_9972);
and U12648 (N_12648,N_10541,N_10761);
nor U12649 (N_12649,N_11716,N_11067);
and U12650 (N_12650,N_11002,N_11070);
or U12651 (N_12651,N_12354,N_9719);
nand U12652 (N_12652,N_10629,N_11856);
or U12653 (N_12653,N_11145,N_11433);
and U12654 (N_12654,N_11836,N_10395);
and U12655 (N_12655,N_9691,N_11206);
nor U12656 (N_12656,N_12407,N_9921);
and U12657 (N_12657,N_9804,N_10437);
nor U12658 (N_12658,N_10391,N_10705);
nor U12659 (N_12659,N_9587,N_9658);
and U12660 (N_12660,N_10745,N_12329);
nor U12661 (N_12661,N_12029,N_10901);
and U12662 (N_12662,N_9710,N_12271);
nor U12663 (N_12663,N_12269,N_9576);
or U12664 (N_12664,N_10456,N_11655);
nand U12665 (N_12665,N_10272,N_11016);
or U12666 (N_12666,N_12234,N_10226);
and U12667 (N_12667,N_9432,N_11712);
or U12668 (N_12668,N_9688,N_11300);
nor U12669 (N_12669,N_11491,N_9456);
nor U12670 (N_12670,N_10835,N_11794);
nor U12671 (N_12671,N_9694,N_11835);
xor U12672 (N_12672,N_10193,N_11105);
nor U12673 (N_12673,N_10396,N_9451);
or U12674 (N_12674,N_12086,N_12110);
and U12675 (N_12675,N_12489,N_11481);
nand U12676 (N_12676,N_12142,N_9589);
nand U12677 (N_12677,N_10583,N_9509);
and U12678 (N_12678,N_9492,N_11601);
and U12679 (N_12679,N_12264,N_9868);
and U12680 (N_12680,N_10220,N_12305);
nand U12681 (N_12681,N_11510,N_12184);
nor U12682 (N_12682,N_9676,N_10006);
nand U12683 (N_12683,N_10043,N_11121);
nor U12684 (N_12684,N_9695,N_10439);
or U12685 (N_12685,N_9942,N_9463);
or U12686 (N_12686,N_11350,N_9853);
or U12687 (N_12687,N_10471,N_12453);
nor U12688 (N_12688,N_11474,N_9521);
nand U12689 (N_12689,N_10608,N_11069);
or U12690 (N_12690,N_12008,N_10859);
or U12691 (N_12691,N_10485,N_11997);
or U12692 (N_12692,N_11839,N_12386);
and U12693 (N_12693,N_11821,N_11153);
nand U12694 (N_12694,N_10074,N_10339);
xor U12695 (N_12695,N_10567,N_11572);
nand U12696 (N_12696,N_9681,N_11301);
nand U12697 (N_12697,N_10219,N_11137);
nand U12698 (N_12698,N_10238,N_10057);
xor U12699 (N_12699,N_11973,N_9789);
nor U12700 (N_12700,N_11127,N_11028);
or U12701 (N_12701,N_9736,N_10634);
or U12702 (N_12702,N_11074,N_9882);
and U12703 (N_12703,N_11392,N_12026);
nand U12704 (N_12704,N_9523,N_11840);
xor U12705 (N_12705,N_12320,N_11809);
nand U12706 (N_12706,N_11104,N_9655);
nand U12707 (N_12707,N_9962,N_11855);
nor U12708 (N_12708,N_12009,N_12162);
or U12709 (N_12709,N_12274,N_9870);
nand U12710 (N_12710,N_10039,N_9380);
nor U12711 (N_12711,N_11059,N_9411);
nand U12712 (N_12712,N_12337,N_10969);
nand U12713 (N_12713,N_9738,N_12318);
and U12714 (N_12714,N_11807,N_11468);
nand U12715 (N_12715,N_12229,N_11092);
and U12716 (N_12716,N_9662,N_10653);
and U12717 (N_12717,N_12176,N_10335);
and U12718 (N_12718,N_11838,N_11719);
xnor U12719 (N_12719,N_10695,N_9917);
or U12720 (N_12720,N_10804,N_12352);
or U12721 (N_12721,N_11302,N_11767);
nor U12722 (N_12722,N_9930,N_9622);
nand U12723 (N_12723,N_12039,N_9639);
nand U12724 (N_12724,N_12332,N_12341);
and U12725 (N_12725,N_11318,N_12042);
or U12726 (N_12726,N_11257,N_9901);
or U12727 (N_12727,N_10640,N_11532);
and U12728 (N_12728,N_9437,N_10465);
nor U12729 (N_12729,N_11361,N_9826);
or U12730 (N_12730,N_11916,N_12335);
and U12731 (N_12731,N_9565,N_10814);
nor U12732 (N_12732,N_10987,N_9728);
and U12733 (N_12733,N_9443,N_9878);
xnor U12734 (N_12734,N_11329,N_10528);
nand U12735 (N_12735,N_11176,N_9726);
or U12736 (N_12736,N_9645,N_11483);
xnor U12737 (N_12737,N_10385,N_11443);
nor U12738 (N_12738,N_11365,N_11774);
nor U12739 (N_12739,N_10199,N_10026);
or U12740 (N_12740,N_10382,N_11178);
and U12741 (N_12741,N_9702,N_9979);
nand U12742 (N_12742,N_11150,N_11924);
xnor U12743 (N_12743,N_11424,N_10686);
or U12744 (N_12744,N_12304,N_12206);
xnor U12745 (N_12745,N_11090,N_12058);
xor U12746 (N_12746,N_12034,N_11489);
or U12747 (N_12747,N_11177,N_9839);
and U12748 (N_12748,N_12446,N_11260);
nand U12749 (N_12749,N_9536,N_10275);
nand U12750 (N_12750,N_9937,N_11871);
or U12751 (N_12751,N_12384,N_11640);
or U12752 (N_12752,N_11700,N_9994);
nor U12753 (N_12753,N_10809,N_9659);
or U12754 (N_12754,N_10412,N_9892);
and U12755 (N_12755,N_10169,N_10494);
nor U12756 (N_12756,N_10590,N_10990);
nor U12757 (N_12757,N_11446,N_11396);
and U12758 (N_12758,N_10971,N_9621);
nor U12759 (N_12759,N_12202,N_11103);
and U12760 (N_12760,N_9522,N_11768);
and U12761 (N_12761,N_11210,N_9713);
and U12762 (N_12762,N_10450,N_9808);
or U12763 (N_12763,N_11412,N_11136);
xnor U12764 (N_12764,N_10972,N_9584);
nor U12765 (N_12765,N_9821,N_12452);
nand U12766 (N_12766,N_9602,N_12357);
nand U12767 (N_12767,N_10210,N_11162);
nor U12768 (N_12768,N_11207,N_12098);
and U12769 (N_12769,N_12198,N_12313);
and U12770 (N_12770,N_12243,N_10111);
and U12771 (N_12771,N_11383,N_12070);
or U12772 (N_12772,N_10449,N_11847);
nand U12773 (N_12773,N_11954,N_10133);
nand U12774 (N_12774,N_10822,N_10674);
and U12775 (N_12775,N_11606,N_10888);
and U12776 (N_12776,N_10016,N_11868);
nand U12777 (N_12777,N_11806,N_10072);
or U12778 (N_12778,N_9428,N_10144);
and U12779 (N_12779,N_10876,N_10989);
and U12780 (N_12780,N_11343,N_11487);
and U12781 (N_12781,N_11098,N_11650);
nand U12782 (N_12782,N_11739,N_10668);
and U12783 (N_12783,N_10134,N_9844);
and U12784 (N_12784,N_11918,N_11330);
xnor U12785 (N_12785,N_10442,N_10036);
nor U12786 (N_12786,N_10916,N_11490);
nor U12787 (N_12787,N_10165,N_10840);
or U12788 (N_12788,N_11935,N_12431);
nand U12789 (N_12789,N_10935,N_10007);
and U12790 (N_12790,N_12191,N_10179);
nor U12791 (N_12791,N_9704,N_10746);
and U12792 (N_12792,N_10289,N_12379);
or U12793 (N_12793,N_10737,N_10340);
and U12794 (N_12794,N_11026,N_10953);
nand U12795 (N_12795,N_10027,N_10941);
nor U12796 (N_12796,N_11106,N_12010);
nand U12797 (N_12797,N_11933,N_11820);
or U12798 (N_12798,N_10857,N_12094);
or U12799 (N_12799,N_10910,N_12132);
nand U12800 (N_12800,N_10407,N_11231);
nor U12801 (N_12801,N_10197,N_10452);
and U12802 (N_12802,N_9407,N_10510);
xnor U12803 (N_12803,N_9747,N_11981);
and U12804 (N_12804,N_12177,N_11036);
nor U12805 (N_12805,N_9383,N_10535);
and U12806 (N_12806,N_11540,N_10578);
and U12807 (N_12807,N_12396,N_11377);
and U12808 (N_12808,N_10358,N_9904);
nand U12809 (N_12809,N_10300,N_11375);
and U12810 (N_12810,N_12093,N_12398);
nor U12811 (N_12811,N_11438,N_10586);
nand U12812 (N_12812,N_12064,N_9740);
nand U12813 (N_12813,N_12056,N_10080);
and U12814 (N_12814,N_11958,N_10406);
and U12815 (N_12815,N_11826,N_10473);
nor U12816 (N_12816,N_10877,N_11175);
xor U12817 (N_12817,N_10195,N_10790);
or U12818 (N_12818,N_11094,N_9470);
or U12819 (N_12819,N_10481,N_9806);
nand U12820 (N_12820,N_9377,N_9968);
nor U12821 (N_12821,N_10292,N_9395);
nor U12822 (N_12822,N_11400,N_11721);
or U12823 (N_12823,N_12122,N_10757);
nand U12824 (N_12824,N_9743,N_11547);
or U12825 (N_12825,N_9653,N_9647);
or U12826 (N_12826,N_10069,N_11544);
and U12827 (N_12827,N_11447,N_12374);
or U12828 (N_12828,N_10823,N_12046);
nor U12829 (N_12829,N_10905,N_9579);
or U12830 (N_12830,N_12217,N_11277);
nand U12831 (N_12831,N_9563,N_11577);
or U12832 (N_12832,N_11116,N_9975);
nor U12833 (N_12833,N_9742,N_10805);
nor U12834 (N_12834,N_11999,N_10170);
and U12835 (N_12835,N_11164,N_11114);
nor U12836 (N_12836,N_9573,N_12321);
nor U12837 (N_12837,N_10834,N_11404);
or U12838 (N_12838,N_10333,N_11506);
nand U12839 (N_12839,N_12164,N_12148);
or U12840 (N_12840,N_12245,N_10324);
xnor U12841 (N_12841,N_12392,N_11494);
nand U12842 (N_12842,N_12371,N_11242);
nor U12843 (N_12843,N_10779,N_11616);
nand U12844 (N_12844,N_11274,N_11118);
nand U12845 (N_12845,N_10271,N_10756);
and U12846 (N_12846,N_12248,N_11571);
or U12847 (N_12847,N_9956,N_9765);
or U12848 (N_12848,N_10438,N_9544);
and U12849 (N_12849,N_12351,N_11147);
and U12850 (N_12850,N_11022,N_9900);
nor U12851 (N_12851,N_11551,N_11041);
nor U12852 (N_12852,N_12095,N_12400);
xnor U12853 (N_12853,N_10694,N_12133);
nand U12854 (N_12854,N_10401,N_10994);
and U12855 (N_12855,N_10393,N_10409);
or U12856 (N_12856,N_9852,N_10236);
and U12857 (N_12857,N_11927,N_11952);
nor U12858 (N_12858,N_9454,N_11187);
nand U12859 (N_12859,N_10100,N_10024);
nand U12860 (N_12860,N_10904,N_10284);
nand U12861 (N_12861,N_11853,N_12152);
and U12862 (N_12862,N_9397,N_11158);
nand U12863 (N_12863,N_12294,N_11442);
nand U12864 (N_12864,N_11382,N_11469);
nor U12865 (N_12865,N_11485,N_12385);
nand U12866 (N_12866,N_11449,N_11073);
or U12867 (N_12867,N_12426,N_9610);
nor U12868 (N_12868,N_9720,N_10417);
or U12869 (N_12869,N_9535,N_10664);
xor U12870 (N_12870,N_10044,N_10164);
nand U12871 (N_12871,N_9698,N_11844);
xor U12872 (N_12872,N_9538,N_10042);
nand U12873 (N_12873,N_10266,N_11414);
nor U12874 (N_12874,N_10907,N_11720);
nor U12875 (N_12875,N_12395,N_12113);
or U12876 (N_12876,N_11578,N_12241);
and U12877 (N_12877,N_11355,N_9585);
nand U12878 (N_12878,N_10176,N_10747);
or U12879 (N_12879,N_10727,N_10555);
and U12880 (N_12880,N_12498,N_9954);
or U12881 (N_12881,N_10546,N_11582);
or U12882 (N_12882,N_11725,N_12282);
nand U12883 (N_12883,N_9391,N_12486);
xnor U12884 (N_12884,N_11511,N_10611);
and U12885 (N_12885,N_11634,N_11144);
xnor U12886 (N_12886,N_12106,N_10301);
nor U12887 (N_12887,N_10315,N_10493);
nand U12888 (N_12888,N_11141,N_11949);
xor U12889 (N_12889,N_9512,N_10280);
or U12890 (N_12890,N_9444,N_11647);
or U12891 (N_12891,N_10019,N_10988);
or U12892 (N_12892,N_11403,N_9706);
nand U12893 (N_12893,N_9918,N_10075);
or U12894 (N_12894,N_9431,N_11126);
and U12895 (N_12895,N_12424,N_10936);
or U12896 (N_12896,N_12073,N_9537);
or U12897 (N_12897,N_10371,N_11917);
or U12898 (N_12898,N_12270,N_11133);
nor U12899 (N_12899,N_10225,N_11146);
nand U12900 (N_12900,N_10628,N_11892);
xnor U12901 (N_12901,N_9863,N_12401);
xnor U12902 (N_12902,N_12240,N_12233);
or U12903 (N_12903,N_11563,N_11520);
nor U12904 (N_12904,N_10648,N_9982);
xnor U12905 (N_12905,N_10189,N_10601);
and U12906 (N_12906,N_10852,N_11991);
nor U12907 (N_12907,N_9941,N_9630);
nor U12908 (N_12908,N_11670,N_11216);
and U12909 (N_12909,N_9559,N_11970);
nand U12910 (N_12910,N_12017,N_11685);
nor U12911 (N_12911,N_11632,N_12327);
nor U12912 (N_12912,N_10314,N_11049);
or U12913 (N_12913,N_10878,N_12018);
nor U12914 (N_12914,N_10302,N_12139);
or U12915 (N_12915,N_12465,N_10318);
nor U12916 (N_12916,N_11526,N_11851);
nand U12917 (N_12917,N_10791,N_10119);
nor U12918 (N_12918,N_11599,N_11600);
and U12919 (N_12919,N_11677,N_10174);
nor U12920 (N_12920,N_9682,N_11730);
xnor U12921 (N_12921,N_9668,N_11160);
nand U12922 (N_12922,N_11931,N_10418);
nand U12923 (N_12923,N_10589,N_11975);
xnor U12924 (N_12924,N_10090,N_9502);
or U12925 (N_12925,N_11321,N_11537);
and U12926 (N_12926,N_9516,N_10196);
nor U12927 (N_12927,N_10577,N_9527);
nand U12928 (N_12928,N_9803,N_11619);
or U12929 (N_12929,N_10921,N_12181);
nand U12930 (N_12930,N_11095,N_9788);
or U12931 (N_12931,N_9636,N_12299);
nor U12932 (N_12932,N_10230,N_12474);
nor U12933 (N_12933,N_10596,N_9888);
nor U12934 (N_12934,N_11038,N_9947);
nor U12935 (N_12935,N_9452,N_9539);
nand U12936 (N_12936,N_12196,N_10730);
xor U12937 (N_12937,N_11278,N_10986);
or U12938 (N_12938,N_10451,N_9842);
nor U12939 (N_12939,N_10741,N_10354);
nand U12940 (N_12940,N_9776,N_10291);
nand U12941 (N_12941,N_9390,N_10491);
and U12942 (N_12942,N_11765,N_11759);
nand U12943 (N_12943,N_11566,N_10841);
or U12944 (N_12944,N_12347,N_11584);
nand U12945 (N_12945,N_10508,N_11248);
and U12946 (N_12946,N_10212,N_11282);
or U12947 (N_12947,N_11271,N_11238);
nand U12948 (N_12948,N_11697,N_12150);
and U12949 (N_12949,N_10998,N_10184);
or U12950 (N_12950,N_11255,N_11051);
nand U12951 (N_12951,N_10265,N_10117);
nor U12952 (N_12952,N_11689,N_10709);
or U12953 (N_12953,N_12065,N_10479);
nor U12954 (N_12954,N_11679,N_12464);
xor U12955 (N_12955,N_10795,N_9696);
nor U12956 (N_12956,N_10922,N_9959);
nand U12957 (N_12957,N_12447,N_9382);
nor U12958 (N_12958,N_11696,N_10233);
nand U12959 (N_12959,N_10152,N_9914);
xor U12960 (N_12960,N_11273,N_9910);
nor U12961 (N_12961,N_10581,N_12130);
and U12962 (N_12962,N_12211,N_11131);
nor U12963 (N_12963,N_11415,N_12307);
nand U12964 (N_12964,N_10415,N_12149);
and U12965 (N_12965,N_10552,N_11876);
or U12966 (N_12966,N_12210,N_10514);
and U12967 (N_12967,N_9699,N_9820);
nand U12968 (N_12968,N_9683,N_11139);
or U12969 (N_12969,N_11501,N_12288);
or U12970 (N_12970,N_11615,N_11308);
nand U12971 (N_12971,N_10194,N_9828);
and U12972 (N_12972,N_12230,N_9907);
and U12973 (N_12973,N_11093,N_12137);
xor U12974 (N_12974,N_9673,N_10869);
nand U12975 (N_12975,N_11340,N_10365);
nor U12976 (N_12976,N_9774,N_12193);
nor U12977 (N_12977,N_11561,N_12302);
and U12978 (N_12978,N_12308,N_11861);
or U12979 (N_12979,N_10311,N_11456);
or U12980 (N_12980,N_11173,N_9697);
nand U12981 (N_12981,N_11285,N_11284);
or U12982 (N_12982,N_11581,N_10298);
or U12983 (N_12983,N_10784,N_11665);
xor U12984 (N_12984,N_11595,N_10862);
or U12985 (N_12985,N_10631,N_11218);
xnor U12986 (N_12986,N_12239,N_9598);
or U12987 (N_12987,N_9986,N_11208);
xnor U12988 (N_12988,N_10929,N_11496);
and U12989 (N_12989,N_12273,N_12151);
and U12990 (N_12990,N_9834,N_9671);
nor U12991 (N_12991,N_11171,N_12279);
and U12992 (N_12992,N_11755,N_10978);
and U12993 (N_12993,N_10351,N_12365);
nand U12994 (N_12994,N_11692,N_10489);
nor U12995 (N_12995,N_11068,N_9777);
and U12996 (N_12996,N_10132,N_11165);
and U12997 (N_12997,N_10269,N_12298);
nor U12998 (N_12998,N_9396,N_11811);
and U12999 (N_12999,N_10037,N_10744);
or U13000 (N_13000,N_9560,N_10181);
xor U13001 (N_13001,N_10553,N_9686);
nand U13002 (N_13002,N_11624,N_11631);
nand U13003 (N_13003,N_9417,N_11653);
nor U13004 (N_13004,N_9430,N_11734);
or U13005 (N_13005,N_11738,N_9542);
and U13006 (N_13006,N_10509,N_9420);
nor U13007 (N_13007,N_9811,N_12226);
or U13008 (N_13008,N_10531,N_9997);
and U13009 (N_13009,N_12268,N_11117);
nor U13010 (N_13010,N_11824,N_12022);
or U13011 (N_13011,N_10537,N_11128);
nor U13012 (N_13012,N_11743,N_10874);
nor U13013 (N_13013,N_10984,N_11541);
nor U13014 (N_13014,N_10828,N_10077);
or U13015 (N_13015,N_11817,N_12195);
or U13016 (N_13016,N_12487,N_11495);
nor U13017 (N_13017,N_9505,N_9468);
and U13018 (N_13018,N_11124,N_12071);
and U13019 (N_13019,N_9423,N_10711);
or U13020 (N_13020,N_10310,N_10663);
nand U13021 (N_13021,N_10378,N_11639);
or U13022 (N_13022,N_11188,N_9379);
nor U13023 (N_13023,N_11316,N_10127);
and U13024 (N_13024,N_12397,N_12303);
xor U13025 (N_13025,N_12420,N_9898);
xor U13026 (N_13026,N_10966,N_12192);
and U13027 (N_13027,N_10930,N_10534);
nor U13028 (N_13028,N_10260,N_11464);
nor U13029 (N_13029,N_11152,N_10476);
xnor U13030 (N_13030,N_10009,N_10356);
or U13031 (N_13031,N_10947,N_12345);
nor U13032 (N_13032,N_12246,N_12209);
and U13033 (N_13033,N_11182,N_10898);
or U13034 (N_13034,N_10996,N_11912);
and U13035 (N_13035,N_11452,N_12348);
and U13036 (N_13036,N_9447,N_11702);
or U13037 (N_13037,N_11948,N_10216);
nand U13038 (N_13038,N_11324,N_11295);
xnor U13039 (N_13039,N_9984,N_10543);
xnor U13040 (N_13040,N_10279,N_12413);
nor U13041 (N_13041,N_11875,N_12389);
and U13042 (N_13042,N_9499,N_9729);
nor U13043 (N_13043,N_11352,N_11185);
or U13044 (N_13044,N_11422,N_10700);
or U13045 (N_13045,N_10463,N_9562);
or U13046 (N_13046,N_12445,N_9378);
nor U13047 (N_13047,N_11980,N_11270);
nor U13048 (N_13048,N_9857,N_10486);
and U13049 (N_13049,N_11134,N_11327);
nor U13050 (N_13050,N_10499,N_10374);
or U13051 (N_13051,N_12250,N_11052);
nand U13052 (N_13052,N_10985,N_9778);
nor U13053 (N_13053,N_12091,N_10002);
nor U13054 (N_13054,N_11405,N_11348);
or U13055 (N_13055,N_9435,N_10124);
and U13056 (N_13056,N_9990,N_12194);
or U13057 (N_13057,N_10171,N_9386);
nor U13058 (N_13058,N_9648,N_11694);
and U13059 (N_13059,N_10445,N_11286);
nand U13060 (N_13060,N_11570,N_9814);
nand U13061 (N_13061,N_10278,N_11550);
xnor U13062 (N_13062,N_12309,N_10123);
nand U13063 (N_13063,N_10453,N_12167);
xor U13064 (N_13064,N_10958,N_10658);
xor U13065 (N_13065,N_11842,N_11907);
or U13066 (N_13066,N_10765,N_11132);
xor U13067 (N_13067,N_11191,N_9650);
nand U13068 (N_13068,N_9519,N_11810);
or U13069 (N_13069,N_11603,N_12494);
and U13070 (N_13070,N_11431,N_11310);
xor U13071 (N_13071,N_12383,N_9469);
nor U13072 (N_13072,N_10525,N_9812);
xor U13073 (N_13073,N_10725,N_12200);
and U13074 (N_13074,N_9413,N_12323);
xnor U13075 (N_13075,N_11683,N_9830);
or U13076 (N_13076,N_11586,N_11642);
or U13077 (N_13077,N_11251,N_11014);
xor U13078 (N_13078,N_11040,N_10515);
and U13079 (N_13079,N_11910,N_11249);
or U13080 (N_13080,N_9800,N_9714);
nand U13081 (N_13081,N_11622,N_10997);
nor U13082 (N_13082,N_10781,N_11227);
nor U13083 (N_13083,N_10529,N_11486);
nor U13084 (N_13084,N_9932,N_11183);
nand U13085 (N_13085,N_11633,N_11845);
and U13086 (N_13086,N_10810,N_10008);
or U13087 (N_13087,N_9394,N_10030);
xnor U13088 (N_13088,N_10576,N_12484);
nor U13089 (N_13089,N_9780,N_12461);
and U13090 (N_13090,N_9618,N_10214);
and U13091 (N_13091,N_11559,N_10294);
nor U13092 (N_13092,N_11370,N_9466);
nand U13093 (N_13093,N_10198,N_12173);
or U13094 (N_13094,N_11120,N_10719);
and U13095 (N_13095,N_11941,N_10480);
and U13096 (N_13096,N_10244,N_11053);
or U13097 (N_13097,N_10866,N_9879);
or U13098 (N_13098,N_9582,N_9511);
nor U13099 (N_13099,N_9547,N_11957);
nand U13100 (N_13100,N_11773,N_11723);
and U13101 (N_13101,N_12450,N_12203);
nand U13102 (N_13102,N_10322,N_9406);
xnor U13103 (N_13103,N_12119,N_11391);
xor U13104 (N_13104,N_12123,N_11859);
nand U13105 (N_13105,N_9506,N_11627);
nand U13106 (N_13106,N_10095,N_11416);
or U13107 (N_13107,N_10708,N_10500);
nand U13108 (N_13108,N_12163,N_10492);
and U13109 (N_13109,N_10221,N_10797);
or U13110 (N_13110,N_11815,N_12428);
nor U13111 (N_13111,N_10440,N_11717);
nor U13112 (N_13112,N_9781,N_10153);
or U13113 (N_13113,N_10870,N_12205);
nand U13114 (N_13114,N_10799,N_12079);
and U13115 (N_13115,N_9805,N_10871);
and U13116 (N_13116,N_12291,N_10082);
nor U13117 (N_13117,N_12051,N_9739);
nand U13118 (N_13118,N_10750,N_11364);
nor U13119 (N_13119,N_11865,N_10667);
xnor U13120 (N_13120,N_11979,N_11198);
or U13121 (N_13121,N_11437,N_11233);
and U13122 (N_13122,N_11525,N_11657);
or U13123 (N_13123,N_12342,N_10665);
xor U13124 (N_13124,N_11664,N_11193);
and U13125 (N_13125,N_11460,N_10038);
xnor U13126 (N_13126,N_10332,N_11013);
or U13127 (N_13127,N_9685,N_11943);
and U13128 (N_13128,N_9541,N_12324);
nor U13129 (N_13129,N_11304,N_11778);
and U13130 (N_13130,N_12049,N_12084);
nor U13131 (N_13131,N_9677,N_11503);
and U13132 (N_13132,N_10636,N_11354);
or U13133 (N_13133,N_10414,N_10639);
nor U13134 (N_13134,N_9855,N_10411);
nor U13135 (N_13135,N_10177,N_10364);
xor U13136 (N_13136,N_9891,N_9961);
or U13137 (N_13137,N_10554,N_11471);
nand U13138 (N_13138,N_11882,N_10071);
and U13139 (N_13139,N_11356,N_11276);
nand U13140 (N_13140,N_11401,N_9405);
and U13141 (N_13141,N_11323,N_10913);
nor U13142 (N_13142,N_10731,N_12378);
or U13143 (N_13143,N_10854,N_11962);
and U13144 (N_13144,N_10556,N_10372);
nand U13145 (N_13145,N_11534,N_9605);
xor U13146 (N_13146,N_11969,N_11678);
nor U13147 (N_13147,N_10642,N_9845);
xnor U13148 (N_13148,N_11039,N_10146);
and U13149 (N_13149,N_10588,N_9938);
nor U13150 (N_13150,N_10368,N_11351);
xor U13151 (N_13151,N_10227,N_11466);
nor U13152 (N_13152,N_9558,N_10999);
nand U13153 (N_13153,N_11326,N_12359);
or U13154 (N_13154,N_9606,N_11881);
or U13155 (N_13155,N_11538,N_10718);
and U13156 (N_13156,N_11946,N_12043);
and U13157 (N_13157,N_11587,N_11896);
or U13158 (N_13158,N_12456,N_9670);
nand U13159 (N_13159,N_10012,N_10974);
and U13160 (N_13160,N_10766,N_11967);
nand U13161 (N_13161,N_11753,N_12185);
nor U13162 (N_13162,N_9940,N_12330);
nor U13163 (N_13163,N_9649,N_11346);
nand U13164 (N_13164,N_12338,N_12325);
nand U13165 (N_13165,N_9922,N_11142);
or U13166 (N_13166,N_10137,N_9429);
or U13167 (N_13167,N_10085,N_11703);
xnor U13168 (N_13168,N_12306,N_10028);
nand U13169 (N_13169,N_10882,N_11000);
or U13170 (N_13170,N_10609,N_10517);
or U13171 (N_13171,N_11684,N_9829);
xor U13172 (N_13172,N_10253,N_9934);
xnor U13173 (N_13173,N_10404,N_10015);
nor U13174 (N_13174,N_10408,N_10939);
nor U13175 (N_13175,N_10135,N_12140);
and U13176 (N_13176,N_9733,N_10390);
nor U13177 (N_13177,N_12367,N_12475);
nand U13178 (N_13178,N_10482,N_10957);
and U13179 (N_13179,N_9441,N_10964);
nand U13180 (N_13180,N_10114,N_11371);
nor U13181 (N_13181,N_10059,N_10655);
nor U13182 (N_13182,N_10388,N_10864);
nand U13183 (N_13183,N_10455,N_10594);
and U13184 (N_13184,N_9619,N_11423);
or U13185 (N_13185,N_12105,N_11775);
nand U13186 (N_13186,N_10863,N_10503);
nor U13187 (N_13187,N_9514,N_10680);
or U13188 (N_13188,N_10420,N_11951);
nor U13189 (N_13189,N_10679,N_11199);
or U13190 (N_13190,N_11384,N_10890);
nor U13191 (N_13191,N_11938,N_10826);
nand U13192 (N_13192,N_10524,N_10362);
nor U13193 (N_13193,N_10070,N_11672);
xor U13194 (N_13194,N_11180,N_10722);
xnor U13195 (N_13195,N_12236,N_9381);
and U13196 (N_13196,N_11706,N_10249);
and U13197 (N_13197,N_9609,N_11475);
nand U13198 (N_13198,N_12145,N_11089);
nand U13199 (N_13199,N_11262,N_11574);
nand U13200 (N_13200,N_9577,N_12144);
and U13201 (N_13201,N_12488,N_10551);
nor U13202 (N_13202,N_11569,N_11425);
and U13203 (N_13203,N_11977,N_12451);
nor U13204 (N_13204,N_12006,N_10295);
or U13205 (N_13205,N_11135,N_11959);
and U13206 (N_13206,N_11592,N_11576);
nand U13207 (N_13207,N_9672,N_9859);
or U13208 (N_13208,N_11883,N_11691);
nand U13209 (N_13209,N_10961,N_11681);
xor U13210 (N_13210,N_10696,N_12468);
nand U13211 (N_13211,N_10635,N_9999);
nor U13212 (N_13212,N_9581,N_11675);
nor U13213 (N_13213,N_9666,N_11825);
and U13214 (N_13214,N_9866,N_12353);
xnor U13215 (N_13215,N_9613,N_10067);
nand U13216 (N_13216,N_9449,N_11480);
and U13217 (N_13217,N_11463,N_9478);
nor U13218 (N_13218,N_12355,N_9495);
nand U13219 (N_13219,N_9410,N_11395);
nor U13220 (N_13220,N_11944,N_11628);
nand U13221 (N_13221,N_11037,N_9750);
xnor U13222 (N_13222,N_11222,N_9944);
and U13223 (N_13223,N_9721,N_12393);
nand U13224 (N_13224,N_11130,N_9689);
and U13225 (N_13225,N_10538,N_11435);
nor U13226 (N_13226,N_10563,N_11770);
nand U13227 (N_13227,N_10115,N_11869);
nor U13228 (N_13228,N_11870,N_9903);
or U13229 (N_13229,N_9575,N_11289);
nor U13230 (N_13230,N_9848,N_9885);
nor U13231 (N_13231,N_11221,N_9642);
nor U13232 (N_13232,N_12175,N_11535);
xnor U13233 (N_13233,N_10749,N_10778);
nor U13234 (N_13234,N_9894,N_11688);
or U13235 (N_13235,N_9458,N_10055);
nand U13236 (N_13236,N_11234,N_11886);
or U13237 (N_13237,N_11484,N_10926);
and U13238 (N_13238,N_11982,N_11822);
xor U13239 (N_13239,N_12289,N_11521);
nand U13240 (N_13240,N_9500,N_10703);
xor U13241 (N_13241,N_11459,N_12023);
nand U13242 (N_13242,N_11740,N_11837);
nor U13243 (N_13243,N_10337,N_11030);
or U13244 (N_13244,N_11303,N_12296);
nor U13245 (N_13245,N_9626,N_12255);
and U13246 (N_13246,N_10001,N_9727);
and U13247 (N_13247,N_9488,N_10106);
and U13248 (N_13248,N_10248,N_9889);
nand U13249 (N_13249,N_9520,N_10687);
nand U13250 (N_13250,N_10353,N_11519);
nand U13251 (N_13251,N_9425,N_12405);
xor U13252 (N_13252,N_9991,N_9489);
or U13253 (N_13253,N_11390,N_10912);
nand U13254 (N_13254,N_10815,N_10512);
xor U13255 (N_13255,N_12490,N_9980);
or U13256 (N_13256,N_10771,N_9816);
nand U13257 (N_13257,N_9628,N_11536);
nand U13258 (N_13258,N_10526,N_11065);
or U13259 (N_13259,N_10618,N_12014);
nand U13260 (N_13260,N_10919,N_10881);
nand U13261 (N_13261,N_11266,N_10617);
nor U13262 (N_13262,N_10151,N_12005);
or U13263 (N_13263,N_10309,N_11729);
or U13264 (N_13264,N_11621,N_10536);
nand U13265 (N_13265,N_10462,N_9679);
or U13266 (N_13266,N_10384,N_10872);
or U13267 (N_13267,N_10054,N_11201);
and U13268 (N_13268,N_10619,N_12050);
nor U13269 (N_13269,N_10460,N_9973);
xor U13270 (N_13270,N_12458,N_11960);
nand U13271 (N_13271,N_11280,N_11024);
or U13272 (N_13272,N_10497,N_11673);
xor U13273 (N_13273,N_12258,N_10022);
nand U13274 (N_13274,N_9401,N_12369);
or U13275 (N_13275,N_11170,N_9498);
nor U13276 (N_13276,N_11154,N_10573);
and U13277 (N_13277,N_11698,N_11841);
nor U13278 (N_13278,N_10751,N_12044);
and U13279 (N_13279,N_11976,N_11265);
and U13280 (N_13280,N_9708,N_11084);
or U13281 (N_13281,N_9731,N_12002);
nor U13282 (N_13282,N_11512,N_12478);
nor U13283 (N_13283,N_11374,N_11007);
nor U13284 (N_13284,N_12448,N_10672);
or U13285 (N_13285,N_9782,N_12469);
or U13286 (N_13286,N_10458,N_11420);
and U13287 (N_13287,N_12075,N_9843);
xor U13288 (N_13288,N_10321,N_12047);
nor U13289 (N_13289,N_10706,N_11830);
and U13290 (N_13290,N_12283,N_10675);
xnor U13291 (N_13291,N_10330,N_11397);
nor U13292 (N_13292,N_10620,N_10830);
xor U13293 (N_13293,N_10793,N_10650);
or U13294 (N_13294,N_10000,N_9795);
nand U13295 (N_13295,N_10928,N_11787);
or U13296 (N_13296,N_10710,N_9955);
nand U13297 (N_13297,N_11388,N_9943);
and U13298 (N_13298,N_12380,N_12012);
nor U13299 (N_13299,N_9692,N_11929);
and U13300 (N_13300,N_11217,N_9656);
nand U13301 (N_13301,N_9758,N_11448);
xnor U13302 (N_13302,N_10405,N_10684);
and U13303 (N_13303,N_9967,N_10803);
or U13304 (N_13304,N_10254,N_11575);
or U13305 (N_13305,N_10247,N_9474);
nand U13306 (N_13306,N_11149,N_12375);
and U13307 (N_13307,N_10924,N_10689);
nand U13308 (N_13308,N_10308,N_12491);
xnor U13309 (N_13309,N_9574,N_9908);
nor U13310 (N_13310,N_9459,N_9684);
and U13311 (N_13311,N_12285,N_10150);
nor U13312 (N_13312,N_11690,N_10942);
and U13313 (N_13313,N_10673,N_10188);
and U13314 (N_13314,N_9376,N_9924);
nand U13315 (N_13315,N_10180,N_12021);
nand U13316 (N_13316,N_10856,N_12346);
xor U13317 (N_13317,N_10434,N_11795);
and U13318 (N_13318,N_12293,N_10845);
or U13319 (N_13319,N_12169,N_9964);
and U13320 (N_13320,N_9835,N_11968);
nor U13321 (N_13321,N_10587,N_12366);
and U13322 (N_13322,N_9518,N_10561);
and U13323 (N_13323,N_10657,N_11023);
nand U13324 (N_13324,N_9513,N_10940);
nor U13325 (N_13325,N_11338,N_10829);
and U13326 (N_13326,N_9746,N_10662);
nor U13327 (N_13327,N_10732,N_10035);
or U13328 (N_13328,N_10021,N_11263);
or U13329 (N_13329,N_11885,N_9919);
or U13330 (N_13330,N_11283,N_10052);
xor U13331 (N_13331,N_10413,N_9772);
and U13332 (N_13332,N_11813,N_9652);
nor U13333 (N_13333,N_11470,N_11782);
nand U13334 (N_13334,N_10422,N_10659);
and U13335 (N_13335,N_12422,N_11925);
and U13336 (N_13336,N_11190,N_10467);
and U13337 (N_13337,N_10261,N_9935);
and U13338 (N_13338,N_11322,N_11482);
or U13339 (N_13339,N_11555,N_11963);
nor U13340 (N_13340,N_11017,N_10511);
and U13341 (N_13341,N_12116,N_10827);
nor U13342 (N_13342,N_12256,N_10400);
xnor U13343 (N_13343,N_11169,N_10931);
or U13344 (N_13344,N_10980,N_10712);
nor U13345 (N_13345,N_12083,N_12404);
nor U13346 (N_13346,N_11196,N_10108);
nand U13347 (N_13347,N_9392,N_9998);
nor U13348 (N_13348,N_10973,N_11097);
and U13349 (N_13349,N_11908,N_11159);
or U13350 (N_13350,N_10287,N_12159);
xor U13351 (N_13351,N_12336,N_11783);
and U13352 (N_13352,N_11629,N_10347);
or U13353 (N_13353,N_11305,N_10092);
and U13354 (N_13354,N_11625,N_12495);
nand U13355 (N_13355,N_10029,N_11953);
nand U13356 (N_13356,N_9926,N_12103);
nand U13357 (N_13357,N_10317,N_9664);
nand U13358 (N_13358,N_10050,N_10457);
nor U13359 (N_13359,N_12031,N_11763);
nor U13360 (N_13360,N_9643,N_11439);
or U13361 (N_13361,N_10410,N_9693);
or U13362 (N_13362,N_12467,N_10258);
xnor U13363 (N_13363,N_12197,N_12160);
xnor U13364 (N_13364,N_9960,N_10505);
nor U13365 (N_13365,N_11197,N_10402);
xnor U13366 (N_13366,N_10542,N_12493);
nor U13367 (N_13367,N_9909,N_12459);
nand U13368 (N_13368,N_9734,N_9815);
nand U13369 (N_13369,N_11367,N_11637);
nand U13370 (N_13370,N_10637,N_10688);
nor U13371 (N_13371,N_12390,N_10215);
or U13372 (N_13372,N_11585,N_9545);
or U13373 (N_13373,N_10477,N_10652);
nand U13374 (N_13374,N_11579,N_12373);
or U13375 (N_13375,N_12216,N_10131);
nor U13376 (N_13376,N_9595,N_9916);
nor U13377 (N_13377,N_10379,N_11656);
nor U13378 (N_13378,N_9607,N_12251);
nand U13379 (N_13379,N_10669,N_11031);
xor U13380 (N_13380,N_12399,N_9987);
xnor U13381 (N_13381,N_10398,N_11213);
nand U13382 (N_13382,N_11219,N_11091);
or U13383 (N_13383,N_10087,N_11297);
or U13384 (N_13384,N_12470,N_12215);
nand U13385 (N_13385,N_10763,N_10086);
nor U13386 (N_13386,N_11108,N_10061);
or U13387 (N_13387,N_11565,N_11204);
nand U13388 (N_13388,N_11252,N_10743);
and U13389 (N_13389,N_12360,N_12003);
nand U13390 (N_13390,N_10993,N_10167);
or U13391 (N_13391,N_10274,N_10521);
or U13392 (N_13392,N_9450,N_9557);
nor U13393 (N_13393,N_10547,N_10387);
xor U13394 (N_13394,N_10794,N_11335);
nand U13395 (N_13395,N_10228,N_11701);
and U13396 (N_13396,N_11344,N_12171);
and U13397 (N_13397,N_10155,N_10892);
xnor U13398 (N_13398,N_9387,N_12463);
nor U13399 (N_13399,N_10299,N_11008);
xnor U13400 (N_13400,N_12037,N_9825);
nor U13401 (N_13401,N_10046,N_10549);
nor U13402 (N_13402,N_9735,N_9913);
nand U13403 (N_13403,N_9977,N_10956);
nor U13404 (N_13404,N_10343,N_10615);
or U13405 (N_13405,N_12112,N_11614);
xor U13406 (N_13406,N_11034,N_10081);
or U13407 (N_13407,N_11659,N_10777);
nand U13408 (N_13408,N_10780,N_9872);
nand U13409 (N_13409,N_11889,N_12425);
nor U13410 (N_13410,N_11987,N_10428);
or U13411 (N_13411,N_11754,N_9427);
and U13412 (N_13412,N_11454,N_9723);
and U13413 (N_13413,N_11990,N_11533);
nor U13414 (N_13414,N_10158,N_10435);
nor U13415 (N_13415,N_12362,N_10595);
nand U13416 (N_13416,N_10677,N_10752);
nor U13417 (N_13417,N_11250,N_11357);
or U13418 (N_13418,N_12317,N_12011);
nand U13419 (N_13419,N_11478,N_11741);
and U13420 (N_13420,N_9497,N_10715);
and U13421 (N_13421,N_10945,N_10156);
and U13422 (N_13422,N_10183,N_11796);
or U13423 (N_13423,N_9426,N_12115);
nor U13424 (N_13424,N_10178,N_12403);
and U13425 (N_13425,N_10915,N_9818);
nor U13426 (N_13426,N_10911,N_10342);
nand U13427 (N_13427,N_9748,N_11756);
nor U13428 (N_13428,N_11748,N_12060);
or U13429 (N_13429,N_9752,N_9665);
nor U13430 (N_13430,N_12297,N_11984);
xnor U13431 (N_13431,N_10213,N_12277);
and U13432 (N_13432,N_11306,N_11288);
nor U13433 (N_13433,N_12063,N_10427);
xor U13434 (N_13434,N_10433,N_10770);
xnor U13435 (N_13435,N_9446,N_10880);
xnor U13436 (N_13436,N_10714,N_11733);
nand U13437 (N_13437,N_11623,N_11732);
nor U13438 (N_13438,N_12129,N_9436);
nand U13439 (N_13439,N_11709,N_9678);
and U13440 (N_13440,N_10624,N_12429);
or U13441 (N_13441,N_10735,N_11080);
or U13442 (N_13442,N_12104,N_11735);
or U13443 (N_13443,N_9737,N_10496);
or U13444 (N_13444,N_10842,N_10048);
nor U13445 (N_13445,N_11695,N_12066);
nand U13446 (N_13446,N_11864,N_12048);
nand U13447 (N_13447,N_9802,N_11552);
xor U13448 (N_13448,N_9501,N_11531);
nor U13449 (N_13449,N_11015,N_11989);
nor U13450 (N_13450,N_11731,N_10903);
nand U13451 (N_13451,N_10352,N_11986);
or U13452 (N_13452,N_12089,N_9883);
or U13453 (N_13453,N_9753,N_12143);
or U13454 (N_13454,N_11966,N_10692);
nor U13455 (N_13455,N_11751,N_11281);
or U13456 (N_13456,N_9836,N_11077);
xnor U13457 (N_13457,N_11879,N_11157);
nor U13458 (N_13458,N_11006,N_11711);
nor U13459 (N_13459,N_10698,N_10101);
nor U13460 (N_13460,N_12088,N_11229);
and U13461 (N_13461,N_11674,N_12382);
or U13462 (N_13462,N_12158,N_9864);
xor U13463 (N_13463,N_12170,N_10792);
nor U13464 (N_13464,N_10091,N_10267);
nor U13465 (N_13465,N_9567,N_12266);
nand U13466 (N_13466,N_10544,N_11597);
and U13467 (N_13467,N_12135,N_10276);
or U13468 (N_13468,N_12244,N_11790);
and U13469 (N_13469,N_10504,N_9796);
or U13470 (N_13470,N_11269,N_10540);
or U13471 (N_13471,N_10991,N_10307);
and U13472 (N_13472,N_10192,N_10954);
and U13473 (N_13473,N_11465,N_11156);
nand U13474 (N_13474,N_10162,N_10789);
nand U13475 (N_13475,N_10345,N_10860);
nor U13476 (N_13476,N_12473,N_11063);
nand U13477 (N_13477,N_11045,N_11961);
nand U13478 (N_13478,N_9965,N_9945);
nand U13479 (N_13479,N_11476,N_11923);
and U13480 (N_13480,N_11044,N_11993);
or U13481 (N_13481,N_12207,N_9555);
or U13482 (N_13482,N_10487,N_10013);
nand U13483 (N_13483,N_10303,N_12178);
or U13484 (N_13484,N_10755,N_12033);
nand U13485 (N_13485,N_12441,N_11858);
nor U13486 (N_13486,N_11939,N_10088);
nor U13487 (N_13487,N_10139,N_11956);
nor U13488 (N_13488,N_11598,N_11373);
or U13489 (N_13489,N_11461,N_12479);
nor U13490 (N_13490,N_11557,N_10867);
xor U13491 (N_13491,N_9419,N_11722);
or U13492 (N_13492,N_10202,N_10049);
or U13493 (N_13493,N_11317,N_10597);
nor U13494 (N_13494,N_9578,N_10824);
nor U13495 (N_13495,N_12295,N_9424);
or U13496 (N_13496,N_9969,N_11457);
nand U13497 (N_13497,N_11331,N_11880);
or U13498 (N_13498,N_12161,N_10760);
xnor U13499 (N_13499,N_11358,N_12343);
nand U13500 (N_13500,N_12449,N_11411);
nor U13501 (N_13501,N_11658,N_10141);
and U13502 (N_13502,N_10959,N_10717);
nor U13503 (N_13503,N_9496,N_10895);
nand U13504 (N_13504,N_9635,N_11035);
nor U13505 (N_13505,N_10564,N_11708);
nor U13506 (N_13506,N_9399,N_11455);
nand U13507 (N_13507,N_12138,N_11850);
and U13508 (N_13508,N_10334,N_10693);
or U13509 (N_13509,N_10932,N_10644);
nor U13510 (N_13510,N_11440,N_10369);
and U13511 (N_13511,N_11589,N_12334);
nand U13512 (N_13512,N_10257,N_10062);
nand U13513 (N_13513,N_10886,N_9992);
nor U13514 (N_13514,N_12328,N_11823);
or U13515 (N_13515,N_10426,N_11724);
nand U13516 (N_13516,N_11873,N_9933);
or U13517 (N_13517,N_11081,N_9880);
and U13518 (N_13518,N_10058,N_12377);
xor U13519 (N_13519,N_10523,N_10357);
or U13520 (N_13520,N_10475,N_10819);
nand U13521 (N_13521,N_10011,N_9983);
nor U13522 (N_13522,N_12444,N_11172);
nand U13523 (N_13523,N_10600,N_12381);
nor U13524 (N_13524,N_9421,N_11522);
and U13525 (N_13525,N_10394,N_9807);
and U13526 (N_13526,N_12368,N_10093);
and U13527 (N_13527,N_10699,N_9775);
and U13528 (N_13528,N_10808,N_9993);
nand U13529 (N_13529,N_9493,N_10873);
nand U13530 (N_13530,N_11713,N_10320);
or U13531 (N_13531,N_10323,N_9766);
nand U13532 (N_13532,N_10855,N_11113);
xor U13533 (N_13533,N_11333,N_10148);
nor U13534 (N_13534,N_10975,N_12165);
and U13535 (N_13535,N_12080,N_11155);
and U13536 (N_13536,N_9923,N_10370);
or U13537 (N_13537,N_10579,N_10900);
or U13538 (N_13538,N_12410,N_11123);
nor U13539 (N_13539,N_10128,N_10593);
nand U13540 (N_13540,N_11852,N_11027);
nor U13541 (N_13541,N_11887,N_10161);
nor U13542 (N_13542,N_12218,N_11298);
xnor U13543 (N_13543,N_9970,N_10377);
nor U13544 (N_13544,N_9756,N_10585);
and U13545 (N_13545,N_11019,N_10582);
nor U13546 (N_13546,N_10513,N_9408);
or U13547 (N_13547,N_11884,N_12437);
or U13548 (N_13548,N_10762,N_10281);
nor U13549 (N_13549,N_11228,N_10914);
nor U13550 (N_13550,N_9762,N_11893);
xnor U13551 (N_13551,N_9475,N_9745);
and U13552 (N_13552,N_11025,N_11430);
and U13553 (N_13553,N_9597,N_10884);
nand U13554 (N_13554,N_9996,N_11542);
xor U13555 (N_13555,N_11115,N_11818);
and U13556 (N_13556,N_11784,N_10160);
and U13557 (N_13557,N_10283,N_9792);
nor U13558 (N_13558,N_9412,N_9634);
nand U13559 (N_13559,N_11513,N_11667);
nand U13560 (N_13560,N_10906,N_10844);
nand U13561 (N_13561,N_10927,N_12154);
and U13562 (N_13562,N_11200,N_11211);
nor U13563 (N_13563,N_9927,N_9504);
xnor U13564 (N_13564,N_9981,N_11771);
nor U13565 (N_13565,N_10360,N_12423);
or U13566 (N_13566,N_12180,N_12001);
or U13567 (N_13567,N_10235,N_10349);
and U13568 (N_13568,N_10103,N_9588);
or U13569 (N_13569,N_10126,N_11253);
nor U13570 (N_13570,N_10083,N_10685);
or U13571 (N_13571,N_9915,N_11978);
nand U13572 (N_13572,N_11140,N_11072);
xor U13573 (N_13573,N_11369,N_10992);
or U13574 (N_13574,N_9442,N_11964);
xor U13575 (N_13575,N_11223,N_9617);
or U13576 (N_13576,N_10031,N_11143);
or U13577 (N_13577,N_9724,N_12134);
xor U13578 (N_13578,N_11381,N_10548);
nand U13579 (N_13579,N_11502,N_12118);
nor U13580 (N_13580,N_12292,N_10105);
or U13581 (N_13581,N_10239,N_9929);
xnor U13582 (N_13582,N_11654,N_11988);
nand U13583 (N_13583,N_11805,N_9486);
xnor U13584 (N_13584,N_10130,N_9849);
nand U13585 (N_13585,N_10702,N_11996);
and U13586 (N_13586,N_9461,N_11867);
nand U13587 (N_13587,N_9669,N_11398);
xor U13588 (N_13588,N_12186,N_10004);
nor U13589 (N_13589,N_9725,N_12406);
xor U13590 (N_13590,N_10136,N_10584);
nor U13591 (N_13591,N_10331,N_12361);
xor U13592 (N_13592,N_10232,N_10798);
or U13593 (N_13593,N_10625,N_10005);
xnor U13594 (N_13594,N_9700,N_10217);
nand U13595 (N_13595,N_9890,N_9741);
nand U13596 (N_13596,N_10252,N_12172);
and U13597 (N_13597,N_10211,N_11504);
or U13598 (N_13598,N_12391,N_11545);
xnor U13599 (N_13599,N_11747,N_10908);
and U13600 (N_13600,N_10545,N_11258);
and U13601 (N_13601,N_10159,N_10386);
and U13602 (N_13602,N_11626,N_11714);
and U13603 (N_13603,N_12201,N_11189);
nand U13604 (N_13604,N_9823,N_10738);
nand U13605 (N_13605,N_10831,N_11919);
nor U13606 (N_13606,N_10200,N_10023);
or U13607 (N_13607,N_11524,N_11387);
and U13608 (N_13608,N_9637,N_11591);
nor U13609 (N_13609,N_11347,N_12280);
nand U13610 (N_13610,N_9414,N_9989);
nand U13611 (N_13611,N_12408,N_12045);
nand U13612 (N_13612,N_11224,N_11386);
or U13613 (N_13613,N_10224,N_9481);
nand U13614 (N_13614,N_12102,N_12004);
xnor U13615 (N_13615,N_9460,N_11660);
xnor U13616 (N_13616,N_11828,N_10575);
and U13617 (N_13617,N_10800,N_11085);
or U13618 (N_13618,N_10424,N_10833);
and U13619 (N_13619,N_9517,N_10754);
xor U13620 (N_13620,N_11906,N_10191);
xor U13621 (N_13621,N_12231,N_12237);
or U13622 (N_13622,N_10952,N_12435);
xnor U13623 (N_13623,N_12100,N_10837);
and U13624 (N_13624,N_9385,N_10304);
and U13625 (N_13625,N_9472,N_11241);
and U13626 (N_13626,N_12028,N_9827);
and U13627 (N_13627,N_11849,N_11379);
nand U13628 (N_13628,N_10361,N_9375);
nor U13629 (N_13629,N_9813,N_11900);
or U13630 (N_13630,N_10602,N_10293);
xnor U13631 (N_13631,N_10431,N_12128);
or U13632 (N_13632,N_11500,N_10723);
xor U13633 (N_13633,N_9939,N_10943);
nor U13634 (N_13634,N_11001,N_11309);
nand U13635 (N_13635,N_11635,N_9715);
nand U13636 (N_13636,N_10574,N_11530);
nor U13637 (N_13637,N_10056,N_11528);
nand U13638 (N_13638,N_12228,N_12126);
or U13639 (N_13639,N_12481,N_11419);
or U13640 (N_13640,N_11800,N_11148);
nor U13641 (N_13641,N_11937,N_11636);
nor U13642 (N_13642,N_10262,N_11651);
or U13643 (N_13643,N_11111,N_11100);
xnor U13644 (N_13644,N_10316,N_12062);
nor U13645 (N_13645,N_9415,N_12322);
nand U13646 (N_13646,N_9953,N_11901);
nand U13647 (N_13647,N_10690,N_10704);
and U13648 (N_13648,N_10149,N_10288);
xnor U13649 (N_13649,N_9473,N_10820);
and U13650 (N_13650,N_11328,N_10421);
and U13651 (N_13651,N_9491,N_11167);
or U13652 (N_13652,N_11902,N_10312);
xor U13653 (N_13653,N_10182,N_9476);
or U13654 (N_13654,N_12300,N_9718);
or U13655 (N_13655,N_10483,N_11746);
nor U13656 (N_13656,N_10187,N_10645);
or U13657 (N_13657,N_9515,N_12101);
nor U13658 (N_13658,N_10107,N_10066);
or U13659 (N_13659,N_10832,N_9906);
nor U13660 (N_13660,N_9612,N_12376);
and U13661 (N_13661,N_11353,N_9641);
or U13662 (N_13662,N_10218,N_10367);
nor U13663 (N_13663,N_11445,N_12019);
nor U13664 (N_13664,N_12316,N_10243);
and U13665 (N_13665,N_11467,N_9730);
and U13666 (N_13666,N_9422,N_9580);
nor U13667 (N_13667,N_9875,N_11921);
or U13668 (N_13668,N_11812,N_11965);
nor U13669 (N_13669,N_9384,N_11237);
nor U13670 (N_13670,N_11078,N_10076);
nor U13671 (N_13671,N_10498,N_10897);
or U13672 (N_13672,N_11610,N_11527);
nand U13673 (N_13673,N_10506,N_11549);
nand U13674 (N_13674,N_11514,N_10701);
and U13675 (N_13675,N_11264,N_10089);
or U13676 (N_13676,N_11750,N_11261);
or U13677 (N_13677,N_11086,N_12417);
or U13678 (N_13678,N_10796,N_9554);
nor U13679 (N_13679,N_11611,N_10336);
and U13680 (N_13680,N_11138,N_11874);
nand U13681 (N_13681,N_10591,N_11742);
nand U13682 (N_13682,N_12082,N_10865);
and U13683 (N_13683,N_9388,N_12174);
or U13684 (N_13684,N_11161,N_11018);
or U13685 (N_13685,N_10383,N_10519);
or U13686 (N_13686,N_10488,N_9548);
xor U13687 (N_13687,N_11558,N_9614);
nor U13688 (N_13688,N_10570,N_10626);
nor U13689 (N_13689,N_9448,N_10060);
nor U13690 (N_13690,N_10768,N_11311);
xnor U13691 (N_13691,N_10163,N_9951);
xnor U13692 (N_13692,N_9591,N_11777);
nand U13693 (N_13693,N_9869,N_11011);
and U13694 (N_13694,N_11666,N_12480);
nand U13695 (N_13695,N_10466,N_9773);
and U13696 (N_13696,N_11909,N_11096);
nor U13697 (N_13697,N_9701,N_11972);
or U13698 (N_13698,N_11071,N_11998);
nand U13699 (N_13699,N_9445,N_9854);
nand U13700 (N_13700,N_12213,N_10887);
and U13701 (N_13701,N_9553,N_9754);
and U13702 (N_13702,N_10607,N_11109);
nand U13703 (N_13703,N_9840,N_12262);
nor U13704 (N_13704,N_11101,N_10568);
nor U13705 (N_13705,N_12460,N_11163);
xor U13706 (N_13706,N_11662,N_11436);
nor U13707 (N_13707,N_11057,N_10120);
nand U13708 (N_13708,N_9896,N_9867);
xnor U13709 (N_13709,N_11930,N_12156);
or U13710 (N_13710,N_9525,N_10017);
and U13711 (N_13711,N_10623,N_9680);
nand U13712 (N_13712,N_10432,N_10256);
xnor U13713 (N_13713,N_12190,N_12153);
nand U13714 (N_13714,N_10338,N_10425);
nand U13715 (N_13715,N_9958,N_11363);
nor U13716 (N_13716,N_10767,N_9403);
and U13717 (N_13717,N_10325,N_9633);
and U13718 (N_13718,N_9851,N_10231);
nand U13719 (N_13719,N_10846,N_11831);
or U13720 (N_13720,N_11808,N_10787);
nor U13721 (N_13721,N_11641,N_12247);
nand U13722 (N_13722,N_11898,N_10282);
nand U13723 (N_13723,N_12344,N_9409);
xnor U13724 (N_13724,N_10788,N_9767);
nor U13725 (N_13725,N_12131,N_11319);
and U13726 (N_13726,N_10592,N_10329);
or U13727 (N_13727,N_11215,N_10769);
nor U13728 (N_13728,N_11897,N_10173);
nand U13729 (N_13729,N_11863,N_10399);
nand U13730 (N_13730,N_12257,N_11760);
nor U13731 (N_13731,N_12409,N_12097);
and U13732 (N_13732,N_12015,N_10392);
and U13733 (N_13733,N_9631,N_9543);
nor U13734 (N_13734,N_11947,N_10416);
and U13735 (N_13735,N_10933,N_10147);
nand U13736 (N_13736,N_10891,N_12496);
nand U13737 (N_13737,N_9832,N_9897);
nand U13738 (N_13738,N_10047,N_11021);
and U13739 (N_13739,N_9440,N_12267);
and U13740 (N_13740,N_12339,N_12326);
and U13741 (N_13741,N_11762,N_11050);
or U13742 (N_13742,N_10807,N_9761);
nor U13743 (N_13743,N_12471,N_11194);
and U13744 (N_13744,N_10776,N_12394);
nand U13745 (N_13745,N_11911,N_10951);
or U13746 (N_13746,N_10539,N_12402);
nor U13747 (N_13747,N_12032,N_12301);
nor U13748 (N_13748,N_11994,N_9533);
or U13749 (N_13749,N_12433,N_10344);
nor U13750 (N_13750,N_10341,N_11604);
and U13751 (N_13751,N_9794,N_10507);
xnor U13752 (N_13752,N_11337,N_11509);
or U13753 (N_13753,N_11058,N_12419);
nand U13754 (N_13754,N_12421,N_12166);
xor U13755 (N_13755,N_9611,N_10967);
and U13756 (N_13756,N_11663,N_10237);
nor U13757 (N_13757,N_11107,N_10670);
nor U13758 (N_13758,N_11259,N_11580);
nor U13759 (N_13759,N_9418,N_11608);
nand U13760 (N_13760,N_9604,N_12024);
nor U13761 (N_13761,N_10516,N_11426);
xor U13762 (N_13762,N_12388,N_11888);
or U13763 (N_13763,N_9393,N_10241);
xor U13764 (N_13764,N_11749,N_10983);
and U13765 (N_13765,N_12030,N_12146);
nor U13766 (N_13766,N_9824,N_9632);
nand U13767 (N_13767,N_9623,N_11737);
nor U13768 (N_13768,N_11903,N_12436);
or U13769 (N_13769,N_11421,N_11779);
nor U13770 (N_13770,N_11920,N_11780);
or U13771 (N_13771,N_10429,N_11498);
xor U13772 (N_13772,N_11110,N_11846);
or U13773 (N_13773,N_11473,N_10734);
nor U13774 (N_13774,N_12187,N_11612);
and U13775 (N_13775,N_10565,N_12287);
nor U13776 (N_13776,N_11776,N_11497);
and U13777 (N_13777,N_10350,N_10436);
nand U13778 (N_13778,N_9572,N_9663);
nand U13779 (N_13779,N_12358,N_11079);
nor U13780 (N_13780,N_11974,N_10459);
and U13781 (N_13781,N_12182,N_12275);
nand U13782 (N_13782,N_12477,N_12284);
and U13783 (N_13783,N_10138,N_11590);
nand U13784 (N_13784,N_9510,N_10622);
nor U13785 (N_13785,N_10883,N_11472);
nor U13786 (N_13786,N_11046,N_10616);
or U13787 (N_13787,N_9540,N_12168);
and U13788 (N_13788,N_10656,N_10326);
nor U13789 (N_13789,N_10366,N_10447);
xnor U13790 (N_13790,N_9583,N_9601);
nand U13791 (N_13791,N_9433,N_11112);
nand U13792 (N_13792,N_9596,N_11630);
and U13793 (N_13793,N_11772,N_12087);
or U13794 (N_13794,N_9988,N_11523);
and U13795 (N_13795,N_10359,N_11617);
and U13796 (N_13796,N_9690,N_10557);
xnor U13797 (N_13797,N_12370,N_10346);
xor U13798 (N_13798,N_9675,N_9529);
nand U13799 (N_13799,N_9884,N_11313);
nor U13800 (N_13800,N_9389,N_11505);
or U13801 (N_13801,N_9404,N_12055);
or U13802 (N_13802,N_11434,N_12099);
nand U13803 (N_13803,N_9625,N_10209);
or U13804 (N_13804,N_10003,N_9707);
nand U13805 (N_13805,N_10613,N_11872);
nand U13806 (N_13806,N_12440,N_11727);
or U13807 (N_13807,N_11451,N_11493);
or U13808 (N_13808,N_9785,N_10979);
and U13809 (N_13809,N_11005,N_11256);
and U13810 (N_13810,N_9978,N_11408);
and U13811 (N_13811,N_11235,N_11362);
and U13812 (N_13812,N_11560,N_11757);
nand U13813 (N_13813,N_11769,N_11299);
nand U13814 (N_13814,N_11042,N_11230);
nand U13815 (N_13815,N_9858,N_10121);
nor U13816 (N_13816,N_10464,N_12418);
or U13817 (N_13817,N_10818,N_12120);
or U13818 (N_13818,N_12069,N_10222);
nor U13819 (N_13819,N_10078,N_11618);
nand U13820 (N_13820,N_11209,N_10893);
nand U13821 (N_13821,N_9465,N_11441);
nand U13822 (N_13822,N_10920,N_11047);
or U13823 (N_13823,N_9566,N_12462);
nand U13824 (N_13824,N_10772,N_11834);
and U13825 (N_13825,N_9787,N_9561);
and U13826 (N_13826,N_11802,N_11345);
and U13827 (N_13827,N_10558,N_11429);
nand U13828 (N_13828,N_10839,N_11056);
nand U13829 (N_13829,N_10397,N_9398);
nor U13830 (N_13830,N_11682,N_11043);
or U13831 (N_13831,N_11268,N_10726);
nand U13832 (N_13832,N_9477,N_10461);
or U13833 (N_13833,N_10109,N_11833);
nor U13834 (N_13834,N_9526,N_11212);
and U13835 (N_13835,N_11644,N_11060);
and U13836 (N_13836,N_11766,N_10097);
nor U13837 (N_13837,N_9638,N_9911);
nand U13838 (N_13838,N_9952,N_10950);
or U13839 (N_13839,N_11378,N_10296);
nand U13840 (N_13840,N_9485,N_10270);
nor U13841 (N_13841,N_9716,N_9764);
and U13842 (N_13842,N_10185,N_11076);
nand U13843 (N_13843,N_12482,N_12016);
nor U13844 (N_13844,N_10102,N_11781);
and U13845 (N_13845,N_12085,N_10894);
xor U13846 (N_13846,N_11366,N_10423);
nor U13847 (N_13847,N_9985,N_11529);
or U13848 (N_13848,N_9556,N_11877);
nor U13849 (N_13849,N_10234,N_11593);
nor U13850 (N_13850,N_9876,N_11671);
or U13851 (N_13851,N_11332,N_11646);
nor U13852 (N_13852,N_10724,N_9995);
or U13853 (N_13853,N_12432,N_11764);
nor U13854 (N_13854,N_9661,N_11294);
nand U13855 (N_13855,N_10569,N_11202);
or U13856 (N_13856,N_11186,N_12223);
nand U13857 (N_13857,N_9571,N_10175);
xnor U13858 (N_13858,N_10885,N_10899);
or U13859 (N_13859,N_11942,N_10879);
nor U13860 (N_13860,N_10375,N_10681);
or U13861 (N_13861,N_11913,N_9798);
or U13862 (N_13862,N_11272,N_11620);
nor U13863 (N_13863,N_10474,N_9768);
and U13864 (N_13864,N_10468,N_10470);
or U13865 (N_13865,N_11726,N_12072);
nand U13866 (N_13866,N_11860,N_11638);
nor U13867 (N_13867,N_11890,N_9817);
and U13868 (N_13868,N_10948,N_11275);
nor U13869 (N_13869,N_9569,N_9532);
nand U13870 (N_13870,N_9966,N_12188);
nor U13871 (N_13871,N_10255,N_12333);
nor U13872 (N_13872,N_11915,N_9760);
nor U13873 (N_13873,N_10683,N_10660);
nor U13874 (N_13874,N_9779,N_11349);
and U13875 (N_13875,N_10363,N_9600);
nand U13876 (N_13876,N_11296,N_11236);
xor U13877 (N_13877,N_10981,N_9717);
nor U13878 (N_13878,N_9651,N_11546);
or U13879 (N_13879,N_10633,N_10251);
or U13880 (N_13880,N_11827,N_11195);
nand U13881 (N_13881,N_9732,N_10562);
nor U13882 (N_13882,N_10938,N_12350);
xor U13883 (N_13883,N_9799,N_11508);
xor U13884 (N_13884,N_11866,N_9912);
xnor U13885 (N_13885,N_12179,N_10286);
nand U13886 (N_13886,N_12260,N_10530);
nand U13887 (N_13887,N_9400,N_10518);
nor U13888 (N_13888,N_11254,N_10122);
nand U13889 (N_13889,N_11668,N_9594);
and U13890 (N_13890,N_10495,N_12254);
xnor U13891 (N_13891,N_12204,N_9759);
nor U13892 (N_13892,N_10014,N_9963);
and U13893 (N_13893,N_9974,N_11761);
nor U13894 (N_13894,N_11099,N_12208);
or U13895 (N_13895,N_9711,N_9744);
or U13896 (N_13896,N_10853,N_12225);
nor U13897 (N_13897,N_12261,N_10774);
and U13898 (N_13898,N_12438,N_11279);
nor U13899 (N_13899,N_12466,N_11320);
and U13900 (N_13900,N_12310,N_10118);
nor U13901 (N_13901,N_11360,N_10073);
and U13902 (N_13902,N_11458,N_10116);
nand U13903 (N_13903,N_11607,N_11801);
and U13904 (N_13904,N_12414,N_11613);
and U13905 (N_13905,N_11372,N_9482);
nand U13906 (N_13906,N_11181,N_11012);
and U13907 (N_13907,N_11032,N_10550);
nor U13908 (N_13908,N_10963,N_10297);
and U13909 (N_13909,N_12331,N_12499);
nor U13910 (N_13910,N_10443,N_11758);
and U13911 (N_13911,N_12349,N_9534);
nand U13912 (N_13912,N_9490,N_10306);
nand U13913 (N_13913,N_9783,N_10889);
or U13914 (N_13914,N_11798,N_9769);
xor U13915 (N_13915,N_11314,N_12020);
nand U13916 (N_13916,N_10034,N_11376);
nor U13917 (N_13917,N_9530,N_10802);
nor U13918 (N_13918,N_10560,N_10328);
or U13919 (N_13919,N_12076,N_9920);
nor U13920 (N_13920,N_12227,N_10327);
or U13921 (N_13921,N_11819,N_10847);
nor U13922 (N_13922,N_9865,N_9946);
and U13923 (N_13923,N_11334,N_10838);
or U13924 (N_13924,N_10110,N_10782);
and U13925 (N_13925,N_10520,N_10527);
and U13926 (N_13926,N_10484,N_9905);
or U13927 (N_13927,N_10955,N_10207);
nand U13928 (N_13928,N_10621,N_11083);
nor U13929 (N_13929,N_12497,N_10172);
nand U13930 (N_13930,N_12457,N_11554);
and U13931 (N_13931,N_11799,N_11009);
xor U13932 (N_13932,N_10785,N_10965);
nor U13933 (N_13933,N_11061,N_9895);
and U13934 (N_13934,N_10960,N_11225);
nor U13935 (N_13935,N_11718,N_12219);
xor U13936 (N_13936,N_11293,N_9480);
nor U13937 (N_13937,N_9790,N_11064);
or U13938 (N_13938,N_10084,N_10759);
or U13939 (N_13939,N_9793,N_10204);
nor U13940 (N_13940,N_9874,N_11583);
xnor U13941 (N_13941,N_12290,N_9483);
and U13942 (N_13942,N_12249,N_12253);
xor U13943 (N_13943,N_12455,N_10566);
or U13944 (N_13944,N_10995,N_11290);
or U13945 (N_13945,N_9457,N_9503);
nor U13946 (N_13946,N_12442,N_11940);
xor U13947 (N_13947,N_10403,N_10812);
nor U13948 (N_13948,N_10096,N_11088);
or U13949 (N_13949,N_9847,N_10934);
nor U13950 (N_13950,N_11075,N_10273);
xnor U13951 (N_13951,N_9928,N_11786);
and U13952 (N_13952,N_10654,N_9592);
nand U13953 (N_13953,N_12476,N_11507);
xor U13954 (N_13954,N_11715,N_9487);
and U13955 (N_13955,N_9438,N_10748);
or U13956 (N_13956,N_10154,N_11710);
or U13957 (N_13957,N_11596,N_11543);
nand U13958 (N_13958,N_11797,N_10816);
nor U13959 (N_13959,N_11479,N_9646);
nand U13960 (N_13960,N_10836,N_11418);
or U13961 (N_13961,N_10858,N_10909);
and U13962 (N_13962,N_11409,N_12356);
nor U13963 (N_13963,N_10786,N_12157);
nand U13964 (N_13964,N_12221,N_11179);
and U13965 (N_13965,N_10454,N_12281);
and U13966 (N_13966,N_11205,N_11945);
and U13967 (N_13967,N_9507,N_10201);
nand U13968 (N_13968,N_10010,N_10290);
nand U13969 (N_13969,N_9531,N_9551);
and U13970 (N_13970,N_10112,N_11226);
nor U13971 (N_13971,N_9791,N_12189);
nor U13972 (N_13972,N_11444,N_10806);
or U13973 (N_13973,N_10068,N_9467);
nor U13974 (N_13974,N_11652,N_12183);
or U13975 (N_13975,N_10753,N_9640);
and U13976 (N_13976,N_11789,N_11936);
nor U13977 (N_13977,N_9797,N_11862);
or U13978 (N_13978,N_9841,N_12276);
or U13979 (N_13979,N_11393,N_12485);
nand U13980 (N_13980,N_11292,N_10502);
nand U13981 (N_13981,N_10099,N_10208);
and U13982 (N_13982,N_9763,N_9599);
nand U13983 (N_13983,N_11518,N_12439);
and U13984 (N_13984,N_11122,N_11192);
xor U13985 (N_13985,N_10063,N_12025);
and U13986 (N_13986,N_9838,N_11905);
nor U13987 (N_13987,N_9936,N_9971);
nand U13988 (N_13988,N_10666,N_11102);
nor U13989 (N_13989,N_10697,N_11119);
or U13990 (N_13990,N_10606,N_9877);
or U13991 (N_13991,N_11857,N_9871);
or U13992 (N_13992,N_10240,N_9552);
xor U13993 (N_13993,N_11539,N_12074);
nand U13994 (N_13994,N_11926,N_12108);
and U13995 (N_13995,N_9508,N_12199);
nand U13996 (N_13996,N_12067,N_11950);
nor U13997 (N_13997,N_11341,N_11728);
nor U13998 (N_13998,N_9593,N_10389);
and U13999 (N_13999,N_11568,N_10532);
or U14000 (N_14000,N_12121,N_9629);
nor U14001 (N_14001,N_11020,N_11033);
nand U14002 (N_14002,N_9667,N_10381);
and U14003 (N_14003,N_11829,N_11410);
and U14004 (N_14004,N_10598,N_11129);
or U14005 (N_14005,N_10773,N_12454);
nand U14006 (N_14006,N_10604,N_10937);
nand U14007 (N_14007,N_11380,N_12315);
and U14008 (N_14008,N_10599,N_12224);
or U14009 (N_14009,N_11556,N_12041);
and U14010 (N_14010,N_10647,N_10612);
or U14011 (N_14011,N_10970,N_9770);
and U14012 (N_14012,N_9455,N_10559);
or U14013 (N_14013,N_12111,N_10851);
xor U14014 (N_14014,N_11899,N_11649);
nand U14015 (N_14015,N_11342,N_10944);
xnor U14016 (N_14016,N_11359,N_12314);
nor U14017 (N_14017,N_11643,N_12415);
nand U14018 (N_14018,N_10065,N_9416);
nor U14019 (N_14019,N_10245,N_12212);
and U14020 (N_14020,N_9925,N_11955);
and U14021 (N_14021,N_9873,N_10868);
or U14022 (N_14022,N_12040,N_9856);
nor U14023 (N_14023,N_12427,N_10025);
or U14024 (N_14024,N_11406,N_10355);
xor U14025 (N_14025,N_9833,N_11934);
nand U14026 (N_14026,N_11686,N_10313);
and U14027 (N_14027,N_11010,N_11661);
or U14028 (N_14028,N_10190,N_9757);
nand U14029 (N_14029,N_10125,N_11203);
and U14030 (N_14030,N_10721,N_9887);
nand U14031 (N_14031,N_10145,N_10875);
xor U14032 (N_14032,N_11573,N_9822);
or U14033 (N_14033,N_11971,N_11736);
xnor U14034 (N_14034,N_11267,N_11785);
nor U14035 (N_14035,N_10603,N_9819);
nand U14036 (N_14036,N_10813,N_10319);
or U14037 (N_14037,N_10707,N_10033);
and U14038 (N_14038,N_11904,N_10739);
or U14039 (N_14039,N_10682,N_10277);
and U14040 (N_14040,N_9709,N_9434);
and U14041 (N_14041,N_9749,N_10641);
and U14042 (N_14042,N_10079,N_10638);
nand U14043 (N_14043,N_12363,N_10713);
or U14044 (N_14044,N_10801,N_11399);
nor U14045 (N_14045,N_11567,N_10430);
nand U14046 (N_14046,N_11816,N_11693);
or U14047 (N_14047,N_11168,N_12000);
nand U14048 (N_14048,N_11932,N_10850);
xor U14049 (N_14049,N_9479,N_10186);
nand U14050 (N_14050,N_11705,N_12319);
and U14051 (N_14051,N_9627,N_10651);
and U14052 (N_14052,N_10917,N_12286);
nor U14053 (N_14053,N_10041,N_10242);
and U14054 (N_14054,N_10157,N_11602);
and U14055 (N_14055,N_9837,N_10446);
and U14056 (N_14056,N_11477,N_9771);
nand U14057 (N_14057,N_12061,N_10849);
xnor U14058 (N_14058,N_10918,N_11247);
nand U14059 (N_14059,N_11151,N_10045);
or U14060 (N_14060,N_9657,N_12109);
nor U14061 (N_14061,N_12263,N_9402);
nor U14062 (N_14062,N_10630,N_9794);
nor U14063 (N_14063,N_9848,N_12141);
xnor U14064 (N_14064,N_12122,N_9447);
and U14065 (N_14065,N_11459,N_11467);
nand U14066 (N_14066,N_11546,N_11008);
nand U14067 (N_14067,N_12463,N_9397);
or U14068 (N_14068,N_10463,N_11137);
or U14069 (N_14069,N_10653,N_11660);
or U14070 (N_14070,N_9504,N_12134);
nor U14071 (N_14071,N_12441,N_11706);
xor U14072 (N_14072,N_10742,N_10104);
and U14073 (N_14073,N_10295,N_11812);
and U14074 (N_14074,N_12100,N_11753);
nand U14075 (N_14075,N_12306,N_9578);
nor U14076 (N_14076,N_12350,N_10299);
nor U14077 (N_14077,N_11015,N_11272);
and U14078 (N_14078,N_10502,N_9671);
nand U14079 (N_14079,N_10940,N_10124);
nand U14080 (N_14080,N_9391,N_11783);
xnor U14081 (N_14081,N_9598,N_10146);
xnor U14082 (N_14082,N_10851,N_12015);
and U14083 (N_14083,N_9931,N_9747);
or U14084 (N_14084,N_11069,N_11584);
nand U14085 (N_14085,N_10614,N_9981);
or U14086 (N_14086,N_11801,N_12088);
or U14087 (N_14087,N_11276,N_10677);
and U14088 (N_14088,N_11033,N_9629);
xnor U14089 (N_14089,N_10394,N_9958);
nand U14090 (N_14090,N_10230,N_11472);
and U14091 (N_14091,N_9689,N_10066);
or U14092 (N_14092,N_10952,N_10268);
nand U14093 (N_14093,N_10264,N_11513);
or U14094 (N_14094,N_10557,N_10536);
nor U14095 (N_14095,N_9843,N_9547);
or U14096 (N_14096,N_10421,N_11730);
or U14097 (N_14097,N_10031,N_9895);
or U14098 (N_14098,N_11434,N_9874);
xor U14099 (N_14099,N_9390,N_11194);
nor U14100 (N_14100,N_12227,N_10736);
nor U14101 (N_14101,N_9524,N_10753);
or U14102 (N_14102,N_12363,N_9749);
nor U14103 (N_14103,N_10559,N_12204);
and U14104 (N_14104,N_11564,N_10743);
and U14105 (N_14105,N_9823,N_10325);
or U14106 (N_14106,N_10235,N_11011);
or U14107 (N_14107,N_11619,N_10407);
or U14108 (N_14108,N_12234,N_10018);
nor U14109 (N_14109,N_9537,N_10862);
nor U14110 (N_14110,N_10343,N_9497);
or U14111 (N_14111,N_9723,N_10709);
nand U14112 (N_14112,N_10999,N_10478);
nor U14113 (N_14113,N_9921,N_10717);
nand U14114 (N_14114,N_11761,N_10191);
and U14115 (N_14115,N_12034,N_11590);
nor U14116 (N_14116,N_9708,N_10046);
nand U14117 (N_14117,N_11698,N_12023);
xor U14118 (N_14118,N_12149,N_12171);
nand U14119 (N_14119,N_10675,N_9669);
nand U14120 (N_14120,N_9748,N_11272);
nor U14121 (N_14121,N_10619,N_11926);
nand U14122 (N_14122,N_12249,N_9615);
nand U14123 (N_14123,N_9384,N_10944);
or U14124 (N_14124,N_12368,N_9483);
and U14125 (N_14125,N_11434,N_12431);
or U14126 (N_14126,N_9639,N_10466);
nand U14127 (N_14127,N_10244,N_11738);
xnor U14128 (N_14128,N_9895,N_10587);
and U14129 (N_14129,N_10794,N_11904);
nor U14130 (N_14130,N_9737,N_10485);
nor U14131 (N_14131,N_9559,N_9557);
and U14132 (N_14132,N_10622,N_11996);
and U14133 (N_14133,N_11854,N_11077);
or U14134 (N_14134,N_11775,N_10326);
xnor U14135 (N_14135,N_10758,N_10935);
and U14136 (N_14136,N_9451,N_9378);
or U14137 (N_14137,N_10889,N_9965);
and U14138 (N_14138,N_10317,N_10561);
and U14139 (N_14139,N_12218,N_11419);
nand U14140 (N_14140,N_9804,N_10719);
and U14141 (N_14141,N_11961,N_10316);
and U14142 (N_14142,N_9471,N_10050);
and U14143 (N_14143,N_11211,N_11395);
nand U14144 (N_14144,N_11831,N_9582);
or U14145 (N_14145,N_10688,N_11705);
nand U14146 (N_14146,N_12012,N_9968);
nand U14147 (N_14147,N_11898,N_12095);
nand U14148 (N_14148,N_9809,N_10349);
nand U14149 (N_14149,N_9853,N_11238);
xnor U14150 (N_14150,N_12348,N_9887);
nand U14151 (N_14151,N_11171,N_10388);
or U14152 (N_14152,N_9445,N_12319);
nor U14153 (N_14153,N_9519,N_12138);
or U14154 (N_14154,N_10732,N_11785);
and U14155 (N_14155,N_10529,N_9533);
nand U14156 (N_14156,N_10915,N_12371);
nor U14157 (N_14157,N_10490,N_9954);
nor U14158 (N_14158,N_9460,N_9931);
nor U14159 (N_14159,N_12250,N_10317);
nand U14160 (N_14160,N_10683,N_9376);
and U14161 (N_14161,N_11237,N_10634);
nand U14162 (N_14162,N_12111,N_10096);
or U14163 (N_14163,N_10176,N_10780);
and U14164 (N_14164,N_12245,N_12119);
and U14165 (N_14165,N_11814,N_11354);
or U14166 (N_14166,N_11455,N_11191);
and U14167 (N_14167,N_10700,N_10663);
and U14168 (N_14168,N_10335,N_11558);
nor U14169 (N_14169,N_12229,N_9726);
nor U14170 (N_14170,N_11124,N_9496);
nand U14171 (N_14171,N_11092,N_12320);
or U14172 (N_14172,N_10575,N_11034);
and U14173 (N_14173,N_10295,N_12159);
nor U14174 (N_14174,N_11045,N_10948);
or U14175 (N_14175,N_11222,N_11443);
nand U14176 (N_14176,N_10708,N_11706);
nand U14177 (N_14177,N_11174,N_11699);
nand U14178 (N_14178,N_10318,N_9450);
or U14179 (N_14179,N_12053,N_9487);
xor U14180 (N_14180,N_11244,N_9735);
nor U14181 (N_14181,N_10826,N_10930);
nand U14182 (N_14182,N_10925,N_11915);
xnor U14183 (N_14183,N_12484,N_11741);
and U14184 (N_14184,N_10035,N_10802);
and U14185 (N_14185,N_10563,N_9551);
and U14186 (N_14186,N_11918,N_12429);
and U14187 (N_14187,N_12499,N_9895);
nand U14188 (N_14188,N_10117,N_11111);
nor U14189 (N_14189,N_10046,N_9659);
or U14190 (N_14190,N_11337,N_9866);
nand U14191 (N_14191,N_11582,N_11647);
nor U14192 (N_14192,N_9866,N_11771);
or U14193 (N_14193,N_10352,N_10698);
or U14194 (N_14194,N_12052,N_10226);
and U14195 (N_14195,N_10364,N_10263);
and U14196 (N_14196,N_11633,N_10669);
or U14197 (N_14197,N_10320,N_11105);
nand U14198 (N_14198,N_12258,N_9470);
nor U14199 (N_14199,N_10341,N_11754);
nor U14200 (N_14200,N_11172,N_11679);
and U14201 (N_14201,N_11102,N_9727);
xor U14202 (N_14202,N_10568,N_10304);
xnor U14203 (N_14203,N_12008,N_11784);
or U14204 (N_14204,N_10577,N_11309);
nor U14205 (N_14205,N_9810,N_10477);
xnor U14206 (N_14206,N_11257,N_10830);
and U14207 (N_14207,N_10955,N_9807);
or U14208 (N_14208,N_11528,N_11286);
or U14209 (N_14209,N_9501,N_11948);
and U14210 (N_14210,N_11678,N_11309);
nand U14211 (N_14211,N_11954,N_11002);
xor U14212 (N_14212,N_11367,N_10772);
or U14213 (N_14213,N_11024,N_11643);
and U14214 (N_14214,N_12265,N_9999);
nand U14215 (N_14215,N_11567,N_12151);
and U14216 (N_14216,N_9936,N_9403);
nand U14217 (N_14217,N_12266,N_11752);
nor U14218 (N_14218,N_11266,N_11943);
nor U14219 (N_14219,N_12437,N_11653);
or U14220 (N_14220,N_9808,N_9636);
and U14221 (N_14221,N_9575,N_11337);
and U14222 (N_14222,N_12344,N_9778);
or U14223 (N_14223,N_11051,N_9955);
xnor U14224 (N_14224,N_11318,N_10260);
and U14225 (N_14225,N_11307,N_11540);
nor U14226 (N_14226,N_10485,N_11232);
or U14227 (N_14227,N_10085,N_10635);
nand U14228 (N_14228,N_10657,N_12114);
xnor U14229 (N_14229,N_12463,N_12415);
nand U14230 (N_14230,N_12353,N_10650);
xor U14231 (N_14231,N_11306,N_11967);
and U14232 (N_14232,N_11186,N_11876);
nor U14233 (N_14233,N_11612,N_10623);
and U14234 (N_14234,N_9474,N_11217);
and U14235 (N_14235,N_12320,N_11872);
xor U14236 (N_14236,N_9487,N_11787);
nand U14237 (N_14237,N_11855,N_10912);
or U14238 (N_14238,N_11000,N_9379);
xor U14239 (N_14239,N_12258,N_11363);
and U14240 (N_14240,N_11211,N_12007);
nor U14241 (N_14241,N_11198,N_11464);
xor U14242 (N_14242,N_10948,N_12067);
nand U14243 (N_14243,N_10913,N_9730);
nand U14244 (N_14244,N_10927,N_11748);
or U14245 (N_14245,N_9807,N_10204);
nand U14246 (N_14246,N_11257,N_11804);
or U14247 (N_14247,N_9964,N_9436);
or U14248 (N_14248,N_10945,N_10621);
nor U14249 (N_14249,N_9970,N_10548);
nand U14250 (N_14250,N_10414,N_10637);
and U14251 (N_14251,N_10931,N_11481);
and U14252 (N_14252,N_11415,N_9980);
and U14253 (N_14253,N_10589,N_10487);
and U14254 (N_14254,N_9416,N_10572);
nand U14255 (N_14255,N_11909,N_11121);
xor U14256 (N_14256,N_11679,N_12294);
or U14257 (N_14257,N_12418,N_11115);
and U14258 (N_14258,N_10687,N_9438);
nor U14259 (N_14259,N_10000,N_11846);
nor U14260 (N_14260,N_11281,N_11834);
and U14261 (N_14261,N_11727,N_9724);
xor U14262 (N_14262,N_9668,N_10723);
nor U14263 (N_14263,N_10887,N_10244);
and U14264 (N_14264,N_11785,N_11226);
nor U14265 (N_14265,N_10505,N_10438);
xor U14266 (N_14266,N_10534,N_12308);
or U14267 (N_14267,N_11425,N_9414);
nor U14268 (N_14268,N_12135,N_9778);
nand U14269 (N_14269,N_10712,N_11191);
or U14270 (N_14270,N_12021,N_9523);
nand U14271 (N_14271,N_11259,N_9572);
and U14272 (N_14272,N_12174,N_10935);
and U14273 (N_14273,N_10982,N_12047);
nor U14274 (N_14274,N_12063,N_12333);
or U14275 (N_14275,N_11119,N_12001);
nor U14276 (N_14276,N_11013,N_10319);
and U14277 (N_14277,N_11435,N_12319);
nor U14278 (N_14278,N_10220,N_12403);
or U14279 (N_14279,N_11078,N_10881);
nor U14280 (N_14280,N_11560,N_10418);
or U14281 (N_14281,N_9402,N_11528);
or U14282 (N_14282,N_9769,N_11275);
and U14283 (N_14283,N_9774,N_9425);
and U14284 (N_14284,N_12464,N_12128);
nor U14285 (N_14285,N_11539,N_12419);
nand U14286 (N_14286,N_11511,N_10639);
and U14287 (N_14287,N_11491,N_12142);
xor U14288 (N_14288,N_9627,N_11955);
and U14289 (N_14289,N_12060,N_11217);
xor U14290 (N_14290,N_11982,N_9980);
and U14291 (N_14291,N_12095,N_10160);
nor U14292 (N_14292,N_11671,N_9961);
nor U14293 (N_14293,N_11167,N_10092);
nor U14294 (N_14294,N_10297,N_11588);
nor U14295 (N_14295,N_9984,N_10883);
nor U14296 (N_14296,N_12027,N_12166);
nand U14297 (N_14297,N_11366,N_12400);
and U14298 (N_14298,N_10916,N_11230);
nand U14299 (N_14299,N_11246,N_11635);
nor U14300 (N_14300,N_12094,N_10273);
or U14301 (N_14301,N_11664,N_11537);
xnor U14302 (N_14302,N_11720,N_10363);
xnor U14303 (N_14303,N_10630,N_9735);
or U14304 (N_14304,N_11279,N_10828);
nor U14305 (N_14305,N_10990,N_10687);
nor U14306 (N_14306,N_11065,N_10588);
nor U14307 (N_14307,N_11801,N_10155);
xor U14308 (N_14308,N_9620,N_9896);
and U14309 (N_14309,N_11491,N_11310);
nor U14310 (N_14310,N_10593,N_10936);
nand U14311 (N_14311,N_11462,N_12323);
and U14312 (N_14312,N_11642,N_11854);
nor U14313 (N_14313,N_10300,N_10949);
nor U14314 (N_14314,N_11615,N_10203);
and U14315 (N_14315,N_9927,N_10641);
and U14316 (N_14316,N_11416,N_11816);
nor U14317 (N_14317,N_11789,N_11210);
or U14318 (N_14318,N_10255,N_10235);
or U14319 (N_14319,N_11114,N_12244);
nor U14320 (N_14320,N_11586,N_12368);
nor U14321 (N_14321,N_12255,N_9825);
and U14322 (N_14322,N_11210,N_10888);
nor U14323 (N_14323,N_11537,N_10826);
nor U14324 (N_14324,N_12174,N_12429);
xnor U14325 (N_14325,N_11913,N_12471);
nand U14326 (N_14326,N_9632,N_11975);
nor U14327 (N_14327,N_9591,N_11281);
or U14328 (N_14328,N_9786,N_9724);
or U14329 (N_14329,N_9684,N_10469);
and U14330 (N_14330,N_12321,N_12058);
nand U14331 (N_14331,N_11878,N_10630);
nand U14332 (N_14332,N_11502,N_9860);
nand U14333 (N_14333,N_9501,N_10408);
nand U14334 (N_14334,N_11129,N_11311);
or U14335 (N_14335,N_10010,N_9898);
or U14336 (N_14336,N_10711,N_10332);
and U14337 (N_14337,N_11760,N_9922);
or U14338 (N_14338,N_11360,N_11175);
nor U14339 (N_14339,N_9466,N_11654);
nand U14340 (N_14340,N_10628,N_9970);
or U14341 (N_14341,N_11958,N_10198);
and U14342 (N_14342,N_11754,N_9718);
nand U14343 (N_14343,N_12124,N_10292);
xnor U14344 (N_14344,N_12491,N_11000);
or U14345 (N_14345,N_11400,N_11545);
and U14346 (N_14346,N_10845,N_9499);
nand U14347 (N_14347,N_10416,N_11938);
and U14348 (N_14348,N_11662,N_9657);
nor U14349 (N_14349,N_9716,N_10292);
nor U14350 (N_14350,N_12259,N_9428);
and U14351 (N_14351,N_11644,N_10778);
and U14352 (N_14352,N_11832,N_11931);
xor U14353 (N_14353,N_11109,N_10146);
and U14354 (N_14354,N_11348,N_10353);
nand U14355 (N_14355,N_10293,N_11886);
nor U14356 (N_14356,N_12085,N_10017);
or U14357 (N_14357,N_9855,N_9869);
nand U14358 (N_14358,N_10482,N_10932);
or U14359 (N_14359,N_11224,N_9923);
nor U14360 (N_14360,N_9699,N_9383);
and U14361 (N_14361,N_11985,N_9703);
nor U14362 (N_14362,N_11966,N_10821);
or U14363 (N_14363,N_9753,N_12402);
or U14364 (N_14364,N_9653,N_12263);
nand U14365 (N_14365,N_12171,N_9417);
and U14366 (N_14366,N_11264,N_10449);
nand U14367 (N_14367,N_12111,N_11291);
and U14368 (N_14368,N_11885,N_12433);
and U14369 (N_14369,N_9967,N_10680);
nor U14370 (N_14370,N_10161,N_9622);
nand U14371 (N_14371,N_10147,N_10992);
or U14372 (N_14372,N_11673,N_11590);
and U14373 (N_14373,N_11964,N_9895);
or U14374 (N_14374,N_9964,N_10835);
and U14375 (N_14375,N_9636,N_11796);
and U14376 (N_14376,N_9740,N_9725);
nand U14377 (N_14377,N_12055,N_10496);
nor U14378 (N_14378,N_11074,N_11280);
and U14379 (N_14379,N_11115,N_11398);
or U14380 (N_14380,N_11389,N_9648);
nor U14381 (N_14381,N_11156,N_10876);
nand U14382 (N_14382,N_9848,N_11754);
and U14383 (N_14383,N_12107,N_9705);
and U14384 (N_14384,N_11435,N_12478);
nand U14385 (N_14385,N_10830,N_9977);
and U14386 (N_14386,N_9757,N_11409);
or U14387 (N_14387,N_12000,N_12345);
nor U14388 (N_14388,N_12248,N_12173);
or U14389 (N_14389,N_11992,N_9783);
and U14390 (N_14390,N_10322,N_9944);
xnor U14391 (N_14391,N_11100,N_10775);
nor U14392 (N_14392,N_9385,N_11740);
and U14393 (N_14393,N_12273,N_10350);
and U14394 (N_14394,N_12175,N_11246);
and U14395 (N_14395,N_10805,N_12025);
and U14396 (N_14396,N_11393,N_10854);
or U14397 (N_14397,N_11125,N_10970);
or U14398 (N_14398,N_11619,N_10341);
nand U14399 (N_14399,N_11850,N_10265);
xor U14400 (N_14400,N_9621,N_9858);
nor U14401 (N_14401,N_9695,N_12161);
nand U14402 (N_14402,N_10721,N_9592);
and U14403 (N_14403,N_10743,N_12239);
or U14404 (N_14404,N_9974,N_10486);
or U14405 (N_14405,N_11500,N_10495);
nand U14406 (N_14406,N_9955,N_10951);
nor U14407 (N_14407,N_9818,N_11285);
or U14408 (N_14408,N_11438,N_10165);
nand U14409 (N_14409,N_10068,N_10034);
nor U14410 (N_14410,N_11315,N_9475);
and U14411 (N_14411,N_10983,N_11528);
nor U14412 (N_14412,N_11286,N_9601);
nor U14413 (N_14413,N_12026,N_9625);
nor U14414 (N_14414,N_10830,N_12389);
nor U14415 (N_14415,N_10206,N_12387);
and U14416 (N_14416,N_11996,N_10773);
or U14417 (N_14417,N_9766,N_9382);
nand U14418 (N_14418,N_12198,N_11285);
and U14419 (N_14419,N_9747,N_10613);
nand U14420 (N_14420,N_12389,N_11229);
nand U14421 (N_14421,N_11767,N_11843);
or U14422 (N_14422,N_11112,N_9710);
xor U14423 (N_14423,N_10482,N_10417);
or U14424 (N_14424,N_11299,N_10832);
and U14425 (N_14425,N_10810,N_9620);
or U14426 (N_14426,N_9616,N_10175);
and U14427 (N_14427,N_11717,N_9720);
or U14428 (N_14428,N_10441,N_11061);
and U14429 (N_14429,N_12408,N_12436);
nand U14430 (N_14430,N_11734,N_11246);
nor U14431 (N_14431,N_10533,N_12423);
nand U14432 (N_14432,N_12392,N_10290);
or U14433 (N_14433,N_11447,N_12428);
nor U14434 (N_14434,N_12414,N_10981);
or U14435 (N_14435,N_9619,N_10551);
and U14436 (N_14436,N_9427,N_11170);
nand U14437 (N_14437,N_12407,N_11101);
xor U14438 (N_14438,N_11426,N_11337);
nor U14439 (N_14439,N_10226,N_9784);
and U14440 (N_14440,N_11444,N_11782);
and U14441 (N_14441,N_10274,N_11159);
or U14442 (N_14442,N_12498,N_11240);
nand U14443 (N_14443,N_9727,N_10475);
and U14444 (N_14444,N_10897,N_11706);
nand U14445 (N_14445,N_9461,N_12228);
and U14446 (N_14446,N_9735,N_11744);
nor U14447 (N_14447,N_9812,N_12145);
nand U14448 (N_14448,N_12048,N_9965);
nor U14449 (N_14449,N_9478,N_10004);
xnor U14450 (N_14450,N_10404,N_11317);
or U14451 (N_14451,N_12415,N_10063);
xor U14452 (N_14452,N_9795,N_11292);
and U14453 (N_14453,N_12331,N_9974);
nor U14454 (N_14454,N_11795,N_10852);
nor U14455 (N_14455,N_9767,N_11214);
nor U14456 (N_14456,N_10484,N_11254);
xor U14457 (N_14457,N_10140,N_12201);
nand U14458 (N_14458,N_10230,N_11519);
xor U14459 (N_14459,N_10200,N_12331);
or U14460 (N_14460,N_12018,N_12393);
nand U14461 (N_14461,N_10264,N_9575);
nor U14462 (N_14462,N_11413,N_9526);
nand U14463 (N_14463,N_12411,N_9563);
nand U14464 (N_14464,N_10475,N_11915);
nand U14465 (N_14465,N_11875,N_11511);
nor U14466 (N_14466,N_11749,N_12096);
and U14467 (N_14467,N_9573,N_11185);
nor U14468 (N_14468,N_9846,N_9912);
nand U14469 (N_14469,N_12023,N_10946);
xnor U14470 (N_14470,N_11552,N_10642);
and U14471 (N_14471,N_10247,N_11061);
nor U14472 (N_14472,N_10616,N_9465);
or U14473 (N_14473,N_12141,N_12321);
nor U14474 (N_14474,N_12244,N_11648);
or U14475 (N_14475,N_12206,N_12177);
xor U14476 (N_14476,N_11551,N_11852);
and U14477 (N_14477,N_11378,N_9912);
and U14478 (N_14478,N_9578,N_10526);
nand U14479 (N_14479,N_11683,N_9980);
nor U14480 (N_14480,N_9761,N_9682);
nand U14481 (N_14481,N_10981,N_9834);
xor U14482 (N_14482,N_11639,N_11925);
nor U14483 (N_14483,N_11088,N_11899);
and U14484 (N_14484,N_12024,N_11585);
xor U14485 (N_14485,N_12014,N_10595);
and U14486 (N_14486,N_12316,N_10895);
or U14487 (N_14487,N_12099,N_11046);
nor U14488 (N_14488,N_10547,N_12114);
or U14489 (N_14489,N_12169,N_12109);
and U14490 (N_14490,N_11888,N_11092);
nor U14491 (N_14491,N_12484,N_10168);
nand U14492 (N_14492,N_10859,N_11730);
nand U14493 (N_14493,N_10795,N_12166);
nand U14494 (N_14494,N_11846,N_11988);
and U14495 (N_14495,N_9784,N_11454);
nor U14496 (N_14496,N_9755,N_12430);
or U14497 (N_14497,N_11846,N_10675);
nor U14498 (N_14498,N_10178,N_10622);
and U14499 (N_14499,N_9620,N_11258);
or U14500 (N_14500,N_11379,N_11260);
and U14501 (N_14501,N_12028,N_10977);
nor U14502 (N_14502,N_11535,N_10021);
and U14503 (N_14503,N_10349,N_10084);
and U14504 (N_14504,N_10052,N_10419);
nand U14505 (N_14505,N_11401,N_10424);
nor U14506 (N_14506,N_11923,N_10558);
nor U14507 (N_14507,N_10773,N_12402);
and U14508 (N_14508,N_9388,N_11187);
or U14509 (N_14509,N_12176,N_10347);
nor U14510 (N_14510,N_10745,N_11491);
xnor U14511 (N_14511,N_10532,N_11311);
and U14512 (N_14512,N_9427,N_12410);
nand U14513 (N_14513,N_9827,N_10379);
or U14514 (N_14514,N_12186,N_11970);
and U14515 (N_14515,N_11858,N_10660);
nand U14516 (N_14516,N_10085,N_11401);
or U14517 (N_14517,N_11495,N_11552);
or U14518 (N_14518,N_11327,N_12228);
nor U14519 (N_14519,N_11296,N_11742);
or U14520 (N_14520,N_11141,N_11021);
nor U14521 (N_14521,N_9914,N_10156);
nand U14522 (N_14522,N_9814,N_10537);
nand U14523 (N_14523,N_10488,N_11258);
nor U14524 (N_14524,N_11790,N_10728);
or U14525 (N_14525,N_11387,N_10849);
nand U14526 (N_14526,N_12214,N_9772);
and U14527 (N_14527,N_12324,N_12486);
nor U14528 (N_14528,N_11694,N_9552);
or U14529 (N_14529,N_11700,N_10140);
and U14530 (N_14530,N_10650,N_10114);
xor U14531 (N_14531,N_12315,N_9876);
xnor U14532 (N_14532,N_10815,N_10263);
or U14533 (N_14533,N_11953,N_11839);
nor U14534 (N_14534,N_10545,N_11376);
nor U14535 (N_14535,N_10061,N_9929);
nand U14536 (N_14536,N_12201,N_10405);
nor U14537 (N_14537,N_11709,N_11568);
or U14538 (N_14538,N_11583,N_10756);
xor U14539 (N_14539,N_11745,N_10189);
or U14540 (N_14540,N_11740,N_11137);
nand U14541 (N_14541,N_10021,N_12487);
or U14542 (N_14542,N_9700,N_11394);
or U14543 (N_14543,N_9809,N_9676);
or U14544 (N_14544,N_9593,N_9784);
or U14545 (N_14545,N_9631,N_11744);
or U14546 (N_14546,N_11107,N_11112);
and U14547 (N_14547,N_10295,N_11834);
nor U14548 (N_14548,N_12302,N_11299);
nor U14549 (N_14549,N_12011,N_10743);
and U14550 (N_14550,N_10451,N_11049);
or U14551 (N_14551,N_10288,N_11616);
and U14552 (N_14552,N_11363,N_10032);
xor U14553 (N_14553,N_12038,N_12002);
and U14554 (N_14554,N_10090,N_10062);
or U14555 (N_14555,N_10707,N_11209);
or U14556 (N_14556,N_10202,N_9700);
nand U14557 (N_14557,N_10898,N_10376);
nand U14558 (N_14558,N_11687,N_10762);
xor U14559 (N_14559,N_11198,N_11125);
or U14560 (N_14560,N_11257,N_11123);
or U14561 (N_14561,N_11860,N_9743);
nor U14562 (N_14562,N_10903,N_9512);
nand U14563 (N_14563,N_10563,N_10152);
xnor U14564 (N_14564,N_11071,N_12246);
and U14565 (N_14565,N_10409,N_10712);
nand U14566 (N_14566,N_9644,N_9582);
nor U14567 (N_14567,N_10392,N_9405);
or U14568 (N_14568,N_11450,N_10498);
xor U14569 (N_14569,N_11285,N_10336);
and U14570 (N_14570,N_11207,N_11341);
and U14571 (N_14571,N_10634,N_12056);
nor U14572 (N_14572,N_10783,N_12338);
or U14573 (N_14573,N_9844,N_12235);
nand U14574 (N_14574,N_10185,N_12108);
and U14575 (N_14575,N_10638,N_9677);
or U14576 (N_14576,N_9599,N_12111);
or U14577 (N_14577,N_11218,N_12048);
and U14578 (N_14578,N_9782,N_11191);
xor U14579 (N_14579,N_10323,N_11666);
or U14580 (N_14580,N_12343,N_11309);
xor U14581 (N_14581,N_11162,N_11595);
and U14582 (N_14582,N_9495,N_10293);
xnor U14583 (N_14583,N_12265,N_10287);
and U14584 (N_14584,N_9721,N_11381);
or U14585 (N_14585,N_9881,N_9878);
or U14586 (N_14586,N_12257,N_10057);
nor U14587 (N_14587,N_11028,N_11808);
nand U14588 (N_14588,N_11172,N_10248);
xnor U14589 (N_14589,N_11938,N_11386);
or U14590 (N_14590,N_10549,N_12143);
nand U14591 (N_14591,N_11032,N_12121);
nor U14592 (N_14592,N_12259,N_9873);
or U14593 (N_14593,N_11585,N_9960);
or U14594 (N_14594,N_10679,N_9887);
and U14595 (N_14595,N_9849,N_10992);
nand U14596 (N_14596,N_9512,N_9429);
and U14597 (N_14597,N_11197,N_12328);
and U14598 (N_14598,N_11436,N_11998);
nor U14599 (N_14599,N_12010,N_10715);
xnor U14600 (N_14600,N_12168,N_9635);
nand U14601 (N_14601,N_10333,N_12403);
xor U14602 (N_14602,N_12156,N_10371);
or U14603 (N_14603,N_10356,N_11293);
xor U14604 (N_14604,N_11739,N_11586);
nand U14605 (N_14605,N_11714,N_10928);
or U14606 (N_14606,N_10501,N_11977);
nor U14607 (N_14607,N_11646,N_11123);
or U14608 (N_14608,N_10420,N_10445);
and U14609 (N_14609,N_9606,N_11068);
xnor U14610 (N_14610,N_9775,N_9993);
xnor U14611 (N_14611,N_10055,N_10842);
nand U14612 (N_14612,N_9805,N_11080);
nor U14613 (N_14613,N_9606,N_10191);
nor U14614 (N_14614,N_12154,N_12127);
and U14615 (N_14615,N_11869,N_10835);
xnor U14616 (N_14616,N_11564,N_11653);
and U14617 (N_14617,N_10076,N_9616);
nand U14618 (N_14618,N_10743,N_9848);
and U14619 (N_14619,N_12494,N_11654);
nand U14620 (N_14620,N_10874,N_9719);
and U14621 (N_14621,N_11433,N_10475);
nand U14622 (N_14622,N_9712,N_12357);
and U14623 (N_14623,N_10939,N_11215);
xor U14624 (N_14624,N_9847,N_11757);
nor U14625 (N_14625,N_10124,N_10347);
nor U14626 (N_14626,N_11110,N_10959);
and U14627 (N_14627,N_11184,N_11218);
nand U14628 (N_14628,N_10092,N_10267);
or U14629 (N_14629,N_10204,N_11179);
nand U14630 (N_14630,N_9896,N_12392);
nor U14631 (N_14631,N_11458,N_10508);
nor U14632 (N_14632,N_12441,N_10832);
or U14633 (N_14633,N_12252,N_10130);
or U14634 (N_14634,N_12483,N_10113);
and U14635 (N_14635,N_12248,N_12038);
nor U14636 (N_14636,N_10436,N_11571);
or U14637 (N_14637,N_10021,N_10476);
or U14638 (N_14638,N_10456,N_10535);
nand U14639 (N_14639,N_12443,N_11894);
nand U14640 (N_14640,N_12024,N_11472);
and U14641 (N_14641,N_10566,N_11622);
xor U14642 (N_14642,N_11882,N_11032);
or U14643 (N_14643,N_11229,N_9636);
and U14644 (N_14644,N_11302,N_11214);
or U14645 (N_14645,N_9898,N_11206);
and U14646 (N_14646,N_12442,N_10689);
and U14647 (N_14647,N_11283,N_11854);
nand U14648 (N_14648,N_11529,N_11768);
or U14649 (N_14649,N_10750,N_11321);
nor U14650 (N_14650,N_11503,N_11329);
nand U14651 (N_14651,N_12447,N_11311);
or U14652 (N_14652,N_10261,N_10614);
nand U14653 (N_14653,N_9587,N_11145);
nor U14654 (N_14654,N_11039,N_10575);
xnor U14655 (N_14655,N_9599,N_9463);
or U14656 (N_14656,N_12243,N_10228);
and U14657 (N_14657,N_10215,N_11635);
xnor U14658 (N_14658,N_11077,N_9731);
xor U14659 (N_14659,N_10253,N_9662);
xnor U14660 (N_14660,N_12057,N_10913);
or U14661 (N_14661,N_12049,N_10468);
nor U14662 (N_14662,N_10215,N_12169);
nor U14663 (N_14663,N_9455,N_11152);
and U14664 (N_14664,N_10843,N_10496);
or U14665 (N_14665,N_10182,N_10240);
and U14666 (N_14666,N_11084,N_9396);
or U14667 (N_14667,N_11264,N_9788);
nand U14668 (N_14668,N_11401,N_9661);
xor U14669 (N_14669,N_12105,N_12319);
or U14670 (N_14670,N_11350,N_11011);
or U14671 (N_14671,N_9827,N_10926);
and U14672 (N_14672,N_10105,N_10123);
nand U14673 (N_14673,N_11404,N_12226);
nand U14674 (N_14674,N_11937,N_10234);
or U14675 (N_14675,N_9955,N_11171);
nand U14676 (N_14676,N_11228,N_12317);
or U14677 (N_14677,N_11099,N_11687);
nor U14678 (N_14678,N_12254,N_12115);
nor U14679 (N_14679,N_9484,N_11387);
nand U14680 (N_14680,N_12479,N_10922);
and U14681 (N_14681,N_12244,N_11357);
nand U14682 (N_14682,N_11126,N_11805);
and U14683 (N_14683,N_11057,N_10735);
and U14684 (N_14684,N_9581,N_10718);
and U14685 (N_14685,N_10120,N_12152);
xnor U14686 (N_14686,N_11033,N_12234);
xnor U14687 (N_14687,N_12069,N_9868);
nor U14688 (N_14688,N_10612,N_12179);
and U14689 (N_14689,N_12401,N_9539);
and U14690 (N_14690,N_12295,N_11427);
or U14691 (N_14691,N_11140,N_11473);
nor U14692 (N_14692,N_9638,N_10400);
xor U14693 (N_14693,N_11515,N_10792);
and U14694 (N_14694,N_10051,N_11790);
nor U14695 (N_14695,N_11816,N_9649);
xnor U14696 (N_14696,N_11638,N_10405);
nor U14697 (N_14697,N_12294,N_9503);
nor U14698 (N_14698,N_9760,N_9603);
nor U14699 (N_14699,N_11558,N_11579);
nand U14700 (N_14700,N_9431,N_10822);
or U14701 (N_14701,N_10228,N_12038);
or U14702 (N_14702,N_10736,N_11251);
or U14703 (N_14703,N_10922,N_9452);
and U14704 (N_14704,N_10807,N_12054);
and U14705 (N_14705,N_11130,N_12475);
and U14706 (N_14706,N_12290,N_12480);
nand U14707 (N_14707,N_9472,N_11477);
and U14708 (N_14708,N_11550,N_10822);
nand U14709 (N_14709,N_11248,N_12498);
nor U14710 (N_14710,N_10221,N_10823);
nand U14711 (N_14711,N_12260,N_11956);
nand U14712 (N_14712,N_12160,N_12180);
xnor U14713 (N_14713,N_11517,N_9802);
nor U14714 (N_14714,N_11471,N_11680);
nor U14715 (N_14715,N_12382,N_12467);
nor U14716 (N_14716,N_9988,N_10020);
nor U14717 (N_14717,N_11919,N_9805);
nand U14718 (N_14718,N_12102,N_10415);
and U14719 (N_14719,N_10707,N_12055);
nor U14720 (N_14720,N_9810,N_12326);
nor U14721 (N_14721,N_11529,N_10645);
and U14722 (N_14722,N_12198,N_9569);
or U14723 (N_14723,N_11563,N_11141);
or U14724 (N_14724,N_10255,N_11726);
or U14725 (N_14725,N_11470,N_11832);
nand U14726 (N_14726,N_11726,N_9384);
nor U14727 (N_14727,N_11315,N_10465);
or U14728 (N_14728,N_12364,N_11070);
or U14729 (N_14729,N_11488,N_11269);
nand U14730 (N_14730,N_11913,N_11422);
and U14731 (N_14731,N_12107,N_10072);
nor U14732 (N_14732,N_10794,N_9571);
or U14733 (N_14733,N_9537,N_12170);
or U14734 (N_14734,N_9749,N_12305);
or U14735 (N_14735,N_10633,N_10716);
xnor U14736 (N_14736,N_10788,N_12115);
xnor U14737 (N_14737,N_9997,N_10480);
or U14738 (N_14738,N_11996,N_10312);
nand U14739 (N_14739,N_10232,N_12295);
and U14740 (N_14740,N_12379,N_11343);
nand U14741 (N_14741,N_10186,N_9589);
and U14742 (N_14742,N_11692,N_10104);
and U14743 (N_14743,N_11639,N_11796);
and U14744 (N_14744,N_11018,N_12009);
and U14745 (N_14745,N_11064,N_12045);
or U14746 (N_14746,N_11162,N_11146);
nand U14747 (N_14747,N_10607,N_12485);
nand U14748 (N_14748,N_9929,N_11812);
and U14749 (N_14749,N_11335,N_11755);
nand U14750 (N_14750,N_11709,N_11385);
or U14751 (N_14751,N_10621,N_11092);
nor U14752 (N_14752,N_9887,N_9957);
or U14753 (N_14753,N_12210,N_10988);
or U14754 (N_14754,N_9786,N_11241);
nand U14755 (N_14755,N_11163,N_9447);
or U14756 (N_14756,N_11567,N_9790);
or U14757 (N_14757,N_11246,N_11261);
nand U14758 (N_14758,N_12209,N_11337);
nor U14759 (N_14759,N_12239,N_9509);
and U14760 (N_14760,N_9617,N_9600);
and U14761 (N_14761,N_10147,N_11353);
and U14762 (N_14762,N_10983,N_9643);
or U14763 (N_14763,N_10420,N_11500);
nand U14764 (N_14764,N_10227,N_12074);
xor U14765 (N_14765,N_9787,N_11124);
and U14766 (N_14766,N_9946,N_10647);
xor U14767 (N_14767,N_9694,N_11685);
nand U14768 (N_14768,N_11423,N_10923);
and U14769 (N_14769,N_12499,N_10803);
nor U14770 (N_14770,N_10355,N_12114);
or U14771 (N_14771,N_12296,N_11037);
or U14772 (N_14772,N_10598,N_9781);
nor U14773 (N_14773,N_10370,N_11627);
or U14774 (N_14774,N_10455,N_11425);
nor U14775 (N_14775,N_11874,N_11429);
or U14776 (N_14776,N_10191,N_9850);
or U14777 (N_14777,N_12312,N_11831);
nor U14778 (N_14778,N_11766,N_11266);
and U14779 (N_14779,N_10927,N_11081);
or U14780 (N_14780,N_10141,N_12481);
nand U14781 (N_14781,N_9704,N_12016);
or U14782 (N_14782,N_10016,N_11050);
nand U14783 (N_14783,N_10509,N_10179);
xor U14784 (N_14784,N_10030,N_11352);
xor U14785 (N_14785,N_9635,N_11646);
and U14786 (N_14786,N_10769,N_10126);
or U14787 (N_14787,N_11427,N_11057);
or U14788 (N_14788,N_12075,N_10468);
or U14789 (N_14789,N_9771,N_12373);
and U14790 (N_14790,N_10309,N_10068);
nand U14791 (N_14791,N_9992,N_10048);
or U14792 (N_14792,N_11152,N_11707);
or U14793 (N_14793,N_10677,N_9549);
nand U14794 (N_14794,N_11320,N_11575);
and U14795 (N_14795,N_11140,N_11413);
nand U14796 (N_14796,N_9859,N_10022);
nor U14797 (N_14797,N_11479,N_10981);
nor U14798 (N_14798,N_9505,N_9979);
nand U14799 (N_14799,N_10063,N_11099);
and U14800 (N_14800,N_9436,N_10762);
xor U14801 (N_14801,N_10129,N_12403);
and U14802 (N_14802,N_11017,N_10819);
or U14803 (N_14803,N_9650,N_12200);
xnor U14804 (N_14804,N_9787,N_9650);
and U14805 (N_14805,N_9510,N_10412);
xnor U14806 (N_14806,N_10593,N_9529);
nor U14807 (N_14807,N_10151,N_10595);
nor U14808 (N_14808,N_11405,N_9921);
or U14809 (N_14809,N_12131,N_11370);
or U14810 (N_14810,N_10787,N_9379);
nand U14811 (N_14811,N_10733,N_9420);
or U14812 (N_14812,N_10000,N_11576);
nand U14813 (N_14813,N_11236,N_11059);
and U14814 (N_14814,N_12332,N_10771);
or U14815 (N_14815,N_10018,N_10061);
nor U14816 (N_14816,N_10327,N_9378);
or U14817 (N_14817,N_12035,N_12320);
and U14818 (N_14818,N_9406,N_10571);
and U14819 (N_14819,N_10349,N_10556);
nand U14820 (N_14820,N_12424,N_10645);
xor U14821 (N_14821,N_12342,N_11117);
nor U14822 (N_14822,N_10729,N_10823);
nor U14823 (N_14823,N_12072,N_9962);
and U14824 (N_14824,N_10608,N_9594);
and U14825 (N_14825,N_10073,N_11573);
xor U14826 (N_14826,N_11889,N_9841);
nor U14827 (N_14827,N_12466,N_10629);
and U14828 (N_14828,N_9955,N_11794);
or U14829 (N_14829,N_10757,N_11380);
and U14830 (N_14830,N_10604,N_12202);
nor U14831 (N_14831,N_10577,N_9601);
and U14832 (N_14832,N_12240,N_12115);
nand U14833 (N_14833,N_9927,N_9699);
xor U14834 (N_14834,N_11157,N_12097);
or U14835 (N_14835,N_10638,N_10106);
nor U14836 (N_14836,N_12367,N_11960);
nor U14837 (N_14837,N_12263,N_11708);
and U14838 (N_14838,N_10580,N_11826);
nand U14839 (N_14839,N_9436,N_10178);
nor U14840 (N_14840,N_10178,N_10302);
nand U14841 (N_14841,N_11266,N_11900);
or U14842 (N_14842,N_9484,N_9834);
nor U14843 (N_14843,N_9455,N_10729);
nor U14844 (N_14844,N_11215,N_11563);
nand U14845 (N_14845,N_10677,N_11286);
xnor U14846 (N_14846,N_11935,N_9650);
nand U14847 (N_14847,N_10245,N_9806);
nand U14848 (N_14848,N_10368,N_12310);
nor U14849 (N_14849,N_10942,N_12105);
or U14850 (N_14850,N_10883,N_10185);
nor U14851 (N_14851,N_12147,N_11240);
or U14852 (N_14852,N_11873,N_11821);
or U14853 (N_14853,N_10479,N_10942);
nand U14854 (N_14854,N_10922,N_10784);
or U14855 (N_14855,N_11617,N_9513);
or U14856 (N_14856,N_10022,N_9502);
nand U14857 (N_14857,N_10269,N_9512);
nand U14858 (N_14858,N_11759,N_12389);
nand U14859 (N_14859,N_12035,N_11821);
nand U14860 (N_14860,N_12373,N_9424);
xor U14861 (N_14861,N_9854,N_10208);
and U14862 (N_14862,N_9967,N_9959);
nor U14863 (N_14863,N_11305,N_9753);
xnor U14864 (N_14864,N_9721,N_10154);
and U14865 (N_14865,N_11350,N_9379);
nor U14866 (N_14866,N_10493,N_11115);
nand U14867 (N_14867,N_11764,N_11627);
and U14868 (N_14868,N_9872,N_11990);
nand U14869 (N_14869,N_11877,N_11345);
nor U14870 (N_14870,N_11741,N_9817);
nor U14871 (N_14871,N_9856,N_11373);
nand U14872 (N_14872,N_10259,N_11435);
nor U14873 (N_14873,N_10047,N_10976);
or U14874 (N_14874,N_10396,N_12164);
or U14875 (N_14875,N_11358,N_10094);
or U14876 (N_14876,N_9944,N_9738);
nand U14877 (N_14877,N_10604,N_11027);
nor U14878 (N_14878,N_11582,N_10229);
and U14879 (N_14879,N_12462,N_10295);
or U14880 (N_14880,N_10113,N_11037);
and U14881 (N_14881,N_11586,N_10711);
nand U14882 (N_14882,N_12347,N_11632);
or U14883 (N_14883,N_11431,N_11787);
or U14884 (N_14884,N_12026,N_11201);
and U14885 (N_14885,N_11197,N_9800);
nand U14886 (N_14886,N_10318,N_10201);
nor U14887 (N_14887,N_12227,N_11711);
nor U14888 (N_14888,N_10376,N_10937);
or U14889 (N_14889,N_10554,N_12047);
or U14890 (N_14890,N_11664,N_9628);
nor U14891 (N_14891,N_10699,N_12001);
nand U14892 (N_14892,N_9737,N_11042);
and U14893 (N_14893,N_11808,N_10203);
and U14894 (N_14894,N_9541,N_10254);
and U14895 (N_14895,N_9751,N_9762);
nor U14896 (N_14896,N_11175,N_11827);
nand U14897 (N_14897,N_10283,N_12335);
nand U14898 (N_14898,N_10460,N_9732);
xor U14899 (N_14899,N_11238,N_9630);
and U14900 (N_14900,N_9577,N_11806);
nand U14901 (N_14901,N_11822,N_10833);
nand U14902 (N_14902,N_9690,N_10787);
or U14903 (N_14903,N_12475,N_12193);
xor U14904 (N_14904,N_10919,N_11514);
nand U14905 (N_14905,N_9380,N_9552);
or U14906 (N_14906,N_9640,N_10881);
nor U14907 (N_14907,N_11759,N_11110);
nor U14908 (N_14908,N_11089,N_11548);
and U14909 (N_14909,N_12131,N_10024);
nand U14910 (N_14910,N_10026,N_10861);
and U14911 (N_14911,N_11520,N_11887);
nand U14912 (N_14912,N_11062,N_10185);
nand U14913 (N_14913,N_11633,N_11263);
nand U14914 (N_14914,N_12419,N_10865);
nor U14915 (N_14915,N_10478,N_10440);
nand U14916 (N_14916,N_9544,N_10559);
or U14917 (N_14917,N_12485,N_9921);
nand U14918 (N_14918,N_11791,N_11743);
nor U14919 (N_14919,N_10633,N_10432);
or U14920 (N_14920,N_12053,N_10147);
and U14921 (N_14921,N_10477,N_10541);
or U14922 (N_14922,N_11656,N_9684);
nand U14923 (N_14923,N_9439,N_10876);
or U14924 (N_14924,N_11562,N_11215);
and U14925 (N_14925,N_10924,N_10101);
or U14926 (N_14926,N_9494,N_11993);
xor U14927 (N_14927,N_10540,N_10680);
and U14928 (N_14928,N_9668,N_11466);
nand U14929 (N_14929,N_9830,N_9376);
and U14930 (N_14930,N_9480,N_11027);
nand U14931 (N_14931,N_10453,N_10695);
or U14932 (N_14932,N_10472,N_11801);
or U14933 (N_14933,N_11463,N_10433);
nor U14934 (N_14934,N_10544,N_12467);
and U14935 (N_14935,N_9592,N_9583);
nor U14936 (N_14936,N_9466,N_10953);
or U14937 (N_14937,N_11012,N_9431);
and U14938 (N_14938,N_12016,N_11628);
nor U14939 (N_14939,N_11048,N_10391);
nand U14940 (N_14940,N_11394,N_12025);
or U14941 (N_14941,N_11640,N_9621);
and U14942 (N_14942,N_11259,N_11858);
xor U14943 (N_14943,N_10800,N_11055);
xnor U14944 (N_14944,N_10894,N_11939);
nand U14945 (N_14945,N_9521,N_11050);
nor U14946 (N_14946,N_11101,N_11726);
nor U14947 (N_14947,N_11166,N_11531);
xor U14948 (N_14948,N_12046,N_10180);
or U14949 (N_14949,N_10024,N_9927);
nor U14950 (N_14950,N_12161,N_11003);
nand U14951 (N_14951,N_10631,N_11305);
and U14952 (N_14952,N_11034,N_10620);
nor U14953 (N_14953,N_12071,N_11922);
nor U14954 (N_14954,N_9793,N_11868);
nor U14955 (N_14955,N_11142,N_12220);
xnor U14956 (N_14956,N_10492,N_10677);
xnor U14957 (N_14957,N_10474,N_10081);
or U14958 (N_14958,N_9670,N_12282);
or U14959 (N_14959,N_9702,N_11199);
and U14960 (N_14960,N_9447,N_9409);
xor U14961 (N_14961,N_12005,N_11628);
nand U14962 (N_14962,N_9424,N_11730);
and U14963 (N_14963,N_9618,N_10743);
and U14964 (N_14964,N_12342,N_12053);
or U14965 (N_14965,N_9440,N_11212);
nor U14966 (N_14966,N_9601,N_12281);
xnor U14967 (N_14967,N_10600,N_10151);
and U14968 (N_14968,N_11979,N_9408);
and U14969 (N_14969,N_12085,N_12323);
nand U14970 (N_14970,N_10777,N_11414);
and U14971 (N_14971,N_11358,N_12009);
nor U14972 (N_14972,N_11080,N_9806);
nand U14973 (N_14973,N_10298,N_9825);
nor U14974 (N_14974,N_11523,N_12035);
and U14975 (N_14975,N_11217,N_9664);
nor U14976 (N_14976,N_9911,N_9482);
nand U14977 (N_14977,N_9481,N_9850);
nand U14978 (N_14978,N_11558,N_11266);
nand U14979 (N_14979,N_11210,N_11836);
nand U14980 (N_14980,N_10225,N_9895);
nand U14981 (N_14981,N_11151,N_10640);
and U14982 (N_14982,N_10010,N_12359);
or U14983 (N_14983,N_9697,N_9416);
and U14984 (N_14984,N_11815,N_10110);
or U14985 (N_14985,N_10930,N_11789);
nand U14986 (N_14986,N_9406,N_11853);
nand U14987 (N_14987,N_11636,N_10970);
and U14988 (N_14988,N_12473,N_11320);
nand U14989 (N_14989,N_9449,N_11804);
or U14990 (N_14990,N_10030,N_11211);
nand U14991 (N_14991,N_10530,N_11377);
nor U14992 (N_14992,N_9941,N_10700);
nor U14993 (N_14993,N_10190,N_11769);
and U14994 (N_14994,N_12162,N_10084);
nand U14995 (N_14995,N_12037,N_9914);
and U14996 (N_14996,N_10990,N_12405);
xor U14997 (N_14997,N_11201,N_10398);
nand U14998 (N_14998,N_12032,N_9529);
and U14999 (N_14999,N_11220,N_9757);
or U15000 (N_15000,N_10176,N_12218);
or U15001 (N_15001,N_11255,N_11589);
and U15002 (N_15002,N_10344,N_11663);
xnor U15003 (N_15003,N_10413,N_12455);
or U15004 (N_15004,N_12149,N_9867);
nand U15005 (N_15005,N_10195,N_10436);
or U15006 (N_15006,N_11857,N_10114);
and U15007 (N_15007,N_11952,N_11175);
nor U15008 (N_15008,N_9403,N_10646);
and U15009 (N_15009,N_10256,N_12042);
nor U15010 (N_15010,N_10911,N_11583);
or U15011 (N_15011,N_11475,N_11674);
or U15012 (N_15012,N_9950,N_10036);
and U15013 (N_15013,N_11470,N_10362);
nand U15014 (N_15014,N_11905,N_9739);
nor U15015 (N_15015,N_9953,N_9485);
and U15016 (N_15016,N_12263,N_11562);
nor U15017 (N_15017,N_11676,N_10533);
and U15018 (N_15018,N_11280,N_12183);
or U15019 (N_15019,N_11837,N_9592);
nand U15020 (N_15020,N_11740,N_10213);
and U15021 (N_15021,N_9419,N_12184);
xnor U15022 (N_15022,N_11167,N_11888);
nor U15023 (N_15023,N_11930,N_11185);
and U15024 (N_15024,N_10234,N_9812);
and U15025 (N_15025,N_10962,N_9684);
and U15026 (N_15026,N_10438,N_10147);
and U15027 (N_15027,N_10725,N_11192);
nor U15028 (N_15028,N_9736,N_12138);
or U15029 (N_15029,N_10061,N_11503);
and U15030 (N_15030,N_10984,N_9664);
or U15031 (N_15031,N_11396,N_11240);
nand U15032 (N_15032,N_11863,N_10429);
or U15033 (N_15033,N_9401,N_9551);
and U15034 (N_15034,N_9877,N_11840);
or U15035 (N_15035,N_10766,N_11406);
and U15036 (N_15036,N_11996,N_10903);
nor U15037 (N_15037,N_11053,N_10886);
or U15038 (N_15038,N_9924,N_11900);
and U15039 (N_15039,N_11884,N_11295);
nor U15040 (N_15040,N_10165,N_11868);
xor U15041 (N_15041,N_10728,N_9815);
xnor U15042 (N_15042,N_12280,N_12299);
xor U15043 (N_15043,N_9690,N_11967);
nand U15044 (N_15044,N_11339,N_10590);
or U15045 (N_15045,N_11926,N_10202);
or U15046 (N_15046,N_12220,N_9791);
or U15047 (N_15047,N_10869,N_10632);
nor U15048 (N_15048,N_12389,N_10488);
and U15049 (N_15049,N_11971,N_10684);
nand U15050 (N_15050,N_12288,N_11919);
nand U15051 (N_15051,N_10759,N_9948);
and U15052 (N_15052,N_11426,N_10888);
xor U15053 (N_15053,N_10278,N_11542);
nand U15054 (N_15054,N_11893,N_10425);
nand U15055 (N_15055,N_11996,N_9459);
nor U15056 (N_15056,N_9399,N_11901);
nand U15057 (N_15057,N_10763,N_10826);
or U15058 (N_15058,N_11816,N_10869);
nand U15059 (N_15059,N_10119,N_11205);
or U15060 (N_15060,N_10119,N_12388);
nand U15061 (N_15061,N_9505,N_12274);
or U15062 (N_15062,N_12314,N_12306);
nor U15063 (N_15063,N_9627,N_10086);
xor U15064 (N_15064,N_9645,N_12355);
or U15065 (N_15065,N_11517,N_11903);
and U15066 (N_15066,N_9391,N_11617);
and U15067 (N_15067,N_10898,N_9643);
or U15068 (N_15068,N_12270,N_12370);
nor U15069 (N_15069,N_9470,N_11603);
nor U15070 (N_15070,N_11505,N_11367);
nor U15071 (N_15071,N_9451,N_10630);
nand U15072 (N_15072,N_11707,N_9834);
nor U15073 (N_15073,N_11718,N_10289);
nand U15074 (N_15074,N_10526,N_9526);
nor U15075 (N_15075,N_9771,N_10106);
nand U15076 (N_15076,N_11204,N_12140);
xor U15077 (N_15077,N_11332,N_11141);
nor U15078 (N_15078,N_10750,N_11424);
or U15079 (N_15079,N_9768,N_9803);
xnor U15080 (N_15080,N_10801,N_10208);
and U15081 (N_15081,N_12317,N_9399);
and U15082 (N_15082,N_9936,N_10747);
and U15083 (N_15083,N_10479,N_9649);
or U15084 (N_15084,N_10071,N_10755);
or U15085 (N_15085,N_12020,N_10156);
and U15086 (N_15086,N_10573,N_9547);
nand U15087 (N_15087,N_10778,N_10606);
nor U15088 (N_15088,N_9965,N_11103);
nand U15089 (N_15089,N_9532,N_9664);
or U15090 (N_15090,N_9727,N_10168);
nand U15091 (N_15091,N_11507,N_10856);
nor U15092 (N_15092,N_11336,N_11143);
nand U15093 (N_15093,N_11181,N_11927);
or U15094 (N_15094,N_12437,N_9467);
nor U15095 (N_15095,N_10700,N_9510);
nand U15096 (N_15096,N_12490,N_9919);
nor U15097 (N_15097,N_10130,N_12341);
nand U15098 (N_15098,N_10975,N_10674);
or U15099 (N_15099,N_10684,N_10527);
nor U15100 (N_15100,N_12063,N_12455);
and U15101 (N_15101,N_11504,N_10828);
nand U15102 (N_15102,N_11457,N_10898);
nand U15103 (N_15103,N_10687,N_9938);
xnor U15104 (N_15104,N_9985,N_11813);
nor U15105 (N_15105,N_10119,N_10747);
and U15106 (N_15106,N_12335,N_10440);
and U15107 (N_15107,N_9619,N_10801);
nor U15108 (N_15108,N_9732,N_10128);
nor U15109 (N_15109,N_12142,N_10584);
or U15110 (N_15110,N_11719,N_12183);
nor U15111 (N_15111,N_9901,N_10432);
and U15112 (N_15112,N_9812,N_11665);
nor U15113 (N_15113,N_11073,N_11214);
or U15114 (N_15114,N_11138,N_10609);
nand U15115 (N_15115,N_9727,N_9970);
nor U15116 (N_15116,N_12312,N_12092);
or U15117 (N_15117,N_10884,N_12303);
or U15118 (N_15118,N_10494,N_11895);
or U15119 (N_15119,N_10210,N_11454);
or U15120 (N_15120,N_9740,N_10086);
or U15121 (N_15121,N_9463,N_11359);
nand U15122 (N_15122,N_10640,N_9835);
or U15123 (N_15123,N_10900,N_10377);
nor U15124 (N_15124,N_11361,N_10021);
and U15125 (N_15125,N_10708,N_11893);
nand U15126 (N_15126,N_10623,N_10265);
xnor U15127 (N_15127,N_10863,N_10956);
or U15128 (N_15128,N_10483,N_9667);
xnor U15129 (N_15129,N_9890,N_9980);
nor U15130 (N_15130,N_11690,N_11747);
and U15131 (N_15131,N_10991,N_12206);
xor U15132 (N_15132,N_11923,N_10589);
and U15133 (N_15133,N_11203,N_10162);
and U15134 (N_15134,N_11334,N_10184);
nor U15135 (N_15135,N_9720,N_10185);
and U15136 (N_15136,N_9752,N_12406);
and U15137 (N_15137,N_10020,N_10765);
and U15138 (N_15138,N_10703,N_11170);
and U15139 (N_15139,N_9427,N_10724);
nand U15140 (N_15140,N_11612,N_9406);
nor U15141 (N_15141,N_11808,N_11066);
nor U15142 (N_15142,N_9806,N_10140);
or U15143 (N_15143,N_11367,N_9720);
xor U15144 (N_15144,N_12351,N_11751);
or U15145 (N_15145,N_9737,N_10976);
and U15146 (N_15146,N_12101,N_11277);
and U15147 (N_15147,N_12236,N_11277);
xnor U15148 (N_15148,N_10314,N_9916);
or U15149 (N_15149,N_9596,N_11066);
and U15150 (N_15150,N_10480,N_10852);
nand U15151 (N_15151,N_11408,N_11126);
nand U15152 (N_15152,N_11806,N_12307);
or U15153 (N_15153,N_11444,N_11631);
nor U15154 (N_15154,N_12109,N_9458);
and U15155 (N_15155,N_10782,N_12440);
and U15156 (N_15156,N_9585,N_11361);
nor U15157 (N_15157,N_12016,N_11399);
and U15158 (N_15158,N_9834,N_10536);
xor U15159 (N_15159,N_11244,N_10444);
nand U15160 (N_15160,N_12495,N_11403);
nand U15161 (N_15161,N_11436,N_10752);
nor U15162 (N_15162,N_12308,N_10457);
nor U15163 (N_15163,N_11120,N_10687);
nand U15164 (N_15164,N_11424,N_9404);
or U15165 (N_15165,N_9660,N_12065);
nor U15166 (N_15166,N_10858,N_11209);
and U15167 (N_15167,N_12049,N_10009);
nand U15168 (N_15168,N_10190,N_9630);
nand U15169 (N_15169,N_12362,N_10608);
and U15170 (N_15170,N_11007,N_11402);
nand U15171 (N_15171,N_12330,N_11494);
nand U15172 (N_15172,N_9507,N_11863);
and U15173 (N_15173,N_9915,N_9375);
nor U15174 (N_15174,N_9586,N_11917);
and U15175 (N_15175,N_10360,N_10670);
and U15176 (N_15176,N_12479,N_10486);
nor U15177 (N_15177,N_12018,N_11006);
nor U15178 (N_15178,N_11203,N_12354);
and U15179 (N_15179,N_12126,N_9690);
nor U15180 (N_15180,N_12066,N_9881);
and U15181 (N_15181,N_9793,N_10745);
nor U15182 (N_15182,N_11104,N_11791);
nor U15183 (N_15183,N_10420,N_11905);
nand U15184 (N_15184,N_10200,N_10858);
nor U15185 (N_15185,N_11800,N_11143);
nand U15186 (N_15186,N_12213,N_12300);
or U15187 (N_15187,N_10825,N_10190);
nand U15188 (N_15188,N_9909,N_11844);
nand U15189 (N_15189,N_10807,N_9731);
nand U15190 (N_15190,N_10055,N_11780);
nand U15191 (N_15191,N_9843,N_9708);
nand U15192 (N_15192,N_11383,N_9499);
or U15193 (N_15193,N_11843,N_11310);
nand U15194 (N_15194,N_12477,N_9519);
and U15195 (N_15195,N_11433,N_11318);
xnor U15196 (N_15196,N_10883,N_9536);
xor U15197 (N_15197,N_12140,N_11845);
and U15198 (N_15198,N_12195,N_10122);
nor U15199 (N_15199,N_10612,N_9946);
nor U15200 (N_15200,N_10190,N_12412);
and U15201 (N_15201,N_12019,N_9501);
nor U15202 (N_15202,N_12197,N_12386);
nand U15203 (N_15203,N_9871,N_9995);
and U15204 (N_15204,N_10316,N_10215);
or U15205 (N_15205,N_11284,N_12327);
nor U15206 (N_15206,N_9909,N_9823);
or U15207 (N_15207,N_12079,N_10064);
nor U15208 (N_15208,N_11598,N_11470);
nand U15209 (N_15209,N_12048,N_11385);
nor U15210 (N_15210,N_12064,N_12095);
xnor U15211 (N_15211,N_11215,N_9428);
nor U15212 (N_15212,N_10896,N_9484);
nand U15213 (N_15213,N_12080,N_11492);
and U15214 (N_15214,N_10177,N_9567);
or U15215 (N_15215,N_11349,N_10854);
nand U15216 (N_15216,N_11019,N_9389);
nor U15217 (N_15217,N_9988,N_10836);
nor U15218 (N_15218,N_11452,N_12027);
nand U15219 (N_15219,N_10603,N_12030);
or U15220 (N_15220,N_11639,N_10609);
or U15221 (N_15221,N_11399,N_11973);
nor U15222 (N_15222,N_10341,N_11447);
nand U15223 (N_15223,N_10186,N_10168);
or U15224 (N_15224,N_12065,N_9780);
and U15225 (N_15225,N_10259,N_10300);
xor U15226 (N_15226,N_11079,N_10233);
or U15227 (N_15227,N_9481,N_11291);
nand U15228 (N_15228,N_11609,N_11078);
xor U15229 (N_15229,N_10536,N_9710);
nand U15230 (N_15230,N_10100,N_10529);
nor U15231 (N_15231,N_12368,N_9399);
and U15232 (N_15232,N_11514,N_11944);
xnor U15233 (N_15233,N_11183,N_9556);
nand U15234 (N_15234,N_11282,N_11548);
nor U15235 (N_15235,N_11361,N_10445);
and U15236 (N_15236,N_10352,N_11021);
or U15237 (N_15237,N_11070,N_10640);
and U15238 (N_15238,N_10399,N_11406);
and U15239 (N_15239,N_10057,N_9775);
and U15240 (N_15240,N_10386,N_12024);
and U15241 (N_15241,N_10227,N_11575);
or U15242 (N_15242,N_11221,N_10548);
and U15243 (N_15243,N_11968,N_11442);
and U15244 (N_15244,N_10568,N_10029);
or U15245 (N_15245,N_11799,N_9689);
nand U15246 (N_15246,N_9849,N_9486);
xor U15247 (N_15247,N_11645,N_9768);
nor U15248 (N_15248,N_9696,N_12382);
or U15249 (N_15249,N_9741,N_10162);
nor U15250 (N_15250,N_10310,N_10215);
or U15251 (N_15251,N_11111,N_10400);
nand U15252 (N_15252,N_11355,N_10285);
or U15253 (N_15253,N_10573,N_10202);
and U15254 (N_15254,N_11798,N_10004);
nor U15255 (N_15255,N_10877,N_10932);
nand U15256 (N_15256,N_11898,N_9798);
or U15257 (N_15257,N_12148,N_10956);
xor U15258 (N_15258,N_10639,N_11468);
and U15259 (N_15259,N_11383,N_10910);
xor U15260 (N_15260,N_10393,N_9804);
nand U15261 (N_15261,N_10692,N_10518);
and U15262 (N_15262,N_12177,N_9901);
or U15263 (N_15263,N_11091,N_11056);
and U15264 (N_15264,N_11763,N_10218);
nand U15265 (N_15265,N_12053,N_9570);
nand U15266 (N_15266,N_12025,N_10591);
or U15267 (N_15267,N_9662,N_9773);
nand U15268 (N_15268,N_10343,N_11902);
nor U15269 (N_15269,N_9414,N_9458);
xor U15270 (N_15270,N_9627,N_11325);
nand U15271 (N_15271,N_9685,N_10385);
xor U15272 (N_15272,N_12335,N_12006);
or U15273 (N_15273,N_9750,N_11645);
xor U15274 (N_15274,N_10615,N_12037);
nor U15275 (N_15275,N_11956,N_10525);
or U15276 (N_15276,N_9680,N_10569);
nand U15277 (N_15277,N_9907,N_12395);
xnor U15278 (N_15278,N_10777,N_10675);
xor U15279 (N_15279,N_9768,N_10705);
nor U15280 (N_15280,N_12010,N_12138);
nor U15281 (N_15281,N_11231,N_11895);
nand U15282 (N_15282,N_11590,N_10211);
and U15283 (N_15283,N_11331,N_10250);
nor U15284 (N_15284,N_11538,N_10922);
nand U15285 (N_15285,N_11085,N_9938);
and U15286 (N_15286,N_10025,N_10895);
xor U15287 (N_15287,N_11691,N_10645);
and U15288 (N_15288,N_11235,N_11941);
or U15289 (N_15289,N_11072,N_12378);
nand U15290 (N_15290,N_9665,N_10913);
xnor U15291 (N_15291,N_9722,N_10188);
nor U15292 (N_15292,N_11170,N_11932);
and U15293 (N_15293,N_12396,N_9724);
nor U15294 (N_15294,N_9634,N_11598);
or U15295 (N_15295,N_10566,N_9625);
or U15296 (N_15296,N_11165,N_9728);
nor U15297 (N_15297,N_11029,N_9658);
nor U15298 (N_15298,N_11979,N_10467);
or U15299 (N_15299,N_12310,N_10014);
or U15300 (N_15300,N_10040,N_9611);
nor U15301 (N_15301,N_10656,N_9897);
nand U15302 (N_15302,N_9675,N_12061);
nand U15303 (N_15303,N_9961,N_10731);
nand U15304 (N_15304,N_10933,N_10954);
nor U15305 (N_15305,N_10261,N_11772);
or U15306 (N_15306,N_11138,N_11780);
xnor U15307 (N_15307,N_10982,N_9769);
or U15308 (N_15308,N_11860,N_9680);
nor U15309 (N_15309,N_10105,N_12113);
and U15310 (N_15310,N_12362,N_11314);
and U15311 (N_15311,N_10500,N_10191);
nand U15312 (N_15312,N_9674,N_12415);
and U15313 (N_15313,N_9992,N_10914);
nand U15314 (N_15314,N_11916,N_12195);
nor U15315 (N_15315,N_9953,N_9729);
xor U15316 (N_15316,N_9471,N_11401);
nand U15317 (N_15317,N_11283,N_11848);
or U15318 (N_15318,N_12463,N_9860);
xnor U15319 (N_15319,N_9450,N_12263);
or U15320 (N_15320,N_9567,N_9713);
nand U15321 (N_15321,N_11440,N_11533);
nor U15322 (N_15322,N_11666,N_12128);
and U15323 (N_15323,N_9977,N_11675);
and U15324 (N_15324,N_10069,N_11538);
nor U15325 (N_15325,N_10066,N_10914);
nor U15326 (N_15326,N_12258,N_10944);
nor U15327 (N_15327,N_9997,N_10623);
or U15328 (N_15328,N_9381,N_12276);
nor U15329 (N_15329,N_9576,N_12449);
nand U15330 (N_15330,N_9413,N_9761);
nor U15331 (N_15331,N_12043,N_10901);
and U15332 (N_15332,N_9462,N_10414);
nor U15333 (N_15333,N_10498,N_11489);
nand U15334 (N_15334,N_11918,N_9475);
nor U15335 (N_15335,N_11454,N_11483);
xor U15336 (N_15336,N_9471,N_9729);
or U15337 (N_15337,N_10065,N_12223);
or U15338 (N_15338,N_11521,N_9803);
nand U15339 (N_15339,N_9676,N_10637);
xnor U15340 (N_15340,N_11370,N_11561);
xor U15341 (N_15341,N_11092,N_10337);
nand U15342 (N_15342,N_9683,N_9667);
nor U15343 (N_15343,N_10880,N_10867);
nor U15344 (N_15344,N_10651,N_12279);
nand U15345 (N_15345,N_10411,N_10961);
and U15346 (N_15346,N_12334,N_10602);
nand U15347 (N_15347,N_10743,N_12485);
xnor U15348 (N_15348,N_10657,N_10216);
nor U15349 (N_15349,N_9549,N_12400);
or U15350 (N_15350,N_11084,N_9692);
and U15351 (N_15351,N_10627,N_11165);
and U15352 (N_15352,N_11839,N_11167);
nand U15353 (N_15353,N_11943,N_9636);
xor U15354 (N_15354,N_9724,N_12063);
and U15355 (N_15355,N_9975,N_12178);
nor U15356 (N_15356,N_10677,N_11617);
or U15357 (N_15357,N_12275,N_12357);
nand U15358 (N_15358,N_12001,N_11776);
and U15359 (N_15359,N_9431,N_10147);
nor U15360 (N_15360,N_11517,N_10187);
or U15361 (N_15361,N_11009,N_9824);
and U15362 (N_15362,N_9470,N_12152);
nor U15363 (N_15363,N_11104,N_12422);
or U15364 (N_15364,N_10063,N_9572);
and U15365 (N_15365,N_11996,N_10519);
or U15366 (N_15366,N_11268,N_9846);
nand U15367 (N_15367,N_10384,N_10706);
nand U15368 (N_15368,N_10737,N_10558);
nand U15369 (N_15369,N_10905,N_10832);
xor U15370 (N_15370,N_9743,N_12398);
nand U15371 (N_15371,N_9903,N_9710);
nor U15372 (N_15372,N_12462,N_10346);
nor U15373 (N_15373,N_10477,N_9460);
nand U15374 (N_15374,N_10746,N_10391);
and U15375 (N_15375,N_11217,N_10014);
xor U15376 (N_15376,N_12294,N_12192);
and U15377 (N_15377,N_10005,N_9550);
or U15378 (N_15378,N_10460,N_11575);
nand U15379 (N_15379,N_9589,N_10684);
and U15380 (N_15380,N_9916,N_9860);
or U15381 (N_15381,N_11948,N_12173);
nand U15382 (N_15382,N_10576,N_9507);
or U15383 (N_15383,N_11372,N_10359);
and U15384 (N_15384,N_9510,N_12238);
and U15385 (N_15385,N_11062,N_12126);
or U15386 (N_15386,N_11735,N_10046);
or U15387 (N_15387,N_10584,N_11041);
nand U15388 (N_15388,N_9644,N_10020);
nor U15389 (N_15389,N_11703,N_9673);
or U15390 (N_15390,N_11490,N_9554);
nor U15391 (N_15391,N_12234,N_11215);
or U15392 (N_15392,N_12245,N_10067);
and U15393 (N_15393,N_9775,N_11130);
nand U15394 (N_15394,N_12409,N_9642);
or U15395 (N_15395,N_12183,N_10218);
nand U15396 (N_15396,N_12029,N_9947);
or U15397 (N_15397,N_11532,N_9873);
nand U15398 (N_15398,N_12300,N_11867);
nand U15399 (N_15399,N_10229,N_11755);
nand U15400 (N_15400,N_10289,N_9833);
nand U15401 (N_15401,N_11846,N_11914);
or U15402 (N_15402,N_11588,N_11343);
nor U15403 (N_15403,N_11684,N_9847);
or U15404 (N_15404,N_12306,N_11234);
nand U15405 (N_15405,N_10129,N_12350);
nand U15406 (N_15406,N_12400,N_9726);
or U15407 (N_15407,N_10399,N_12411);
xor U15408 (N_15408,N_11248,N_11329);
nand U15409 (N_15409,N_9956,N_9771);
or U15410 (N_15410,N_10712,N_9480);
or U15411 (N_15411,N_12482,N_9691);
nand U15412 (N_15412,N_10268,N_9584);
or U15413 (N_15413,N_10796,N_12145);
nor U15414 (N_15414,N_12010,N_10419);
nand U15415 (N_15415,N_11383,N_9818);
nand U15416 (N_15416,N_10792,N_11927);
nand U15417 (N_15417,N_11203,N_11373);
nand U15418 (N_15418,N_9561,N_11513);
or U15419 (N_15419,N_10268,N_11220);
nor U15420 (N_15420,N_10011,N_10121);
or U15421 (N_15421,N_11304,N_11323);
or U15422 (N_15422,N_11799,N_10233);
nor U15423 (N_15423,N_9753,N_12288);
nand U15424 (N_15424,N_11285,N_11880);
or U15425 (N_15425,N_10715,N_11064);
and U15426 (N_15426,N_10414,N_11672);
nand U15427 (N_15427,N_10186,N_12442);
and U15428 (N_15428,N_12355,N_11461);
or U15429 (N_15429,N_11206,N_11658);
nand U15430 (N_15430,N_11775,N_12278);
or U15431 (N_15431,N_10325,N_12228);
and U15432 (N_15432,N_12441,N_11239);
and U15433 (N_15433,N_10807,N_11483);
and U15434 (N_15434,N_12082,N_9781);
nor U15435 (N_15435,N_11414,N_11422);
nand U15436 (N_15436,N_10327,N_11415);
xor U15437 (N_15437,N_11440,N_9684);
or U15438 (N_15438,N_9631,N_9446);
nor U15439 (N_15439,N_9984,N_12218);
xnor U15440 (N_15440,N_10709,N_9607);
and U15441 (N_15441,N_11429,N_12335);
nand U15442 (N_15442,N_10410,N_12377);
nand U15443 (N_15443,N_12045,N_9386);
nand U15444 (N_15444,N_10617,N_9799);
nor U15445 (N_15445,N_12443,N_10242);
nor U15446 (N_15446,N_12271,N_11241);
nor U15447 (N_15447,N_11157,N_12279);
nor U15448 (N_15448,N_12214,N_12017);
or U15449 (N_15449,N_11776,N_12233);
nand U15450 (N_15450,N_11055,N_10916);
nor U15451 (N_15451,N_12383,N_12461);
nor U15452 (N_15452,N_10735,N_9759);
nor U15453 (N_15453,N_11554,N_9439);
or U15454 (N_15454,N_11048,N_11762);
and U15455 (N_15455,N_12004,N_11421);
nand U15456 (N_15456,N_10680,N_10500);
nand U15457 (N_15457,N_9801,N_11452);
xnor U15458 (N_15458,N_12041,N_10459);
nor U15459 (N_15459,N_9915,N_11569);
nand U15460 (N_15460,N_11317,N_10883);
xor U15461 (N_15461,N_10923,N_12090);
nor U15462 (N_15462,N_9642,N_11669);
nand U15463 (N_15463,N_9914,N_9933);
xnor U15464 (N_15464,N_10610,N_11371);
or U15465 (N_15465,N_12143,N_12108);
xor U15466 (N_15466,N_10583,N_11333);
and U15467 (N_15467,N_10512,N_11307);
nor U15468 (N_15468,N_10390,N_9577);
nand U15469 (N_15469,N_10438,N_11249);
nand U15470 (N_15470,N_11520,N_9377);
or U15471 (N_15471,N_10924,N_9918);
nand U15472 (N_15472,N_10477,N_11711);
or U15473 (N_15473,N_12189,N_11549);
nand U15474 (N_15474,N_10020,N_10879);
and U15475 (N_15475,N_10584,N_10777);
and U15476 (N_15476,N_9542,N_9642);
or U15477 (N_15477,N_9998,N_11259);
xnor U15478 (N_15478,N_9879,N_9732);
nand U15479 (N_15479,N_10987,N_11100);
nand U15480 (N_15480,N_11689,N_10637);
nand U15481 (N_15481,N_9421,N_9916);
nor U15482 (N_15482,N_9586,N_12024);
nor U15483 (N_15483,N_10518,N_10292);
xor U15484 (N_15484,N_10733,N_12002);
or U15485 (N_15485,N_10144,N_10440);
or U15486 (N_15486,N_11739,N_10978);
nand U15487 (N_15487,N_10506,N_10539);
and U15488 (N_15488,N_12471,N_12217);
or U15489 (N_15489,N_11008,N_12081);
and U15490 (N_15490,N_11974,N_11945);
and U15491 (N_15491,N_10138,N_11549);
and U15492 (N_15492,N_12442,N_9571);
xor U15493 (N_15493,N_11514,N_10913);
and U15494 (N_15494,N_10852,N_10618);
nor U15495 (N_15495,N_9414,N_9987);
nand U15496 (N_15496,N_12287,N_10718);
and U15497 (N_15497,N_12026,N_11299);
and U15498 (N_15498,N_11197,N_9662);
xnor U15499 (N_15499,N_9407,N_9837);
nor U15500 (N_15500,N_12323,N_10060);
and U15501 (N_15501,N_10080,N_11780);
nand U15502 (N_15502,N_12089,N_9663);
xor U15503 (N_15503,N_11123,N_10888);
nand U15504 (N_15504,N_9901,N_10338);
and U15505 (N_15505,N_10940,N_11421);
nor U15506 (N_15506,N_9831,N_10907);
nor U15507 (N_15507,N_11822,N_10838);
nor U15508 (N_15508,N_12194,N_11194);
nand U15509 (N_15509,N_11931,N_11855);
xor U15510 (N_15510,N_10002,N_11235);
nor U15511 (N_15511,N_9565,N_9471);
or U15512 (N_15512,N_9492,N_11567);
or U15513 (N_15513,N_10904,N_10541);
nand U15514 (N_15514,N_10190,N_10073);
or U15515 (N_15515,N_11166,N_10832);
nor U15516 (N_15516,N_10931,N_10537);
nor U15517 (N_15517,N_10359,N_11909);
and U15518 (N_15518,N_9865,N_11834);
nor U15519 (N_15519,N_10701,N_10240);
or U15520 (N_15520,N_11610,N_10051);
nor U15521 (N_15521,N_11675,N_9693);
nand U15522 (N_15522,N_10132,N_9890);
or U15523 (N_15523,N_10520,N_11994);
or U15524 (N_15524,N_10858,N_12465);
or U15525 (N_15525,N_10864,N_12404);
nor U15526 (N_15526,N_10815,N_10262);
or U15527 (N_15527,N_10803,N_10496);
nand U15528 (N_15528,N_12350,N_10418);
and U15529 (N_15529,N_12315,N_12425);
and U15530 (N_15530,N_10126,N_11999);
nor U15531 (N_15531,N_11156,N_9606);
xor U15532 (N_15532,N_12214,N_11816);
and U15533 (N_15533,N_12067,N_10897);
or U15534 (N_15534,N_12041,N_11469);
or U15535 (N_15535,N_9871,N_10501);
or U15536 (N_15536,N_11521,N_12233);
and U15537 (N_15537,N_9468,N_12400);
nor U15538 (N_15538,N_12454,N_10087);
nor U15539 (N_15539,N_11418,N_10561);
nor U15540 (N_15540,N_10474,N_10773);
or U15541 (N_15541,N_10515,N_11700);
nor U15542 (N_15542,N_11787,N_9810);
and U15543 (N_15543,N_9799,N_12238);
nor U15544 (N_15544,N_11675,N_10344);
xnor U15545 (N_15545,N_11293,N_9795);
and U15546 (N_15546,N_11429,N_10961);
xor U15547 (N_15547,N_11745,N_10731);
or U15548 (N_15548,N_9461,N_9996);
and U15549 (N_15549,N_12431,N_10453);
or U15550 (N_15550,N_11578,N_9884);
nor U15551 (N_15551,N_10197,N_10572);
xnor U15552 (N_15552,N_11786,N_9840);
nand U15553 (N_15553,N_12413,N_10435);
or U15554 (N_15554,N_11037,N_12293);
nor U15555 (N_15555,N_10975,N_11485);
nand U15556 (N_15556,N_9906,N_12439);
or U15557 (N_15557,N_11358,N_11584);
and U15558 (N_15558,N_11138,N_11816);
nor U15559 (N_15559,N_12412,N_11270);
or U15560 (N_15560,N_12281,N_10624);
nor U15561 (N_15561,N_10209,N_10526);
nor U15562 (N_15562,N_11780,N_9845);
nand U15563 (N_15563,N_9437,N_10440);
xnor U15564 (N_15564,N_10570,N_11541);
and U15565 (N_15565,N_10655,N_10351);
or U15566 (N_15566,N_10747,N_9889);
nor U15567 (N_15567,N_12135,N_12168);
and U15568 (N_15568,N_11330,N_10150);
nor U15569 (N_15569,N_11401,N_11869);
and U15570 (N_15570,N_11725,N_9869);
nor U15571 (N_15571,N_10530,N_10533);
or U15572 (N_15572,N_10950,N_10436);
nor U15573 (N_15573,N_10691,N_11399);
and U15574 (N_15574,N_12148,N_10798);
xor U15575 (N_15575,N_11461,N_10968);
nand U15576 (N_15576,N_9621,N_12418);
and U15577 (N_15577,N_10017,N_9968);
or U15578 (N_15578,N_10793,N_9766);
nor U15579 (N_15579,N_9838,N_10097);
and U15580 (N_15580,N_12403,N_12365);
or U15581 (N_15581,N_9424,N_11689);
and U15582 (N_15582,N_11909,N_9605);
or U15583 (N_15583,N_11962,N_12428);
xor U15584 (N_15584,N_10991,N_10059);
nand U15585 (N_15585,N_9962,N_12441);
or U15586 (N_15586,N_10101,N_9934);
or U15587 (N_15587,N_10344,N_11244);
and U15588 (N_15588,N_12242,N_9568);
xor U15589 (N_15589,N_10935,N_10887);
nor U15590 (N_15590,N_10966,N_11681);
nand U15591 (N_15591,N_11328,N_9483);
nand U15592 (N_15592,N_12449,N_12484);
and U15593 (N_15593,N_11861,N_9621);
nor U15594 (N_15594,N_11826,N_11100);
and U15595 (N_15595,N_11231,N_10625);
and U15596 (N_15596,N_10473,N_10557);
and U15597 (N_15597,N_11245,N_9543);
nand U15598 (N_15598,N_12281,N_9848);
nand U15599 (N_15599,N_11393,N_11997);
and U15600 (N_15600,N_9916,N_10708);
and U15601 (N_15601,N_11943,N_9440);
nor U15602 (N_15602,N_10125,N_10198);
and U15603 (N_15603,N_11471,N_10799);
nor U15604 (N_15604,N_9489,N_11285);
nand U15605 (N_15605,N_11215,N_10445);
or U15606 (N_15606,N_10205,N_12458);
nand U15607 (N_15607,N_10227,N_12179);
or U15608 (N_15608,N_9522,N_9786);
nand U15609 (N_15609,N_11119,N_10237);
nand U15610 (N_15610,N_10379,N_10167);
nand U15611 (N_15611,N_9982,N_11943);
nand U15612 (N_15612,N_9831,N_10296);
and U15613 (N_15613,N_11766,N_12032);
or U15614 (N_15614,N_12127,N_11491);
or U15615 (N_15615,N_9566,N_12219);
nand U15616 (N_15616,N_10824,N_11091);
nor U15617 (N_15617,N_9503,N_10681);
nand U15618 (N_15618,N_11521,N_11973);
or U15619 (N_15619,N_10636,N_10945);
and U15620 (N_15620,N_9727,N_11949);
and U15621 (N_15621,N_11561,N_9526);
nand U15622 (N_15622,N_10720,N_12280);
and U15623 (N_15623,N_12052,N_11270);
nor U15624 (N_15624,N_10725,N_12490);
nor U15625 (N_15625,N_13045,N_14989);
and U15626 (N_15626,N_13617,N_14920);
nand U15627 (N_15627,N_14395,N_13179);
nand U15628 (N_15628,N_12625,N_14518);
nand U15629 (N_15629,N_13297,N_15173);
or U15630 (N_15630,N_13715,N_12973);
and U15631 (N_15631,N_14414,N_13275);
and U15632 (N_15632,N_13340,N_15584);
or U15633 (N_15633,N_13492,N_14440);
or U15634 (N_15634,N_12514,N_14788);
nor U15635 (N_15635,N_15414,N_14619);
or U15636 (N_15636,N_15140,N_12700);
or U15637 (N_15637,N_14351,N_15486);
xnor U15638 (N_15638,N_15258,N_14429);
and U15639 (N_15639,N_14531,N_14138);
nand U15640 (N_15640,N_14391,N_14460);
nor U15641 (N_15641,N_13674,N_14940);
xnor U15642 (N_15642,N_12989,N_15399);
or U15643 (N_15643,N_14929,N_15532);
or U15644 (N_15644,N_14037,N_13050);
xor U15645 (N_15645,N_12770,N_12596);
nand U15646 (N_15646,N_12569,N_14262);
and U15647 (N_15647,N_13768,N_13676);
nor U15648 (N_15648,N_15282,N_15426);
nand U15649 (N_15649,N_13299,N_15189);
xor U15650 (N_15650,N_14828,N_12898);
or U15651 (N_15651,N_14645,N_13111);
or U15652 (N_15652,N_13413,N_13270);
xor U15653 (N_15653,N_14729,N_13563);
or U15654 (N_15654,N_15116,N_13473);
and U15655 (N_15655,N_15395,N_15440);
nand U15656 (N_15656,N_13288,N_14546);
nor U15657 (N_15657,N_12693,N_12997);
and U15658 (N_15658,N_15385,N_14325);
or U15659 (N_15659,N_14789,N_13843);
nand U15660 (N_15660,N_13550,N_14353);
nor U15661 (N_15661,N_12921,N_12577);
nor U15662 (N_15662,N_13228,N_12870);
and U15663 (N_15663,N_15576,N_14100);
nand U15664 (N_15664,N_14694,N_14346);
or U15665 (N_15665,N_13744,N_14995);
or U15666 (N_15666,N_14404,N_14715);
xor U15667 (N_15667,N_15005,N_14664);
or U15668 (N_15668,N_12803,N_14448);
nor U15669 (N_15669,N_13580,N_14219);
nor U15670 (N_15670,N_12623,N_12772);
nand U15671 (N_15671,N_12923,N_14135);
nand U15672 (N_15672,N_13221,N_15245);
or U15673 (N_15673,N_12946,N_12594);
nand U15674 (N_15674,N_14466,N_12834);
nor U15675 (N_15675,N_14807,N_13669);
nand U15676 (N_15676,N_13528,N_13258);
nor U15677 (N_15677,N_15289,N_15138);
nand U15678 (N_15678,N_13975,N_15037);
or U15679 (N_15679,N_14381,N_12971);
and U15680 (N_15680,N_14710,N_14363);
nand U15681 (N_15681,N_13914,N_13578);
and U15682 (N_15682,N_14109,N_14380);
xnor U15683 (N_15683,N_13173,N_13274);
and U15684 (N_15684,N_14957,N_12882);
xnor U15685 (N_15685,N_12788,N_15531);
nor U15686 (N_15686,N_13495,N_15236);
nor U15687 (N_15687,N_13039,N_15230);
nand U15688 (N_15688,N_14134,N_13398);
xnor U15689 (N_15689,N_15066,N_12779);
and U15690 (N_15690,N_13420,N_13241);
and U15691 (N_15691,N_15203,N_13476);
and U15692 (N_15692,N_13349,N_14055);
nor U15693 (N_15693,N_12793,N_13396);
nor U15694 (N_15694,N_15192,N_15604);
nor U15695 (N_15695,N_12512,N_13763);
nor U15696 (N_15696,N_13936,N_13403);
xor U15697 (N_15697,N_14066,N_15535);
nor U15698 (N_15698,N_15057,N_15432);
xor U15699 (N_15699,N_15571,N_14476);
nand U15700 (N_15700,N_12888,N_14865);
and U15701 (N_15701,N_14804,N_13874);
nor U15702 (N_15702,N_14961,N_14969);
and U15703 (N_15703,N_15483,N_15216);
nor U15704 (N_15704,N_15158,N_13280);
or U15705 (N_15705,N_14912,N_13102);
nor U15706 (N_15706,N_14427,N_12697);
nand U15707 (N_15707,N_13816,N_14901);
or U15708 (N_15708,N_12904,N_13229);
and U15709 (N_15709,N_14772,N_13348);
nor U15710 (N_15710,N_14170,N_15614);
nand U15711 (N_15711,N_12631,N_14663);
nor U15712 (N_15712,N_15046,N_14107);
nand U15713 (N_15713,N_12566,N_15335);
or U15714 (N_15714,N_15132,N_12843);
and U15715 (N_15715,N_14647,N_14375);
nand U15716 (N_15716,N_12502,N_13222);
nand U15717 (N_15717,N_15585,N_13155);
or U15718 (N_15718,N_15315,N_13732);
and U15719 (N_15719,N_14399,N_15525);
and U15720 (N_15720,N_15554,N_14354);
nor U15721 (N_15721,N_12580,N_12727);
and U15722 (N_15722,N_14153,N_14332);
nor U15723 (N_15723,N_13485,N_12523);
xnor U15724 (N_15724,N_14626,N_14913);
nand U15725 (N_15725,N_13205,N_14463);
nand U15726 (N_15726,N_12829,N_14622);
and U15727 (N_15727,N_13860,N_13959);
or U15728 (N_15728,N_13519,N_14874);
and U15729 (N_15729,N_13167,N_13516);
xor U15730 (N_15730,N_13211,N_13067);
or U15731 (N_15731,N_12524,N_14348);
and U15732 (N_15732,N_15229,N_12785);
nand U15733 (N_15733,N_14509,N_12984);
xnor U15734 (N_15734,N_15000,N_14556);
or U15735 (N_15735,N_15179,N_13367);
or U15736 (N_15736,N_14437,N_13592);
nor U15737 (N_15737,N_14295,N_15023);
nand U15738 (N_15738,N_15187,N_13264);
nand U15739 (N_15739,N_15354,N_14385);
nor U15740 (N_15740,N_13298,N_12783);
and U15741 (N_15741,N_12953,N_14403);
xor U15742 (N_15742,N_13951,N_13438);
and U15743 (N_15743,N_13699,N_13074);
and U15744 (N_15744,N_13197,N_13265);
xor U15745 (N_15745,N_13670,N_15266);
nand U15746 (N_15746,N_13786,N_14606);
or U15747 (N_15747,N_13242,N_14759);
or U15748 (N_15748,N_12696,N_13933);
nand U15749 (N_15749,N_12741,N_15361);
or U15750 (N_15750,N_13190,N_13220);
or U15751 (N_15751,N_14272,N_13481);
and U15752 (N_15752,N_15445,N_12646);
or U15753 (N_15753,N_12748,N_13741);
nor U15754 (N_15754,N_13375,N_14058);
nand U15755 (N_15755,N_12603,N_14624);
and U15756 (N_15756,N_12585,N_13341);
xnor U15757 (N_15757,N_13463,N_12551);
or U15758 (N_15758,N_15468,N_12660);
nor U15759 (N_15759,N_13455,N_14895);
xnor U15760 (N_15760,N_15590,N_14733);
nand U15761 (N_15761,N_15367,N_13870);
and U15762 (N_15762,N_14162,N_14205);
xor U15763 (N_15763,N_14330,N_12819);
nor U15764 (N_15764,N_13273,N_15154);
xnor U15765 (N_15765,N_15123,N_14255);
nand U15766 (N_15766,N_13177,N_13238);
nand U15767 (N_15767,N_14934,N_13588);
nor U15768 (N_15768,N_14638,N_13657);
xor U15769 (N_15769,N_15301,N_13480);
xor U15770 (N_15770,N_12977,N_14666);
and U15771 (N_15771,N_14061,N_13129);
xor U15772 (N_15772,N_13650,N_15155);
and U15773 (N_15773,N_13654,N_14453);
nor U15774 (N_15774,N_13140,N_12600);
nor U15775 (N_15775,N_12992,N_13754);
nand U15776 (N_15776,N_12722,N_12543);
and U15777 (N_15777,N_13200,N_14569);
nor U15778 (N_15778,N_13047,N_13098);
or U15779 (N_15779,N_15586,N_12507);
or U15780 (N_15780,N_15613,N_13802);
or U15781 (N_15781,N_12568,N_14358);
nor U15782 (N_15782,N_15074,N_13989);
nor U15783 (N_15783,N_13240,N_14001);
xor U15784 (N_15784,N_13753,N_15064);
or U15785 (N_15785,N_15600,N_15522);
nand U15786 (N_15786,N_13643,N_14616);
or U15787 (N_15787,N_14840,N_14247);
nor U15788 (N_15788,N_12664,N_15540);
nand U15789 (N_15789,N_14266,N_15444);
and U15790 (N_15790,N_14852,N_14470);
and U15791 (N_15791,N_14250,N_13004);
nand U15792 (N_15792,N_12915,N_12941);
and U15793 (N_15793,N_15506,N_13862);
nor U15794 (N_15794,N_13712,N_14716);
and U15795 (N_15795,N_14725,N_13922);
and U15796 (N_15796,N_13479,N_14667);
and U15797 (N_15797,N_13976,N_15561);
and U15798 (N_15798,N_15325,N_15006);
nor U15799 (N_15799,N_14323,N_13154);
nand U15800 (N_15800,N_13210,N_13764);
nand U15801 (N_15801,N_13419,N_12517);
or U15802 (N_15802,N_13044,N_13108);
and U15803 (N_15803,N_14273,N_14079);
and U15804 (N_15804,N_12613,N_14415);
or U15805 (N_15805,N_14233,N_13306);
nor U15806 (N_15806,N_14514,N_13257);
xnor U15807 (N_15807,N_14076,N_14141);
and U15808 (N_15808,N_13705,N_14821);
nand U15809 (N_15809,N_12736,N_14500);
xor U15810 (N_15810,N_15172,N_13981);
nor U15811 (N_15811,N_14782,N_13491);
nor U15812 (N_15812,N_13424,N_15151);
or U15813 (N_15813,N_13621,N_14342);
nor U15814 (N_15814,N_14428,N_15547);
nand U15815 (N_15815,N_15371,N_15208);
nand U15816 (N_15816,N_15602,N_14411);
and U15817 (N_15817,N_15277,N_14712);
nand U15818 (N_15818,N_13460,N_12970);
and U15819 (N_15819,N_15303,N_13377);
nor U15820 (N_15820,N_12542,N_15487);
nor U15821 (N_15821,N_12976,N_13692);
and U15822 (N_15822,N_15152,N_15213);
and U15823 (N_15823,N_13902,N_15254);
nand U15824 (N_15824,N_14580,N_12728);
nand U15825 (N_15825,N_13005,N_14423);
nand U15826 (N_15826,N_13149,N_13958);
nand U15827 (N_15827,N_13189,N_15346);
or U15828 (N_15828,N_14090,N_14767);
and U15829 (N_15829,N_15275,N_12546);
and U15830 (N_15830,N_14560,N_14537);
and U15831 (N_15831,N_12821,N_14595);
nand U15832 (N_15832,N_13466,N_14340);
and U15833 (N_15833,N_13170,N_13648);
and U15834 (N_15834,N_14454,N_12545);
and U15835 (N_15835,N_15523,N_12581);
and U15836 (N_15836,N_13890,N_13204);
and U15837 (N_15837,N_12804,N_12868);
nor U15838 (N_15838,N_14693,N_13016);
nor U15839 (N_15839,N_13095,N_14457);
nor U15840 (N_15840,N_13746,N_12895);
and U15841 (N_15841,N_13104,N_13472);
nand U15842 (N_15842,N_13858,N_15541);
nor U15843 (N_15843,N_14139,N_13832);
nand U15844 (N_15844,N_13689,N_14925);
nand U15845 (N_15845,N_15366,N_14630);
and U15846 (N_15846,N_12647,N_14536);
and U15847 (N_15847,N_15476,N_15271);
nand U15848 (N_15848,N_14589,N_13641);
or U15849 (N_15849,N_14486,N_12798);
nor U15850 (N_15850,N_13518,N_13691);
nand U15851 (N_15851,N_14129,N_12726);
nor U15852 (N_15852,N_13123,N_13686);
or U15853 (N_15853,N_15169,N_12814);
nand U15854 (N_15854,N_13295,N_14433);
xor U15855 (N_15855,N_13751,N_13660);
nor U15856 (N_15856,N_13148,N_15012);
or U15857 (N_15857,N_12812,N_14704);
nand U15858 (N_15858,N_12958,N_13401);
nand U15859 (N_15859,N_14841,N_13086);
xnor U15860 (N_15860,N_15422,N_14697);
xnor U15861 (N_15861,N_13162,N_14345);
nand U15862 (N_15862,N_14053,N_14213);
or U15863 (N_15863,N_12828,N_15459);
and U15864 (N_15864,N_12961,N_13351);
nand U15865 (N_15865,N_13214,N_12630);
or U15866 (N_15866,N_13174,N_14150);
nand U15867 (N_15867,N_12972,N_13247);
and U15868 (N_15868,N_14728,N_15609);
nor U15869 (N_15869,N_15329,N_12506);
or U15870 (N_15870,N_14128,N_14899);
and U15871 (N_15871,N_14242,N_14094);
xnor U15872 (N_15872,N_12947,N_13064);
and U15873 (N_15873,N_12940,N_15092);
nand U15874 (N_15874,N_14274,N_12872);
or U15875 (N_15875,N_12745,N_14130);
nor U15876 (N_15876,N_14409,N_13335);
and U15877 (N_15877,N_12878,N_15134);
and U15878 (N_15878,N_13028,N_15125);
nor U15879 (N_15879,N_14636,N_13607);
nor U15880 (N_15880,N_13327,N_12756);
and U15881 (N_15881,N_13219,N_15355);
xnor U15882 (N_15882,N_13445,N_13964);
nor U15883 (N_15883,N_13459,N_13730);
or U15884 (N_15884,N_14850,N_14349);
or U15885 (N_15885,N_15048,N_12739);
nor U15886 (N_15886,N_14319,N_14963);
or U15887 (N_15887,N_12801,N_14620);
or U15888 (N_15888,N_15078,N_14573);
or U15889 (N_15889,N_15442,N_15067);
nand U15890 (N_15890,N_12747,N_15159);
and U15891 (N_15891,N_13760,N_14171);
xnor U15892 (N_15892,N_13840,N_14953);
or U15893 (N_15893,N_14072,N_14123);
xnor U15894 (N_15894,N_15246,N_12652);
nand U15895 (N_15895,N_12561,N_12764);
nor U15896 (N_15896,N_13255,N_15574);
nand U15897 (N_15897,N_15466,N_14571);
and U15898 (N_15898,N_15339,N_14683);
nor U15899 (N_15899,N_15130,N_14558);
and U15900 (N_15900,N_13777,N_13344);
nand U15901 (N_15901,N_13234,N_12761);
and U15902 (N_15902,N_13866,N_13488);
and U15903 (N_15903,N_13049,N_13404);
and U15904 (N_15904,N_13017,N_14112);
nor U15905 (N_15905,N_15474,N_13794);
and U15906 (N_15906,N_14956,N_15220);
nor U15907 (N_15907,N_14629,N_15077);
and U15908 (N_15908,N_13346,N_12824);
nor U15909 (N_15909,N_14048,N_14148);
xnor U15910 (N_15910,N_13993,N_15249);
nor U15911 (N_15911,N_15370,N_14191);
nand U15912 (N_15912,N_14062,N_13355);
nand U15913 (N_15913,N_14018,N_15307);
nor U15914 (N_15914,N_13576,N_12692);
xor U15915 (N_15915,N_14826,N_15477);
nand U15916 (N_15916,N_14180,N_13608);
or U15917 (N_15917,N_14591,N_13879);
nand U15918 (N_15918,N_13628,N_12808);
nand U15919 (N_15919,N_14830,N_12570);
or U15920 (N_15920,N_13869,N_13791);
nor U15921 (N_15921,N_15100,N_14501);
or U15922 (N_15922,N_14227,N_12638);
nor U15923 (N_15923,N_14504,N_14115);
nor U15924 (N_15924,N_14189,N_14464);
or U15925 (N_15925,N_12780,N_14027);
nor U15926 (N_15926,N_13015,N_15148);
and U15927 (N_15927,N_13623,N_13319);
or U15928 (N_15928,N_14758,N_13508);
or U15929 (N_15929,N_12908,N_14216);
nand U15930 (N_15930,N_12671,N_15126);
nand U15931 (N_15931,N_15436,N_14907);
xor U15932 (N_15932,N_14442,N_13597);
and U15933 (N_15933,N_12679,N_14540);
xnor U15934 (N_15934,N_14761,N_14204);
nand U15935 (N_15935,N_13066,N_13366);
and U15936 (N_15936,N_15461,N_15496);
nor U15937 (N_15937,N_13977,N_14831);
or U15938 (N_15938,N_14284,N_12691);
nor U15939 (N_15939,N_13897,N_14705);
or U15940 (N_15940,N_14905,N_14069);
nor U15941 (N_15941,N_15133,N_15475);
nand U15942 (N_15942,N_14125,N_13995);
nor U15943 (N_15943,N_14401,N_15566);
xor U15944 (N_15944,N_13939,N_14254);
nand U15945 (N_15945,N_14658,N_14034);
or U15946 (N_15946,N_15076,N_12730);
or U15947 (N_15947,N_15588,N_15558);
nor U15948 (N_15948,N_13245,N_13325);
and U15949 (N_15949,N_13567,N_13765);
or U15950 (N_15950,N_14101,N_12667);
or U15951 (N_15951,N_13176,N_14373);
or U15952 (N_15952,N_13790,N_13304);
or U15953 (N_15953,N_14283,N_14007);
nand U15954 (N_15954,N_14416,N_13291);
xnor U15955 (N_15955,N_12707,N_13590);
or U15956 (N_15956,N_12985,N_15330);
nand U15957 (N_15957,N_12720,N_15562);
or U15958 (N_15958,N_13192,N_12945);
or U15959 (N_15959,N_12645,N_12871);
and U15960 (N_15960,N_14074,N_13896);
nand U15961 (N_15961,N_12505,N_13996);
xnor U15962 (N_15962,N_14757,N_14842);
nand U15963 (N_15963,N_13252,N_13236);
or U15964 (N_15964,N_13296,N_12621);
nor U15965 (N_15965,N_12784,N_14182);
or U15966 (N_15966,N_13166,N_15272);
or U15967 (N_15967,N_12800,N_14853);
and U15968 (N_15968,N_12637,N_14530);
or U15969 (N_15969,N_14095,N_14393);
or U15970 (N_15970,N_13187,N_13653);
nor U15971 (N_15971,N_14851,N_13143);
nand U15972 (N_15972,N_15162,N_14121);
and U15973 (N_15973,N_14145,N_14859);
and U15974 (N_15974,N_15093,N_14088);
or U15975 (N_15975,N_13469,N_13061);
or U15976 (N_15976,N_13458,N_14517);
and U15977 (N_15977,N_12677,N_13530);
xnor U15978 (N_15978,N_12557,N_13119);
and U15979 (N_15979,N_15267,N_13723);
nand U15980 (N_15980,N_15441,N_15139);
nor U15981 (N_15981,N_14993,N_15167);
and U15982 (N_15982,N_15353,N_15081);
nor U15983 (N_15983,N_13714,N_12737);
nand U15984 (N_15984,N_13090,N_13717);
and U15985 (N_15985,N_12522,N_13497);
or U15986 (N_15986,N_15357,N_14080);
and U15987 (N_15987,N_13815,N_13708);
nand U15988 (N_15988,N_14714,N_12591);
nand U15989 (N_15989,N_15113,N_14231);
or U15990 (N_15990,N_14120,N_13467);
or U15991 (N_15991,N_13664,N_15580);
and U15992 (N_15992,N_12610,N_13990);
xor U15993 (N_15993,N_12740,N_13268);
or U15994 (N_15994,N_12765,N_13068);
nand U15995 (N_15995,N_15292,N_13758);
and U15996 (N_15996,N_15238,N_15494);
and U15997 (N_15997,N_14555,N_14986);
nor U15998 (N_15998,N_13907,N_13911);
and U15999 (N_15999,N_12620,N_13729);
nand U16000 (N_16000,N_14494,N_14339);
xor U16001 (N_16001,N_14557,N_13805);
xnor U16002 (N_16002,N_12714,N_13147);
or U16003 (N_16003,N_14023,N_14286);
nand U16004 (N_16004,N_14175,N_14485);
nand U16005 (N_16005,N_14524,N_12969);
nand U16006 (N_16006,N_14784,N_15623);
and U16007 (N_16007,N_12820,N_14376);
and U16008 (N_16008,N_14168,N_13957);
nand U16009 (N_16009,N_13126,N_15402);
or U16010 (N_16010,N_15143,N_13449);
nand U16011 (N_16011,N_12914,N_14660);
or U16012 (N_16012,N_13888,N_15406);
nand U16013 (N_16013,N_12964,N_13727);
nand U16014 (N_16014,N_12862,N_15110);
and U16015 (N_16015,N_12500,N_13545);
and U16016 (N_16016,N_13948,N_12684);
nor U16017 (N_16017,N_15534,N_13787);
and U16018 (N_16018,N_12823,N_13638);
and U16019 (N_16019,N_15250,N_14156);
nand U16020 (N_16020,N_14498,N_12974);
nor U16021 (N_16021,N_13822,N_14910);
or U16022 (N_16022,N_14310,N_13253);
and U16023 (N_16023,N_14880,N_15288);
or U16024 (N_16024,N_14838,N_13812);
or U16025 (N_16025,N_13083,N_15281);
and U16026 (N_16026,N_15075,N_12586);
nor U16027 (N_16027,N_14975,N_13570);
nor U16028 (N_16028,N_12587,N_15407);
nand U16029 (N_16029,N_12817,N_14818);
or U16030 (N_16030,N_14964,N_14118);
nor U16031 (N_16031,N_13793,N_14817);
or U16032 (N_16032,N_14009,N_14078);
and U16033 (N_16033,N_13839,N_13702);
and U16034 (N_16034,N_13885,N_14679);
nor U16035 (N_16035,N_13282,N_12752);
and U16036 (N_16036,N_15501,N_13901);
or U16037 (N_16037,N_13314,N_15350);
nor U16038 (N_16038,N_13289,N_12896);
nand U16039 (N_16039,N_14482,N_14366);
nand U16040 (N_16040,N_14802,N_15349);
xor U16041 (N_16041,N_14402,N_13360);
xor U16042 (N_16042,N_15392,N_14331);
or U16043 (N_16043,N_15340,N_13213);
or U16044 (N_16044,N_12583,N_14408);
nor U16045 (N_16045,N_14045,N_13984);
nor U16046 (N_16046,N_14424,N_12893);
and U16047 (N_16047,N_15018,N_12641);
nor U16048 (N_16048,N_12782,N_15156);
or U16049 (N_16049,N_14695,N_12889);
xor U16050 (N_16050,N_13818,N_14869);
nand U16051 (N_16051,N_13548,N_14378);
and U16052 (N_16052,N_14970,N_12848);
nand U16053 (N_16053,N_13855,N_13747);
or U16054 (N_16054,N_14535,N_15136);
nand U16055 (N_16055,N_14008,N_15103);
or U16056 (N_16056,N_13019,N_14032);
or U16057 (N_16057,N_15039,N_13523);
or U16058 (N_16058,N_15176,N_13644);
or U16059 (N_16059,N_13603,N_15336);
nand U16060 (N_16060,N_13376,N_13748);
or U16061 (N_16061,N_14474,N_12609);
or U16062 (N_16062,N_14028,N_13407);
xnor U16063 (N_16063,N_12927,N_15570);
nor U16064 (N_16064,N_13854,N_15099);
and U16065 (N_16065,N_14631,N_13771);
and U16066 (N_16066,N_13949,N_15322);
and U16067 (N_16067,N_15280,N_13631);
or U16068 (N_16068,N_15378,N_13347);
and U16069 (N_16069,N_15543,N_13916);
nand U16070 (N_16070,N_14673,N_13906);
and U16071 (N_16071,N_15135,N_12774);
or U16072 (N_16072,N_15231,N_14152);
nor U16073 (N_16073,N_15268,N_13501);
xnor U16074 (N_16074,N_13233,N_14258);
nand U16075 (N_16075,N_13188,N_13937);
xnor U16076 (N_16076,N_14894,N_13400);
nor U16077 (N_16077,N_14014,N_15131);
xnor U16078 (N_16078,N_14878,N_13439);
nor U16079 (N_16079,N_14199,N_15393);
and U16080 (N_16080,N_14748,N_14406);
and U16081 (N_16081,N_15400,N_14598);
and U16082 (N_16082,N_13085,N_13030);
and U16083 (N_16083,N_15387,N_13733);
xor U16084 (N_16084,N_13584,N_13573);
and U16085 (N_16085,N_15528,N_12532);
or U16086 (N_16086,N_14091,N_12869);
nor U16087 (N_16087,N_15343,N_14985);
nor U16088 (N_16088,N_15054,N_15401);
and U16089 (N_16089,N_12916,N_13795);
and U16090 (N_16090,N_13020,N_13533);
nor U16091 (N_16091,N_14126,N_14483);
or U16092 (N_16092,N_15086,N_13946);
or U16093 (N_16093,N_13096,N_15513);
or U16094 (N_16094,N_13353,N_14682);
and U16095 (N_16095,N_13710,N_15233);
and U16096 (N_16096,N_12884,N_13372);
or U16097 (N_16097,N_12951,N_13369);
nor U16098 (N_16098,N_15111,N_12642);
nand U16099 (N_16099,N_14523,N_14994);
and U16100 (N_16100,N_14525,N_14978);
and U16101 (N_16101,N_14774,N_14825);
or U16102 (N_16102,N_13359,N_15413);
or U16103 (N_16103,N_15484,N_13320);
nand U16104 (N_16104,N_13262,N_15222);
and U16105 (N_16105,N_12666,N_15223);
nor U16106 (N_16106,N_15326,N_15175);
nand U16107 (N_16107,N_14073,N_14703);
and U16108 (N_16108,N_13071,N_14099);
or U16109 (N_16109,N_15021,N_15384);
xnor U16110 (N_16110,N_13809,N_14471);
xor U16111 (N_16111,N_13322,N_14756);
nor U16112 (N_16112,N_14549,N_15454);
nor U16113 (N_16113,N_12879,N_13053);
xnor U16114 (N_16114,N_13427,N_12687);
nor U16115 (N_16115,N_13859,N_12575);
nor U16116 (N_16116,N_13800,N_15293);
or U16117 (N_16117,N_14766,N_14279);
and U16118 (N_16118,N_13405,N_13378);
and U16119 (N_16119,N_14713,N_14361);
xnor U16120 (N_16120,N_14740,N_12703);
nor U16121 (N_16121,N_14367,N_13184);
nand U16122 (N_16122,N_14585,N_15607);
or U16123 (N_16123,N_12509,N_14696);
and U16124 (N_16124,N_14608,N_13417);
nor U16125 (N_16125,N_15546,N_15026);
and U16126 (N_16126,N_15089,N_15470);
or U16127 (N_16127,N_15583,N_15161);
nand U16128 (N_16128,N_13055,N_13810);
nand U16129 (N_16129,N_13769,N_13863);
nor U16130 (N_16130,N_15451,N_14699);
xor U16131 (N_16131,N_14618,N_15283);
and U16132 (N_16132,N_12539,N_14944);
and U16133 (N_16133,N_13811,N_14848);
nand U16134 (N_16134,N_15482,N_14593);
nor U16135 (N_16135,N_14783,N_13196);
and U16136 (N_16136,N_13720,N_13358);
or U16137 (N_16137,N_12831,N_12792);
nor U16138 (N_16138,N_12516,N_12682);
nor U16139 (N_16139,N_13450,N_13529);
nor U16140 (N_16140,N_12883,N_14217);
and U16141 (N_16141,N_14522,N_14006);
nor U16142 (N_16142,N_14060,N_14924);
and U16143 (N_16143,N_14312,N_14891);
nand U16144 (N_16144,N_13452,N_12866);
or U16145 (N_16145,N_12886,N_12781);
or U16146 (N_16146,N_12695,N_13742);
and U16147 (N_16147,N_12712,N_15569);
and U16148 (N_16148,N_13826,N_13574);
nor U16149 (N_16149,N_14904,N_12525);
or U16150 (N_16150,N_14326,N_12887);
nor U16151 (N_16151,N_13909,N_13172);
or U16152 (N_16152,N_12822,N_13898);
nor U16153 (N_16153,N_15373,N_12622);
nand U16154 (N_16154,N_13626,N_13736);
or U16155 (N_16155,N_12939,N_13113);
nor U16156 (N_16156,N_13175,N_13482);
or U16157 (N_16157,N_13127,N_12504);
nor U16158 (N_16158,N_14211,N_14562);
or U16159 (N_16159,N_14547,N_12806);
or U16160 (N_16160,N_14159,N_13986);
or U16161 (N_16161,N_14475,N_13605);
and U16162 (N_16162,N_13987,N_14106);
or U16163 (N_16163,N_14019,N_14566);
and U16164 (N_16164,N_15559,N_14275);
and U16165 (N_16165,N_15219,N_15334);
nor U16166 (N_16166,N_14997,N_15405);
nor U16167 (N_16167,N_13315,N_12968);
or U16168 (N_16168,N_12673,N_14301);
xor U16169 (N_16169,N_12578,N_14808);
or U16170 (N_16170,N_15104,N_12510);
nor U16171 (N_16171,N_14183,N_15259);
xor U16172 (N_16172,N_12852,N_12918);
nand U16173 (N_16173,N_14815,N_14867);
and U16174 (N_16174,N_13613,N_13505);
and U16175 (N_16175,N_15080,N_12704);
or U16176 (N_16176,N_13834,N_12653);
xor U16177 (N_16177,N_15253,N_14033);
and U16178 (N_16178,N_15164,N_14384);
nand U16179 (N_16179,N_13766,N_13535);
or U16180 (N_16180,N_13543,N_13180);
and U16181 (N_16181,N_14021,N_12833);
or U16182 (N_16182,N_14155,N_15300);
nand U16183 (N_16183,N_14394,N_15548);
nand U16184 (N_16184,N_14508,N_13731);
xor U16185 (N_16185,N_13772,N_15212);
xnor U16186 (N_16186,N_15165,N_14372);
and U16187 (N_16187,N_13934,N_13272);
or U16188 (N_16188,N_15564,N_13169);
nor U16189 (N_16189,N_14335,N_15419);
xor U16190 (N_16190,N_13364,N_12929);
or U16191 (N_16191,N_12619,N_14462);
nor U16192 (N_16192,N_14928,N_15255);
and U16193 (N_16193,N_13825,N_14281);
nor U16194 (N_16194,N_13624,N_14506);
and U16195 (N_16195,N_12503,N_12742);
xor U16196 (N_16196,N_13380,N_15356);
nand U16197 (N_16197,N_12676,N_14669);
nand U16198 (N_16198,N_15311,N_13554);
and U16199 (N_16199,N_15338,N_14392);
nand U16200 (N_16200,N_14539,N_13817);
nand U16201 (N_16201,N_13558,N_12689);
and U16202 (N_16202,N_13634,N_15269);
nand U16203 (N_16203,N_13178,N_15538);
xor U16204 (N_16204,N_13097,N_14723);
nand U16205 (N_16205,N_14257,N_13988);
or U16206 (N_16206,N_14056,N_12759);
nor U16207 (N_16207,N_15109,N_14110);
nand U16208 (N_16208,N_12885,N_14976);
or U16209 (N_16209,N_13814,N_14996);
or U16210 (N_16210,N_12599,N_15510);
or U16211 (N_16211,N_14024,N_13437);
nor U16212 (N_16212,N_14396,N_14116);
nor U16213 (N_16213,N_13673,N_13381);
nor U16214 (N_16214,N_12705,N_13761);
nor U16215 (N_16215,N_12633,N_12659);
or U16216 (N_16216,N_15205,N_13365);
or U16217 (N_16217,N_14550,N_13249);
xnor U16218 (N_16218,N_13551,N_13018);
and U16219 (N_16219,N_14998,N_12851);
nand U16220 (N_16220,N_14249,N_12636);
or U16221 (N_16221,N_12526,N_13433);
or U16222 (N_16222,N_12794,N_13464);
xnor U16223 (N_16223,N_13559,N_14977);
xnor U16224 (N_16224,N_13447,N_14410);
and U16225 (N_16225,N_13397,N_13770);
nand U16226 (N_16226,N_15019,N_13035);
nand U16227 (N_16227,N_14496,N_14265);
nand U16228 (N_16228,N_14397,N_15491);
xnor U16229 (N_16229,N_14149,N_13239);
nor U16230 (N_16230,N_13538,N_14980);
or U16231 (N_16231,N_14382,N_15593);
and U16232 (N_16232,N_14672,N_15198);
or U16233 (N_16233,N_14897,N_12813);
and U16234 (N_16234,N_14553,N_15294);
nor U16235 (N_16235,N_14253,N_14600);
or U16236 (N_16236,N_15327,N_15425);
nand U16237 (N_16237,N_15043,N_13294);
nand U16238 (N_16238,N_13198,N_13967);
nand U16239 (N_16239,N_14218,N_13577);
nand U16240 (N_16240,N_13217,N_13606);
nand U16241 (N_16241,N_13612,N_15471);
or U16242 (N_16242,N_15318,N_12830);
nand U16243 (N_16243,N_15575,N_15239);
and U16244 (N_16244,N_14529,N_14369);
and U16245 (N_16245,N_15463,N_12826);
and U16246 (N_16246,N_14796,N_13849);
and U16247 (N_16247,N_14596,N_12565);
xnor U16248 (N_16248,N_15352,N_15097);
nand U16249 (N_16249,N_13410,N_15030);
and U16250 (N_16250,N_14089,N_14133);
or U16251 (N_16251,N_13021,N_13225);
nand U16252 (N_16252,N_14749,N_15060);
nor U16253 (N_16253,N_15443,N_13923);
nand U16254 (N_16254,N_13985,N_15264);
xnor U16255 (N_16255,N_12668,N_14579);
and U16256 (N_16256,N_14844,N_13312);
nor U16257 (N_16257,N_14441,N_13560);
and U16258 (N_16258,N_15410,N_15171);
or U16259 (N_16259,N_13412,N_14164);
nor U16260 (N_16260,N_13940,N_13442);
and U16261 (N_16261,N_13738,N_15617);
xnor U16262 (N_16262,N_15622,N_14794);
nand U16263 (N_16263,N_15191,N_12987);
or U16264 (N_16264,N_13683,N_14568);
and U16265 (N_16265,N_15417,N_14386);
nand U16266 (N_16266,N_13847,N_13737);
or U16267 (N_16267,N_15608,N_13785);
or U16268 (N_16268,N_14131,N_14479);
nor U16269 (N_16269,N_14889,N_13830);
nand U16270 (N_16270,N_14082,N_15297);
and U16271 (N_16271,N_14293,N_13872);
and U16272 (N_16272,N_12521,N_15185);
nand U16273 (N_16273,N_13589,N_13968);
or U16274 (N_16274,N_13684,N_13414);
nand U16275 (N_16275,N_15377,N_12979);
and U16276 (N_16276,N_14552,N_13677);
or U16277 (N_16277,N_13971,N_14544);
nand U16278 (N_16278,N_13444,N_13201);
nand U16279 (N_16279,N_12654,N_14574);
or U16280 (N_16280,N_14225,N_15119);
nand U16281 (N_16281,N_14751,N_13784);
and U16282 (N_16282,N_13780,N_14157);
xnor U16283 (N_16283,N_14921,N_14046);
nor U16284 (N_16284,N_12952,N_14011);
nor U16285 (N_16285,N_13675,N_13889);
or U16286 (N_16286,N_15478,N_13339);
or U16287 (N_16287,N_13629,N_14734);
nand U16288 (N_16288,N_14356,N_15605);
or U16289 (N_16289,N_12665,N_14083);
nor U16290 (N_16290,N_15069,N_14086);
nor U16291 (N_16291,N_14864,N_12554);
and U16292 (N_16292,N_14350,N_13596);
nor U16293 (N_16293,N_14786,N_15505);
and U16294 (N_16294,N_12550,N_14736);
nor U16295 (N_16295,N_12982,N_14461);
nand U16296 (N_16296,N_13598,N_15530);
and U16297 (N_16297,N_13828,N_13602);
or U16298 (N_16298,N_12640,N_15007);
and U16299 (N_16299,N_13311,N_12912);
nor U16300 (N_16300,N_12787,N_13230);
and U16301 (N_16301,N_12579,N_13796);
xnor U16302 (N_16302,N_14617,N_12991);
and U16303 (N_16303,N_14186,N_12797);
nand U16304 (N_16304,N_13781,N_12754);
nand U16305 (N_16305,N_14586,N_13048);
nor U16306 (N_16306,N_13227,N_14707);
nand U16307 (N_16307,N_14644,N_12937);
and U16308 (N_16308,N_14816,N_15016);
and U16309 (N_16309,N_15383,N_13637);
nand U16310 (N_16310,N_12861,N_15295);
or U16311 (N_16311,N_13121,N_14824);
nor U16312 (N_16312,N_15449,N_12688);
nand U16313 (N_16313,N_14105,N_15615);
xor U16314 (N_16314,N_14806,N_13982);
nand U16315 (N_16315,N_15121,N_13969);
nand U16316 (N_16316,N_15563,N_12864);
nand U16317 (N_16317,N_13337,N_12536);
and U16318 (N_16318,N_15279,N_13593);
and U16319 (N_16319,N_14472,N_12573);
nor U16320 (N_16320,N_12905,N_14035);
and U16321 (N_16321,N_13195,N_14065);
nand U16322 (N_16322,N_14103,N_13212);
or U16323 (N_16323,N_13992,N_14179);
and U16324 (N_16324,N_14640,N_13130);
and U16325 (N_16325,N_13081,N_14434);
nor U16326 (N_16326,N_14984,N_14854);
or U16327 (N_16327,N_13426,N_13886);
and U16328 (N_16328,N_15029,N_13423);
or U16329 (N_16329,N_15616,N_13552);
nor U16330 (N_16330,N_13357,N_13775);
or U16331 (N_16331,N_13483,N_13057);
nor U16332 (N_16332,N_15041,N_12928);
nand U16333 (N_16333,N_15166,N_15195);
nor U16334 (N_16334,N_14203,N_13137);
and U16335 (N_16335,N_15469,N_14775);
nand U16336 (N_16336,N_14291,N_13008);
or U16337 (N_16337,N_13711,N_15221);
or U16338 (N_16338,N_14041,N_14497);
nand U16339 (N_16339,N_14887,N_14839);
nand U16340 (N_16340,N_15070,N_13938);
and U16341 (N_16341,N_15553,N_13917);
or U16342 (N_16342,N_12930,N_15011);
nand U16343 (N_16343,N_13248,N_15042);
nand U16344 (N_16344,N_14922,N_14962);
nor U16345 (N_16345,N_13059,N_15380);
and U16346 (N_16346,N_13313,N_12909);
and U16347 (N_16347,N_15286,N_14900);
xnor U16348 (N_16348,N_14206,N_13256);
or U16349 (N_16349,N_12894,N_14063);
xor U16350 (N_16350,N_13037,N_14419);
nand U16351 (N_16351,N_13991,N_14285);
nor U16352 (N_16352,N_13837,N_13106);
nand U16353 (N_16353,N_14857,N_15218);
and U16354 (N_16354,N_13406,N_15296);
xor U16355 (N_16355,N_12818,N_14701);
nor U16356 (N_16356,N_14140,N_12571);
and U16357 (N_16357,N_13667,N_14898);
or U16358 (N_16358,N_13719,N_13418);
and U16359 (N_16359,N_15324,N_14792);
nor U16360 (N_16360,N_13191,N_13181);
nor U16361 (N_16361,N_13435,N_13952);
and U16362 (N_16362,N_13599,N_12651);
nor U16363 (N_16363,N_12686,N_15518);
nor U16364 (N_16364,N_13089,N_14003);
or U16365 (N_16365,N_15201,N_12559);
nand U16366 (N_16366,N_15124,N_14495);
or U16367 (N_16367,N_12706,N_14868);
and U16368 (N_16368,N_15226,N_12920);
xor U16369 (N_16369,N_13402,N_14309);
and U16370 (N_16370,N_15508,N_15544);
or U16371 (N_16371,N_13461,N_13453);
nor U16372 (N_16372,N_13443,N_15582);
or U16373 (N_16373,N_13395,N_14503);
and U16374 (N_16374,N_15240,N_13141);
and U16375 (N_16375,N_13203,N_15369);
and U16376 (N_16376,N_13159,N_14163);
nor U16377 (N_16377,N_13224,N_15098);
and U16378 (N_16378,N_14684,N_15073);
and U16379 (N_16379,N_12533,N_12612);
nor U16380 (N_16380,N_12897,N_13681);
nor U16381 (N_16381,N_14246,N_14198);
and U16382 (N_16382,N_14567,N_12511);
nor U16383 (N_16383,N_13051,N_12709);
or U16384 (N_16384,N_12966,N_15375);
and U16385 (N_16385,N_13215,N_14668);
nor U16386 (N_16386,N_13163,N_13619);
or U16387 (N_16387,N_15129,N_14311);
nand U16388 (N_16388,N_14676,N_14143);
and U16389 (N_16389,N_15430,N_12924);
nor U16390 (N_16390,N_12746,N_13630);
or U16391 (N_16391,N_13878,N_13694);
nor U16392 (N_16392,N_12996,N_13279);
nor U16393 (N_16393,N_15473,N_15423);
nor U16394 (N_16394,N_15079,N_15310);
nor U16395 (N_16395,N_13774,N_12832);
nor U16396 (N_16396,N_14188,N_15492);
or U16397 (N_16397,N_15287,N_13011);
nor U16398 (N_16398,N_12875,N_12999);
xor U16399 (N_16399,N_15504,N_13956);
or U16400 (N_16400,N_14320,N_13942);
nor U16401 (N_16401,N_14344,N_14548);
and U16402 (N_16402,N_15497,N_13513);
xor U16403 (N_16403,N_15363,N_15592);
xnor U16404 (N_16404,N_14154,N_12716);
nand U16405 (N_16405,N_15256,N_13185);
and U16406 (N_16406,N_13945,N_13076);
xnor U16407 (N_16407,N_14967,N_15305);
or U16408 (N_16408,N_14908,N_14491);
nor U16409 (N_16409,N_14181,N_14059);
and U16410 (N_16410,N_15596,N_12750);
nand U16411 (N_16411,N_12582,N_13905);
xnor U16412 (N_16412,N_14559,N_14421);
or U16413 (N_16413,N_15050,N_14685);
or U16414 (N_16414,N_13755,N_14013);
nand U16415 (N_16415,N_13371,N_15184);
nor U16416 (N_16416,N_15087,N_13379);
nand U16417 (N_16417,N_12855,N_12917);
or U16418 (N_16418,N_13801,N_14719);
nor U16419 (N_16419,N_14691,N_14307);
xnor U16420 (N_16420,N_13520,N_13208);
nand U16421 (N_16421,N_14114,N_14732);
or U16422 (N_16422,N_14881,N_12670);
nor U16423 (N_16423,N_15341,N_14753);
xor U16424 (N_16424,N_14754,N_14541);
or U16425 (N_16425,N_12900,N_13564);
nand U16426 (N_16426,N_15128,N_14268);
nor U16427 (N_16427,N_12593,N_15557);
and U16428 (N_16428,N_14379,N_14407);
nand U16429 (N_16429,N_14771,N_12880);
and U16430 (N_16430,N_12632,N_14147);
xor U16431 (N_16431,N_15031,N_15418);
or U16432 (N_16432,N_15278,N_12562);
or U16433 (N_16433,N_14108,N_13514);
nor U16434 (N_16434,N_14777,N_12644);
and U16435 (N_16435,N_12838,N_12807);
and U16436 (N_16436,N_13656,N_13451);
nand U16437 (N_16437,N_15034,N_14337);
xor U16438 (N_16438,N_14999,N_13713);
and U16439 (N_16439,N_14972,N_15404);
nor U16440 (N_16440,N_13652,N_13431);
xor U16441 (N_16441,N_15437,N_15560);
and U16442 (N_16442,N_14360,N_12639);
or U16443 (N_16443,N_12513,N_12572);
nand U16444 (N_16444,N_13853,N_13486);
or U16445 (N_16445,N_12865,N_12935);
and U16446 (N_16446,N_13750,N_14930);
and U16447 (N_16447,N_15433,N_13246);
or U16448 (N_16448,N_15170,N_14863);
or U16449 (N_16449,N_15519,N_15002);
and U16450 (N_16450,N_14526,N_15493);
nor U16451 (N_16451,N_15498,N_15550);
and U16452 (N_16452,N_13374,N_13151);
or U16453 (N_16453,N_12574,N_15577);
or U16454 (N_16454,N_15025,N_15263);
nor U16455 (N_16455,N_12541,N_15321);
nor U16456 (N_16456,N_15337,N_13666);
or U16457 (N_16457,N_14174,N_14688);
or U16458 (N_16458,N_13361,N_14879);
nor U16459 (N_16459,N_15137,N_14654);
and U16460 (N_16460,N_15345,N_15479);
or U16461 (N_16461,N_13000,N_14377);
or U16462 (N_16462,N_14735,N_13920);
and U16463 (N_16463,N_14260,N_13052);
nand U16464 (N_16464,N_14870,N_15102);
or U16465 (N_16465,N_14251,N_12846);
or U16466 (N_16466,N_15331,N_15047);
or U16467 (N_16467,N_15056,N_15145);
nand U16468 (N_16468,N_14221,N_15348);
and U16469 (N_16469,N_13510,N_15052);
nor U16470 (N_16470,N_13915,N_15603);
nor U16471 (N_16471,N_13649,N_13328);
or U16472 (N_16472,N_13133,N_13009);
nor U16473 (N_16473,N_13725,N_13700);
nand U16474 (N_16474,N_13352,N_13073);
nor U16475 (N_16475,N_14235,N_13829);
nand U16476 (N_16476,N_14468,N_13640);
xnor U16477 (N_16477,N_15452,N_13383);
and U16478 (N_16478,N_13583,N_14689);
xor U16479 (N_16479,N_15068,N_14931);
or U16480 (N_16480,N_13425,N_13415);
and U16481 (N_16481,N_14604,N_14861);
or U16482 (N_16482,N_14671,N_13070);
nand U16483 (N_16483,N_13693,N_15106);
nand U16484 (N_16484,N_14516,N_14302);
nor U16485 (N_16485,N_14722,N_14374);
and U16486 (N_16486,N_14264,N_14465);
nor U16487 (N_16487,N_12777,N_14439);
nor U16488 (N_16488,N_13877,N_13604);
xnor U16489 (N_16489,N_14952,N_14942);
or U16490 (N_16490,N_14791,N_15127);
nor U16491 (N_16491,N_15013,N_13160);
nor U16492 (N_16492,N_14819,N_14230);
nand U16493 (N_16493,N_14317,N_14456);
nor U16494 (N_16494,N_15397,N_14973);
nand U16495 (N_16495,N_14570,N_14741);
and U16496 (N_16496,N_15247,N_13983);
or U16497 (N_16497,N_15027,N_13724);
nor U16498 (N_16498,N_15232,N_14561);
and U16499 (N_16499,N_13266,N_14743);
nand U16500 (N_16500,N_14820,N_15228);
and U16501 (N_16501,N_13846,N_14277);
or U16502 (N_16502,N_14030,N_14711);
nand U16503 (N_16503,N_12606,N_15038);
and U16504 (N_16504,N_13082,N_14228);
or U16505 (N_16505,N_13506,N_15509);
nand U16506 (N_16506,N_14239,N_13591);
nand U16507 (N_16507,N_13031,N_14632);
or U16508 (N_16508,N_13884,N_14941);
or U16509 (N_16509,N_13146,N_14760);
nor U16510 (N_16510,N_13892,N_15347);
nand U16511 (N_16511,N_14160,N_14588);
xor U16512 (N_16512,N_13487,N_14877);
and U16513 (N_16513,N_13421,N_14092);
nor U16514 (N_16514,N_13152,N_14883);
or U16515 (N_16515,N_14935,N_15512);
nand U16516 (N_16516,N_13099,N_14983);
xor U16517 (N_16517,N_14303,N_13135);
or U16518 (N_16518,N_13027,N_15391);
xor U16519 (N_16519,N_12508,N_13254);
xor U16520 (N_16520,N_13921,N_12773);
nand U16521 (N_16521,N_15434,N_14481);
or U16522 (N_16522,N_15091,N_12589);
or U16523 (N_16523,N_14849,N_12860);
and U16524 (N_16524,N_14039,N_15227);
nor U16525 (N_16525,N_13117,N_13918);
or U16526 (N_16526,N_14447,N_15364);
or U16527 (N_16527,N_15180,N_13561);
or U16528 (N_16528,N_13093,N_13807);
nand U16529 (N_16529,N_14621,N_14142);
nor U16530 (N_16530,N_13783,N_13285);
or U16531 (N_16531,N_13493,N_14538);
and U16532 (N_16532,N_14790,N_12723);
nand U16533 (N_16533,N_13354,N_15061);
nand U16534 (N_16534,N_15529,N_14178);
and U16535 (N_16535,N_13851,N_15457);
nand U16536 (N_16536,N_12735,N_14731);
nand U16537 (N_16537,N_14718,N_13757);
nand U16538 (N_16538,N_13250,N_14520);
nand U16539 (N_16539,N_14151,N_14431);
and U16540 (N_16540,N_13532,N_13284);
or U16541 (N_16541,N_15096,N_12881);
nor U16542 (N_16542,N_14690,N_12919);
nand U16543 (N_16543,N_12675,N_14084);
nor U16544 (N_16544,N_12802,N_15146);
nor U16545 (N_16545,N_14328,N_14117);
xor U16546 (N_16546,N_13281,N_13441);
nor U16547 (N_16547,N_14810,N_14214);
and U16548 (N_16548,N_15200,N_13056);
nor U16549 (N_16549,N_14680,N_14015);
and U16550 (N_16550,N_13084,N_15365);
and U16551 (N_16551,N_12711,N_15235);
nor U16552 (N_16552,N_14750,N_15526);
nor U16553 (N_16553,N_14659,N_13542);
and U16554 (N_16554,N_15465,N_12590);
nand U16555 (N_16555,N_14208,N_14909);
xnor U16556 (N_16556,N_12629,N_12960);
or U16557 (N_16557,N_14333,N_13831);
and U16558 (N_16558,N_15314,N_15527);
nand U16559 (N_16559,N_12849,N_15049);
nor U16560 (N_16560,N_13566,N_13517);
nand U16561 (N_16561,N_14044,N_13079);
nor U16562 (N_16562,N_14296,N_14981);
and U16563 (N_16563,N_14202,N_15033);
nor U16564 (N_16564,N_13171,N_13698);
xor U16565 (N_16565,N_12549,N_12911);
or U16566 (N_16566,N_14510,N_15599);
nand U16567 (N_16567,N_13323,N_13537);
and U16568 (N_16568,N_15209,N_12790);
or U16569 (N_16569,N_12713,N_14389);
nor U16570 (N_16570,N_13931,N_12520);
nor U16571 (N_16571,N_13136,N_12699);
nand U16572 (N_16572,N_12617,N_13672);
nor U16573 (N_16573,N_14611,N_13503);
nor U16574 (N_16574,N_13662,N_13883);
and U16575 (N_16575,N_14678,N_13300);
and U16576 (N_16576,N_14308,N_15085);
nor U16577 (N_16577,N_14686,N_12853);
nand U16578 (N_16578,N_13614,N_14959);
nand U16579 (N_16579,N_12799,N_13868);
xor U16580 (N_16580,N_15252,N_15429);
xor U16581 (N_16581,N_14122,N_13054);
nor U16582 (N_16582,N_15549,N_15511);
and U16583 (N_16583,N_12624,N_14004);
nand U16584 (N_16584,N_15120,N_13820);
and U16585 (N_16585,N_15036,N_14241);
nand U16586 (N_16586,N_12558,N_13474);
nand U16587 (N_16587,N_14893,N_12598);
or U16588 (N_16588,N_14603,N_13161);
or U16589 (N_16589,N_13023,N_14581);
nand U16590 (N_16590,N_12840,N_15084);
nor U16591 (N_16591,N_12717,N_12563);
and U16592 (N_16592,N_13739,N_13880);
nor U16593 (N_16593,N_13087,N_14294);
or U16594 (N_16594,N_13362,N_12749);
xnor U16595 (N_16595,N_14269,N_15168);
and U16596 (N_16596,N_13861,N_13363);
and U16597 (N_16597,N_14812,N_13490);
xor U16598 (N_16598,N_13269,N_15122);
and U16599 (N_16599,N_14584,N_15193);
nand U16600 (N_16600,N_14383,N_15024);
and U16601 (N_16601,N_13887,N_13194);
or U16602 (N_16602,N_15408,N_14661);
nor U16603 (N_16603,N_15290,N_13894);
or U16604 (N_16604,N_13072,N_13701);
or U16605 (N_16605,N_13504,N_14137);
or U16606 (N_16606,N_15573,N_14846);
or U16607 (N_16607,N_15182,N_14167);
nor U16608 (N_16608,N_12540,N_14390);
and U16609 (N_16609,N_14425,N_15316);
xor U16610 (N_16610,N_12537,N_12611);
nand U16611 (N_16611,N_13370,N_13540);
or U16612 (N_16612,N_12796,N_15424);
nor U16613 (N_16613,N_13223,N_14971);
nand U16614 (N_16614,N_14229,N_13876);
nand U16615 (N_16615,N_14780,N_15480);
and U16616 (N_16616,N_15524,N_14515);
and U16617 (N_16617,N_15242,N_13799);
nor U16618 (N_16618,N_14036,N_12845);
xor U16619 (N_16619,N_14936,N_13521);
nor U16620 (N_16620,N_15495,N_13881);
and U16621 (N_16621,N_14809,N_15153);
nand U16622 (N_16622,N_15196,N_12547);
and U16623 (N_16623,N_13283,N_12988);
or U16624 (N_16624,N_14306,N_14017);
nor U16625 (N_16625,N_14240,N_13836);
or U16626 (N_16626,N_13199,N_14698);
nor U16627 (N_16627,N_13804,N_12584);
and U16628 (N_16628,N_14519,N_15421);
nor U16629 (N_16629,N_14443,N_15536);
nor U16630 (N_16630,N_13509,N_12701);
or U16631 (N_16631,N_12715,N_13317);
nor U16632 (N_16632,N_14837,N_12615);
and U16633 (N_16633,N_13531,N_15114);
nor U16634 (N_16634,N_13536,N_15008);
nand U16635 (N_16635,N_13069,N_14651);
or U16636 (N_16636,N_12901,N_15517);
and U16637 (N_16637,N_12962,N_14347);
nand U16638 (N_16638,N_15556,N_14590);
and U16639 (N_16639,N_12743,N_14958);
nor U16640 (N_16640,N_14398,N_14951);
nor U16641 (N_16641,N_14594,N_15595);
or U16642 (N_16642,N_12597,N_12933);
nand U16643 (N_16643,N_14511,N_13500);
or U16644 (N_16644,N_12993,N_14960);
or U16645 (N_16645,N_12643,N_14950);
or U16646 (N_16646,N_13206,N_13806);
and U16647 (N_16647,N_15516,N_15225);
nand U16648 (N_16648,N_13900,N_13120);
nor U16649 (N_16649,N_12877,N_15460);
nand U16650 (N_16650,N_14276,N_13544);
nand U16651 (N_16651,N_13150,N_14762);
and U16652 (N_16652,N_14955,N_13972);
nor U16653 (N_16653,N_14146,N_15462);
xnor U16654 (N_16654,N_13385,N_14918);
nor U16655 (N_16655,N_14641,N_12708);
nand U16656 (N_16656,N_15427,N_13209);
or U16657 (N_16657,N_13819,N_14650);
and U16658 (N_16658,N_14551,N_13182);
nor U16659 (N_16659,N_13646,N_13103);
or U16660 (N_16660,N_14327,N_13636);
nor U16661 (N_16661,N_13430,N_12601);
and U16662 (N_16662,N_15521,N_14322);
nand U16663 (N_16663,N_13088,N_14210);
xor U16664 (N_16664,N_14220,N_13980);
or U16665 (N_16665,N_14172,N_13867);
or U16666 (N_16666,N_13507,N_12980);
or U16667 (N_16667,N_13962,N_13697);
and U16668 (N_16668,N_13813,N_13022);
nor U16669 (N_16669,N_13436,N_15612);
and U16670 (N_16670,N_15028,N_14365);
and U16671 (N_16671,N_15555,N_12942);
nand U16672 (N_16672,N_14124,N_15183);
nand U16673 (N_16673,N_12627,N_13671);
and U16674 (N_16674,N_14607,N_12955);
nor U16675 (N_16675,N_14633,N_12850);
or U16676 (N_16676,N_13321,N_14236);
nand U16677 (N_16677,N_13092,N_14420);
or U16678 (N_16678,N_14002,N_15186);
nand U16679 (N_16679,N_12614,N_15333);
nor U16680 (N_16680,N_15499,N_14299);
and U16681 (N_16681,N_13399,N_14763);
nor U16682 (N_16682,N_14057,N_15500);
nor U16683 (N_16683,N_14670,N_13661);
nand U16684 (N_16684,N_14417,N_13316);
or U16685 (N_16685,N_13575,N_13308);
nor U16686 (N_16686,N_14533,N_14026);
nand U16687 (N_16687,N_13808,N_14954);
nand U16688 (N_16688,N_15309,N_15503);
nand U16689 (N_16689,N_14244,N_13448);
xor U16690 (N_16690,N_14822,N_13525);
nand U16691 (N_16691,N_12724,N_12534);
or U16692 (N_16692,N_14843,N_15362);
nor U16693 (N_16693,N_13118,N_13556);
and U16694 (N_16694,N_15446,N_13953);
nor U16695 (N_16695,N_12931,N_15105);
or U16696 (N_16696,N_14195,N_12678);
xnor U16697 (N_16697,N_13305,N_13124);
or U16698 (N_16698,N_13338,N_14634);
nand U16699 (N_16699,N_12531,N_13462);
nand U16700 (N_16700,N_14102,N_12721);
nor U16701 (N_16701,N_13040,N_15117);
nor U16702 (N_16702,N_12891,N_14359);
xnor U16703 (N_16703,N_14259,N_14127);
xnor U16704 (N_16704,N_12825,N_14436);
nor U16705 (N_16705,N_15435,N_14991);
and U16706 (N_16706,N_15304,N_13726);
or U16707 (N_16707,N_13434,N_14637);
nand U16708 (N_16708,N_13342,N_15260);
nor U16709 (N_16709,N_12626,N_13334);
and U16710 (N_16710,N_12753,N_14628);
xnor U16711 (N_16711,N_14770,N_14798);
and U16712 (N_16712,N_13036,N_13622);
xor U16713 (N_16713,N_13446,N_12902);
nand U16714 (N_16714,N_13526,N_14692);
or U16715 (N_16715,N_13696,N_13112);
and U16716 (N_16716,N_14764,N_13025);
nor U16717 (N_16717,N_13632,N_15257);
nor U16718 (N_16718,N_13688,N_14119);
or U16719 (N_16719,N_13075,N_14316);
and U16720 (N_16720,N_15372,N_12778);
and U16721 (N_16721,N_13292,N_15481);
nand U16722 (N_16722,N_14769,N_13006);
nand U16723 (N_16723,N_13679,N_12859);
xor U16724 (N_16724,N_13158,N_13063);
and U16725 (N_16725,N_14813,N_15273);
nor U16726 (N_16726,N_13910,N_13373);
nor U16727 (N_16727,N_12515,N_14012);
nand U16728 (N_16728,N_15181,N_13961);
nand U16729 (N_16729,N_13331,N_12634);
and U16730 (N_16730,N_13032,N_12702);
and U16731 (N_16731,N_14717,N_15302);
xor U16732 (N_16732,N_15112,N_14648);
nor U16733 (N_16733,N_14646,N_15389);
xnor U16734 (N_16734,N_12925,N_15359);
and U16735 (N_16735,N_14487,N_13635);
nand U16736 (N_16736,N_14261,N_15053);
and U16737 (N_16737,N_14990,N_13131);
nand U16738 (N_16738,N_13065,N_14814);
nor U16739 (N_16739,N_14917,N_15177);
nand U16740 (N_16740,N_15598,N_13663);
or U16741 (N_16741,N_14554,N_13307);
or U16742 (N_16742,N_14610,N_13935);
or U16743 (N_16743,N_15261,N_14298);
nor U16744 (N_16744,N_12535,N_12948);
and U16745 (N_16745,N_13803,N_13924);
xor U16746 (N_16746,N_12816,N_14866);
and U16747 (N_16747,N_14505,N_14368);
and U16748 (N_16748,N_14563,N_14270);
or U16749 (N_16749,N_13620,N_12903);
nand U16750 (N_16750,N_15320,N_13963);
or U16751 (N_16751,N_13290,N_12858);
nand U16752 (N_16752,N_13202,N_13511);
nand U16753 (N_16753,N_13218,N_12954);
and U16754 (N_16754,N_14933,N_14029);
and U16755 (N_16755,N_13594,N_14797);
nand U16756 (N_16756,N_13454,N_14300);
xnor U16757 (N_16757,N_15157,N_13168);
and U16758 (N_16758,N_15274,N_15379);
nor U16759 (N_16759,N_13778,N_14085);
nor U16760 (N_16760,N_13498,N_13293);
and U16761 (N_16761,N_14077,N_14161);
or U16762 (N_16762,N_14860,N_13156);
xnor U16763 (N_16763,N_15390,N_14405);
nor U16764 (N_16764,N_12950,N_15386);
nor U16765 (N_16765,N_13833,N_15234);
and U16766 (N_16766,N_12922,N_13107);
or U16767 (N_16767,N_13844,N_14700);
xor U16768 (N_16768,N_14823,N_14836);
nand U16769 (N_16769,N_14966,N_13642);
or U16770 (N_16770,N_13838,N_13243);
nor U16771 (N_16771,N_13827,N_14988);
or U16772 (N_16772,N_15244,N_14974);
nor U16773 (N_16773,N_14071,N_14068);
or U16774 (N_16774,N_15083,N_15332);
nor U16775 (N_16775,N_15537,N_14040);
nand U16776 (N_16776,N_15396,N_12944);
or U16777 (N_16777,N_15456,N_14502);
xnor U16778 (N_16778,N_12811,N_14165);
nand U16779 (N_16779,N_13471,N_13534);
and U16780 (N_16780,N_12719,N_14847);
and U16781 (N_16781,N_14832,N_15040);
or U16782 (N_16782,N_13645,N_13303);
nand U16783 (N_16783,N_13014,N_15062);
or U16784 (N_16784,N_13394,N_14104);
and U16785 (N_16785,N_12932,N_14111);
nor U16786 (N_16786,N_12873,N_14400);
nand U16787 (N_16787,N_15115,N_14582);
xnor U16788 (N_16788,N_14097,N_13568);
and U16789 (N_16789,N_12662,N_12981);
nand U16790 (N_16790,N_15485,N_12669);
nor U16791 (N_16791,N_15539,N_15381);
nor U16792 (N_16792,N_12965,N_14289);
and U16793 (N_16793,N_13001,N_14343);
nand U16794 (N_16794,N_13565,N_15472);
or U16795 (N_16795,N_15224,N_14625);
or U16796 (N_16796,N_12835,N_14043);
nand U16797 (N_16797,N_13324,N_15063);
or U16798 (N_16798,N_14965,N_13024);
and U16799 (N_16799,N_14856,N_12527);
nor U16800 (N_16800,N_13302,N_12926);
nor U16801 (N_16801,N_13930,N_13929);
xor U16802 (N_16802,N_13391,N_12983);
or U16803 (N_16803,N_14675,N_13908);
and U16804 (N_16804,N_14720,N_12874);
and U16805 (N_16805,N_15141,N_13042);
or U16806 (N_16806,N_13848,N_13857);
and U16807 (N_16807,N_14336,N_13411);
nor U16808 (N_16808,N_15308,N_13329);
and U16809 (N_16809,N_13899,N_13581);
nor U16810 (N_16810,N_14426,N_13026);
or U16811 (N_16811,N_15515,N_12967);
or U16812 (N_16812,N_13745,N_13393);
nor U16813 (N_16813,N_15299,N_12564);
or U16814 (N_16814,N_15015,N_13232);
nand U16815 (N_16815,N_12656,N_13706);
nor U16816 (N_16816,N_12595,N_13572);
nand U16817 (N_16817,N_14801,N_12815);
or U16818 (N_16818,N_14833,N_15312);
and U16819 (N_16819,N_14793,N_13571);
xnor U16820 (N_16820,N_14914,N_14545);
nand U16821 (N_16821,N_13287,N_12836);
nand U16822 (N_16822,N_13633,N_14612);
nor U16823 (N_16823,N_14305,N_14042);
or U16824 (N_16824,N_14943,N_14215);
and U16825 (N_16825,N_13767,N_13041);
nand U16826 (N_16826,N_15448,N_14081);
or U16827 (N_16827,N_13286,N_13350);
or U16828 (N_16828,N_12844,N_12769);
nand U16829 (N_16829,N_13835,N_13046);
and U16830 (N_16830,N_13625,N_15624);
or U16831 (N_16831,N_12501,N_13913);
nor U16832 (N_16832,N_13549,N_13610);
and U16833 (N_16833,N_13382,N_14642);
nor U16834 (N_16834,N_14896,N_13010);
or U16835 (N_16835,N_12733,N_12847);
nor U16836 (N_16836,N_13502,N_14875);
xnor U16837 (N_16837,N_13336,N_14785);
nor U16838 (N_16838,N_14709,N_14196);
or U16839 (N_16839,N_14212,N_14050);
nor U16840 (N_16840,N_14313,N_14742);
and U16841 (N_16841,N_13078,N_13582);
nand U16842 (N_16842,N_14020,N_15428);
nand U16843 (N_16843,N_15545,N_14000);
or U16844 (N_16844,N_13226,N_13003);
or U16845 (N_16845,N_13718,N_14639);
nand U16846 (N_16846,N_12729,N_13216);
nand U16847 (N_16847,N_13356,N_12648);
xor U16848 (N_16848,N_12994,N_14263);
xor U16849 (N_16849,N_14458,N_13125);
or U16850 (N_16850,N_14542,N_13615);
xnor U16851 (N_16851,N_14388,N_14444);
xnor U16852 (N_16852,N_13722,N_14882);
and U16853 (N_16853,N_13387,N_15215);
nand U16854 (N_16854,N_14016,N_14687);
and U16855 (N_16855,N_13392,N_14025);
or U16856 (N_16856,N_13609,N_13231);
nor U16857 (N_16857,N_12734,N_13409);
or U16858 (N_16858,N_13659,N_15344);
nor U16859 (N_16859,N_15094,N_12906);
and U16860 (N_16860,N_15313,N_12867);
and U16861 (N_16861,N_15058,N_13332);
xor U16862 (N_16862,N_15001,N_15578);
and U16863 (N_16863,N_15597,N_15358);
and U16864 (N_16864,N_13721,N_13428);
nor U16865 (N_16865,N_15591,N_15017);
and U16866 (N_16866,N_14919,N_14341);
nand U16867 (N_16867,N_14412,N_14051);
and U16868 (N_16868,N_13965,N_14173);
nand U16869 (N_16869,N_14064,N_13244);
and U16870 (N_16870,N_12618,N_14324);
or U16871 (N_16871,N_13944,N_14674);
nor U16872 (N_16872,N_15174,N_15368);
or U16873 (N_16873,N_14906,N_14738);
or U16874 (N_16874,N_12751,N_13138);
nor U16875 (N_16875,N_13585,N_13144);
xnor U16876 (N_16876,N_14177,N_14968);
nand U16877 (N_16877,N_15323,N_14169);
nor U16878 (N_16878,N_14499,N_14450);
and U16879 (N_16879,N_13309,N_15490);
nand U16880 (N_16880,N_13033,N_15420);
nand U16881 (N_16881,N_13782,N_15488);
or U16882 (N_16882,N_14721,N_15606);
nand U16883 (N_16883,N_14665,N_14627);
and U16884 (N_16884,N_13145,N_14492);
nor U16885 (N_16885,N_13776,N_15160);
and U16886 (N_16886,N_14902,N_15150);
and U16887 (N_16887,N_13494,N_13060);
xnor U16888 (N_16888,N_13034,N_14010);
and U16889 (N_16889,N_15144,N_15568);
or U16890 (N_16890,N_15285,N_13527);
and U16891 (N_16891,N_12655,N_12518);
or U16892 (N_16892,N_14926,N_13547);
and U16893 (N_16893,N_15035,N_15149);
nand U16894 (N_16894,N_14903,N_14005);
xor U16895 (N_16895,N_12605,N_14467);
nand U16896 (N_16896,N_14022,N_13749);
nand U16897 (N_16897,N_14271,N_12934);
and U16898 (N_16898,N_14739,N_15374);
and U16899 (N_16899,N_15552,N_13235);
and U16900 (N_16900,N_14132,N_14432);
nand U16901 (N_16901,N_14532,N_14946);
nor U16902 (N_16902,N_15217,N_15455);
nor U16903 (N_16903,N_14602,N_13926);
or U16904 (N_16904,N_13865,N_14334);
nor U16905 (N_16905,N_12995,N_13384);
or U16906 (N_16906,N_15107,N_12795);
and U16907 (N_16907,N_12957,N_14609);
nor U16908 (N_16908,N_13601,N_14884);
or U16909 (N_16909,N_14755,N_15621);
or U16910 (N_16910,N_13390,N_15579);
nand U16911 (N_16911,N_15065,N_15489);
and U16912 (N_16912,N_14649,N_13277);
nor U16913 (N_16913,N_13728,N_14587);
and U16914 (N_16914,N_15589,N_13142);
nand U16915 (N_16915,N_14098,N_13927);
nor U16916 (N_16916,N_13668,N_14613);
nand U16917 (N_16917,N_13260,N_12592);
and U16918 (N_16918,N_13994,N_13013);
and U16919 (N_16919,N_14597,N_13655);
nand U16920 (N_16920,N_14982,N_12616);
nand U16921 (N_16921,N_13925,N_15101);
and U16922 (N_16922,N_12938,N_15319);
nand U16923 (N_16923,N_14948,N_12544);
and U16924 (N_16924,N_14445,N_13276);
nor U16925 (N_16925,N_13627,N_12661);
and U16926 (N_16926,N_15248,N_13555);
nand U16927 (N_16927,N_12552,N_14200);
and U16928 (N_16928,N_14493,N_12762);
nand U16929 (N_16929,N_12528,N_14194);
xor U16930 (N_16930,N_12732,N_12760);
or U16931 (N_16931,N_15360,N_14677);
nor U16932 (N_16932,N_14939,N_15388);
nand U16933 (N_16933,N_13259,N_15207);
nand U16934 (N_16934,N_13386,N_13389);
or U16935 (N_16935,N_14643,N_13422);
and U16936 (N_16936,N_13207,N_13978);
nor U16937 (N_16937,N_15188,N_15004);
or U16938 (N_16938,N_15197,N_13345);
nor U16939 (N_16939,N_14192,N_14543);
nor U16940 (N_16940,N_14592,N_13091);
nand U16941 (N_16941,N_12604,N_13310);
or U16942 (N_16942,N_12978,N_13798);
nor U16943 (N_16943,N_14583,N_13735);
nor U16944 (N_16944,N_13893,N_13973);
nand U16945 (N_16945,N_13077,N_13388);
or U16946 (N_16946,N_15202,N_13716);
nor U16947 (N_16947,N_15003,N_12755);
nor U16948 (N_16948,N_12791,N_14237);
and U16949 (N_16949,N_15565,N_15142);
nand U16950 (N_16950,N_12663,N_14614);
and U16951 (N_16951,N_13237,N_14572);
nor U16952 (N_16952,N_13600,N_15438);
and U16953 (N_16953,N_15206,N_14773);
nor U16954 (N_16954,N_13465,N_12710);
nand U16955 (N_16955,N_15382,N_13752);
nor U16956 (N_16956,N_13904,N_14226);
nand U16957 (N_16957,N_14190,N_14803);
nor U16958 (N_16958,N_14355,N_14949);
or U16959 (N_16959,N_12744,N_12548);
xor U16960 (N_16960,N_12805,N_12698);
and U16961 (N_16961,N_13271,N_14615);
or U16962 (N_16962,N_13512,N_14987);
nor U16963 (N_16963,N_13457,N_13416);
and U16964 (N_16964,N_14038,N_14480);
nand U16965 (N_16965,N_13489,N_14702);
nand U16966 (N_16966,N_13164,N_13470);
and U16967 (N_16967,N_14252,N_13966);
or U16968 (N_16968,N_13997,N_13955);
nor U16969 (N_16969,N_15032,N_12560);
nand U16970 (N_16970,N_13440,N_13094);
nor U16971 (N_16971,N_14737,N_12876);
or U16972 (N_16972,N_13682,N_14575);
nor U16973 (N_16973,N_12567,N_14534);
xnor U16974 (N_16974,N_13432,N_12680);
or U16975 (N_16975,N_12758,N_15453);
and U16976 (N_16976,N_15409,N_14834);
or U16977 (N_16977,N_14778,N_13647);
or U16978 (N_16978,N_15620,N_14438);
nand U16979 (N_16979,N_13707,N_12943);
and U16980 (N_16980,N_14449,N_14287);
xor U16981 (N_16981,N_13478,N_15210);
nor U16982 (N_16982,N_14681,N_14197);
xnor U16983 (N_16983,N_15619,N_14362);
xnor U16984 (N_16984,N_14927,N_13703);
nand U16985 (N_16985,N_14031,N_14800);
or U16986 (N_16986,N_14708,N_15241);
nand U16987 (N_16987,N_14827,N_13824);
or U16988 (N_16988,N_12576,N_14245);
or U16989 (N_16989,N_14727,N_14113);
nand U16990 (N_16990,N_14490,N_14876);
nand U16991 (N_16991,N_13263,N_13562);
nand U16992 (N_16992,N_12907,N_14418);
and U16993 (N_16993,N_12681,N_13852);
nor U16994 (N_16994,N_13954,N_15416);
or U16995 (N_16995,N_14248,N_14862);
or U16996 (N_16996,N_12529,N_12998);
or U16997 (N_16997,N_14726,N_14187);
nand U16998 (N_16998,N_15581,N_12683);
nand U16999 (N_16999,N_13553,N_15020);
nand U17000 (N_17000,N_13875,N_15090);
or U17001 (N_17001,N_13165,N_14656);
or U17002 (N_17002,N_14923,N_14201);
or U17003 (N_17003,N_14238,N_15317);
nand U17004 (N_17004,N_14992,N_14623);
or U17005 (N_17005,N_13261,N_15587);
or U17006 (N_17006,N_13029,N_12650);
and U17007 (N_17007,N_14724,N_13616);
nand U17008 (N_17008,N_13100,N_14765);
nand U17009 (N_17009,N_13475,N_12767);
and U17010 (N_17010,N_14745,N_12538);
nor U17011 (N_17011,N_14352,N_15190);
or U17012 (N_17012,N_15276,N_13109);
or U17013 (N_17013,N_13999,N_14136);
and U17014 (N_17014,N_13928,N_13734);
nor U17015 (N_17015,N_12963,N_14811);
and U17016 (N_17016,N_13105,N_13579);
nand U17017 (N_17017,N_14489,N_14835);
xor U17018 (N_17018,N_13970,N_13456);
xor U17019 (N_17019,N_14528,N_15411);
and U17020 (N_17020,N_14527,N_14446);
nand U17021 (N_17021,N_14911,N_14290);
nor U17022 (N_17022,N_14422,N_12810);
nand U17023 (N_17023,N_15045,N_14477);
nor U17024 (N_17024,N_13639,N_13740);
or U17025 (N_17025,N_14657,N_15412);
nand U17026 (N_17026,N_14779,N_15163);
or U17027 (N_17027,N_14280,N_13038);
nand U17028 (N_17028,N_14371,N_14890);
nand U17029 (N_17029,N_14185,N_13139);
or U17030 (N_17030,N_15306,N_14795);
xor U17031 (N_17031,N_14047,N_12555);
or U17032 (N_17032,N_14364,N_14484);
nand U17033 (N_17033,N_14730,N_15458);
xnor U17034 (N_17034,N_15072,N_14232);
and U17035 (N_17035,N_14054,N_14599);
or U17036 (N_17036,N_13932,N_14513);
xor U17037 (N_17037,N_12607,N_12766);
and U17038 (N_17038,N_12763,N_12857);
nor U17039 (N_17039,N_13941,N_15199);
or U17040 (N_17040,N_13841,N_13665);
and U17041 (N_17041,N_12910,N_14855);
or U17042 (N_17042,N_13193,N_13823);
xnor U17043 (N_17043,N_12556,N_13484);
nor U17044 (N_17044,N_13788,N_14781);
nor U17045 (N_17045,N_13586,N_15051);
or U17046 (N_17046,N_13998,N_14605);
nand U17047 (N_17047,N_12694,N_12936);
or U17048 (N_17048,N_13522,N_12530);
and U17049 (N_17049,N_15431,N_14652);
nand U17050 (N_17050,N_14653,N_13789);
and U17051 (N_17051,N_12553,N_15551);
and U17052 (N_17052,N_14184,N_13058);
or U17053 (N_17053,N_15095,N_14787);
nor U17054 (N_17054,N_15178,N_14292);
and U17055 (N_17055,N_15071,N_13762);
nand U17056 (N_17056,N_14752,N_13524);
nor U17057 (N_17057,N_15342,N_14635);
or U17058 (N_17058,N_14234,N_13301);
or U17059 (N_17059,N_13882,N_13043);
nor U17060 (N_17060,N_14451,N_13797);
xnor U17061 (N_17061,N_14845,N_14932);
nor U17062 (N_17062,N_13116,N_14744);
xnor U17063 (N_17063,N_13950,N_14267);
nor U17064 (N_17064,N_15467,N_13704);
xor U17065 (N_17065,N_12899,N_12863);
xnor U17066 (N_17066,N_14224,N_14413);
nor U17067 (N_17067,N_14979,N_14488);
nand U17068 (N_17068,N_13569,N_15542);
xnor U17069 (N_17069,N_12588,N_14565);
and U17070 (N_17070,N_14338,N_15618);
or U17071 (N_17071,N_13122,N_15398);
nand U17072 (N_17072,N_15010,N_13695);
nand U17073 (N_17073,N_14662,N_13080);
xnor U17074 (N_17074,N_14938,N_15108);
and U17075 (N_17075,N_14746,N_15291);
or U17076 (N_17076,N_14288,N_14314);
and U17077 (N_17077,N_15533,N_14507);
nor U17078 (N_17078,N_15502,N_12959);
or U17079 (N_17079,N_14873,N_12768);
nor U17080 (N_17080,N_14945,N_13101);
xnor U17081 (N_17081,N_12789,N_13546);
nand U17082 (N_17082,N_15514,N_14577);
and U17083 (N_17083,N_12628,N_14370);
or U17084 (N_17084,N_12519,N_14158);
nand U17085 (N_17085,N_14387,N_14304);
and U17086 (N_17086,N_12657,N_12608);
nor U17087 (N_17087,N_15439,N_13850);
or U17088 (N_17088,N_15464,N_14075);
or U17089 (N_17089,N_13690,N_13368);
nand U17090 (N_17090,N_15082,N_14256);
or U17091 (N_17091,N_14243,N_14318);
nor U17092 (N_17092,N_12602,N_13974);
xor U17093 (N_17093,N_14564,N_12986);
nor U17094 (N_17094,N_13842,N_14049);
and U17095 (N_17095,N_14067,N_13856);
nand U17096 (N_17096,N_13110,N_13943);
or U17097 (N_17097,N_13012,N_13658);
nand U17098 (N_17098,N_12956,N_15351);
nor U17099 (N_17099,N_15376,N_14888);
and U17100 (N_17100,N_12854,N_15265);
and U17101 (N_17101,N_12674,N_13759);
nor U17102 (N_17102,N_13330,N_12738);
and U17103 (N_17103,N_13153,N_15610);
or U17104 (N_17104,N_13183,N_13912);
or U17105 (N_17105,N_13002,N_14655);
nor U17106 (N_17106,N_13007,N_13468);
and U17107 (N_17107,N_14601,N_14315);
xnor U17108 (N_17108,N_14087,N_15450);
nand U17109 (N_17109,N_13267,N_14747);
nor U17110 (N_17110,N_13114,N_12718);
or U17111 (N_17111,N_13128,N_13343);
nor U17112 (N_17112,N_13318,N_14278);
xor U17113 (N_17113,N_15507,N_13134);
nor U17114 (N_17114,N_12725,N_13979);
nor U17115 (N_17115,N_15447,N_14805);
nor U17116 (N_17116,N_13873,N_13919);
nand U17117 (N_17117,N_15055,N_13864);
or U17118 (N_17118,N_14886,N_13157);
and U17119 (N_17119,N_13333,N_14829);
or U17120 (N_17120,N_15328,N_15394);
and U17121 (N_17121,N_12839,N_13891);
xor U17122 (N_17122,N_13709,N_12635);
nand U17123 (N_17123,N_14193,N_12856);
nor U17124 (N_17124,N_14166,N_14459);
nor U17125 (N_17125,N_15403,N_15194);
nor U17126 (N_17126,N_14858,N_15298);
and U17127 (N_17127,N_12690,N_12913);
and U17128 (N_17128,N_15147,N_12658);
or U17129 (N_17129,N_15520,N_13871);
nand U17130 (N_17130,N_15251,N_15611);
and U17131 (N_17131,N_15243,N_14916);
or U17132 (N_17132,N_13115,N_14947);
and U17133 (N_17133,N_13678,N_12786);
nand U17134 (N_17134,N_13680,N_15014);
nor U17135 (N_17135,N_14176,N_15211);
or U17136 (N_17136,N_14357,N_14452);
nand U17137 (N_17137,N_12841,N_13773);
nand U17138 (N_17138,N_12649,N_14435);
nor U17139 (N_17139,N_14096,N_12975);
xnor U17140 (N_17140,N_12892,N_15204);
nor U17141 (N_17141,N_12890,N_14799);
nand U17142 (N_17142,N_13408,N_12837);
nand U17143 (N_17143,N_13595,N_14297);
or U17144 (N_17144,N_13651,N_13539);
and U17145 (N_17145,N_15118,N_14321);
or U17146 (N_17146,N_14282,N_12775);
and U17147 (N_17147,N_13845,N_14937);
nand U17148 (N_17148,N_14915,N_15572);
nor U17149 (N_17149,N_15044,N_15214);
nor U17150 (N_17150,N_15262,N_12731);
or U17151 (N_17151,N_13557,N_12827);
or U17152 (N_17152,N_13326,N_14478);
and U17153 (N_17153,N_12771,N_13587);
or U17154 (N_17154,N_14222,N_14455);
or U17155 (N_17155,N_14768,N_13251);
xnor U17156 (N_17156,N_12672,N_14144);
nor U17157 (N_17157,N_14052,N_13429);
nor U17158 (N_17158,N_13541,N_12990);
nor U17159 (N_17159,N_14576,N_13132);
or U17160 (N_17160,N_14473,N_14885);
nor U17161 (N_17161,N_15022,N_12809);
or U17162 (N_17162,N_14223,N_13618);
nand U17163 (N_17163,N_14892,N_13685);
or U17164 (N_17164,N_13496,N_13062);
nand U17165 (N_17165,N_15088,N_13743);
nand U17166 (N_17166,N_15270,N_13779);
or U17167 (N_17167,N_13960,N_14209);
or U17168 (N_17168,N_14329,N_14776);
nand U17169 (N_17169,N_13186,N_14871);
xnor U17170 (N_17170,N_13756,N_15567);
nand U17171 (N_17171,N_12757,N_14093);
or U17172 (N_17172,N_15009,N_13477);
nor U17173 (N_17173,N_12949,N_15415);
nor U17174 (N_17174,N_13947,N_13821);
xor U17175 (N_17175,N_13278,N_12776);
nand U17176 (N_17176,N_15594,N_15237);
xnor U17177 (N_17177,N_14578,N_13515);
or U17178 (N_17178,N_14706,N_13895);
nand U17179 (N_17179,N_13792,N_12685);
or U17180 (N_17180,N_13611,N_14070);
and U17181 (N_17181,N_12842,N_15284);
or U17182 (N_17182,N_14872,N_14512);
and U17183 (N_17183,N_15601,N_13903);
and U17184 (N_17184,N_14430,N_13687);
nand U17185 (N_17185,N_15059,N_14207);
or U17186 (N_17186,N_13499,N_14469);
or U17187 (N_17187,N_14521,N_14372);
nor U17188 (N_17188,N_13400,N_12877);
or U17189 (N_17189,N_14447,N_13302);
or U17190 (N_17190,N_14660,N_13889);
or U17191 (N_17191,N_14407,N_14601);
and U17192 (N_17192,N_13885,N_13583);
and U17193 (N_17193,N_14725,N_14414);
and U17194 (N_17194,N_14056,N_12517);
xor U17195 (N_17195,N_12576,N_12717);
nand U17196 (N_17196,N_15445,N_14682);
or U17197 (N_17197,N_12536,N_15082);
nand U17198 (N_17198,N_13269,N_13353);
and U17199 (N_17199,N_13772,N_12950);
or U17200 (N_17200,N_15481,N_14268);
nand U17201 (N_17201,N_13875,N_14469);
or U17202 (N_17202,N_14913,N_15401);
nand U17203 (N_17203,N_13417,N_12790);
or U17204 (N_17204,N_13964,N_14646);
xnor U17205 (N_17205,N_15374,N_12609);
xor U17206 (N_17206,N_12934,N_15357);
nand U17207 (N_17207,N_13512,N_15064);
nand U17208 (N_17208,N_15520,N_15305);
nand U17209 (N_17209,N_13313,N_12516);
nor U17210 (N_17210,N_14505,N_14942);
or U17211 (N_17211,N_15264,N_12829);
and U17212 (N_17212,N_14206,N_14178);
nor U17213 (N_17213,N_14592,N_12750);
nand U17214 (N_17214,N_13600,N_14034);
and U17215 (N_17215,N_13868,N_14231);
nor U17216 (N_17216,N_12969,N_14054);
and U17217 (N_17217,N_13843,N_14314);
nor U17218 (N_17218,N_13594,N_13439);
or U17219 (N_17219,N_14003,N_13653);
and U17220 (N_17220,N_15003,N_14551);
and U17221 (N_17221,N_15039,N_13531);
and U17222 (N_17222,N_15539,N_14946);
xnor U17223 (N_17223,N_13093,N_12793);
nor U17224 (N_17224,N_12846,N_13480);
nor U17225 (N_17225,N_13483,N_13019);
nand U17226 (N_17226,N_14072,N_14435);
or U17227 (N_17227,N_15443,N_13135);
nand U17228 (N_17228,N_12796,N_15559);
or U17229 (N_17229,N_14187,N_13663);
xnor U17230 (N_17230,N_14316,N_14792);
nor U17231 (N_17231,N_13537,N_13500);
nand U17232 (N_17232,N_14692,N_12905);
and U17233 (N_17233,N_15295,N_13145);
xor U17234 (N_17234,N_13756,N_13840);
or U17235 (N_17235,N_14205,N_12876);
nor U17236 (N_17236,N_14066,N_13664);
or U17237 (N_17237,N_13519,N_12780);
nand U17238 (N_17238,N_14183,N_13942);
nor U17239 (N_17239,N_14676,N_15276);
or U17240 (N_17240,N_13554,N_15220);
and U17241 (N_17241,N_13680,N_14974);
and U17242 (N_17242,N_15025,N_15136);
or U17243 (N_17243,N_13683,N_13580);
or U17244 (N_17244,N_14242,N_14813);
and U17245 (N_17245,N_15520,N_14941);
and U17246 (N_17246,N_14087,N_14636);
nor U17247 (N_17247,N_12927,N_15318);
and U17248 (N_17248,N_15047,N_13561);
nand U17249 (N_17249,N_13452,N_13780);
nand U17250 (N_17250,N_14678,N_12674);
or U17251 (N_17251,N_14847,N_14892);
nor U17252 (N_17252,N_13492,N_13224);
nand U17253 (N_17253,N_14310,N_13361);
nor U17254 (N_17254,N_12934,N_13284);
nor U17255 (N_17255,N_13772,N_13103);
nand U17256 (N_17256,N_13583,N_14796);
or U17257 (N_17257,N_14583,N_15274);
nand U17258 (N_17258,N_12909,N_15031);
nand U17259 (N_17259,N_14403,N_13303);
nand U17260 (N_17260,N_14151,N_13693);
and U17261 (N_17261,N_15552,N_14003);
nand U17262 (N_17262,N_12705,N_14014);
nor U17263 (N_17263,N_15281,N_15442);
or U17264 (N_17264,N_15154,N_14211);
and U17265 (N_17265,N_14412,N_13835);
xor U17266 (N_17266,N_13034,N_15355);
and U17267 (N_17267,N_13011,N_15178);
nor U17268 (N_17268,N_14902,N_14633);
xnor U17269 (N_17269,N_13651,N_15541);
and U17270 (N_17270,N_14800,N_15424);
or U17271 (N_17271,N_14993,N_14419);
or U17272 (N_17272,N_12692,N_14165);
and U17273 (N_17273,N_13702,N_14660);
or U17274 (N_17274,N_13972,N_15110);
xor U17275 (N_17275,N_15031,N_14712);
or U17276 (N_17276,N_12604,N_14962);
nand U17277 (N_17277,N_15582,N_14331);
xor U17278 (N_17278,N_14577,N_13232);
and U17279 (N_17279,N_14121,N_12907);
nor U17280 (N_17280,N_12664,N_12559);
nand U17281 (N_17281,N_13610,N_13804);
nor U17282 (N_17282,N_15488,N_15096);
or U17283 (N_17283,N_12906,N_14964);
or U17284 (N_17284,N_15132,N_13042);
and U17285 (N_17285,N_13401,N_12920);
nor U17286 (N_17286,N_14746,N_12789);
and U17287 (N_17287,N_14680,N_15061);
or U17288 (N_17288,N_13306,N_12568);
nor U17289 (N_17289,N_14125,N_14665);
nand U17290 (N_17290,N_13151,N_12818);
or U17291 (N_17291,N_12719,N_13138);
nand U17292 (N_17292,N_12593,N_15125);
or U17293 (N_17293,N_12823,N_12759);
xnor U17294 (N_17294,N_13874,N_14935);
nor U17295 (N_17295,N_13134,N_15605);
nand U17296 (N_17296,N_13872,N_13942);
and U17297 (N_17297,N_15076,N_15227);
nor U17298 (N_17298,N_14667,N_15234);
or U17299 (N_17299,N_15044,N_12984);
nand U17300 (N_17300,N_14403,N_15472);
nand U17301 (N_17301,N_14488,N_14018);
and U17302 (N_17302,N_13635,N_12805);
or U17303 (N_17303,N_14507,N_13754);
and U17304 (N_17304,N_13040,N_13607);
and U17305 (N_17305,N_14250,N_13844);
or U17306 (N_17306,N_14388,N_13955);
and U17307 (N_17307,N_14306,N_14096);
and U17308 (N_17308,N_14537,N_14593);
nand U17309 (N_17309,N_13609,N_15169);
xor U17310 (N_17310,N_14033,N_14624);
nor U17311 (N_17311,N_14326,N_15560);
and U17312 (N_17312,N_12956,N_15315);
or U17313 (N_17313,N_15035,N_14496);
nor U17314 (N_17314,N_14908,N_13032);
nand U17315 (N_17315,N_14787,N_14783);
nor U17316 (N_17316,N_13149,N_14336);
nand U17317 (N_17317,N_15138,N_13739);
nand U17318 (N_17318,N_13873,N_14801);
nand U17319 (N_17319,N_13760,N_14883);
nor U17320 (N_17320,N_13859,N_13813);
nand U17321 (N_17321,N_15048,N_13568);
or U17322 (N_17322,N_14654,N_13203);
and U17323 (N_17323,N_14008,N_14572);
nand U17324 (N_17324,N_14696,N_14748);
or U17325 (N_17325,N_14077,N_14025);
or U17326 (N_17326,N_14257,N_12862);
nand U17327 (N_17327,N_14057,N_13705);
nor U17328 (N_17328,N_15314,N_13761);
or U17329 (N_17329,N_12551,N_14556);
nand U17330 (N_17330,N_15342,N_13132);
or U17331 (N_17331,N_12541,N_14746);
and U17332 (N_17332,N_14243,N_14476);
nand U17333 (N_17333,N_13721,N_15576);
nor U17334 (N_17334,N_13953,N_13409);
nor U17335 (N_17335,N_13417,N_13816);
or U17336 (N_17336,N_14533,N_14678);
nor U17337 (N_17337,N_15239,N_14749);
nor U17338 (N_17338,N_13172,N_15607);
and U17339 (N_17339,N_14555,N_14238);
xor U17340 (N_17340,N_13009,N_12510);
nand U17341 (N_17341,N_12540,N_15208);
nor U17342 (N_17342,N_15448,N_14532);
and U17343 (N_17343,N_13475,N_13946);
nand U17344 (N_17344,N_14769,N_15559);
and U17345 (N_17345,N_14194,N_13434);
or U17346 (N_17346,N_13211,N_12933);
and U17347 (N_17347,N_14725,N_13676);
nand U17348 (N_17348,N_13280,N_13975);
or U17349 (N_17349,N_12648,N_14704);
or U17350 (N_17350,N_13356,N_12752);
xnor U17351 (N_17351,N_12715,N_15001);
or U17352 (N_17352,N_14213,N_14292);
or U17353 (N_17353,N_15099,N_12856);
nor U17354 (N_17354,N_15202,N_13084);
nor U17355 (N_17355,N_13604,N_15620);
or U17356 (N_17356,N_14113,N_14500);
nand U17357 (N_17357,N_13390,N_13720);
nor U17358 (N_17358,N_14575,N_15069);
or U17359 (N_17359,N_14222,N_12683);
and U17360 (N_17360,N_15070,N_12774);
nor U17361 (N_17361,N_15279,N_14078);
nand U17362 (N_17362,N_12901,N_14702);
nor U17363 (N_17363,N_14331,N_12735);
or U17364 (N_17364,N_12587,N_14191);
and U17365 (N_17365,N_15607,N_14100);
or U17366 (N_17366,N_15575,N_13018);
xnor U17367 (N_17367,N_13155,N_14412);
or U17368 (N_17368,N_13808,N_15598);
nand U17369 (N_17369,N_15233,N_13359);
and U17370 (N_17370,N_15445,N_13403);
and U17371 (N_17371,N_14272,N_15304);
or U17372 (N_17372,N_13626,N_14903);
nor U17373 (N_17373,N_15541,N_14449);
nor U17374 (N_17374,N_12710,N_13186);
nor U17375 (N_17375,N_13426,N_15486);
nand U17376 (N_17376,N_14941,N_14224);
nand U17377 (N_17377,N_12590,N_14715);
xnor U17378 (N_17378,N_14922,N_15532);
or U17379 (N_17379,N_13166,N_14649);
nor U17380 (N_17380,N_12865,N_14931);
or U17381 (N_17381,N_14095,N_12579);
nor U17382 (N_17382,N_12777,N_12880);
xor U17383 (N_17383,N_13084,N_12537);
nand U17384 (N_17384,N_14771,N_13664);
nand U17385 (N_17385,N_14659,N_15070);
nand U17386 (N_17386,N_12907,N_15192);
and U17387 (N_17387,N_14201,N_12536);
xnor U17388 (N_17388,N_14262,N_15565);
nor U17389 (N_17389,N_13900,N_13917);
and U17390 (N_17390,N_14882,N_15031);
nand U17391 (N_17391,N_14584,N_13849);
nor U17392 (N_17392,N_12676,N_13141);
nand U17393 (N_17393,N_14587,N_13354);
and U17394 (N_17394,N_14431,N_14452);
and U17395 (N_17395,N_14468,N_12924);
nand U17396 (N_17396,N_12826,N_13397);
nor U17397 (N_17397,N_15156,N_14613);
and U17398 (N_17398,N_13703,N_14948);
and U17399 (N_17399,N_12671,N_13341);
xor U17400 (N_17400,N_13830,N_15466);
and U17401 (N_17401,N_13763,N_12664);
nor U17402 (N_17402,N_14270,N_13791);
xnor U17403 (N_17403,N_13430,N_13155);
nand U17404 (N_17404,N_13415,N_15331);
and U17405 (N_17405,N_13976,N_14162);
nand U17406 (N_17406,N_13414,N_15314);
xnor U17407 (N_17407,N_13429,N_14639);
nor U17408 (N_17408,N_13380,N_15601);
and U17409 (N_17409,N_14830,N_14583);
and U17410 (N_17410,N_13738,N_14981);
xnor U17411 (N_17411,N_14823,N_15038);
nand U17412 (N_17412,N_15312,N_14289);
xor U17413 (N_17413,N_12541,N_13799);
nand U17414 (N_17414,N_12748,N_12784);
and U17415 (N_17415,N_14112,N_12502);
nand U17416 (N_17416,N_14529,N_14651);
nor U17417 (N_17417,N_12590,N_13542);
nor U17418 (N_17418,N_14723,N_12806);
and U17419 (N_17419,N_14644,N_13375);
nand U17420 (N_17420,N_12741,N_13737);
nor U17421 (N_17421,N_12627,N_14057);
nor U17422 (N_17422,N_13136,N_15488);
nor U17423 (N_17423,N_15620,N_13339);
or U17424 (N_17424,N_14476,N_14606);
nand U17425 (N_17425,N_14406,N_14232);
xor U17426 (N_17426,N_12800,N_13486);
nor U17427 (N_17427,N_13102,N_14479);
nand U17428 (N_17428,N_12658,N_12686);
xor U17429 (N_17429,N_14970,N_13512);
nand U17430 (N_17430,N_13538,N_14883);
nand U17431 (N_17431,N_13752,N_14695);
or U17432 (N_17432,N_13383,N_13232);
and U17433 (N_17433,N_13026,N_14608);
or U17434 (N_17434,N_13952,N_14069);
or U17435 (N_17435,N_15216,N_13228);
and U17436 (N_17436,N_13571,N_15345);
or U17437 (N_17437,N_15187,N_13501);
nand U17438 (N_17438,N_12771,N_13894);
nand U17439 (N_17439,N_13892,N_13257);
or U17440 (N_17440,N_15340,N_14328);
and U17441 (N_17441,N_15271,N_14004);
xnor U17442 (N_17442,N_15451,N_13225);
nor U17443 (N_17443,N_14543,N_15256);
nand U17444 (N_17444,N_14555,N_13967);
nand U17445 (N_17445,N_13710,N_14406);
xnor U17446 (N_17446,N_14834,N_13203);
and U17447 (N_17447,N_12720,N_14353);
nor U17448 (N_17448,N_14761,N_14984);
nand U17449 (N_17449,N_14281,N_12620);
nor U17450 (N_17450,N_14608,N_14097);
and U17451 (N_17451,N_12524,N_14098);
or U17452 (N_17452,N_15554,N_13738);
xor U17453 (N_17453,N_15084,N_15342);
nand U17454 (N_17454,N_14680,N_13591);
nor U17455 (N_17455,N_13493,N_12983);
or U17456 (N_17456,N_12620,N_13486);
nor U17457 (N_17457,N_13893,N_15350);
nand U17458 (N_17458,N_14299,N_15450);
or U17459 (N_17459,N_15074,N_12838);
nor U17460 (N_17460,N_13497,N_15398);
nand U17461 (N_17461,N_14724,N_14139);
nand U17462 (N_17462,N_15007,N_14448);
and U17463 (N_17463,N_13888,N_15469);
nand U17464 (N_17464,N_12947,N_15472);
and U17465 (N_17465,N_14536,N_14945);
or U17466 (N_17466,N_12910,N_13201);
or U17467 (N_17467,N_13094,N_12821);
nor U17468 (N_17468,N_13798,N_15231);
nand U17469 (N_17469,N_13151,N_13806);
nor U17470 (N_17470,N_14629,N_15055);
nor U17471 (N_17471,N_13647,N_12850);
or U17472 (N_17472,N_14313,N_14038);
nand U17473 (N_17473,N_14885,N_15143);
nor U17474 (N_17474,N_14002,N_13233);
and U17475 (N_17475,N_15089,N_14949);
nand U17476 (N_17476,N_15215,N_13802);
and U17477 (N_17477,N_14406,N_13774);
or U17478 (N_17478,N_13901,N_13133);
nand U17479 (N_17479,N_14357,N_13418);
or U17480 (N_17480,N_15507,N_14732);
and U17481 (N_17481,N_14622,N_14075);
xor U17482 (N_17482,N_12673,N_15236);
nor U17483 (N_17483,N_14648,N_15242);
or U17484 (N_17484,N_14650,N_14782);
or U17485 (N_17485,N_13519,N_14829);
nor U17486 (N_17486,N_14036,N_14927);
nor U17487 (N_17487,N_12512,N_14012);
or U17488 (N_17488,N_13979,N_13925);
nand U17489 (N_17489,N_12834,N_13514);
nand U17490 (N_17490,N_14727,N_15340);
nand U17491 (N_17491,N_13456,N_12668);
nor U17492 (N_17492,N_13551,N_13533);
nand U17493 (N_17493,N_13049,N_13561);
nor U17494 (N_17494,N_12514,N_13911);
nand U17495 (N_17495,N_15232,N_12781);
and U17496 (N_17496,N_13989,N_12519);
nor U17497 (N_17497,N_13322,N_13946);
or U17498 (N_17498,N_13139,N_14786);
and U17499 (N_17499,N_14525,N_13577);
or U17500 (N_17500,N_14532,N_13911);
nand U17501 (N_17501,N_14651,N_15619);
nor U17502 (N_17502,N_13521,N_13441);
and U17503 (N_17503,N_13847,N_15108);
xnor U17504 (N_17504,N_15014,N_14169);
nor U17505 (N_17505,N_14704,N_15410);
and U17506 (N_17506,N_13466,N_14309);
and U17507 (N_17507,N_14913,N_14274);
nand U17508 (N_17508,N_13179,N_15083);
xnor U17509 (N_17509,N_12722,N_15343);
nor U17510 (N_17510,N_13853,N_13651);
nor U17511 (N_17511,N_13870,N_15029);
and U17512 (N_17512,N_15162,N_14370);
or U17513 (N_17513,N_12932,N_13389);
and U17514 (N_17514,N_14101,N_15256);
nand U17515 (N_17515,N_13014,N_14785);
nand U17516 (N_17516,N_13824,N_15391);
or U17517 (N_17517,N_14359,N_13712);
nand U17518 (N_17518,N_13753,N_15295);
nand U17519 (N_17519,N_15506,N_14936);
or U17520 (N_17520,N_14131,N_13152);
nand U17521 (N_17521,N_14728,N_13306);
nand U17522 (N_17522,N_13895,N_14814);
nand U17523 (N_17523,N_13049,N_15224);
nor U17524 (N_17524,N_14891,N_14404);
nor U17525 (N_17525,N_13355,N_13679);
nor U17526 (N_17526,N_14866,N_15093);
nor U17527 (N_17527,N_12549,N_13187);
and U17528 (N_17528,N_14323,N_13119);
xnor U17529 (N_17529,N_14166,N_13575);
nand U17530 (N_17530,N_15458,N_14867);
or U17531 (N_17531,N_15325,N_15316);
or U17532 (N_17532,N_13090,N_14793);
and U17533 (N_17533,N_13670,N_13621);
xor U17534 (N_17534,N_14512,N_12631);
or U17535 (N_17535,N_13965,N_12771);
nand U17536 (N_17536,N_15400,N_15143);
xnor U17537 (N_17537,N_14366,N_14977);
or U17538 (N_17538,N_13397,N_14751);
nand U17539 (N_17539,N_12831,N_13455);
nor U17540 (N_17540,N_13039,N_12505);
or U17541 (N_17541,N_13438,N_14184);
or U17542 (N_17542,N_15482,N_14919);
or U17543 (N_17543,N_14985,N_13060);
xor U17544 (N_17544,N_14047,N_13746);
xor U17545 (N_17545,N_15317,N_12975);
or U17546 (N_17546,N_14840,N_15352);
or U17547 (N_17547,N_15433,N_13971);
or U17548 (N_17548,N_13503,N_14209);
nor U17549 (N_17549,N_15111,N_13986);
nor U17550 (N_17550,N_14288,N_12744);
and U17551 (N_17551,N_14448,N_13404);
and U17552 (N_17552,N_15455,N_14044);
or U17553 (N_17553,N_15299,N_15571);
or U17554 (N_17554,N_13071,N_14046);
nand U17555 (N_17555,N_15181,N_13048);
nand U17556 (N_17556,N_15045,N_13082);
nand U17557 (N_17557,N_13410,N_13302);
and U17558 (N_17558,N_15317,N_15373);
nand U17559 (N_17559,N_14531,N_14649);
or U17560 (N_17560,N_15478,N_13502);
nor U17561 (N_17561,N_12636,N_15012);
or U17562 (N_17562,N_14992,N_15497);
nand U17563 (N_17563,N_13580,N_14593);
and U17564 (N_17564,N_13701,N_15103);
xnor U17565 (N_17565,N_14614,N_14513);
nor U17566 (N_17566,N_15170,N_13098);
xor U17567 (N_17567,N_12669,N_14013);
xnor U17568 (N_17568,N_13136,N_15422);
nor U17569 (N_17569,N_14472,N_14085);
nand U17570 (N_17570,N_15475,N_13271);
or U17571 (N_17571,N_14926,N_14897);
or U17572 (N_17572,N_15402,N_13172);
nor U17573 (N_17573,N_13673,N_12748);
nor U17574 (N_17574,N_14075,N_14104);
nand U17575 (N_17575,N_12632,N_14156);
and U17576 (N_17576,N_14637,N_13059);
nor U17577 (N_17577,N_15052,N_14770);
nand U17578 (N_17578,N_13254,N_12675);
nor U17579 (N_17579,N_13879,N_13141);
nand U17580 (N_17580,N_14101,N_13859);
xor U17581 (N_17581,N_13913,N_14170);
nand U17582 (N_17582,N_12787,N_15029);
nand U17583 (N_17583,N_15332,N_13260);
nor U17584 (N_17584,N_15017,N_12511);
xor U17585 (N_17585,N_15481,N_15137);
or U17586 (N_17586,N_12694,N_14443);
nand U17587 (N_17587,N_13359,N_12721);
and U17588 (N_17588,N_15374,N_14566);
and U17589 (N_17589,N_12902,N_14142);
nor U17590 (N_17590,N_12697,N_15145);
and U17591 (N_17591,N_12645,N_15266);
or U17592 (N_17592,N_14827,N_14545);
nand U17593 (N_17593,N_12575,N_13170);
nor U17594 (N_17594,N_15183,N_13709);
nor U17595 (N_17595,N_13480,N_15279);
xnor U17596 (N_17596,N_12619,N_14271);
nand U17597 (N_17597,N_13763,N_13010);
nor U17598 (N_17598,N_12744,N_14795);
nor U17599 (N_17599,N_14029,N_14591);
nor U17600 (N_17600,N_15155,N_13084);
nor U17601 (N_17601,N_13136,N_14955);
and U17602 (N_17602,N_15226,N_14593);
and U17603 (N_17603,N_14924,N_14339);
and U17604 (N_17604,N_12721,N_14248);
nand U17605 (N_17605,N_13216,N_14163);
and U17606 (N_17606,N_15623,N_15394);
and U17607 (N_17607,N_15418,N_12995);
nor U17608 (N_17608,N_15270,N_14377);
xnor U17609 (N_17609,N_15361,N_12883);
xnor U17610 (N_17610,N_14938,N_15077);
nand U17611 (N_17611,N_14795,N_13640);
and U17612 (N_17612,N_14759,N_13191);
and U17613 (N_17613,N_13945,N_13525);
xor U17614 (N_17614,N_15499,N_13926);
nor U17615 (N_17615,N_13773,N_14079);
or U17616 (N_17616,N_13417,N_15082);
nor U17617 (N_17617,N_13392,N_15463);
nor U17618 (N_17618,N_14839,N_14181);
xnor U17619 (N_17619,N_14130,N_12502);
nand U17620 (N_17620,N_12782,N_13544);
and U17621 (N_17621,N_12922,N_12974);
xnor U17622 (N_17622,N_15109,N_14008);
and U17623 (N_17623,N_15477,N_15362);
xor U17624 (N_17624,N_14052,N_15003);
and U17625 (N_17625,N_13808,N_13328);
nor U17626 (N_17626,N_12868,N_14935);
nand U17627 (N_17627,N_15141,N_15226);
or U17628 (N_17628,N_14490,N_12817);
and U17629 (N_17629,N_15340,N_12567);
or U17630 (N_17630,N_15362,N_14197);
or U17631 (N_17631,N_13096,N_13766);
nand U17632 (N_17632,N_12505,N_14951);
or U17633 (N_17633,N_13275,N_13484);
or U17634 (N_17634,N_14954,N_13363);
nand U17635 (N_17635,N_14632,N_15610);
nand U17636 (N_17636,N_12629,N_14579);
and U17637 (N_17637,N_12802,N_14317);
and U17638 (N_17638,N_15062,N_14455);
and U17639 (N_17639,N_14310,N_13697);
or U17640 (N_17640,N_13998,N_13165);
xor U17641 (N_17641,N_13944,N_15037);
and U17642 (N_17642,N_15117,N_13193);
nand U17643 (N_17643,N_14235,N_12966);
and U17644 (N_17644,N_13298,N_12881);
nor U17645 (N_17645,N_13073,N_15545);
nor U17646 (N_17646,N_14999,N_13661);
and U17647 (N_17647,N_15120,N_15177);
nand U17648 (N_17648,N_15153,N_13826);
and U17649 (N_17649,N_14660,N_14574);
nor U17650 (N_17650,N_12931,N_13945);
xor U17651 (N_17651,N_13413,N_14431);
or U17652 (N_17652,N_15420,N_14454);
and U17653 (N_17653,N_13374,N_12919);
xnor U17654 (N_17654,N_12986,N_14473);
nor U17655 (N_17655,N_15181,N_13142);
nand U17656 (N_17656,N_13810,N_13048);
and U17657 (N_17657,N_14923,N_12683);
nor U17658 (N_17658,N_13491,N_14359);
or U17659 (N_17659,N_12660,N_13689);
nand U17660 (N_17660,N_13652,N_14945);
nor U17661 (N_17661,N_14104,N_12588);
nor U17662 (N_17662,N_14902,N_14244);
xnor U17663 (N_17663,N_13121,N_15489);
and U17664 (N_17664,N_15317,N_13526);
and U17665 (N_17665,N_12971,N_15259);
and U17666 (N_17666,N_13673,N_13248);
or U17667 (N_17667,N_12983,N_13041);
nor U17668 (N_17668,N_13076,N_12957);
or U17669 (N_17669,N_14085,N_13577);
nand U17670 (N_17670,N_14502,N_13375);
nand U17671 (N_17671,N_13986,N_14489);
or U17672 (N_17672,N_13042,N_13122);
xor U17673 (N_17673,N_13869,N_12514);
or U17674 (N_17674,N_14173,N_13923);
nor U17675 (N_17675,N_13033,N_15614);
or U17676 (N_17676,N_13532,N_13422);
and U17677 (N_17677,N_15326,N_12804);
xor U17678 (N_17678,N_12794,N_13330);
nand U17679 (N_17679,N_13518,N_15030);
or U17680 (N_17680,N_14849,N_15260);
nand U17681 (N_17681,N_14800,N_14313);
nand U17682 (N_17682,N_13187,N_13523);
or U17683 (N_17683,N_13534,N_14135);
nand U17684 (N_17684,N_14740,N_13866);
and U17685 (N_17685,N_15287,N_14404);
nor U17686 (N_17686,N_14077,N_14744);
or U17687 (N_17687,N_14837,N_14318);
nand U17688 (N_17688,N_15408,N_15538);
xor U17689 (N_17689,N_14935,N_14596);
nor U17690 (N_17690,N_12635,N_13536);
or U17691 (N_17691,N_14788,N_15508);
nor U17692 (N_17692,N_14260,N_14501);
and U17693 (N_17693,N_12928,N_15196);
xor U17694 (N_17694,N_12645,N_12797);
nor U17695 (N_17695,N_13557,N_13724);
nor U17696 (N_17696,N_13157,N_15257);
and U17697 (N_17697,N_15105,N_14201);
and U17698 (N_17698,N_12745,N_15287);
nor U17699 (N_17699,N_14220,N_13817);
nand U17700 (N_17700,N_12864,N_13594);
xor U17701 (N_17701,N_15211,N_15118);
or U17702 (N_17702,N_14110,N_15423);
and U17703 (N_17703,N_14412,N_13735);
nor U17704 (N_17704,N_14740,N_14896);
xor U17705 (N_17705,N_14944,N_12792);
and U17706 (N_17706,N_12988,N_13372);
nand U17707 (N_17707,N_13037,N_14082);
nor U17708 (N_17708,N_14254,N_13477);
or U17709 (N_17709,N_13076,N_13465);
nand U17710 (N_17710,N_12996,N_12620);
nor U17711 (N_17711,N_14855,N_14484);
and U17712 (N_17712,N_13514,N_15471);
or U17713 (N_17713,N_13256,N_14525);
and U17714 (N_17714,N_13515,N_14299);
nor U17715 (N_17715,N_14730,N_13993);
nor U17716 (N_17716,N_15082,N_15436);
xnor U17717 (N_17717,N_14661,N_14671);
and U17718 (N_17718,N_14321,N_13810);
nand U17719 (N_17719,N_14046,N_15390);
or U17720 (N_17720,N_14893,N_14548);
and U17721 (N_17721,N_14112,N_14094);
nand U17722 (N_17722,N_13553,N_13693);
and U17723 (N_17723,N_13343,N_13377);
nor U17724 (N_17724,N_14405,N_15172);
nand U17725 (N_17725,N_14104,N_15249);
and U17726 (N_17726,N_14112,N_14147);
or U17727 (N_17727,N_15336,N_15083);
nor U17728 (N_17728,N_14926,N_13119);
or U17729 (N_17729,N_14962,N_15163);
nand U17730 (N_17730,N_13306,N_13369);
and U17731 (N_17731,N_13096,N_12696);
and U17732 (N_17732,N_15586,N_14333);
or U17733 (N_17733,N_15363,N_12929);
nand U17734 (N_17734,N_13368,N_14016);
xor U17735 (N_17735,N_12697,N_14715);
nor U17736 (N_17736,N_13059,N_13026);
and U17737 (N_17737,N_12561,N_15209);
nand U17738 (N_17738,N_13528,N_14146);
or U17739 (N_17739,N_15270,N_15505);
nand U17740 (N_17740,N_14725,N_15364);
or U17741 (N_17741,N_15360,N_12635);
and U17742 (N_17742,N_15539,N_13789);
and U17743 (N_17743,N_14597,N_14167);
nand U17744 (N_17744,N_14238,N_14247);
or U17745 (N_17745,N_14203,N_13324);
xor U17746 (N_17746,N_15369,N_13118);
nand U17747 (N_17747,N_13137,N_13015);
and U17748 (N_17748,N_14448,N_15170);
or U17749 (N_17749,N_14336,N_14158);
or U17750 (N_17750,N_13041,N_14065);
or U17751 (N_17751,N_15336,N_13914);
nor U17752 (N_17752,N_13131,N_15169);
nor U17753 (N_17753,N_13242,N_13455);
and U17754 (N_17754,N_13306,N_14945);
and U17755 (N_17755,N_15163,N_12694);
and U17756 (N_17756,N_14624,N_13789);
nand U17757 (N_17757,N_13697,N_13482);
or U17758 (N_17758,N_15343,N_14359);
and U17759 (N_17759,N_12868,N_13191);
nand U17760 (N_17760,N_14997,N_14449);
nor U17761 (N_17761,N_15301,N_13353);
and U17762 (N_17762,N_13329,N_15519);
or U17763 (N_17763,N_14899,N_13599);
nand U17764 (N_17764,N_13771,N_13557);
nor U17765 (N_17765,N_14500,N_14670);
or U17766 (N_17766,N_13712,N_14174);
nand U17767 (N_17767,N_12972,N_13699);
or U17768 (N_17768,N_15420,N_14276);
nor U17769 (N_17769,N_13776,N_13793);
and U17770 (N_17770,N_15384,N_14730);
and U17771 (N_17771,N_14325,N_13949);
and U17772 (N_17772,N_14682,N_15382);
nand U17773 (N_17773,N_14213,N_13685);
nand U17774 (N_17774,N_12733,N_13507);
nand U17775 (N_17775,N_14865,N_15226);
and U17776 (N_17776,N_12679,N_15387);
and U17777 (N_17777,N_15196,N_15353);
nand U17778 (N_17778,N_14500,N_14910);
nand U17779 (N_17779,N_14997,N_15236);
nor U17780 (N_17780,N_13530,N_13852);
xor U17781 (N_17781,N_12687,N_14044);
or U17782 (N_17782,N_14497,N_12588);
xor U17783 (N_17783,N_14985,N_13357);
xor U17784 (N_17784,N_14723,N_12668);
nand U17785 (N_17785,N_14279,N_14909);
nand U17786 (N_17786,N_14694,N_12842);
nor U17787 (N_17787,N_14858,N_12547);
or U17788 (N_17788,N_15074,N_15310);
nor U17789 (N_17789,N_14371,N_14025);
or U17790 (N_17790,N_12676,N_14708);
and U17791 (N_17791,N_15604,N_15522);
or U17792 (N_17792,N_15482,N_13591);
nor U17793 (N_17793,N_12788,N_12637);
nor U17794 (N_17794,N_13817,N_14032);
nand U17795 (N_17795,N_13409,N_13864);
xnor U17796 (N_17796,N_12910,N_15134);
and U17797 (N_17797,N_15251,N_14804);
and U17798 (N_17798,N_13063,N_13781);
or U17799 (N_17799,N_14433,N_13937);
nand U17800 (N_17800,N_14696,N_13241);
xnor U17801 (N_17801,N_15178,N_15209);
nor U17802 (N_17802,N_13789,N_14687);
nor U17803 (N_17803,N_14354,N_14513);
and U17804 (N_17804,N_15368,N_12899);
nand U17805 (N_17805,N_13601,N_15413);
xnor U17806 (N_17806,N_13151,N_15113);
nor U17807 (N_17807,N_15017,N_12707);
and U17808 (N_17808,N_13929,N_14825);
nor U17809 (N_17809,N_12811,N_14853);
xor U17810 (N_17810,N_14541,N_13105);
or U17811 (N_17811,N_15354,N_14331);
nand U17812 (N_17812,N_12564,N_15552);
or U17813 (N_17813,N_15609,N_13643);
nor U17814 (N_17814,N_14489,N_13410);
nand U17815 (N_17815,N_13082,N_15248);
or U17816 (N_17816,N_13899,N_12873);
xor U17817 (N_17817,N_13486,N_12862);
nor U17818 (N_17818,N_14846,N_15203);
and U17819 (N_17819,N_14284,N_13682);
nor U17820 (N_17820,N_12539,N_13485);
nand U17821 (N_17821,N_13906,N_13902);
nand U17822 (N_17822,N_14784,N_14577);
nor U17823 (N_17823,N_15217,N_13513);
and U17824 (N_17824,N_13778,N_13873);
nand U17825 (N_17825,N_14833,N_12941);
nand U17826 (N_17826,N_14947,N_14726);
xnor U17827 (N_17827,N_15216,N_14583);
nand U17828 (N_17828,N_13832,N_13645);
nand U17829 (N_17829,N_13339,N_14818);
nor U17830 (N_17830,N_13823,N_14242);
nand U17831 (N_17831,N_12965,N_12801);
nand U17832 (N_17832,N_13056,N_12665);
or U17833 (N_17833,N_13346,N_12835);
and U17834 (N_17834,N_15230,N_14236);
nor U17835 (N_17835,N_14760,N_13351);
nand U17836 (N_17836,N_13615,N_13611);
nand U17837 (N_17837,N_12983,N_14721);
or U17838 (N_17838,N_12841,N_14177);
and U17839 (N_17839,N_15196,N_13837);
and U17840 (N_17840,N_13152,N_14862);
and U17841 (N_17841,N_12909,N_15610);
nor U17842 (N_17842,N_15007,N_14560);
and U17843 (N_17843,N_14130,N_14936);
or U17844 (N_17844,N_13353,N_15437);
nor U17845 (N_17845,N_15114,N_13314);
nand U17846 (N_17846,N_13453,N_14186);
and U17847 (N_17847,N_12592,N_13744);
and U17848 (N_17848,N_12707,N_13265);
or U17849 (N_17849,N_15371,N_15005);
nor U17850 (N_17850,N_12526,N_15005);
or U17851 (N_17851,N_13593,N_13895);
or U17852 (N_17852,N_12882,N_13349);
or U17853 (N_17853,N_13072,N_15365);
xor U17854 (N_17854,N_13297,N_15225);
nand U17855 (N_17855,N_14749,N_15090);
and U17856 (N_17856,N_12607,N_12804);
or U17857 (N_17857,N_13977,N_14276);
nor U17858 (N_17858,N_15492,N_13349);
nor U17859 (N_17859,N_15544,N_15451);
nand U17860 (N_17860,N_14655,N_15395);
nand U17861 (N_17861,N_12932,N_15295);
nand U17862 (N_17862,N_13651,N_13357);
nand U17863 (N_17863,N_14636,N_13984);
or U17864 (N_17864,N_14152,N_14001);
and U17865 (N_17865,N_13585,N_13982);
nor U17866 (N_17866,N_12504,N_13773);
nor U17867 (N_17867,N_12547,N_14332);
xnor U17868 (N_17868,N_13455,N_14664);
nand U17869 (N_17869,N_14809,N_12658);
nor U17870 (N_17870,N_13821,N_14193);
nor U17871 (N_17871,N_15060,N_14632);
nor U17872 (N_17872,N_15035,N_14314);
nand U17873 (N_17873,N_14127,N_15495);
nand U17874 (N_17874,N_14448,N_15612);
nand U17875 (N_17875,N_12818,N_13873);
nand U17876 (N_17876,N_13023,N_14251);
nor U17877 (N_17877,N_13503,N_13604);
and U17878 (N_17878,N_12595,N_13381);
or U17879 (N_17879,N_13310,N_12943);
nand U17880 (N_17880,N_13380,N_12682);
nand U17881 (N_17881,N_14906,N_14383);
nor U17882 (N_17882,N_12542,N_14829);
nor U17883 (N_17883,N_12850,N_12713);
nand U17884 (N_17884,N_13902,N_13414);
and U17885 (N_17885,N_13830,N_12678);
nand U17886 (N_17886,N_14811,N_13471);
nor U17887 (N_17887,N_15071,N_14401);
or U17888 (N_17888,N_14583,N_15089);
and U17889 (N_17889,N_13416,N_13621);
nor U17890 (N_17890,N_15459,N_13750);
nand U17891 (N_17891,N_15040,N_13384);
and U17892 (N_17892,N_14799,N_14402);
xnor U17893 (N_17893,N_13826,N_15586);
nor U17894 (N_17894,N_13758,N_15291);
or U17895 (N_17895,N_12890,N_15002);
or U17896 (N_17896,N_12842,N_12751);
nor U17897 (N_17897,N_13654,N_12604);
nand U17898 (N_17898,N_13469,N_12705);
and U17899 (N_17899,N_13947,N_13238);
xor U17900 (N_17900,N_13812,N_12753);
nor U17901 (N_17901,N_13658,N_14428);
nor U17902 (N_17902,N_13515,N_12904);
nand U17903 (N_17903,N_13805,N_15455);
or U17904 (N_17904,N_15587,N_15233);
xor U17905 (N_17905,N_14895,N_13300);
and U17906 (N_17906,N_15466,N_15121);
xor U17907 (N_17907,N_14168,N_13302);
nor U17908 (N_17908,N_15464,N_12531);
nand U17909 (N_17909,N_14438,N_14303);
and U17910 (N_17910,N_15602,N_14250);
and U17911 (N_17911,N_13259,N_13068);
or U17912 (N_17912,N_14983,N_12602);
or U17913 (N_17913,N_14774,N_12978);
nand U17914 (N_17914,N_13364,N_14357);
and U17915 (N_17915,N_12686,N_14887);
nor U17916 (N_17916,N_15210,N_14987);
xnor U17917 (N_17917,N_12696,N_13658);
and U17918 (N_17918,N_15290,N_15451);
nand U17919 (N_17919,N_13724,N_13307);
nor U17920 (N_17920,N_13357,N_12841);
xor U17921 (N_17921,N_14022,N_12796);
xor U17922 (N_17922,N_14523,N_14748);
xor U17923 (N_17923,N_15013,N_12916);
and U17924 (N_17924,N_14341,N_14916);
or U17925 (N_17925,N_14808,N_13034);
nor U17926 (N_17926,N_14328,N_14448);
nor U17927 (N_17927,N_13498,N_14787);
nor U17928 (N_17928,N_13497,N_12538);
nor U17929 (N_17929,N_14136,N_13282);
and U17930 (N_17930,N_13273,N_13760);
nor U17931 (N_17931,N_15228,N_14596);
or U17932 (N_17932,N_12704,N_12854);
and U17933 (N_17933,N_15457,N_12868);
nand U17934 (N_17934,N_14746,N_15459);
nor U17935 (N_17935,N_13766,N_14634);
or U17936 (N_17936,N_14945,N_14446);
or U17937 (N_17937,N_15500,N_13876);
or U17938 (N_17938,N_12501,N_14197);
nor U17939 (N_17939,N_15477,N_14662);
or U17940 (N_17940,N_12731,N_15252);
or U17941 (N_17941,N_15201,N_13124);
and U17942 (N_17942,N_15059,N_14151);
or U17943 (N_17943,N_13479,N_12552);
xnor U17944 (N_17944,N_14705,N_14181);
and U17945 (N_17945,N_12575,N_15368);
nand U17946 (N_17946,N_12607,N_14139);
or U17947 (N_17947,N_13048,N_14556);
or U17948 (N_17948,N_15233,N_14227);
and U17949 (N_17949,N_14249,N_14894);
nand U17950 (N_17950,N_14036,N_14274);
nand U17951 (N_17951,N_15296,N_14092);
and U17952 (N_17952,N_13101,N_15094);
nor U17953 (N_17953,N_14606,N_15470);
nor U17954 (N_17954,N_14715,N_13399);
nor U17955 (N_17955,N_14130,N_12926);
nor U17956 (N_17956,N_12620,N_15103);
xnor U17957 (N_17957,N_13226,N_13758);
xnor U17958 (N_17958,N_13835,N_13712);
and U17959 (N_17959,N_12526,N_13049);
nor U17960 (N_17960,N_13327,N_15615);
and U17961 (N_17961,N_13972,N_13054);
and U17962 (N_17962,N_14809,N_12874);
or U17963 (N_17963,N_15540,N_12804);
nor U17964 (N_17964,N_13214,N_14801);
nor U17965 (N_17965,N_13268,N_13853);
xor U17966 (N_17966,N_14845,N_13170);
and U17967 (N_17967,N_14788,N_13746);
xor U17968 (N_17968,N_13282,N_14259);
xor U17969 (N_17969,N_13014,N_14871);
nand U17970 (N_17970,N_13748,N_13853);
nor U17971 (N_17971,N_15142,N_13124);
xnor U17972 (N_17972,N_15321,N_14397);
and U17973 (N_17973,N_14540,N_14177);
nand U17974 (N_17974,N_13415,N_13917);
or U17975 (N_17975,N_13058,N_14792);
and U17976 (N_17976,N_14509,N_12921);
nand U17977 (N_17977,N_14230,N_14735);
nor U17978 (N_17978,N_14967,N_12871);
nor U17979 (N_17979,N_13737,N_12835);
nand U17980 (N_17980,N_13987,N_12713);
nor U17981 (N_17981,N_14687,N_12947);
xnor U17982 (N_17982,N_14649,N_12838);
nand U17983 (N_17983,N_14503,N_13066);
and U17984 (N_17984,N_13753,N_13149);
and U17985 (N_17985,N_14413,N_15510);
nor U17986 (N_17986,N_12910,N_12998);
and U17987 (N_17987,N_13398,N_13987);
nor U17988 (N_17988,N_15365,N_14399);
and U17989 (N_17989,N_14276,N_12780);
nand U17990 (N_17990,N_14179,N_15560);
or U17991 (N_17991,N_13626,N_13229);
or U17992 (N_17992,N_13481,N_15427);
and U17993 (N_17993,N_14767,N_14371);
nor U17994 (N_17994,N_13847,N_15123);
or U17995 (N_17995,N_14458,N_15423);
xnor U17996 (N_17996,N_14020,N_13078);
xnor U17997 (N_17997,N_13588,N_14416);
and U17998 (N_17998,N_14503,N_14735);
or U17999 (N_17999,N_14588,N_14886);
and U18000 (N_18000,N_12852,N_13282);
and U18001 (N_18001,N_14185,N_13741);
xnor U18002 (N_18002,N_12870,N_14453);
or U18003 (N_18003,N_12523,N_12601);
nor U18004 (N_18004,N_12788,N_13491);
xnor U18005 (N_18005,N_13366,N_14657);
xor U18006 (N_18006,N_13919,N_15146);
nor U18007 (N_18007,N_14675,N_15029);
nor U18008 (N_18008,N_13772,N_12646);
nand U18009 (N_18009,N_14451,N_13907);
and U18010 (N_18010,N_14552,N_14443);
and U18011 (N_18011,N_13747,N_15217);
nor U18012 (N_18012,N_13844,N_13894);
nand U18013 (N_18013,N_14112,N_13730);
and U18014 (N_18014,N_13385,N_14464);
nand U18015 (N_18015,N_13617,N_12851);
and U18016 (N_18016,N_12616,N_12858);
or U18017 (N_18017,N_14886,N_13982);
or U18018 (N_18018,N_14496,N_14644);
nand U18019 (N_18019,N_14616,N_15158);
nand U18020 (N_18020,N_12859,N_15255);
nand U18021 (N_18021,N_15581,N_14936);
and U18022 (N_18022,N_15093,N_13793);
xnor U18023 (N_18023,N_15182,N_15041);
nor U18024 (N_18024,N_13499,N_14401);
or U18025 (N_18025,N_12788,N_13198);
nand U18026 (N_18026,N_14007,N_13595);
xor U18027 (N_18027,N_13778,N_14701);
nand U18028 (N_18028,N_13070,N_15100);
nand U18029 (N_18029,N_15171,N_13488);
nand U18030 (N_18030,N_14634,N_15104);
nor U18031 (N_18031,N_15239,N_14157);
nor U18032 (N_18032,N_13744,N_14099);
xor U18033 (N_18033,N_13274,N_13799);
nand U18034 (N_18034,N_14481,N_13304);
nor U18035 (N_18035,N_13591,N_13838);
nor U18036 (N_18036,N_13276,N_13280);
and U18037 (N_18037,N_15388,N_14996);
and U18038 (N_18038,N_15137,N_13293);
or U18039 (N_18039,N_14771,N_14190);
and U18040 (N_18040,N_15039,N_14768);
or U18041 (N_18041,N_12940,N_13308);
nor U18042 (N_18042,N_14176,N_13911);
or U18043 (N_18043,N_14378,N_13968);
and U18044 (N_18044,N_12596,N_13536);
and U18045 (N_18045,N_13137,N_15405);
nand U18046 (N_18046,N_14428,N_13000);
xnor U18047 (N_18047,N_14813,N_12857);
and U18048 (N_18048,N_15214,N_15300);
or U18049 (N_18049,N_14555,N_15403);
nor U18050 (N_18050,N_15051,N_14139);
xor U18051 (N_18051,N_14335,N_14686);
and U18052 (N_18052,N_15209,N_15391);
and U18053 (N_18053,N_13265,N_13609);
nor U18054 (N_18054,N_14486,N_14149);
and U18055 (N_18055,N_13104,N_15109);
nor U18056 (N_18056,N_13719,N_13481);
or U18057 (N_18057,N_13005,N_13503);
nand U18058 (N_18058,N_13203,N_13866);
nor U18059 (N_18059,N_12681,N_13920);
or U18060 (N_18060,N_13206,N_13080);
and U18061 (N_18061,N_14917,N_13492);
or U18062 (N_18062,N_13356,N_14231);
xor U18063 (N_18063,N_13157,N_15405);
nor U18064 (N_18064,N_15478,N_13518);
nor U18065 (N_18065,N_12870,N_13116);
nor U18066 (N_18066,N_12950,N_13040);
nand U18067 (N_18067,N_13040,N_13860);
nor U18068 (N_18068,N_15550,N_13282);
nand U18069 (N_18069,N_15077,N_14669);
and U18070 (N_18070,N_15586,N_14526);
or U18071 (N_18071,N_14115,N_14124);
or U18072 (N_18072,N_15030,N_12549);
nand U18073 (N_18073,N_14300,N_12977);
and U18074 (N_18074,N_12904,N_12842);
or U18075 (N_18075,N_13944,N_12743);
and U18076 (N_18076,N_12974,N_12952);
nor U18077 (N_18077,N_12887,N_14749);
and U18078 (N_18078,N_14289,N_15053);
nand U18079 (N_18079,N_14596,N_13710);
xnor U18080 (N_18080,N_15316,N_13008);
and U18081 (N_18081,N_12658,N_12652);
and U18082 (N_18082,N_13284,N_13326);
nand U18083 (N_18083,N_12780,N_15473);
nor U18084 (N_18084,N_14773,N_13814);
nor U18085 (N_18085,N_12874,N_14095);
and U18086 (N_18086,N_14783,N_14212);
xor U18087 (N_18087,N_12754,N_12888);
nor U18088 (N_18088,N_13597,N_13807);
nor U18089 (N_18089,N_15268,N_14635);
or U18090 (N_18090,N_14282,N_14464);
nor U18091 (N_18091,N_13165,N_12914);
and U18092 (N_18092,N_14518,N_13160);
nand U18093 (N_18093,N_14301,N_13230);
nand U18094 (N_18094,N_14810,N_15427);
and U18095 (N_18095,N_15165,N_12524);
and U18096 (N_18096,N_13689,N_12627);
nand U18097 (N_18097,N_15126,N_13398);
and U18098 (N_18098,N_15195,N_14810);
nor U18099 (N_18099,N_13640,N_15179);
or U18100 (N_18100,N_12685,N_14648);
nor U18101 (N_18101,N_14762,N_12887);
nor U18102 (N_18102,N_14555,N_13912);
nor U18103 (N_18103,N_14935,N_14475);
nand U18104 (N_18104,N_13461,N_13978);
or U18105 (N_18105,N_14724,N_14741);
nor U18106 (N_18106,N_14044,N_13026);
nor U18107 (N_18107,N_15599,N_13220);
nand U18108 (N_18108,N_13920,N_14165);
and U18109 (N_18109,N_14112,N_13219);
nor U18110 (N_18110,N_13161,N_13001);
or U18111 (N_18111,N_14250,N_15081);
and U18112 (N_18112,N_12603,N_13846);
nand U18113 (N_18113,N_14521,N_12658);
and U18114 (N_18114,N_14421,N_15077);
nand U18115 (N_18115,N_13356,N_14250);
nor U18116 (N_18116,N_14147,N_14133);
nor U18117 (N_18117,N_13504,N_14215);
or U18118 (N_18118,N_14483,N_15598);
nor U18119 (N_18119,N_14944,N_14624);
or U18120 (N_18120,N_12918,N_13233);
nand U18121 (N_18121,N_14908,N_13006);
nor U18122 (N_18122,N_13007,N_13919);
nor U18123 (N_18123,N_12919,N_15275);
or U18124 (N_18124,N_15223,N_12623);
nor U18125 (N_18125,N_13640,N_12653);
or U18126 (N_18126,N_14281,N_14499);
and U18127 (N_18127,N_13710,N_13379);
xor U18128 (N_18128,N_14131,N_13074);
nor U18129 (N_18129,N_13454,N_12957);
nand U18130 (N_18130,N_14825,N_15038);
or U18131 (N_18131,N_14378,N_12948);
and U18132 (N_18132,N_14137,N_12625);
or U18133 (N_18133,N_12691,N_14659);
xor U18134 (N_18134,N_15289,N_13696);
nand U18135 (N_18135,N_14561,N_14070);
nor U18136 (N_18136,N_13839,N_13827);
xnor U18137 (N_18137,N_13848,N_12784);
xor U18138 (N_18138,N_13363,N_13494);
nor U18139 (N_18139,N_14224,N_13236);
xnor U18140 (N_18140,N_13518,N_13912);
nor U18141 (N_18141,N_13286,N_14979);
or U18142 (N_18142,N_15480,N_12937);
and U18143 (N_18143,N_15458,N_15048);
or U18144 (N_18144,N_13604,N_12644);
xor U18145 (N_18145,N_15212,N_12586);
or U18146 (N_18146,N_14008,N_13709);
nor U18147 (N_18147,N_14234,N_15442);
or U18148 (N_18148,N_15119,N_13204);
and U18149 (N_18149,N_14083,N_13010);
or U18150 (N_18150,N_14584,N_13457);
and U18151 (N_18151,N_14867,N_13899);
nor U18152 (N_18152,N_15111,N_15017);
xor U18153 (N_18153,N_15586,N_15361);
nor U18154 (N_18154,N_13120,N_13759);
nand U18155 (N_18155,N_13989,N_15166);
nand U18156 (N_18156,N_15276,N_13734);
nand U18157 (N_18157,N_13808,N_14014);
nor U18158 (N_18158,N_12890,N_12682);
nand U18159 (N_18159,N_13091,N_14618);
and U18160 (N_18160,N_13739,N_14584);
nor U18161 (N_18161,N_12930,N_13700);
or U18162 (N_18162,N_13904,N_13710);
and U18163 (N_18163,N_15265,N_13872);
or U18164 (N_18164,N_14413,N_12833);
and U18165 (N_18165,N_14119,N_15342);
xnor U18166 (N_18166,N_12971,N_13120);
and U18167 (N_18167,N_14001,N_12917);
nor U18168 (N_18168,N_12623,N_12948);
or U18169 (N_18169,N_14202,N_14129);
nand U18170 (N_18170,N_13715,N_14152);
or U18171 (N_18171,N_13345,N_14166);
nand U18172 (N_18172,N_13264,N_13760);
nand U18173 (N_18173,N_15023,N_13179);
xnor U18174 (N_18174,N_13965,N_13628);
nand U18175 (N_18175,N_14781,N_15124);
nand U18176 (N_18176,N_14994,N_14148);
or U18177 (N_18177,N_12524,N_14650);
nand U18178 (N_18178,N_14781,N_15597);
nand U18179 (N_18179,N_13803,N_15237);
and U18180 (N_18180,N_13012,N_13079);
nor U18181 (N_18181,N_15240,N_14403);
and U18182 (N_18182,N_13895,N_14892);
nand U18183 (N_18183,N_14247,N_15448);
nor U18184 (N_18184,N_14769,N_14695);
or U18185 (N_18185,N_15169,N_12594);
nor U18186 (N_18186,N_14458,N_13219);
and U18187 (N_18187,N_12586,N_15314);
and U18188 (N_18188,N_12805,N_14574);
and U18189 (N_18189,N_14486,N_12847);
nand U18190 (N_18190,N_14582,N_14348);
and U18191 (N_18191,N_13109,N_13864);
and U18192 (N_18192,N_13554,N_14130);
and U18193 (N_18193,N_13023,N_14041);
or U18194 (N_18194,N_14947,N_14869);
xnor U18195 (N_18195,N_13026,N_14917);
and U18196 (N_18196,N_15428,N_15209);
nand U18197 (N_18197,N_13307,N_13500);
and U18198 (N_18198,N_13286,N_14610);
nand U18199 (N_18199,N_13538,N_13583);
and U18200 (N_18200,N_15139,N_15526);
and U18201 (N_18201,N_12848,N_14922);
nor U18202 (N_18202,N_12626,N_15571);
nand U18203 (N_18203,N_15288,N_15464);
and U18204 (N_18204,N_13237,N_14281);
or U18205 (N_18205,N_14442,N_15416);
and U18206 (N_18206,N_14767,N_15085);
nor U18207 (N_18207,N_14658,N_14316);
xor U18208 (N_18208,N_14378,N_13015);
nand U18209 (N_18209,N_12545,N_13364);
nor U18210 (N_18210,N_14805,N_13573);
nand U18211 (N_18211,N_14296,N_13383);
nor U18212 (N_18212,N_15079,N_13055);
xnor U18213 (N_18213,N_13007,N_12904);
nand U18214 (N_18214,N_15322,N_14091);
and U18215 (N_18215,N_14015,N_14064);
nand U18216 (N_18216,N_12819,N_14129);
or U18217 (N_18217,N_12917,N_14702);
or U18218 (N_18218,N_13403,N_13122);
and U18219 (N_18219,N_12940,N_14436);
nor U18220 (N_18220,N_14684,N_14056);
or U18221 (N_18221,N_14018,N_14315);
nor U18222 (N_18222,N_13666,N_13159);
and U18223 (N_18223,N_13039,N_14962);
or U18224 (N_18224,N_15556,N_14699);
or U18225 (N_18225,N_14539,N_14094);
xnor U18226 (N_18226,N_14254,N_12680);
nand U18227 (N_18227,N_15306,N_13446);
and U18228 (N_18228,N_14830,N_13861);
nand U18229 (N_18229,N_12663,N_14042);
and U18230 (N_18230,N_14466,N_14168);
nor U18231 (N_18231,N_12935,N_12880);
nor U18232 (N_18232,N_13045,N_15260);
or U18233 (N_18233,N_14833,N_14463);
or U18234 (N_18234,N_15202,N_15581);
nand U18235 (N_18235,N_13063,N_15509);
or U18236 (N_18236,N_13985,N_13866);
nor U18237 (N_18237,N_13484,N_14508);
or U18238 (N_18238,N_14514,N_13097);
and U18239 (N_18239,N_13438,N_13867);
nor U18240 (N_18240,N_13116,N_12505);
nor U18241 (N_18241,N_15112,N_12765);
or U18242 (N_18242,N_12643,N_14107);
or U18243 (N_18243,N_14363,N_12568);
xnor U18244 (N_18244,N_13834,N_15589);
and U18245 (N_18245,N_13133,N_13315);
nand U18246 (N_18246,N_13378,N_15127);
xnor U18247 (N_18247,N_13706,N_13728);
nor U18248 (N_18248,N_15136,N_13559);
nand U18249 (N_18249,N_13806,N_15215);
nand U18250 (N_18250,N_14240,N_14227);
or U18251 (N_18251,N_13051,N_12983);
nand U18252 (N_18252,N_12883,N_12812);
nor U18253 (N_18253,N_15510,N_13827);
or U18254 (N_18254,N_13779,N_14623);
or U18255 (N_18255,N_13829,N_13505);
xnor U18256 (N_18256,N_14595,N_13537);
and U18257 (N_18257,N_14835,N_15433);
nand U18258 (N_18258,N_13950,N_12896);
or U18259 (N_18259,N_14811,N_12718);
nand U18260 (N_18260,N_13904,N_13361);
or U18261 (N_18261,N_15125,N_14671);
and U18262 (N_18262,N_14774,N_13396);
nor U18263 (N_18263,N_12889,N_14876);
and U18264 (N_18264,N_13950,N_15334);
nor U18265 (N_18265,N_14784,N_14081);
nor U18266 (N_18266,N_13427,N_13108);
nor U18267 (N_18267,N_14127,N_12835);
nand U18268 (N_18268,N_14417,N_15487);
xnor U18269 (N_18269,N_15413,N_13785);
nor U18270 (N_18270,N_15245,N_15561);
nand U18271 (N_18271,N_15077,N_15324);
or U18272 (N_18272,N_13440,N_13050);
xnor U18273 (N_18273,N_13641,N_14123);
and U18274 (N_18274,N_12838,N_13026);
and U18275 (N_18275,N_15519,N_15449);
or U18276 (N_18276,N_13572,N_13398);
or U18277 (N_18277,N_15534,N_14284);
and U18278 (N_18278,N_15533,N_13119);
nand U18279 (N_18279,N_14458,N_14836);
and U18280 (N_18280,N_14959,N_14117);
nor U18281 (N_18281,N_13944,N_12707);
nand U18282 (N_18282,N_14023,N_13528);
nand U18283 (N_18283,N_14354,N_15021);
or U18284 (N_18284,N_15274,N_14793);
or U18285 (N_18285,N_13815,N_12501);
and U18286 (N_18286,N_15104,N_12776);
nor U18287 (N_18287,N_12748,N_13247);
nor U18288 (N_18288,N_14232,N_14953);
xnor U18289 (N_18289,N_15199,N_13227);
nand U18290 (N_18290,N_13060,N_12513);
nor U18291 (N_18291,N_15169,N_15363);
nand U18292 (N_18292,N_13153,N_13324);
nor U18293 (N_18293,N_14257,N_14493);
and U18294 (N_18294,N_12859,N_14677);
nand U18295 (N_18295,N_15378,N_14567);
nand U18296 (N_18296,N_14615,N_14950);
nand U18297 (N_18297,N_15285,N_12702);
or U18298 (N_18298,N_14119,N_12610);
and U18299 (N_18299,N_13439,N_14385);
and U18300 (N_18300,N_14372,N_13846);
and U18301 (N_18301,N_14439,N_12950);
nor U18302 (N_18302,N_14708,N_15303);
xnor U18303 (N_18303,N_13948,N_12811);
or U18304 (N_18304,N_14152,N_13240);
xnor U18305 (N_18305,N_13911,N_15035);
nand U18306 (N_18306,N_14643,N_13442);
or U18307 (N_18307,N_14997,N_12915);
xnor U18308 (N_18308,N_13754,N_14008);
or U18309 (N_18309,N_14995,N_15572);
xnor U18310 (N_18310,N_15472,N_12788);
nor U18311 (N_18311,N_15119,N_14263);
and U18312 (N_18312,N_13376,N_14894);
nor U18313 (N_18313,N_15501,N_13808);
or U18314 (N_18314,N_14611,N_12539);
nand U18315 (N_18315,N_13943,N_13850);
nand U18316 (N_18316,N_13862,N_15239);
or U18317 (N_18317,N_14485,N_15254);
and U18318 (N_18318,N_13603,N_15013);
nand U18319 (N_18319,N_14456,N_15211);
nand U18320 (N_18320,N_13970,N_13371);
xor U18321 (N_18321,N_14590,N_12514);
nor U18322 (N_18322,N_15242,N_12846);
and U18323 (N_18323,N_13763,N_12626);
nor U18324 (N_18324,N_15612,N_15311);
nor U18325 (N_18325,N_14352,N_12788);
nor U18326 (N_18326,N_15004,N_14581);
nand U18327 (N_18327,N_13820,N_14978);
and U18328 (N_18328,N_14424,N_14256);
and U18329 (N_18329,N_13907,N_15589);
or U18330 (N_18330,N_14229,N_12833);
or U18331 (N_18331,N_14628,N_15578);
or U18332 (N_18332,N_15489,N_13393);
nor U18333 (N_18333,N_13123,N_14933);
or U18334 (N_18334,N_12794,N_14425);
nor U18335 (N_18335,N_13499,N_13217);
nor U18336 (N_18336,N_13019,N_13488);
nand U18337 (N_18337,N_13709,N_15400);
nand U18338 (N_18338,N_14048,N_13329);
or U18339 (N_18339,N_14911,N_14921);
nor U18340 (N_18340,N_12823,N_14091);
and U18341 (N_18341,N_12971,N_15248);
nand U18342 (N_18342,N_14411,N_14770);
or U18343 (N_18343,N_14051,N_13808);
or U18344 (N_18344,N_13941,N_13810);
nor U18345 (N_18345,N_13255,N_14690);
nor U18346 (N_18346,N_13352,N_13226);
nand U18347 (N_18347,N_12643,N_13792);
nand U18348 (N_18348,N_13167,N_13788);
nand U18349 (N_18349,N_13295,N_14294);
or U18350 (N_18350,N_12700,N_12696);
or U18351 (N_18351,N_14196,N_13868);
nor U18352 (N_18352,N_15513,N_15047);
nand U18353 (N_18353,N_15281,N_12615);
xor U18354 (N_18354,N_13501,N_15324);
or U18355 (N_18355,N_15540,N_15062);
nand U18356 (N_18356,N_15496,N_12818);
nor U18357 (N_18357,N_13804,N_14766);
or U18358 (N_18358,N_14179,N_15255);
nor U18359 (N_18359,N_13870,N_14086);
nand U18360 (N_18360,N_13584,N_14332);
xnor U18361 (N_18361,N_15350,N_13482);
and U18362 (N_18362,N_14444,N_13926);
nor U18363 (N_18363,N_13258,N_14064);
nor U18364 (N_18364,N_13648,N_15386);
and U18365 (N_18365,N_15192,N_12616);
and U18366 (N_18366,N_13770,N_13101);
nor U18367 (N_18367,N_12802,N_12753);
nand U18368 (N_18368,N_13492,N_15059);
or U18369 (N_18369,N_14589,N_14719);
and U18370 (N_18370,N_14433,N_13019);
nand U18371 (N_18371,N_12792,N_15197);
or U18372 (N_18372,N_14249,N_13571);
nor U18373 (N_18373,N_15192,N_15110);
and U18374 (N_18374,N_12519,N_14939);
or U18375 (N_18375,N_12743,N_15336);
nor U18376 (N_18376,N_13424,N_14237);
or U18377 (N_18377,N_14681,N_14907);
nand U18378 (N_18378,N_13978,N_12546);
nand U18379 (N_18379,N_13134,N_13302);
nor U18380 (N_18380,N_14171,N_14365);
nand U18381 (N_18381,N_12865,N_15378);
or U18382 (N_18382,N_13050,N_15489);
or U18383 (N_18383,N_13175,N_13559);
and U18384 (N_18384,N_12537,N_14390);
nor U18385 (N_18385,N_12546,N_13898);
nand U18386 (N_18386,N_14609,N_14910);
and U18387 (N_18387,N_14181,N_15136);
xnor U18388 (N_18388,N_15358,N_14032);
nand U18389 (N_18389,N_15181,N_15139);
or U18390 (N_18390,N_12506,N_15426);
nor U18391 (N_18391,N_13752,N_13783);
or U18392 (N_18392,N_13962,N_13483);
and U18393 (N_18393,N_13921,N_14121);
nand U18394 (N_18394,N_13739,N_12534);
or U18395 (N_18395,N_14285,N_12519);
or U18396 (N_18396,N_15031,N_15201);
and U18397 (N_18397,N_13063,N_15241);
nand U18398 (N_18398,N_12567,N_12920);
or U18399 (N_18399,N_12731,N_13514);
or U18400 (N_18400,N_13948,N_12623);
or U18401 (N_18401,N_15452,N_13757);
or U18402 (N_18402,N_12506,N_12914);
nand U18403 (N_18403,N_14071,N_13939);
or U18404 (N_18404,N_14885,N_14889);
nor U18405 (N_18405,N_14421,N_13868);
and U18406 (N_18406,N_14801,N_13354);
nor U18407 (N_18407,N_13974,N_14466);
nor U18408 (N_18408,N_14051,N_14253);
and U18409 (N_18409,N_15189,N_13367);
nand U18410 (N_18410,N_12596,N_14565);
or U18411 (N_18411,N_13878,N_12918);
and U18412 (N_18412,N_14193,N_14210);
and U18413 (N_18413,N_15189,N_14515);
nand U18414 (N_18414,N_12576,N_15112);
nand U18415 (N_18415,N_14649,N_15489);
xnor U18416 (N_18416,N_13595,N_13207);
and U18417 (N_18417,N_13141,N_14281);
nor U18418 (N_18418,N_12561,N_13389);
and U18419 (N_18419,N_13877,N_15491);
and U18420 (N_18420,N_13151,N_14018);
or U18421 (N_18421,N_13107,N_13586);
or U18422 (N_18422,N_13915,N_13372);
or U18423 (N_18423,N_14968,N_15588);
and U18424 (N_18424,N_14086,N_14340);
nand U18425 (N_18425,N_14160,N_13839);
nor U18426 (N_18426,N_13996,N_15584);
xnor U18427 (N_18427,N_13857,N_14116);
nand U18428 (N_18428,N_15361,N_15271);
or U18429 (N_18429,N_13447,N_15330);
nand U18430 (N_18430,N_13949,N_15388);
or U18431 (N_18431,N_14815,N_13888);
or U18432 (N_18432,N_12588,N_12637);
nor U18433 (N_18433,N_13479,N_14416);
and U18434 (N_18434,N_13134,N_12588);
xor U18435 (N_18435,N_14322,N_12709);
or U18436 (N_18436,N_13196,N_12723);
nor U18437 (N_18437,N_15535,N_13557);
nor U18438 (N_18438,N_15171,N_13114);
nand U18439 (N_18439,N_15551,N_14061);
or U18440 (N_18440,N_12610,N_14832);
or U18441 (N_18441,N_15604,N_13868);
and U18442 (N_18442,N_13649,N_14554);
nand U18443 (N_18443,N_15196,N_13278);
and U18444 (N_18444,N_13148,N_12508);
nor U18445 (N_18445,N_12523,N_14016);
nand U18446 (N_18446,N_13591,N_14824);
nor U18447 (N_18447,N_13995,N_15542);
nand U18448 (N_18448,N_15053,N_15178);
or U18449 (N_18449,N_12921,N_15095);
or U18450 (N_18450,N_13317,N_12674);
nand U18451 (N_18451,N_13280,N_12959);
or U18452 (N_18452,N_15422,N_14979);
or U18453 (N_18453,N_12736,N_14167);
xor U18454 (N_18454,N_12748,N_15387);
or U18455 (N_18455,N_12767,N_12928);
nor U18456 (N_18456,N_15088,N_15199);
xor U18457 (N_18457,N_13727,N_14209);
and U18458 (N_18458,N_15523,N_13827);
nand U18459 (N_18459,N_13097,N_15185);
nor U18460 (N_18460,N_13400,N_14622);
nand U18461 (N_18461,N_15317,N_13055);
nand U18462 (N_18462,N_13335,N_14982);
and U18463 (N_18463,N_13597,N_14203);
or U18464 (N_18464,N_15484,N_14661);
nor U18465 (N_18465,N_13174,N_13802);
nand U18466 (N_18466,N_13013,N_13950);
nand U18467 (N_18467,N_13882,N_13483);
nand U18468 (N_18468,N_13577,N_15066);
xnor U18469 (N_18469,N_15350,N_15174);
nand U18470 (N_18470,N_14105,N_15187);
and U18471 (N_18471,N_14520,N_14029);
nor U18472 (N_18472,N_13104,N_14512);
nand U18473 (N_18473,N_14445,N_12968);
nor U18474 (N_18474,N_14505,N_13991);
and U18475 (N_18475,N_13468,N_12855);
nor U18476 (N_18476,N_12528,N_14713);
nor U18477 (N_18477,N_14636,N_13264);
or U18478 (N_18478,N_14253,N_14367);
nor U18479 (N_18479,N_13098,N_14147);
nand U18480 (N_18480,N_13541,N_14339);
nand U18481 (N_18481,N_14641,N_15144);
and U18482 (N_18482,N_12682,N_14371);
and U18483 (N_18483,N_13067,N_13274);
or U18484 (N_18484,N_14127,N_14231);
and U18485 (N_18485,N_13770,N_13662);
nor U18486 (N_18486,N_14439,N_15149);
and U18487 (N_18487,N_15167,N_13069);
or U18488 (N_18488,N_14922,N_14806);
and U18489 (N_18489,N_15032,N_13698);
nand U18490 (N_18490,N_14298,N_12979);
or U18491 (N_18491,N_12993,N_13803);
nor U18492 (N_18492,N_13763,N_12962);
xor U18493 (N_18493,N_13965,N_12533);
nor U18494 (N_18494,N_15346,N_14174);
or U18495 (N_18495,N_15531,N_13695);
nand U18496 (N_18496,N_15282,N_14610);
or U18497 (N_18497,N_13663,N_13618);
and U18498 (N_18498,N_13165,N_14053);
and U18499 (N_18499,N_15605,N_13243);
nand U18500 (N_18500,N_14489,N_14895);
and U18501 (N_18501,N_14775,N_15428);
nor U18502 (N_18502,N_15361,N_14762);
and U18503 (N_18503,N_15291,N_15091);
or U18504 (N_18504,N_15183,N_14299);
nand U18505 (N_18505,N_13832,N_15568);
and U18506 (N_18506,N_14853,N_14868);
and U18507 (N_18507,N_13777,N_15080);
or U18508 (N_18508,N_13994,N_13133);
nand U18509 (N_18509,N_13031,N_14550);
nor U18510 (N_18510,N_14375,N_12563);
or U18511 (N_18511,N_14700,N_13888);
and U18512 (N_18512,N_13928,N_14975);
or U18513 (N_18513,N_15294,N_14145);
and U18514 (N_18514,N_13016,N_15038);
nand U18515 (N_18515,N_14969,N_13391);
or U18516 (N_18516,N_13548,N_14730);
and U18517 (N_18517,N_15195,N_15425);
nor U18518 (N_18518,N_13770,N_14366);
or U18519 (N_18519,N_12940,N_14356);
nand U18520 (N_18520,N_14897,N_14483);
nor U18521 (N_18521,N_14033,N_14418);
nor U18522 (N_18522,N_13574,N_15047);
nand U18523 (N_18523,N_14132,N_13687);
nand U18524 (N_18524,N_13171,N_13229);
xnor U18525 (N_18525,N_13010,N_13841);
nor U18526 (N_18526,N_13230,N_14264);
nand U18527 (N_18527,N_14476,N_14226);
nand U18528 (N_18528,N_12938,N_13507);
nor U18529 (N_18529,N_15151,N_13396);
and U18530 (N_18530,N_14360,N_15396);
nor U18531 (N_18531,N_14480,N_14319);
nand U18532 (N_18532,N_14447,N_15222);
nor U18533 (N_18533,N_15210,N_14577);
or U18534 (N_18534,N_15167,N_15058);
xor U18535 (N_18535,N_15247,N_15371);
and U18536 (N_18536,N_13207,N_14635);
nand U18537 (N_18537,N_13846,N_13181);
xor U18538 (N_18538,N_14888,N_14748);
nand U18539 (N_18539,N_14220,N_15529);
nor U18540 (N_18540,N_14179,N_13138);
nor U18541 (N_18541,N_13868,N_14530);
or U18542 (N_18542,N_13046,N_12878);
or U18543 (N_18543,N_15449,N_15214);
nor U18544 (N_18544,N_13231,N_13211);
nor U18545 (N_18545,N_13426,N_13656);
nor U18546 (N_18546,N_12874,N_15249);
xor U18547 (N_18547,N_14733,N_12835);
nand U18548 (N_18548,N_13467,N_15356);
and U18549 (N_18549,N_12988,N_13340);
nand U18550 (N_18550,N_13163,N_15119);
nand U18551 (N_18551,N_13970,N_15585);
and U18552 (N_18552,N_14293,N_14417);
nor U18553 (N_18553,N_13872,N_14613);
and U18554 (N_18554,N_14269,N_14002);
nor U18555 (N_18555,N_14239,N_12641);
nor U18556 (N_18556,N_14741,N_12827);
nand U18557 (N_18557,N_15016,N_13316);
and U18558 (N_18558,N_13154,N_14767);
or U18559 (N_18559,N_13107,N_15006);
xnor U18560 (N_18560,N_12922,N_14415);
nor U18561 (N_18561,N_13475,N_14728);
nand U18562 (N_18562,N_12891,N_13858);
nor U18563 (N_18563,N_13143,N_12791);
and U18564 (N_18564,N_15364,N_12996);
or U18565 (N_18565,N_13348,N_15171);
xor U18566 (N_18566,N_12507,N_13902);
nor U18567 (N_18567,N_14408,N_15567);
nand U18568 (N_18568,N_14339,N_15217);
and U18569 (N_18569,N_15480,N_14080);
or U18570 (N_18570,N_14439,N_14221);
nor U18571 (N_18571,N_12745,N_15104);
nand U18572 (N_18572,N_13078,N_14994);
xor U18573 (N_18573,N_15171,N_14636);
or U18574 (N_18574,N_15109,N_14172);
or U18575 (N_18575,N_13075,N_15510);
nand U18576 (N_18576,N_14210,N_14602);
and U18577 (N_18577,N_14402,N_14947);
and U18578 (N_18578,N_13495,N_13377);
or U18579 (N_18579,N_13248,N_13874);
and U18580 (N_18580,N_12809,N_14510);
nand U18581 (N_18581,N_14851,N_15238);
nand U18582 (N_18582,N_15383,N_13483);
nor U18583 (N_18583,N_15262,N_13822);
and U18584 (N_18584,N_14923,N_13106);
nand U18585 (N_18585,N_13673,N_13666);
nand U18586 (N_18586,N_13113,N_13191);
nand U18587 (N_18587,N_14881,N_15003);
nor U18588 (N_18588,N_13367,N_13746);
or U18589 (N_18589,N_15176,N_13387);
and U18590 (N_18590,N_15412,N_15203);
nor U18591 (N_18591,N_15264,N_14578);
or U18592 (N_18592,N_13032,N_13515);
xor U18593 (N_18593,N_14017,N_13725);
and U18594 (N_18594,N_15398,N_13722);
nand U18595 (N_18595,N_15571,N_13219);
nor U18596 (N_18596,N_13084,N_14601);
or U18597 (N_18597,N_14116,N_13689);
and U18598 (N_18598,N_14272,N_15139);
and U18599 (N_18599,N_15051,N_13487);
xor U18600 (N_18600,N_13421,N_12801);
and U18601 (N_18601,N_13834,N_14419);
and U18602 (N_18602,N_13795,N_14156);
or U18603 (N_18603,N_15327,N_13616);
or U18604 (N_18604,N_14804,N_14972);
or U18605 (N_18605,N_15159,N_15104);
nand U18606 (N_18606,N_13629,N_12626);
nor U18607 (N_18607,N_14902,N_15440);
nor U18608 (N_18608,N_13255,N_14980);
nand U18609 (N_18609,N_13233,N_12577);
and U18610 (N_18610,N_15402,N_13344);
or U18611 (N_18611,N_14995,N_14589);
nor U18612 (N_18612,N_12956,N_15061);
or U18613 (N_18613,N_13381,N_14921);
and U18614 (N_18614,N_12805,N_13908);
nor U18615 (N_18615,N_13902,N_14893);
nor U18616 (N_18616,N_14825,N_14964);
and U18617 (N_18617,N_15571,N_13127);
and U18618 (N_18618,N_14141,N_14003);
or U18619 (N_18619,N_13779,N_13624);
nor U18620 (N_18620,N_14382,N_15422);
xor U18621 (N_18621,N_14292,N_13474);
nand U18622 (N_18622,N_14459,N_14593);
or U18623 (N_18623,N_15435,N_15490);
or U18624 (N_18624,N_13100,N_13509);
nor U18625 (N_18625,N_13973,N_14467);
nor U18626 (N_18626,N_13262,N_15003);
and U18627 (N_18627,N_14622,N_14830);
nand U18628 (N_18628,N_13542,N_12591);
and U18629 (N_18629,N_14979,N_13024);
and U18630 (N_18630,N_15133,N_14225);
nor U18631 (N_18631,N_15497,N_14142);
nor U18632 (N_18632,N_13839,N_14043);
xor U18633 (N_18633,N_13501,N_14928);
nand U18634 (N_18634,N_12580,N_12712);
and U18635 (N_18635,N_14810,N_13228);
or U18636 (N_18636,N_13007,N_14012);
and U18637 (N_18637,N_14498,N_14609);
and U18638 (N_18638,N_12976,N_13753);
nand U18639 (N_18639,N_12525,N_12895);
nor U18640 (N_18640,N_14862,N_15490);
and U18641 (N_18641,N_14910,N_12957);
and U18642 (N_18642,N_15106,N_15331);
nor U18643 (N_18643,N_15529,N_13797);
and U18644 (N_18644,N_14519,N_15441);
nor U18645 (N_18645,N_15300,N_13926);
nor U18646 (N_18646,N_15415,N_14969);
or U18647 (N_18647,N_13674,N_14013);
nand U18648 (N_18648,N_13211,N_15492);
nor U18649 (N_18649,N_14247,N_14450);
or U18650 (N_18650,N_13730,N_13184);
nor U18651 (N_18651,N_13860,N_14802);
xnor U18652 (N_18652,N_14286,N_14809);
nor U18653 (N_18653,N_14499,N_14568);
nand U18654 (N_18654,N_14363,N_13395);
or U18655 (N_18655,N_13233,N_13492);
and U18656 (N_18656,N_12741,N_13241);
nor U18657 (N_18657,N_15057,N_14803);
or U18658 (N_18658,N_14360,N_15522);
or U18659 (N_18659,N_14826,N_14727);
or U18660 (N_18660,N_13807,N_14074);
or U18661 (N_18661,N_13188,N_12745);
or U18662 (N_18662,N_12913,N_12697);
and U18663 (N_18663,N_14704,N_13443);
or U18664 (N_18664,N_14241,N_12569);
nor U18665 (N_18665,N_13517,N_13875);
or U18666 (N_18666,N_13886,N_15024);
xor U18667 (N_18667,N_15244,N_14957);
and U18668 (N_18668,N_13348,N_13411);
xnor U18669 (N_18669,N_15115,N_14070);
nand U18670 (N_18670,N_14476,N_13871);
and U18671 (N_18671,N_12657,N_14743);
nor U18672 (N_18672,N_13127,N_14936);
or U18673 (N_18673,N_14186,N_13330);
and U18674 (N_18674,N_12922,N_15475);
or U18675 (N_18675,N_12788,N_15114);
xor U18676 (N_18676,N_13580,N_14829);
or U18677 (N_18677,N_15159,N_15384);
and U18678 (N_18678,N_13855,N_15033);
and U18679 (N_18679,N_13260,N_15587);
or U18680 (N_18680,N_12605,N_14088);
nand U18681 (N_18681,N_14987,N_14740);
or U18682 (N_18682,N_14486,N_14566);
or U18683 (N_18683,N_14532,N_13364);
nor U18684 (N_18684,N_15519,N_14729);
nand U18685 (N_18685,N_13920,N_13277);
and U18686 (N_18686,N_12838,N_14005);
nand U18687 (N_18687,N_14656,N_14538);
and U18688 (N_18688,N_13160,N_15598);
nor U18689 (N_18689,N_14963,N_15050);
nand U18690 (N_18690,N_13831,N_13707);
or U18691 (N_18691,N_15214,N_14681);
nand U18692 (N_18692,N_14152,N_13371);
and U18693 (N_18693,N_12590,N_13521);
nor U18694 (N_18694,N_13204,N_12682);
xor U18695 (N_18695,N_15160,N_14747);
nand U18696 (N_18696,N_12782,N_15601);
or U18697 (N_18697,N_12964,N_14142);
and U18698 (N_18698,N_13073,N_15232);
and U18699 (N_18699,N_14485,N_13700);
or U18700 (N_18700,N_14609,N_14001);
nand U18701 (N_18701,N_14508,N_12735);
and U18702 (N_18702,N_13775,N_15140);
xor U18703 (N_18703,N_14878,N_14711);
nand U18704 (N_18704,N_13931,N_14539);
nor U18705 (N_18705,N_15270,N_12621);
nand U18706 (N_18706,N_13281,N_15373);
xnor U18707 (N_18707,N_13424,N_12560);
or U18708 (N_18708,N_15469,N_13310);
or U18709 (N_18709,N_13436,N_13350);
and U18710 (N_18710,N_13361,N_14885);
nand U18711 (N_18711,N_12626,N_15184);
and U18712 (N_18712,N_15510,N_15554);
or U18713 (N_18713,N_13360,N_14890);
and U18714 (N_18714,N_14904,N_12953);
nand U18715 (N_18715,N_15387,N_13919);
or U18716 (N_18716,N_14055,N_14461);
nor U18717 (N_18717,N_15111,N_13268);
nand U18718 (N_18718,N_14325,N_13159);
nor U18719 (N_18719,N_15298,N_14774);
nor U18720 (N_18720,N_15206,N_15615);
nor U18721 (N_18721,N_13388,N_13460);
or U18722 (N_18722,N_14002,N_13926);
nand U18723 (N_18723,N_13985,N_13376);
xnor U18724 (N_18724,N_13109,N_12556);
nand U18725 (N_18725,N_14101,N_13321);
and U18726 (N_18726,N_13041,N_15170);
nor U18727 (N_18727,N_13241,N_13505);
xnor U18728 (N_18728,N_14772,N_15512);
or U18729 (N_18729,N_14368,N_13418);
or U18730 (N_18730,N_13064,N_12917);
nor U18731 (N_18731,N_12826,N_15102);
nand U18732 (N_18732,N_13226,N_15549);
nor U18733 (N_18733,N_14251,N_12729);
or U18734 (N_18734,N_14211,N_13223);
nor U18735 (N_18735,N_14047,N_13751);
or U18736 (N_18736,N_13950,N_15391);
nor U18737 (N_18737,N_15392,N_13510);
nand U18738 (N_18738,N_12653,N_14220);
nor U18739 (N_18739,N_15197,N_14119);
nor U18740 (N_18740,N_13605,N_14282);
and U18741 (N_18741,N_15432,N_13260);
nor U18742 (N_18742,N_15154,N_13711);
nand U18743 (N_18743,N_13071,N_14250);
nor U18744 (N_18744,N_12819,N_15319);
and U18745 (N_18745,N_13686,N_13723);
or U18746 (N_18746,N_15329,N_14608);
nor U18747 (N_18747,N_14271,N_12843);
xor U18748 (N_18748,N_13296,N_15292);
nand U18749 (N_18749,N_14125,N_13994);
nor U18750 (N_18750,N_15965,N_18424);
nor U18751 (N_18751,N_16664,N_16399);
or U18752 (N_18752,N_17156,N_16343);
xor U18753 (N_18753,N_17455,N_16159);
nand U18754 (N_18754,N_16445,N_16708);
and U18755 (N_18755,N_17054,N_16505);
xor U18756 (N_18756,N_17074,N_17789);
or U18757 (N_18757,N_17110,N_17702);
or U18758 (N_18758,N_17095,N_18552);
nor U18759 (N_18759,N_18721,N_16068);
xnor U18760 (N_18760,N_18266,N_16265);
nand U18761 (N_18761,N_15658,N_18065);
and U18762 (N_18762,N_15715,N_18637);
nor U18763 (N_18763,N_18548,N_17986);
and U18764 (N_18764,N_16342,N_17280);
nor U18765 (N_18765,N_16299,N_16800);
nor U18766 (N_18766,N_16689,N_18503);
or U18767 (N_18767,N_15968,N_15687);
or U18768 (N_18768,N_16564,N_16997);
nand U18769 (N_18769,N_17570,N_16697);
and U18770 (N_18770,N_17884,N_18416);
nand U18771 (N_18771,N_17299,N_17154);
nor U18772 (N_18772,N_16570,N_15857);
and U18773 (N_18773,N_17676,N_18563);
or U18774 (N_18774,N_17498,N_16055);
and U18775 (N_18775,N_16527,N_17984);
nor U18776 (N_18776,N_17288,N_17893);
and U18777 (N_18777,N_16216,N_16157);
nand U18778 (N_18778,N_16455,N_16001);
nor U18779 (N_18779,N_18110,N_17077);
and U18780 (N_18780,N_18694,N_18437);
nor U18781 (N_18781,N_16734,N_16281);
xnor U18782 (N_18782,N_17452,N_18665);
nand U18783 (N_18783,N_18556,N_15826);
nor U18784 (N_18784,N_16757,N_16073);
nand U18785 (N_18785,N_18641,N_17963);
nor U18786 (N_18786,N_18335,N_16475);
nand U18787 (N_18787,N_16306,N_18484);
and U18788 (N_18788,N_17257,N_15856);
nor U18789 (N_18789,N_17476,N_17086);
nor U18790 (N_18790,N_18032,N_17786);
or U18791 (N_18791,N_15911,N_17582);
nand U18792 (N_18792,N_18570,N_16197);
or U18793 (N_18793,N_18398,N_16899);
nand U18794 (N_18794,N_17733,N_18425);
or U18795 (N_18795,N_16992,N_16226);
or U18796 (N_18796,N_18175,N_16155);
or U18797 (N_18797,N_18452,N_16245);
or U18798 (N_18798,N_18649,N_16900);
or U18799 (N_18799,N_16132,N_17489);
or U18800 (N_18800,N_17849,N_17309);
or U18801 (N_18801,N_17898,N_18714);
nand U18802 (N_18802,N_18667,N_18729);
xnor U18803 (N_18803,N_17001,N_16628);
nor U18804 (N_18804,N_15957,N_18114);
xnor U18805 (N_18805,N_16936,N_18281);
xnor U18806 (N_18806,N_17332,N_17279);
nand U18807 (N_18807,N_18577,N_16759);
nor U18808 (N_18808,N_17401,N_18487);
nor U18809 (N_18809,N_17347,N_17363);
nand U18810 (N_18810,N_16507,N_17266);
nor U18811 (N_18811,N_16685,N_17615);
and U18812 (N_18812,N_16098,N_16634);
nor U18813 (N_18813,N_17329,N_16890);
or U18814 (N_18814,N_17989,N_17715);
nor U18815 (N_18815,N_15932,N_18274);
xnor U18816 (N_18816,N_15811,N_17404);
nor U18817 (N_18817,N_17620,N_16533);
nor U18818 (N_18818,N_17837,N_15812);
or U18819 (N_18819,N_16893,N_18012);
and U18820 (N_18820,N_18346,N_16136);
nor U18821 (N_18821,N_16450,N_17527);
and U18822 (N_18822,N_18286,N_18597);
nor U18823 (N_18823,N_17794,N_17284);
or U18824 (N_18824,N_17604,N_16538);
or U18825 (N_18825,N_16926,N_16665);
nand U18826 (N_18826,N_16719,N_15706);
nor U18827 (N_18827,N_17291,N_18308);
nor U18828 (N_18828,N_18463,N_16416);
or U18829 (N_18829,N_18609,N_15922);
or U18830 (N_18830,N_17999,N_16753);
nand U18831 (N_18831,N_18476,N_18048);
nand U18832 (N_18832,N_15738,N_17477);
nand U18833 (N_18833,N_17651,N_17803);
or U18834 (N_18834,N_17449,N_18426);
nor U18835 (N_18835,N_16693,N_17448);
nand U18836 (N_18836,N_17192,N_18304);
and U18837 (N_18837,N_18368,N_18344);
nor U18838 (N_18838,N_18545,N_18671);
or U18839 (N_18839,N_15888,N_17507);
nand U18840 (N_18840,N_16508,N_16384);
and U18841 (N_18841,N_18373,N_18250);
nor U18842 (N_18842,N_18525,N_17729);
nand U18843 (N_18843,N_15972,N_15651);
xor U18844 (N_18844,N_18047,N_18633);
nand U18845 (N_18845,N_16004,N_17305);
nand U18846 (N_18846,N_17857,N_17464);
or U18847 (N_18847,N_18343,N_18064);
and U18848 (N_18848,N_18294,N_18388);
and U18849 (N_18849,N_16637,N_17487);
nand U18850 (N_18850,N_17160,N_16646);
nor U18851 (N_18851,N_17630,N_17890);
nor U18852 (N_18852,N_18247,N_18567);
nor U18853 (N_18853,N_17688,N_16441);
and U18854 (N_18854,N_16189,N_18735);
xnor U18855 (N_18855,N_16577,N_18385);
nor U18856 (N_18856,N_16559,N_18334);
nand U18857 (N_18857,N_17956,N_17506);
nor U18858 (N_18858,N_15809,N_17435);
and U18859 (N_18859,N_17317,N_17508);
or U18860 (N_18860,N_16710,N_16582);
or U18861 (N_18861,N_16949,N_18349);
nor U18862 (N_18862,N_18742,N_17005);
and U18863 (N_18863,N_15966,N_17550);
nor U18864 (N_18864,N_18302,N_17597);
or U18865 (N_18865,N_18131,N_18283);
or U18866 (N_18866,N_18038,N_17365);
nand U18867 (N_18867,N_16295,N_16186);
or U18868 (N_18868,N_18521,N_16539);
or U18869 (N_18869,N_18477,N_18256);
nand U18870 (N_18870,N_17191,N_18236);
or U18871 (N_18871,N_17722,N_17995);
or U18872 (N_18872,N_18314,N_15976);
nand U18873 (N_18873,N_18449,N_17566);
nand U18874 (N_18874,N_18044,N_18643);
and U18875 (N_18875,N_16609,N_18025);
nor U18876 (N_18876,N_16297,N_18178);
and U18877 (N_18877,N_16263,N_17020);
and U18878 (N_18878,N_16131,N_16581);
nand U18879 (N_18879,N_16781,N_16790);
nor U18880 (N_18880,N_15998,N_18124);
and U18881 (N_18881,N_15853,N_17934);
nand U18882 (N_18882,N_16077,N_17410);
nor U18883 (N_18883,N_18046,N_17018);
nor U18884 (N_18884,N_18713,N_15654);
nand U18885 (N_18885,N_16133,N_17343);
or U18886 (N_18886,N_16464,N_17824);
nor U18887 (N_18887,N_16712,N_16687);
nor U18888 (N_18888,N_17345,N_16544);
nand U18889 (N_18889,N_17783,N_17817);
or U18890 (N_18890,N_18541,N_16663);
nor U18891 (N_18891,N_17013,N_17606);
and U18892 (N_18892,N_18033,N_16522);
nor U18893 (N_18893,N_16404,N_17631);
and U18894 (N_18894,N_16597,N_16983);
and U18895 (N_18895,N_18214,N_16830);
xnor U18896 (N_18896,N_17927,N_18153);
and U18897 (N_18897,N_18093,N_16094);
and U18898 (N_18898,N_15884,N_15883);
and U18899 (N_18899,N_15784,N_18389);
xor U18900 (N_18900,N_16877,N_18305);
and U18901 (N_18901,N_17777,N_18573);
nor U18902 (N_18902,N_18352,N_15690);
and U18903 (N_18903,N_16692,N_16779);
nor U18904 (N_18904,N_17860,N_16161);
and U18905 (N_18905,N_16383,N_17264);
or U18906 (N_18906,N_18387,N_16035);
xor U18907 (N_18907,N_16876,N_16914);
nand U18908 (N_18908,N_15930,N_15807);
nand U18909 (N_18909,N_18075,N_18000);
or U18910 (N_18910,N_18074,N_17744);
and U18911 (N_18911,N_17248,N_15788);
xnor U18912 (N_18912,N_16504,N_18692);
xnor U18913 (N_18913,N_17058,N_18138);
nor U18914 (N_18914,N_15837,N_16961);
or U18915 (N_18915,N_16179,N_15937);
or U18916 (N_18916,N_17321,N_17384);
nand U18917 (N_18917,N_17953,N_17395);
nand U18918 (N_18918,N_16206,N_18696);
and U18919 (N_18919,N_17928,N_17009);
nand U18920 (N_18920,N_16232,N_17308);
or U18921 (N_18921,N_17938,N_17896);
and U18922 (N_18922,N_16082,N_15744);
nor U18923 (N_18923,N_18052,N_16229);
and U18924 (N_18924,N_18470,N_16408);
xnor U18925 (N_18925,N_16502,N_16390);
nand U18926 (N_18926,N_16543,N_15644);
and U18927 (N_18927,N_18260,N_17823);
nand U18928 (N_18928,N_15944,N_16878);
nor U18929 (N_18929,N_16151,N_16561);
xnor U18930 (N_18930,N_15885,N_17149);
and U18931 (N_18931,N_18037,N_17627);
nor U18932 (N_18932,N_17381,N_18181);
and U18933 (N_18933,N_16081,N_18510);
nand U18934 (N_18934,N_17352,N_18288);
nand U18935 (N_18935,N_16501,N_18591);
nand U18936 (N_18936,N_18013,N_17840);
or U18937 (N_18937,N_16647,N_17705);
or U18938 (N_18938,N_18413,N_17866);
nand U18939 (N_18939,N_17011,N_15909);
or U18940 (N_18940,N_15716,N_16856);
xor U18941 (N_18941,N_16468,N_18489);
nor U18942 (N_18942,N_18170,N_17208);
nand U18943 (N_18943,N_18396,N_18727);
nand U18944 (N_18944,N_16492,N_16848);
xnor U18945 (N_18945,N_16407,N_17788);
nor U18946 (N_18946,N_16086,N_16403);
nor U18947 (N_18947,N_18122,N_15795);
and U18948 (N_18948,N_18318,N_18595);
or U18949 (N_18949,N_16520,N_16929);
nor U18950 (N_18950,N_18369,N_17976);
nand U18951 (N_18951,N_17116,N_18420);
nor U18952 (N_18952,N_15996,N_18007);
nand U18953 (N_18953,N_17377,N_15820);
nor U18954 (N_18954,N_17559,N_17367);
and U18955 (N_18955,N_16181,N_16436);
nor U18956 (N_18956,N_18513,N_17406);
and U18957 (N_18957,N_15951,N_15823);
nand U18958 (N_18958,N_17580,N_17856);
nor U18959 (N_18959,N_18345,N_17358);
or U18960 (N_18960,N_16050,N_17808);
nand U18961 (N_18961,N_16957,N_18472);
nand U18962 (N_18962,N_15803,N_18002);
nand U18963 (N_18963,N_18241,N_17717);
xor U18964 (N_18964,N_17617,N_18540);
and U18965 (N_18965,N_18496,N_17790);
nand U18966 (N_18966,N_15630,N_16023);
nor U18967 (N_18967,N_17344,N_15844);
and U18968 (N_18968,N_16944,N_17601);
xnor U18969 (N_18969,N_17174,N_18277);
and U18970 (N_18970,N_17387,N_16818);
or U18971 (N_18971,N_17323,N_18378);
nand U18972 (N_18972,N_17542,N_16483);
or U18973 (N_18973,N_18354,N_18623);
or U18974 (N_18974,N_16472,N_17441);
xnor U18975 (N_18975,N_17867,N_16458);
xnor U18976 (N_18976,N_16648,N_16409);
xor U18977 (N_18977,N_17669,N_15890);
nand U18978 (N_18978,N_17776,N_18140);
nand U18979 (N_18979,N_17211,N_18723);
or U18980 (N_18980,N_17543,N_17481);
nand U18981 (N_18981,N_16242,N_18135);
xor U18982 (N_18982,N_17947,N_17787);
and U18983 (N_18983,N_16274,N_15833);
and U18984 (N_18984,N_16851,N_16661);
nand U18985 (N_18985,N_15950,N_17240);
or U18986 (N_18986,N_16309,N_17621);
nand U18987 (N_18987,N_15747,N_18417);
nand U18988 (N_18988,N_15628,N_17206);
nor U18989 (N_18989,N_15882,N_17534);
nor U18990 (N_18990,N_17662,N_16715);
xnor U18991 (N_18991,N_16378,N_16487);
and U18992 (N_18992,N_18231,N_16578);
nor U18993 (N_18993,N_18392,N_18180);
and U18994 (N_18994,N_16204,N_18251);
nor U18995 (N_18995,N_16304,N_16454);
or U18996 (N_18996,N_16529,N_18056);
or U18997 (N_18997,N_15871,N_18126);
or U18998 (N_18998,N_18681,N_17017);
xor U18999 (N_18999,N_16188,N_18116);
xnor U19000 (N_19000,N_16747,N_15785);
nor U19001 (N_19001,N_18078,N_15652);
and U19002 (N_19002,N_16447,N_18450);
or U19003 (N_19003,N_16739,N_16496);
nand U19004 (N_19004,N_18339,N_16735);
nor U19005 (N_19005,N_16118,N_15880);
nand U19006 (N_19006,N_15799,N_17034);
nor U19007 (N_19007,N_16981,N_15717);
or U19008 (N_19008,N_18526,N_16532);
nand U19009 (N_19009,N_17515,N_15735);
nor U19010 (N_19010,N_16208,N_17210);
nor U19011 (N_19011,N_16334,N_16150);
and U19012 (N_19012,N_18159,N_18071);
and U19013 (N_19013,N_17518,N_18278);
nand U19014 (N_19014,N_17212,N_15660);
and U19015 (N_19015,N_17125,N_16859);
and U19016 (N_19016,N_16398,N_15679);
nand U19017 (N_19017,N_16725,N_16224);
or U19018 (N_19018,N_18559,N_17497);
or U19019 (N_19019,N_18148,N_18726);
and U19020 (N_19020,N_16410,N_18401);
or U19021 (N_19021,N_17030,N_16461);
nor U19022 (N_19022,N_16785,N_16322);
and U19023 (N_19023,N_17663,N_18357);
nand U19024 (N_19024,N_17331,N_18341);
xor U19025 (N_19025,N_17207,N_16430);
or U19026 (N_19026,N_16928,N_16874);
nand U19027 (N_19027,N_16824,N_16531);
xnor U19028 (N_19028,N_17892,N_17251);
nor U19029 (N_19029,N_16655,N_17623);
nor U19030 (N_19030,N_16889,N_17739);
xnor U19031 (N_19031,N_17392,N_15742);
nand U19032 (N_19032,N_15991,N_17727);
or U19033 (N_19033,N_15924,N_16215);
nand U19034 (N_19034,N_17104,N_17393);
and U19035 (N_19035,N_17761,N_16626);
xor U19036 (N_19036,N_17502,N_17460);
nand U19037 (N_19037,N_17238,N_18495);
nor U19038 (N_19038,N_17573,N_17523);
nor U19039 (N_19039,N_16995,N_16110);
nand U19040 (N_19040,N_17980,N_16421);
xnor U19041 (N_19041,N_15761,N_18100);
or U19042 (N_19042,N_17258,N_18230);
nor U19043 (N_19043,N_17142,N_16090);
or U19044 (N_19044,N_15855,N_16194);
or U19045 (N_19045,N_16611,N_17260);
nand U19046 (N_19046,N_16971,N_16250);
nand U19047 (N_19047,N_18393,N_17848);
nor U19048 (N_19048,N_16317,N_16310);
xor U19049 (N_19049,N_15946,N_18394);
xor U19050 (N_19050,N_16528,N_17960);
nor U19051 (N_19051,N_17126,N_18136);
nand U19052 (N_19052,N_17895,N_16121);
nor U19053 (N_19053,N_16395,N_15737);
nand U19054 (N_19054,N_16838,N_16970);
or U19055 (N_19055,N_16463,N_16249);
and U19056 (N_19056,N_16964,N_18087);
nor U19057 (N_19057,N_15867,N_17673);
xnor U19058 (N_19058,N_17970,N_16515);
or U19059 (N_19059,N_15943,N_16761);
nor U19060 (N_19060,N_18598,N_16059);
nor U19061 (N_19061,N_16037,N_16462);
nor U19062 (N_19062,N_16752,N_18362);
or U19063 (N_19063,N_16006,N_15659);
nor U19064 (N_19064,N_17851,N_16172);
xnor U19065 (N_19065,N_16010,N_16868);
or U19066 (N_19066,N_17170,N_16488);
nor U19067 (N_19067,N_16241,N_17233);
nor U19068 (N_19068,N_16572,N_15763);
nor U19069 (N_19069,N_16256,N_18740);
and U19070 (N_19070,N_16567,N_17549);
nand U19071 (N_19071,N_18182,N_16335);
nand U19072 (N_19072,N_16580,N_17157);
and U19073 (N_19073,N_17637,N_18421);
and U19074 (N_19074,N_18199,N_18383);
xor U19075 (N_19075,N_16788,N_17403);
or U19076 (N_19076,N_17021,N_16311);
nand U19077 (N_19077,N_16716,N_17419);
nand U19078 (N_19078,N_15645,N_16415);
xor U19079 (N_19079,N_17762,N_16610);
or U19080 (N_19080,N_18174,N_15663);
nand U19081 (N_19081,N_18298,N_17270);
xor U19082 (N_19082,N_17581,N_18678);
and U19083 (N_19083,N_16321,N_16174);
nand U19084 (N_19084,N_16481,N_17906);
or U19085 (N_19085,N_16221,N_16866);
nor U19086 (N_19086,N_18269,N_17526);
or U19087 (N_19087,N_18123,N_18455);
nor U19088 (N_19088,N_16205,N_18379);
xor U19089 (N_19089,N_17708,N_18118);
or U19090 (N_19090,N_18322,N_16618);
and U19091 (N_19091,N_16932,N_17841);
nand U19092 (N_19092,N_16474,N_16579);
nor U19093 (N_19093,N_15668,N_16828);
and U19094 (N_19094,N_18143,N_16773);
nand U19095 (N_19095,N_16545,N_16969);
nand U19096 (N_19096,N_18720,N_18458);
or U19097 (N_19097,N_18222,N_17665);
nand U19098 (N_19098,N_18235,N_16809);
nand U19099 (N_19099,N_18034,N_18683);
and U19100 (N_19100,N_16018,N_17902);
nor U19101 (N_19101,N_17805,N_15649);
nand U19102 (N_19102,N_16509,N_18265);
nand U19103 (N_19103,N_17852,N_18493);
or U19104 (N_19104,N_18200,N_17929);
or U19105 (N_19105,N_16099,N_16540);
or U19106 (N_19106,N_15889,N_17535);
nand U19107 (N_19107,N_16910,N_18359);
nor U19108 (N_19108,N_16816,N_16602);
xor U19109 (N_19109,N_16742,N_16775);
or U19110 (N_19110,N_17796,N_16290);
and U19111 (N_19111,N_17073,N_15635);
nor U19112 (N_19112,N_17706,N_15854);
nor U19113 (N_19113,N_16794,N_17473);
or U19114 (N_19114,N_17505,N_17775);
nor U19115 (N_19115,N_18254,N_18168);
nor U19116 (N_19116,N_18042,N_18730);
and U19117 (N_19117,N_17565,N_17672);
nand U19118 (N_19118,N_17296,N_15755);
xnor U19119 (N_19119,N_17613,N_17194);
xor U19120 (N_19120,N_18519,N_18478);
and U19121 (N_19121,N_17988,N_17561);
or U19122 (N_19122,N_18099,N_18672);
or U19123 (N_19123,N_16175,N_17002);
xor U19124 (N_19124,N_17289,N_16705);
nor U19125 (N_19125,N_17735,N_16593);
or U19126 (N_19126,N_16095,N_16392);
or U19127 (N_19127,N_16111,N_17484);
nand U19128 (N_19128,N_17184,N_17568);
and U19129 (N_19129,N_16147,N_17065);
nor U19130 (N_19130,N_17319,N_15886);
nor U19131 (N_19131,N_18707,N_16296);
nand U19132 (N_19132,N_16514,N_17548);
or U19133 (N_19133,N_18512,N_15859);
nor U19134 (N_19134,N_18480,N_18246);
and U19135 (N_19135,N_16884,N_18043);
xnor U19136 (N_19136,N_18252,N_17052);
xor U19137 (N_19137,N_17080,N_17300);
nor U19138 (N_19138,N_18055,N_18491);
nor U19139 (N_19139,N_18360,N_17802);
nand U19140 (N_19140,N_16337,N_16134);
nand U19141 (N_19141,N_16998,N_18511);
xnor U19142 (N_19142,N_16521,N_16280);
nor U19143 (N_19143,N_16016,N_18611);
nand U19144 (N_19144,N_18716,N_17063);
and U19145 (N_19145,N_16019,N_17391);
and U19146 (N_19146,N_18160,N_18021);
or U19147 (N_19147,N_15987,N_18482);
nor U19148 (N_19148,N_18337,N_15653);
nor U19149 (N_19149,N_17180,N_16126);
and U19150 (N_19150,N_16353,N_18375);
or U19151 (N_19151,N_16801,N_17353);
xor U19152 (N_19152,N_16733,N_16990);
nand U19153 (N_19153,N_17780,N_18332);
or U19154 (N_19154,N_16918,N_17166);
and U19155 (N_19155,N_17726,N_16369);
nand U19156 (N_19156,N_16085,N_17610);
and U19157 (N_19157,N_17055,N_15749);
or U19158 (N_19158,N_16960,N_18045);
nand U19159 (N_19159,N_17218,N_18376);
xnor U19160 (N_19160,N_15764,N_16479);
nor U19161 (N_19161,N_17853,N_15860);
or U19162 (N_19162,N_16873,N_18494);
and U19163 (N_19163,N_15891,N_17977);
and U19164 (N_19164,N_15810,N_16033);
or U19165 (N_19165,N_17112,N_18586);
or U19166 (N_19166,N_15895,N_16104);
nor U19167 (N_19167,N_17333,N_16113);
nand U19168 (N_19168,N_16560,N_16114);
nor U19169 (N_19169,N_15956,N_17835);
nand U19170 (N_19170,N_16328,N_16935);
nand U19171 (N_19171,N_15636,N_18647);
or U19172 (N_19172,N_17129,N_18745);
nand U19173 (N_19173,N_16552,N_18121);
or U19174 (N_19174,N_15787,N_17197);
or U19175 (N_19175,N_16273,N_16102);
nor U19176 (N_19176,N_17390,N_16677);
or U19177 (N_19177,N_18028,N_18502);
and U19178 (N_19178,N_15695,N_18197);
or U19179 (N_19179,N_15999,N_17509);
or U19180 (N_19180,N_18558,N_18657);
or U19181 (N_19181,N_17680,N_18749);
or U19182 (N_19182,N_16105,N_15701);
xnor U19183 (N_19183,N_15846,N_17081);
or U19184 (N_19184,N_17492,N_17622);
nor U19185 (N_19185,N_17532,N_17459);
and U19186 (N_19186,N_17290,N_17096);
or U19187 (N_19187,N_16805,N_17701);
or U19188 (N_19188,N_17774,N_16727);
nand U19189 (N_19189,N_15769,N_17538);
or U19190 (N_19190,N_15835,N_16200);
or U19191 (N_19191,N_17742,N_17176);
and U19192 (N_19192,N_18418,N_15813);
xor U19193 (N_19193,N_15915,N_18529);
nand U19194 (N_19194,N_15754,N_16456);
nand U19195 (N_19195,N_16420,N_17626);
or U19196 (N_19196,N_16275,N_18731);
nor U19197 (N_19197,N_18640,N_15863);
and U19198 (N_19198,N_18361,N_17119);
and U19199 (N_19199,N_17059,N_17342);
nor U19200 (N_19200,N_18460,N_17696);
nand U19201 (N_19201,N_16239,N_18473);
or U19202 (N_19202,N_16429,N_17640);
and U19203 (N_19203,N_17262,N_15758);
xnor U19204 (N_19204,N_18439,N_18432);
nor U19205 (N_19205,N_17457,N_16282);
nor U19206 (N_19206,N_16075,N_16919);
and U19207 (N_19207,N_17148,N_16798);
or U19208 (N_19208,N_16007,N_18355);
nand U19209 (N_19209,N_16236,N_15851);
and U19210 (N_19210,N_18268,N_18498);
nor U19211 (N_19211,N_17983,N_16302);
xor U19212 (N_19212,N_18475,N_16437);
and U19213 (N_19213,N_16924,N_16840);
nand U19214 (N_19214,N_16649,N_18677);
nand U19215 (N_19215,N_17415,N_16193);
nand U19216 (N_19216,N_17799,N_16259);
and U19217 (N_19217,N_16225,N_18132);
nor U19218 (N_19218,N_17341,N_18506);
xor U19219 (N_19219,N_17655,N_17730);
nor U19220 (N_19220,N_18184,N_18625);
nor U19221 (N_19221,N_17765,N_16030);
and U19222 (N_19222,N_16883,N_17227);
and U19223 (N_19223,N_16489,N_16839);
nor U19224 (N_19224,N_15732,N_15776);
and U19225 (N_19225,N_15815,N_16278);
nor U19226 (N_19226,N_15993,N_16366);
nand U19227 (N_19227,N_15678,N_17528);
and U19228 (N_19228,N_16888,N_16344);
and U19229 (N_19229,N_16015,N_18005);
or U19230 (N_19230,N_16927,N_17355);
nand U19231 (N_19231,N_17757,N_18638);
and U19232 (N_19232,N_18732,N_17529);
and U19233 (N_19233,N_16323,N_18019);
nand U19234 (N_19234,N_18736,N_17402);
nand U19235 (N_19235,N_16815,N_18436);
and U19236 (N_19236,N_18682,N_17829);
xnor U19237 (N_19237,N_16553,N_18627);
xor U19238 (N_19238,N_17195,N_16285);
and U19239 (N_19239,N_16536,N_15816);
nor U19240 (N_19240,N_17027,N_16402);
nor U19241 (N_19241,N_15825,N_17022);
xnor U19242 (N_19242,N_16619,N_17249);
or U19243 (N_19243,N_16031,N_16203);
and U19244 (N_19244,N_16558,N_18205);
or U19245 (N_19245,N_16040,N_15722);
nor U19246 (N_19246,N_16541,N_15865);
or U19247 (N_19247,N_17771,N_18146);
and U19248 (N_19248,N_15961,N_16101);
and U19249 (N_19249,N_17854,N_16897);
and U19250 (N_19250,N_18722,N_17911);
and U19251 (N_19251,N_16300,N_15675);
nand U19252 (N_19252,N_16557,N_18534);
nand U19253 (N_19253,N_16700,N_17397);
xnor U19254 (N_19254,N_16651,N_18660);
nand U19255 (N_19255,N_17028,N_16516);
and U19256 (N_19256,N_18306,N_17553);
and U19257 (N_19257,N_17436,N_18654);
nand U19258 (N_19258,N_18725,N_16347);
or U19259 (N_19259,N_16303,N_17599);
nand U19260 (N_19260,N_17920,N_18023);
or U19261 (N_19261,N_17768,N_16562);
nand U19262 (N_19262,N_15960,N_16534);
nand U19263 (N_19263,N_15648,N_17093);
nand U19264 (N_19264,N_16305,N_17577);
nor U19265 (N_19265,N_16791,N_16738);
and U19266 (N_19266,N_17127,N_15817);
nor U19267 (N_19267,N_16896,N_15704);
or U19268 (N_19268,N_18066,N_16758);
nor U19269 (N_19269,N_16744,N_16594);
nor U19270 (N_19270,N_17026,N_16079);
nand U19271 (N_19271,N_18655,N_18468);
and U19272 (N_19272,N_18271,N_17709);
xor U19273 (N_19273,N_17193,N_17949);
or U19274 (N_19274,N_16128,N_16683);
or U19275 (N_19275,N_16371,N_16268);
or U19276 (N_19276,N_16762,N_16550);
and U19277 (N_19277,N_18594,N_17552);
nand U19278 (N_19278,N_17990,N_17921);
and U19279 (N_19279,N_16026,N_15739);
nor U19280 (N_19280,N_16062,N_17217);
nand U19281 (N_19281,N_18347,N_17265);
and U19282 (N_19282,N_17271,N_17973);
nor U19283 (N_19283,N_17687,N_15757);
and U19284 (N_19284,N_16627,N_17275);
nor U19285 (N_19285,N_17121,N_17686);
nor U19286 (N_19286,N_16227,N_16267);
and U19287 (N_19287,N_16365,N_18670);
or U19288 (N_19288,N_18515,N_17728);
and U19289 (N_19289,N_16833,N_18212);
nand U19290 (N_19290,N_18546,N_17753);
nand U19291 (N_19291,N_17135,N_17618);
nand U19292 (N_19292,N_18203,N_17634);
nor U19293 (N_19293,N_15935,N_18448);
nand U19294 (N_19294,N_16041,N_17714);
and U19295 (N_19295,N_16590,N_18656);
and U19296 (N_19296,N_17008,N_18141);
and U19297 (N_19297,N_17716,N_15638);
or U19298 (N_19298,N_17671,N_16325);
xor U19299 (N_19299,N_18202,N_16247);
or U19300 (N_19300,N_18538,N_15709);
nor U19301 (N_19301,N_16478,N_15901);
xor U19302 (N_19302,N_18050,N_18291);
nand U19303 (N_19303,N_17752,N_16364);
or U19304 (N_19304,N_15681,N_16737);
nand U19305 (N_19305,N_16279,N_16704);
nand U19306 (N_19306,N_17587,N_16196);
nand U19307 (N_19307,N_16948,N_17304);
and U19308 (N_19308,N_18719,N_17778);
or U19309 (N_19309,N_16803,N_16832);
nand U19310 (N_19310,N_16620,N_18547);
or U19311 (N_19311,N_16153,N_16373);
and U19312 (N_19312,N_17442,N_18467);
nand U19313 (N_19313,N_16036,N_16451);
and U19314 (N_19314,N_16490,N_17483);
nand U19315 (N_19315,N_17940,N_17231);
nor U19316 (N_19316,N_16435,N_16694);
nor U19317 (N_19317,N_18664,N_17915);
and U19318 (N_19318,N_17816,N_16943);
or U19319 (N_19319,N_18686,N_16326);
nor U19320 (N_19320,N_18327,N_17000);
or U19321 (N_19321,N_16714,N_17379);
and U19322 (N_19322,N_17274,N_16152);
and U19323 (N_19323,N_17648,N_15666);
nor U19324 (N_19324,N_18465,N_18399);
and U19325 (N_19325,N_17120,N_18451);
nor U19326 (N_19326,N_17061,N_18275);
or U19327 (N_19327,N_18698,N_17209);
nand U19328 (N_19328,N_16167,N_17636);
nor U19329 (N_19329,N_15703,N_15745);
and U19330 (N_19330,N_17873,N_16027);
or U19331 (N_19331,N_18371,N_15879);
or U19332 (N_19332,N_17370,N_15942);
nand U19333 (N_19333,N_16787,N_18488);
nor U19334 (N_19334,N_16670,N_17198);
nor U19335 (N_19335,N_17165,N_18741);
nand U19336 (N_19336,N_17605,N_15724);
nand U19337 (N_19337,N_18057,N_18699);
and U19338 (N_19338,N_18070,N_16333);
and U19339 (N_19339,N_18384,N_16246);
and U19340 (N_19340,N_17607,N_17968);
nor U19341 (N_19341,N_17368,N_17846);
and U19342 (N_19342,N_17724,N_18111);
nor U19343 (N_19343,N_17516,N_18580);
and U19344 (N_19344,N_18086,N_16695);
or U19345 (N_19345,N_18119,N_18325);
or U19346 (N_19346,N_15876,N_17306);
xnor U19347 (N_19347,N_16741,N_17653);
or U19348 (N_19348,N_16804,N_15711);
and U19349 (N_19349,N_16690,N_16212);
or U19350 (N_19350,N_16158,N_18063);
nor U19351 (N_19351,N_16257,N_15927);
nor U19352 (N_19352,N_17974,N_16341);
nand U19353 (N_19353,N_16202,N_17312);
and U19354 (N_19354,N_16807,N_17068);
nor U19355 (N_19355,N_17608,N_15980);
nand U19356 (N_19356,N_18645,N_18622);
and U19357 (N_19357,N_16974,N_17010);
nand U19358 (N_19358,N_16183,N_15656);
and U19359 (N_19359,N_17554,N_16352);
or U19360 (N_19360,N_16940,N_16166);
nand U19361 (N_19361,N_17691,N_16171);
nand U19362 (N_19362,N_16187,N_17475);
nand U19363 (N_19363,N_15798,N_16604);
nand U19364 (N_19364,N_18520,N_18669);
xor U19365 (N_19365,N_16038,N_18014);
nand U19366 (N_19366,N_17012,N_17763);
or U19367 (N_19367,N_18718,N_17113);
nand U19368 (N_19368,N_16754,N_17939);
or U19369 (N_19369,N_17732,N_17996);
nand U19370 (N_19370,N_17967,N_17993);
nand U19371 (N_19371,N_18444,N_17302);
or U19372 (N_19372,N_15805,N_18551);
nor U19373 (N_19373,N_17278,N_16898);
nor U19374 (N_19374,N_16934,N_18588);
or U19375 (N_19375,N_15849,N_18370);
nor U19376 (N_19376,N_18317,N_15832);
nor U19377 (N_19377,N_18315,N_18187);
and U19378 (N_19378,N_16668,N_17751);
nand U19379 (N_19379,N_17668,N_17641);
nand U19380 (N_19380,N_18501,N_17879);
nor U19381 (N_19381,N_15766,N_16013);
and U19382 (N_19382,N_17657,N_18062);
and U19383 (N_19383,N_15664,N_16598);
nand U19384 (N_19384,N_17595,N_16397);
or U19385 (N_19385,N_18676,N_17602);
xor U19386 (N_19386,N_16684,N_18364);
nor U19387 (N_19387,N_16823,N_16069);
nand U19388 (N_19388,N_15978,N_16530);
nor U19389 (N_19389,N_16011,N_18176);
xor U19390 (N_19390,N_18367,N_16360);
nor U19391 (N_19391,N_16401,N_16449);
nand U19392 (N_19392,N_15940,N_16138);
or U19393 (N_19393,N_17253,N_18001);
nand U19394 (N_19394,N_16387,N_16391);
nor U19395 (N_19395,N_17781,N_17048);
nor U19396 (N_19396,N_16494,N_16941);
or U19397 (N_19397,N_16457,N_16054);
nand U19398 (N_19398,N_16662,N_16034);
nand U19399 (N_19399,N_17295,N_17877);
nand U19400 (N_19400,N_15800,N_18117);
and U19401 (N_19401,N_16645,N_18579);
nor U19402 (N_19402,N_17140,N_15874);
nand U19403 (N_19403,N_16721,N_16547);
nand U19404 (N_19404,N_16862,N_17427);
and U19405 (N_19405,N_18113,N_17132);
or U19406 (N_19406,N_16308,N_16376);
and U19407 (N_19407,N_17087,N_17220);
or U19408 (N_19408,N_16729,N_17831);
nand U19409 (N_19409,N_16144,N_16565);
and U19410 (N_19410,N_16291,N_17698);
and U19411 (N_19411,N_18365,N_15903);
and U19412 (N_19412,N_16443,N_16657);
nand U19413 (N_19413,N_17050,N_16400);
and U19414 (N_19414,N_17072,N_18192);
nand U19415 (N_19415,N_18693,N_16860);
and U19416 (N_19416,N_18372,N_17682);
or U19417 (N_19417,N_17181,N_18668);
nand U19418 (N_19418,N_18333,N_15802);
nand U19419 (N_19419,N_16962,N_18560);
nor U19420 (N_19420,N_18382,N_18446);
nor U19421 (N_19421,N_17313,N_16510);
and U19422 (N_19422,N_18581,N_17958);
and U19423 (N_19423,N_17178,N_15955);
or U19424 (N_19424,N_16993,N_17588);
and U19425 (N_19425,N_17242,N_16316);
nor U19426 (N_19426,N_15625,N_17431);
xnor U19427 (N_19427,N_17519,N_17695);
nand U19428 (N_19428,N_17556,N_15793);
or U19429 (N_19429,N_17707,N_16906);
and U19430 (N_19430,N_17188,N_15939);
and U19431 (N_19431,N_16573,N_16091);
nand U19432 (N_19432,N_15657,N_17979);
or U19433 (N_19433,N_16615,N_17413);
or U19434 (N_19434,N_17083,N_17629);
nor U19435 (N_19435,N_16652,N_17910);
nand U19436 (N_19436,N_18280,N_18215);
nor U19437 (N_19437,N_17825,N_16603);
or U19438 (N_19438,N_15954,N_15714);
nand U19439 (N_19439,N_17677,N_17479);
or U19440 (N_19440,N_17703,N_17177);
or U19441 (N_19441,N_18300,N_16209);
xnor U19442 (N_19442,N_15740,N_15781);
nor U19443 (N_19443,N_18020,N_17244);
xnor U19444 (N_19444,N_16931,N_18103);
or U19445 (N_19445,N_18724,N_17689);
or U19446 (N_19446,N_17830,N_16760);
or U19447 (N_19447,N_18342,N_17085);
and U19448 (N_19448,N_17115,N_16307);
nor U19449 (N_19449,N_18419,N_18219);
or U19450 (N_19450,N_18431,N_17868);
nand U19451 (N_19451,N_15824,N_16327);
nand U19452 (N_19452,N_18008,N_18128);
and U19453 (N_19453,N_16836,N_18237);
nand U19454 (N_19454,N_17040,N_16165);
and U19455 (N_19455,N_16847,N_17499);
and U19456 (N_19456,N_17023,N_16324);
and U19457 (N_19457,N_16088,N_18127);
or U19458 (N_19458,N_16470,N_15834);
or U19459 (N_19459,N_17740,N_18412);
nor U19460 (N_19460,N_17122,N_18504);
or U19461 (N_19461,N_16853,N_16954);
nand U19462 (N_19462,N_17434,N_15780);
nor U19463 (N_19463,N_18109,N_16219);
nand U19464 (N_19464,N_15898,N_16639);
and U19465 (N_19465,N_16732,N_16298);
nand U19466 (N_19466,N_18225,N_17062);
and U19467 (N_19467,N_16673,N_15639);
or U19468 (N_19468,N_17360,N_17082);
nor U19469 (N_19469,N_18706,N_16731);
nand U19470 (N_19470,N_16792,N_18115);
or U19471 (N_19471,N_16713,N_18616);
nor U19472 (N_19472,N_17100,N_18410);
xnor U19473 (N_19473,N_17490,N_16772);
nor U19474 (N_19474,N_17200,N_18150);
and U19475 (N_19475,N_16484,N_17281);
xnor U19476 (N_19476,N_17092,N_18555);
nor U19477 (N_19477,N_16092,N_17504);
nor U19478 (N_19478,N_16829,N_16122);
or U19479 (N_19479,N_17943,N_17838);
nor U19480 (N_19480,N_16585,N_16419);
or U19481 (N_19481,N_18629,N_16237);
nand U19482 (N_19482,N_16852,N_17916);
or U19483 (N_19483,N_16002,N_16372);
or U19484 (N_19484,N_16958,N_18453);
nor U19485 (N_19485,N_16043,N_18703);
or U19486 (N_19486,N_18620,N_18533);
nor U19487 (N_19487,N_16937,N_16264);
nor U19488 (N_19488,N_18041,N_17524);
or U19489 (N_19489,N_17043,N_17766);
nand U19490 (N_19490,N_16681,N_17670);
nor U19491 (N_19491,N_18612,N_18299);
nand U19492 (N_19492,N_16051,N_16438);
nand U19493 (N_19493,N_15725,N_16386);
or U19494 (N_19494,N_17810,N_17223);
or U19495 (N_19495,N_17006,N_17600);
xor U19496 (N_19496,N_15723,N_16930);
nor U19497 (N_19497,N_16802,N_18107);
nand U19498 (N_19498,N_18196,N_18310);
or U19499 (N_19499,N_17821,N_15753);
nand U19500 (N_19500,N_17667,N_15997);
nor U19501 (N_19501,N_17301,N_17496);
and U19502 (N_19502,N_18734,N_17446);
xor U19503 (N_19503,N_18218,N_15905);
xor U19504 (N_19504,N_17320,N_15670);
nor U19505 (N_19505,N_16154,N_16089);
or U19506 (N_19506,N_16977,N_16524);
nand U19507 (N_19507,N_18172,N_16546);
nand U19508 (N_19508,N_16750,N_17375);
or U19509 (N_19509,N_17583,N_16827);
nand U19510 (N_19510,N_17865,N_15804);
nor U19511 (N_19511,N_18249,N_17952);
xor U19512 (N_19512,N_15692,N_17151);
nor U19513 (N_19513,N_18440,N_17155);
nor U19514 (N_19514,N_18217,N_17738);
or U19515 (N_19515,N_16568,N_16422);
and U19516 (N_19516,N_16112,N_16755);
nand U19517 (N_19517,N_18326,N_16912);
nor U19518 (N_19518,N_17241,N_18232);
nor U19519 (N_19519,N_17470,N_16431);
xor U19520 (N_19520,N_18574,N_17230);
nor U19521 (N_19521,N_17462,N_16952);
nand U19522 (N_19522,N_17106,N_17562);
or U19523 (N_19523,N_16482,N_17272);
xnor U19524 (N_19524,N_15902,N_16723);
nand U19525 (N_19525,N_18733,N_17699);
nor U19526 (N_19526,N_18242,N_16426);
nor U19527 (N_19527,N_17111,N_17520);
and U19528 (N_19528,N_15641,N_16812);
xnor U19529 (N_19529,N_17679,N_16831);
nor U19530 (N_19530,N_17388,N_16555);
nor U19531 (N_19531,N_17985,N_16491);
or U19532 (N_19532,N_18051,N_18689);
and U19533 (N_19533,N_16107,N_15914);
nor U19534 (N_19534,N_18572,N_18517);
or U19535 (N_19535,N_16999,N_18120);
and U19536 (N_19536,N_18666,N_17219);
and U19537 (N_19537,N_16198,N_16135);
or U19538 (N_19538,N_17014,N_18457);
xnor U19539 (N_19539,N_17226,N_17972);
or U19540 (N_19540,N_18565,N_16920);
or U19541 (N_19541,N_17029,N_15878);
and U19542 (N_19542,N_18213,N_17316);
nor U19543 (N_19543,N_18243,N_18164);
or U19544 (N_19544,N_17638,N_16767);
and U19545 (N_19545,N_17889,N_16586);
nor U19546 (N_19546,N_16076,N_15818);
nand U19547 (N_19547,N_16886,N_17749);
nor U19548 (N_19548,N_18596,N_16793);
nand U19549 (N_19549,N_17758,N_16056);
and U19550 (N_19550,N_16140,N_17189);
nand U19551 (N_19551,N_18466,N_18613);
nor U19552 (N_19552,N_16676,N_17924);
nor U19553 (N_19553,N_17845,N_15685);
and U19554 (N_19554,N_15938,N_16797);
nand U19555 (N_19555,N_18085,N_15702);
nor U19556 (N_19556,N_16837,N_15982);
or U19557 (N_19557,N_16340,N_16656);
nand U19558 (N_19558,N_17134,N_16053);
nand U19559 (N_19559,N_16123,N_16117);
or U19560 (N_19560,N_15850,N_16423);
and U19561 (N_19561,N_15762,N_18177);
and U19562 (N_19562,N_17334,N_17571);
or U19563 (N_19563,N_15642,N_15748);
nand U19564 (N_19564,N_18009,N_16871);
nand U19565 (N_19565,N_16591,N_16743);
nor U19566 (N_19566,N_16162,N_18330);
nand U19567 (N_19567,N_16115,N_18680);
nor U19568 (N_19568,N_17429,N_17287);
and U19569 (N_19569,N_18036,N_17560);
or U19570 (N_19570,N_17069,N_18578);
and U19571 (N_19571,N_15929,N_16549);
or U19572 (N_19572,N_17346,N_16933);
or U19573 (N_19573,N_17997,N_17678);
and U19574 (N_19574,N_17168,N_16633);
nor U19575 (N_19575,N_17833,N_15897);
nand U19576 (N_19576,N_18191,N_16336);
nand U19577 (N_19577,N_18091,N_18209);
nand U19578 (N_19578,N_17660,N_17243);
nor U19579 (N_19579,N_17297,N_16052);
nor U19580 (N_19580,N_17478,N_15887);
or U19581 (N_19581,N_16244,N_16819);
or U19582 (N_19582,N_17158,N_17366);
nand U19583 (N_19583,N_17038,N_15952);
and U19584 (N_19584,N_17899,N_18321);
and U19585 (N_19585,N_17042,N_17812);
and U19586 (N_19586,N_17204,N_15990);
and U19587 (N_19587,N_15746,N_16588);
or U19588 (N_19588,N_18522,N_17461);
or U19589 (N_19589,N_18662,N_17850);
and U19590 (N_19590,N_18499,N_17882);
nor U19591 (N_19591,N_18208,N_17779);
nor U19592 (N_19592,N_18599,N_17324);
and U19593 (N_19593,N_16223,N_17495);
nor U19594 (N_19594,N_18194,N_18130);
nor U19595 (N_19595,N_17819,N_16368);
nand U19596 (N_19596,N_18039,N_18646);
and U19597 (N_19597,N_17611,N_17737);
or U19598 (N_19598,N_15989,N_16778);
and U19599 (N_19599,N_18324,N_18185);
or U19600 (N_19600,N_16465,N_18031);
xor U19601 (N_19601,N_17917,N_18292);
nor U19602 (N_19602,N_15868,N_18264);
nand U19603 (N_19603,N_18391,N_17330);
nand U19604 (N_19604,N_17133,N_17881);
nor U19605 (N_19605,N_16922,N_16213);
and U19606 (N_19606,N_17971,N_17136);
nand U19607 (N_19607,N_18459,N_17511);
xor U19608 (N_19608,N_18397,N_17386);
and U19609 (N_19609,N_17237,N_16600);
and U19610 (N_19610,N_17175,N_17572);
and U19611 (N_19611,N_16542,N_17031);
nor U19612 (N_19612,N_17146,N_16024);
nand U19613 (N_19613,N_17147,N_16012);
or U19614 (N_19614,N_18687,N_17900);
nor U19615 (N_19615,N_16511,N_18161);
nand U19616 (N_19616,N_17521,N_16808);
nor U19617 (N_19617,N_16339,N_16584);
or U19618 (N_19618,N_18583,N_17930);
or U19619 (N_19619,N_18691,N_18701);
nand U19620 (N_19620,N_16506,N_15768);
nand U19621 (N_19621,N_17832,N_16178);
and U19622 (N_19622,N_16182,N_16987);
nor U19623 (N_19623,N_17664,N_17937);
and U19624 (N_19624,N_16706,N_18626);
and U19625 (N_19625,N_17510,N_17339);
xor U19626 (N_19626,N_17255,N_18568);
nand U19627 (N_19627,N_16503,N_17094);
nand U19628 (N_19628,N_16959,N_16469);
nor U19629 (N_19629,N_16965,N_16356);
and U19630 (N_19630,N_17650,N_15862);
or U19631 (N_19631,N_16806,N_18348);
nand U19632 (N_19632,N_16605,N_18585);
nor U19633 (N_19633,N_16277,N_16370);
nor U19634 (N_19634,N_17932,N_17992);
and U19635 (N_19635,N_16348,N_17408);
nor U19636 (N_19636,N_18228,N_17123);
or U19637 (N_19637,N_18447,N_15721);
nor U19638 (N_19638,N_17551,N_16865);
nand U19639 (N_19639,N_16381,N_17245);
and U19640 (N_19640,N_17820,N_17325);
and U19641 (N_19641,N_17918,N_18183);
and U19642 (N_19642,N_15974,N_17246);
nand U19643 (N_19643,N_17533,N_17187);
or U19644 (N_19644,N_18282,N_16640);
nand U19645 (N_19645,N_17414,N_18738);
nand U19646 (N_19646,N_18528,N_16184);
nand U19647 (N_19647,N_18427,N_15845);
nand U19648 (N_19648,N_15686,N_16214);
nor U19649 (N_19649,N_18562,N_18090);
or U19650 (N_19650,N_16210,N_16003);
nand U19651 (N_19651,N_15917,N_17144);
nor U19652 (N_19652,N_16084,N_17721);
nor U19653 (N_19653,N_17978,N_17897);
nand U19654 (N_19654,N_15841,N_17371);
xnor U19655 (N_19655,N_17293,N_16217);
nand U19656 (N_19656,N_17957,N_17405);
nand U19657 (N_19657,N_18518,N_17075);
nor U19658 (N_19658,N_15906,N_17469);
nor U19659 (N_19659,N_16923,N_16968);
and U19660 (N_19660,N_17114,N_17046);
xor U19661 (N_19661,N_15680,N_18635);
and U19662 (N_19662,N_17931,N_18366);
nor U19663 (N_19663,N_18523,N_16351);
or U19664 (N_19664,N_18112,N_16939);
and U19665 (N_19665,N_16284,N_18423);
nand U19666 (N_19666,N_17964,N_18190);
and U19667 (N_19667,N_17847,N_17173);
nor U19668 (N_19668,N_17522,N_15773);
nor U19669 (N_19669,N_18747,N_15731);
xnor U19670 (N_19670,N_16766,N_18134);
nor U19671 (N_19671,N_18632,N_16671);
nor U19672 (N_19672,N_17474,N_17089);
and U19673 (N_19673,N_18077,N_16446);
xor U19674 (N_19674,N_17143,N_17007);
nor U19675 (N_19675,N_15673,N_18234);
nand U19676 (N_19676,N_18211,N_16795);
or U19677 (N_19677,N_18653,N_17683);
nand U19678 (N_19678,N_18244,N_18084);
nand U19679 (N_19679,N_16844,N_17863);
nor U19680 (N_19680,N_17809,N_17770);
xor U19681 (N_19681,N_16248,N_18303);
nand U19682 (N_19682,N_18651,N_15637);
and U19683 (N_19683,N_16880,N_16746);
and U19684 (N_19684,N_15858,N_18312);
or U19685 (N_19685,N_18601,N_16362);
nor U19686 (N_19686,N_18380,N_16776);
and U19687 (N_19687,N_15775,N_17035);
nand U19688 (N_19688,N_18454,N_17268);
xor U19689 (N_19689,N_18261,N_16813);
nor U19690 (N_19690,N_17885,N_16177);
and U19691 (N_19691,N_16338,N_15985);
and U19692 (N_19692,N_18500,N_16523);
nor U19693 (N_19693,N_15729,N_17221);
xor U19694 (N_19694,N_15840,N_18248);
and U19695 (N_19695,N_18293,N_16207);
and U19696 (N_19696,N_17959,N_17322);
or U19697 (N_19697,N_17969,N_17545);
nand U19698 (N_19698,N_17417,N_15975);
nand U19699 (N_19699,N_16556,N_18267);
nor U19700 (N_19700,N_18618,N_18040);
nor U19701 (N_19701,N_15830,N_16740);
nand U19702 (N_19702,N_18537,N_17247);
xnor U19703 (N_19703,N_18221,N_15778);
nand U19704 (N_19704,N_17167,N_16956);
or U19705 (N_19705,N_16230,N_17105);
nand U19706 (N_19706,N_16985,N_15984);
nand U19707 (N_19707,N_17137,N_15691);
or U19708 (N_19708,N_16160,N_15870);
nand U19709 (N_19709,N_17015,N_16411);
and U19710 (N_19710,N_16440,N_18486);
or U19711 (N_19711,N_17372,N_18356);
nor U19712 (N_19712,N_15655,N_17056);
or U19713 (N_19713,N_16168,N_18340);
nand U19714 (N_19714,N_16822,N_17466);
or U19715 (N_19715,N_17886,N_18129);
nand U19716 (N_19716,N_17169,N_18026);
nand U19717 (N_19717,N_16825,N_17179);
nor U19718 (N_19718,N_17693,N_17674);
or U19719 (N_19719,N_16260,N_17152);
nand U19720 (N_19720,N_15866,N_17463);
nand U19721 (N_19721,N_16771,N_16885);
or U19722 (N_19722,N_17369,N_16978);
or U19723 (N_19723,N_16587,N_16060);
or U19724 (N_19724,N_18320,N_18571);
nor U19725 (N_19725,N_17045,N_16720);
and U19726 (N_19726,N_18527,N_15632);
and U19727 (N_19727,N_16810,N_15892);
xor U19728 (N_19728,N_18443,N_17084);
and U19729 (N_19729,N_16519,N_17383);
and U19730 (N_19730,N_15693,N_17385);
nand U19731 (N_19731,N_17700,N_17044);
nor U19732 (N_19732,N_17070,N_16916);
nor U19733 (N_19733,N_16176,N_17760);
nor U19734 (N_19734,N_17239,N_15783);
xnor U19735 (N_19735,N_17644,N_18089);
or U19736 (N_19736,N_16163,N_17862);
xnor U19737 (N_19737,N_15633,N_15705);
and U19738 (N_19738,N_18059,N_18471);
nor U19739 (N_19739,N_18272,N_15770);
nor U19740 (N_19740,N_15779,N_16406);
and U19741 (N_19741,N_17950,N_18390);
or U19742 (N_19742,N_18049,N_18566);
and U19743 (N_19743,N_16870,N_15988);
nor U19744 (N_19744,N_15634,N_16863);
nand U19745 (N_19745,N_17767,N_17904);
and U19746 (N_19746,N_16909,N_16129);
or U19747 (N_19747,N_16414,N_17164);
nor U19748 (N_19748,N_16575,N_18289);
xnor U19749 (N_19749,N_17389,N_18102);
nand U19750 (N_19750,N_17454,N_16047);
xnor U19751 (N_19751,N_16975,N_15751);
nand U19752 (N_19752,N_18624,N_16374);
xor U19753 (N_19753,N_16835,N_17201);
nor U19754 (N_19754,N_17941,N_18536);
nor U19755 (N_19755,N_16141,N_16354);
nor U19756 (N_19756,N_18462,N_16363);
nand U19757 (N_19757,N_15912,N_16439);
or U19758 (N_19758,N_17797,N_16945);
nor U19759 (N_19759,N_17103,N_15875);
nand U19760 (N_19760,N_15672,N_15683);
and U19761 (N_19761,N_15697,N_17349);
nor U19762 (N_19762,N_18587,N_17632);
and U19763 (N_19763,N_17225,N_17801);
nor U19764 (N_19764,N_18016,N_17101);
or U19765 (N_19765,N_16614,N_15643);
or U19766 (N_19766,N_17813,N_16320);
nand U19767 (N_19767,N_18018,N_18679);
xnor U19768 (N_19768,N_16846,N_18395);
and U19769 (N_19769,N_18239,N_16625);
or U19770 (N_19770,N_16471,N_17944);
or U19771 (N_19771,N_15720,N_17004);
and U19772 (N_19772,N_18593,N_15931);
nand U19773 (N_19773,N_15741,N_16137);
nor U19774 (N_19774,N_17684,N_18216);
or U19775 (N_19775,N_17443,N_17576);
and U19776 (N_19776,N_17185,N_17416);
and U19777 (N_19777,N_17501,N_17874);
nand U19778 (N_19778,N_15676,N_15688);
or U19779 (N_19779,N_16269,N_16972);
nand U19780 (N_19780,N_15794,N_18162);
nand U19781 (N_19781,N_17649,N_18030);
xnor U19782 (N_19782,N_18381,N_16288);
nand U19783 (N_19783,N_16057,N_16459);
nand U19784 (N_19784,N_16629,N_17946);
and U19785 (N_19785,N_17337,N_16709);
nor U19786 (N_19786,N_15831,N_17718);
and U19787 (N_19787,N_18386,N_18606);
and U19788 (N_19788,N_18659,N_17426);
nand U19789 (N_19789,N_18461,N_18377);
and U19790 (N_19790,N_18605,N_18072);
and U19791 (N_19791,N_18220,N_18076);
and U19792 (N_19792,N_17117,N_17933);
nand U19793 (N_19793,N_16170,N_17710);
and U19794 (N_19794,N_18147,N_18569);
and U19795 (N_19795,N_16989,N_17183);
nand U19796 (N_19796,N_18279,N_16228);
nor U19797 (N_19797,N_18189,N_17839);
or U19798 (N_19798,N_15689,N_17574);
and U19799 (N_19799,N_17544,N_17756);
xor U19800 (N_19800,N_17536,N_16826);
nand U19801 (N_19801,N_17424,N_16518);
and U19802 (N_19802,N_17252,N_17359);
nor U19803 (N_19803,N_18492,N_17869);
nand U19804 (N_19804,N_17712,N_17172);
nand U19805 (N_19805,N_18301,N_16039);
or U19806 (N_19806,N_15838,N_18433);
or U19807 (N_19807,N_16904,N_16385);
nand U19808 (N_19808,N_18708,N_16967);
nor U19809 (N_19809,N_16493,N_15796);
nand U19810 (N_19810,N_18313,N_16601);
or U19811 (N_19811,N_16892,N_16921);
and U19812 (N_19812,N_15822,N_16606);
or U19813 (N_19813,N_17348,N_18024);
or U19814 (N_19814,N_16393,N_18374);
nand U19815 (N_19815,N_17994,N_16592);
nand U19816 (N_19816,N_16020,N_16313);
and U19817 (N_19817,N_17376,N_17328);
or U19818 (N_19818,N_16432,N_15923);
nand U19819 (N_19819,N_17471,N_18685);
xnor U19820 (N_19820,N_17338,N_15727);
nor U19821 (N_19821,N_16080,N_15712);
and U19822 (N_19822,N_17962,N_16703);
nor U19823 (N_19823,N_17590,N_17557);
and U19824 (N_19824,N_17891,N_17685);
or U19825 (N_19825,N_18092,N_18479);
xor U19826 (N_19826,N_16330,N_17828);
or U19827 (N_19827,N_17876,N_16984);
and U19828 (N_19828,N_17880,N_17834);
and U19829 (N_19829,N_16976,N_18224);
or U19830 (N_19830,N_17382,N_15777);
nand U19831 (N_19831,N_17256,N_15904);
or U19832 (N_19832,N_17033,N_17569);
and U19833 (N_19833,N_17575,N_17609);
or U19834 (N_19834,N_16894,N_16017);
and U19835 (N_19835,N_17190,N_16500);
and U19836 (N_19836,N_17064,N_16201);
or U19837 (N_19837,N_16329,N_17656);
and U19838 (N_19838,N_18415,N_16612);
nor U19839 (N_19839,N_16405,N_17987);
and U19840 (N_19840,N_17003,N_16707);
nand U19841 (N_19841,N_17261,N_16143);
nor U19842 (N_19842,N_16907,N_18592);
xor U19843 (N_19843,N_17720,N_16951);
xnor U19844 (N_19844,N_17250,N_18497);
nor U19845 (N_19845,N_18549,N_16786);
nand U19846 (N_19846,N_17159,N_18193);
or U19847 (N_19847,N_15696,N_17336);
xor U19848 (N_19848,N_16096,N_17394);
xor U19849 (N_19849,N_18351,N_16164);
and U19850 (N_19850,N_15926,N_15910);
nand U19851 (N_19851,N_18336,N_17827);
or U19852 (N_19852,N_17731,N_16551);
and U19853 (N_19853,N_17558,N_16025);
or U19854 (N_19854,N_18363,N_18445);
nand U19855 (N_19855,N_15790,N_17539);
xor U19856 (N_19856,N_15925,N_16711);
or U19857 (N_19857,N_16641,N_15674);
or U19858 (N_19858,N_17150,N_16495);
or U19859 (N_19859,N_16589,N_17283);
or U19860 (N_19860,N_16817,N_18673);
nand U19861 (N_19861,N_18053,N_16009);
or U19862 (N_19862,N_17310,N_16537);
nor U19863 (N_19863,N_15772,N_18505);
nor U19864 (N_19864,N_16535,N_16000);
and U19865 (N_19865,N_18253,N_18434);
nand U19866 (N_19866,N_16388,N_15963);
nor U19867 (N_19867,N_17815,N_15847);
nor U19868 (N_19868,N_15964,N_17485);
xnor U19869 (N_19869,N_16266,N_15967);
nand U19870 (N_19870,N_18704,N_18133);
and U19871 (N_19871,N_17991,N_17814);
nor U19872 (N_19872,N_16146,N_15936);
xnor U19873 (N_19873,N_16389,N_15629);
and U19874 (N_19874,N_17955,N_17563);
nor U19875 (N_19875,N_17362,N_17923);
nor U19876 (N_19876,N_15861,N_17350);
nand U19877 (N_19877,N_16243,N_17642);
or U19878 (N_19878,N_18650,N_18144);
nand U19879 (N_19879,N_17273,N_15726);
or U19880 (N_19880,N_17203,N_18711);
nor U19881 (N_19881,N_18553,N_15767);
nand U19882 (N_19882,N_16120,N_17888);
or U19883 (N_19883,N_17335,N_18663);
nor U19884 (N_19884,N_18564,N_15921);
and U19885 (N_19885,N_17465,N_16350);
and U19886 (N_19886,N_18490,N_18469);
nand U19887 (N_19887,N_15918,N_16169);
nand U19888 (N_19888,N_18508,N_17628);
or U19889 (N_19889,N_16258,N_17051);
and U19890 (N_19890,N_17259,N_15661);
or U19891 (N_19891,N_17163,N_16234);
xor U19892 (N_19892,N_18408,N_16980);
or U19893 (N_19893,N_15814,N_18652);
and U19894 (N_19894,N_17396,N_18589);
nand U19895 (N_19895,N_17594,N_16654);
nor U19896 (N_19896,N_17584,N_16358);
nand U19897 (N_19897,N_17440,N_17661);
nand U19898 (N_19898,N_16749,N_18309);
nand U19899 (N_19899,N_17690,N_18323);
xnor U19900 (N_19900,N_17421,N_16728);
nand U19901 (N_19901,N_17468,N_16905);
nand U19902 (N_19902,N_16595,N_15992);
nand U19903 (N_19903,N_18011,N_15752);
or U19904 (N_19904,N_16563,N_18238);
nand U19905 (N_19905,N_16173,N_17141);
nand U19906 (N_19906,N_15986,N_15713);
and U19907 (N_19907,N_18430,N_16621);
nand U19908 (N_19908,N_15728,N_16499);
nand U19909 (N_19909,N_16218,N_16008);
or U19910 (N_19910,N_16028,N_15941);
nand U19911 (N_19911,N_16251,N_17267);
and U19912 (N_19912,N_16751,N_17216);
or U19913 (N_19913,N_15973,N_16355);
nand U19914 (N_19914,N_18263,N_16240);
or U19915 (N_19915,N_16382,N_17901);
or U19916 (N_19916,N_16841,N_18151);
nand U19917 (N_19917,N_17942,N_16071);
or U19918 (N_19918,N_15801,N_16624);
or U19919 (N_19919,N_16380,N_18441);
or U19920 (N_19920,N_18270,N_17422);
or U19921 (N_19921,N_15647,N_17254);
nand U19922 (N_19922,N_17482,N_18201);
nand U19923 (N_19923,N_16881,N_17919);
or U19924 (N_19924,N_16517,N_17719);
nor U19925 (N_19925,N_18158,N_17925);
and U19926 (N_19926,N_16879,N_16911);
or U19927 (N_19927,N_16902,N_15869);
and U19928 (N_19928,N_17438,N_18006);
and U19929 (N_19929,N_18297,N_17579);
or U19930 (N_19930,N_16698,N_18338);
or U19931 (N_19931,N_16195,N_15718);
or U19932 (N_19932,N_16412,N_15677);
nor U19933 (N_19933,N_16220,N_18353);
and U19934 (N_19934,N_16834,N_16083);
or U19935 (N_19935,N_18082,N_16736);
nor U19936 (N_19936,N_17199,N_16650);
nand U19937 (N_19937,N_16724,N_16292);
nand U19938 (N_19938,N_17723,N_17131);
nor U19939 (N_19939,N_16124,N_16127);
and U19940 (N_19940,N_18067,N_16675);
nand U19941 (N_19941,N_18186,N_17697);
and U19942 (N_19942,N_17130,N_16596);
nor U19943 (N_19943,N_17224,N_16413);
and U19944 (N_19944,N_18179,N_17975);
nor U19945 (N_19945,N_18101,N_16048);
nor U19946 (N_19946,N_17450,N_18088);
nor U19947 (N_19947,N_16666,N_16780);
nand U19948 (N_19948,N_16525,N_15896);
or U19949 (N_19949,N_17741,N_16211);
nor U19950 (N_19950,N_18712,N_18311);
nor U19951 (N_19951,N_15827,N_17633);
or U19952 (N_19952,N_16901,N_18634);
and U19953 (N_19953,N_17513,N_16345);
nand U19954 (N_19954,N_18083,N_17842);
and U19955 (N_19955,N_16276,N_17124);
and U19956 (N_19956,N_17894,N_16130);
nor U19957 (N_19957,N_18688,N_17567);
nor U19958 (N_19958,N_17318,N_17843);
nand U19959 (N_19959,N_18073,N_18507);
nor U19960 (N_19960,N_17161,N_16072);
nand U19961 (N_19961,N_18295,N_17844);
nand U19962 (N_19962,N_16014,N_17784);
nor U19963 (N_19963,N_15881,N_18149);
or U19964 (N_19964,N_16301,N_18474);
or U19965 (N_19965,N_17659,N_15981);
nand U19966 (N_19966,N_17315,N_18296);
and U19967 (N_19967,N_18173,N_16722);
and U19968 (N_19968,N_18636,N_16674);
and U19969 (N_19969,N_18106,N_17412);
nor U19970 (N_19970,N_17769,N_17612);
nand U19971 (N_19971,N_18285,N_18145);
or U19972 (N_19972,N_18409,N_16145);
or U19973 (N_19973,N_16185,N_17603);
nor U19974 (N_19974,N_17024,N_17982);
nand U19975 (N_19975,N_18210,N_16367);
nand U19976 (N_19976,N_16453,N_17782);
or U19977 (N_19977,N_15786,N_17811);
nand U19978 (N_19978,N_15983,N_16252);
and U19979 (N_19979,N_17598,N_16087);
or U19980 (N_19980,N_18607,N_18644);
and U19981 (N_19981,N_17725,N_17097);
nand U19982 (N_19982,N_18481,N_16680);
and U19983 (N_19983,N_15958,N_16867);
and U19984 (N_19984,N_16855,N_18108);
and U19985 (N_19985,N_16480,N_18483);
and U19986 (N_19986,N_17635,N_17472);
and U19987 (N_19987,N_17423,N_17537);
xor U19988 (N_19988,N_16467,N_16065);
and U19989 (N_19989,N_18702,N_16864);
and U19990 (N_19990,N_18642,N_18514);
xnor U19991 (N_19991,N_16764,N_17547);
and U19992 (N_19992,N_17098,N_18329);
or U19993 (N_19993,N_17409,N_16433);
xnor U19994 (N_19994,N_15934,N_16607);
xor U19995 (N_19995,N_15631,N_15970);
or U19996 (N_19996,N_15994,N_18022);
or U19997 (N_19997,N_18188,N_17049);
and U19998 (N_19998,N_17277,N_15650);
or U19999 (N_19999,N_17503,N_17711);
nor U20000 (N_20000,N_16782,N_15843);
and U20001 (N_20001,N_18690,N_16796);
or U20002 (N_20002,N_17759,N_16947);
and U20003 (N_20003,N_17540,N_17453);
xor U20004 (N_20004,N_17214,N_16021);
or U20005 (N_20005,N_16925,N_17798);
nor U20006 (N_20006,N_17444,N_15948);
or U20007 (N_20007,N_17060,N_17704);
or U20008 (N_20008,N_17694,N_17286);
nand U20009 (N_20009,N_17864,N_18464);
or U20010 (N_20010,N_17411,N_16074);
nand U20011 (N_20011,N_16108,N_16199);
nor U20012 (N_20012,N_17981,N_17138);
nor U20013 (N_20013,N_17773,N_16843);
nor U20014 (N_20014,N_17378,N_15665);
and U20015 (N_20015,N_16425,N_16861);
and U20016 (N_20016,N_17750,N_16950);
nor U20017 (N_20017,N_16357,N_17307);
nand U20018 (N_20018,N_17456,N_17032);
and U20019 (N_20019,N_17314,N_17909);
and U20020 (N_20020,N_18276,N_15684);
and U20021 (N_20021,N_18717,N_17373);
nor U20022 (N_20022,N_16109,N_15873);
nand U20023 (N_20023,N_15949,N_16222);
nand U20024 (N_20024,N_17420,N_16638);
and U20025 (N_20025,N_17836,N_16346);
and U20026 (N_20026,N_18610,N_15828);
or U20027 (N_20027,N_18029,N_16255);
nand U20028 (N_20028,N_16005,N_18171);
or U20029 (N_20029,N_17139,N_18658);
nand U20030 (N_20030,N_17747,N_16669);
and U20031 (N_20031,N_16045,N_15662);
or U20032 (N_20032,N_16717,N_16473);
nor U20033 (N_20033,N_16858,N_17213);
nand U20034 (N_20034,N_16272,N_16106);
or U20035 (N_20035,N_17327,N_16066);
and U20036 (N_20036,N_16608,N_18226);
or U20037 (N_20037,N_17905,N_17903);
and U20038 (N_20038,N_15627,N_18319);
and U20039 (N_20039,N_17681,N_15821);
nand U20040 (N_20040,N_16253,N_17855);
nor U20041 (N_20041,N_17755,N_17822);
nand U20042 (N_20042,N_18539,N_16361);
nand U20043 (N_20043,N_17263,N_17041);
nor U20044 (N_20044,N_16029,N_16769);
xor U20045 (N_20045,N_16616,N_18411);
or U20046 (N_20046,N_16063,N_17596);
or U20047 (N_20047,N_17858,N_16768);
nand U20048 (N_20048,N_17340,N_17745);
or U20049 (N_20049,N_17145,N_17525);
xor U20050 (N_20050,N_18157,N_17079);
and U20051 (N_20051,N_18142,N_17433);
nand U20052 (N_20052,N_16583,N_17564);
nor U20053 (N_20053,N_16119,N_17912);
or U20054 (N_20054,N_16444,N_18350);
nor U20055 (N_20055,N_18054,N_15829);
nor U20056 (N_20056,N_16667,N_18554);
xor U20057 (N_20057,N_17439,N_15792);
nor U20058 (N_20058,N_17458,N_15947);
and U20059 (N_20059,N_17361,N_18535);
nor U20060 (N_20060,N_17875,N_16799);
nor U20061 (N_20061,N_17451,N_18530);
and U20062 (N_20062,N_16942,N_16630);
nand U20063 (N_20063,N_17546,N_17380);
nor U20064 (N_20064,N_15808,N_17800);
or U20065 (N_20065,N_18003,N_16377);
and U20066 (N_20066,N_17872,N_15848);
and U20067 (N_20067,N_16821,N_18137);
and U20068 (N_20068,N_16116,N_18422);
xnor U20069 (N_20069,N_16498,N_15919);
nand U20070 (N_20070,N_18287,N_18404);
or U20071 (N_20071,N_17878,N_18240);
or U20072 (N_20072,N_18257,N_17541);
nor U20073 (N_20073,N_18094,N_16294);
and U20074 (N_20074,N_15928,N_17861);
nand U20075 (N_20075,N_16679,N_17235);
or U20076 (N_20076,N_17792,N_16891);
xor U20077 (N_20077,N_18080,N_16427);
nor U20078 (N_20078,N_17530,N_18060);
or U20079 (N_20079,N_17486,N_15791);
or U20080 (N_20080,N_16653,N_16599);
and U20081 (N_20081,N_16093,N_17428);
nor U20082 (N_20082,N_17202,N_16125);
xnor U20083 (N_20083,N_16917,N_17675);
nor U20084 (N_20084,N_16982,N_18631);
nor U20085 (N_20085,N_17500,N_16417);
nand U20086 (N_20086,N_18630,N_16763);
nor U20087 (N_20087,N_16748,N_18245);
nand U20088 (N_20088,N_17785,N_16097);
and U20089 (N_20089,N_16678,N_16617);
nand U20090 (N_20090,N_16571,N_16233);
nor U20091 (N_20091,N_15640,N_17804);
and U20092 (N_20092,N_17205,N_16067);
or U20093 (N_20093,N_16042,N_16682);
nand U20094 (N_20094,N_16100,N_16988);
nand U20095 (N_20095,N_17591,N_17555);
nand U20096 (N_20096,N_18604,N_16811);
nor U20097 (N_20097,N_15907,N_16908);
and U20098 (N_20098,N_18509,N_17067);
nand U20099 (N_20099,N_18017,N_16262);
xnor U20100 (N_20100,N_15698,N_18204);
nor U20101 (N_20101,N_17914,N_16938);
nand U20102 (N_20102,N_16460,N_15760);
and U20103 (N_20103,N_16895,N_16696);
or U20104 (N_20104,N_16448,N_18600);
and U20105 (N_20105,N_17228,N_16623);
or U20106 (N_20106,N_15669,N_18125);
nor U20107 (N_20107,N_18531,N_16428);
nor U20108 (N_20108,N_18674,N_16991);
nor U20109 (N_20109,N_16418,N_18081);
and U20110 (N_20110,N_17826,N_18328);
and U20111 (N_20111,N_16777,N_17019);
or U20112 (N_20112,N_17276,N_17039);
nor U20113 (N_20113,N_16293,N_16554);
and U20114 (N_20114,N_16442,N_16632);
or U20115 (N_20115,N_15667,N_17961);
and U20116 (N_20116,N_18068,N_16574);
and U20117 (N_20117,N_18010,N_18715);
nand U20118 (N_20118,N_17234,N_16476);
nand U20119 (N_20119,N_18561,N_16064);
or U20120 (N_20120,N_17998,N_18255);
or U20121 (N_20121,N_18198,N_17859);
nand U20122 (N_20122,N_17531,N_15852);
or U20123 (N_20123,N_16452,N_18621);
nor U20124 (N_20124,N_15908,N_16270);
nor U20125 (N_20125,N_17351,N_16424);
or U20126 (N_20126,N_18004,N_15959);
xnor U20127 (N_20127,N_18744,N_16963);
or U20128 (N_20128,N_16869,N_18139);
and U20129 (N_20129,N_18628,N_16953);
nand U20130 (N_20130,N_17488,N_18165);
and U20131 (N_20131,N_18602,N_17418);
and U20132 (N_20132,N_16774,N_16850);
xor U20133 (N_20133,N_18156,N_18227);
nand U20134 (N_20134,N_18709,N_17746);
or U20135 (N_20135,N_16635,N_18576);
nor U20136 (N_20136,N_17425,N_16238);
xnor U20137 (N_20137,N_17806,N_16148);
or U20138 (N_20138,N_17791,N_16915);
or U20139 (N_20139,N_16569,N_18619);
nand U20140 (N_20140,N_15962,N_18316);
nor U20141 (N_20141,N_18456,N_15995);
nand U20142 (N_20142,N_18058,N_16349);
nand U20143 (N_20143,N_15671,N_15734);
nor U20144 (N_20144,N_18273,N_15719);
nand U20145 (N_20145,N_16996,N_16396);
or U20146 (N_20146,N_16644,N_16946);
or U20147 (N_20147,N_18104,N_17282);
or U20148 (N_20148,N_16466,N_17922);
nor U20149 (N_20149,N_17736,N_18661);
or U20150 (N_20150,N_18154,N_17647);
and U20151 (N_20151,N_18614,N_15694);
and U20152 (N_20152,N_16070,N_17091);
nor U20153 (N_20153,N_18695,N_16702);
nor U20154 (N_20154,N_15979,N_17053);
and U20155 (N_20155,N_15700,N_17652);
or U20156 (N_20156,N_16394,N_16359);
or U20157 (N_20157,N_16814,N_16658);
nor U20158 (N_20158,N_18543,N_18258);
nand U20159 (N_20159,N_16966,N_16688);
nand U20160 (N_20160,N_15969,N_17430);
nand U20161 (N_20161,N_18163,N_18584);
nor U20162 (N_20162,N_17713,N_17578);
nor U20163 (N_20163,N_18557,N_18358);
nand U20164 (N_20164,N_18639,N_16312);
nor U20165 (N_20165,N_17593,N_18259);
and U20166 (N_20166,N_17517,N_16875);
xor U20167 (N_20167,N_16659,N_17057);
nand U20168 (N_20168,N_17445,N_17036);
nor U20169 (N_20169,N_17356,N_17743);
or U20170 (N_20170,N_16315,N_17871);
xor U20171 (N_20171,N_17818,N_15920);
or U20172 (N_20172,N_17400,N_17624);
and U20173 (N_20173,N_16022,N_17748);
nand U20174 (N_20174,N_16142,N_16512);
or U20175 (N_20175,N_18608,N_17951);
or U20176 (N_20176,N_16283,N_18262);
nand U20177 (N_20177,N_17639,N_17493);
and U20178 (N_20178,N_15933,N_18429);
nand U20179 (N_20179,N_16566,N_17480);
or U20180 (N_20180,N_17586,N_15953);
or U20181 (N_20181,N_15977,N_17229);
and U20182 (N_20182,N_16379,N_16699);
nor U20183 (N_20183,N_15743,N_17047);
or U20184 (N_20184,N_17643,N_18069);
nor U20185 (N_20185,N_18728,N_18615);
nand U20186 (N_20186,N_15756,N_16044);
or U20187 (N_20187,N_17326,N_18575);
nor U20188 (N_20188,N_15916,N_18428);
nand U20189 (N_20189,N_16286,N_16180);
and U20190 (N_20190,N_17303,N_16319);
nor U20191 (N_20191,N_17945,N_17215);
nand U20192 (N_20192,N_16046,N_16986);
nand U20193 (N_20193,N_15971,N_18524);
nand U20194 (N_20194,N_18155,N_16718);
nor U20195 (N_20195,N_17222,N_17407);
nor U20196 (N_20196,N_17099,N_15759);
or U20197 (N_20197,N_15771,N_17066);
or U20198 (N_20198,N_17294,N_18229);
nor U20199 (N_20199,N_17088,N_17883);
nor U20200 (N_20200,N_17908,N_16032);
or U20201 (N_20201,N_16756,N_16691);
xnor U20202 (N_20202,N_17666,N_15699);
nor U20203 (N_20203,N_15877,N_16231);
nand U20204 (N_20204,N_17585,N_15708);
or U20205 (N_20205,N_18166,N_17658);
nor U20206 (N_20206,N_17108,N_17926);
nand U20207 (N_20207,N_18438,N_16854);
nor U20208 (N_20208,N_15836,N_18648);
nand U20209 (N_20209,N_18290,N_15797);
nor U20210 (N_20210,N_15945,N_16548);
and U20211 (N_20211,N_16434,N_18405);
nand U20212 (N_20212,N_17935,N_17153);
nand U20213 (N_20213,N_17646,N_17196);
nand U20214 (N_20214,N_17491,N_17398);
nand U20215 (N_20215,N_18167,N_16477);
and U20216 (N_20216,N_18532,N_17102);
nand U20217 (N_20217,N_16331,N_15707);
xnor U20218 (N_20218,N_17625,N_17374);
and U20219 (N_20219,N_18414,N_15682);
xor U20220 (N_20220,N_16849,N_17589);
nor U20221 (N_20221,N_15782,N_18096);
nor U20222 (N_20222,N_18402,N_15789);
nor U20223 (N_20223,N_16513,N_16049);
nand U20224 (N_20224,N_16903,N_18195);
nand U20225 (N_20225,N_16660,N_15913);
nand U20226 (N_20226,N_16486,N_17182);
nand U20227 (N_20227,N_18403,N_17171);
nand U20228 (N_20228,N_17965,N_16191);
xnor U20229 (N_20229,N_16156,N_16058);
or U20230 (N_20230,N_16622,N_18705);
nor U20231 (N_20231,N_18590,N_18400);
nor U20232 (N_20232,N_17269,N_17793);
and U20233 (N_20233,N_18675,N_18550);
or U20234 (N_20234,N_17285,N_17107);
nand U20235 (N_20235,N_18684,N_17936);
and U20236 (N_20236,N_17186,N_16318);
nand U20237 (N_20237,N_16765,N_16820);
nand U20238 (N_20238,N_17399,N_17764);
nor U20239 (N_20239,N_17447,N_16103);
or U20240 (N_20240,N_18739,N_15765);
or U20241 (N_20241,N_17754,N_17512);
nand U20242 (N_20242,N_17118,N_17807);
or U20243 (N_20243,N_16287,N_17795);
nor U20244 (N_20244,N_18307,N_17645);
nand U20245 (N_20245,N_17232,N_16149);
xnor U20246 (N_20246,N_16636,N_17236);
and U20247 (N_20247,N_16845,N_15900);
nand U20248 (N_20248,N_18582,N_17592);
and U20249 (N_20249,N_16994,N_18284);
and U20250 (N_20250,N_17954,N_17298);
nand U20251 (N_20251,N_17494,N_17037);
nor U20252 (N_20252,N_18105,N_17966);
nor U20253 (N_20253,N_16576,N_18015);
or U20254 (N_20254,N_17162,N_16882);
and U20255 (N_20255,N_18435,N_18207);
or U20256 (N_20256,N_16857,N_17734);
and U20257 (N_20257,N_16254,N_15819);
or U20258 (N_20258,N_15626,N_17090);
nand U20259 (N_20259,N_16789,N_16314);
nor U20260 (N_20260,N_16613,N_16955);
nand U20261 (N_20261,N_18097,N_16642);
or U20262 (N_20262,N_18331,N_16672);
nand U20263 (N_20263,N_16139,N_16061);
or U20264 (N_20264,N_18743,N_16872);
or U20265 (N_20265,N_18169,N_16979);
xor U20266 (N_20266,N_15774,N_18035);
and U20267 (N_20267,N_17614,N_16190);
nand U20268 (N_20268,N_18407,N_18098);
nand U20269 (N_20269,N_17109,N_16078);
or U20270 (N_20270,N_16526,N_16631);
nor U20271 (N_20271,N_18544,N_16375);
or U20272 (N_20272,N_17292,N_17364);
xnor U20273 (N_20273,N_18027,N_15894);
nor U20274 (N_20274,N_18223,N_16235);
and U20275 (N_20275,N_18079,N_15750);
nand U20276 (N_20276,N_18542,N_17692);
nand U20277 (N_20277,N_17619,N_15730);
nand U20278 (N_20278,N_15839,N_17948);
nor U20279 (N_20279,N_16730,N_16192);
nor U20280 (N_20280,N_18406,N_17311);
nor U20281 (N_20281,N_16784,N_16726);
nor U20282 (N_20282,N_16783,N_17071);
nand U20283 (N_20283,N_16745,N_16289);
nand U20284 (N_20284,N_15893,N_16770);
and U20285 (N_20285,N_15646,N_17772);
nor U20286 (N_20286,N_17432,N_15899);
or U20287 (N_20287,N_17357,N_18603);
and U20288 (N_20288,N_16973,N_17887);
nand U20289 (N_20289,N_18442,N_15872);
nor U20290 (N_20290,N_17514,N_15733);
and U20291 (N_20291,N_15736,N_16332);
xnor U20292 (N_20292,N_16497,N_15710);
xnor U20293 (N_20293,N_17913,N_16887);
nand U20294 (N_20294,N_18233,N_16913);
nand U20295 (N_20295,N_18485,N_18061);
and U20296 (N_20296,N_18748,N_17025);
or U20297 (N_20297,N_17907,N_18710);
nor U20298 (N_20298,N_16261,N_17078);
or U20299 (N_20299,N_17654,N_17437);
and U20300 (N_20300,N_16485,N_18095);
nor U20301 (N_20301,N_16842,N_17467);
and U20302 (N_20302,N_18206,N_17128);
nor U20303 (N_20303,N_17016,N_18617);
or U20304 (N_20304,N_16271,N_17354);
and U20305 (N_20305,N_16643,N_15842);
and U20306 (N_20306,N_16701,N_18516);
or U20307 (N_20307,N_17870,N_18697);
nor U20308 (N_20308,N_16686,N_17616);
and U20309 (N_20309,N_18700,N_15864);
or U20310 (N_20310,N_15806,N_17076);
or U20311 (N_20311,N_18746,N_18737);
or U20312 (N_20312,N_18152,N_17390);
or U20313 (N_20313,N_17173,N_17044);
nand U20314 (N_20314,N_16752,N_18241);
xor U20315 (N_20315,N_16957,N_16870);
nor U20316 (N_20316,N_16379,N_17828);
nor U20317 (N_20317,N_17139,N_16446);
and U20318 (N_20318,N_16964,N_17844);
nor U20319 (N_20319,N_17266,N_18341);
nand U20320 (N_20320,N_15710,N_17993);
nand U20321 (N_20321,N_18023,N_17724);
nand U20322 (N_20322,N_18031,N_18396);
nand U20323 (N_20323,N_18388,N_17505);
or U20324 (N_20324,N_15921,N_18260);
and U20325 (N_20325,N_16536,N_16197);
nor U20326 (N_20326,N_17526,N_18579);
and U20327 (N_20327,N_17017,N_16802);
and U20328 (N_20328,N_15909,N_18368);
nand U20329 (N_20329,N_17114,N_18325);
or U20330 (N_20330,N_16850,N_17349);
nand U20331 (N_20331,N_18403,N_17301);
xnor U20332 (N_20332,N_17334,N_15644);
or U20333 (N_20333,N_15692,N_18473);
nand U20334 (N_20334,N_15625,N_17619);
or U20335 (N_20335,N_15737,N_16265);
and U20336 (N_20336,N_17321,N_16095);
and U20337 (N_20337,N_18295,N_18139);
nand U20338 (N_20338,N_18598,N_18015);
nand U20339 (N_20339,N_17255,N_16723);
nand U20340 (N_20340,N_18082,N_16521);
or U20341 (N_20341,N_15797,N_18161);
and U20342 (N_20342,N_17717,N_15857);
or U20343 (N_20343,N_17581,N_16933);
or U20344 (N_20344,N_16214,N_17726);
nor U20345 (N_20345,N_16176,N_17147);
nand U20346 (N_20346,N_18156,N_18171);
and U20347 (N_20347,N_16100,N_18017);
or U20348 (N_20348,N_17671,N_15814);
or U20349 (N_20349,N_16847,N_15840);
xor U20350 (N_20350,N_18558,N_16836);
and U20351 (N_20351,N_16139,N_18582);
and U20352 (N_20352,N_16831,N_16184);
nor U20353 (N_20353,N_16740,N_17783);
nor U20354 (N_20354,N_16803,N_16472);
and U20355 (N_20355,N_16529,N_17525);
nor U20356 (N_20356,N_16388,N_17989);
and U20357 (N_20357,N_16644,N_16848);
nand U20358 (N_20358,N_17793,N_16680);
and U20359 (N_20359,N_16759,N_15786);
or U20360 (N_20360,N_16161,N_17494);
and U20361 (N_20361,N_17729,N_16265);
or U20362 (N_20362,N_17835,N_18465);
and U20363 (N_20363,N_17497,N_16586);
and U20364 (N_20364,N_16273,N_16124);
nand U20365 (N_20365,N_16035,N_17080);
or U20366 (N_20366,N_17690,N_17723);
and U20367 (N_20367,N_15885,N_16149);
and U20368 (N_20368,N_17410,N_18436);
xor U20369 (N_20369,N_17441,N_18344);
or U20370 (N_20370,N_17665,N_15774);
xnor U20371 (N_20371,N_16087,N_16933);
or U20372 (N_20372,N_16642,N_17683);
or U20373 (N_20373,N_17088,N_15745);
nor U20374 (N_20374,N_16995,N_18270);
nor U20375 (N_20375,N_16113,N_16082);
and U20376 (N_20376,N_18498,N_15860);
nor U20377 (N_20377,N_18294,N_16582);
nor U20378 (N_20378,N_16648,N_15709);
or U20379 (N_20379,N_17638,N_16411);
or U20380 (N_20380,N_16393,N_18644);
nor U20381 (N_20381,N_15919,N_15686);
xnor U20382 (N_20382,N_17580,N_16679);
and U20383 (N_20383,N_17936,N_17161);
nor U20384 (N_20384,N_16336,N_16941);
and U20385 (N_20385,N_18672,N_16883);
xor U20386 (N_20386,N_18430,N_17822);
nor U20387 (N_20387,N_18269,N_15989);
nand U20388 (N_20388,N_15833,N_17406);
nor U20389 (N_20389,N_15991,N_16687);
nor U20390 (N_20390,N_17564,N_18153);
nor U20391 (N_20391,N_17193,N_17545);
nand U20392 (N_20392,N_15884,N_17672);
nor U20393 (N_20393,N_16457,N_16055);
nand U20394 (N_20394,N_17557,N_16272);
nand U20395 (N_20395,N_17395,N_15694);
nand U20396 (N_20396,N_18469,N_15859);
nand U20397 (N_20397,N_17214,N_17797);
nor U20398 (N_20398,N_17014,N_18164);
nand U20399 (N_20399,N_18718,N_17607);
and U20400 (N_20400,N_16776,N_18159);
nand U20401 (N_20401,N_18152,N_17553);
nor U20402 (N_20402,N_17710,N_17052);
nand U20403 (N_20403,N_15979,N_15939);
xnor U20404 (N_20404,N_17997,N_18050);
xor U20405 (N_20405,N_18309,N_16079);
or U20406 (N_20406,N_16437,N_18462);
and U20407 (N_20407,N_18515,N_15870);
or U20408 (N_20408,N_16583,N_17951);
nand U20409 (N_20409,N_18452,N_17104);
and U20410 (N_20410,N_18370,N_16347);
nor U20411 (N_20411,N_16582,N_18524);
nor U20412 (N_20412,N_18477,N_17625);
nor U20413 (N_20413,N_18041,N_18197);
or U20414 (N_20414,N_17098,N_18263);
and U20415 (N_20415,N_15980,N_18409);
nor U20416 (N_20416,N_16989,N_16547);
nand U20417 (N_20417,N_16376,N_15906);
and U20418 (N_20418,N_16105,N_18556);
or U20419 (N_20419,N_17255,N_17520);
or U20420 (N_20420,N_17077,N_17770);
or U20421 (N_20421,N_16395,N_18654);
nor U20422 (N_20422,N_17696,N_17979);
or U20423 (N_20423,N_16458,N_18667);
nor U20424 (N_20424,N_16951,N_17787);
or U20425 (N_20425,N_18481,N_17364);
and U20426 (N_20426,N_17285,N_18267);
and U20427 (N_20427,N_18186,N_18073);
nor U20428 (N_20428,N_17187,N_15959);
nor U20429 (N_20429,N_16131,N_17240);
and U20430 (N_20430,N_16089,N_15627);
nor U20431 (N_20431,N_17365,N_16634);
and U20432 (N_20432,N_16292,N_18068);
nand U20433 (N_20433,N_16016,N_17703);
or U20434 (N_20434,N_17874,N_16085);
or U20435 (N_20435,N_15768,N_15935);
nor U20436 (N_20436,N_18351,N_16849);
or U20437 (N_20437,N_17722,N_18389);
nand U20438 (N_20438,N_17164,N_16675);
and U20439 (N_20439,N_18306,N_17748);
and U20440 (N_20440,N_16472,N_16478);
and U20441 (N_20441,N_15750,N_17962);
nor U20442 (N_20442,N_15928,N_16470);
and U20443 (N_20443,N_15808,N_15873);
or U20444 (N_20444,N_17905,N_15844);
nand U20445 (N_20445,N_16317,N_18656);
or U20446 (N_20446,N_17331,N_16996);
nor U20447 (N_20447,N_17933,N_16398);
nand U20448 (N_20448,N_15889,N_16970);
nand U20449 (N_20449,N_18655,N_16627);
and U20450 (N_20450,N_18134,N_18614);
nand U20451 (N_20451,N_17450,N_18154);
and U20452 (N_20452,N_17476,N_16362);
and U20453 (N_20453,N_17575,N_17726);
nor U20454 (N_20454,N_16261,N_16495);
and U20455 (N_20455,N_16581,N_16154);
nand U20456 (N_20456,N_15949,N_17987);
nand U20457 (N_20457,N_17670,N_16634);
or U20458 (N_20458,N_15666,N_18262);
or U20459 (N_20459,N_16255,N_16195);
nor U20460 (N_20460,N_17094,N_16233);
nor U20461 (N_20461,N_18053,N_17455);
and U20462 (N_20462,N_17192,N_15949);
nor U20463 (N_20463,N_18566,N_16116);
and U20464 (N_20464,N_16866,N_16482);
nor U20465 (N_20465,N_16013,N_15867);
or U20466 (N_20466,N_17289,N_15808);
or U20467 (N_20467,N_18486,N_18257);
nand U20468 (N_20468,N_15954,N_15873);
xnor U20469 (N_20469,N_16340,N_17160);
and U20470 (N_20470,N_17234,N_18014);
nor U20471 (N_20471,N_16836,N_17396);
xor U20472 (N_20472,N_18512,N_17294);
nor U20473 (N_20473,N_17577,N_16415);
xnor U20474 (N_20474,N_15904,N_15932);
nor U20475 (N_20475,N_17111,N_17973);
nor U20476 (N_20476,N_18251,N_16865);
nor U20477 (N_20477,N_17066,N_16491);
and U20478 (N_20478,N_18175,N_16713);
and U20479 (N_20479,N_17920,N_17520);
xor U20480 (N_20480,N_18177,N_16162);
and U20481 (N_20481,N_18358,N_16549);
and U20482 (N_20482,N_18343,N_15684);
nor U20483 (N_20483,N_18070,N_16480);
nand U20484 (N_20484,N_16468,N_17819);
and U20485 (N_20485,N_17135,N_18181);
xor U20486 (N_20486,N_17894,N_17651);
nand U20487 (N_20487,N_17149,N_17043);
nand U20488 (N_20488,N_18491,N_16500);
or U20489 (N_20489,N_16344,N_17201);
or U20490 (N_20490,N_16404,N_16965);
and U20491 (N_20491,N_18574,N_16711);
nor U20492 (N_20492,N_16052,N_16897);
nand U20493 (N_20493,N_15706,N_18352);
and U20494 (N_20494,N_17725,N_17383);
and U20495 (N_20495,N_18057,N_16697);
nor U20496 (N_20496,N_18725,N_17846);
xor U20497 (N_20497,N_17037,N_18395);
nand U20498 (N_20498,N_18469,N_17005);
and U20499 (N_20499,N_16933,N_16007);
and U20500 (N_20500,N_17458,N_16552);
and U20501 (N_20501,N_18644,N_15743);
nor U20502 (N_20502,N_16454,N_15850);
or U20503 (N_20503,N_15895,N_18055);
and U20504 (N_20504,N_17236,N_16060);
and U20505 (N_20505,N_18056,N_16090);
nor U20506 (N_20506,N_18411,N_17140);
nand U20507 (N_20507,N_15854,N_17365);
or U20508 (N_20508,N_17158,N_17284);
nor U20509 (N_20509,N_16702,N_18461);
nand U20510 (N_20510,N_17881,N_15872);
or U20511 (N_20511,N_16457,N_18347);
nor U20512 (N_20512,N_17287,N_16084);
and U20513 (N_20513,N_17169,N_16558);
nor U20514 (N_20514,N_17475,N_17606);
nor U20515 (N_20515,N_15635,N_16296);
or U20516 (N_20516,N_17394,N_15731);
nor U20517 (N_20517,N_16247,N_17408);
and U20518 (N_20518,N_17984,N_16489);
nand U20519 (N_20519,N_17157,N_18359);
xnor U20520 (N_20520,N_17567,N_17349);
and U20521 (N_20521,N_15716,N_16672);
and U20522 (N_20522,N_16853,N_16453);
xnor U20523 (N_20523,N_18151,N_16797);
nor U20524 (N_20524,N_16838,N_15687);
or U20525 (N_20525,N_18439,N_18594);
nand U20526 (N_20526,N_17068,N_18672);
or U20527 (N_20527,N_17497,N_17286);
nand U20528 (N_20528,N_18461,N_16527);
and U20529 (N_20529,N_16614,N_15963);
nor U20530 (N_20530,N_17248,N_17029);
nand U20531 (N_20531,N_18368,N_17008);
xnor U20532 (N_20532,N_17081,N_15987);
and U20533 (N_20533,N_17886,N_16211);
xnor U20534 (N_20534,N_16593,N_16096);
or U20535 (N_20535,N_17934,N_18504);
and U20536 (N_20536,N_16891,N_16972);
nor U20537 (N_20537,N_16488,N_15876);
or U20538 (N_20538,N_16529,N_16931);
nand U20539 (N_20539,N_16741,N_16098);
nor U20540 (N_20540,N_18737,N_16826);
or U20541 (N_20541,N_17803,N_15854);
or U20542 (N_20542,N_16023,N_17082);
and U20543 (N_20543,N_18406,N_18575);
nor U20544 (N_20544,N_15867,N_15837);
and U20545 (N_20545,N_16625,N_17342);
or U20546 (N_20546,N_17222,N_15652);
nor U20547 (N_20547,N_18724,N_17085);
nand U20548 (N_20548,N_17241,N_18516);
and U20549 (N_20549,N_16037,N_16882);
or U20550 (N_20550,N_18642,N_15846);
or U20551 (N_20551,N_18479,N_18062);
and U20552 (N_20552,N_15660,N_18169);
and U20553 (N_20553,N_16307,N_17350);
xnor U20554 (N_20554,N_17275,N_16874);
and U20555 (N_20555,N_18197,N_17505);
or U20556 (N_20556,N_17977,N_18150);
nor U20557 (N_20557,N_16661,N_16207);
or U20558 (N_20558,N_17290,N_18610);
nand U20559 (N_20559,N_18555,N_16811);
or U20560 (N_20560,N_18186,N_16553);
and U20561 (N_20561,N_18091,N_17592);
and U20562 (N_20562,N_16564,N_16120);
and U20563 (N_20563,N_17285,N_15848);
and U20564 (N_20564,N_17453,N_17026);
nand U20565 (N_20565,N_17102,N_18174);
nand U20566 (N_20566,N_18406,N_18445);
nor U20567 (N_20567,N_15963,N_16904);
nand U20568 (N_20568,N_17157,N_16091);
or U20569 (N_20569,N_18178,N_16638);
xnor U20570 (N_20570,N_16726,N_18186);
or U20571 (N_20571,N_17237,N_18194);
nor U20572 (N_20572,N_16643,N_18394);
nor U20573 (N_20573,N_15961,N_16004);
nand U20574 (N_20574,N_16733,N_16433);
and U20575 (N_20575,N_16602,N_16458);
nor U20576 (N_20576,N_17845,N_18590);
nor U20577 (N_20577,N_17626,N_17382);
nor U20578 (N_20578,N_15803,N_16220);
or U20579 (N_20579,N_17959,N_17663);
and U20580 (N_20580,N_16415,N_16164);
nor U20581 (N_20581,N_17406,N_16802);
nor U20582 (N_20582,N_15992,N_16488);
nor U20583 (N_20583,N_18008,N_17944);
and U20584 (N_20584,N_16663,N_16323);
nand U20585 (N_20585,N_18319,N_16929);
nand U20586 (N_20586,N_18339,N_18178);
or U20587 (N_20587,N_16048,N_16842);
and U20588 (N_20588,N_17865,N_16660);
nor U20589 (N_20589,N_17757,N_18143);
nand U20590 (N_20590,N_17393,N_17758);
nor U20591 (N_20591,N_17234,N_18019);
and U20592 (N_20592,N_18383,N_16845);
and U20593 (N_20593,N_18238,N_17220);
xor U20594 (N_20594,N_18310,N_18046);
nand U20595 (N_20595,N_17005,N_16084);
and U20596 (N_20596,N_16483,N_18362);
nand U20597 (N_20597,N_17200,N_16278);
nor U20598 (N_20598,N_15972,N_18417);
or U20599 (N_20599,N_16091,N_16914);
and U20600 (N_20600,N_15655,N_17674);
nand U20601 (N_20601,N_16273,N_18563);
and U20602 (N_20602,N_15643,N_17632);
and U20603 (N_20603,N_15653,N_15985);
nand U20604 (N_20604,N_18448,N_16280);
nor U20605 (N_20605,N_16588,N_17241);
nand U20606 (N_20606,N_18381,N_16973);
nor U20607 (N_20607,N_16832,N_17693);
and U20608 (N_20608,N_18335,N_16578);
and U20609 (N_20609,N_18423,N_16368);
xnor U20610 (N_20610,N_17284,N_17774);
xor U20611 (N_20611,N_18381,N_17882);
or U20612 (N_20612,N_17889,N_16983);
and U20613 (N_20613,N_16240,N_18156);
nand U20614 (N_20614,N_16560,N_15673);
and U20615 (N_20615,N_18469,N_16311);
and U20616 (N_20616,N_17364,N_17913);
or U20617 (N_20617,N_17916,N_18121);
or U20618 (N_20618,N_16405,N_15953);
and U20619 (N_20619,N_16916,N_16016);
nand U20620 (N_20620,N_17666,N_18084);
or U20621 (N_20621,N_17069,N_16783);
nand U20622 (N_20622,N_16188,N_18671);
and U20623 (N_20623,N_16409,N_17554);
nor U20624 (N_20624,N_18156,N_17647);
nand U20625 (N_20625,N_18287,N_15891);
and U20626 (N_20626,N_16178,N_16702);
nor U20627 (N_20627,N_18419,N_16418);
or U20628 (N_20628,N_17993,N_16041);
or U20629 (N_20629,N_17120,N_18321);
and U20630 (N_20630,N_17908,N_18240);
nand U20631 (N_20631,N_16805,N_16367);
and U20632 (N_20632,N_17274,N_17911);
nand U20633 (N_20633,N_17315,N_17878);
nor U20634 (N_20634,N_18162,N_18379);
and U20635 (N_20635,N_16397,N_18151);
xor U20636 (N_20636,N_16764,N_15869);
or U20637 (N_20637,N_16730,N_17024);
or U20638 (N_20638,N_18669,N_16644);
or U20639 (N_20639,N_16494,N_18012);
or U20640 (N_20640,N_18136,N_16212);
nor U20641 (N_20641,N_16826,N_17858);
nor U20642 (N_20642,N_18212,N_15799);
and U20643 (N_20643,N_17126,N_18016);
or U20644 (N_20644,N_18282,N_16257);
or U20645 (N_20645,N_17161,N_17371);
and U20646 (N_20646,N_16488,N_16811);
and U20647 (N_20647,N_18490,N_17360);
xnor U20648 (N_20648,N_16876,N_15741);
nor U20649 (N_20649,N_18113,N_16760);
nor U20650 (N_20650,N_18179,N_16304);
and U20651 (N_20651,N_17652,N_15902);
nand U20652 (N_20652,N_15951,N_16030);
nand U20653 (N_20653,N_16808,N_15890);
nor U20654 (N_20654,N_18412,N_18668);
and U20655 (N_20655,N_15952,N_17739);
nor U20656 (N_20656,N_18407,N_18028);
nand U20657 (N_20657,N_17952,N_17556);
nor U20658 (N_20658,N_17694,N_15648);
nor U20659 (N_20659,N_17912,N_15872);
and U20660 (N_20660,N_18596,N_18248);
nor U20661 (N_20661,N_17459,N_17849);
nor U20662 (N_20662,N_16321,N_16714);
and U20663 (N_20663,N_16010,N_16093);
or U20664 (N_20664,N_17691,N_15755);
nand U20665 (N_20665,N_18643,N_17116);
nand U20666 (N_20666,N_16060,N_17605);
nor U20667 (N_20667,N_16104,N_17384);
nand U20668 (N_20668,N_17691,N_18173);
xnor U20669 (N_20669,N_17504,N_17759);
and U20670 (N_20670,N_18447,N_16682);
or U20671 (N_20671,N_18287,N_18575);
nand U20672 (N_20672,N_17560,N_18101);
nand U20673 (N_20673,N_16111,N_15919);
and U20674 (N_20674,N_18200,N_15894);
and U20675 (N_20675,N_17412,N_18321);
nor U20676 (N_20676,N_18282,N_16102);
or U20677 (N_20677,N_16396,N_16898);
nor U20678 (N_20678,N_16265,N_16443);
nand U20679 (N_20679,N_17262,N_18221);
nand U20680 (N_20680,N_17605,N_17895);
nor U20681 (N_20681,N_17815,N_16003);
nor U20682 (N_20682,N_18252,N_18596);
nand U20683 (N_20683,N_17925,N_18141);
and U20684 (N_20684,N_18061,N_18699);
nand U20685 (N_20685,N_18002,N_17908);
and U20686 (N_20686,N_17127,N_15814);
xnor U20687 (N_20687,N_16539,N_17823);
and U20688 (N_20688,N_17184,N_17593);
nor U20689 (N_20689,N_16993,N_18596);
or U20690 (N_20690,N_16880,N_16527);
and U20691 (N_20691,N_18130,N_18277);
nand U20692 (N_20692,N_16617,N_17623);
nand U20693 (N_20693,N_18312,N_18014);
and U20694 (N_20694,N_16471,N_16923);
nand U20695 (N_20695,N_16072,N_18443);
or U20696 (N_20696,N_17387,N_17471);
or U20697 (N_20697,N_16319,N_16151);
xnor U20698 (N_20698,N_15747,N_17609);
or U20699 (N_20699,N_16104,N_16997);
nor U20700 (N_20700,N_16000,N_17259);
nor U20701 (N_20701,N_17188,N_18682);
nor U20702 (N_20702,N_16588,N_16872);
nor U20703 (N_20703,N_16676,N_16595);
and U20704 (N_20704,N_15880,N_16776);
xnor U20705 (N_20705,N_16452,N_15899);
or U20706 (N_20706,N_17078,N_17985);
or U20707 (N_20707,N_18038,N_16119);
nand U20708 (N_20708,N_17695,N_17668);
xnor U20709 (N_20709,N_18117,N_16099);
or U20710 (N_20710,N_17728,N_16349);
or U20711 (N_20711,N_17947,N_17642);
nor U20712 (N_20712,N_18422,N_15764);
nor U20713 (N_20713,N_15754,N_16178);
or U20714 (N_20714,N_16900,N_16459);
nand U20715 (N_20715,N_18553,N_16156);
nor U20716 (N_20716,N_16558,N_17867);
xnor U20717 (N_20717,N_15929,N_16417);
and U20718 (N_20718,N_17898,N_15955);
and U20719 (N_20719,N_16436,N_18158);
nor U20720 (N_20720,N_16587,N_18069);
nand U20721 (N_20721,N_16765,N_16898);
and U20722 (N_20722,N_17047,N_16754);
xnor U20723 (N_20723,N_17368,N_17411);
and U20724 (N_20724,N_15732,N_16681);
or U20725 (N_20725,N_17756,N_17562);
nor U20726 (N_20726,N_16962,N_16842);
or U20727 (N_20727,N_16462,N_16893);
and U20728 (N_20728,N_17709,N_17577);
nand U20729 (N_20729,N_15727,N_18225);
nand U20730 (N_20730,N_16004,N_18626);
nand U20731 (N_20731,N_17260,N_18198);
nand U20732 (N_20732,N_18519,N_18069);
or U20733 (N_20733,N_17353,N_18156);
and U20734 (N_20734,N_18375,N_15719);
and U20735 (N_20735,N_16481,N_15933);
nand U20736 (N_20736,N_16288,N_18651);
or U20737 (N_20737,N_17958,N_18032);
or U20738 (N_20738,N_17745,N_17929);
and U20739 (N_20739,N_17108,N_16177);
nand U20740 (N_20740,N_15860,N_16590);
nor U20741 (N_20741,N_17121,N_17657);
nand U20742 (N_20742,N_18722,N_17532);
or U20743 (N_20743,N_16584,N_17827);
nand U20744 (N_20744,N_16683,N_16478);
and U20745 (N_20745,N_17932,N_16424);
or U20746 (N_20746,N_15767,N_15797);
nor U20747 (N_20747,N_16942,N_17207);
and U20748 (N_20748,N_17434,N_16968);
and U20749 (N_20749,N_16557,N_16195);
nor U20750 (N_20750,N_17452,N_18024);
and U20751 (N_20751,N_16574,N_18349);
and U20752 (N_20752,N_17774,N_15679);
and U20753 (N_20753,N_16549,N_17829);
or U20754 (N_20754,N_18001,N_16860);
nand U20755 (N_20755,N_18745,N_18680);
or U20756 (N_20756,N_17888,N_16457);
nor U20757 (N_20757,N_15735,N_18494);
nand U20758 (N_20758,N_18235,N_18083);
nor U20759 (N_20759,N_17343,N_15944);
or U20760 (N_20760,N_17917,N_17216);
xnor U20761 (N_20761,N_16867,N_18303);
nor U20762 (N_20762,N_16959,N_16788);
xor U20763 (N_20763,N_15784,N_17060);
and U20764 (N_20764,N_18339,N_18535);
or U20765 (N_20765,N_18465,N_17609);
and U20766 (N_20766,N_15905,N_18485);
or U20767 (N_20767,N_17626,N_16197);
nand U20768 (N_20768,N_17883,N_17783);
or U20769 (N_20769,N_16689,N_17736);
or U20770 (N_20770,N_16892,N_16789);
and U20771 (N_20771,N_18473,N_16391);
nand U20772 (N_20772,N_17047,N_18428);
nor U20773 (N_20773,N_18515,N_18324);
or U20774 (N_20774,N_17087,N_18150);
nand U20775 (N_20775,N_16174,N_17673);
xor U20776 (N_20776,N_16244,N_16161);
nor U20777 (N_20777,N_18254,N_18377);
and U20778 (N_20778,N_17874,N_16237);
or U20779 (N_20779,N_17958,N_16678);
or U20780 (N_20780,N_16293,N_17146);
xor U20781 (N_20781,N_17148,N_17943);
xor U20782 (N_20782,N_17221,N_18483);
nor U20783 (N_20783,N_18542,N_17430);
or U20784 (N_20784,N_18425,N_15844);
or U20785 (N_20785,N_16849,N_18663);
nor U20786 (N_20786,N_18157,N_16956);
nor U20787 (N_20787,N_17991,N_15974);
xnor U20788 (N_20788,N_16512,N_18652);
nor U20789 (N_20789,N_16874,N_18442);
and U20790 (N_20790,N_18640,N_15849);
and U20791 (N_20791,N_16001,N_18041);
nor U20792 (N_20792,N_18336,N_16516);
xnor U20793 (N_20793,N_16118,N_17670);
nand U20794 (N_20794,N_17337,N_16903);
nand U20795 (N_20795,N_16448,N_18039);
nor U20796 (N_20796,N_16930,N_16029);
nor U20797 (N_20797,N_17576,N_18464);
or U20798 (N_20798,N_17895,N_17102);
xnor U20799 (N_20799,N_17448,N_17373);
and U20800 (N_20800,N_17169,N_17009);
and U20801 (N_20801,N_16548,N_16046);
nand U20802 (N_20802,N_17015,N_17948);
nand U20803 (N_20803,N_16382,N_16754);
xor U20804 (N_20804,N_16013,N_16234);
or U20805 (N_20805,N_17080,N_17795);
and U20806 (N_20806,N_17388,N_16123);
nor U20807 (N_20807,N_17537,N_16192);
and U20808 (N_20808,N_16456,N_16200);
nand U20809 (N_20809,N_16218,N_17215);
nand U20810 (N_20810,N_15650,N_18075);
or U20811 (N_20811,N_16298,N_15850);
nor U20812 (N_20812,N_16963,N_17703);
and U20813 (N_20813,N_16755,N_18219);
nand U20814 (N_20814,N_18491,N_17357);
nand U20815 (N_20815,N_16460,N_17680);
nand U20816 (N_20816,N_18427,N_16609);
and U20817 (N_20817,N_16763,N_18402);
or U20818 (N_20818,N_15879,N_17630);
or U20819 (N_20819,N_17452,N_17551);
nand U20820 (N_20820,N_16986,N_17566);
and U20821 (N_20821,N_18436,N_15742);
nor U20822 (N_20822,N_17940,N_18504);
nor U20823 (N_20823,N_18527,N_16932);
and U20824 (N_20824,N_18572,N_18665);
nor U20825 (N_20825,N_18697,N_17816);
nand U20826 (N_20826,N_17908,N_18443);
or U20827 (N_20827,N_17998,N_15898);
nor U20828 (N_20828,N_18435,N_18388);
nor U20829 (N_20829,N_16567,N_17550);
xor U20830 (N_20830,N_17576,N_16805);
nor U20831 (N_20831,N_17341,N_15881);
or U20832 (N_20832,N_16537,N_18347);
nand U20833 (N_20833,N_18428,N_16094);
nor U20834 (N_20834,N_16251,N_18548);
or U20835 (N_20835,N_16335,N_17022);
or U20836 (N_20836,N_15810,N_16498);
nand U20837 (N_20837,N_18699,N_16949);
nand U20838 (N_20838,N_17980,N_16019);
and U20839 (N_20839,N_17101,N_18078);
and U20840 (N_20840,N_18002,N_17486);
nand U20841 (N_20841,N_16028,N_17974);
nand U20842 (N_20842,N_17090,N_17623);
xnor U20843 (N_20843,N_17094,N_15991);
nor U20844 (N_20844,N_16207,N_17724);
nor U20845 (N_20845,N_15757,N_17379);
and U20846 (N_20846,N_17873,N_16226);
nor U20847 (N_20847,N_16397,N_18032);
or U20848 (N_20848,N_15999,N_16166);
or U20849 (N_20849,N_18134,N_16966);
nor U20850 (N_20850,N_16899,N_16256);
xnor U20851 (N_20851,N_15657,N_16718);
and U20852 (N_20852,N_17074,N_16257);
nand U20853 (N_20853,N_17541,N_18541);
and U20854 (N_20854,N_17527,N_16225);
nand U20855 (N_20855,N_18638,N_15728);
nor U20856 (N_20856,N_16850,N_16164);
or U20857 (N_20857,N_15806,N_18689);
nor U20858 (N_20858,N_18238,N_16830);
or U20859 (N_20859,N_18259,N_16021);
nor U20860 (N_20860,N_16838,N_16846);
and U20861 (N_20861,N_18481,N_17840);
and U20862 (N_20862,N_18339,N_17270);
nand U20863 (N_20863,N_15930,N_16979);
or U20864 (N_20864,N_17106,N_17430);
or U20865 (N_20865,N_17699,N_15942);
or U20866 (N_20866,N_16725,N_17731);
and U20867 (N_20867,N_16036,N_16779);
and U20868 (N_20868,N_16199,N_18533);
xnor U20869 (N_20869,N_18404,N_17766);
and U20870 (N_20870,N_17241,N_16290);
or U20871 (N_20871,N_17101,N_17016);
nor U20872 (N_20872,N_17858,N_16400);
nor U20873 (N_20873,N_16947,N_16398);
nand U20874 (N_20874,N_17749,N_18497);
and U20875 (N_20875,N_17042,N_17739);
xor U20876 (N_20876,N_17408,N_15908);
nor U20877 (N_20877,N_17245,N_16226);
xnor U20878 (N_20878,N_15823,N_17966);
xnor U20879 (N_20879,N_17487,N_17548);
and U20880 (N_20880,N_18735,N_15736);
xor U20881 (N_20881,N_17964,N_16988);
and U20882 (N_20882,N_15703,N_16083);
or U20883 (N_20883,N_17199,N_16680);
nor U20884 (N_20884,N_17944,N_15910);
nand U20885 (N_20885,N_15731,N_18661);
and U20886 (N_20886,N_18467,N_16758);
or U20887 (N_20887,N_16038,N_18663);
nand U20888 (N_20888,N_18322,N_18146);
nor U20889 (N_20889,N_16715,N_17437);
and U20890 (N_20890,N_15711,N_16789);
and U20891 (N_20891,N_17209,N_18677);
and U20892 (N_20892,N_18379,N_18467);
nor U20893 (N_20893,N_16950,N_18534);
and U20894 (N_20894,N_18467,N_16807);
or U20895 (N_20895,N_16178,N_16753);
and U20896 (N_20896,N_16823,N_18276);
and U20897 (N_20897,N_17580,N_16700);
nand U20898 (N_20898,N_16663,N_16620);
nand U20899 (N_20899,N_16309,N_18069);
nand U20900 (N_20900,N_17894,N_16478);
or U20901 (N_20901,N_18020,N_15860);
nor U20902 (N_20902,N_17064,N_17317);
or U20903 (N_20903,N_15710,N_16281);
nor U20904 (N_20904,N_18655,N_15827);
nor U20905 (N_20905,N_18724,N_17263);
and U20906 (N_20906,N_15818,N_16140);
nor U20907 (N_20907,N_18264,N_16222);
nand U20908 (N_20908,N_18037,N_18601);
or U20909 (N_20909,N_16303,N_17680);
or U20910 (N_20910,N_16147,N_16932);
nor U20911 (N_20911,N_17103,N_17890);
nand U20912 (N_20912,N_17092,N_17670);
or U20913 (N_20913,N_16545,N_15960);
and U20914 (N_20914,N_15942,N_17543);
or U20915 (N_20915,N_16612,N_17257);
or U20916 (N_20916,N_18397,N_18671);
nand U20917 (N_20917,N_18731,N_18233);
xor U20918 (N_20918,N_17629,N_17011);
nor U20919 (N_20919,N_18018,N_18558);
nor U20920 (N_20920,N_16973,N_17342);
nand U20921 (N_20921,N_17884,N_18683);
or U20922 (N_20922,N_16035,N_16984);
nand U20923 (N_20923,N_18652,N_18402);
nor U20924 (N_20924,N_16036,N_15768);
nor U20925 (N_20925,N_17793,N_18620);
or U20926 (N_20926,N_18463,N_18630);
nor U20927 (N_20927,N_16618,N_18661);
and U20928 (N_20928,N_17735,N_16127);
or U20929 (N_20929,N_16300,N_17501);
nor U20930 (N_20930,N_18690,N_18647);
nand U20931 (N_20931,N_16650,N_16160);
nand U20932 (N_20932,N_17408,N_16959);
and U20933 (N_20933,N_15921,N_16620);
or U20934 (N_20934,N_16272,N_17933);
xnor U20935 (N_20935,N_18723,N_15821);
nand U20936 (N_20936,N_17868,N_15992);
nor U20937 (N_20937,N_18685,N_18228);
and U20938 (N_20938,N_15741,N_16086);
and U20939 (N_20939,N_17565,N_15948);
nor U20940 (N_20940,N_18648,N_17421);
nor U20941 (N_20941,N_17767,N_15942);
and U20942 (N_20942,N_18551,N_17504);
nand U20943 (N_20943,N_17174,N_18684);
and U20944 (N_20944,N_15926,N_16746);
nand U20945 (N_20945,N_16006,N_16846);
xor U20946 (N_20946,N_16169,N_17662);
xor U20947 (N_20947,N_16157,N_17104);
nor U20948 (N_20948,N_17547,N_16113);
nand U20949 (N_20949,N_17062,N_16716);
and U20950 (N_20950,N_18631,N_17525);
and U20951 (N_20951,N_17143,N_18466);
or U20952 (N_20952,N_16049,N_15781);
xor U20953 (N_20953,N_17845,N_16171);
or U20954 (N_20954,N_18312,N_16116);
xor U20955 (N_20955,N_18107,N_16036);
and U20956 (N_20956,N_16333,N_16501);
nor U20957 (N_20957,N_18435,N_17611);
and U20958 (N_20958,N_17557,N_16435);
and U20959 (N_20959,N_18192,N_15904);
nand U20960 (N_20960,N_17480,N_16233);
or U20961 (N_20961,N_15965,N_15651);
nand U20962 (N_20962,N_16669,N_18161);
or U20963 (N_20963,N_18117,N_17718);
nand U20964 (N_20964,N_15634,N_18736);
nor U20965 (N_20965,N_17943,N_18048);
or U20966 (N_20966,N_16150,N_18579);
or U20967 (N_20967,N_17815,N_15817);
xnor U20968 (N_20968,N_16763,N_17648);
xnor U20969 (N_20969,N_18549,N_17466);
or U20970 (N_20970,N_17641,N_18062);
nor U20971 (N_20971,N_17485,N_15844);
and U20972 (N_20972,N_15637,N_16678);
or U20973 (N_20973,N_16392,N_15861);
xor U20974 (N_20974,N_17401,N_18265);
xnor U20975 (N_20975,N_17329,N_18669);
nor U20976 (N_20976,N_18133,N_15900);
and U20977 (N_20977,N_17543,N_15648);
nor U20978 (N_20978,N_15782,N_18109);
and U20979 (N_20979,N_18225,N_18627);
nand U20980 (N_20980,N_16070,N_16763);
nand U20981 (N_20981,N_18307,N_18654);
or U20982 (N_20982,N_15789,N_18736);
nand U20983 (N_20983,N_17344,N_16037);
or U20984 (N_20984,N_17510,N_16699);
nor U20985 (N_20985,N_17622,N_16896);
xor U20986 (N_20986,N_17838,N_18266);
or U20987 (N_20987,N_16022,N_17980);
nor U20988 (N_20988,N_15959,N_18223);
nor U20989 (N_20989,N_15941,N_16452);
or U20990 (N_20990,N_17856,N_16353);
xor U20991 (N_20991,N_17786,N_18161);
and U20992 (N_20992,N_18721,N_16640);
nand U20993 (N_20993,N_17553,N_17775);
nand U20994 (N_20994,N_15999,N_17198);
nor U20995 (N_20995,N_17968,N_18739);
and U20996 (N_20996,N_17805,N_16799);
and U20997 (N_20997,N_16740,N_18365);
or U20998 (N_20998,N_17477,N_18242);
or U20999 (N_20999,N_16655,N_17361);
nor U21000 (N_21000,N_17701,N_18566);
nand U21001 (N_21001,N_18058,N_18194);
or U21002 (N_21002,N_17867,N_17203);
and U21003 (N_21003,N_17028,N_16454);
or U21004 (N_21004,N_18075,N_16875);
nor U21005 (N_21005,N_16972,N_16695);
nand U21006 (N_21006,N_15746,N_15895);
nand U21007 (N_21007,N_17824,N_18253);
and U21008 (N_21008,N_18319,N_16654);
xor U21009 (N_21009,N_17270,N_18205);
and U21010 (N_21010,N_17265,N_17246);
xor U21011 (N_21011,N_16319,N_17521);
and U21012 (N_21012,N_17170,N_16023);
or U21013 (N_21013,N_18219,N_16517);
and U21014 (N_21014,N_18175,N_15928);
nand U21015 (N_21015,N_16131,N_15839);
nand U21016 (N_21016,N_16760,N_18216);
xor U21017 (N_21017,N_16113,N_18334);
and U21018 (N_21018,N_16654,N_15799);
or U21019 (N_21019,N_17507,N_17777);
nor U21020 (N_21020,N_16454,N_16203);
nand U21021 (N_21021,N_18279,N_15988);
nand U21022 (N_21022,N_18461,N_17948);
or U21023 (N_21023,N_17936,N_18720);
and U21024 (N_21024,N_17070,N_16188);
nor U21025 (N_21025,N_15704,N_16125);
and U21026 (N_21026,N_17463,N_18407);
xor U21027 (N_21027,N_16818,N_15729);
nor U21028 (N_21028,N_18319,N_16155);
and U21029 (N_21029,N_15763,N_17333);
nor U21030 (N_21030,N_17355,N_16290);
and U21031 (N_21031,N_15688,N_17961);
or U21032 (N_21032,N_16002,N_17853);
nand U21033 (N_21033,N_16220,N_16598);
nand U21034 (N_21034,N_18502,N_16303);
and U21035 (N_21035,N_17935,N_16990);
nor U21036 (N_21036,N_17460,N_18695);
and U21037 (N_21037,N_17434,N_17925);
nor U21038 (N_21038,N_16982,N_18337);
or U21039 (N_21039,N_17761,N_17341);
or U21040 (N_21040,N_17938,N_16944);
nor U21041 (N_21041,N_15631,N_15673);
and U21042 (N_21042,N_16776,N_18322);
nor U21043 (N_21043,N_17911,N_16756);
xnor U21044 (N_21044,N_17680,N_18664);
xnor U21045 (N_21045,N_18370,N_18247);
and U21046 (N_21046,N_18434,N_16589);
or U21047 (N_21047,N_16707,N_16871);
nor U21048 (N_21048,N_16078,N_18546);
and U21049 (N_21049,N_17372,N_17188);
or U21050 (N_21050,N_15928,N_18217);
or U21051 (N_21051,N_17431,N_16399);
nand U21052 (N_21052,N_18109,N_15765);
xor U21053 (N_21053,N_17724,N_15956);
xor U21054 (N_21054,N_18182,N_16884);
nand U21055 (N_21055,N_16889,N_18240);
or U21056 (N_21056,N_17513,N_16518);
nand U21057 (N_21057,N_15632,N_18591);
nand U21058 (N_21058,N_18655,N_18443);
nand U21059 (N_21059,N_17291,N_17509);
nor U21060 (N_21060,N_16790,N_16809);
nor U21061 (N_21061,N_16907,N_16230);
nand U21062 (N_21062,N_15882,N_17384);
xnor U21063 (N_21063,N_16332,N_18092);
or U21064 (N_21064,N_18002,N_18435);
nor U21065 (N_21065,N_16885,N_16305);
nand U21066 (N_21066,N_15762,N_16754);
or U21067 (N_21067,N_16471,N_15817);
nand U21068 (N_21068,N_15710,N_15723);
and U21069 (N_21069,N_16834,N_17320);
nand U21070 (N_21070,N_16575,N_18115);
or U21071 (N_21071,N_17916,N_16137);
and U21072 (N_21072,N_18279,N_16064);
xnor U21073 (N_21073,N_18615,N_16799);
or U21074 (N_21074,N_16276,N_15724);
nand U21075 (N_21075,N_17514,N_16145);
and U21076 (N_21076,N_15892,N_18496);
nand U21077 (N_21077,N_16323,N_16109);
and U21078 (N_21078,N_17630,N_16448);
or U21079 (N_21079,N_18487,N_16598);
xor U21080 (N_21080,N_17621,N_16032);
nor U21081 (N_21081,N_18074,N_18191);
nand U21082 (N_21082,N_18729,N_17179);
xor U21083 (N_21083,N_18275,N_17232);
and U21084 (N_21084,N_18331,N_18665);
xor U21085 (N_21085,N_15701,N_18672);
and U21086 (N_21086,N_17611,N_18350);
and U21087 (N_21087,N_17983,N_15722);
nand U21088 (N_21088,N_16868,N_15676);
nand U21089 (N_21089,N_16807,N_17626);
xnor U21090 (N_21090,N_16643,N_18116);
nand U21091 (N_21091,N_17991,N_18405);
or U21092 (N_21092,N_16352,N_18718);
or U21093 (N_21093,N_16214,N_15687);
and U21094 (N_21094,N_17517,N_16709);
or U21095 (N_21095,N_15819,N_17462);
nand U21096 (N_21096,N_18107,N_15865);
xor U21097 (N_21097,N_17643,N_15860);
nor U21098 (N_21098,N_17849,N_18686);
nor U21099 (N_21099,N_17005,N_16851);
or U21100 (N_21100,N_17520,N_17377);
or U21101 (N_21101,N_17487,N_17437);
or U21102 (N_21102,N_15807,N_18539);
nand U21103 (N_21103,N_18216,N_17884);
nor U21104 (N_21104,N_16204,N_17055);
nor U21105 (N_21105,N_17882,N_18171);
and U21106 (N_21106,N_18646,N_18224);
and U21107 (N_21107,N_16917,N_17994);
nor U21108 (N_21108,N_16193,N_17315);
nand U21109 (N_21109,N_16821,N_17643);
and U21110 (N_21110,N_17122,N_16655);
nand U21111 (N_21111,N_17427,N_17926);
and U21112 (N_21112,N_16851,N_16765);
or U21113 (N_21113,N_18720,N_17506);
nand U21114 (N_21114,N_17522,N_18384);
or U21115 (N_21115,N_18235,N_18161);
nor U21116 (N_21116,N_18733,N_16956);
or U21117 (N_21117,N_16394,N_17762);
nand U21118 (N_21118,N_15649,N_18280);
or U21119 (N_21119,N_15796,N_17778);
or U21120 (N_21120,N_16905,N_15731);
nor U21121 (N_21121,N_16768,N_16438);
and U21122 (N_21122,N_16790,N_16454);
nor U21123 (N_21123,N_17459,N_17470);
or U21124 (N_21124,N_18689,N_15796);
nand U21125 (N_21125,N_16704,N_18173);
nand U21126 (N_21126,N_17940,N_18401);
nand U21127 (N_21127,N_17009,N_16422);
xor U21128 (N_21128,N_16351,N_17085);
or U21129 (N_21129,N_17099,N_18471);
nor U21130 (N_21130,N_18123,N_16835);
nand U21131 (N_21131,N_17584,N_16659);
nor U21132 (N_21132,N_18119,N_17944);
and U21133 (N_21133,N_17010,N_18399);
nand U21134 (N_21134,N_18545,N_18457);
nor U21135 (N_21135,N_18654,N_18029);
and U21136 (N_21136,N_17870,N_18344);
and U21137 (N_21137,N_16507,N_17642);
nor U21138 (N_21138,N_17010,N_16011);
or U21139 (N_21139,N_15803,N_18163);
or U21140 (N_21140,N_17767,N_16858);
and U21141 (N_21141,N_17367,N_17342);
and U21142 (N_21142,N_16801,N_17923);
and U21143 (N_21143,N_18087,N_18723);
nor U21144 (N_21144,N_15951,N_15827);
and U21145 (N_21145,N_16638,N_17673);
nand U21146 (N_21146,N_17353,N_16074);
nand U21147 (N_21147,N_16049,N_17454);
nand U21148 (N_21148,N_15844,N_16002);
nor U21149 (N_21149,N_16242,N_17864);
nor U21150 (N_21150,N_15710,N_17745);
nand U21151 (N_21151,N_18287,N_17571);
nand U21152 (N_21152,N_18483,N_16317);
or U21153 (N_21153,N_16543,N_16880);
or U21154 (N_21154,N_18095,N_17808);
xnor U21155 (N_21155,N_17995,N_18559);
nor U21156 (N_21156,N_16681,N_16990);
xor U21157 (N_21157,N_17065,N_18687);
xnor U21158 (N_21158,N_16412,N_16421);
nor U21159 (N_21159,N_17630,N_18480);
nor U21160 (N_21160,N_17701,N_15636);
nor U21161 (N_21161,N_16121,N_16502);
or U21162 (N_21162,N_18036,N_16390);
or U21163 (N_21163,N_15825,N_16177);
nor U21164 (N_21164,N_17900,N_16743);
or U21165 (N_21165,N_16254,N_16111);
or U21166 (N_21166,N_16480,N_17621);
and U21167 (N_21167,N_17531,N_15962);
or U21168 (N_21168,N_16065,N_18322);
nor U21169 (N_21169,N_18146,N_17930);
xor U21170 (N_21170,N_18631,N_16047);
nand U21171 (N_21171,N_18503,N_18369);
or U21172 (N_21172,N_17372,N_16391);
or U21173 (N_21173,N_17556,N_15670);
or U21174 (N_21174,N_17796,N_18268);
xnor U21175 (N_21175,N_17222,N_16728);
and U21176 (N_21176,N_18351,N_17419);
nor U21177 (N_21177,N_17095,N_18350);
or U21178 (N_21178,N_16615,N_15876);
or U21179 (N_21179,N_18440,N_17743);
nor U21180 (N_21180,N_17203,N_18326);
or U21181 (N_21181,N_16181,N_16409);
xnor U21182 (N_21182,N_17884,N_17355);
nor U21183 (N_21183,N_17500,N_17952);
nand U21184 (N_21184,N_16530,N_16808);
and U21185 (N_21185,N_18045,N_17084);
xor U21186 (N_21186,N_16780,N_16062);
and U21187 (N_21187,N_17534,N_16530);
or U21188 (N_21188,N_18366,N_18488);
nor U21189 (N_21189,N_18201,N_18613);
or U21190 (N_21190,N_18705,N_17874);
xor U21191 (N_21191,N_15943,N_17492);
nand U21192 (N_21192,N_16074,N_18607);
or U21193 (N_21193,N_17613,N_16646);
nand U21194 (N_21194,N_18354,N_16516);
and U21195 (N_21195,N_16216,N_18445);
nor U21196 (N_21196,N_17745,N_15959);
and U21197 (N_21197,N_17546,N_17847);
or U21198 (N_21198,N_17351,N_16964);
nand U21199 (N_21199,N_17409,N_17916);
and U21200 (N_21200,N_17358,N_16367);
nor U21201 (N_21201,N_17646,N_15857);
nor U21202 (N_21202,N_16744,N_17497);
nor U21203 (N_21203,N_16360,N_18422);
nand U21204 (N_21204,N_18651,N_17098);
or U21205 (N_21205,N_16775,N_18518);
or U21206 (N_21206,N_15744,N_17034);
and U21207 (N_21207,N_16961,N_15878);
nor U21208 (N_21208,N_16665,N_15888);
or U21209 (N_21209,N_17010,N_17727);
nor U21210 (N_21210,N_18298,N_18521);
xnor U21211 (N_21211,N_17792,N_17098);
nor U21212 (N_21212,N_17114,N_16506);
and U21213 (N_21213,N_18684,N_16486);
and U21214 (N_21214,N_18044,N_18040);
and U21215 (N_21215,N_17817,N_16313);
or U21216 (N_21216,N_15771,N_17515);
and U21217 (N_21217,N_16022,N_16485);
nor U21218 (N_21218,N_17901,N_18511);
nor U21219 (N_21219,N_17184,N_17595);
and U21220 (N_21220,N_16418,N_16932);
or U21221 (N_21221,N_15765,N_16566);
or U21222 (N_21222,N_16705,N_17051);
xor U21223 (N_21223,N_15987,N_17961);
xnor U21224 (N_21224,N_18691,N_18298);
nor U21225 (N_21225,N_16144,N_16193);
nor U21226 (N_21226,N_16732,N_18187);
and U21227 (N_21227,N_17674,N_16258);
or U21228 (N_21228,N_18635,N_17444);
nor U21229 (N_21229,N_18521,N_16556);
and U21230 (N_21230,N_16383,N_17179);
nand U21231 (N_21231,N_17193,N_15791);
nor U21232 (N_21232,N_17799,N_18487);
or U21233 (N_21233,N_16917,N_18428);
xor U21234 (N_21234,N_17029,N_18414);
nor U21235 (N_21235,N_15700,N_17426);
xnor U21236 (N_21236,N_16919,N_18217);
or U21237 (N_21237,N_17770,N_16013);
xnor U21238 (N_21238,N_15856,N_16504);
and U21239 (N_21239,N_16334,N_17283);
and U21240 (N_21240,N_17182,N_16293);
and U21241 (N_21241,N_18275,N_17105);
xor U21242 (N_21242,N_17563,N_17122);
and U21243 (N_21243,N_16920,N_16978);
nand U21244 (N_21244,N_17141,N_18217);
nand U21245 (N_21245,N_16470,N_18716);
xor U21246 (N_21246,N_15929,N_16371);
xor U21247 (N_21247,N_17511,N_18121);
and U21248 (N_21248,N_17920,N_17883);
nor U21249 (N_21249,N_17902,N_15995);
nor U21250 (N_21250,N_16028,N_16763);
and U21251 (N_21251,N_16093,N_18202);
nor U21252 (N_21252,N_16735,N_17910);
nand U21253 (N_21253,N_17142,N_18079);
nor U21254 (N_21254,N_16564,N_18347);
xor U21255 (N_21255,N_15873,N_18554);
nor U21256 (N_21256,N_16529,N_18378);
nand U21257 (N_21257,N_18359,N_18183);
nor U21258 (N_21258,N_18651,N_18630);
xnor U21259 (N_21259,N_17438,N_17324);
or U21260 (N_21260,N_18272,N_18653);
nor U21261 (N_21261,N_17462,N_18656);
nor U21262 (N_21262,N_18145,N_15743);
nand U21263 (N_21263,N_17065,N_16416);
nand U21264 (N_21264,N_18595,N_18479);
nand U21265 (N_21265,N_17269,N_16854);
nand U21266 (N_21266,N_18217,N_16161);
nand U21267 (N_21267,N_16860,N_18530);
nand U21268 (N_21268,N_16085,N_18411);
nor U21269 (N_21269,N_15746,N_16597);
and U21270 (N_21270,N_16821,N_17434);
nor U21271 (N_21271,N_15952,N_16903);
and U21272 (N_21272,N_18164,N_16443);
xor U21273 (N_21273,N_16829,N_15834);
nor U21274 (N_21274,N_17970,N_18420);
and U21275 (N_21275,N_18353,N_17816);
and U21276 (N_21276,N_18014,N_17366);
nor U21277 (N_21277,N_18106,N_16387);
nor U21278 (N_21278,N_16005,N_18683);
xor U21279 (N_21279,N_16437,N_17456);
nor U21280 (N_21280,N_16936,N_15870);
nor U21281 (N_21281,N_18527,N_16572);
or U21282 (N_21282,N_17630,N_18486);
or U21283 (N_21283,N_17300,N_18482);
or U21284 (N_21284,N_15847,N_16679);
xnor U21285 (N_21285,N_16750,N_15922);
and U21286 (N_21286,N_16236,N_17902);
nand U21287 (N_21287,N_16217,N_18221);
nor U21288 (N_21288,N_16833,N_17527);
nand U21289 (N_21289,N_17593,N_18273);
and U21290 (N_21290,N_15947,N_17644);
and U21291 (N_21291,N_17265,N_18584);
nor U21292 (N_21292,N_15796,N_17244);
nor U21293 (N_21293,N_16224,N_17701);
or U21294 (N_21294,N_17354,N_15775);
xor U21295 (N_21295,N_17047,N_17312);
nand U21296 (N_21296,N_15975,N_16400);
nand U21297 (N_21297,N_18599,N_18449);
and U21298 (N_21298,N_16878,N_16590);
and U21299 (N_21299,N_17435,N_17156);
nor U21300 (N_21300,N_18595,N_16764);
nor U21301 (N_21301,N_16572,N_16282);
or U21302 (N_21302,N_18220,N_15634);
and U21303 (N_21303,N_17782,N_16105);
and U21304 (N_21304,N_18327,N_18049);
nand U21305 (N_21305,N_17064,N_17094);
and U21306 (N_21306,N_16952,N_17402);
nand U21307 (N_21307,N_16376,N_16120);
nor U21308 (N_21308,N_15803,N_18433);
or U21309 (N_21309,N_17778,N_16757);
nor U21310 (N_21310,N_18034,N_18195);
nand U21311 (N_21311,N_16289,N_17123);
nand U21312 (N_21312,N_17517,N_16426);
nor U21313 (N_21313,N_17578,N_16744);
nor U21314 (N_21314,N_17875,N_17903);
nand U21315 (N_21315,N_18247,N_16746);
nand U21316 (N_21316,N_18296,N_18621);
xor U21317 (N_21317,N_15768,N_16221);
nand U21318 (N_21318,N_17056,N_16127);
nor U21319 (N_21319,N_16866,N_15964);
nor U21320 (N_21320,N_15903,N_18501);
or U21321 (N_21321,N_17294,N_17983);
nand U21322 (N_21322,N_17279,N_17338);
or U21323 (N_21323,N_17400,N_18185);
or U21324 (N_21324,N_18085,N_15770);
and U21325 (N_21325,N_18587,N_16641);
or U21326 (N_21326,N_16152,N_18519);
nor U21327 (N_21327,N_16548,N_15851);
nand U21328 (N_21328,N_16419,N_17392);
nand U21329 (N_21329,N_16022,N_16529);
or U21330 (N_21330,N_16305,N_17822);
and U21331 (N_21331,N_16521,N_17684);
and U21332 (N_21332,N_16982,N_18501);
nor U21333 (N_21333,N_18183,N_17790);
or U21334 (N_21334,N_16200,N_17757);
nand U21335 (N_21335,N_15704,N_18160);
or U21336 (N_21336,N_18014,N_16255);
or U21337 (N_21337,N_16941,N_16032);
and U21338 (N_21338,N_16192,N_16536);
xnor U21339 (N_21339,N_15890,N_17621);
and U21340 (N_21340,N_16320,N_16392);
nand U21341 (N_21341,N_18559,N_17818);
nand U21342 (N_21342,N_18369,N_15885);
nor U21343 (N_21343,N_16842,N_16017);
xnor U21344 (N_21344,N_16261,N_17168);
or U21345 (N_21345,N_16050,N_16817);
and U21346 (N_21346,N_16446,N_16064);
or U21347 (N_21347,N_16785,N_15658);
nor U21348 (N_21348,N_18495,N_16068);
nor U21349 (N_21349,N_17664,N_18070);
nor U21350 (N_21350,N_16846,N_15741);
and U21351 (N_21351,N_17715,N_16372);
or U21352 (N_21352,N_18092,N_17680);
nor U21353 (N_21353,N_17553,N_18709);
nand U21354 (N_21354,N_18667,N_17202);
nand U21355 (N_21355,N_16387,N_15976);
nor U21356 (N_21356,N_15843,N_18035);
or U21357 (N_21357,N_16089,N_15983);
or U21358 (N_21358,N_16608,N_18426);
nor U21359 (N_21359,N_17469,N_18671);
nand U21360 (N_21360,N_17289,N_18625);
and U21361 (N_21361,N_17005,N_16293);
nand U21362 (N_21362,N_17133,N_17122);
nor U21363 (N_21363,N_17418,N_17150);
nor U21364 (N_21364,N_15655,N_15943);
or U21365 (N_21365,N_18339,N_17811);
nand U21366 (N_21366,N_16508,N_16502);
nor U21367 (N_21367,N_15829,N_16445);
and U21368 (N_21368,N_16283,N_16336);
or U21369 (N_21369,N_18615,N_16561);
or U21370 (N_21370,N_17249,N_18414);
nand U21371 (N_21371,N_17729,N_17042);
and U21372 (N_21372,N_18664,N_17491);
or U21373 (N_21373,N_17465,N_16242);
or U21374 (N_21374,N_17382,N_18525);
xnor U21375 (N_21375,N_16564,N_15727);
nand U21376 (N_21376,N_17811,N_17413);
nand U21377 (N_21377,N_17225,N_17884);
nand U21378 (N_21378,N_15625,N_18404);
nor U21379 (N_21379,N_18727,N_18212);
and U21380 (N_21380,N_16578,N_15981);
or U21381 (N_21381,N_17632,N_17025);
and U21382 (N_21382,N_16173,N_18628);
nor U21383 (N_21383,N_17498,N_16456);
nand U21384 (N_21384,N_16412,N_17980);
nand U21385 (N_21385,N_17122,N_17130);
or U21386 (N_21386,N_17216,N_16617);
and U21387 (N_21387,N_18100,N_17513);
nor U21388 (N_21388,N_15822,N_18024);
nand U21389 (N_21389,N_17605,N_16498);
nor U21390 (N_21390,N_17606,N_17609);
nand U21391 (N_21391,N_15887,N_16769);
nand U21392 (N_21392,N_18065,N_16080);
nor U21393 (N_21393,N_16862,N_18704);
or U21394 (N_21394,N_18272,N_17797);
and U21395 (N_21395,N_15775,N_17044);
nor U21396 (N_21396,N_16549,N_16941);
and U21397 (N_21397,N_16661,N_15993);
and U21398 (N_21398,N_17942,N_15628);
or U21399 (N_21399,N_16325,N_16729);
xnor U21400 (N_21400,N_17143,N_16289);
nor U21401 (N_21401,N_17100,N_17162);
nand U21402 (N_21402,N_16462,N_16106);
or U21403 (N_21403,N_16248,N_16979);
xnor U21404 (N_21404,N_16813,N_16482);
nor U21405 (N_21405,N_17599,N_17682);
and U21406 (N_21406,N_17815,N_16213);
xor U21407 (N_21407,N_17473,N_16042);
nand U21408 (N_21408,N_18741,N_17447);
nor U21409 (N_21409,N_18008,N_18017);
xor U21410 (N_21410,N_18346,N_15882);
nand U21411 (N_21411,N_17551,N_16511);
nand U21412 (N_21412,N_17534,N_17006);
nor U21413 (N_21413,N_17662,N_16154);
nor U21414 (N_21414,N_16859,N_16326);
and U21415 (N_21415,N_16344,N_17555);
nor U21416 (N_21416,N_16149,N_16945);
nor U21417 (N_21417,N_16834,N_16805);
nor U21418 (N_21418,N_15957,N_16261);
or U21419 (N_21419,N_15949,N_18491);
or U21420 (N_21420,N_17976,N_16839);
and U21421 (N_21421,N_18165,N_16888);
nand U21422 (N_21422,N_17234,N_17655);
or U21423 (N_21423,N_16846,N_17857);
xor U21424 (N_21424,N_16788,N_18392);
nor U21425 (N_21425,N_18258,N_18547);
nor U21426 (N_21426,N_17171,N_16118);
and U21427 (N_21427,N_18456,N_18525);
nor U21428 (N_21428,N_16984,N_15731);
or U21429 (N_21429,N_17232,N_17486);
nor U21430 (N_21430,N_16105,N_17615);
or U21431 (N_21431,N_16797,N_18186);
nand U21432 (N_21432,N_17125,N_18366);
nor U21433 (N_21433,N_17407,N_17614);
and U21434 (N_21434,N_18463,N_18647);
and U21435 (N_21435,N_18635,N_17122);
nor U21436 (N_21436,N_17128,N_16126);
and U21437 (N_21437,N_16804,N_16678);
and U21438 (N_21438,N_17815,N_17447);
xor U21439 (N_21439,N_15850,N_18463);
and U21440 (N_21440,N_17476,N_16991);
nor U21441 (N_21441,N_15670,N_18542);
nand U21442 (N_21442,N_18072,N_18029);
or U21443 (N_21443,N_16899,N_17228);
and U21444 (N_21444,N_18725,N_17587);
nor U21445 (N_21445,N_15627,N_18370);
and U21446 (N_21446,N_17238,N_15908);
or U21447 (N_21447,N_15638,N_18362);
and U21448 (N_21448,N_17536,N_17685);
xnor U21449 (N_21449,N_17652,N_16840);
or U21450 (N_21450,N_17865,N_17001);
and U21451 (N_21451,N_18370,N_17651);
or U21452 (N_21452,N_15681,N_15635);
or U21453 (N_21453,N_15720,N_17993);
xor U21454 (N_21454,N_16374,N_16451);
and U21455 (N_21455,N_17661,N_18602);
or U21456 (N_21456,N_16045,N_18628);
and U21457 (N_21457,N_17327,N_17456);
nor U21458 (N_21458,N_17582,N_18587);
xnor U21459 (N_21459,N_15637,N_18586);
xor U21460 (N_21460,N_18732,N_18458);
xor U21461 (N_21461,N_15807,N_15784);
or U21462 (N_21462,N_17056,N_15848);
nor U21463 (N_21463,N_16714,N_16820);
nand U21464 (N_21464,N_17440,N_16786);
or U21465 (N_21465,N_17888,N_18038);
nor U21466 (N_21466,N_16997,N_16289);
xnor U21467 (N_21467,N_18493,N_17453);
nand U21468 (N_21468,N_18731,N_15878);
nor U21469 (N_21469,N_16676,N_15705);
or U21470 (N_21470,N_18053,N_18341);
nor U21471 (N_21471,N_17235,N_16531);
or U21472 (N_21472,N_18328,N_18082);
nor U21473 (N_21473,N_16211,N_18480);
nand U21474 (N_21474,N_16233,N_16513);
nand U21475 (N_21475,N_16807,N_16177);
nand U21476 (N_21476,N_17046,N_16701);
and U21477 (N_21477,N_16759,N_17697);
or U21478 (N_21478,N_16527,N_18524);
and U21479 (N_21479,N_15962,N_15737);
and U21480 (N_21480,N_16315,N_17856);
nand U21481 (N_21481,N_18132,N_16360);
xor U21482 (N_21482,N_18218,N_17305);
or U21483 (N_21483,N_17933,N_17978);
nor U21484 (N_21484,N_18601,N_16417);
and U21485 (N_21485,N_16764,N_17245);
nor U21486 (N_21486,N_18387,N_18240);
or U21487 (N_21487,N_15736,N_16939);
or U21488 (N_21488,N_15818,N_17344);
and U21489 (N_21489,N_17063,N_15947);
nor U21490 (N_21490,N_16146,N_15755);
nand U21491 (N_21491,N_18197,N_18508);
xnor U21492 (N_21492,N_16853,N_17063);
or U21493 (N_21493,N_15679,N_17877);
nand U21494 (N_21494,N_15682,N_18167);
nand U21495 (N_21495,N_17368,N_17939);
nand U21496 (N_21496,N_15825,N_15729);
and U21497 (N_21497,N_18437,N_16900);
nor U21498 (N_21498,N_18357,N_18312);
or U21499 (N_21499,N_17429,N_15884);
and U21500 (N_21500,N_16295,N_17666);
nand U21501 (N_21501,N_16949,N_17814);
nor U21502 (N_21502,N_16456,N_17998);
nor U21503 (N_21503,N_18577,N_15823);
or U21504 (N_21504,N_17692,N_15999);
or U21505 (N_21505,N_16290,N_17987);
and U21506 (N_21506,N_16551,N_16561);
and U21507 (N_21507,N_17350,N_16537);
nor U21508 (N_21508,N_17744,N_16664);
and U21509 (N_21509,N_15867,N_16198);
or U21510 (N_21510,N_15756,N_17290);
and U21511 (N_21511,N_17859,N_16533);
or U21512 (N_21512,N_18291,N_17919);
nand U21513 (N_21513,N_18620,N_17680);
nor U21514 (N_21514,N_18616,N_17871);
nand U21515 (N_21515,N_17231,N_16715);
and U21516 (N_21516,N_15631,N_17145);
nand U21517 (N_21517,N_15916,N_18341);
nor U21518 (N_21518,N_17399,N_16822);
and U21519 (N_21519,N_15895,N_18185);
or U21520 (N_21520,N_17767,N_17164);
and U21521 (N_21521,N_18042,N_16212);
nor U21522 (N_21522,N_16176,N_16662);
or U21523 (N_21523,N_17465,N_17389);
nor U21524 (N_21524,N_17274,N_16691);
xnor U21525 (N_21525,N_18064,N_15684);
or U21526 (N_21526,N_15971,N_17951);
and U21527 (N_21527,N_17335,N_18011);
or U21528 (N_21528,N_16225,N_15833);
and U21529 (N_21529,N_17115,N_16011);
nor U21530 (N_21530,N_17502,N_16648);
and U21531 (N_21531,N_18664,N_16992);
or U21532 (N_21532,N_16553,N_18016);
xnor U21533 (N_21533,N_16442,N_16832);
nor U21534 (N_21534,N_18278,N_18121);
nand U21535 (N_21535,N_15877,N_18473);
or U21536 (N_21536,N_16165,N_18234);
xnor U21537 (N_21537,N_15879,N_16740);
nor U21538 (N_21538,N_16733,N_17926);
nand U21539 (N_21539,N_15884,N_17969);
and U21540 (N_21540,N_15687,N_18585);
nand U21541 (N_21541,N_17480,N_15709);
xor U21542 (N_21542,N_16735,N_15799);
or U21543 (N_21543,N_18469,N_16085);
nand U21544 (N_21544,N_16105,N_18492);
xor U21545 (N_21545,N_17274,N_17860);
or U21546 (N_21546,N_15652,N_17959);
and U21547 (N_21547,N_15750,N_17311);
xnor U21548 (N_21548,N_16794,N_17196);
or U21549 (N_21549,N_16753,N_16695);
and U21550 (N_21550,N_17730,N_16189);
or U21551 (N_21551,N_18483,N_17453);
or U21552 (N_21552,N_16353,N_16296);
and U21553 (N_21553,N_16429,N_18336);
xor U21554 (N_21554,N_17456,N_15657);
and U21555 (N_21555,N_15634,N_16761);
and U21556 (N_21556,N_15947,N_16811);
xnor U21557 (N_21557,N_16491,N_15760);
xor U21558 (N_21558,N_17634,N_16233);
nand U21559 (N_21559,N_17444,N_18112);
nand U21560 (N_21560,N_18270,N_17133);
nand U21561 (N_21561,N_17905,N_18399);
and U21562 (N_21562,N_17306,N_18364);
nand U21563 (N_21563,N_15653,N_18296);
or U21564 (N_21564,N_15838,N_16113);
and U21565 (N_21565,N_16309,N_17541);
nor U21566 (N_21566,N_17490,N_18438);
or U21567 (N_21567,N_15774,N_16168);
nand U21568 (N_21568,N_16976,N_17561);
and U21569 (N_21569,N_16254,N_17945);
or U21570 (N_21570,N_18402,N_18171);
nand U21571 (N_21571,N_16590,N_17661);
and U21572 (N_21572,N_15662,N_18099);
and U21573 (N_21573,N_16721,N_17955);
xnor U21574 (N_21574,N_18655,N_16529);
and U21575 (N_21575,N_15957,N_15882);
nand U21576 (N_21576,N_15877,N_17207);
nor U21577 (N_21577,N_17875,N_17931);
or U21578 (N_21578,N_17725,N_16144);
nand U21579 (N_21579,N_17775,N_15769);
xor U21580 (N_21580,N_15946,N_15738);
or U21581 (N_21581,N_16067,N_17471);
xnor U21582 (N_21582,N_17305,N_18494);
nor U21583 (N_21583,N_16017,N_17646);
or U21584 (N_21584,N_16479,N_17882);
or U21585 (N_21585,N_15877,N_17454);
or U21586 (N_21586,N_17538,N_17670);
xor U21587 (N_21587,N_18744,N_17423);
xor U21588 (N_21588,N_17592,N_16176);
xnor U21589 (N_21589,N_15783,N_18425);
and U21590 (N_21590,N_18392,N_17225);
or U21591 (N_21591,N_17564,N_17578);
or U21592 (N_21592,N_16659,N_15983);
nand U21593 (N_21593,N_16679,N_18238);
nand U21594 (N_21594,N_18350,N_18601);
nor U21595 (N_21595,N_18203,N_16269);
or U21596 (N_21596,N_17379,N_18277);
xnor U21597 (N_21597,N_16646,N_18413);
and U21598 (N_21598,N_17326,N_15702);
nand U21599 (N_21599,N_18579,N_16244);
nand U21600 (N_21600,N_16909,N_16741);
and U21601 (N_21601,N_17558,N_16532);
nand U21602 (N_21602,N_15784,N_17287);
nand U21603 (N_21603,N_16004,N_16153);
or U21604 (N_21604,N_18047,N_18056);
or U21605 (N_21605,N_17482,N_18395);
nor U21606 (N_21606,N_17771,N_17133);
and U21607 (N_21607,N_18477,N_16129);
nand U21608 (N_21608,N_17930,N_17450);
nor U21609 (N_21609,N_17917,N_18104);
nor U21610 (N_21610,N_16785,N_16352);
or U21611 (N_21611,N_16581,N_16708);
nand U21612 (N_21612,N_17784,N_16591);
nand U21613 (N_21613,N_17143,N_16630);
and U21614 (N_21614,N_15826,N_17315);
xor U21615 (N_21615,N_16458,N_18538);
or U21616 (N_21616,N_17869,N_17412);
nand U21617 (N_21617,N_17186,N_16202);
or U21618 (N_21618,N_16126,N_17523);
xor U21619 (N_21619,N_15722,N_15991);
nand U21620 (N_21620,N_17661,N_17120);
nand U21621 (N_21621,N_18625,N_18741);
nand U21622 (N_21622,N_16709,N_16253);
or U21623 (N_21623,N_17582,N_17246);
xor U21624 (N_21624,N_15769,N_17812);
and U21625 (N_21625,N_15925,N_17095);
nand U21626 (N_21626,N_16277,N_17872);
nor U21627 (N_21627,N_17883,N_17584);
nor U21628 (N_21628,N_15838,N_18000);
xnor U21629 (N_21629,N_18739,N_18516);
and U21630 (N_21630,N_17678,N_17566);
or U21631 (N_21631,N_16836,N_17283);
or U21632 (N_21632,N_17041,N_16852);
nor U21633 (N_21633,N_17865,N_15782);
xor U21634 (N_21634,N_16013,N_16913);
xnor U21635 (N_21635,N_15828,N_15906);
nor U21636 (N_21636,N_17855,N_16222);
nand U21637 (N_21637,N_18154,N_17499);
and U21638 (N_21638,N_16632,N_16535);
nor U21639 (N_21639,N_16142,N_16952);
nand U21640 (N_21640,N_17325,N_15741);
or U21641 (N_21641,N_17621,N_16366);
or U21642 (N_21642,N_16904,N_16805);
nor U21643 (N_21643,N_17226,N_17478);
and U21644 (N_21644,N_18529,N_16162);
or U21645 (N_21645,N_16321,N_17668);
nor U21646 (N_21646,N_17623,N_16728);
xor U21647 (N_21647,N_16356,N_18276);
and U21648 (N_21648,N_18601,N_17155);
and U21649 (N_21649,N_17595,N_16824);
or U21650 (N_21650,N_16397,N_17914);
nor U21651 (N_21651,N_16135,N_18628);
and U21652 (N_21652,N_17803,N_18082);
and U21653 (N_21653,N_18179,N_18382);
nand U21654 (N_21654,N_16436,N_16423);
nand U21655 (N_21655,N_17513,N_15855);
nand U21656 (N_21656,N_17871,N_18681);
nor U21657 (N_21657,N_18548,N_16832);
and U21658 (N_21658,N_18282,N_17229);
and U21659 (N_21659,N_18046,N_18361);
xnor U21660 (N_21660,N_18282,N_16963);
nand U21661 (N_21661,N_16943,N_15636);
or U21662 (N_21662,N_18435,N_16324);
nand U21663 (N_21663,N_18105,N_17993);
or U21664 (N_21664,N_17403,N_17136);
and U21665 (N_21665,N_15861,N_18196);
and U21666 (N_21666,N_16625,N_16035);
xor U21667 (N_21667,N_16483,N_15900);
or U21668 (N_21668,N_15955,N_16457);
nand U21669 (N_21669,N_18048,N_16687);
nand U21670 (N_21670,N_16622,N_16137);
nand U21671 (N_21671,N_17047,N_16159);
nand U21672 (N_21672,N_17730,N_17506);
nor U21673 (N_21673,N_18371,N_17410);
nand U21674 (N_21674,N_16073,N_17674);
nand U21675 (N_21675,N_18637,N_16750);
or U21676 (N_21676,N_18134,N_16300);
and U21677 (N_21677,N_16614,N_18058);
or U21678 (N_21678,N_18513,N_16899);
or U21679 (N_21679,N_15961,N_16275);
and U21680 (N_21680,N_16637,N_18114);
nand U21681 (N_21681,N_16024,N_17986);
and U21682 (N_21682,N_17784,N_17641);
or U21683 (N_21683,N_17264,N_18689);
and U21684 (N_21684,N_17511,N_15671);
and U21685 (N_21685,N_15931,N_16696);
nor U21686 (N_21686,N_15745,N_17859);
nor U21687 (N_21687,N_16936,N_16660);
nand U21688 (N_21688,N_15943,N_16739);
nand U21689 (N_21689,N_16158,N_17999);
or U21690 (N_21690,N_15817,N_17472);
nor U21691 (N_21691,N_17420,N_16342);
or U21692 (N_21692,N_17989,N_17406);
nand U21693 (N_21693,N_16481,N_16508);
or U21694 (N_21694,N_16575,N_16506);
nand U21695 (N_21695,N_17050,N_18140);
or U21696 (N_21696,N_15698,N_17249);
nor U21697 (N_21697,N_18237,N_17594);
or U21698 (N_21698,N_16464,N_18031);
nand U21699 (N_21699,N_18045,N_16563);
nand U21700 (N_21700,N_15786,N_16869);
and U21701 (N_21701,N_17447,N_16116);
and U21702 (N_21702,N_17676,N_18390);
nand U21703 (N_21703,N_15918,N_16749);
nor U21704 (N_21704,N_16771,N_17945);
nor U21705 (N_21705,N_16533,N_17054);
or U21706 (N_21706,N_18152,N_15818);
or U21707 (N_21707,N_16467,N_17436);
nor U21708 (N_21708,N_17558,N_18699);
and U21709 (N_21709,N_15748,N_18211);
and U21710 (N_21710,N_16276,N_17412);
and U21711 (N_21711,N_16470,N_17819);
and U21712 (N_21712,N_16541,N_15888);
and U21713 (N_21713,N_18746,N_17327);
and U21714 (N_21714,N_17743,N_16673);
and U21715 (N_21715,N_16636,N_17574);
nor U21716 (N_21716,N_18169,N_15678);
xor U21717 (N_21717,N_17167,N_16540);
and U21718 (N_21718,N_16820,N_18318);
nor U21719 (N_21719,N_18233,N_16798);
or U21720 (N_21720,N_17166,N_15916);
xnor U21721 (N_21721,N_17329,N_18636);
nand U21722 (N_21722,N_18060,N_16995);
or U21723 (N_21723,N_17122,N_17988);
and U21724 (N_21724,N_18566,N_17944);
nor U21725 (N_21725,N_18710,N_16143);
or U21726 (N_21726,N_16869,N_18549);
nor U21727 (N_21727,N_15787,N_18173);
and U21728 (N_21728,N_17874,N_16754);
nand U21729 (N_21729,N_16394,N_17768);
nor U21730 (N_21730,N_16733,N_16105);
nor U21731 (N_21731,N_16852,N_16223);
or U21732 (N_21732,N_16500,N_17703);
or U21733 (N_21733,N_16609,N_16361);
nand U21734 (N_21734,N_17291,N_18168);
and U21735 (N_21735,N_17130,N_17465);
nor U21736 (N_21736,N_18387,N_15719);
nor U21737 (N_21737,N_17990,N_16551);
or U21738 (N_21738,N_17092,N_16152);
nor U21739 (N_21739,N_16996,N_18330);
or U21740 (N_21740,N_18494,N_18462);
nand U21741 (N_21741,N_18418,N_18598);
nor U21742 (N_21742,N_16522,N_15949);
and U21743 (N_21743,N_18700,N_17025);
nor U21744 (N_21744,N_16221,N_16203);
nand U21745 (N_21745,N_17360,N_18646);
and U21746 (N_21746,N_16814,N_18286);
nand U21747 (N_21747,N_15747,N_18203);
xor U21748 (N_21748,N_17422,N_18252);
xor U21749 (N_21749,N_17460,N_17313);
xnor U21750 (N_21750,N_17163,N_15981);
nor U21751 (N_21751,N_17074,N_18302);
or U21752 (N_21752,N_16875,N_17341);
nor U21753 (N_21753,N_16938,N_17291);
and U21754 (N_21754,N_16686,N_18596);
nor U21755 (N_21755,N_17888,N_15662);
nor U21756 (N_21756,N_16735,N_16107);
nor U21757 (N_21757,N_18491,N_17750);
or U21758 (N_21758,N_16538,N_15645);
nand U21759 (N_21759,N_16601,N_16139);
nor U21760 (N_21760,N_18481,N_16708);
or U21761 (N_21761,N_17299,N_16979);
nor U21762 (N_21762,N_16904,N_18459);
nor U21763 (N_21763,N_15823,N_17426);
or U21764 (N_21764,N_17749,N_15721);
nand U21765 (N_21765,N_16207,N_17144);
and U21766 (N_21766,N_18730,N_17748);
nand U21767 (N_21767,N_17217,N_17286);
or U21768 (N_21768,N_16959,N_18021);
and U21769 (N_21769,N_16267,N_17629);
nand U21770 (N_21770,N_17555,N_16175);
xnor U21771 (N_21771,N_16959,N_18638);
nand U21772 (N_21772,N_17220,N_16123);
nand U21773 (N_21773,N_17284,N_17613);
nor U21774 (N_21774,N_15983,N_17871);
nand U21775 (N_21775,N_16761,N_16685);
or U21776 (N_21776,N_17569,N_17113);
xor U21777 (N_21777,N_16967,N_18524);
or U21778 (N_21778,N_17061,N_15954);
nand U21779 (N_21779,N_15957,N_16217);
or U21780 (N_21780,N_18502,N_15895);
xnor U21781 (N_21781,N_16489,N_17954);
or U21782 (N_21782,N_18193,N_16706);
xor U21783 (N_21783,N_16093,N_16228);
nor U21784 (N_21784,N_18007,N_17905);
nand U21785 (N_21785,N_17357,N_18253);
nand U21786 (N_21786,N_15972,N_16878);
or U21787 (N_21787,N_18569,N_15969);
nor U21788 (N_21788,N_16887,N_16043);
nand U21789 (N_21789,N_17981,N_16390);
nand U21790 (N_21790,N_17557,N_16588);
xnor U21791 (N_21791,N_16914,N_18452);
nor U21792 (N_21792,N_17039,N_17469);
or U21793 (N_21793,N_18217,N_18486);
and U21794 (N_21794,N_17882,N_17337);
nor U21795 (N_21795,N_17038,N_17293);
or U21796 (N_21796,N_18732,N_17149);
nor U21797 (N_21797,N_16282,N_17578);
or U21798 (N_21798,N_17076,N_17496);
nor U21799 (N_21799,N_18236,N_16319);
xnor U21800 (N_21800,N_15960,N_16168);
or U21801 (N_21801,N_18253,N_17956);
xor U21802 (N_21802,N_16871,N_16040);
nand U21803 (N_21803,N_17840,N_15821);
or U21804 (N_21804,N_16401,N_16950);
and U21805 (N_21805,N_16164,N_15995);
nor U21806 (N_21806,N_17190,N_17775);
nand U21807 (N_21807,N_16792,N_16219);
and U21808 (N_21808,N_15808,N_16839);
nor U21809 (N_21809,N_16025,N_15900);
nor U21810 (N_21810,N_18360,N_15951);
or U21811 (N_21811,N_17232,N_17093);
nand U21812 (N_21812,N_16023,N_18120);
or U21813 (N_21813,N_16882,N_17059);
or U21814 (N_21814,N_17793,N_17198);
or U21815 (N_21815,N_17540,N_16457);
or U21816 (N_21816,N_18744,N_18060);
nand U21817 (N_21817,N_16542,N_16964);
and U21818 (N_21818,N_18080,N_16735);
nor U21819 (N_21819,N_17107,N_16754);
and U21820 (N_21820,N_17451,N_18351);
or U21821 (N_21821,N_18034,N_16584);
or U21822 (N_21822,N_16636,N_16986);
nor U21823 (N_21823,N_16650,N_18023);
xnor U21824 (N_21824,N_17280,N_17506);
and U21825 (N_21825,N_15974,N_17155);
xor U21826 (N_21826,N_17316,N_18337);
nor U21827 (N_21827,N_17301,N_17662);
nor U21828 (N_21828,N_18063,N_18436);
or U21829 (N_21829,N_15640,N_18006);
or U21830 (N_21830,N_17001,N_18635);
xor U21831 (N_21831,N_18642,N_18674);
or U21832 (N_21832,N_17759,N_16218);
nand U21833 (N_21833,N_17201,N_18106);
nand U21834 (N_21834,N_17877,N_17197);
nor U21835 (N_21835,N_16465,N_17909);
xnor U21836 (N_21836,N_16508,N_16374);
nand U21837 (N_21837,N_17431,N_16128);
and U21838 (N_21838,N_16611,N_16170);
or U21839 (N_21839,N_16210,N_15775);
xor U21840 (N_21840,N_15930,N_15997);
nand U21841 (N_21841,N_17533,N_16255);
or U21842 (N_21842,N_17556,N_17239);
or U21843 (N_21843,N_17852,N_18102);
nand U21844 (N_21844,N_18077,N_16013);
nor U21845 (N_21845,N_18191,N_17629);
xor U21846 (N_21846,N_17229,N_17537);
and U21847 (N_21847,N_17916,N_17396);
and U21848 (N_21848,N_16128,N_18338);
and U21849 (N_21849,N_16664,N_17551);
nor U21850 (N_21850,N_18402,N_15709);
and U21851 (N_21851,N_18269,N_18562);
and U21852 (N_21852,N_17131,N_16367);
nor U21853 (N_21853,N_17859,N_16481);
nor U21854 (N_21854,N_17396,N_18394);
or U21855 (N_21855,N_16992,N_17013);
nand U21856 (N_21856,N_18453,N_17999);
xor U21857 (N_21857,N_17854,N_17965);
xor U21858 (N_21858,N_16317,N_15744);
nor U21859 (N_21859,N_16756,N_16570);
nand U21860 (N_21860,N_15747,N_17865);
nor U21861 (N_21861,N_18263,N_17268);
and U21862 (N_21862,N_17550,N_17073);
nand U21863 (N_21863,N_16475,N_17465);
nand U21864 (N_21864,N_17714,N_16840);
nor U21865 (N_21865,N_16267,N_16853);
and U21866 (N_21866,N_17066,N_17908);
nor U21867 (N_21867,N_16717,N_18171);
nand U21868 (N_21868,N_18132,N_17350);
nand U21869 (N_21869,N_18655,N_17849);
nand U21870 (N_21870,N_17738,N_16103);
nand U21871 (N_21871,N_17387,N_18685);
and U21872 (N_21872,N_17807,N_18235);
nor U21873 (N_21873,N_17761,N_18376);
or U21874 (N_21874,N_18362,N_17442);
xor U21875 (N_21875,N_19840,N_19345);
nand U21876 (N_21876,N_21758,N_21714);
nor U21877 (N_21877,N_18783,N_21302);
nand U21878 (N_21878,N_20564,N_20499);
xnor U21879 (N_21879,N_21207,N_19419);
xor U21880 (N_21880,N_19178,N_20467);
nor U21881 (N_21881,N_18926,N_19738);
or U21882 (N_21882,N_19444,N_21501);
nor U21883 (N_21883,N_20038,N_20712);
nand U21884 (N_21884,N_19778,N_18979);
and U21885 (N_21885,N_19571,N_19906);
and U21886 (N_21886,N_19295,N_21829);
and U21887 (N_21887,N_19651,N_19940);
nand U21888 (N_21888,N_20341,N_19806);
and U21889 (N_21889,N_20761,N_21414);
xnor U21890 (N_21890,N_19889,N_21103);
xor U21891 (N_21891,N_20222,N_19809);
nand U21892 (N_21892,N_20822,N_21323);
and U21893 (N_21893,N_18974,N_20209);
xor U21894 (N_21894,N_20674,N_20690);
nand U21895 (N_21895,N_19144,N_19274);
nor U21896 (N_21896,N_19681,N_21218);
or U21897 (N_21897,N_19740,N_21183);
and U21898 (N_21898,N_19358,N_21263);
nand U21899 (N_21899,N_21299,N_21461);
nand U21900 (N_21900,N_20724,N_21537);
nor U21901 (N_21901,N_19500,N_19510);
xnor U21902 (N_21902,N_21647,N_19393);
xor U21903 (N_21903,N_21097,N_20930);
and U21904 (N_21904,N_18796,N_21431);
nand U21905 (N_21905,N_21617,N_19316);
and U21906 (N_21906,N_20161,N_20884);
and U21907 (N_21907,N_19464,N_21716);
nor U21908 (N_21908,N_21860,N_20781);
xor U21909 (N_21909,N_21707,N_19229);
or U21910 (N_21910,N_20278,N_21249);
nor U21911 (N_21911,N_18860,N_19818);
or U21912 (N_21912,N_20173,N_21834);
nor U21913 (N_21913,N_20502,N_20292);
xnor U21914 (N_21914,N_18751,N_19783);
nor U21915 (N_21915,N_19534,N_21423);
nor U21916 (N_21916,N_20907,N_20892);
or U21917 (N_21917,N_20537,N_21418);
or U21918 (N_21918,N_21490,N_19607);
nor U21919 (N_21919,N_19337,N_19196);
nand U21920 (N_21920,N_18940,N_19282);
nand U21921 (N_21921,N_21228,N_21402);
and U21922 (N_21922,N_20236,N_21140);
nor U21923 (N_21923,N_21477,N_21327);
and U21924 (N_21924,N_18971,N_19433);
xor U21925 (N_21925,N_19851,N_21099);
or U21926 (N_21926,N_21870,N_19844);
nand U21927 (N_21927,N_21817,N_19080);
and U21928 (N_21928,N_21050,N_18970);
or U21929 (N_21929,N_19952,N_19539);
nor U21930 (N_21930,N_20858,N_19453);
and U21931 (N_21931,N_20333,N_21400);
xor U21932 (N_21932,N_20553,N_21137);
nand U21933 (N_21933,N_21457,N_19710);
nand U21934 (N_21934,N_21657,N_19723);
nor U21935 (N_21935,N_21038,N_20993);
or U21936 (N_21936,N_20691,N_20729);
nand U21937 (N_21937,N_21417,N_19614);
nand U21938 (N_21938,N_21086,N_20579);
xor U21939 (N_21939,N_19819,N_19114);
xor U21940 (N_21940,N_21795,N_20381);
nand U21941 (N_21941,N_21363,N_19276);
nand U21942 (N_21942,N_21138,N_20475);
or U21943 (N_21943,N_19373,N_21284);
or U21944 (N_21944,N_21694,N_20626);
or U21945 (N_21945,N_19149,N_19252);
or U21946 (N_21946,N_21648,N_19175);
nand U21947 (N_21947,N_20837,N_21724);
nand U21948 (N_21948,N_19777,N_19462);
and U21949 (N_21949,N_20082,N_18877);
nor U21950 (N_21950,N_19645,N_21785);
and U21951 (N_21951,N_20942,N_19918);
nand U21952 (N_21952,N_19027,N_21411);
or U21953 (N_21953,N_20565,N_20665);
nand U21954 (N_21954,N_19850,N_21736);
or U21955 (N_21955,N_21008,N_21229);
and U21956 (N_21956,N_21010,N_19398);
xor U21957 (N_21957,N_19306,N_20253);
nor U21958 (N_21958,N_19064,N_21822);
nand U21959 (N_21959,N_21389,N_19245);
nor U21960 (N_21960,N_19468,N_21452);
nand U21961 (N_21961,N_21044,N_20747);
or U21962 (N_21962,N_20523,N_21230);
nor U21963 (N_21963,N_20067,N_21326);
or U21964 (N_21964,N_21799,N_20142);
nor U21965 (N_21965,N_21342,N_21238);
or U21966 (N_21966,N_20198,N_20513);
and U21967 (N_21967,N_20969,N_21282);
nand U21968 (N_21968,N_19670,N_21319);
or U21969 (N_21969,N_20768,N_18827);
or U21970 (N_21970,N_20493,N_19895);
nand U21971 (N_21971,N_21195,N_20262);
nand U21972 (N_21972,N_21126,N_20979);
nand U21973 (N_21973,N_20878,N_21114);
nand U21974 (N_21974,N_20807,N_19982);
nand U21975 (N_21975,N_20752,N_20977);
or U21976 (N_21976,N_18881,N_21318);
or U21977 (N_21977,N_20051,N_20189);
and U21978 (N_21978,N_20025,N_18938);
or U21979 (N_21979,N_20211,N_20525);
or U21980 (N_21980,N_19097,N_21732);
nor U21981 (N_21981,N_19516,N_21051);
nand U21982 (N_21982,N_19112,N_20479);
or U21983 (N_21983,N_19056,N_20461);
nand U21984 (N_21984,N_20370,N_20149);
or U21985 (N_21985,N_19242,N_19969);
and U21986 (N_21986,N_20423,N_20938);
nand U21987 (N_21987,N_20257,N_18954);
nand U21988 (N_21988,N_20451,N_20687);
or U21989 (N_21989,N_21059,N_20744);
or U21990 (N_21990,N_20374,N_19101);
nand U21991 (N_21991,N_19440,N_19380);
xor U21992 (N_21992,N_21562,N_20542);
and U21993 (N_21993,N_20965,N_20304);
nand U21994 (N_21994,N_21488,N_19221);
and U21995 (N_21995,N_21508,N_20489);
or U21996 (N_21996,N_19737,N_21035);
or U21997 (N_21997,N_19300,N_19362);
or U21998 (N_21998,N_20165,N_21200);
and U21999 (N_21999,N_20477,N_21854);
or U22000 (N_22000,N_21046,N_21398);
nor U22001 (N_22001,N_18843,N_20442);
and U22002 (N_22002,N_20737,N_19456);
xnor U22003 (N_22003,N_20995,N_19567);
and U22004 (N_22004,N_21320,N_21330);
or U22005 (N_22005,N_18917,N_19657);
nand U22006 (N_22006,N_21243,N_19622);
nor U22007 (N_22007,N_18785,N_21026);
and U22008 (N_22008,N_20345,N_19547);
nor U22009 (N_22009,N_20599,N_20195);
nor U22010 (N_22010,N_19794,N_19824);
or U22011 (N_22011,N_20830,N_19748);
and U22012 (N_22012,N_20091,N_21312);
or U22013 (N_22013,N_21575,N_18956);
nand U22014 (N_22014,N_19963,N_20355);
nand U22015 (N_22015,N_19105,N_20206);
and U22016 (N_22016,N_20642,N_21491);
nand U22017 (N_22017,N_20276,N_21394);
and U22018 (N_22018,N_20934,N_19275);
or U22019 (N_22019,N_21281,N_20436);
nor U22020 (N_22020,N_21703,N_19003);
nand U22021 (N_22021,N_19726,N_21741);
or U22022 (N_22022,N_18951,N_21237);
nand U22023 (N_22023,N_21679,N_20678);
and U22024 (N_22024,N_20433,N_19368);
or U22025 (N_22025,N_18975,N_21427);
and U22026 (N_22026,N_21581,N_20032);
nand U22027 (N_22027,N_21075,N_20462);
or U22028 (N_22028,N_19904,N_19074);
or U22029 (N_22029,N_21310,N_21467);
nand U22030 (N_22030,N_21279,N_20087);
or U22031 (N_22031,N_18855,N_20578);
nor U22032 (N_22032,N_21025,N_19503);
or U22033 (N_22033,N_20793,N_20816);
nor U22034 (N_22034,N_19210,N_21015);
or U22035 (N_22035,N_19513,N_20920);
and U22036 (N_22036,N_21801,N_21698);
or U22037 (N_22037,N_20636,N_19529);
nor U22038 (N_22038,N_20811,N_21303);
nor U22039 (N_22039,N_20193,N_19587);
nor U22040 (N_22040,N_20702,N_19219);
and U22041 (N_22041,N_21609,N_19787);
and U22042 (N_22042,N_18905,N_20071);
and U22043 (N_22043,N_21864,N_21257);
or U22044 (N_22044,N_21256,N_21278);
or U22045 (N_22045,N_21524,N_21123);
and U22046 (N_22046,N_20365,N_20283);
or U22047 (N_22047,N_19448,N_21840);
and U22048 (N_22048,N_19744,N_21831);
and U22049 (N_22049,N_19447,N_21339);
and U22050 (N_22050,N_20170,N_21353);
or U22051 (N_22051,N_20711,N_19939);
xnor U22052 (N_22052,N_19304,N_21098);
xor U22053 (N_22053,N_20927,N_19466);
xor U22054 (N_22054,N_21232,N_19664);
nand U22055 (N_22055,N_20758,N_19685);
nor U22056 (N_22056,N_19115,N_19186);
nor U22057 (N_22057,N_21204,N_19881);
or U22058 (N_22058,N_20096,N_20776);
or U22059 (N_22059,N_20814,N_18791);
or U22060 (N_22060,N_18770,N_19404);
or U22061 (N_22061,N_18910,N_21513);
nand U22062 (N_22062,N_18798,N_21317);
xor U22063 (N_22063,N_21573,N_20469);
nor U22064 (N_22064,N_20454,N_19294);
and U22065 (N_22065,N_19153,N_19773);
xor U22066 (N_22066,N_20215,N_18826);
or U22067 (N_22067,N_20728,N_19353);
nor U22068 (N_22068,N_21749,N_21773);
nor U22069 (N_22069,N_19451,N_20673);
or U22070 (N_22070,N_19845,N_20464);
or U22071 (N_22071,N_19649,N_19912);
nand U22072 (N_22072,N_20108,N_20347);
and U22073 (N_22073,N_20414,N_21796);
xnor U22074 (N_22074,N_21246,N_21533);
or U22075 (N_22075,N_21315,N_19564);
nand U22076 (N_22076,N_19790,N_19885);
nand U22077 (N_22077,N_18838,N_21787);
nand U22078 (N_22078,N_21819,N_20901);
nand U22079 (N_22079,N_21780,N_20074);
or U22080 (N_22080,N_20289,N_21376);
or U22081 (N_22081,N_20180,N_18840);
and U22082 (N_22082,N_21135,N_21157);
nor U22083 (N_22083,N_20845,N_19188);
or U22084 (N_22084,N_21553,N_21442);
or U22085 (N_22085,N_21606,N_21045);
or U22086 (N_22086,N_20364,N_19687);
xnor U22087 (N_22087,N_20679,N_21273);
nand U22088 (N_22088,N_20988,N_20548);
nand U22089 (N_22089,N_21753,N_19767);
nor U22090 (N_22090,N_20085,N_18831);
nor U22091 (N_22091,N_20535,N_20006);
nand U22092 (N_22092,N_21636,N_20632);
nand U22093 (N_22093,N_18908,N_18930);
nor U22094 (N_22094,N_20202,N_19619);
nor U22095 (N_22095,N_20321,N_20978);
or U22096 (N_22096,N_20847,N_18807);
xor U22097 (N_22097,N_20270,N_21779);
and U22098 (N_22098,N_21337,N_20771);
nor U22099 (N_22099,N_21776,N_20131);
nor U22100 (N_22100,N_21316,N_20280);
and U22101 (N_22101,N_20366,N_20998);
xor U22102 (N_22102,N_20964,N_20957);
nand U22103 (N_22103,N_21151,N_21055);
or U22104 (N_22104,N_19719,N_20031);
xnor U22105 (N_22105,N_20800,N_21681);
or U22106 (N_22106,N_21410,N_19933);
and U22107 (N_22107,N_19759,N_19347);
nor U22108 (N_22108,N_19267,N_21286);
nand U22109 (N_22109,N_21441,N_19887);
nand U22110 (N_22110,N_19590,N_18750);
nor U22111 (N_22111,N_20218,N_20492);
xnor U22112 (N_22112,N_19960,N_21224);
nand U22113 (N_22113,N_20088,N_18773);
nor U22114 (N_22114,N_18849,N_20664);
and U22115 (N_22115,N_21709,N_18965);
nand U22116 (N_22116,N_19869,N_19349);
or U22117 (N_22117,N_20151,N_20315);
or U22118 (N_22118,N_20398,N_19332);
nor U22119 (N_22119,N_21345,N_19452);
and U22120 (N_22120,N_21445,N_20171);
or U22121 (N_22121,N_21409,N_19580);
nand U22122 (N_22122,N_19165,N_20812);
nand U22123 (N_22123,N_19926,N_19174);
nor U22124 (N_22124,N_20913,N_21557);
xnor U22125 (N_22125,N_19335,N_20540);
nand U22126 (N_22126,N_19682,N_20438);
or U22127 (N_22127,N_21838,N_20107);
nand U22128 (N_22128,N_20294,N_19297);
nand U22129 (N_22129,N_19560,N_18962);
xnor U22130 (N_22130,N_19709,N_19754);
or U22131 (N_22131,N_19011,N_19660);
nor U22132 (N_22132,N_19382,N_19197);
nor U22133 (N_22133,N_19099,N_21661);
and U22134 (N_22134,N_19793,N_19264);
nand U22135 (N_22135,N_19040,N_19813);
nor U22136 (N_22136,N_20187,N_20163);
or U22137 (N_22137,N_18861,N_19820);
or U22138 (N_22138,N_20385,N_21769);
and U22139 (N_22139,N_19270,N_20972);
nor U22140 (N_22140,N_20232,N_19477);
or U22141 (N_22141,N_18958,N_18886);
nand U22142 (N_22142,N_19268,N_20675);
or U22143 (N_22143,N_21746,N_19713);
and U22144 (N_22144,N_19224,N_21415);
nand U22145 (N_22145,N_20899,N_19834);
nor U22146 (N_22146,N_19078,N_21863);
nand U22147 (N_22147,N_19296,N_20886);
nand U22148 (N_22148,N_19086,N_21872);
nand U22149 (N_22149,N_20521,N_21288);
and U22150 (N_22150,N_19727,N_19739);
nand U22151 (N_22151,N_19030,N_19507);
and U22152 (N_22152,N_19354,N_21509);
xor U22153 (N_22153,N_19746,N_20119);
or U22154 (N_22154,N_20953,N_19232);
nand U22155 (N_22155,N_20146,N_18776);
nand U22156 (N_22156,N_21133,N_20468);
nand U22157 (N_22157,N_19254,N_19044);
and U22158 (N_22158,N_18866,N_18848);
or U22159 (N_22159,N_21324,N_18766);
or U22160 (N_22160,N_20966,N_21434);
nor U22161 (N_22161,N_19965,N_20445);
xor U22162 (N_22162,N_19430,N_20806);
and U22163 (N_22163,N_21397,N_19018);
or U22164 (N_22164,N_20444,N_20945);
and U22165 (N_22165,N_19629,N_21836);
or U22166 (N_22166,N_21483,N_20939);
nand U22167 (N_22167,N_19623,N_19652);
or U22168 (N_22168,N_21560,N_19095);
or U22169 (N_22169,N_20405,N_20080);
nor U22170 (N_22170,N_21077,N_21569);
nand U22171 (N_22171,N_21106,N_21644);
nand U22172 (N_22172,N_20795,N_20646);
nand U22173 (N_22173,N_18913,N_19515);
nor U22174 (N_22174,N_19495,N_20943);
nor U22175 (N_22175,N_20813,N_20298);
nor U22176 (N_22176,N_20547,N_19072);
and U22177 (N_22177,N_21865,N_18959);
xnor U22178 (N_22178,N_19522,N_21390);
and U22179 (N_22179,N_21125,N_21742);
xor U22180 (N_22180,N_21605,N_18927);
or U22181 (N_22181,N_19407,N_20853);
or U22182 (N_22182,N_19311,N_19523);
nor U22183 (N_22183,N_20035,N_19230);
and U22184 (N_22184,N_19890,N_19949);
xnor U22185 (N_22185,N_19667,N_20362);
or U22186 (N_22186,N_18875,N_21520);
xor U22187 (N_22187,N_21514,N_21270);
and U22188 (N_22188,N_19801,N_21039);
and U22189 (N_22189,N_20072,N_19298);
and U22190 (N_22190,N_19676,N_18756);
or U22191 (N_22191,N_21668,N_20157);
and U22192 (N_22192,N_19053,N_19484);
xor U22193 (N_22193,N_19046,N_20472);
nor U22194 (N_22194,N_20497,N_19130);
xnor U22195 (N_22195,N_18775,N_20680);
xnor U22196 (N_22196,N_19572,N_21518);
or U22197 (N_22197,N_21146,N_19140);
and U22198 (N_22198,N_19803,N_19392);
or U22199 (N_22199,N_19920,N_19519);
or U22200 (N_22200,N_20179,N_20710);
nand U22201 (N_22201,N_19081,N_19944);
nor U22202 (N_22202,N_19035,N_18936);
and U22203 (N_22203,N_19796,N_21240);
nand U22204 (N_22204,N_19742,N_21460);
and U22205 (N_22205,N_21305,N_20478);
nand U22206 (N_22206,N_19909,N_20951);
or U22207 (N_22207,N_18999,N_18857);
or U22208 (N_22208,N_21735,N_21767);
nor U22209 (N_22209,N_19073,N_21188);
and U22210 (N_22210,N_19026,N_20490);
nand U22211 (N_22211,N_21480,N_20217);
or U22212 (N_22212,N_20174,N_20463);
and U22213 (N_22213,N_18844,N_19108);
nor U22214 (N_22214,N_19415,N_20358);
nand U22215 (N_22215,N_20427,N_21021);
nor U22216 (N_22216,N_19677,N_21651);
or U22217 (N_22217,N_19181,N_20243);
nor U22218 (N_22218,N_20740,N_20282);
nor U22219 (N_22219,N_19322,N_18893);
and U22220 (N_22220,N_19568,N_18876);
xnor U22221 (N_22221,N_20573,N_21778);
or U22222 (N_22222,N_21579,N_18898);
nor U22223 (N_22223,N_21202,N_21869);
nand U22224 (N_22224,N_21671,N_20319);
nand U22225 (N_22225,N_20104,N_20344);
and U22226 (N_22226,N_19518,N_21163);
nand U22227 (N_22227,N_19163,N_20120);
nor U22228 (N_22228,N_21815,N_18797);
and U22229 (N_22229,N_20430,N_20918);
xor U22230 (N_22230,N_19594,N_20620);
nand U22231 (N_22231,N_19542,N_19546);
xor U22232 (N_22232,N_20852,N_19494);
or U22233 (N_22233,N_20220,N_19853);
or U22234 (N_22234,N_20407,N_21626);
or U22235 (N_22235,N_18878,N_21206);
or U22236 (N_22236,N_20757,N_21184);
nand U22237 (N_22237,N_20621,N_20326);
and U22238 (N_22238,N_19665,N_20630);
nor U22239 (N_22239,N_20567,N_18937);
or U22240 (N_22240,N_19233,N_20248);
and U22241 (N_22241,N_18784,N_20459);
and U22242 (N_22242,N_18977,N_19107);
nor U22243 (N_22243,N_19479,N_21331);
xnor U22244 (N_22244,N_19291,N_20068);
or U22245 (N_22245,N_19371,N_19336);
and U22246 (N_22246,N_21812,N_18836);
nand U22247 (N_22247,N_19562,N_20688);
or U22248 (N_22248,N_18889,N_20301);
nor U22249 (N_22249,N_19873,N_19902);
nand U22250 (N_22250,N_20961,N_20734);
or U22251 (N_22251,N_19122,N_18897);
xnor U22252 (N_22252,N_18765,N_21283);
nand U22253 (N_22253,N_21275,N_21094);
or U22254 (N_22254,N_19488,N_21692);
nor U22255 (N_22255,N_19816,N_19799);
nand U22256 (N_22256,N_20306,N_21547);
and U22257 (N_22257,N_19690,N_21851);
or U22258 (N_22258,N_21242,N_20867);
and U22259 (N_22259,N_21845,N_19000);
or U22260 (N_22260,N_19735,N_20101);
nor U22261 (N_22261,N_20968,N_21091);
or U22262 (N_22262,N_19948,N_21166);
or U22263 (N_22263,N_19171,N_20584);
or U22264 (N_22264,N_21057,N_20639);
or U22265 (N_22265,N_19006,N_21676);
and U22266 (N_22266,N_20075,N_21631);
and U22267 (N_22267,N_19992,N_20821);
and U22268 (N_22268,N_20199,N_21593);
nand U22269 (N_22269,N_20139,N_20507);
nor U22270 (N_22270,N_20586,N_20879);
nor U22271 (N_22271,N_21567,N_18955);
or U22272 (N_22272,N_19339,N_19090);
nor U22273 (N_22273,N_21190,N_21771);
and U22274 (N_22274,N_20695,N_20487);
nand U22275 (N_22275,N_21058,N_19941);
nor U22276 (N_22276,N_21842,N_20058);
nand U22277 (N_22277,N_19170,N_21515);
and U22278 (N_22278,N_20495,N_21723);
nor U22279 (N_22279,N_21293,N_21497);
and U22280 (N_22280,N_18782,N_19636);
and U22281 (N_22281,N_19931,N_21482);
or U22282 (N_22282,N_19289,N_20554);
and U22283 (N_22283,N_19583,N_21843);
nand U22284 (N_22284,N_19953,N_21236);
nand U22285 (N_22285,N_19865,N_20457);
nand U22286 (N_22286,N_21107,N_21622);
and U22287 (N_22287,N_20371,N_19603);
nand U22288 (N_22288,N_18824,N_20560);
nand U22289 (N_22289,N_21726,N_20588);
and U22290 (N_22290,N_20485,N_18903);
or U22291 (N_22291,N_18948,N_20699);
and U22292 (N_22292,N_20572,N_19967);
nand U22293 (N_22293,N_20352,N_19138);
nor U22294 (N_22294,N_20054,N_19505);
and U22295 (N_22295,N_19187,N_21718);
nor U22296 (N_22296,N_21674,N_21344);
or U22297 (N_22297,N_21447,N_21465);
and U22298 (N_22298,N_20030,N_21377);
nor U22299 (N_22299,N_19863,N_20707);
nor U22300 (N_22300,N_19555,N_19891);
nand U22301 (N_22301,N_21115,N_19679);
xnor U22302 (N_22302,N_21489,N_20532);
or U22303 (N_22303,N_19067,N_18909);
nand U22304 (N_22304,N_18935,N_19009);
xnor U22305 (N_22305,N_20153,N_19884);
nand U22306 (N_22306,N_20991,N_19693);
nand U22307 (N_22307,N_20359,N_18806);
and U22308 (N_22308,N_20623,N_19247);
nand U22309 (N_22309,N_21646,N_20917);
nor U22310 (N_22310,N_20980,N_20904);
nand U22311 (N_22311,N_19714,N_19786);
and U22312 (N_22312,N_21209,N_21401);
or U22313 (N_22313,N_20518,N_20406);
xnor U22314 (N_22314,N_19262,N_20106);
nor U22315 (N_22315,N_18879,N_21159);
nor U22316 (N_22316,N_19697,N_20216);
xor U22317 (N_22317,N_20860,N_19450);
nor U22318 (N_22318,N_19037,N_19925);
nor U22319 (N_22319,N_21523,N_20424);
and U22320 (N_22320,N_20862,N_20871);
xor U22321 (N_22321,N_19728,N_18894);
nor U22322 (N_22322,N_20150,N_19303);
nand U22323 (N_22323,N_20342,N_21462);
nor U22324 (N_22324,N_18973,N_21600);
nor U22325 (N_22325,N_19753,N_20911);
nand U22326 (N_22326,N_19432,N_19577);
or U22327 (N_22327,N_20287,N_20603);
nand U22328 (N_22328,N_20127,N_19628);
or U22329 (N_22329,N_20115,N_19722);
and U22330 (N_22330,N_20615,N_20797);
nand U22331 (N_22331,N_20439,N_19277);
nand U22332 (N_22332,N_21544,N_20159);
nor U22333 (N_22333,N_21788,N_21124);
nand U22334 (N_22334,N_21612,N_19841);
nor U22335 (N_22335,N_21635,N_21689);
or U22336 (N_22336,N_19769,N_19049);
or U22337 (N_22337,N_19467,N_19543);
or U22338 (N_22338,N_18795,N_21837);
or U22339 (N_22339,N_20923,N_21352);
nor U22340 (N_22340,N_18993,N_19278);
xor U22341 (N_22341,N_19864,N_20903);
and U22342 (N_22342,N_18858,N_20251);
and U22343 (N_22343,N_19050,N_19932);
or U22344 (N_22344,N_20817,N_19913);
and U22345 (N_22345,N_21485,N_21476);
nand U22346 (N_22346,N_19261,N_19103);
and U22347 (N_22347,N_19550,N_19146);
nand U22348 (N_22348,N_18901,N_18814);
nand U22349 (N_22349,N_21100,N_19117);
or U22350 (N_22350,N_20017,N_20536);
and U22351 (N_22351,N_18829,N_18980);
or U22352 (N_22352,N_19898,N_18786);
nand U22353 (N_22353,N_20376,N_20268);
and U22354 (N_22354,N_21857,N_21634);
nor U22355 (N_22355,N_21068,N_20741);
or U22356 (N_22356,N_21357,N_19314);
nand U22357 (N_22357,N_19566,N_21627);
nor U22358 (N_22358,N_19194,N_18768);
nor U22359 (N_22359,N_21155,N_21858);
nor U22360 (N_22360,N_20196,N_21502);
and U22361 (N_22361,N_21274,N_19259);
and U22362 (N_22362,N_21154,N_19996);
nand U22363 (N_22363,N_21525,N_20435);
or U22364 (N_22364,N_21255,N_20004);
nor U22365 (N_22365,N_19549,N_21454);
nand U22366 (N_22366,N_21307,N_20905);
or U22367 (N_22367,N_20098,N_18819);
and U22368 (N_22368,N_19048,N_19413);
or U22369 (N_22369,N_18969,N_19329);
nand U22370 (N_22370,N_20876,N_21790);
nand U22371 (N_22371,N_19075,N_19089);
nor U22372 (N_22372,N_21027,N_19051);
nand U22373 (N_22373,N_21061,N_20133);
nand U22374 (N_22374,N_20823,N_19648);
and U22375 (N_22375,N_21253,N_19193);
xnor U22376 (N_22376,N_21664,N_20078);
nor U22377 (N_22377,N_19743,N_20310);
and U22378 (N_22378,N_21004,N_19758);
and U22379 (N_22379,N_19708,N_21487);
nand U22380 (N_22380,N_20722,N_19326);
nand U22381 (N_22381,N_19975,N_19508);
nand U22382 (N_22382,N_20001,N_20838);
and U22383 (N_22383,N_21412,N_19290);
nand U22384 (N_22384,N_19692,N_19379);
and U22385 (N_22385,N_21542,N_20895);
and U22386 (N_22386,N_21507,N_20869);
or U22387 (N_22387,N_19706,N_20973);
nand U22388 (N_22388,N_21290,N_19721);
xor U22389 (N_22389,N_18933,N_21458);
or U22390 (N_22390,N_19002,N_18957);
xnor U22391 (N_22391,N_20308,N_20984);
nand U22392 (N_22392,N_20191,N_20081);
nand U22393 (N_22393,N_21564,N_21583);
nor U22394 (N_22394,N_19131,N_21696);
and U22395 (N_22395,N_19608,N_21733);
nor U22396 (N_22396,N_19837,N_21132);
nand U22397 (N_22397,N_21652,N_20786);
or U22398 (N_22398,N_21789,N_19586);
nor U22399 (N_22399,N_19601,N_19375);
nand U22400 (N_22400,N_19497,N_21695);
nor U22401 (N_22401,N_21504,N_21313);
nor U22402 (N_22402,N_20896,N_20130);
or U22403 (N_22403,N_21291,N_21519);
nor U22404 (N_22404,N_20826,N_20135);
or U22405 (N_22405,N_18859,N_18982);
nand U22406 (N_22406,N_20643,N_19642);
or U22407 (N_22407,N_18952,N_21591);
nand U22408 (N_22408,N_18764,N_21496);
and U22409 (N_22409,N_18981,N_20527);
or U22410 (N_22410,N_19167,N_21640);
and U22411 (N_22411,N_21203,N_21081);
and U22412 (N_22412,N_20732,N_20458);
nand U22413 (N_22413,N_18890,N_21639);
nor U22414 (N_22414,N_21551,N_21131);
or U22415 (N_22415,N_19079,N_19439);
nand U22416 (N_22416,N_21570,N_20802);
and U22417 (N_22417,N_20210,N_19183);
nor U22418 (N_22418,N_21380,N_18774);
nand U22419 (N_22419,N_20986,N_20307);
nand U22420 (N_22420,N_21079,N_21474);
nor U22421 (N_22421,N_19499,N_19025);
nand U22422 (N_22422,N_20541,N_18900);
or U22423 (N_22423,N_20624,N_21031);
or U22424 (N_22424,N_21594,N_18932);
nor U22425 (N_22425,N_20790,N_19065);
and U22426 (N_22426,N_20390,N_20552);
or U22427 (N_22427,N_19124,N_21715);
nand U22428 (N_22428,N_21556,N_20419);
and U22429 (N_22429,N_19880,N_20701);
nor U22430 (N_22430,N_19350,N_20716);
nand U22431 (N_22431,N_18793,N_19658);
or U22432 (N_22432,N_21208,N_21161);
nand U22433 (N_22433,N_20657,N_19087);
nor U22434 (N_22434,N_21432,N_19214);
xor U22435 (N_22435,N_21472,N_21366);
or U22436 (N_22436,N_19490,N_19128);
nor U22437 (N_22437,N_21017,N_19663);
or U22438 (N_22438,N_20520,N_21322);
and U22439 (N_22439,N_19272,N_21540);
or U22440 (N_22440,N_21470,N_21731);
xor U22441 (N_22441,N_20955,N_19386);
or U22442 (N_22442,N_19678,N_19414);
or U22443 (N_22443,N_21076,N_20866);
nand U22444 (N_22444,N_21334,N_20835);
or U22445 (N_22445,N_20967,N_18771);
nand U22446 (N_22446,N_21765,N_21793);
or U22447 (N_22447,N_21393,N_19180);
or U22448 (N_22448,N_20663,N_18961);
and U22449 (N_22449,N_19511,N_19191);
or U22450 (N_22450,N_20348,N_20910);
or U22451 (N_22451,N_19689,N_20799);
and U22452 (N_22452,N_21453,N_20929);
xnor U22453 (N_22453,N_19400,N_19200);
or U22454 (N_22454,N_20595,N_19937);
nand U22455 (N_22455,N_21478,N_20997);
nor U22456 (N_22456,N_21269,N_21568);
xnor U22457 (N_22457,N_18868,N_21656);
nor U22458 (N_22458,N_21750,N_21529);
nand U22459 (N_22459,N_21448,N_19936);
nor U22460 (N_22460,N_21770,N_19892);
or U22461 (N_22461,N_20960,N_18854);
nand U22462 (N_22462,N_21728,N_21374);
or U22463 (N_22463,N_21552,N_20726);
nand U22464 (N_22464,N_21000,N_19016);
and U22465 (N_22465,N_21003,N_19469);
xnor U22466 (N_22466,N_19997,N_21451);
xnor U22467 (N_22467,N_19579,N_21247);
xor U22468 (N_22468,N_19985,N_19524);
nor U22469 (N_22469,N_21721,N_20909);
and U22470 (N_22470,N_21030,N_20043);
or U22471 (N_22471,N_20831,N_20975);
xor U22472 (N_22472,N_19866,N_19872);
or U22473 (N_22473,N_19255,N_19184);
nor U22474 (N_22474,N_21308,N_20890);
and U22475 (N_22475,N_20143,N_20073);
nor U22476 (N_22476,N_21625,N_19847);
or U22477 (N_22477,N_19116,N_20227);
nand U22478 (N_22478,N_20394,N_20999);
or U22479 (N_22479,N_20613,N_20194);
nand U22480 (N_22480,N_19039,N_19235);
and U22481 (N_22481,N_21748,N_19504);
and U22482 (N_22482,N_20221,N_20203);
nand U22483 (N_22483,N_20047,N_19227);
nand U22484 (N_22484,N_20005,N_21102);
nor U22485 (N_22485,N_19166,N_19609);
or U22486 (N_22486,N_19119,N_18816);
nor U22487 (N_22487,N_21510,N_21085);
nor U22488 (N_22488,N_21332,N_19620);
and U22489 (N_22489,N_20944,N_20368);
nor U22490 (N_22490,N_20166,N_19070);
and U22491 (N_22491,N_21020,N_18953);
nor U22492 (N_22492,N_21704,N_19190);
or U22493 (N_22493,N_21650,N_18853);
nand U22494 (N_22494,N_20829,N_18852);
nand U22495 (N_22495,N_19251,N_20897);
nand U22496 (N_22496,N_19616,N_20545);
and U22497 (N_22497,N_19092,N_19973);
or U22498 (N_22498,N_20340,N_21655);
nor U22499 (N_22499,N_21272,N_19805);
and U22500 (N_22500,N_18991,N_21846);
nor U22501 (N_22501,N_19541,N_20042);
nand U22502 (N_22502,N_21212,N_19109);
nor U22503 (N_22503,N_20295,N_20851);
and U22504 (N_22504,N_21713,N_21550);
or U22505 (N_22505,N_20856,N_19638);
nor U22506 (N_22506,N_21343,N_20598);
xor U22507 (N_22507,N_19442,N_20600);
nand U22508 (N_22508,N_19388,N_19653);
nor U22509 (N_22509,N_20610,N_19317);
xor U22510 (N_22510,N_19526,N_21364);
nor U22511 (N_22511,N_20668,N_21802);
and U22512 (N_22512,N_19279,N_21484);
nand U22513 (N_22513,N_19383,N_19323);
nor U22514 (N_22514,N_19797,N_20372);
nand U22515 (N_22515,N_19701,N_20828);
or U22516 (N_22516,N_21792,N_20184);
nand U22517 (N_22517,N_19088,N_19705);
nor U22518 (N_22518,N_19397,N_21740);
xnor U22519 (N_22519,N_20048,N_21150);
xor U22520 (N_22520,N_19403,N_20128);
nand U22521 (N_22521,N_20314,N_19308);
nor U22522 (N_22522,N_20136,N_18924);
xnor U22523 (N_22523,N_19360,N_21545);
and U22524 (N_22524,N_19113,N_20175);
xnor U22525 (N_22525,N_21222,N_21589);
and U22526 (N_22526,N_19563,N_19273);
or U22527 (N_22527,N_21136,N_19024);
xnor U22528 (N_22528,N_21614,N_21645);
nand U22529 (N_22529,N_18788,N_21090);
nand U22530 (N_22530,N_20916,N_21177);
nand U22531 (N_22531,N_20570,N_19346);
nand U22532 (N_22532,N_20291,N_18772);
nor U22533 (N_22533,N_19780,N_21586);
or U22534 (N_22534,N_20962,N_20097);
nor U22535 (N_22535,N_20456,N_19410);
nor U22536 (N_22536,N_19951,N_20483);
xor U22537 (N_22537,N_19731,N_19201);
xnor U22538 (N_22538,N_20237,N_21641);
nand U22539 (N_22539,N_18994,N_19900);
or U22540 (N_22540,N_21424,N_21747);
nand U22541 (N_22541,N_21311,N_19256);
nand U22542 (N_22542,N_21251,N_19792);
and U22543 (N_22543,N_20870,N_20297);
nand U22544 (N_22544,N_20055,N_19894);
nor U22545 (N_22545,N_18851,N_19123);
and U22546 (N_22546,N_21444,N_19699);
nand U22547 (N_22547,N_20958,N_20609);
or U22548 (N_22548,N_19390,N_19475);
xor U22549 (N_22549,N_21259,N_19644);
and U22550 (N_22550,N_19972,N_19457);
nor U22551 (N_22551,N_21381,N_19137);
and U22552 (N_22552,N_20225,N_20733);
nor U22553 (N_22553,N_21403,N_19928);
nand U22554 (N_22554,N_20486,N_21682);
or U22555 (N_22555,N_21120,N_20915);
and U22556 (N_22556,N_19305,N_20760);
and U22557 (N_22557,N_20571,N_21037);
and U22558 (N_22558,N_18987,N_19010);
nand U22559 (N_22559,N_19655,N_18821);
nand U22560 (N_22560,N_21104,N_20488);
or U22561 (N_22561,N_18787,N_19671);
and U22562 (N_22562,N_21811,N_19443);
xor U22563 (N_22563,N_19899,N_20705);
nand U22564 (N_22564,N_19647,N_20256);
or U22565 (N_22565,N_21420,N_19441);
nor U22566 (N_22566,N_19310,N_21093);
nor U22567 (N_22567,N_19159,N_19287);
xor U22568 (N_22568,N_20614,N_20420);
nor U22569 (N_22569,N_20476,N_19096);
or U22570 (N_22570,N_20040,N_21219);
xor U22571 (N_22571,N_21162,N_18767);
or U22572 (N_22572,N_20683,N_20281);
and U22573 (N_22573,N_19923,N_21642);
or U22574 (N_22574,N_21808,N_20775);
xor U22575 (N_22575,N_19176,N_21761);
nor U22576 (N_22576,N_19416,N_21365);
and U22577 (N_22577,N_19066,N_19650);
xnor U22578 (N_22578,N_19857,N_20470);
nand U22579 (N_22579,N_20448,N_20810);
nand U22580 (N_22580,N_20881,N_21144);
nand U22581 (N_22581,N_19833,N_21379);
or U22582 (N_22582,N_20787,N_19589);
and U22583 (N_22583,N_19552,N_20739);
or U22584 (N_22584,N_19987,N_21359);
xnor U22585 (N_22585,N_19344,N_20138);
or U22586 (N_22586,N_19148,N_19883);
nor U22587 (N_22587,N_19718,N_20956);
or U22588 (N_22588,N_20887,N_19424);
nand U22589 (N_22589,N_19882,N_21176);
xnor U22590 (N_22590,N_21328,N_20212);
and U22591 (N_22591,N_20672,N_19082);
and U22592 (N_22592,N_21349,N_20498);
nand U22593 (N_22593,N_21853,N_19971);
nand U22594 (N_22594,N_19668,N_20526);
and U22595 (N_22595,N_21063,N_20322);
nor U22596 (N_22596,N_21571,N_19271);
nand U22597 (N_22597,N_19859,N_20667);
or U22598 (N_22598,N_19266,N_19532);
and U22599 (N_22599,N_19656,N_19288);
xnor U22600 (N_22600,N_19807,N_20018);
nor U22601 (N_22601,N_19406,N_18803);
or U22602 (N_22602,N_19763,N_21369);
or U22603 (N_22603,N_21597,N_18871);
nor U22604 (N_22604,N_21407,N_19540);
nor U22605 (N_22605,N_21455,N_21034);
xor U22606 (N_22606,N_19950,N_19063);
nor U22607 (N_22607,N_18808,N_20046);
xor U22608 (N_22608,N_21543,N_20583);
nor U22609 (N_22609,N_19212,N_20948);
and U22610 (N_22610,N_21436,N_19356);
or U22611 (N_22611,N_20279,N_19207);
or U22612 (N_22612,N_19772,N_21665);
or U22613 (N_22613,N_19637,N_19470);
or U22614 (N_22614,N_18950,N_21258);
and U22615 (N_22615,N_20985,N_19666);
and U22616 (N_22616,N_20387,N_21630);
and U22617 (N_22617,N_18789,N_19164);
and U22618 (N_22618,N_19372,N_19150);
or U22619 (N_22619,N_20748,N_19438);
and U22620 (N_22620,N_20354,N_20743);
or U22621 (N_22621,N_20924,N_19968);
nand U22622 (N_22622,N_21762,N_20264);
and U22623 (N_22623,N_20079,N_19151);
xor U22624 (N_22624,N_21446,N_19582);
and U22625 (N_22625,N_19812,N_19173);
or U22626 (N_22626,N_19831,N_19395);
or U22627 (N_22627,N_21248,N_21416);
nor U22628 (N_22628,N_19617,N_20605);
and U22629 (N_22629,N_19280,N_21422);
or U22630 (N_22630,N_20403,N_19045);
and U22631 (N_22631,N_21637,N_21755);
xor U22632 (N_22632,N_20258,N_18990);
nor U22633 (N_22633,N_21355,N_19043);
nand U22634 (N_22634,N_21654,N_21033);
xnor U22635 (N_22635,N_21503,N_20704);
or U22636 (N_22636,N_21559,N_20693);
nand U22637 (N_22637,N_19558,N_19654);
and U22638 (N_22638,N_21814,N_21830);
and U22639 (N_22639,N_20591,N_19964);
xnor U22640 (N_22640,N_20230,N_21500);
nor U22641 (N_22641,N_18845,N_21372);
nand U22642 (N_22642,N_18818,N_18880);
nor U22643 (N_22643,N_19893,N_21850);
nand U22644 (N_22644,N_20604,N_18882);
and U22645 (N_22645,N_19745,N_19659);
and U22646 (N_22646,N_20197,N_18779);
nand U22647 (N_22647,N_20316,N_21169);
nor U22648 (N_22648,N_21373,N_20883);
and U22649 (N_22649,N_19058,N_21777);
or U22650 (N_22650,N_19085,N_20023);
or U22651 (N_22651,N_20912,N_18966);
or U22652 (N_22652,N_19185,N_20627);
or U22653 (N_22653,N_19662,N_18825);
nor U22654 (N_22654,N_20284,N_19094);
and U22655 (N_22655,N_19911,N_19394);
nor U22656 (N_22656,N_20530,N_20063);
nand U22657 (N_22657,N_20954,N_20825);
or U22658 (N_22658,N_19955,N_20399);
or U22659 (N_22659,N_20379,N_19057);
nor U22660 (N_22660,N_21193,N_20027);
nand U22661 (N_22661,N_19449,N_21172);
nor U22662 (N_22662,N_21336,N_21235);
nand U22663 (N_22663,N_21683,N_19795);
and U22664 (N_22664,N_21032,N_19237);
nor U22665 (N_22665,N_19369,N_21471);
xor U22666 (N_22666,N_20789,N_21325);
nor U22667 (N_22667,N_19588,N_20762);
or U22668 (N_22668,N_21794,N_19215);
and U22669 (N_22669,N_21672,N_20434);
nor U22670 (N_22670,N_20516,N_20780);
or U22671 (N_22671,N_19418,N_21697);
nand U22672 (N_22672,N_20325,N_19352);
and U22673 (N_22673,N_19343,N_19600);
xnor U22674 (N_22674,N_20026,N_21706);
nand U22675 (N_22675,N_20581,N_20231);
or U22676 (N_22676,N_20854,N_20186);
or U22677 (N_22677,N_19849,N_19355);
or U22678 (N_22678,N_21859,N_19454);
or U22679 (N_22679,N_20848,N_21826);
nor U22680 (N_22680,N_20859,N_19189);
nor U22681 (N_22681,N_20234,N_21179);
nor U22682 (N_22682,N_20706,N_20612);
and U22683 (N_22683,N_21388,N_19528);
or U22684 (N_22684,N_19602,N_21528);
nor U22685 (N_22685,N_19301,N_20192);
or U22686 (N_22686,N_20123,N_18906);
nor U22687 (N_22687,N_19320,N_20501);
nor U22688 (N_22688,N_20449,N_21592);
nand U22689 (N_22689,N_20057,N_19423);
nor U22690 (N_22690,N_19313,N_21066);
nand U22691 (N_22691,N_20009,N_21347);
and U22692 (N_22692,N_20069,N_19132);
xor U22693 (N_22693,N_19425,N_21295);
xnor U22694 (N_22694,N_21720,N_19008);
and U22695 (N_22695,N_21862,N_21145);
or U22696 (N_22696,N_21861,N_21693);
and U22697 (N_22697,N_19788,N_21584);
and U22698 (N_22698,N_21348,N_19592);
nand U22699 (N_22699,N_19396,N_18949);
nand U22700 (N_22700,N_21475,N_19633);
and U22701 (N_22701,N_20155,N_18997);
and U22702 (N_22702,N_18911,N_21511);
xor U22703 (N_22703,N_19007,N_19958);
and U22704 (N_22704,N_20033,N_21268);
or U22705 (N_22705,N_20730,N_19389);
and U22706 (N_22706,N_21582,N_21147);
and U22707 (N_22707,N_18884,N_21012);
nor U22708 (N_22708,N_20655,N_20410);
and U22709 (N_22709,N_21439,N_20576);
nand U22710 (N_22710,N_19312,N_19736);
or U22711 (N_22711,N_19120,N_20028);
nand U22712 (N_22712,N_20843,N_21217);
nand U22713 (N_22713,N_21526,N_18995);
xnor U22714 (N_22714,N_20401,N_21825);
and U22715 (N_22715,N_20963,N_20577);
xnor U22716 (N_22716,N_19704,N_18834);
nor U22717 (N_22717,N_19798,N_19979);
nor U22718 (N_22718,N_19771,N_19331);
or U22719 (N_22719,N_21666,N_21466);
or U22720 (N_22720,N_21111,N_18891);
nand U22721 (N_22721,N_21007,N_21049);
nand U22722 (N_22722,N_21156,N_20849);
and U22723 (N_22723,N_20246,N_20767);
and U22724 (N_22724,N_21186,N_20094);
nor U22725 (N_22725,N_20546,N_19741);
nor U22726 (N_22726,N_19340,N_20763);
or U22727 (N_22727,N_20323,N_21754);
nand U22728 (N_22728,N_18989,N_19250);
or U22729 (N_22729,N_19990,N_20788);
and U22730 (N_22730,N_18976,N_20059);
nor U22731 (N_22731,N_21127,N_20003);
and U22732 (N_22732,N_21074,N_18810);
and U22733 (N_22733,N_19604,N_20053);
nor U22734 (N_22734,N_19502,N_20592);
nor U22735 (N_22735,N_19474,N_21375);
nor U22736 (N_22736,N_19624,N_20402);
and U22737 (N_22737,N_21371,N_18839);
nor U22738 (N_22738,N_21618,N_19104);
xor U22739 (N_22739,N_18963,N_21048);
nand U22740 (N_22740,N_21522,N_20622);
or U22741 (N_22741,N_21244,N_21009);
and U22742 (N_22742,N_20351,N_20167);
nor U22743 (N_22743,N_19606,N_18781);
nor U22744 (N_22744,N_18811,N_19755);
nand U22745 (N_22745,N_20178,N_20111);
nor U22746 (N_22746,N_21534,N_20118);
or U22747 (N_22747,N_19222,N_21233);
or U22748 (N_22748,N_20770,N_21223);
nand U22749 (N_22749,N_18863,N_19020);
xnor U22750 (N_22750,N_20395,N_21276);
nand U22751 (N_22751,N_21760,N_19364);
and U22752 (N_22752,N_19012,N_21304);
or U22753 (N_22753,N_21578,N_21421);
xnor U22754 (N_22754,N_20772,N_21677);
nand U22755 (N_22755,N_21092,N_21110);
nor U22756 (N_22756,N_20378,N_19994);
xnor U22757 (N_22757,N_20919,N_21404);
nor U22758 (N_22758,N_20408,N_20116);
or U22759 (N_22759,N_21759,N_20036);
nor U22760 (N_22760,N_19292,N_19129);
and U22761 (N_22761,N_20303,N_20393);
nand U22762 (N_22762,N_20908,N_19732);
xnor U22763 (N_22763,N_20606,N_20383);
nor U22764 (N_22764,N_18988,N_19553);
nor U22765 (N_22765,N_21370,N_20714);
or U22766 (N_22766,N_21662,N_20204);
nor U22767 (N_22767,N_21435,N_18867);
xor U22768 (N_22768,N_21165,N_20103);
or U22769 (N_22769,N_21153,N_19198);
nand U22770 (N_22770,N_18799,N_20661);
and U22771 (N_22771,N_19071,N_19943);
and U22772 (N_22772,N_20207,N_19341);
nor U22773 (N_22773,N_21546,N_21001);
nand U22774 (N_22774,N_19875,N_19711);
or U22775 (N_22775,N_19399,N_19260);
and U22776 (N_22776,N_20529,N_20266);
xnor U22777 (N_22777,N_18752,N_20696);
xnor U22778 (N_22778,N_20145,N_20659);
xnor U22779 (N_22779,N_21383,N_20666);
xnor U22780 (N_22780,N_20801,N_19223);
or U22781 (N_22781,N_20992,N_21191);
nand U22782 (N_22782,N_18792,N_20798);
nand U22783 (N_22783,N_21297,N_21130);
nor U22784 (N_22784,N_20601,N_21340);
and U22785 (N_22785,N_21737,N_20555);
nor U22786 (N_22786,N_18925,N_20839);
or U22787 (N_22787,N_20937,N_19716);
nand U22788 (N_22788,N_20313,N_19986);
or U22789 (N_22789,N_19217,N_20052);
and U22790 (N_22790,N_21226,N_20124);
and U22791 (N_22791,N_20233,N_19461);
nand U22792 (N_22792,N_21548,N_20353);
or U22793 (N_22793,N_19995,N_21675);
xor U22794 (N_22794,N_20441,N_18833);
and U22795 (N_22795,N_19782,N_21833);
nor U22796 (N_22796,N_20160,N_20267);
or U22797 (N_22797,N_20329,N_19781);
and U22798 (N_22798,N_21006,N_19750);
and U22799 (N_22799,N_19409,N_20785);
nand U22800 (N_22800,N_19139,N_18983);
nand U22801 (N_22801,N_18755,N_21494);
and U22802 (N_22802,N_19042,N_19752);
and U22803 (N_22803,N_19570,N_19618);
nor U22804 (N_22804,N_19919,N_20750);
nand U22805 (N_22805,N_18992,N_19133);
nor U22806 (N_22806,N_21596,N_20921);
nand U22807 (N_22807,N_18922,N_20561);
nor U22808 (N_22808,N_19022,N_20421);
and U22809 (N_22809,N_21623,N_21067);
nor U22810 (N_22810,N_19557,N_21231);
and U22811 (N_22811,N_21109,N_21699);
and U22812 (N_22812,N_21601,N_20249);
nand U22813 (N_22813,N_19236,N_20803);
nand U22814 (N_22814,N_19556,N_20050);
and U22815 (N_22815,N_21214,N_19054);
nand U22816 (N_22816,N_21820,N_21440);
nor U22817 (N_22817,N_19734,N_19286);
or U22818 (N_22818,N_19897,N_21225);
nor U22819 (N_22819,N_20926,N_19001);
or U22820 (N_22820,N_20989,N_21459);
and U22821 (N_22821,N_20637,N_19208);
nand U22822 (N_22822,N_19768,N_21516);
and U22823 (N_22823,N_19307,N_21512);
nand U22824 (N_22824,N_20563,N_19225);
nor U22825 (N_22825,N_21585,N_18945);
or U22826 (N_22826,N_19209,N_20041);
nand U22827 (N_22827,N_20818,N_21744);
xor U22828 (N_22828,N_19378,N_19363);
and U22829 (N_22829,N_19381,N_21185);
or U22830 (N_22830,N_20317,N_19465);
nand U22831 (N_22831,N_20265,N_20242);
nand U22832 (N_22832,N_19981,N_18943);
nor U22833 (N_22833,N_19896,N_20428);
and U22834 (N_22834,N_21554,N_18869);
xor U22835 (N_22835,N_18780,N_18912);
nand U22836 (N_22836,N_20369,N_20528);
and U22837 (N_22837,N_20755,N_18986);
xnor U22838 (N_22838,N_20723,N_21129);
and U22839 (N_22839,N_19330,N_21088);
nand U22840 (N_22840,N_19605,N_21595);
nor U22841 (N_22841,N_19411,N_20671);
nand U22842 (N_22842,N_21563,N_19702);
nor U22843 (N_22843,N_20971,N_19324);
nor U22844 (N_22844,N_19530,N_21042);
nand U22845 (N_22845,N_20152,N_19436);
or U22846 (N_22846,N_19538,N_21739);
or U22847 (N_22847,N_20377,N_21149);
and U22848 (N_22848,N_19977,N_19244);
nand U22849 (N_22849,N_19861,N_19724);
or U22850 (N_22850,N_19402,N_19800);
and U22851 (N_22851,N_21292,N_19161);
and U22852 (N_22852,N_20616,N_19626);
xor U22853 (N_22853,N_20259,N_20935);
and U22854 (N_22854,N_21856,N_20275);
and U22855 (N_22855,N_21189,N_19569);
and U22856 (N_22856,N_21611,N_21289);
and U22857 (N_22857,N_20952,N_19551);
nor U22858 (N_22858,N_20484,N_20147);
nor U22859 (N_22859,N_20429,N_21216);
nand U22860 (N_22860,N_19169,N_18778);
nand U22861 (N_22861,N_20482,N_20777);
nand U22862 (N_22862,N_21686,N_20121);
nor U22863 (N_22863,N_19431,N_20007);
nor U22864 (N_22864,N_19135,N_21824);
or U22865 (N_22865,N_19525,N_19429);
and U22866 (N_22866,N_20865,N_20650);
xnor U22867 (N_22867,N_21069,N_19076);
nor U22868 (N_22868,N_20183,N_19342);
nand U22869 (N_22869,N_20841,N_21687);
or U22870 (N_22870,N_20891,N_20397);
or U22871 (N_22871,N_21473,N_20662);
and U22872 (N_22872,N_19680,N_20746);
and U22873 (N_22873,N_19240,N_19033);
nand U22874 (N_22874,N_19019,N_20473);
and U22875 (N_22875,N_19695,N_20363);
or U22876 (N_22876,N_20508,N_21354);
and U22877 (N_22877,N_21060,N_21378);
or U22878 (N_22878,N_20582,N_19930);
or U22879 (N_22879,N_19204,N_19641);
or U22880 (N_22880,N_20889,N_18923);
and U22881 (N_22881,N_20062,N_20736);
nand U22882 (N_22882,N_19265,N_21072);
or U22883 (N_22883,N_18946,N_21362);
and U22884 (N_22884,N_20974,N_19574);
and U22885 (N_22885,N_18842,N_20708);
nand U22886 (N_22886,N_20411,N_18802);
nor U22887 (N_22887,N_20404,N_19961);
and U22888 (N_22888,N_19684,N_19761);
nor U22889 (N_22889,N_21041,N_21078);
xnor U22890 (N_22890,N_19717,N_19827);
nor U22891 (N_22891,N_21531,N_20778);
or U22892 (N_22892,N_20677,N_19527);
or U22893 (N_22893,N_19729,N_20361);
and U22894 (N_22894,N_21019,N_21196);
nor U22895 (N_22895,N_19575,N_21690);
or U22896 (N_22896,N_20684,N_19068);
xor U22897 (N_22897,N_19683,N_20188);
nor U22898 (N_22898,N_19206,N_19179);
and U22899 (N_22899,N_19458,N_20846);
nand U22900 (N_22900,N_20158,N_20244);
and U22901 (N_22901,N_19565,N_19083);
and U22902 (N_22902,N_20827,N_20796);
nor U22903 (N_22903,N_20205,N_20872);
and U22904 (N_22904,N_21598,N_21164);
and U22905 (N_22905,N_20644,N_21873);
xnor U22906 (N_22906,N_19694,N_19988);
or U22907 (N_22907,N_20894,N_20641);
nand U22908 (N_22908,N_18762,N_18823);
nand U22909 (N_22909,N_21866,N_21708);
and U22910 (N_22910,N_21018,N_21558);
nor U22911 (N_22911,N_18919,N_20766);
nor U22912 (N_22912,N_19970,N_20338);
or U22913 (N_22913,N_18947,N_21527);
or U22914 (N_22914,N_21620,N_19257);
nand U22915 (N_22915,N_20773,N_19032);
xor U22916 (N_22916,N_19168,N_19991);
nor U22917 (N_22917,N_19843,N_21684);
xor U22918 (N_22918,N_19412,N_19536);
or U22919 (N_22919,N_20898,N_20932);
xnor U22920 (N_22920,N_19238,N_21029);
or U22921 (N_22921,N_20618,N_21711);
nor U22922 (N_22922,N_20976,N_20360);
xnor U22923 (N_22923,N_20481,N_20725);
and U22924 (N_22924,N_21729,N_20654);
xnor U22925 (N_22925,N_20022,N_20320);
xnor U22926 (N_22926,N_18873,N_21572);
xnor U22927 (N_22927,N_19669,N_20686);
nand U22928 (N_22928,N_19802,N_19593);
xor U22929 (N_22929,N_20496,N_20446);
xor U22930 (N_22930,N_21112,N_21181);
nor U22931 (N_22931,N_19318,N_20709);
or U22932 (N_22932,N_19069,N_21670);
nand U22933 (N_22933,N_20631,N_18895);
or U22934 (N_22934,N_19093,N_21234);
or U22935 (N_22935,N_20083,N_18800);
nor U22936 (N_22936,N_21408,N_19234);
nor U22937 (N_22937,N_21167,N_20113);
xnor U22938 (N_22938,N_20093,N_19632);
nand U22939 (N_22939,N_20629,N_20334);
or U22940 (N_22940,N_19815,N_20805);
nor U22941 (N_22941,N_19646,N_21469);
nand U22942 (N_22942,N_20596,N_21321);
and U22943 (N_22943,N_21624,N_18758);
or U22944 (N_22944,N_20089,N_21013);
or U22945 (N_22945,N_20260,N_20453);
nor U22946 (N_22946,N_19052,N_21752);
xor U22947 (N_22947,N_21629,N_19635);
nand U22948 (N_22948,N_21036,N_20717);
or U22949 (N_22949,N_20522,N_20431);
nand U22950 (N_22950,N_19611,N_18899);
and U22951 (N_22951,N_21122,N_21194);
or U22952 (N_22952,N_18809,N_21395);
or U22953 (N_22953,N_19489,N_21358);
xnor U22954 (N_22954,N_19839,N_19916);
xor U22955 (N_22955,N_19999,N_19463);
nand U22956 (N_22956,N_20426,N_19060);
nor U22957 (N_22957,N_20350,N_21803);
nor U22958 (N_22958,N_20416,N_21160);
nand U22959 (N_22959,N_20110,N_21505);
nor U22960 (N_22960,N_21227,N_21285);
nor U22961 (N_22961,N_21602,N_20602);
nor U22962 (N_22962,N_21486,N_21479);
or U22963 (N_22963,N_18769,N_21221);
nand U22964 (N_22964,N_18883,N_19098);
nand U22965 (N_22965,N_21073,N_20271);
nand U22966 (N_22966,N_19385,N_19034);
and U22967 (N_22967,N_19195,N_20274);
nand U22968 (N_22968,N_19573,N_21712);
nor U22969 (N_22969,N_21852,N_19293);
nand U22970 (N_22970,N_19814,N_20959);
or U22971 (N_22971,N_19976,N_19698);
nor U22972 (N_22972,N_20804,N_20465);
nor U22973 (N_22973,N_21252,N_21016);
nor U22974 (N_22974,N_19152,N_20201);
nor U22975 (N_22975,N_19249,N_19760);
or U22976 (N_22976,N_21786,N_21095);
nand U22977 (N_22977,N_19959,N_21087);
and U22978 (N_22978,N_20357,N_20182);
and U22979 (N_22979,N_21329,N_20335);
and U22980 (N_22980,N_19517,N_21101);
nand U22981 (N_22981,N_20240,N_21298);
or U22982 (N_22982,N_19365,N_21023);
xnor U22983 (N_22983,N_19091,N_21603);
nor U22984 (N_22984,N_21673,N_19707);
nor U22985 (N_22985,N_21306,N_20273);
and U22986 (N_22986,N_21710,N_20517);
or U22987 (N_22987,N_21782,N_20011);
nor U22988 (N_22988,N_21658,N_19747);
nand U22989 (N_22989,N_21530,N_20169);
nand U22990 (N_22990,N_19226,N_20002);
nor U22991 (N_22991,N_18754,N_21613);
nand U22992 (N_22992,N_19929,N_19830);
nor U22993 (N_22993,N_18998,N_19826);
xnor U22994 (N_22994,N_19888,N_21743);
nand U22995 (N_22995,N_19061,N_20288);
nand U22996 (N_22996,N_21784,N_20471);
xor U22997 (N_22997,N_20021,N_19625);
or U22998 (N_22998,N_19686,N_19775);
nor U22999 (N_22999,N_19205,N_20494);
and U23000 (N_23000,N_19766,N_18934);
nand U23001 (N_23001,N_20981,N_21071);
and U23002 (N_23002,N_18862,N_21638);
and U23003 (N_23003,N_18892,N_20100);
and U23004 (N_23004,N_21368,N_19263);
and U23005 (N_23005,N_21599,N_20735);
nand U23006 (N_23006,N_19485,N_19493);
nand U23007 (N_23007,N_20885,N_21800);
or U23008 (N_23008,N_21868,N_19023);
nand U23009 (N_23009,N_19634,N_19156);
nor U23010 (N_23010,N_20873,N_20718);
nand U23011 (N_23011,N_21426,N_19473);
nand U23012 (N_23012,N_21096,N_20783);
nand U23013 (N_23013,N_19765,N_20855);
nor U23014 (N_23014,N_21823,N_19915);
nor U23015 (N_23015,N_20524,N_20049);
or U23016 (N_23016,N_18960,N_21178);
or U23017 (N_23017,N_20092,N_19876);
and U23018 (N_23018,N_20531,N_19136);
or U23019 (N_23019,N_20255,N_19435);
or U23020 (N_23020,N_18939,N_21267);
nor U23021 (N_23021,N_20941,N_18914);
xnor U23022 (N_23022,N_20241,N_20742);
and U23023 (N_23023,N_21121,N_21056);
nor U23024 (N_23024,N_21254,N_20415);
nor U23025 (N_23025,N_20474,N_20020);
or U23026 (N_23026,N_20443,N_20346);
and U23027 (N_23027,N_21024,N_21464);
nor U23028 (N_23028,N_21763,N_19924);
nor U23029 (N_23029,N_19299,N_21685);
or U23030 (N_23030,N_21430,N_20689);
nand U23031 (N_23031,N_19871,N_18805);
nor U23032 (N_23032,N_20922,N_18920);
or U23033 (N_23033,N_21141,N_20765);
nand U23034 (N_23034,N_20105,N_18865);
and U23035 (N_23035,N_21517,N_21818);
or U23036 (N_23036,N_19427,N_21119);
nand U23037 (N_23037,N_20694,N_21797);
nor U23038 (N_23038,N_21495,N_19455);
nor U23039 (N_23039,N_21751,N_19712);
or U23040 (N_23040,N_21774,N_19203);
nand U23041 (N_23041,N_20034,N_19535);
nand U23042 (N_23042,N_19155,N_19978);
and U23043 (N_23043,N_19846,N_20164);
and U23044 (N_23044,N_19733,N_20681);
and U23045 (N_23045,N_19501,N_21561);
nand U23046 (N_23046,N_20375,N_21588);
or U23047 (N_23047,N_19036,N_19829);
and U23048 (N_23048,N_20882,N_20906);
nand U23049 (N_23049,N_21734,N_21338);
nor U23050 (N_23050,N_18874,N_19357);
nor U23051 (N_23051,N_19613,N_21213);
and U23052 (N_23052,N_20562,N_19774);
and U23053 (N_23053,N_20721,N_20794);
and U23054 (N_23054,N_21148,N_20252);
nor U23055 (N_23055,N_20245,N_19867);
nor U23056 (N_23056,N_19269,N_18972);
or U23057 (N_23057,N_20720,N_21539);
nand U23058 (N_23058,N_19808,N_20228);
nand U23059 (N_23059,N_21565,N_20066);
nand U23060 (N_23060,N_21798,N_20648);
nor U23061 (N_23061,N_20983,N_19391);
and U23062 (N_23062,N_21810,N_21350);
or U23063 (N_23063,N_18968,N_19281);
nor U23064 (N_23064,N_20933,N_20713);
nor U23065 (N_23065,N_20914,N_20349);
nor U23066 (N_23066,N_21382,N_20512);
nor U23067 (N_23067,N_21535,N_19231);
nand U23068 (N_23068,N_20324,N_21197);
nand U23069 (N_23069,N_19284,N_19387);
and U23070 (N_23070,N_21813,N_21438);
or U23071 (N_23071,N_18837,N_19367);
and U23072 (N_23072,N_21738,N_18902);
xnor U23073 (N_23073,N_20099,N_21205);
xnor U23074 (N_23074,N_20012,N_20290);
or U23075 (N_23075,N_20931,N_19810);
xnor U23076 (N_23076,N_19591,N_20389);
nand U23077 (N_23077,N_19561,N_19514);
nor U23078 (N_23078,N_19302,N_20000);
nor U23079 (N_23079,N_19537,N_20154);
or U23080 (N_23080,N_20396,N_19674);
nand U23081 (N_23081,N_20990,N_19966);
and U23082 (N_23082,N_19954,N_19239);
and U23083 (N_23083,N_21052,N_19921);
and U23084 (N_23084,N_18753,N_21855);
xnor U23085 (N_23085,N_21576,N_20263);
or U23086 (N_23086,N_20719,N_18804);
and U23087 (N_23087,N_20102,N_19491);
xnor U23088 (N_23088,N_19585,N_20384);
and U23089 (N_23089,N_19521,N_19121);
or U23090 (N_23090,N_21002,N_21429);
nand U23091 (N_23091,N_19836,N_20700);
nor U23092 (N_23092,N_20056,N_18887);
nand U23093 (N_23093,N_18967,N_21632);
nand U23094 (N_23094,N_18760,N_21680);
xnor U23095 (N_23095,N_20534,N_19055);
and U23096 (N_23096,N_20137,N_20808);
or U23097 (N_23097,N_19832,N_20589);
nand U23098 (N_23098,N_20792,N_20208);
or U23099 (N_23099,N_21725,N_21385);
and U23100 (N_23100,N_20060,N_19366);
or U23101 (N_23101,N_19597,N_20024);
nor U23102 (N_23102,N_20880,N_20651);
and U23103 (N_23103,N_19855,N_20455);
nor U23104 (N_23104,N_18763,N_21113);
or U23105 (N_23105,N_19460,N_21406);
and U23106 (N_23106,N_21841,N_19160);
and U23107 (N_23107,N_19630,N_19804);
nand U23108 (N_23108,N_18832,N_21549);
and U23109 (N_23109,N_21499,N_20392);
and U23110 (N_23110,N_18907,N_20224);
and U23111 (N_23111,N_20893,N_19325);
or U23112 (N_23112,N_21871,N_21005);
or U23113 (N_23113,N_20144,N_20625);
nand U23114 (N_23114,N_21089,N_20190);
xnor U23115 (N_23115,N_19141,N_19848);
or U23116 (N_23116,N_21781,N_21450);
or U23117 (N_23117,N_21821,N_21391);
and U23118 (N_23118,N_20950,N_20229);
nand U23119 (N_23119,N_21587,N_20682);
nor U23120 (N_23120,N_18941,N_20356);
nor U23121 (N_23121,N_20649,N_19947);
xor U23122 (N_23122,N_18820,N_21180);
or U23123 (N_23123,N_18835,N_19509);
nor U23124 (N_23124,N_20703,N_21384);
nor U23125 (N_23125,N_19361,N_19154);
nand U23126 (N_23126,N_20996,N_19835);
xor U23127 (N_23127,N_21387,N_21210);
nor U23128 (N_23128,N_18812,N_20437);
nor U23129 (N_23129,N_19957,N_19492);
nand U23130 (N_23130,N_20367,N_20388);
nand U23131 (N_23131,N_19145,N_19862);
or U23132 (N_23132,N_19328,N_18931);
or U23133 (N_23133,N_21607,N_21809);
and U23134 (N_23134,N_20857,N_20382);
or U23135 (N_23135,N_19828,N_20925);
or U23136 (N_23136,N_20640,N_21577);
nor U23137 (N_23137,N_20809,N_20753);
xor U23138 (N_23138,N_19599,N_20638);
or U23139 (N_23139,N_20874,N_19309);
nor U23140 (N_23140,N_20660,N_20947);
or U23141 (N_23141,N_20409,N_21874);
nor U23142 (N_23142,N_21168,N_18761);
nor U23143 (N_23143,N_21702,N_21341);
nand U23144 (N_23144,N_19483,N_18830);
or U23145 (N_23145,N_20731,N_18929);
or U23146 (N_23146,N_18964,N_20769);
nand U23147 (N_23147,N_19478,N_20756);
or U23148 (N_23148,N_20076,N_21498);
or U23149 (N_23149,N_18896,N_19544);
nor U23150 (N_23150,N_21610,N_20782);
xnor U23151 (N_23151,N_20466,N_20619);
or U23152 (N_23152,N_21745,N_20511);
nand U23153 (N_23153,N_20440,N_20109);
and U23154 (N_23154,N_20658,N_21615);
and U23155 (N_23155,N_19874,N_20086);
nand U23156 (N_23156,N_20936,N_20293);
nor U23157 (N_23157,N_19084,N_20590);
nand U23158 (N_23158,N_21449,N_19595);
nand U23159 (N_23159,N_21351,N_21011);
nor U23160 (N_23160,N_19910,N_20647);
nor U23161 (N_23161,N_20820,N_20844);
nand U23162 (N_23162,N_20970,N_20318);
nor U23163 (N_23163,N_20272,N_20332);
nand U23164 (N_23164,N_21117,N_21580);
or U23165 (N_23165,N_20652,N_20269);
and U23166 (N_23166,N_20834,N_20791);
xor U23167 (N_23167,N_20432,N_21143);
nor U23168 (N_23168,N_21717,N_21128);
nor U23169 (N_23169,N_20418,N_20064);
nor U23170 (N_23170,N_19348,N_19715);
nor U23171 (N_23171,N_19047,N_19993);
nand U23172 (N_23172,N_21722,N_20219);
and U23173 (N_23173,N_21294,N_21768);
and U23174 (N_23174,N_19220,N_19856);
nand U23175 (N_23175,N_21783,N_21492);
and U23176 (N_23176,N_21022,N_21628);
xor U23177 (N_23177,N_19333,N_19627);
and U23178 (N_23178,N_19059,N_21264);
nand U23179 (N_23179,N_20656,N_20875);
nor U23180 (N_23180,N_20296,N_21835);
nor U23181 (N_23181,N_21506,N_19376);
nor U23182 (N_23182,N_21807,N_20061);
nand U23183 (N_23183,N_18759,N_20685);
and U23184 (N_23184,N_21730,N_21839);
nor U23185 (N_23185,N_20328,N_19253);
nor U23186 (N_23186,N_19158,N_21084);
and U23187 (N_23187,N_20112,N_19615);
nand U23188 (N_23188,N_20764,N_18801);
or U23189 (N_23189,N_18841,N_18777);
nor U23190 (N_23190,N_21521,N_19821);
and U23191 (N_23191,N_21791,N_18794);
and U23192 (N_23192,N_20185,N_21287);
nor U23193 (N_23193,N_20380,N_20300);
nand U23194 (N_23194,N_19471,N_20330);
nand U23195 (N_23195,N_20611,N_19445);
or U23196 (N_23196,N_19334,N_19531);
nand U23197 (N_23197,N_21386,N_20129);
and U23198 (N_23198,N_20460,N_18822);
nand U23199 (N_23199,N_19021,N_19817);
xor U23200 (N_23200,N_19980,N_19878);
nor U23201 (N_23201,N_19903,N_20013);
or U23202 (N_23202,N_21139,N_20861);
or U23203 (N_23203,N_18813,N_18984);
xor U23204 (N_23204,N_21250,N_21827);
nor U23205 (N_23205,N_19696,N_20597);
or U23206 (N_23206,N_19914,N_20645);
nand U23207 (N_23207,N_20594,N_21277);
nand U23208 (N_23208,N_19405,N_19472);
or U23209 (N_23209,N_20946,N_19811);
xor U23210 (N_23210,N_21280,N_21080);
nor U23211 (N_23211,N_21536,N_20557);
nand U23212 (N_23212,N_21083,N_19408);
xnor U23213 (N_23213,N_21705,N_20277);
nand U23214 (N_23214,N_19578,N_19228);
or U23215 (N_23215,N_19860,N_21756);
nor U23216 (N_23216,N_20148,N_19216);
or U23217 (N_23217,N_20181,N_21691);
nor U23218 (N_23218,N_19938,N_21201);
nand U23219 (N_23219,N_19854,N_20751);
nor U23220 (N_23220,N_19870,N_21175);
nand U23221 (N_23221,N_20504,N_20168);
nand U23222 (N_23222,N_19017,N_19559);
nor U23223 (N_23223,N_20863,N_19533);
and U23224 (N_23224,N_20029,N_18978);
nor U23225 (N_23225,N_20888,N_20285);
xnor U23226 (N_23226,N_19258,N_18864);
or U23227 (N_23227,N_20698,N_19749);
or U23228 (N_23228,N_19428,N_19211);
or U23229 (N_23229,N_19157,N_20842);
nand U23230 (N_23230,N_21688,N_19283);
and U23231 (N_23231,N_21241,N_20122);
nand U23232 (N_23232,N_20559,N_20114);
xnor U23233 (N_23233,N_19581,N_19673);
xor U23234 (N_23234,N_21392,N_21399);
nand U23235 (N_23235,N_19401,N_20286);
nand U23236 (N_23236,N_21260,N_21867);
or U23237 (N_23237,N_19838,N_18850);
nor U23238 (N_23238,N_21182,N_19672);
xnor U23239 (N_23239,N_21463,N_20556);
and U23240 (N_23240,N_20617,N_20162);
or U23241 (N_23241,N_18942,N_19520);
and U23242 (N_23242,N_19730,N_21633);
nor U23243 (N_23243,N_19248,N_20928);
or U23244 (N_23244,N_19127,N_21574);
and U23245 (N_23245,N_20759,N_19935);
nor U23246 (N_23246,N_21727,N_19100);
or U23247 (N_23247,N_19789,N_19825);
or U23248 (N_23248,N_19480,N_21766);
nor U23249 (N_23249,N_19374,N_18847);
nor U23250 (N_23250,N_19486,N_21192);
nor U23251 (N_23251,N_18916,N_19989);
nor U23252 (N_23252,N_21806,N_18921);
and U23253 (N_23253,N_19512,N_21804);
nor U23254 (N_23254,N_20176,N_20019);
nor U23255 (N_23255,N_20039,N_20331);
xnor U23256 (N_23256,N_21309,N_19321);
or U23257 (N_23257,N_21555,N_20593);
or U23258 (N_23258,N_19106,N_21643);
or U23259 (N_23259,N_19013,N_20015);
or U23260 (N_23260,N_20065,N_21700);
nand U23261 (N_23261,N_19496,N_19162);
xnor U23262 (N_23262,N_20900,N_20226);
nand U23263 (N_23263,N_19720,N_20784);
or U23264 (N_23264,N_19610,N_20819);
nor U23265 (N_23265,N_19506,N_21211);
or U23266 (N_23266,N_19285,N_20633);
xnor U23267 (N_23267,N_21070,N_21215);
and U23268 (N_23268,N_21433,N_19147);
and U23269 (N_23269,N_19192,N_21047);
or U23270 (N_23270,N_20447,N_20538);
and U23271 (N_23271,N_19791,N_21832);
nand U23272 (N_23272,N_19751,N_19125);
or U23273 (N_23273,N_19062,N_20247);
or U23274 (N_23274,N_20132,N_20815);
xor U23275 (N_23275,N_19922,N_21413);
or U23276 (N_23276,N_19908,N_19917);
nand U23277 (N_23277,N_18928,N_21532);
or U23278 (N_23278,N_19974,N_19434);
nor U23279 (N_23279,N_21775,N_19886);
nand U23280 (N_23280,N_20738,N_20140);
or U23281 (N_23281,N_19554,N_20311);
xor U23282 (N_23282,N_19422,N_20774);
and U23283 (N_23283,N_20587,N_20506);
nand U23284 (N_23284,N_21062,N_21054);
nand U23285 (N_23285,N_19182,N_21719);
nor U23286 (N_23286,N_20868,N_18757);
or U23287 (N_23287,N_21653,N_21772);
nand U23288 (N_23288,N_20413,N_18888);
nand U23289 (N_23289,N_21621,N_20141);
or U23290 (N_23290,N_21265,N_19621);
or U23291 (N_23291,N_20670,N_21333);
xnor U23292 (N_23292,N_20480,N_20669);
and U23293 (N_23293,N_20510,N_19359);
and U23294 (N_23294,N_19907,N_20877);
xor U23295 (N_23295,N_18918,N_19776);
nor U23296 (N_23296,N_21158,N_19661);
or U23297 (N_23297,N_19243,N_19134);
and U23298 (N_23298,N_20533,N_20309);
or U23299 (N_23299,N_20400,N_18856);
nor U23300 (N_23300,N_21105,N_20223);
and U23301 (N_23301,N_21608,N_19612);
or U23302 (N_23302,N_18817,N_19420);
nor U23303 (N_23303,N_19927,N_20254);
nor U23304 (N_23304,N_20500,N_18885);
nand U23305 (N_23305,N_20568,N_20779);
and U23306 (N_23306,N_19901,N_21437);
nand U23307 (N_23307,N_21425,N_19038);
and U23308 (N_23308,N_21538,N_19041);
nor U23309 (N_23309,N_18944,N_19762);
or U23310 (N_23310,N_19984,N_21541);
and U23311 (N_23311,N_19675,N_20299);
nand U23312 (N_23312,N_21199,N_21678);
nand U23313 (N_23313,N_19377,N_21667);
or U23314 (N_23314,N_20697,N_20084);
nand U23315 (N_23315,N_18996,N_19487);
nand U23316 (N_23316,N_21152,N_19142);
or U23317 (N_23317,N_21816,N_19126);
xor U23318 (N_23318,N_20037,N_19446);
and U23319 (N_23319,N_18790,N_19028);
nor U23320 (N_23320,N_19700,N_19338);
nor U23321 (N_23321,N_21663,N_20715);
nand U23322 (N_23322,N_20090,N_19199);
nor U23323 (N_23323,N_19213,N_21360);
xnor U23324 (N_23324,N_20417,N_18846);
nor U23325 (N_23325,N_20077,N_19177);
xor U23326 (N_23326,N_19576,N_19437);
nor U23327 (N_23327,N_20450,N_19868);
and U23328 (N_23328,N_18828,N_20008);
nor U23329 (N_23329,N_21262,N_18872);
nand U23330 (N_23330,N_21356,N_19172);
and U23331 (N_23331,N_19118,N_20994);
and U23332 (N_23332,N_20544,N_21649);
nand U23333 (N_23333,N_20949,N_20505);
nand U23334 (N_23334,N_21468,N_20327);
nor U23335 (N_23335,N_20543,N_21616);
and U23336 (N_23336,N_21456,N_20238);
nor U23337 (N_23337,N_21300,N_20452);
or U23338 (N_23338,N_21669,N_19459);
and U23339 (N_23339,N_20134,N_20200);
or U23340 (N_23340,N_19421,N_19983);
or U23341 (N_23341,N_20987,N_21660);
nor U23342 (N_23342,N_20519,N_19482);
nand U23343 (N_23343,N_21335,N_21043);
and U23344 (N_23344,N_21844,N_21239);
nand U23345 (N_23345,N_20607,N_19476);
or U23346 (N_23346,N_19945,N_21053);
nor U23347 (N_23347,N_20117,N_19643);
nor U23348 (N_23348,N_21118,N_19596);
and U23349 (N_23349,N_19640,N_20343);
nor U23350 (N_23350,N_20515,N_21367);
nor U23351 (N_23351,N_20850,N_19942);
xor U23352 (N_23352,N_21198,N_20503);
or U23353 (N_23353,N_19241,N_20214);
nor U23354 (N_23354,N_19498,N_19639);
or U23355 (N_23355,N_19029,N_20010);
nand U23356 (N_23356,N_20239,N_20580);
nand U23357 (N_23357,N_19384,N_21659);
nor U23358 (N_23358,N_19842,N_20305);
or U23359 (N_23359,N_20235,N_20864);
and U23360 (N_23360,N_21296,N_20412);
or U23361 (N_23361,N_19962,N_19327);
nand U23362 (N_23362,N_21443,N_20749);
and U23363 (N_23363,N_21481,N_21566);
or U23364 (N_23364,N_21028,N_20491);
xor U23365 (N_23365,N_19822,N_20558);
nor U23366 (N_23366,N_19764,N_21261);
and U23367 (N_23367,N_21396,N_19102);
nand U23368 (N_23368,N_20514,N_19879);
or U23369 (N_23369,N_21805,N_20653);
nor U23370 (N_23370,N_20312,N_19111);
nand U23371 (N_23371,N_21220,N_19757);
nand U23372 (N_23372,N_19688,N_20339);
and U23373 (N_23373,N_19246,N_21828);
nor U23374 (N_23374,N_20045,N_21848);
nand U23375 (N_23375,N_21065,N_20391);
nand U23376 (N_23376,N_20574,N_19598);
xnor U23377 (N_23377,N_19584,N_20635);
nand U23378 (N_23378,N_20628,N_18904);
and U23379 (N_23379,N_19319,N_21142);
nand U23380 (N_23380,N_19703,N_20982);
and U23381 (N_23381,N_21361,N_21619);
and U23382 (N_23382,N_19998,N_19545);
or U23383 (N_23383,N_20302,N_20044);
or U23384 (N_23384,N_20172,N_20692);
nor U23385 (N_23385,N_19548,N_20566);
xnor U23386 (N_23386,N_21171,N_19015);
nand U23387 (N_23387,N_19725,N_21134);
nand U23388 (N_23388,N_21346,N_19785);
nor U23389 (N_23389,N_19956,N_21108);
and U23390 (N_23390,N_20836,N_19417);
xnor U23391 (N_23391,N_20095,N_21187);
nand U23392 (N_23392,N_19852,N_20070);
xnor U23393 (N_23393,N_20745,N_19143);
nor U23394 (N_23394,N_20425,N_20575);
and U23395 (N_23395,N_20585,N_19351);
nor U23396 (N_23396,N_20373,N_19770);
and U23397 (N_23397,N_18985,N_18815);
and U23398 (N_23398,N_20569,N_21849);
or U23399 (N_23399,N_21170,N_21082);
nor U23400 (N_23400,N_19014,N_20177);
and U23401 (N_23401,N_20833,N_21428);
nor U23402 (N_23402,N_20156,N_19202);
nor U23403 (N_23403,N_19426,N_20676);
or U23404 (N_23404,N_21040,N_21301);
nand U23405 (N_23405,N_19784,N_21405);
and U23406 (N_23406,N_18915,N_20634);
nor U23407 (N_23407,N_20727,N_19756);
and U23408 (N_23408,N_20250,N_20126);
or U23409 (N_23409,N_21174,N_20125);
and U23410 (N_23410,N_19823,N_21764);
nor U23411 (N_23411,N_21266,N_19934);
nand U23412 (N_23412,N_19905,N_19077);
or U23413 (N_23413,N_20422,N_20551);
or U23414 (N_23414,N_19877,N_21314);
and U23415 (N_23415,N_18870,N_20014);
and U23416 (N_23416,N_20902,N_19315);
or U23417 (N_23417,N_20539,N_20549);
xnor U23418 (N_23418,N_20608,N_19858);
or U23419 (N_23419,N_19005,N_21493);
or U23420 (N_23420,N_21064,N_20336);
nor U23421 (N_23421,N_21604,N_19691);
and U23422 (N_23422,N_21590,N_20509);
xor U23423 (N_23423,N_21701,N_20261);
nand U23424 (N_23424,N_20940,N_19110);
nor U23425 (N_23425,N_21245,N_21014);
nor U23426 (N_23426,N_21173,N_20550);
and U23427 (N_23427,N_19031,N_20824);
nand U23428 (N_23428,N_21419,N_21847);
and U23429 (N_23429,N_21116,N_20754);
and U23430 (N_23430,N_21757,N_20016);
and U23431 (N_23431,N_19779,N_19946);
and U23432 (N_23432,N_20337,N_19481);
and U23433 (N_23433,N_21271,N_19218);
xor U23434 (N_23434,N_20832,N_19370);
and U23435 (N_23435,N_20840,N_19004);
and U23436 (N_23436,N_20213,N_20386);
nor U23437 (N_23437,N_19631,N_19522);
and U23438 (N_23438,N_19162,N_18849);
nor U23439 (N_23439,N_19463,N_21486);
and U23440 (N_23440,N_20943,N_21262);
nand U23441 (N_23441,N_20553,N_19874);
nand U23442 (N_23442,N_19246,N_20431);
nand U23443 (N_23443,N_20112,N_20784);
xnor U23444 (N_23444,N_19726,N_19753);
or U23445 (N_23445,N_20455,N_18830);
or U23446 (N_23446,N_19685,N_21407);
or U23447 (N_23447,N_21005,N_20607);
nor U23448 (N_23448,N_20555,N_19056);
and U23449 (N_23449,N_18947,N_20617);
xor U23450 (N_23450,N_21834,N_21027);
and U23451 (N_23451,N_19199,N_21706);
nand U23452 (N_23452,N_21434,N_21486);
nor U23453 (N_23453,N_20068,N_21448);
or U23454 (N_23454,N_20775,N_20201);
and U23455 (N_23455,N_21035,N_19289);
or U23456 (N_23456,N_19149,N_20456);
and U23457 (N_23457,N_20926,N_19844);
nor U23458 (N_23458,N_20065,N_19723);
or U23459 (N_23459,N_18849,N_20666);
nor U23460 (N_23460,N_21350,N_20473);
nor U23461 (N_23461,N_19304,N_20564);
or U23462 (N_23462,N_19939,N_20714);
nor U23463 (N_23463,N_19168,N_21393);
and U23464 (N_23464,N_19006,N_19798);
and U23465 (N_23465,N_20132,N_18760);
and U23466 (N_23466,N_21740,N_21029);
nand U23467 (N_23467,N_21787,N_21825);
xor U23468 (N_23468,N_20013,N_21300);
and U23469 (N_23469,N_20098,N_20573);
nand U23470 (N_23470,N_18991,N_19011);
and U23471 (N_23471,N_19632,N_20918);
or U23472 (N_23472,N_21080,N_20632);
xnor U23473 (N_23473,N_20489,N_20994);
and U23474 (N_23474,N_19513,N_18779);
xor U23475 (N_23475,N_19072,N_20388);
xor U23476 (N_23476,N_20002,N_19775);
and U23477 (N_23477,N_20956,N_21665);
nand U23478 (N_23478,N_21338,N_20554);
nor U23479 (N_23479,N_20812,N_20496);
nand U23480 (N_23480,N_21546,N_20840);
or U23481 (N_23481,N_21312,N_21113);
nand U23482 (N_23482,N_19345,N_21752);
or U23483 (N_23483,N_20910,N_20051);
or U23484 (N_23484,N_20830,N_20277);
nor U23485 (N_23485,N_20386,N_21153);
or U23486 (N_23486,N_19401,N_19439);
and U23487 (N_23487,N_19067,N_18865);
nor U23488 (N_23488,N_20221,N_21112);
nor U23489 (N_23489,N_20451,N_21020);
nand U23490 (N_23490,N_19652,N_19390);
and U23491 (N_23491,N_20253,N_20782);
and U23492 (N_23492,N_19864,N_20640);
nand U23493 (N_23493,N_20622,N_19262);
or U23494 (N_23494,N_20786,N_20867);
and U23495 (N_23495,N_18900,N_19459);
and U23496 (N_23496,N_19781,N_20672);
xnor U23497 (N_23497,N_19167,N_19938);
or U23498 (N_23498,N_21297,N_20515);
nor U23499 (N_23499,N_19967,N_19410);
nand U23500 (N_23500,N_21598,N_21658);
nand U23501 (N_23501,N_18869,N_20709);
and U23502 (N_23502,N_21219,N_21588);
or U23503 (N_23503,N_21100,N_20378);
nor U23504 (N_23504,N_20446,N_19978);
and U23505 (N_23505,N_21162,N_19296);
and U23506 (N_23506,N_21775,N_19734);
nor U23507 (N_23507,N_20347,N_19489);
nand U23508 (N_23508,N_18909,N_18777);
nor U23509 (N_23509,N_19528,N_20875);
nor U23510 (N_23510,N_19201,N_19633);
or U23511 (N_23511,N_21650,N_19246);
or U23512 (N_23512,N_21283,N_19870);
and U23513 (N_23513,N_18927,N_21484);
and U23514 (N_23514,N_20219,N_21003);
xnor U23515 (N_23515,N_20204,N_20718);
xnor U23516 (N_23516,N_18981,N_20022);
or U23517 (N_23517,N_21222,N_20452);
and U23518 (N_23518,N_19814,N_18991);
and U23519 (N_23519,N_19255,N_20932);
or U23520 (N_23520,N_19039,N_21081);
nor U23521 (N_23521,N_19524,N_21787);
nand U23522 (N_23522,N_21441,N_19267);
and U23523 (N_23523,N_20378,N_20240);
nand U23524 (N_23524,N_19453,N_21182);
or U23525 (N_23525,N_19001,N_20415);
and U23526 (N_23526,N_21698,N_19133);
nand U23527 (N_23527,N_19608,N_20428);
and U23528 (N_23528,N_19982,N_20491);
xnor U23529 (N_23529,N_19943,N_19379);
or U23530 (N_23530,N_20452,N_21645);
and U23531 (N_23531,N_19968,N_21652);
nand U23532 (N_23532,N_21068,N_20267);
and U23533 (N_23533,N_21679,N_20606);
xnor U23534 (N_23534,N_21153,N_20346);
or U23535 (N_23535,N_20724,N_19612);
xnor U23536 (N_23536,N_18751,N_19560);
nand U23537 (N_23537,N_20651,N_19875);
nor U23538 (N_23538,N_18790,N_21170);
nor U23539 (N_23539,N_18902,N_21482);
and U23540 (N_23540,N_20445,N_19860);
nor U23541 (N_23541,N_21189,N_21727);
or U23542 (N_23542,N_20191,N_19369);
nand U23543 (N_23543,N_20182,N_20530);
nand U23544 (N_23544,N_21103,N_19212);
or U23545 (N_23545,N_18923,N_20768);
nor U23546 (N_23546,N_19293,N_19590);
and U23547 (N_23547,N_18842,N_20302);
or U23548 (N_23548,N_21256,N_21048);
or U23549 (N_23549,N_21501,N_19864);
or U23550 (N_23550,N_20971,N_21750);
nand U23551 (N_23551,N_19431,N_18758);
and U23552 (N_23552,N_20874,N_19814);
or U23553 (N_23553,N_19228,N_19355);
xnor U23554 (N_23554,N_18889,N_20440);
xor U23555 (N_23555,N_20638,N_21809);
nor U23556 (N_23556,N_21486,N_21610);
nand U23557 (N_23557,N_19708,N_20255);
nand U23558 (N_23558,N_20140,N_19840);
nor U23559 (N_23559,N_20701,N_21778);
and U23560 (N_23560,N_19334,N_20501);
nand U23561 (N_23561,N_21682,N_18890);
nor U23562 (N_23562,N_19900,N_21385);
or U23563 (N_23563,N_19120,N_21212);
nand U23564 (N_23564,N_21500,N_19858);
nand U23565 (N_23565,N_21580,N_21029);
or U23566 (N_23566,N_21401,N_20188);
xnor U23567 (N_23567,N_20626,N_21477);
or U23568 (N_23568,N_20763,N_19502);
and U23569 (N_23569,N_20429,N_21860);
or U23570 (N_23570,N_20267,N_18989);
and U23571 (N_23571,N_21764,N_20240);
or U23572 (N_23572,N_20222,N_21202);
and U23573 (N_23573,N_20987,N_19778);
nor U23574 (N_23574,N_20395,N_21005);
xor U23575 (N_23575,N_21213,N_19043);
nor U23576 (N_23576,N_21834,N_19308);
or U23577 (N_23577,N_20798,N_21811);
or U23578 (N_23578,N_20724,N_20055);
nor U23579 (N_23579,N_19436,N_20225);
and U23580 (N_23580,N_20769,N_20799);
and U23581 (N_23581,N_20490,N_21076);
xnor U23582 (N_23582,N_19653,N_18973);
or U23583 (N_23583,N_20924,N_21653);
xor U23584 (N_23584,N_19442,N_18892);
nand U23585 (N_23585,N_19154,N_19888);
or U23586 (N_23586,N_19325,N_18979);
xor U23587 (N_23587,N_21383,N_19100);
and U23588 (N_23588,N_19470,N_21094);
nor U23589 (N_23589,N_21547,N_20253);
xor U23590 (N_23590,N_19871,N_19395);
or U23591 (N_23591,N_21756,N_21446);
xnor U23592 (N_23592,N_20762,N_21515);
nor U23593 (N_23593,N_20579,N_20677);
and U23594 (N_23594,N_20372,N_21378);
xnor U23595 (N_23595,N_21603,N_21067);
and U23596 (N_23596,N_21856,N_20031);
nor U23597 (N_23597,N_19877,N_18989);
or U23598 (N_23598,N_20326,N_20063);
nor U23599 (N_23599,N_20410,N_21497);
nand U23600 (N_23600,N_20344,N_20888);
and U23601 (N_23601,N_20890,N_21669);
or U23602 (N_23602,N_19895,N_21260);
and U23603 (N_23603,N_20052,N_20724);
nor U23604 (N_23604,N_20180,N_20504);
or U23605 (N_23605,N_19238,N_19915);
xor U23606 (N_23606,N_20202,N_21386);
or U23607 (N_23607,N_21556,N_20350);
or U23608 (N_23608,N_20179,N_20290);
nand U23609 (N_23609,N_21699,N_20605);
and U23610 (N_23610,N_21814,N_21625);
nor U23611 (N_23611,N_20871,N_21276);
and U23612 (N_23612,N_20580,N_19355);
or U23613 (N_23613,N_19775,N_19102);
nor U23614 (N_23614,N_19456,N_21225);
or U23615 (N_23615,N_20530,N_19992);
nand U23616 (N_23616,N_19036,N_20728);
and U23617 (N_23617,N_20934,N_19290);
and U23618 (N_23618,N_19758,N_21534);
nor U23619 (N_23619,N_19131,N_21569);
xor U23620 (N_23620,N_19973,N_19014);
xnor U23621 (N_23621,N_20817,N_19577);
or U23622 (N_23622,N_19161,N_20538);
and U23623 (N_23623,N_19832,N_20300);
and U23624 (N_23624,N_19858,N_18932);
or U23625 (N_23625,N_21346,N_19177);
nor U23626 (N_23626,N_21633,N_19946);
and U23627 (N_23627,N_18767,N_19847);
or U23628 (N_23628,N_20608,N_20976);
or U23629 (N_23629,N_18949,N_20459);
and U23630 (N_23630,N_18892,N_21670);
nor U23631 (N_23631,N_21740,N_19682);
nand U23632 (N_23632,N_19459,N_20139);
or U23633 (N_23633,N_18920,N_20678);
nor U23634 (N_23634,N_20876,N_19454);
nor U23635 (N_23635,N_20986,N_21188);
nand U23636 (N_23636,N_19229,N_19601);
and U23637 (N_23637,N_21423,N_19668);
nand U23638 (N_23638,N_21463,N_21672);
nand U23639 (N_23639,N_19358,N_20040);
and U23640 (N_23640,N_19822,N_20624);
or U23641 (N_23641,N_21132,N_21758);
nand U23642 (N_23642,N_18923,N_20622);
or U23643 (N_23643,N_19327,N_19576);
nor U23644 (N_23644,N_21406,N_19776);
nor U23645 (N_23645,N_20718,N_21789);
and U23646 (N_23646,N_19562,N_20786);
nor U23647 (N_23647,N_19588,N_21810);
xor U23648 (N_23648,N_20626,N_21684);
nand U23649 (N_23649,N_21116,N_20379);
nand U23650 (N_23650,N_19224,N_20920);
nor U23651 (N_23651,N_20197,N_20709);
or U23652 (N_23652,N_21000,N_21699);
xor U23653 (N_23653,N_19106,N_18930);
and U23654 (N_23654,N_19231,N_20608);
nand U23655 (N_23655,N_20589,N_20093);
nor U23656 (N_23656,N_21117,N_18907);
nand U23657 (N_23657,N_21342,N_19282);
and U23658 (N_23658,N_19362,N_19275);
nor U23659 (N_23659,N_21141,N_21065);
or U23660 (N_23660,N_21545,N_18835);
nor U23661 (N_23661,N_19595,N_21217);
or U23662 (N_23662,N_20096,N_19242);
nand U23663 (N_23663,N_20678,N_19426);
or U23664 (N_23664,N_20219,N_19861);
xor U23665 (N_23665,N_19461,N_19852);
and U23666 (N_23666,N_18922,N_19607);
nor U23667 (N_23667,N_20607,N_20745);
nand U23668 (N_23668,N_19569,N_20403);
and U23669 (N_23669,N_19218,N_20359);
or U23670 (N_23670,N_19537,N_19309);
nor U23671 (N_23671,N_19384,N_19440);
nand U23672 (N_23672,N_20496,N_18800);
or U23673 (N_23673,N_21853,N_21750);
nor U23674 (N_23674,N_19311,N_19320);
and U23675 (N_23675,N_20250,N_19043);
nor U23676 (N_23676,N_18893,N_19824);
nand U23677 (N_23677,N_18955,N_21358);
or U23678 (N_23678,N_20995,N_21399);
or U23679 (N_23679,N_20430,N_21452);
nand U23680 (N_23680,N_19492,N_21079);
or U23681 (N_23681,N_19902,N_21575);
nand U23682 (N_23682,N_19151,N_21450);
nor U23683 (N_23683,N_18815,N_20533);
and U23684 (N_23684,N_20165,N_19682);
xnor U23685 (N_23685,N_19103,N_19591);
nand U23686 (N_23686,N_21047,N_20604);
xor U23687 (N_23687,N_19961,N_19947);
or U23688 (N_23688,N_19644,N_19881);
nand U23689 (N_23689,N_21063,N_20614);
nor U23690 (N_23690,N_19138,N_20342);
nand U23691 (N_23691,N_20989,N_18751);
nor U23692 (N_23692,N_21586,N_20841);
nand U23693 (N_23693,N_19080,N_19119);
xor U23694 (N_23694,N_18933,N_20732);
nand U23695 (N_23695,N_21578,N_20904);
or U23696 (N_23696,N_21259,N_19153);
and U23697 (N_23697,N_20051,N_19712);
nor U23698 (N_23698,N_20778,N_19547);
or U23699 (N_23699,N_19599,N_20594);
or U23700 (N_23700,N_19944,N_19476);
nor U23701 (N_23701,N_20508,N_21356);
or U23702 (N_23702,N_21746,N_18836);
nor U23703 (N_23703,N_19423,N_18912);
and U23704 (N_23704,N_21034,N_21397);
nor U23705 (N_23705,N_21157,N_19918);
nand U23706 (N_23706,N_19250,N_18752);
nor U23707 (N_23707,N_19118,N_21160);
or U23708 (N_23708,N_19933,N_21258);
or U23709 (N_23709,N_21493,N_19688);
nand U23710 (N_23710,N_20970,N_21087);
nor U23711 (N_23711,N_19789,N_21232);
and U23712 (N_23712,N_21034,N_21765);
xnor U23713 (N_23713,N_19541,N_19150);
xnor U23714 (N_23714,N_18801,N_19707);
nand U23715 (N_23715,N_19798,N_20620);
or U23716 (N_23716,N_21070,N_21335);
and U23717 (N_23717,N_19238,N_20540);
xor U23718 (N_23718,N_20494,N_19985);
nand U23719 (N_23719,N_19859,N_20593);
nand U23720 (N_23720,N_20410,N_20841);
or U23721 (N_23721,N_20554,N_19543);
nor U23722 (N_23722,N_20432,N_21514);
or U23723 (N_23723,N_19597,N_21019);
nand U23724 (N_23724,N_21829,N_21579);
or U23725 (N_23725,N_20097,N_19112);
or U23726 (N_23726,N_20967,N_19268);
or U23727 (N_23727,N_19976,N_19101);
and U23728 (N_23728,N_20186,N_20309);
and U23729 (N_23729,N_21242,N_20638);
nor U23730 (N_23730,N_21463,N_20041);
nand U23731 (N_23731,N_18883,N_20105);
xor U23732 (N_23732,N_21325,N_20521);
or U23733 (N_23733,N_20994,N_19536);
and U23734 (N_23734,N_20835,N_20907);
xnor U23735 (N_23735,N_21873,N_19282);
nand U23736 (N_23736,N_19242,N_20627);
nand U23737 (N_23737,N_20801,N_21732);
nor U23738 (N_23738,N_21517,N_20090);
nor U23739 (N_23739,N_19352,N_20430);
and U23740 (N_23740,N_21383,N_20437);
and U23741 (N_23741,N_20038,N_19771);
or U23742 (N_23742,N_19557,N_19299);
nor U23743 (N_23743,N_18931,N_19354);
nor U23744 (N_23744,N_21127,N_20477);
nor U23745 (N_23745,N_21595,N_20841);
nand U23746 (N_23746,N_19423,N_20731);
xor U23747 (N_23747,N_20229,N_21076);
nor U23748 (N_23748,N_18811,N_19370);
nor U23749 (N_23749,N_21461,N_19221);
xor U23750 (N_23750,N_21508,N_21724);
nor U23751 (N_23751,N_21297,N_20024);
nand U23752 (N_23752,N_21755,N_21418);
nand U23753 (N_23753,N_18780,N_21658);
nor U23754 (N_23754,N_18870,N_21046);
nor U23755 (N_23755,N_20401,N_20936);
nor U23756 (N_23756,N_21305,N_19957);
or U23757 (N_23757,N_19437,N_20381);
nand U23758 (N_23758,N_21371,N_21171);
nor U23759 (N_23759,N_20831,N_20632);
nand U23760 (N_23760,N_21737,N_19645);
nor U23761 (N_23761,N_19235,N_21803);
nand U23762 (N_23762,N_21802,N_19562);
or U23763 (N_23763,N_21284,N_20337);
and U23764 (N_23764,N_21334,N_21499);
or U23765 (N_23765,N_21844,N_19316);
nor U23766 (N_23766,N_20116,N_18783);
nand U23767 (N_23767,N_20604,N_20904);
nor U23768 (N_23768,N_19926,N_20606);
or U23769 (N_23769,N_21864,N_19732);
or U23770 (N_23770,N_21631,N_19123);
or U23771 (N_23771,N_19754,N_18956);
nand U23772 (N_23772,N_21246,N_21265);
and U23773 (N_23773,N_20361,N_19932);
or U23774 (N_23774,N_20517,N_19266);
nand U23775 (N_23775,N_21130,N_18921);
or U23776 (N_23776,N_19376,N_20552);
nand U23777 (N_23777,N_19724,N_21093);
nor U23778 (N_23778,N_18755,N_19359);
nor U23779 (N_23779,N_19264,N_19356);
and U23780 (N_23780,N_21501,N_21339);
or U23781 (N_23781,N_19853,N_21476);
or U23782 (N_23782,N_21290,N_20997);
nand U23783 (N_23783,N_21526,N_20543);
xor U23784 (N_23784,N_19181,N_18957);
nor U23785 (N_23785,N_18855,N_18902);
nor U23786 (N_23786,N_19457,N_20680);
and U23787 (N_23787,N_20915,N_20790);
or U23788 (N_23788,N_20870,N_20052);
or U23789 (N_23789,N_19798,N_20960);
nor U23790 (N_23790,N_20773,N_20242);
and U23791 (N_23791,N_20471,N_18786);
nand U23792 (N_23792,N_21662,N_19460);
and U23793 (N_23793,N_20636,N_21388);
xnor U23794 (N_23794,N_20717,N_19034);
nand U23795 (N_23795,N_21621,N_19246);
or U23796 (N_23796,N_19649,N_21613);
or U23797 (N_23797,N_19932,N_19356);
or U23798 (N_23798,N_20990,N_21424);
or U23799 (N_23799,N_19639,N_19019);
nor U23800 (N_23800,N_21158,N_20216);
and U23801 (N_23801,N_19907,N_20791);
and U23802 (N_23802,N_21110,N_21057);
nand U23803 (N_23803,N_19904,N_20333);
nand U23804 (N_23804,N_19041,N_18893);
nand U23805 (N_23805,N_20345,N_20639);
xor U23806 (N_23806,N_20024,N_20794);
nand U23807 (N_23807,N_19986,N_20243);
or U23808 (N_23808,N_19497,N_19208);
or U23809 (N_23809,N_19852,N_19486);
or U23810 (N_23810,N_21526,N_21038);
nand U23811 (N_23811,N_20663,N_20007);
or U23812 (N_23812,N_19245,N_20914);
or U23813 (N_23813,N_18826,N_18784);
nand U23814 (N_23814,N_19056,N_20290);
or U23815 (N_23815,N_20813,N_19723);
and U23816 (N_23816,N_20764,N_19362);
or U23817 (N_23817,N_19428,N_19567);
or U23818 (N_23818,N_20633,N_19838);
and U23819 (N_23819,N_21458,N_18876);
nor U23820 (N_23820,N_20926,N_21111);
or U23821 (N_23821,N_19237,N_20234);
nand U23822 (N_23822,N_21243,N_18821);
nor U23823 (N_23823,N_19221,N_19347);
xor U23824 (N_23824,N_20972,N_20863);
nand U23825 (N_23825,N_19750,N_21272);
or U23826 (N_23826,N_21210,N_20061);
nand U23827 (N_23827,N_20275,N_19560);
and U23828 (N_23828,N_21261,N_18989);
nand U23829 (N_23829,N_20949,N_18768);
nor U23830 (N_23830,N_19805,N_20824);
or U23831 (N_23831,N_21652,N_20330);
and U23832 (N_23832,N_20456,N_21422);
nand U23833 (N_23833,N_20177,N_18911);
or U23834 (N_23834,N_20205,N_20866);
and U23835 (N_23835,N_19324,N_21710);
and U23836 (N_23836,N_21509,N_20369);
or U23837 (N_23837,N_20788,N_20499);
nor U23838 (N_23838,N_19168,N_20368);
and U23839 (N_23839,N_20306,N_19836);
nand U23840 (N_23840,N_18889,N_20005);
nor U23841 (N_23841,N_21228,N_21334);
nor U23842 (N_23842,N_21560,N_19749);
and U23843 (N_23843,N_21563,N_19532);
xor U23844 (N_23844,N_20958,N_20953);
and U23845 (N_23845,N_21054,N_21424);
and U23846 (N_23846,N_21069,N_19159);
nand U23847 (N_23847,N_20783,N_20766);
nor U23848 (N_23848,N_19010,N_19155);
xor U23849 (N_23849,N_21114,N_19766);
or U23850 (N_23850,N_21102,N_19687);
nor U23851 (N_23851,N_20069,N_20408);
or U23852 (N_23852,N_19177,N_19301);
nand U23853 (N_23853,N_20128,N_19993);
or U23854 (N_23854,N_19109,N_20746);
or U23855 (N_23855,N_19262,N_20052);
or U23856 (N_23856,N_20303,N_20986);
nand U23857 (N_23857,N_21655,N_19612);
and U23858 (N_23858,N_19920,N_19161);
and U23859 (N_23859,N_19296,N_20382);
or U23860 (N_23860,N_21643,N_21557);
nand U23861 (N_23861,N_20033,N_18775);
nand U23862 (N_23862,N_21681,N_21004);
nor U23863 (N_23863,N_20577,N_19852);
xnor U23864 (N_23864,N_21796,N_20016);
nor U23865 (N_23865,N_20575,N_20094);
nand U23866 (N_23866,N_19300,N_20323);
nand U23867 (N_23867,N_21598,N_20945);
and U23868 (N_23868,N_19062,N_20936);
xnor U23869 (N_23869,N_18894,N_18840);
xor U23870 (N_23870,N_20497,N_19658);
and U23871 (N_23871,N_20108,N_21166);
or U23872 (N_23872,N_20695,N_19077);
and U23873 (N_23873,N_20002,N_19491);
nor U23874 (N_23874,N_19422,N_20123);
or U23875 (N_23875,N_21488,N_20661);
or U23876 (N_23876,N_18831,N_20951);
or U23877 (N_23877,N_21639,N_19456);
nor U23878 (N_23878,N_21137,N_21548);
or U23879 (N_23879,N_20047,N_18836);
or U23880 (N_23880,N_20773,N_19012);
nor U23881 (N_23881,N_18760,N_21233);
nor U23882 (N_23882,N_19138,N_19777);
nor U23883 (N_23883,N_20520,N_20419);
and U23884 (N_23884,N_20324,N_20525);
or U23885 (N_23885,N_20843,N_21581);
and U23886 (N_23886,N_19697,N_20887);
or U23887 (N_23887,N_20134,N_19046);
or U23888 (N_23888,N_20508,N_20215);
and U23889 (N_23889,N_19174,N_20989);
and U23890 (N_23890,N_20227,N_19694);
or U23891 (N_23891,N_21645,N_20322);
or U23892 (N_23892,N_20511,N_21855);
xnor U23893 (N_23893,N_18892,N_19515);
and U23894 (N_23894,N_21802,N_21258);
nand U23895 (N_23895,N_19829,N_21047);
nor U23896 (N_23896,N_21135,N_20032);
nand U23897 (N_23897,N_21167,N_20964);
xor U23898 (N_23898,N_19383,N_20623);
and U23899 (N_23899,N_21506,N_21202);
and U23900 (N_23900,N_20436,N_19104);
or U23901 (N_23901,N_21766,N_19382);
nor U23902 (N_23902,N_20105,N_19290);
or U23903 (N_23903,N_21864,N_19368);
nand U23904 (N_23904,N_20967,N_21815);
nor U23905 (N_23905,N_18928,N_20667);
and U23906 (N_23906,N_19390,N_21561);
or U23907 (N_23907,N_21280,N_20362);
xnor U23908 (N_23908,N_19478,N_20044);
nand U23909 (N_23909,N_19630,N_20956);
and U23910 (N_23910,N_21537,N_20376);
nand U23911 (N_23911,N_19761,N_21464);
xnor U23912 (N_23912,N_20154,N_20960);
or U23913 (N_23913,N_19310,N_21346);
nor U23914 (N_23914,N_20855,N_21175);
or U23915 (N_23915,N_20420,N_20705);
or U23916 (N_23916,N_19700,N_19725);
or U23917 (N_23917,N_20623,N_20766);
nand U23918 (N_23918,N_19869,N_20351);
and U23919 (N_23919,N_20665,N_21849);
or U23920 (N_23920,N_19523,N_20199);
or U23921 (N_23921,N_20834,N_19192);
nand U23922 (N_23922,N_19674,N_21020);
and U23923 (N_23923,N_19135,N_21461);
and U23924 (N_23924,N_20849,N_19072);
nand U23925 (N_23925,N_20740,N_21051);
or U23926 (N_23926,N_21726,N_19679);
or U23927 (N_23927,N_18801,N_21810);
or U23928 (N_23928,N_20588,N_21755);
and U23929 (N_23929,N_18978,N_20942);
nor U23930 (N_23930,N_19880,N_20055);
or U23931 (N_23931,N_19433,N_19997);
or U23932 (N_23932,N_20259,N_21101);
nand U23933 (N_23933,N_21236,N_19556);
nor U23934 (N_23934,N_21864,N_21562);
nor U23935 (N_23935,N_18912,N_18984);
and U23936 (N_23936,N_20649,N_21108);
and U23937 (N_23937,N_21419,N_20177);
xor U23938 (N_23938,N_20276,N_21366);
nor U23939 (N_23939,N_20866,N_21028);
xor U23940 (N_23940,N_20244,N_18840);
or U23941 (N_23941,N_21625,N_21641);
nor U23942 (N_23942,N_20843,N_19516);
and U23943 (N_23943,N_21282,N_19971);
and U23944 (N_23944,N_20725,N_18967);
nor U23945 (N_23945,N_18766,N_21087);
nor U23946 (N_23946,N_21741,N_19926);
and U23947 (N_23947,N_19430,N_19075);
nand U23948 (N_23948,N_19129,N_19647);
and U23949 (N_23949,N_20486,N_21225);
xnor U23950 (N_23950,N_19567,N_20940);
xor U23951 (N_23951,N_20605,N_21437);
or U23952 (N_23952,N_18790,N_20000);
and U23953 (N_23953,N_19120,N_21274);
nor U23954 (N_23954,N_21579,N_19693);
nand U23955 (N_23955,N_21409,N_21207);
nor U23956 (N_23956,N_20443,N_18900);
nor U23957 (N_23957,N_20598,N_20904);
and U23958 (N_23958,N_20369,N_21733);
and U23959 (N_23959,N_19647,N_21480);
nand U23960 (N_23960,N_20307,N_20567);
xnor U23961 (N_23961,N_18842,N_20775);
or U23962 (N_23962,N_19741,N_18934);
and U23963 (N_23963,N_20700,N_21782);
and U23964 (N_23964,N_19766,N_19548);
or U23965 (N_23965,N_20261,N_21840);
and U23966 (N_23966,N_20878,N_20630);
xnor U23967 (N_23967,N_19362,N_20069);
nor U23968 (N_23968,N_21304,N_19478);
nor U23969 (N_23969,N_21553,N_19952);
nor U23970 (N_23970,N_20369,N_20756);
nand U23971 (N_23971,N_19053,N_19206);
and U23972 (N_23972,N_20068,N_19230);
xor U23973 (N_23973,N_19675,N_18798);
and U23974 (N_23974,N_20498,N_20167);
or U23975 (N_23975,N_18840,N_19891);
or U23976 (N_23976,N_19065,N_19680);
nor U23977 (N_23977,N_19571,N_21808);
nor U23978 (N_23978,N_19826,N_21040);
nand U23979 (N_23979,N_21698,N_19519);
nor U23980 (N_23980,N_19037,N_21750);
or U23981 (N_23981,N_20369,N_20175);
or U23982 (N_23982,N_19156,N_21558);
or U23983 (N_23983,N_20620,N_20262);
or U23984 (N_23984,N_19347,N_19025);
nand U23985 (N_23985,N_21114,N_21562);
nand U23986 (N_23986,N_19758,N_19567);
and U23987 (N_23987,N_19047,N_21125);
and U23988 (N_23988,N_19343,N_20052);
or U23989 (N_23989,N_19776,N_19605);
and U23990 (N_23990,N_21415,N_21476);
or U23991 (N_23991,N_19905,N_19144);
xnor U23992 (N_23992,N_21472,N_19303);
nand U23993 (N_23993,N_20983,N_19219);
nor U23994 (N_23994,N_21216,N_20951);
nand U23995 (N_23995,N_21173,N_20150);
nor U23996 (N_23996,N_18840,N_20735);
and U23997 (N_23997,N_20776,N_20228);
and U23998 (N_23998,N_19249,N_21547);
nand U23999 (N_23999,N_21297,N_21797);
nor U24000 (N_24000,N_21866,N_19831);
or U24001 (N_24001,N_20610,N_20688);
and U24002 (N_24002,N_19383,N_19268);
nand U24003 (N_24003,N_19669,N_21736);
or U24004 (N_24004,N_21379,N_20267);
nor U24005 (N_24005,N_19304,N_20438);
and U24006 (N_24006,N_21782,N_20815);
and U24007 (N_24007,N_20159,N_19079);
nand U24008 (N_24008,N_21201,N_19438);
xor U24009 (N_24009,N_21148,N_21608);
nand U24010 (N_24010,N_19784,N_20652);
nand U24011 (N_24011,N_20412,N_20981);
nand U24012 (N_24012,N_20215,N_19679);
xor U24013 (N_24013,N_21727,N_21287);
or U24014 (N_24014,N_21860,N_20720);
nor U24015 (N_24015,N_19289,N_18866);
nand U24016 (N_24016,N_20427,N_20620);
nor U24017 (N_24017,N_19195,N_19012);
and U24018 (N_24018,N_18909,N_21224);
and U24019 (N_24019,N_20758,N_20706);
nand U24020 (N_24020,N_18876,N_21675);
and U24021 (N_24021,N_20482,N_19228);
nand U24022 (N_24022,N_21689,N_19070);
or U24023 (N_24023,N_21123,N_19045);
nor U24024 (N_24024,N_20143,N_20450);
and U24025 (N_24025,N_21198,N_19877);
and U24026 (N_24026,N_19533,N_20473);
nand U24027 (N_24027,N_19011,N_18932);
nand U24028 (N_24028,N_19873,N_20785);
nor U24029 (N_24029,N_20573,N_19501);
or U24030 (N_24030,N_20286,N_21670);
xor U24031 (N_24031,N_21571,N_19659);
nand U24032 (N_24032,N_21059,N_20580);
nor U24033 (N_24033,N_19694,N_18915);
or U24034 (N_24034,N_19678,N_19730);
nor U24035 (N_24035,N_19446,N_20699);
or U24036 (N_24036,N_20776,N_19733);
nand U24037 (N_24037,N_20281,N_20943);
xnor U24038 (N_24038,N_21755,N_21702);
and U24039 (N_24039,N_21823,N_19165);
and U24040 (N_24040,N_21019,N_18794);
xor U24041 (N_24041,N_20059,N_21509);
nor U24042 (N_24042,N_18822,N_20174);
xnor U24043 (N_24043,N_19871,N_21715);
or U24044 (N_24044,N_19256,N_18817);
or U24045 (N_24045,N_20578,N_20338);
and U24046 (N_24046,N_21262,N_19378);
nor U24047 (N_24047,N_20037,N_19581);
nor U24048 (N_24048,N_20086,N_19718);
nor U24049 (N_24049,N_19621,N_21438);
nand U24050 (N_24050,N_20248,N_19909);
and U24051 (N_24051,N_19807,N_21415);
or U24052 (N_24052,N_18960,N_19277);
and U24053 (N_24053,N_19957,N_20577);
and U24054 (N_24054,N_20710,N_19793);
nand U24055 (N_24055,N_19431,N_19772);
xnor U24056 (N_24056,N_21230,N_18880);
nand U24057 (N_24057,N_19419,N_20529);
nor U24058 (N_24058,N_20750,N_20209);
nand U24059 (N_24059,N_18791,N_21355);
nor U24060 (N_24060,N_21043,N_20668);
or U24061 (N_24061,N_20043,N_21339);
or U24062 (N_24062,N_18922,N_20658);
nor U24063 (N_24063,N_19495,N_18811);
xor U24064 (N_24064,N_20522,N_19632);
and U24065 (N_24065,N_20405,N_21044);
nor U24066 (N_24066,N_21583,N_18917);
nor U24067 (N_24067,N_21590,N_18961);
and U24068 (N_24068,N_21294,N_19955);
nor U24069 (N_24069,N_21130,N_19503);
nand U24070 (N_24070,N_19800,N_19836);
and U24071 (N_24071,N_21401,N_18796);
and U24072 (N_24072,N_21791,N_18807);
or U24073 (N_24073,N_20132,N_20174);
nand U24074 (N_24074,N_19622,N_21150);
or U24075 (N_24075,N_21197,N_20201);
xor U24076 (N_24076,N_20652,N_19749);
nand U24077 (N_24077,N_19164,N_21165);
or U24078 (N_24078,N_21810,N_19956);
and U24079 (N_24079,N_20927,N_20529);
nor U24080 (N_24080,N_20146,N_21200);
and U24081 (N_24081,N_20696,N_20205);
xor U24082 (N_24082,N_18981,N_21445);
or U24083 (N_24083,N_20045,N_20188);
nor U24084 (N_24084,N_20040,N_21107);
and U24085 (N_24085,N_19928,N_20179);
nor U24086 (N_24086,N_21019,N_20026);
or U24087 (N_24087,N_21472,N_19411);
or U24088 (N_24088,N_20389,N_18865);
or U24089 (N_24089,N_19336,N_21349);
and U24090 (N_24090,N_19814,N_21254);
xnor U24091 (N_24091,N_19570,N_21283);
and U24092 (N_24092,N_21712,N_19562);
or U24093 (N_24093,N_19697,N_21199);
or U24094 (N_24094,N_20126,N_19695);
nor U24095 (N_24095,N_21746,N_18905);
nand U24096 (N_24096,N_20271,N_19047);
nor U24097 (N_24097,N_20435,N_20814);
xor U24098 (N_24098,N_20958,N_20766);
or U24099 (N_24099,N_21820,N_19478);
or U24100 (N_24100,N_20952,N_21133);
nor U24101 (N_24101,N_19344,N_20168);
nor U24102 (N_24102,N_21648,N_20947);
or U24103 (N_24103,N_19490,N_21495);
nor U24104 (N_24104,N_19486,N_20562);
nor U24105 (N_24105,N_19746,N_21120);
xor U24106 (N_24106,N_20204,N_21441);
nand U24107 (N_24107,N_20261,N_21143);
nor U24108 (N_24108,N_19687,N_21137);
or U24109 (N_24109,N_20944,N_19325);
and U24110 (N_24110,N_20343,N_19714);
and U24111 (N_24111,N_19080,N_19238);
nand U24112 (N_24112,N_21727,N_19103);
nand U24113 (N_24113,N_19477,N_20166);
or U24114 (N_24114,N_19173,N_19025);
nand U24115 (N_24115,N_18954,N_20189);
and U24116 (N_24116,N_21649,N_21224);
and U24117 (N_24117,N_19837,N_18928);
and U24118 (N_24118,N_21071,N_19994);
nand U24119 (N_24119,N_19564,N_21162);
nor U24120 (N_24120,N_19553,N_20942);
or U24121 (N_24121,N_20398,N_20215);
and U24122 (N_24122,N_19871,N_19034);
and U24123 (N_24123,N_19606,N_20335);
or U24124 (N_24124,N_20277,N_19305);
nand U24125 (N_24125,N_19944,N_20262);
or U24126 (N_24126,N_20514,N_21497);
nor U24127 (N_24127,N_20805,N_21217);
nor U24128 (N_24128,N_20918,N_20311);
nand U24129 (N_24129,N_21778,N_19061);
or U24130 (N_24130,N_21454,N_18832);
or U24131 (N_24131,N_19341,N_19694);
nor U24132 (N_24132,N_20589,N_21283);
nand U24133 (N_24133,N_18800,N_20824);
nand U24134 (N_24134,N_19219,N_20252);
and U24135 (N_24135,N_19275,N_19044);
nor U24136 (N_24136,N_20507,N_19339);
and U24137 (N_24137,N_20074,N_20426);
nand U24138 (N_24138,N_20468,N_20820);
nor U24139 (N_24139,N_19232,N_20467);
or U24140 (N_24140,N_18765,N_19056);
nor U24141 (N_24141,N_20944,N_19768);
nor U24142 (N_24142,N_21442,N_18863);
and U24143 (N_24143,N_19766,N_21415);
nand U24144 (N_24144,N_21064,N_18761);
and U24145 (N_24145,N_21296,N_20507);
or U24146 (N_24146,N_20410,N_20950);
and U24147 (N_24147,N_19893,N_19295);
and U24148 (N_24148,N_20850,N_19175);
nor U24149 (N_24149,N_19748,N_21188);
nand U24150 (N_24150,N_21335,N_18877);
or U24151 (N_24151,N_21423,N_18834);
or U24152 (N_24152,N_20330,N_20788);
and U24153 (N_24153,N_20915,N_19160);
or U24154 (N_24154,N_21341,N_19570);
nor U24155 (N_24155,N_20124,N_20070);
and U24156 (N_24156,N_19017,N_19845);
nand U24157 (N_24157,N_19474,N_20855);
nand U24158 (N_24158,N_20902,N_18865);
and U24159 (N_24159,N_19748,N_20479);
nand U24160 (N_24160,N_20517,N_19134);
nor U24161 (N_24161,N_19504,N_21821);
and U24162 (N_24162,N_21787,N_20412);
nor U24163 (N_24163,N_20899,N_18783);
xor U24164 (N_24164,N_21064,N_21212);
xor U24165 (N_24165,N_18784,N_19532);
and U24166 (N_24166,N_20646,N_21135);
and U24167 (N_24167,N_19595,N_20758);
nor U24168 (N_24168,N_20322,N_21408);
nor U24169 (N_24169,N_20788,N_20678);
nand U24170 (N_24170,N_21752,N_20632);
and U24171 (N_24171,N_19542,N_21455);
or U24172 (N_24172,N_21780,N_18919);
or U24173 (N_24173,N_19846,N_20554);
nor U24174 (N_24174,N_18795,N_21095);
and U24175 (N_24175,N_19279,N_20988);
or U24176 (N_24176,N_19473,N_19891);
nand U24177 (N_24177,N_21705,N_18752);
or U24178 (N_24178,N_21186,N_19044);
and U24179 (N_24179,N_19854,N_20975);
and U24180 (N_24180,N_21323,N_20315);
and U24181 (N_24181,N_18928,N_21109);
xor U24182 (N_24182,N_20156,N_18929);
nand U24183 (N_24183,N_21647,N_19051);
or U24184 (N_24184,N_20536,N_20323);
nor U24185 (N_24185,N_19344,N_18809);
or U24186 (N_24186,N_21873,N_19494);
or U24187 (N_24187,N_21344,N_21457);
and U24188 (N_24188,N_19216,N_21332);
and U24189 (N_24189,N_20772,N_19812);
or U24190 (N_24190,N_20461,N_21633);
nor U24191 (N_24191,N_19438,N_21031);
and U24192 (N_24192,N_19045,N_20630);
xnor U24193 (N_24193,N_19862,N_20784);
and U24194 (N_24194,N_20315,N_18807);
and U24195 (N_24195,N_20120,N_19292);
xnor U24196 (N_24196,N_20331,N_21443);
and U24197 (N_24197,N_19517,N_21451);
and U24198 (N_24198,N_21447,N_20583);
and U24199 (N_24199,N_21151,N_19641);
nor U24200 (N_24200,N_18783,N_20252);
xnor U24201 (N_24201,N_20411,N_20866);
nor U24202 (N_24202,N_19033,N_21732);
nor U24203 (N_24203,N_21024,N_19416);
and U24204 (N_24204,N_21319,N_19849);
or U24205 (N_24205,N_19629,N_21189);
nor U24206 (N_24206,N_20976,N_20265);
nor U24207 (N_24207,N_19302,N_21180);
nor U24208 (N_24208,N_19279,N_21465);
nor U24209 (N_24209,N_20139,N_21236);
and U24210 (N_24210,N_21735,N_20269);
nor U24211 (N_24211,N_20139,N_21745);
nor U24212 (N_24212,N_20977,N_20911);
nand U24213 (N_24213,N_19105,N_19274);
nand U24214 (N_24214,N_20542,N_19056);
or U24215 (N_24215,N_18894,N_20865);
xnor U24216 (N_24216,N_20298,N_18933);
or U24217 (N_24217,N_20509,N_20599);
and U24218 (N_24218,N_19088,N_21515);
or U24219 (N_24219,N_20529,N_21606);
xor U24220 (N_24220,N_19424,N_18999);
nor U24221 (N_24221,N_21515,N_21301);
and U24222 (N_24222,N_19057,N_21708);
or U24223 (N_24223,N_20439,N_21707);
and U24224 (N_24224,N_19528,N_19035);
nor U24225 (N_24225,N_19110,N_18780);
nand U24226 (N_24226,N_20278,N_21070);
xnor U24227 (N_24227,N_20713,N_19229);
nand U24228 (N_24228,N_20127,N_19363);
nor U24229 (N_24229,N_19940,N_20291);
or U24230 (N_24230,N_19992,N_21124);
and U24231 (N_24231,N_20478,N_20055);
and U24232 (N_24232,N_19184,N_21022);
nor U24233 (N_24233,N_20815,N_19383);
nand U24234 (N_24234,N_21238,N_19632);
and U24235 (N_24235,N_19129,N_19459);
or U24236 (N_24236,N_21810,N_20162);
and U24237 (N_24237,N_20888,N_21221);
xor U24238 (N_24238,N_20686,N_19675);
or U24239 (N_24239,N_20307,N_20674);
or U24240 (N_24240,N_18810,N_21679);
or U24241 (N_24241,N_20875,N_20528);
nand U24242 (N_24242,N_20932,N_20679);
nand U24243 (N_24243,N_20487,N_18795);
nand U24244 (N_24244,N_21078,N_19868);
nand U24245 (N_24245,N_21754,N_21020);
nor U24246 (N_24246,N_20281,N_21227);
nand U24247 (N_24247,N_21854,N_18805);
nor U24248 (N_24248,N_19537,N_21278);
xnor U24249 (N_24249,N_21451,N_19810);
nand U24250 (N_24250,N_21325,N_20747);
xor U24251 (N_24251,N_20081,N_20907);
nand U24252 (N_24252,N_21524,N_20953);
and U24253 (N_24253,N_20706,N_19525);
nand U24254 (N_24254,N_19051,N_20419);
or U24255 (N_24255,N_21022,N_20914);
nand U24256 (N_24256,N_20679,N_21193);
and U24257 (N_24257,N_19213,N_19953);
or U24258 (N_24258,N_19442,N_20045);
xor U24259 (N_24259,N_21425,N_18938);
nor U24260 (N_24260,N_20400,N_20593);
or U24261 (N_24261,N_18913,N_21163);
nor U24262 (N_24262,N_19818,N_20304);
or U24263 (N_24263,N_20665,N_20619);
or U24264 (N_24264,N_19314,N_20324);
nor U24265 (N_24265,N_19826,N_18938);
or U24266 (N_24266,N_19325,N_19572);
or U24267 (N_24267,N_21795,N_18957);
or U24268 (N_24268,N_20523,N_21726);
xor U24269 (N_24269,N_19547,N_20409);
and U24270 (N_24270,N_21108,N_21834);
and U24271 (N_24271,N_18882,N_20735);
nor U24272 (N_24272,N_20392,N_19214);
nand U24273 (N_24273,N_19206,N_20364);
and U24274 (N_24274,N_20958,N_19528);
nand U24275 (N_24275,N_20763,N_20490);
nor U24276 (N_24276,N_20047,N_20146);
and U24277 (N_24277,N_21497,N_19343);
nand U24278 (N_24278,N_19083,N_21144);
nor U24279 (N_24279,N_20780,N_20301);
and U24280 (N_24280,N_21573,N_21290);
and U24281 (N_24281,N_19811,N_20635);
and U24282 (N_24282,N_21187,N_19123);
nor U24283 (N_24283,N_20296,N_20300);
nor U24284 (N_24284,N_21280,N_19831);
or U24285 (N_24285,N_21560,N_19287);
nand U24286 (N_24286,N_18784,N_21729);
nand U24287 (N_24287,N_20065,N_21683);
nand U24288 (N_24288,N_19547,N_19681);
and U24289 (N_24289,N_20338,N_21556);
or U24290 (N_24290,N_21282,N_19888);
xnor U24291 (N_24291,N_18782,N_21432);
and U24292 (N_24292,N_18984,N_21052);
and U24293 (N_24293,N_19073,N_20393);
nor U24294 (N_24294,N_19111,N_19733);
nor U24295 (N_24295,N_19873,N_21692);
nor U24296 (N_24296,N_19907,N_20880);
nor U24297 (N_24297,N_19510,N_20801);
nor U24298 (N_24298,N_19905,N_20961);
or U24299 (N_24299,N_21416,N_19148);
nand U24300 (N_24300,N_19920,N_19731);
or U24301 (N_24301,N_20605,N_21557);
or U24302 (N_24302,N_20564,N_18760);
nor U24303 (N_24303,N_21755,N_19827);
or U24304 (N_24304,N_20576,N_20412);
nand U24305 (N_24305,N_21709,N_19304);
nand U24306 (N_24306,N_19749,N_19860);
or U24307 (N_24307,N_21682,N_19772);
and U24308 (N_24308,N_21396,N_19700);
nor U24309 (N_24309,N_20229,N_21686);
or U24310 (N_24310,N_20171,N_21745);
xor U24311 (N_24311,N_21410,N_21184);
xor U24312 (N_24312,N_21713,N_20613);
nand U24313 (N_24313,N_19504,N_18772);
or U24314 (N_24314,N_21749,N_20896);
or U24315 (N_24315,N_19140,N_20035);
nand U24316 (N_24316,N_19912,N_21246);
nand U24317 (N_24317,N_20716,N_21784);
nor U24318 (N_24318,N_18918,N_19910);
or U24319 (N_24319,N_20560,N_19097);
nand U24320 (N_24320,N_19167,N_21493);
or U24321 (N_24321,N_20116,N_19619);
or U24322 (N_24322,N_19450,N_20665);
nor U24323 (N_24323,N_19153,N_20992);
nor U24324 (N_24324,N_21207,N_20463);
xnor U24325 (N_24325,N_20612,N_21315);
nand U24326 (N_24326,N_19592,N_19953);
nand U24327 (N_24327,N_21724,N_19622);
nand U24328 (N_24328,N_19170,N_20457);
or U24329 (N_24329,N_19170,N_20802);
or U24330 (N_24330,N_19953,N_21845);
nor U24331 (N_24331,N_20802,N_19752);
or U24332 (N_24332,N_19175,N_20257);
nor U24333 (N_24333,N_19284,N_21596);
or U24334 (N_24334,N_21373,N_19962);
nor U24335 (N_24335,N_19184,N_20884);
nand U24336 (N_24336,N_20555,N_20969);
nand U24337 (N_24337,N_20775,N_20289);
and U24338 (N_24338,N_19962,N_21472);
nor U24339 (N_24339,N_20283,N_20026);
or U24340 (N_24340,N_19517,N_21011);
and U24341 (N_24341,N_21874,N_19672);
nor U24342 (N_24342,N_20155,N_19352);
or U24343 (N_24343,N_19041,N_19373);
nor U24344 (N_24344,N_20647,N_19663);
nor U24345 (N_24345,N_20047,N_21705);
xnor U24346 (N_24346,N_21704,N_21591);
xor U24347 (N_24347,N_20390,N_19349);
or U24348 (N_24348,N_19051,N_18869);
nor U24349 (N_24349,N_19030,N_20022);
and U24350 (N_24350,N_21716,N_21781);
nand U24351 (N_24351,N_18781,N_20357);
nand U24352 (N_24352,N_18802,N_20704);
nor U24353 (N_24353,N_19832,N_21364);
or U24354 (N_24354,N_20099,N_21643);
nand U24355 (N_24355,N_19507,N_20739);
nand U24356 (N_24356,N_20901,N_20289);
xnor U24357 (N_24357,N_19600,N_20010);
or U24358 (N_24358,N_18766,N_18847);
xor U24359 (N_24359,N_19449,N_19781);
and U24360 (N_24360,N_21268,N_18882);
or U24361 (N_24361,N_20874,N_19291);
nor U24362 (N_24362,N_18863,N_19335);
and U24363 (N_24363,N_19742,N_20434);
nand U24364 (N_24364,N_20903,N_19566);
nor U24365 (N_24365,N_20723,N_20919);
nand U24366 (N_24366,N_21395,N_19269);
or U24367 (N_24367,N_20136,N_20783);
nor U24368 (N_24368,N_20582,N_20171);
xnor U24369 (N_24369,N_20971,N_21346);
nor U24370 (N_24370,N_19796,N_21469);
xor U24371 (N_24371,N_20638,N_20995);
or U24372 (N_24372,N_20431,N_19325);
nand U24373 (N_24373,N_19138,N_19165);
nand U24374 (N_24374,N_18987,N_21334);
and U24375 (N_24375,N_19828,N_20006);
xnor U24376 (N_24376,N_18982,N_20543);
xor U24377 (N_24377,N_19343,N_21375);
xor U24378 (N_24378,N_20241,N_21218);
and U24379 (N_24379,N_21075,N_20159);
nand U24380 (N_24380,N_21496,N_19283);
nor U24381 (N_24381,N_20034,N_21228);
or U24382 (N_24382,N_18821,N_19751);
nand U24383 (N_24383,N_20092,N_20366);
nor U24384 (N_24384,N_20236,N_19912);
and U24385 (N_24385,N_20856,N_18925);
xnor U24386 (N_24386,N_20170,N_20652);
or U24387 (N_24387,N_21777,N_19691);
and U24388 (N_24388,N_21048,N_21288);
nand U24389 (N_24389,N_19190,N_19027);
or U24390 (N_24390,N_19211,N_19011);
xor U24391 (N_24391,N_19955,N_20456);
xor U24392 (N_24392,N_20265,N_20290);
xnor U24393 (N_24393,N_20565,N_21220);
nor U24394 (N_24394,N_21498,N_19320);
and U24395 (N_24395,N_19339,N_21591);
or U24396 (N_24396,N_21131,N_21106);
and U24397 (N_24397,N_20147,N_19171);
xor U24398 (N_24398,N_21266,N_21177);
nand U24399 (N_24399,N_19212,N_21507);
nand U24400 (N_24400,N_19948,N_20025);
and U24401 (N_24401,N_21067,N_20809);
or U24402 (N_24402,N_19534,N_21310);
or U24403 (N_24403,N_21270,N_21158);
and U24404 (N_24404,N_18961,N_18806);
or U24405 (N_24405,N_21790,N_21071);
or U24406 (N_24406,N_19237,N_20814);
or U24407 (N_24407,N_20223,N_19204);
nand U24408 (N_24408,N_19741,N_21516);
nand U24409 (N_24409,N_19361,N_20421);
nand U24410 (N_24410,N_21463,N_18796);
and U24411 (N_24411,N_20801,N_19553);
and U24412 (N_24412,N_20992,N_20704);
and U24413 (N_24413,N_19062,N_21093);
and U24414 (N_24414,N_20156,N_21521);
nor U24415 (N_24415,N_21246,N_19767);
nand U24416 (N_24416,N_18998,N_19475);
nand U24417 (N_24417,N_20510,N_19863);
or U24418 (N_24418,N_18776,N_20401);
nor U24419 (N_24419,N_20698,N_19210);
nor U24420 (N_24420,N_19684,N_19651);
and U24421 (N_24421,N_18872,N_20105);
nor U24422 (N_24422,N_19448,N_18913);
and U24423 (N_24423,N_19321,N_20866);
or U24424 (N_24424,N_20237,N_19263);
xor U24425 (N_24425,N_18815,N_19778);
or U24426 (N_24426,N_19045,N_21307);
nor U24427 (N_24427,N_21759,N_21164);
xor U24428 (N_24428,N_20097,N_20269);
nor U24429 (N_24429,N_21015,N_21356);
nor U24430 (N_24430,N_18929,N_19330);
and U24431 (N_24431,N_20650,N_19377);
or U24432 (N_24432,N_18794,N_19375);
nand U24433 (N_24433,N_20180,N_21220);
and U24434 (N_24434,N_21190,N_20454);
or U24435 (N_24435,N_19664,N_20610);
xor U24436 (N_24436,N_19142,N_20832);
and U24437 (N_24437,N_20206,N_21758);
nand U24438 (N_24438,N_19613,N_21207);
or U24439 (N_24439,N_20990,N_19018);
nand U24440 (N_24440,N_20313,N_20682);
or U24441 (N_24441,N_21700,N_20488);
nor U24442 (N_24442,N_21504,N_19150);
or U24443 (N_24443,N_19279,N_19221);
or U24444 (N_24444,N_21181,N_18979);
nor U24445 (N_24445,N_21139,N_21010);
nor U24446 (N_24446,N_20434,N_19737);
nor U24447 (N_24447,N_20709,N_18856);
nor U24448 (N_24448,N_20781,N_21099);
nand U24449 (N_24449,N_19800,N_21530);
and U24450 (N_24450,N_21622,N_19798);
and U24451 (N_24451,N_20131,N_20162);
or U24452 (N_24452,N_20465,N_18774);
nor U24453 (N_24453,N_20238,N_19746);
nor U24454 (N_24454,N_18935,N_19966);
nand U24455 (N_24455,N_20554,N_20546);
or U24456 (N_24456,N_21098,N_20742);
and U24457 (N_24457,N_21649,N_20320);
and U24458 (N_24458,N_19230,N_19590);
or U24459 (N_24459,N_19242,N_20889);
or U24460 (N_24460,N_20927,N_20153);
nor U24461 (N_24461,N_18915,N_19465);
nor U24462 (N_24462,N_21734,N_21036);
nor U24463 (N_24463,N_19824,N_20364);
or U24464 (N_24464,N_21814,N_21349);
and U24465 (N_24465,N_19188,N_21835);
or U24466 (N_24466,N_18903,N_20461);
nand U24467 (N_24467,N_21568,N_21504);
xor U24468 (N_24468,N_19525,N_20183);
and U24469 (N_24469,N_20381,N_21480);
or U24470 (N_24470,N_19707,N_21337);
or U24471 (N_24471,N_20261,N_20076);
nor U24472 (N_24472,N_19841,N_20824);
nor U24473 (N_24473,N_21430,N_21509);
or U24474 (N_24474,N_19733,N_19884);
nor U24475 (N_24475,N_21393,N_21757);
nand U24476 (N_24476,N_20027,N_20676);
nor U24477 (N_24477,N_19041,N_20390);
or U24478 (N_24478,N_21091,N_20546);
and U24479 (N_24479,N_19260,N_21241);
nor U24480 (N_24480,N_19649,N_21868);
and U24481 (N_24481,N_20073,N_19699);
nand U24482 (N_24482,N_21042,N_19434);
and U24483 (N_24483,N_19454,N_21066);
or U24484 (N_24484,N_18943,N_19955);
nor U24485 (N_24485,N_21441,N_20411);
nand U24486 (N_24486,N_18884,N_21803);
xor U24487 (N_24487,N_20908,N_19232);
nand U24488 (N_24488,N_21587,N_19812);
nor U24489 (N_24489,N_18793,N_20122);
or U24490 (N_24490,N_19927,N_18943);
nand U24491 (N_24491,N_21393,N_20396);
nor U24492 (N_24492,N_19794,N_20349);
nor U24493 (N_24493,N_19514,N_21335);
and U24494 (N_24494,N_19884,N_20699);
nand U24495 (N_24495,N_19087,N_19097);
nand U24496 (N_24496,N_19668,N_21062);
xor U24497 (N_24497,N_20448,N_18850);
nor U24498 (N_24498,N_20606,N_21586);
nor U24499 (N_24499,N_19093,N_21029);
nor U24500 (N_24500,N_19395,N_21481);
or U24501 (N_24501,N_19668,N_20693);
xor U24502 (N_24502,N_20781,N_19895);
nor U24503 (N_24503,N_21508,N_19207);
nand U24504 (N_24504,N_19194,N_20632);
and U24505 (N_24505,N_18780,N_20953);
xor U24506 (N_24506,N_20306,N_20894);
or U24507 (N_24507,N_21260,N_19927);
and U24508 (N_24508,N_20767,N_20855);
nand U24509 (N_24509,N_20028,N_21466);
nor U24510 (N_24510,N_21391,N_20034);
nor U24511 (N_24511,N_19728,N_21521);
nand U24512 (N_24512,N_19639,N_19177);
and U24513 (N_24513,N_21716,N_20005);
and U24514 (N_24514,N_20680,N_20634);
and U24515 (N_24515,N_21449,N_20863);
nor U24516 (N_24516,N_20858,N_20711);
nand U24517 (N_24517,N_21013,N_20115);
nand U24518 (N_24518,N_21074,N_19654);
nand U24519 (N_24519,N_19097,N_18992);
or U24520 (N_24520,N_20872,N_20403);
or U24521 (N_24521,N_21640,N_20290);
nor U24522 (N_24522,N_19439,N_19575);
or U24523 (N_24523,N_21794,N_19962);
nand U24524 (N_24524,N_20899,N_18814);
xor U24525 (N_24525,N_19343,N_20930);
and U24526 (N_24526,N_20633,N_19936);
nor U24527 (N_24527,N_20545,N_20832);
nor U24528 (N_24528,N_20759,N_20508);
and U24529 (N_24529,N_19888,N_19007);
or U24530 (N_24530,N_21185,N_19480);
or U24531 (N_24531,N_20281,N_21063);
nand U24532 (N_24532,N_19465,N_19012);
nand U24533 (N_24533,N_19800,N_20429);
nor U24534 (N_24534,N_21368,N_19631);
or U24535 (N_24535,N_20906,N_19156);
xnor U24536 (N_24536,N_20165,N_20404);
nor U24537 (N_24537,N_19425,N_18857);
or U24538 (N_24538,N_21288,N_21616);
or U24539 (N_24539,N_21355,N_19148);
and U24540 (N_24540,N_19842,N_20748);
xor U24541 (N_24541,N_20889,N_21134);
or U24542 (N_24542,N_20867,N_21155);
or U24543 (N_24543,N_18793,N_21629);
or U24544 (N_24544,N_21123,N_18975);
or U24545 (N_24545,N_19061,N_19007);
or U24546 (N_24546,N_20121,N_20359);
nand U24547 (N_24547,N_20830,N_19109);
nor U24548 (N_24548,N_18967,N_20178);
nand U24549 (N_24549,N_21035,N_21307);
and U24550 (N_24550,N_20045,N_21116);
xnor U24551 (N_24551,N_21836,N_20447);
or U24552 (N_24552,N_20844,N_21048);
and U24553 (N_24553,N_19995,N_19470);
or U24554 (N_24554,N_20782,N_20693);
nor U24555 (N_24555,N_19593,N_20971);
nor U24556 (N_24556,N_20429,N_20080);
and U24557 (N_24557,N_19044,N_18893);
and U24558 (N_24558,N_21833,N_20654);
and U24559 (N_24559,N_19007,N_18824);
nand U24560 (N_24560,N_19086,N_20813);
or U24561 (N_24561,N_20422,N_20618);
and U24562 (N_24562,N_21735,N_19275);
or U24563 (N_24563,N_19894,N_21340);
or U24564 (N_24564,N_20996,N_19318);
nor U24565 (N_24565,N_20508,N_20498);
nand U24566 (N_24566,N_19291,N_20807);
or U24567 (N_24567,N_19362,N_19317);
or U24568 (N_24568,N_21771,N_19012);
nand U24569 (N_24569,N_18946,N_20270);
nand U24570 (N_24570,N_18753,N_21849);
nand U24571 (N_24571,N_21601,N_20030);
nand U24572 (N_24572,N_21399,N_20507);
nand U24573 (N_24573,N_19098,N_18979);
xor U24574 (N_24574,N_20584,N_21546);
or U24575 (N_24575,N_19504,N_21632);
and U24576 (N_24576,N_18861,N_19098);
or U24577 (N_24577,N_20864,N_20223);
xor U24578 (N_24578,N_21117,N_18787);
nand U24579 (N_24579,N_20315,N_19441);
nor U24580 (N_24580,N_21606,N_19974);
nand U24581 (N_24581,N_21677,N_20100);
and U24582 (N_24582,N_21162,N_21769);
and U24583 (N_24583,N_20984,N_20141);
or U24584 (N_24584,N_20212,N_19061);
nand U24585 (N_24585,N_21381,N_18768);
or U24586 (N_24586,N_20768,N_19104);
or U24587 (N_24587,N_20729,N_19586);
and U24588 (N_24588,N_21587,N_20530);
and U24589 (N_24589,N_20421,N_21761);
nand U24590 (N_24590,N_21166,N_20658);
or U24591 (N_24591,N_19777,N_21657);
nor U24592 (N_24592,N_19919,N_21597);
nand U24593 (N_24593,N_21403,N_21300);
nand U24594 (N_24594,N_21038,N_21111);
and U24595 (N_24595,N_20484,N_19725);
or U24596 (N_24596,N_19089,N_20037);
nor U24597 (N_24597,N_18768,N_19324);
nand U24598 (N_24598,N_19626,N_19971);
nand U24599 (N_24599,N_21682,N_19096);
nand U24600 (N_24600,N_21608,N_20174);
and U24601 (N_24601,N_20848,N_19998);
and U24602 (N_24602,N_20264,N_19637);
nand U24603 (N_24603,N_20004,N_21576);
nand U24604 (N_24604,N_21017,N_20656);
xor U24605 (N_24605,N_19448,N_19293);
or U24606 (N_24606,N_19163,N_19356);
or U24607 (N_24607,N_19797,N_19683);
and U24608 (N_24608,N_19253,N_20871);
nor U24609 (N_24609,N_19588,N_20878);
and U24610 (N_24610,N_21009,N_21620);
xnor U24611 (N_24611,N_19002,N_20601);
nor U24612 (N_24612,N_20006,N_21657);
or U24613 (N_24613,N_21685,N_21392);
or U24614 (N_24614,N_20910,N_20106);
or U24615 (N_24615,N_20513,N_21611);
nor U24616 (N_24616,N_19820,N_20181);
and U24617 (N_24617,N_21547,N_18823);
and U24618 (N_24618,N_20485,N_20478);
and U24619 (N_24619,N_21764,N_21086);
and U24620 (N_24620,N_21568,N_21108);
xor U24621 (N_24621,N_21164,N_21634);
and U24622 (N_24622,N_20847,N_19182);
xor U24623 (N_24623,N_21481,N_18987);
nor U24624 (N_24624,N_20001,N_18836);
or U24625 (N_24625,N_20671,N_21466);
or U24626 (N_24626,N_21044,N_19137);
or U24627 (N_24627,N_20699,N_20189);
nor U24628 (N_24628,N_20778,N_21375);
xnor U24629 (N_24629,N_19255,N_19199);
and U24630 (N_24630,N_21859,N_20661);
or U24631 (N_24631,N_20638,N_20707);
or U24632 (N_24632,N_20308,N_20735);
nand U24633 (N_24633,N_20133,N_19676);
xnor U24634 (N_24634,N_21649,N_20247);
or U24635 (N_24635,N_20347,N_21859);
nand U24636 (N_24636,N_21325,N_19408);
nand U24637 (N_24637,N_19245,N_18880);
and U24638 (N_24638,N_19157,N_19860);
and U24639 (N_24639,N_20686,N_20915);
and U24640 (N_24640,N_21667,N_19515);
nor U24641 (N_24641,N_20834,N_19782);
nand U24642 (N_24642,N_21781,N_21082);
and U24643 (N_24643,N_21116,N_20778);
xor U24644 (N_24644,N_20599,N_20460);
xor U24645 (N_24645,N_19212,N_20024);
xor U24646 (N_24646,N_19499,N_19660);
xor U24647 (N_24647,N_19311,N_20536);
and U24648 (N_24648,N_20169,N_19231);
xnor U24649 (N_24649,N_21261,N_20793);
or U24650 (N_24650,N_20901,N_20836);
nand U24651 (N_24651,N_19860,N_21614);
or U24652 (N_24652,N_20461,N_19364);
nand U24653 (N_24653,N_21622,N_20836);
nand U24654 (N_24654,N_19279,N_19113);
or U24655 (N_24655,N_18780,N_21625);
and U24656 (N_24656,N_20235,N_20413);
nand U24657 (N_24657,N_20140,N_19528);
nand U24658 (N_24658,N_21737,N_18764);
and U24659 (N_24659,N_21538,N_21799);
nand U24660 (N_24660,N_20907,N_20137);
nor U24661 (N_24661,N_19975,N_20019);
nor U24662 (N_24662,N_20311,N_19727);
nor U24663 (N_24663,N_19937,N_21874);
or U24664 (N_24664,N_19593,N_19761);
xor U24665 (N_24665,N_20030,N_21647);
and U24666 (N_24666,N_21292,N_19246);
nor U24667 (N_24667,N_21324,N_19648);
xnor U24668 (N_24668,N_20915,N_19464);
nor U24669 (N_24669,N_21215,N_19825);
or U24670 (N_24670,N_20115,N_19236);
nand U24671 (N_24671,N_19111,N_19980);
and U24672 (N_24672,N_21147,N_19862);
or U24673 (N_24673,N_19466,N_20470);
nand U24674 (N_24674,N_21397,N_21867);
or U24675 (N_24675,N_19224,N_21114);
or U24676 (N_24676,N_21670,N_19777);
nor U24677 (N_24677,N_19521,N_20739);
or U24678 (N_24678,N_21215,N_19891);
nor U24679 (N_24679,N_19565,N_21129);
xnor U24680 (N_24680,N_21311,N_21073);
and U24681 (N_24681,N_21515,N_21355);
nand U24682 (N_24682,N_19063,N_19257);
xnor U24683 (N_24683,N_20229,N_21462);
nor U24684 (N_24684,N_21828,N_21854);
xnor U24685 (N_24685,N_20452,N_19987);
or U24686 (N_24686,N_20348,N_20953);
nor U24687 (N_24687,N_21377,N_20893);
nor U24688 (N_24688,N_21291,N_21202);
nor U24689 (N_24689,N_21250,N_21758);
or U24690 (N_24690,N_21858,N_19585);
nor U24691 (N_24691,N_21025,N_21652);
and U24692 (N_24692,N_20100,N_20166);
nand U24693 (N_24693,N_19679,N_21251);
xnor U24694 (N_24694,N_19401,N_21647);
or U24695 (N_24695,N_19567,N_21823);
or U24696 (N_24696,N_19113,N_21474);
nor U24697 (N_24697,N_19768,N_20418);
nor U24698 (N_24698,N_20119,N_20259);
and U24699 (N_24699,N_20714,N_21341);
or U24700 (N_24700,N_21809,N_20058);
nand U24701 (N_24701,N_20486,N_20358);
or U24702 (N_24702,N_19866,N_21589);
xor U24703 (N_24703,N_19237,N_21659);
or U24704 (N_24704,N_20189,N_19677);
or U24705 (N_24705,N_21250,N_21086);
nor U24706 (N_24706,N_20397,N_20748);
nor U24707 (N_24707,N_20252,N_20381);
nor U24708 (N_24708,N_19092,N_18847);
or U24709 (N_24709,N_19761,N_21685);
nand U24710 (N_24710,N_19690,N_20151);
nand U24711 (N_24711,N_19150,N_21402);
and U24712 (N_24712,N_19176,N_19036);
nand U24713 (N_24713,N_20786,N_18863);
nor U24714 (N_24714,N_19997,N_20405);
or U24715 (N_24715,N_21645,N_20575);
or U24716 (N_24716,N_20493,N_21768);
or U24717 (N_24717,N_20156,N_20784);
nand U24718 (N_24718,N_20084,N_20290);
xnor U24719 (N_24719,N_21095,N_21543);
nand U24720 (N_24720,N_21284,N_18902);
nor U24721 (N_24721,N_20945,N_20789);
nor U24722 (N_24722,N_21673,N_21451);
nand U24723 (N_24723,N_19637,N_20231);
nand U24724 (N_24724,N_21310,N_20354);
nand U24725 (N_24725,N_20063,N_19203);
and U24726 (N_24726,N_21715,N_19806);
and U24727 (N_24727,N_19119,N_21097);
nand U24728 (N_24728,N_19960,N_21547);
nor U24729 (N_24729,N_21536,N_21792);
nor U24730 (N_24730,N_21827,N_21850);
xor U24731 (N_24731,N_21037,N_20069);
or U24732 (N_24732,N_19455,N_21222);
nand U24733 (N_24733,N_18920,N_21794);
and U24734 (N_24734,N_20792,N_18951);
nor U24735 (N_24735,N_21157,N_21742);
nand U24736 (N_24736,N_19564,N_18897);
and U24737 (N_24737,N_21246,N_21745);
or U24738 (N_24738,N_21011,N_19365);
nor U24739 (N_24739,N_19961,N_21516);
or U24740 (N_24740,N_19577,N_20220);
xor U24741 (N_24741,N_20746,N_20779);
xnor U24742 (N_24742,N_19147,N_21108);
or U24743 (N_24743,N_20711,N_21624);
nor U24744 (N_24744,N_20406,N_18904);
nand U24745 (N_24745,N_21071,N_19299);
or U24746 (N_24746,N_20761,N_20195);
or U24747 (N_24747,N_20941,N_19395);
nand U24748 (N_24748,N_20694,N_20497);
nand U24749 (N_24749,N_21617,N_19182);
or U24750 (N_24750,N_19599,N_20384);
or U24751 (N_24751,N_21740,N_19705);
and U24752 (N_24752,N_20733,N_19869);
or U24753 (N_24753,N_21329,N_20242);
xor U24754 (N_24754,N_20282,N_21094);
and U24755 (N_24755,N_21788,N_20803);
or U24756 (N_24756,N_21173,N_21508);
and U24757 (N_24757,N_20067,N_20721);
or U24758 (N_24758,N_20213,N_19477);
or U24759 (N_24759,N_18990,N_20964);
nor U24760 (N_24760,N_20462,N_21317);
and U24761 (N_24761,N_18817,N_21802);
and U24762 (N_24762,N_19247,N_20275);
and U24763 (N_24763,N_20919,N_19581);
or U24764 (N_24764,N_21696,N_21016);
nor U24765 (N_24765,N_20438,N_19790);
nor U24766 (N_24766,N_21411,N_21220);
and U24767 (N_24767,N_18795,N_20116);
nor U24768 (N_24768,N_19545,N_21215);
or U24769 (N_24769,N_18974,N_21725);
or U24770 (N_24770,N_20444,N_19933);
nor U24771 (N_24771,N_21392,N_21458);
or U24772 (N_24772,N_21647,N_20043);
nor U24773 (N_24773,N_20140,N_20487);
nor U24774 (N_24774,N_20185,N_20806);
or U24775 (N_24775,N_20500,N_21235);
xnor U24776 (N_24776,N_21487,N_20494);
nand U24777 (N_24777,N_20934,N_19709);
nor U24778 (N_24778,N_20763,N_20772);
and U24779 (N_24779,N_21112,N_20372);
xor U24780 (N_24780,N_19416,N_21851);
and U24781 (N_24781,N_21035,N_19778);
xnor U24782 (N_24782,N_20315,N_21489);
nor U24783 (N_24783,N_20021,N_20441);
nor U24784 (N_24784,N_19999,N_20624);
nor U24785 (N_24785,N_19107,N_21653);
xor U24786 (N_24786,N_21587,N_18883);
and U24787 (N_24787,N_19206,N_20074);
and U24788 (N_24788,N_19103,N_21273);
nor U24789 (N_24789,N_21650,N_19025);
nor U24790 (N_24790,N_21443,N_20079);
nand U24791 (N_24791,N_20768,N_18974);
or U24792 (N_24792,N_21200,N_20506);
and U24793 (N_24793,N_21667,N_21040);
nand U24794 (N_24794,N_20288,N_19692);
and U24795 (N_24795,N_20197,N_19233);
nand U24796 (N_24796,N_21320,N_19790);
or U24797 (N_24797,N_20351,N_20575);
xnor U24798 (N_24798,N_21034,N_18766);
nand U24799 (N_24799,N_19363,N_20289);
or U24800 (N_24800,N_19905,N_20850);
and U24801 (N_24801,N_19977,N_21584);
and U24802 (N_24802,N_19195,N_21318);
or U24803 (N_24803,N_18890,N_19624);
and U24804 (N_24804,N_20214,N_21655);
and U24805 (N_24805,N_20948,N_19153);
nand U24806 (N_24806,N_19559,N_19580);
nand U24807 (N_24807,N_20382,N_20191);
or U24808 (N_24808,N_21136,N_20468);
nor U24809 (N_24809,N_21480,N_19984);
nand U24810 (N_24810,N_19099,N_18757);
or U24811 (N_24811,N_21305,N_19260);
nor U24812 (N_24812,N_21430,N_20283);
or U24813 (N_24813,N_19056,N_18791);
and U24814 (N_24814,N_18899,N_20957);
nor U24815 (N_24815,N_21077,N_21185);
nand U24816 (N_24816,N_19247,N_19424);
nor U24817 (N_24817,N_20442,N_18833);
nand U24818 (N_24818,N_19145,N_21045);
and U24819 (N_24819,N_19325,N_20263);
or U24820 (N_24820,N_20832,N_19411);
and U24821 (N_24821,N_19277,N_20027);
nor U24822 (N_24822,N_19446,N_20073);
and U24823 (N_24823,N_19672,N_21454);
or U24824 (N_24824,N_20212,N_20449);
xor U24825 (N_24825,N_21122,N_21852);
or U24826 (N_24826,N_21212,N_19019);
nor U24827 (N_24827,N_20181,N_19326);
and U24828 (N_24828,N_19117,N_20011);
or U24829 (N_24829,N_20788,N_20070);
or U24830 (N_24830,N_20468,N_20285);
nand U24831 (N_24831,N_20112,N_19226);
and U24832 (N_24832,N_18807,N_18887);
nand U24833 (N_24833,N_20430,N_19673);
nand U24834 (N_24834,N_18803,N_19922);
and U24835 (N_24835,N_20906,N_20377);
nand U24836 (N_24836,N_21268,N_20138);
or U24837 (N_24837,N_19848,N_21469);
nor U24838 (N_24838,N_19837,N_20325);
nor U24839 (N_24839,N_21125,N_19489);
nand U24840 (N_24840,N_20134,N_19479);
and U24841 (N_24841,N_21454,N_19669);
nor U24842 (N_24842,N_21087,N_19142);
nor U24843 (N_24843,N_19193,N_21046);
and U24844 (N_24844,N_21816,N_19390);
nor U24845 (N_24845,N_21015,N_19953);
xor U24846 (N_24846,N_20542,N_21416);
and U24847 (N_24847,N_20735,N_20300);
nand U24848 (N_24848,N_21472,N_21117);
nand U24849 (N_24849,N_19470,N_20179);
xor U24850 (N_24850,N_19323,N_19641);
or U24851 (N_24851,N_21486,N_20548);
or U24852 (N_24852,N_21546,N_21859);
nand U24853 (N_24853,N_21621,N_20923);
nand U24854 (N_24854,N_20938,N_19301);
nand U24855 (N_24855,N_20087,N_19375);
or U24856 (N_24856,N_18854,N_20324);
nor U24857 (N_24857,N_21551,N_19973);
xor U24858 (N_24858,N_19815,N_19969);
xor U24859 (N_24859,N_19075,N_21704);
nand U24860 (N_24860,N_21473,N_19517);
nand U24861 (N_24861,N_21498,N_20785);
or U24862 (N_24862,N_19684,N_19516);
nor U24863 (N_24863,N_20196,N_19818);
nor U24864 (N_24864,N_19168,N_20677);
or U24865 (N_24865,N_20817,N_19535);
or U24866 (N_24866,N_20400,N_20263);
nor U24867 (N_24867,N_21383,N_20027);
nor U24868 (N_24868,N_20380,N_19383);
nor U24869 (N_24869,N_19646,N_19446);
or U24870 (N_24870,N_20954,N_18914);
nand U24871 (N_24871,N_21530,N_20387);
nor U24872 (N_24872,N_20090,N_21706);
or U24873 (N_24873,N_19807,N_19333);
nor U24874 (N_24874,N_19782,N_19949);
nand U24875 (N_24875,N_19765,N_21482);
nor U24876 (N_24876,N_21325,N_20993);
and U24877 (N_24877,N_21854,N_19870);
nor U24878 (N_24878,N_20827,N_20612);
xor U24879 (N_24879,N_21607,N_19995);
nand U24880 (N_24880,N_19630,N_20670);
xor U24881 (N_24881,N_20294,N_21165);
nor U24882 (N_24882,N_19722,N_20212);
nand U24883 (N_24883,N_21279,N_19894);
or U24884 (N_24884,N_20731,N_21119);
nand U24885 (N_24885,N_21155,N_19603);
nor U24886 (N_24886,N_19930,N_19027);
or U24887 (N_24887,N_19525,N_21860);
nor U24888 (N_24888,N_20542,N_20697);
or U24889 (N_24889,N_18796,N_20953);
nor U24890 (N_24890,N_20662,N_19120);
or U24891 (N_24891,N_19606,N_20732);
and U24892 (N_24892,N_20297,N_19593);
or U24893 (N_24893,N_20603,N_19580);
nand U24894 (N_24894,N_18936,N_19041);
nand U24895 (N_24895,N_19467,N_20164);
nor U24896 (N_24896,N_20792,N_20123);
or U24897 (N_24897,N_20908,N_19064);
or U24898 (N_24898,N_18912,N_19021);
nor U24899 (N_24899,N_20263,N_20095);
or U24900 (N_24900,N_21156,N_19897);
and U24901 (N_24901,N_19581,N_21173);
nand U24902 (N_24902,N_19806,N_20080);
nand U24903 (N_24903,N_20904,N_20918);
and U24904 (N_24904,N_21295,N_19573);
nand U24905 (N_24905,N_20660,N_20969);
or U24906 (N_24906,N_18775,N_19810);
nor U24907 (N_24907,N_19939,N_19959);
nand U24908 (N_24908,N_19896,N_20487);
and U24909 (N_24909,N_21232,N_18940);
nand U24910 (N_24910,N_21154,N_20270);
nor U24911 (N_24911,N_18812,N_19140);
nor U24912 (N_24912,N_20023,N_20359);
nand U24913 (N_24913,N_19229,N_21177);
xnor U24914 (N_24914,N_19536,N_20972);
and U24915 (N_24915,N_21453,N_21775);
nor U24916 (N_24916,N_20395,N_21120);
nor U24917 (N_24917,N_19140,N_21336);
and U24918 (N_24918,N_19710,N_19725);
or U24919 (N_24919,N_21443,N_21364);
nand U24920 (N_24920,N_21468,N_21534);
or U24921 (N_24921,N_20348,N_19851);
nand U24922 (N_24922,N_20322,N_19930);
nand U24923 (N_24923,N_21765,N_20549);
xnor U24924 (N_24924,N_19844,N_20112);
or U24925 (N_24925,N_20277,N_19587);
and U24926 (N_24926,N_21464,N_18945);
and U24927 (N_24927,N_20179,N_21107);
nor U24928 (N_24928,N_21628,N_20570);
or U24929 (N_24929,N_20588,N_19048);
or U24930 (N_24930,N_20685,N_19937);
or U24931 (N_24931,N_20438,N_19331);
nor U24932 (N_24932,N_20334,N_20550);
and U24933 (N_24933,N_20677,N_21549);
and U24934 (N_24934,N_20204,N_19633);
nand U24935 (N_24935,N_21548,N_19090);
nand U24936 (N_24936,N_20896,N_20494);
nor U24937 (N_24937,N_19799,N_20677);
xnor U24938 (N_24938,N_19084,N_21634);
nor U24939 (N_24939,N_19265,N_21371);
nand U24940 (N_24940,N_19783,N_18795);
nand U24941 (N_24941,N_19459,N_19332);
nor U24942 (N_24942,N_19398,N_21532);
nand U24943 (N_24943,N_21124,N_19552);
nor U24944 (N_24944,N_18864,N_21522);
xnor U24945 (N_24945,N_19038,N_19557);
nor U24946 (N_24946,N_19703,N_19281);
nand U24947 (N_24947,N_19002,N_20453);
and U24948 (N_24948,N_18767,N_21120);
nor U24949 (N_24949,N_19777,N_21015);
and U24950 (N_24950,N_19518,N_20458);
xor U24951 (N_24951,N_19015,N_21522);
nor U24952 (N_24952,N_19792,N_19332);
and U24953 (N_24953,N_19758,N_20536);
or U24954 (N_24954,N_20673,N_19698);
xnor U24955 (N_24955,N_20786,N_18956);
or U24956 (N_24956,N_20853,N_21126);
nor U24957 (N_24957,N_20754,N_21411);
and U24958 (N_24958,N_19935,N_20368);
and U24959 (N_24959,N_19753,N_19486);
and U24960 (N_24960,N_21739,N_20673);
nor U24961 (N_24961,N_20991,N_18890);
or U24962 (N_24962,N_19168,N_19160);
or U24963 (N_24963,N_20765,N_20481);
nand U24964 (N_24964,N_21129,N_19693);
and U24965 (N_24965,N_20110,N_19174);
or U24966 (N_24966,N_20510,N_20558);
and U24967 (N_24967,N_20946,N_21242);
nand U24968 (N_24968,N_18806,N_20183);
or U24969 (N_24969,N_20551,N_19587);
nor U24970 (N_24970,N_21069,N_19856);
nor U24971 (N_24971,N_21783,N_21585);
or U24972 (N_24972,N_20131,N_20251);
or U24973 (N_24973,N_19411,N_19352);
xnor U24974 (N_24974,N_21113,N_20306);
and U24975 (N_24975,N_20309,N_21660);
or U24976 (N_24976,N_20570,N_18844);
or U24977 (N_24977,N_20505,N_19791);
xor U24978 (N_24978,N_20174,N_19564);
nor U24979 (N_24979,N_19056,N_21424);
and U24980 (N_24980,N_21746,N_21267);
nor U24981 (N_24981,N_19164,N_19521);
and U24982 (N_24982,N_21575,N_19608);
and U24983 (N_24983,N_20158,N_21808);
and U24984 (N_24984,N_21406,N_21703);
nand U24985 (N_24985,N_19546,N_19406);
nand U24986 (N_24986,N_20169,N_20892);
nand U24987 (N_24987,N_20657,N_18998);
nand U24988 (N_24988,N_19459,N_20679);
or U24989 (N_24989,N_20827,N_20561);
xnor U24990 (N_24990,N_21126,N_19154);
nor U24991 (N_24991,N_20653,N_19031);
nand U24992 (N_24992,N_21729,N_21322);
nor U24993 (N_24993,N_18869,N_21656);
nor U24994 (N_24994,N_21158,N_20709);
nor U24995 (N_24995,N_19730,N_21000);
xor U24996 (N_24996,N_20839,N_19052);
nand U24997 (N_24997,N_20387,N_19600);
or U24998 (N_24998,N_19770,N_19553);
and U24999 (N_24999,N_19600,N_20506);
and UO_0 (O_0,N_24564,N_23580);
xnor UO_1 (O_1,N_23205,N_23500);
and UO_2 (O_2,N_21973,N_22318);
or UO_3 (O_3,N_24774,N_22872);
and UO_4 (O_4,N_24841,N_24311);
nor UO_5 (O_5,N_22635,N_24281);
nand UO_6 (O_6,N_22191,N_24130);
nor UO_7 (O_7,N_24648,N_22567);
xor UO_8 (O_8,N_22895,N_24953);
nand UO_9 (O_9,N_22585,N_24951);
and UO_10 (O_10,N_23346,N_22480);
and UO_11 (O_11,N_24116,N_22432);
or UO_12 (O_12,N_22897,N_24520);
or UO_13 (O_13,N_23540,N_21928);
xor UO_14 (O_14,N_22364,N_23495);
nand UO_15 (O_15,N_24965,N_23379);
nand UO_16 (O_16,N_23093,N_24274);
and UO_17 (O_17,N_23323,N_24479);
nor UO_18 (O_18,N_23218,N_24940);
and UO_19 (O_19,N_23034,N_22050);
or UO_20 (O_20,N_22173,N_24844);
nand UO_21 (O_21,N_24155,N_24166);
and UO_22 (O_22,N_22052,N_23698);
nand UO_23 (O_23,N_23526,N_23122);
nand UO_24 (O_24,N_23378,N_22516);
nor UO_25 (O_25,N_22892,N_23282);
and UO_26 (O_26,N_23940,N_24602);
xnor UO_27 (O_27,N_22581,N_22182);
nand UO_28 (O_28,N_24179,N_23476);
nor UO_29 (O_29,N_24044,N_23833);
and UO_30 (O_30,N_22643,N_22808);
and UO_31 (O_31,N_21983,N_24813);
xor UO_32 (O_32,N_24859,N_24535);
nand UO_33 (O_33,N_22231,N_22030);
nand UO_34 (O_34,N_24306,N_23200);
nand UO_35 (O_35,N_23679,N_22865);
and UO_36 (O_36,N_23197,N_22188);
and UO_37 (O_37,N_22984,N_23621);
or UO_38 (O_38,N_22909,N_23689);
or UO_39 (O_39,N_22092,N_21945);
and UO_40 (O_40,N_24241,N_22180);
nor UO_41 (O_41,N_23944,N_22309);
xor UO_42 (O_42,N_23842,N_22398);
nor UO_43 (O_43,N_24639,N_22236);
or UO_44 (O_44,N_22438,N_23141);
nand UO_45 (O_45,N_22484,N_22389);
and UO_46 (O_46,N_24038,N_24443);
or UO_47 (O_47,N_22574,N_22443);
and UO_48 (O_48,N_24878,N_24171);
or UO_49 (O_49,N_24504,N_23954);
nand UO_50 (O_50,N_22982,N_23193);
nor UO_51 (O_51,N_24925,N_24091);
xnor UO_52 (O_52,N_22072,N_24012);
nor UO_53 (O_53,N_23752,N_23992);
or UO_54 (O_54,N_24890,N_24789);
nand UO_55 (O_55,N_22562,N_23489);
nor UO_56 (O_56,N_24750,N_23825);
nand UO_57 (O_57,N_24669,N_24384);
nand UO_58 (O_58,N_23174,N_24194);
nand UO_59 (O_59,N_24661,N_23538);
and UO_60 (O_60,N_22492,N_22442);
or UO_61 (O_61,N_23380,N_23979);
nand UO_62 (O_62,N_22810,N_23359);
nor UO_63 (O_63,N_24884,N_22434);
nor UO_64 (O_64,N_23659,N_23397);
xor UO_65 (O_65,N_22162,N_23294);
and UO_66 (O_66,N_24956,N_24411);
nor UO_67 (O_67,N_22864,N_23901);
xnor UO_68 (O_68,N_23360,N_24374);
or UO_69 (O_69,N_24278,N_22007);
and UO_70 (O_70,N_23103,N_23573);
or UO_71 (O_71,N_24621,N_24335);
nor UO_72 (O_72,N_24704,N_24871);
or UO_73 (O_73,N_24518,N_23233);
nand UO_74 (O_74,N_24713,N_24201);
nand UO_75 (O_75,N_24214,N_24578);
nand UO_76 (O_76,N_24096,N_24053);
nor UO_77 (O_77,N_22147,N_23860);
or UO_78 (O_78,N_22378,N_24132);
and UO_79 (O_79,N_22120,N_22408);
nand UO_80 (O_80,N_24126,N_24446);
and UO_81 (O_81,N_24711,N_22557);
nand UO_82 (O_82,N_22177,N_23232);
or UO_83 (O_83,N_23691,N_24316);
or UO_84 (O_84,N_23681,N_22522);
and UO_85 (O_85,N_24865,N_23337);
nor UO_86 (O_86,N_23613,N_24204);
and UO_87 (O_87,N_22747,N_21905);
or UO_88 (O_88,N_23917,N_23432);
nor UO_89 (O_89,N_23016,N_24500);
or UO_90 (O_90,N_23366,N_23809);
and UO_91 (O_91,N_23302,N_24935);
nand UO_92 (O_92,N_24183,N_23182);
and UO_93 (O_93,N_23334,N_22705);
or UO_94 (O_94,N_24366,N_23095);
and UO_95 (O_95,N_22657,N_22680);
or UO_96 (O_96,N_22765,N_23411);
and UO_97 (O_97,N_22273,N_23822);
nand UO_98 (O_98,N_22812,N_22337);
and UO_99 (O_99,N_22326,N_23038);
or UO_100 (O_100,N_24026,N_22329);
nor UO_101 (O_101,N_24560,N_24418);
nand UO_102 (O_102,N_23968,N_21916);
and UO_103 (O_103,N_24459,N_24478);
or UO_104 (O_104,N_22768,N_23853);
nor UO_105 (O_105,N_22366,N_23999);
nand UO_106 (O_106,N_22740,N_22627);
nor UO_107 (O_107,N_22604,N_23738);
nor UO_108 (O_108,N_22234,N_23271);
nand UO_109 (O_109,N_23072,N_22928);
or UO_110 (O_110,N_22429,N_22418);
or UO_111 (O_111,N_24185,N_22140);
nand UO_112 (O_112,N_24815,N_23053);
and UO_113 (O_113,N_22462,N_23322);
nor UO_114 (O_114,N_23123,N_24991);
and UO_115 (O_115,N_23648,N_22658);
nor UO_116 (O_116,N_24203,N_23471);
or UO_117 (O_117,N_23354,N_24162);
nor UO_118 (O_118,N_24315,N_24002);
xor UO_119 (O_119,N_24681,N_22776);
or UO_120 (O_120,N_23768,N_21990);
or UO_121 (O_121,N_22850,N_23417);
nor UO_122 (O_122,N_22965,N_24133);
nand UO_123 (O_123,N_23481,N_22158);
or UO_124 (O_124,N_21965,N_24342);
and UO_125 (O_125,N_22525,N_23245);
nand UO_126 (O_126,N_23907,N_24557);
or UO_127 (O_127,N_22206,N_22750);
or UO_128 (O_128,N_22951,N_22226);
nor UO_129 (O_129,N_24405,N_22196);
and UO_130 (O_130,N_24348,N_23001);
and UO_131 (O_131,N_23957,N_22683);
and UO_132 (O_132,N_23563,N_23591);
nand UO_133 (O_133,N_23514,N_24656);
and UO_134 (O_134,N_22999,N_22457);
or UO_135 (O_135,N_23083,N_23480);
and UO_136 (O_136,N_22430,N_24093);
nand UO_137 (O_137,N_22908,N_22717);
nand UO_138 (O_138,N_23088,N_22261);
or UO_139 (O_139,N_24157,N_22542);
nor UO_140 (O_140,N_22874,N_23823);
and UO_141 (O_141,N_22762,N_21920);
xor UO_142 (O_142,N_24483,N_23544);
nor UO_143 (O_143,N_22724,N_24165);
and UO_144 (O_144,N_23576,N_23382);
nor UO_145 (O_145,N_22844,N_23438);
and UO_146 (O_146,N_22617,N_21909);
or UO_147 (O_147,N_23778,N_22912);
nor UO_148 (O_148,N_23509,N_24037);
or UO_149 (O_149,N_22757,N_24706);
nand UO_150 (O_150,N_22902,N_23423);
or UO_151 (O_151,N_24234,N_23325);
or UO_152 (O_152,N_23238,N_24533);
nor UO_153 (O_153,N_22539,N_24187);
and UO_154 (O_154,N_24303,N_24523);
or UO_155 (O_155,N_24840,N_23781);
nor UO_156 (O_156,N_22433,N_23894);
nor UO_157 (O_157,N_24473,N_21879);
nand UO_158 (O_158,N_24728,N_22898);
or UO_159 (O_159,N_21885,N_24738);
or UO_160 (O_160,N_23064,N_23059);
or UO_161 (O_161,N_23821,N_22699);
nand UO_162 (O_162,N_22978,N_24539);
or UO_163 (O_163,N_23473,N_24904);
nand UO_164 (O_164,N_22666,N_24690);
nand UO_165 (O_165,N_22216,N_21966);
nor UO_166 (O_166,N_23706,N_24702);
nand UO_167 (O_167,N_22736,N_22256);
nor UO_168 (O_168,N_24849,N_22315);
xor UO_169 (O_169,N_23726,N_23270);
or UO_170 (O_170,N_24931,N_22953);
or UO_171 (O_171,N_23863,N_24510);
and UO_172 (O_172,N_24231,N_24784);
nor UO_173 (O_173,N_23080,N_22858);
or UO_174 (O_174,N_24779,N_22956);
nand UO_175 (O_175,N_23865,N_22424);
nor UO_176 (O_176,N_24642,N_23568);
or UO_177 (O_177,N_22533,N_24016);
or UO_178 (O_178,N_23522,N_22820);
and UO_179 (O_179,N_24667,N_24822);
xor UO_180 (O_180,N_24641,N_22126);
or UO_181 (O_181,N_24470,N_23994);
nor UO_182 (O_182,N_23923,N_22100);
and UO_183 (O_183,N_23654,N_22787);
nand UO_184 (O_184,N_21956,N_23602);
and UO_185 (O_185,N_23880,N_23463);
nand UO_186 (O_186,N_24022,N_23479);
xnor UO_187 (O_187,N_24593,N_23040);
nor UO_188 (O_188,N_22145,N_23265);
nand UO_189 (O_189,N_22625,N_22381);
xnor UO_190 (O_190,N_24679,N_24146);
or UO_191 (O_191,N_24371,N_23344);
or UO_192 (O_192,N_22425,N_22107);
or UO_193 (O_193,N_24762,N_22507);
nor UO_194 (O_194,N_23523,N_24379);
nand UO_195 (O_195,N_24363,N_24174);
nand UO_196 (O_196,N_24970,N_23100);
nand UO_197 (O_197,N_23737,N_24867);
or UO_198 (O_198,N_24168,N_24806);
nor UO_199 (O_199,N_22062,N_22132);
nand UO_200 (O_200,N_23876,N_23277);
and UO_201 (O_201,N_22804,N_23457);
xor UO_202 (O_202,N_21919,N_21995);
nand UO_203 (O_203,N_24000,N_23308);
nand UO_204 (O_204,N_23811,N_21932);
nand UO_205 (O_205,N_24513,N_22554);
or UO_206 (O_206,N_22654,N_23700);
or UO_207 (O_207,N_24190,N_24941);
and UO_208 (O_208,N_23623,N_24885);
nand UO_209 (O_209,N_24527,N_22043);
and UO_210 (O_210,N_22940,N_23560);
and UO_211 (O_211,N_22482,N_23600);
and UO_212 (O_212,N_24647,N_24979);
or UO_213 (O_213,N_23009,N_24652);
or UO_214 (O_214,N_22000,N_22346);
nor UO_215 (O_215,N_24524,N_22916);
and UO_216 (O_216,N_24842,N_22644);
nor UO_217 (O_217,N_22726,N_22678);
and UO_218 (O_218,N_24192,N_23369);
xnor UO_219 (O_219,N_22606,N_22921);
and UO_220 (O_220,N_24958,N_24402);
nor UO_221 (O_221,N_23903,N_24975);
nand UO_222 (O_222,N_24660,N_22298);
or UO_223 (O_223,N_24553,N_23662);
nor UO_224 (O_224,N_23456,N_23579);
nor UO_225 (O_225,N_24501,N_22568);
and UO_226 (O_226,N_23467,N_23029);
nor UO_227 (O_227,N_23742,N_23686);
nand UO_228 (O_228,N_21876,N_22607);
nand UO_229 (O_229,N_23176,N_23864);
and UO_230 (O_230,N_22624,N_22278);
xnor UO_231 (O_231,N_24901,N_22818);
and UO_232 (O_232,N_22690,N_23594);
nor UO_233 (O_233,N_24356,N_24177);
and UO_234 (O_234,N_22466,N_22615);
nand UO_235 (O_235,N_23527,N_24139);
nand UO_236 (O_236,N_22105,N_22501);
nor UO_237 (O_237,N_23057,N_24296);
and UO_238 (O_238,N_23584,N_22193);
nand UO_239 (O_239,N_22536,N_23446);
and UO_240 (O_240,N_24571,N_22521);
or UO_241 (O_241,N_24228,N_23065);
and UO_242 (O_242,N_24034,N_23785);
nand UO_243 (O_243,N_22045,N_23291);
nor UO_244 (O_244,N_22491,N_22927);
or UO_245 (O_245,N_23362,N_24989);
and UO_246 (O_246,N_22409,N_24930);
nand UO_247 (O_247,N_24294,N_24905);
or UO_248 (O_248,N_24515,N_22697);
nor UO_249 (O_249,N_23272,N_23985);
nand UO_250 (O_250,N_22569,N_24614);
and UO_251 (O_251,N_22709,N_23950);
and UO_252 (O_252,N_24927,N_24236);
or UO_253 (O_253,N_22384,N_23442);
or UO_254 (O_254,N_23076,N_22753);
nor UO_255 (O_255,N_23771,N_23827);
nand UO_256 (O_256,N_24361,N_22650);
and UO_257 (O_257,N_23299,N_24343);
or UO_258 (O_258,N_23020,N_24039);
nand UO_259 (O_259,N_24328,N_23050);
or UO_260 (O_260,N_24532,N_24007);
or UO_261 (O_261,N_23530,N_22171);
and UO_262 (O_262,N_24154,N_23775);
nor UO_263 (O_263,N_22413,N_23431);
or UO_264 (O_264,N_24707,N_23084);
nand UO_265 (O_265,N_24301,N_24549);
nand UO_266 (O_266,N_22013,N_24655);
nor UO_267 (O_267,N_22512,N_24529);
or UO_268 (O_268,N_24734,N_24065);
or UO_269 (O_269,N_22485,N_23424);
nand UO_270 (O_270,N_23967,N_22215);
or UO_271 (O_271,N_23339,N_22117);
nand UO_272 (O_272,N_24741,N_21944);
nand UO_273 (O_273,N_22478,N_24757);
nand UO_274 (O_274,N_23228,N_24934);
and UO_275 (O_275,N_22859,N_23307);
nand UO_276 (O_276,N_22879,N_22086);
and UO_277 (O_277,N_23725,N_22547);
or UO_278 (O_278,N_24386,N_23906);
nand UO_279 (O_279,N_24577,N_23843);
nand UO_280 (O_280,N_24993,N_23871);
and UO_281 (O_281,N_24684,N_22260);
nor UO_282 (O_282,N_22189,N_24280);
or UO_283 (O_283,N_22125,N_22556);
and UO_284 (O_284,N_24814,N_22041);
nor UO_285 (O_285,N_23212,N_22875);
and UO_286 (O_286,N_24926,N_22802);
nand UO_287 (O_287,N_24612,N_23414);
or UO_288 (O_288,N_22842,N_23230);
or UO_289 (O_289,N_22934,N_24457);
nor UO_290 (O_290,N_22047,N_24454);
and UO_291 (O_291,N_21962,N_22590);
nand UO_292 (O_292,N_24898,N_22632);
nand UO_293 (O_293,N_24059,N_23969);
or UO_294 (O_294,N_24914,N_22620);
xnor UO_295 (O_295,N_23902,N_22407);
and UO_296 (O_296,N_23852,N_24864);
nand UO_297 (O_297,N_22944,N_23834);
nor UO_298 (O_298,N_23795,N_24505);
or UO_299 (O_299,N_24997,N_24696);
nand UO_300 (O_300,N_21948,N_23023);
nand UO_301 (O_301,N_23484,N_24887);
nor UO_302 (O_302,N_23956,N_23383);
or UO_303 (O_303,N_22969,N_24739);
nor UO_304 (O_304,N_23996,N_23861);
or UO_305 (O_305,N_23543,N_24138);
and UO_306 (O_306,N_24309,N_23598);
nand UO_307 (O_307,N_23502,N_22955);
and UO_308 (O_308,N_23914,N_22852);
nor UO_309 (O_309,N_24327,N_24131);
nand UO_310 (O_310,N_24731,N_21934);
nand UO_311 (O_311,N_21964,N_24438);
nor UO_312 (O_312,N_24793,N_22076);
and UO_313 (O_313,N_23089,N_24486);
nand UO_314 (O_314,N_23435,N_22689);
nand UO_315 (O_315,N_22185,N_24536);
nor UO_316 (O_316,N_23046,N_23104);
or UO_317 (O_317,N_23296,N_22653);
nand UO_318 (O_318,N_22376,N_23352);
xnor UO_319 (O_319,N_22130,N_23234);
nand UO_320 (O_320,N_24896,N_23485);
nand UO_321 (O_321,N_23276,N_23891);
and UO_322 (O_322,N_23552,N_22400);
nor UO_323 (O_323,N_24765,N_24752);
nand UO_324 (O_324,N_23711,N_22454);
nand UO_325 (O_325,N_22741,N_23330);
and UO_326 (O_326,N_23697,N_22305);
xor UO_327 (O_327,N_22455,N_23603);
and UO_328 (O_328,N_24142,N_24047);
nand UO_329 (O_329,N_23257,N_23358);
or UO_330 (O_330,N_23557,N_23942);
or UO_331 (O_331,N_24125,N_24419);
nand UO_332 (O_332,N_24066,N_24819);
nor UO_333 (O_333,N_24409,N_22073);
or UO_334 (O_334,N_23610,N_24899);
nand UO_335 (O_335,N_23764,N_23839);
xnor UO_336 (O_336,N_24633,N_23281);
nor UO_337 (O_337,N_23086,N_24922);
and UO_338 (O_338,N_24484,N_23644);
nand UO_339 (O_339,N_22899,N_22770);
or UO_340 (O_340,N_24238,N_24101);
nor UO_341 (O_341,N_22113,N_23963);
nor UO_342 (O_342,N_24924,N_23805);
nand UO_343 (O_343,N_23889,N_24703);
nor UO_344 (O_344,N_24268,N_24095);
or UO_345 (O_345,N_22958,N_24746);
nor UO_346 (O_346,N_23769,N_22352);
and UO_347 (O_347,N_24950,N_21969);
nor UO_348 (O_348,N_24198,N_22813);
nand UO_349 (O_349,N_24364,N_23614);
nor UO_350 (O_350,N_22319,N_22532);
or UO_351 (O_351,N_22719,N_24556);
or UO_352 (O_352,N_24099,N_24148);
nand UO_353 (O_353,N_22194,N_24476);
and UO_354 (O_354,N_23849,N_22936);
or UO_355 (O_355,N_24029,N_23581);
nor UO_356 (O_356,N_22519,N_24832);
nor UO_357 (O_357,N_24243,N_22333);
nor UO_358 (O_358,N_24251,N_23246);
nand UO_359 (O_359,N_24824,N_22098);
or UO_360 (O_360,N_22289,N_23306);
and UO_361 (O_361,N_23845,N_24427);
and UO_362 (O_362,N_23721,N_23753);
or UO_363 (O_363,N_24623,N_23041);
or UO_364 (O_364,N_23135,N_24253);
or UO_365 (O_365,N_23735,N_23178);
xnor UO_366 (O_366,N_23810,N_23702);
or UO_367 (O_367,N_22471,N_24981);
nand UO_368 (O_368,N_23247,N_22027);
nor UO_369 (O_369,N_22168,N_23608);
and UO_370 (O_370,N_24978,N_22028);
or UO_371 (O_371,N_22637,N_23788);
nand UO_372 (O_372,N_24213,N_23412);
and UO_373 (O_373,N_23625,N_23260);
nor UO_374 (O_374,N_23553,N_23287);
and UO_375 (O_375,N_23129,N_23762);
nand UO_376 (O_376,N_22332,N_24413);
and UO_377 (O_377,N_24319,N_24465);
nor UO_378 (O_378,N_23813,N_24879);
nor UO_379 (O_379,N_23012,N_22561);
and UO_380 (O_380,N_24735,N_23073);
and UO_381 (O_381,N_21978,N_21884);
nor UO_382 (O_382,N_22947,N_22174);
nor UO_383 (O_383,N_22641,N_24389);
nor UO_384 (O_384,N_23459,N_24946);
and UO_385 (O_385,N_23590,N_24452);
and UO_386 (O_386,N_24163,N_23096);
and UO_387 (O_387,N_22394,N_24225);
and UO_388 (O_388,N_22629,N_22553);
and UO_389 (O_389,N_22016,N_23637);
nand UO_390 (O_390,N_24610,N_23286);
xor UO_391 (O_391,N_23405,N_22887);
and UO_392 (O_392,N_24908,N_23973);
nand UO_393 (O_393,N_24267,N_21913);
or UO_394 (O_394,N_23003,N_22684);
or UO_395 (O_395,N_22870,N_22488);
and UO_396 (O_396,N_22592,N_21899);
xor UO_397 (O_397,N_21963,N_24748);
or UO_398 (O_398,N_22550,N_22386);
nand UO_399 (O_399,N_24687,N_24954);
and UO_400 (O_400,N_23011,N_22775);
nor UO_401 (O_401,N_22640,N_23355);
nand UO_402 (O_402,N_24011,N_22692);
and UO_403 (O_403,N_22816,N_23545);
nand UO_404 (O_404,N_24709,N_22150);
nor UO_405 (O_405,N_23960,N_22758);
xnor UO_406 (O_406,N_24257,N_22192);
and UO_407 (O_407,N_23541,N_23517);
nand UO_408 (O_408,N_23367,N_23268);
xnor UO_409 (O_409,N_24569,N_22826);
nand UO_410 (O_410,N_24522,N_22819);
and UO_411 (O_411,N_24851,N_24299);
nor UO_412 (O_412,N_22919,N_22610);
nand UO_413 (O_413,N_22970,N_22118);
xnor UO_414 (O_414,N_22505,N_24786);
nor UO_415 (O_415,N_22367,N_23665);
and UO_416 (O_416,N_24700,N_22451);
and UO_417 (O_417,N_23211,N_24780);
nand UO_418 (O_418,N_21971,N_23874);
xnor UO_419 (O_419,N_24902,N_22328);
xnor UO_420 (O_420,N_24440,N_22973);
nand UO_421 (O_421,N_22359,N_24086);
nand UO_422 (O_422,N_22530,N_22221);
and UO_423 (O_423,N_24193,N_24329);
or UO_424 (O_424,N_23381,N_24423);
nand UO_425 (O_425,N_22166,N_23185);
xnor UO_426 (O_426,N_23534,N_23207);
nor UO_427 (O_427,N_22004,N_23928);
nor UO_428 (O_428,N_23519,N_23696);
or UO_429 (O_429,N_22044,N_23628);
or UO_430 (O_430,N_23645,N_24158);
or UO_431 (O_431,N_21904,N_22402);
xor UO_432 (O_432,N_23067,N_23748);
nor UO_433 (O_433,N_24377,N_23289);
nand UO_434 (O_434,N_21997,N_23136);
xnor UO_435 (O_435,N_22760,N_23121);
nor UO_436 (O_436,N_24994,N_22152);
and UO_437 (O_437,N_24891,N_22184);
and UO_438 (O_438,N_24874,N_23856);
nor UO_439 (O_439,N_23159,N_22931);
nand UO_440 (O_440,N_24083,N_22972);
and UO_441 (O_441,N_23342,N_21999);
nand UO_442 (O_442,N_24369,N_23714);
and UO_443 (O_443,N_23828,N_24692);
nor UO_444 (O_444,N_24759,N_23508);
nor UO_445 (O_445,N_23324,N_24792);
or UO_446 (O_446,N_23014,N_24937);
nand UO_447 (O_447,N_24128,N_22222);
nand UO_448 (O_448,N_22938,N_22849);
or UO_449 (O_449,N_23437,N_22253);
xnor UO_450 (O_450,N_23137,N_23044);
xnor UO_451 (O_451,N_23806,N_23173);
nand UO_452 (O_452,N_24949,N_23784);
xnor UO_453 (O_453,N_23847,N_22911);
nor UO_454 (O_454,N_24071,N_23450);
nor UO_455 (O_455,N_23461,N_22963);
or UO_456 (O_456,N_23496,N_22576);
and UO_457 (O_457,N_22081,N_23814);
or UO_458 (O_458,N_24474,N_22672);
or UO_459 (O_459,N_23829,N_22211);
nand UO_460 (O_460,N_24237,N_22183);
or UO_461 (O_461,N_24033,N_22179);
nor UO_462 (O_462,N_22095,N_23728);
nand UO_463 (O_463,N_22773,N_23528);
nand UO_464 (O_464,N_21984,N_23692);
nor UO_465 (O_465,N_24622,N_22939);
nor UO_466 (O_466,N_21914,N_24090);
nor UO_467 (O_467,N_23984,N_24649);
or UO_468 (O_468,N_24355,N_22365);
xor UO_469 (O_469,N_24785,N_23075);
nor UO_470 (O_470,N_23593,N_23377);
nor UO_471 (O_471,N_22621,N_24200);
nor UO_472 (O_472,N_24428,N_22885);
or UO_473 (O_473,N_22578,N_24432);
or UO_474 (O_474,N_21898,N_22061);
or UO_475 (O_475,N_23684,N_24718);
and UO_476 (O_476,N_22914,N_21949);
nor UO_477 (O_477,N_22540,N_23761);
or UO_478 (O_478,N_23877,N_22954);
nand UO_479 (O_479,N_23490,N_22878);
nand UO_480 (O_480,N_23227,N_24665);
or UO_481 (O_481,N_24396,N_24598);
nand UO_482 (O_482,N_23491,N_22905);
nor UO_483 (O_483,N_22420,N_24045);
and UO_484 (O_484,N_23866,N_23333);
and UO_485 (O_485,N_22468,N_24848);
and UO_486 (O_486,N_24042,N_23201);
nand UO_487 (O_487,N_23243,N_21959);
or UO_488 (O_488,N_22021,N_22243);
nor UO_489 (O_489,N_22731,N_24399);
nor UO_490 (O_490,N_23152,N_23167);
or UO_491 (O_491,N_23172,N_24347);
and UO_492 (O_492,N_24782,N_22210);
or UO_493 (O_493,N_22738,N_22918);
nand UO_494 (O_494,N_24073,N_23225);
and UO_495 (O_495,N_24948,N_22199);
or UO_496 (O_496,N_24751,N_24290);
nand UO_497 (O_497,N_24818,N_22930);
or UO_498 (O_498,N_23391,N_24447);
nand UO_499 (O_499,N_22350,N_22814);
or UO_500 (O_500,N_22014,N_22985);
nor UO_501 (O_501,N_24103,N_22702);
or UO_502 (O_502,N_24098,N_22703);
nor UO_503 (O_503,N_22138,N_23747);
or UO_504 (O_504,N_24629,N_22993);
and UO_505 (O_505,N_22509,N_22325);
nor UO_506 (O_506,N_22474,N_23816);
or UO_507 (O_507,N_23503,N_22403);
or UO_508 (O_508,N_24252,N_23612);
xor UO_509 (O_509,N_23163,N_23441);
nand UO_510 (O_510,N_22404,N_22608);
xor UO_511 (O_511,N_23585,N_22756);
xor UO_512 (O_512,N_24811,N_23777);
or UO_513 (O_513,N_23712,N_23946);
and UO_514 (O_514,N_24057,N_23309);
xor UO_515 (O_515,N_23030,N_23629);
and UO_516 (O_516,N_24056,N_22851);
nor UO_517 (O_517,N_24341,N_22725);
and UO_518 (O_518,N_22876,N_22447);
and UO_519 (O_519,N_23786,N_21938);
and UO_520 (O_520,N_22040,N_22960);
or UO_521 (O_521,N_23642,N_22687);
and UO_522 (O_522,N_23021,N_24397);
and UO_523 (O_523,N_22698,N_22589);
nand UO_524 (O_524,N_23203,N_21881);
nor UO_525 (O_525,N_24595,N_24712);
nor UO_526 (O_526,N_24048,N_24352);
nand UO_527 (O_527,N_23554,N_22380);
nand UO_528 (O_528,N_21958,N_22307);
and UO_529 (O_529,N_24023,N_22669);
nand UO_530 (O_530,N_23112,N_23069);
nor UO_531 (O_531,N_23596,N_22372);
nand UO_532 (O_532,N_23624,N_24113);
or UO_533 (O_533,N_23445,N_23087);
xnor UO_534 (O_534,N_24917,N_21918);
and UO_535 (O_535,N_23913,N_24102);
nand UO_536 (O_536,N_23869,N_23798);
or UO_537 (O_537,N_24425,N_24464);
and UO_538 (O_538,N_22513,N_22119);
and UO_539 (O_539,N_23638,N_22334);
and UO_540 (O_540,N_22116,N_22647);
nand UO_541 (O_541,N_23550,N_23179);
and UO_542 (O_542,N_22838,N_22571);
xor UO_543 (O_543,N_24747,N_24382);
or UO_544 (O_544,N_22161,N_24151);
nor UO_545 (O_545,N_22419,N_23730);
nor UO_546 (O_546,N_22611,N_24172);
xor UO_547 (O_547,N_22983,N_22312);
nor UO_548 (O_548,N_22601,N_22792);
and UO_549 (O_549,N_23949,N_24666);
nand UO_550 (O_550,N_24567,N_23746);
nor UO_551 (O_551,N_23932,N_23547);
nor UO_552 (O_552,N_24525,N_24273);
nand UO_553 (O_553,N_23532,N_22057);
and UO_554 (O_554,N_22439,N_23953);
and UO_555 (O_555,N_24035,N_23259);
and UO_556 (O_556,N_24512,N_24777);
or UO_557 (O_557,N_23987,N_24370);
nand UO_558 (O_558,N_24336,N_23466);
or UO_559 (O_559,N_24876,N_22143);
or UO_560 (O_560,N_24829,N_22796);
or UO_561 (O_561,N_23108,N_23043);
nor UO_562 (O_562,N_22393,N_22437);
and UO_563 (O_563,N_24743,N_24835);
nor UO_564 (O_564,N_24223,N_24118);
and UO_565 (O_565,N_23066,N_24742);
nor UO_566 (O_566,N_22382,N_24952);
nand UO_567 (O_567,N_23202,N_24318);
xnor UO_568 (O_568,N_23206,N_23908);
nor UO_569 (O_569,N_23660,N_24216);
xor UO_570 (O_570,N_24469,N_23357);
and UO_571 (O_571,N_24724,N_24678);
xnor UO_572 (O_572,N_22575,N_24680);
nand UO_573 (O_573,N_23930,N_24078);
nand UO_574 (O_574,N_22529,N_22285);
nand UO_575 (O_575,N_22283,N_22803);
and UO_576 (O_576,N_22809,N_22361);
nand UO_577 (O_577,N_22019,N_21926);
nor UO_578 (O_578,N_23574,N_21993);
nand UO_579 (O_579,N_22603,N_23551);
and UO_580 (O_580,N_24928,N_22323);
nand UO_581 (O_581,N_22935,N_22101);
and UO_582 (O_582,N_22880,N_22992);
and UO_583 (O_583,N_23005,N_22154);
nand UO_584 (O_584,N_24340,N_22498);
nor UO_585 (O_585,N_22906,N_22287);
and UO_586 (O_586,N_22531,N_22495);
or UO_587 (O_587,N_23241,N_24826);
nand UO_588 (O_588,N_23279,N_24631);
or UO_589 (O_589,N_23340,N_24860);
or UO_590 (O_590,N_22626,N_21989);
nor UO_591 (O_591,N_22240,N_24816);
nand UO_592 (O_592,N_24769,N_24670);
and UO_593 (O_593,N_23663,N_24060);
and UO_594 (O_594,N_22784,N_23755);
and UO_595 (O_595,N_24036,N_24094);
nor UO_596 (O_596,N_24189,N_21951);
nor UO_597 (O_597,N_23110,N_24845);
nor UO_598 (O_598,N_23298,N_24674);
nor UO_599 (O_599,N_21921,N_23331);
nor UO_600 (O_600,N_23139,N_22618);
nand UO_601 (O_601,N_24365,N_21976);
nand UO_602 (O_602,N_22129,N_22868);
nor UO_603 (O_603,N_23948,N_23464);
xnor UO_604 (O_604,N_23240,N_24675);
nand UO_605 (O_605,N_21894,N_24291);
and UO_606 (O_606,N_23204,N_23909);
or UO_607 (O_607,N_24005,N_22831);
or UO_608 (O_608,N_21998,N_22783);
or UO_609 (O_609,N_22244,N_22353);
xnor UO_610 (O_610,N_23261,N_22414);
nor UO_611 (O_611,N_24519,N_24834);
or UO_612 (O_612,N_23911,N_24322);
nand UO_613 (O_613,N_23792,N_22195);
or UO_614 (O_614,N_22078,N_22548);
nand UO_615 (O_615,N_21975,N_23192);
nand UO_616 (O_616,N_23373,N_23661);
nand UO_617 (O_617,N_21908,N_23264);
nand UO_618 (O_618,N_23939,N_24517);
or UO_619 (O_619,N_23421,N_24685);
and UO_620 (O_620,N_22494,N_23444);
or UO_621 (O_621,N_24232,N_23506);
or UO_622 (O_622,N_23868,N_22001);
and UO_623 (O_623,N_22583,N_24627);
and UO_624 (O_624,N_24913,N_24224);
and UO_625 (O_625,N_23643,N_22133);
and UO_626 (O_626,N_24049,N_23171);
and UO_627 (O_627,N_23601,N_21875);
or UO_628 (O_628,N_22815,N_24416);
and UO_629 (O_629,N_24490,N_24976);
and UO_630 (O_630,N_23292,N_22558);
nor UO_631 (O_631,N_24120,N_24528);
nand UO_632 (O_632,N_24420,N_24624);
or UO_633 (O_633,N_24770,N_23835);
nand UO_634 (O_634,N_21979,N_22456);
nor UO_635 (O_635,N_23916,N_23831);
or UO_636 (O_636,N_24987,N_22735);
and UO_637 (O_637,N_23905,N_22127);
nor UO_638 (O_638,N_24830,N_24395);
nor UO_639 (O_639,N_22048,N_24089);
or UO_640 (O_640,N_21924,N_24084);
nor UO_641 (O_641,N_23743,N_23542);
nand UO_642 (O_642,N_24485,N_24805);
and UO_643 (O_643,N_24698,N_22470);
nor UO_644 (O_644,N_23151,N_22102);
and UO_645 (O_645,N_23921,N_24636);
and UO_646 (O_646,N_24897,N_22170);
nand UO_647 (O_647,N_23236,N_22579);
and UO_648 (O_648,N_22123,N_22122);
or UO_649 (O_649,N_24393,N_23605);
nor UO_650 (O_650,N_23478,N_23109);
nor UO_651 (O_651,N_24767,N_24112);
or UO_652 (O_652,N_23966,N_24415);
and UO_653 (O_653,N_23422,N_22493);
and UO_654 (O_654,N_22039,N_23499);
or UO_655 (O_655,N_22920,N_24563);
or UO_656 (O_656,N_23611,N_24310);
nand UO_657 (O_657,N_24592,N_22230);
and UO_658 (O_658,N_24541,N_23092);
nand UO_659 (O_659,N_23142,N_22681);
or UO_660 (O_660,N_22917,N_22467);
nand UO_661 (O_661,N_24507,N_23733);
nor UO_662 (O_662,N_24233,N_21923);
nand UO_663 (O_663,N_24599,N_22998);
and UO_664 (O_664,N_24080,N_24572);
nor UO_665 (O_665,N_22002,N_22588);
nor UO_666 (O_666,N_24430,N_23310);
nor UO_667 (O_667,N_23826,N_23794);
or UO_668 (O_668,N_24076,N_24544);
nor UO_669 (O_669,N_23703,N_22883);
xor UO_670 (O_670,N_22469,N_24284);
or UO_671 (O_671,N_23231,N_22347);
or UO_672 (O_672,N_23055,N_23732);
and UO_673 (O_673,N_22237,N_22517);
nor UO_674 (O_674,N_22015,N_24961);
nand UO_675 (O_675,N_22250,N_24613);
and UO_676 (O_676,N_24337,N_24716);
or UO_677 (O_677,N_24797,N_23562);
and UO_678 (O_678,N_24803,N_22659);
nand UO_679 (O_679,N_22282,N_22713);
or UO_680 (O_680,N_22896,N_23844);
or UO_681 (O_681,N_24962,N_24282);
nor UO_682 (O_682,N_24799,N_24653);
xor UO_683 (O_683,N_24367,N_23754);
and UO_684 (O_684,N_23818,N_22058);
nand UO_685 (O_685,N_24740,N_23273);
and UO_686 (O_686,N_23150,N_24442);
or UO_687 (O_687,N_22570,N_24074);
xnor UO_688 (O_688,N_23669,N_24695);
or UO_689 (O_689,N_21992,N_23375);
or UO_690 (O_690,N_22830,N_23217);
nor UO_691 (O_691,N_21877,N_22990);
and UO_692 (O_692,N_22566,N_22961);
or UO_693 (O_693,N_24604,N_23888);
and UO_694 (O_694,N_22631,N_21953);
and UO_695 (O_695,N_22528,N_22079);
nand UO_696 (O_696,N_22268,N_22662);
nand UO_697 (O_697,N_23328,N_22218);
nand UO_698 (O_698,N_23469,N_22131);
nor UO_699 (O_699,N_22093,N_24561);
nand UO_700 (O_700,N_22144,N_22176);
xor UO_701 (O_701,N_22806,N_24063);
nand UO_702 (O_702,N_23392,N_24753);
and UO_703 (O_703,N_23105,N_24910);
or UO_704 (O_704,N_23361,N_23404);
nand UO_705 (O_705,N_21968,N_24873);
xnor UO_706 (O_706,N_23668,N_24325);
xnor UO_707 (O_707,N_24353,N_24597);
nor UO_708 (O_708,N_24985,N_22786);
and UO_709 (O_709,N_23873,N_23214);
and UO_710 (O_710,N_24761,N_24938);
nand UO_711 (O_711,N_22213,N_22141);
nor UO_712 (O_712,N_22869,N_23434);
or UO_713 (O_713,N_23620,N_22846);
nor UO_714 (O_714,N_24825,N_22392);
and UO_715 (O_715,N_24265,N_22190);
or UO_716 (O_716,N_23015,N_22075);
and UO_717 (O_717,N_22991,N_24691);
nand UO_718 (O_718,N_24375,N_23389);
and UO_719 (O_719,N_23263,N_22097);
nand UO_720 (O_720,N_23487,N_24877);
or UO_721 (O_721,N_23993,N_22351);
nor UO_722 (O_722,N_22054,N_22798);
xor UO_723 (O_723,N_21907,N_24221);
xor UO_724 (O_724,N_23952,N_22096);
nor UO_725 (O_725,N_21937,N_24247);
or UO_726 (O_726,N_23408,N_22339);
and UO_727 (O_727,N_23820,N_24040);
nand UO_728 (O_728,N_23031,N_23451);
nand UO_729 (O_729,N_22785,N_22676);
or UO_730 (O_730,N_22159,N_22239);
and UO_731 (O_731,N_22308,N_22988);
nor UO_732 (O_732,N_22822,N_23071);
nand UO_733 (O_733,N_22727,N_22124);
and UO_734 (O_734,N_24390,N_23327);
nand UO_735 (O_735,N_23314,N_23962);
nand UO_736 (O_736,N_23555,N_22458);
and UO_737 (O_737,N_24068,N_24827);
or UO_738 (O_738,N_23959,N_21930);
nand UO_739 (O_739,N_24387,N_23924);
nor UO_740 (O_740,N_24497,N_24439);
nor UO_741 (O_741,N_22088,N_22114);
and UO_742 (O_742,N_24772,N_23199);
nand UO_743 (O_743,N_22623,N_23937);
or UO_744 (O_744,N_23664,N_24657);
nor UO_745 (O_745,N_23415,N_22198);
nor UO_746 (O_746,N_23518,N_23674);
or UO_747 (O_747,N_24050,N_22441);
nand UO_748 (O_748,N_23688,N_24903);
or UO_749 (O_749,N_24467,N_24839);
nor UO_750 (O_750,N_23039,N_23345);
nor UO_751 (O_751,N_24275,N_22257);
nor UO_752 (O_752,N_24980,N_23893);
and UO_753 (O_753,N_23651,N_22134);
nand UO_754 (O_754,N_22017,N_23229);
and UO_755 (O_755,N_24381,N_23419);
nand UO_756 (O_756,N_23745,N_22893);
and UO_757 (O_757,N_23220,N_22755);
and UO_758 (O_758,N_24414,N_22544);
xnor UO_759 (O_759,N_23975,N_23537);
nor UO_760 (O_760,N_22089,N_22440);
nor UO_761 (O_761,N_22656,N_22732);
nor UO_762 (O_762,N_23918,N_24437);
and UO_763 (O_763,N_23125,N_22573);
xor UO_764 (O_764,N_22913,N_21892);
nor UO_765 (O_765,N_22084,N_22475);
and UO_766 (O_766,N_24717,N_24354);
or UO_767 (O_767,N_24616,N_23505);
nor UO_768 (O_768,N_24339,N_24401);
and UO_769 (O_769,N_24605,N_22744);
nand UO_770 (O_770,N_22835,N_22242);
and UO_771 (O_771,N_24534,N_21936);
and UO_772 (O_772,N_22449,N_24180);
and UO_773 (O_773,N_23531,N_23002);
nor UO_774 (O_774,N_23400,N_23215);
and UO_775 (O_775,N_22294,N_24972);
nand UO_776 (O_776,N_23722,N_22600);
or UO_777 (O_777,N_23394,N_22271);
and UO_778 (O_778,N_24106,N_22799);
or UO_779 (O_779,N_24121,N_22008);
nand UO_780 (O_780,N_22857,N_23284);
or UO_781 (O_781,N_23060,N_23132);
nor UO_782 (O_782,N_22511,N_23494);
nor UO_783 (O_783,N_24109,N_22009);
nand UO_784 (O_784,N_24004,N_23312);
or UO_785 (O_785,N_24986,N_23025);
nand UO_786 (O_786,N_23222,N_22465);
or UO_787 (O_787,N_23980,N_22336);
and UO_788 (O_788,N_23349,N_22060);
xor UO_789 (O_789,N_23787,N_21927);
and UO_790 (O_790,N_24788,N_22460);
nor UO_791 (O_791,N_22591,N_22749);
or UO_792 (O_792,N_24566,N_24448);
nor UO_793 (O_793,N_22761,N_23507);
nand UO_794 (O_794,N_22706,N_23196);
xnor UO_795 (O_795,N_24537,N_22805);
and UO_796 (O_796,N_23210,N_23160);
nand UO_797 (O_797,N_23138,N_21957);
nor UO_798 (O_798,N_24552,N_23329);
and UO_799 (O_799,N_23920,N_23976);
and UO_800 (O_800,N_23347,N_23102);
and UO_801 (O_801,N_24672,N_24008);
nor UO_802 (O_802,N_24892,N_23757);
and UO_803 (O_803,N_23033,N_22108);
and UO_804 (O_804,N_23635,N_22110);
nand UO_805 (O_805,N_23255,N_23875);
and UO_806 (O_806,N_22981,N_23990);
xor UO_807 (O_807,N_22412,N_22941);
or UO_808 (O_808,N_23401,N_23564);
and UO_809 (O_809,N_23175,N_22103);
nor UO_810 (O_810,N_24289,N_23676);
and UO_811 (O_811,N_24883,N_23520);
and UO_812 (O_812,N_23119,N_24266);
xnor UO_813 (O_813,N_23403,N_24495);
and UO_814 (O_814,N_23704,N_24015);
nand UO_815 (O_815,N_24235,N_22169);
xnor UO_816 (O_816,N_23049,N_24651);
or UO_817 (O_817,N_22866,N_23406);
and UO_818 (O_818,N_24570,N_24140);
nor UO_819 (O_819,N_23858,N_23841);
or UO_820 (O_820,N_24188,N_23376);
or UO_821 (O_821,N_24408,N_21994);
or UO_822 (O_822,N_22891,N_24287);
and UO_823 (O_823,N_22357,N_22952);
and UO_824 (O_824,N_24820,N_22197);
nor UO_825 (O_825,N_23791,N_23237);
and UO_826 (O_826,N_23758,N_22267);
nand UO_827 (O_827,N_23370,N_24277);
nand UO_828 (O_828,N_22807,N_23326);
or UO_829 (O_829,N_23751,N_24160);
nor UO_830 (O_830,N_23895,N_22163);
nand UO_831 (O_831,N_22871,N_24020);
and UO_832 (O_832,N_23455,N_23028);
and UO_833 (O_833,N_23830,N_24293);
and UO_834 (O_834,N_23022,N_22949);
nand UO_835 (O_835,N_22745,N_23126);
or UO_836 (O_836,N_22609,N_22674);
nand UO_837 (O_837,N_22436,N_22764);
nor UO_838 (O_838,N_22771,N_22614);
nor UO_839 (O_839,N_23998,N_23254);
nand UO_840 (O_840,N_23678,N_22545);
or UO_841 (O_841,N_24947,N_23558);
nor UO_842 (O_842,N_23300,N_22029);
or UO_843 (O_843,N_21889,N_24175);
and UO_844 (O_844,N_23512,N_24219);
nand UO_845 (O_845,N_22628,N_22715);
nand UO_846 (O_846,N_22619,N_23991);
nor UO_847 (O_847,N_23285,N_22083);
nand UO_848 (O_848,N_22099,N_24889);
nand UO_849 (O_849,N_23958,N_23626);
nand UO_850 (O_850,N_22966,N_24182);
and UO_851 (O_851,N_24582,N_22767);
or UO_852 (O_852,N_23677,N_24514);
or UO_853 (O_853,N_24334,N_23717);
and UO_854 (O_854,N_22053,N_24344);
nand UO_855 (O_855,N_23616,N_23857);
or UO_856 (O_856,N_24790,N_23797);
or UO_857 (O_857,N_23221,N_24141);
nor UO_858 (O_858,N_24373,N_24846);
nand UO_859 (O_859,N_22203,N_24046);
or UO_860 (O_860,N_24856,N_24758);
xnor UO_861 (O_861,N_22622,N_23007);
and UO_862 (O_862,N_22957,N_24600);
nor UO_863 (O_863,N_22115,N_23156);
or UO_864 (O_864,N_24417,N_22527);
nand UO_865 (O_865,N_22371,N_24461);
and UO_866 (O_866,N_24715,N_22486);
or UO_867 (O_867,N_23927,N_22612);
or UO_868 (O_868,N_23143,N_24129);
nand UO_869 (O_869,N_22406,N_24332);
and UO_870 (O_870,N_22506,N_23604);
nand UO_871 (O_871,N_22155,N_22461);
nor UO_872 (O_872,N_22225,N_22518);
or UO_873 (O_873,N_22301,N_21981);
nand UO_874 (O_874,N_24850,N_23186);
and UO_875 (O_875,N_22167,N_24638);
nor UO_876 (O_876,N_23164,N_22444);
nor UO_877 (O_877,N_24955,N_22316);
or UO_878 (O_878,N_23074,N_23010);
xor UO_879 (O_879,N_24967,N_23854);
nand UO_880 (O_880,N_24509,N_23398);
nand UO_881 (O_881,N_22565,N_24957);
nand UO_882 (O_882,N_23709,N_24493);
nor UO_883 (O_883,N_24067,N_22032);
nor UO_884 (O_884,N_22233,N_21931);
nor UO_885 (O_885,N_24307,N_22790);
or UO_886 (O_886,N_23036,N_24810);
or UO_887 (O_887,N_24918,N_24618);
and UO_888 (O_888,N_23559,N_22258);
nor UO_889 (O_889,N_23208,N_22843);
nor UO_890 (O_890,N_22894,N_22721);
and UO_891 (O_891,N_24722,N_23249);
or UO_892 (O_892,N_23153,N_22863);
xor UO_893 (O_893,N_22344,N_23162);
nor UO_894 (O_894,N_24176,N_24321);
and UO_895 (O_895,N_23318,N_23449);
nor UO_896 (O_896,N_22220,N_22157);
nor UO_897 (O_897,N_24671,N_24330);
nor UO_898 (O_898,N_24960,N_24843);
nand UO_899 (O_899,N_24654,N_22049);
or UO_900 (O_900,N_24436,N_23890);
nand UO_901 (O_901,N_24526,N_24124);
xnor UO_902 (O_902,N_24242,N_23900);
or UO_903 (O_903,N_22452,N_24359);
nand UO_904 (O_904,N_22840,N_23592);
or UO_905 (O_905,N_24323,N_24362);
and UO_906 (O_906,N_22711,N_22314);
or UO_907 (O_907,N_22383,N_23195);
or UO_908 (O_908,N_23705,N_22265);
and UO_909 (O_909,N_22847,N_23759);
or UO_910 (O_910,N_21996,N_24590);
and UO_911 (O_911,N_24285,N_24983);
and UO_912 (O_912,N_22766,N_21987);
nand UO_913 (O_913,N_22489,N_22251);
or UO_914 (O_914,N_24609,N_24923);
nand UO_915 (O_915,N_22450,N_24801);
nor UO_916 (O_916,N_23885,N_24013);
nand UO_917 (O_917,N_23566,N_23776);
and UO_918 (O_918,N_22510,N_23147);
and UO_919 (O_919,N_24487,N_22526);
or UO_920 (O_920,N_22153,N_24249);
and UO_921 (O_921,N_24153,N_24650);
or UO_922 (O_922,N_22080,N_22330);
and UO_923 (O_923,N_22675,N_23133);
or UO_924 (O_924,N_22018,N_23462);
xnor UO_925 (O_925,N_22272,N_23091);
nand UO_926 (O_926,N_22397,N_22861);
or UO_927 (O_927,N_24115,N_22148);
nor UO_928 (O_928,N_23169,N_24246);
and UO_929 (O_929,N_23416,N_23097);
and UO_930 (O_930,N_22793,N_23372);
nor UO_931 (O_931,N_24998,N_23556);
nor UO_932 (O_932,N_23051,N_23037);
or UO_933 (O_933,N_24838,N_24853);
or UO_934 (O_934,N_24804,N_24220);
nand UO_935 (O_935,N_21974,N_22636);
nor UO_936 (O_936,N_23630,N_24345);
or UO_937 (O_937,N_23013,N_22205);
or UO_938 (O_938,N_24866,N_23511);
and UO_939 (O_939,N_24869,N_23079);
and UO_940 (O_940,N_23439,N_21878);
or UO_941 (O_941,N_23803,N_21991);
nand UO_942 (O_942,N_22249,N_23335);
xor UO_943 (O_943,N_23850,N_24683);
and UO_944 (O_944,N_23513,N_24888);
nor UO_945 (O_945,N_23180,N_21946);
or UO_946 (O_946,N_23667,N_22164);
nor UO_947 (O_947,N_23773,N_22274);
and UO_948 (O_948,N_23718,N_22778);
nor UO_949 (O_949,N_22924,N_22327);
and UO_950 (O_950,N_24149,N_24764);
xnor UO_951 (O_951,N_23068,N_22693);
nor UO_952 (O_952,N_22321,N_24852);
and UO_953 (O_953,N_22660,N_22889);
nand UO_954 (O_954,N_23483,N_23658);
or UO_955 (O_955,N_24032,N_24317);
nand UO_956 (O_956,N_24471,N_23765);
or UO_957 (O_957,N_24477,N_23407);
nor UO_958 (O_958,N_21901,N_22500);
nor UO_959 (O_959,N_23170,N_23219);
nor UO_960 (O_960,N_23653,N_22582);
or UO_961 (O_961,N_23128,N_22151);
nor UO_962 (O_962,N_24261,N_24137);
or UO_963 (O_963,N_21952,N_24754);
nor UO_964 (O_964,N_23146,N_23363);
or UO_965 (O_965,N_22979,N_22910);
xor UO_966 (O_966,N_24550,N_24543);
nand UO_967 (O_967,N_23736,N_23707);
nand UO_968 (O_968,N_23978,N_24400);
and UO_969 (O_969,N_23165,N_24147);
and UO_970 (O_970,N_23336,N_23915);
or UO_971 (O_971,N_23693,N_22297);
or UO_972 (O_972,N_23561,N_24594);
nand UO_973 (O_973,N_23042,N_22026);
xnor UO_974 (O_974,N_22355,N_24244);
nand UO_975 (O_975,N_23815,N_23430);
nand UO_976 (O_976,N_24943,N_22602);
and UO_977 (O_977,N_23546,N_23904);
and UO_978 (O_978,N_22246,N_24916);
and UO_979 (O_979,N_23731,N_23879);
nand UO_980 (O_980,N_23650,N_24721);
xnor UO_981 (O_981,N_22929,N_23283);
nand UO_982 (O_982,N_24617,N_24136);
or UO_983 (O_983,N_23655,N_22791);
xnor UO_984 (O_984,N_23609,N_23615);
and UO_985 (O_985,N_23018,N_22996);
nor UO_986 (O_986,N_22670,N_24585);
nor UO_987 (O_987,N_24615,N_24051);
xnor UO_988 (O_988,N_24429,N_22563);
or UO_989 (O_989,N_22855,N_24929);
xor UO_990 (O_990,N_22111,N_22667);
nor UO_991 (O_991,N_24499,N_22020);
nor UO_992 (O_992,N_24186,N_24184);
and UO_993 (O_993,N_23078,N_22320);
and UO_994 (O_994,N_21902,N_24017);
and UO_995 (O_995,N_22358,N_23235);
nor UO_996 (O_996,N_22259,N_24596);
and UO_997 (O_997,N_24635,N_24404);
nand UO_998 (O_998,N_24156,N_24215);
nand UO_999 (O_999,N_23599,N_23744);
or UO_1000 (O_1000,N_24861,N_22085);
or UO_1001 (O_1001,N_22223,N_22284);
and UO_1002 (O_1002,N_23492,N_24714);
xor UO_1003 (O_1003,N_23288,N_24333);
nand UO_1004 (O_1004,N_23734,N_21883);
nor UO_1005 (O_1005,N_21970,N_24807);
nor UO_1006 (O_1006,N_24058,N_23713);
or UO_1007 (O_1007,N_22362,N_24920);
nor UO_1008 (O_1008,N_24407,N_22035);
nand UO_1009 (O_1009,N_23618,N_22248);
and UO_1010 (O_1010,N_23793,N_23977);
and UO_1011 (O_1011,N_24462,N_23586);
nand UO_1012 (O_1012,N_24403,N_22395);
nand UO_1013 (O_1013,N_22416,N_22288);
nor UO_1014 (O_1014,N_22254,N_22751);
nor UO_1015 (O_1015,N_24969,N_23770);
or UO_1016 (O_1016,N_22873,N_22677);
xor UO_1017 (O_1017,N_24449,N_24385);
or UO_1018 (O_1018,N_23242,N_22695);
nor UO_1019 (O_1019,N_22739,N_22201);
nor UO_1020 (O_1020,N_22633,N_24489);
nand UO_1021 (O_1021,N_24167,N_22668);
xnor UO_1022 (O_1022,N_23409,N_24210);
nor UO_1023 (O_1023,N_24603,N_24458);
nand UO_1024 (O_1024,N_24122,N_24568);
and UO_1025 (O_1025,N_22411,N_24725);
and UO_1026 (O_1026,N_24854,N_21915);
and UO_1027 (O_1027,N_23189,N_23453);
nor UO_1028 (O_1028,N_22598,N_23315);
xnor UO_1029 (O_1029,N_22024,N_24324);
nor UO_1030 (O_1030,N_22340,N_24009);
or UO_1031 (O_1031,N_23935,N_22405);
and UO_1032 (O_1032,N_24195,N_24276);
or UO_1033 (O_1033,N_22795,N_23343);
nand UO_1034 (O_1034,N_24766,N_23113);
nand UO_1035 (O_1035,N_24664,N_23774);
nor UO_1036 (O_1036,N_23321,N_22270);
nand UO_1037 (O_1037,N_23597,N_23951);
nand UO_1038 (O_1038,N_22277,N_24795);
and UO_1039 (O_1039,N_22824,N_24733);
xnor UO_1040 (O_1040,N_23683,N_23448);
or UO_1041 (O_1041,N_22209,N_24240);
xnor UO_1042 (O_1042,N_24435,N_22789);
nand UO_1043 (O_1043,N_24263,N_24248);
nor UO_1044 (O_1044,N_24542,N_21912);
or UO_1045 (O_1045,N_24398,N_23188);
or UO_1046 (O_1046,N_24547,N_21897);
and UO_1047 (O_1047,N_21890,N_22701);
nand UO_1048 (O_1048,N_24250,N_24431);
nand UO_1049 (O_1049,N_24475,N_22823);
nand UO_1050 (O_1050,N_23524,N_24498);
or UO_1051 (O_1051,N_22774,N_24502);
nor UO_1052 (O_1052,N_23428,N_23386);
nor UO_1053 (O_1053,N_22446,N_23077);
nand UO_1054 (O_1054,N_21935,N_22856);
or UO_1055 (O_1055,N_23120,N_24775);
nand UO_1056 (O_1056,N_23396,N_23127);
nand UO_1057 (O_1057,N_23836,N_23955);
nand UO_1058 (O_1058,N_22005,N_23447);
or UO_1059 (O_1059,N_24010,N_24077);
and UO_1060 (O_1060,N_23789,N_24862);
xor UO_1061 (O_1061,N_24906,N_23672);
and UO_1062 (O_1062,N_23687,N_23313);
xor UO_1063 (O_1063,N_23115,N_24771);
and UO_1064 (O_1064,N_22580,N_22682);
or UO_1065 (O_1065,N_24516,N_22160);
nand UO_1066 (O_1066,N_23569,N_24959);
nand UO_1067 (O_1067,N_22186,N_22022);
nand UO_1068 (O_1068,N_22010,N_24338);
nand UO_1069 (O_1069,N_22903,N_22794);
or UO_1070 (O_1070,N_24018,N_24346);
nor UO_1071 (O_1071,N_24075,N_22087);
or UO_1072 (O_1072,N_22833,N_23749);
and UO_1073 (O_1073,N_24262,N_23058);
xor UO_1074 (O_1074,N_22299,N_23988);
and UO_1075 (O_1075,N_22729,N_22104);
nand UO_1076 (O_1076,N_23756,N_22187);
nand UO_1077 (O_1077,N_23341,N_23947);
or UO_1078 (O_1078,N_23157,N_24919);
nand UO_1079 (O_1079,N_24737,N_23131);
nor UO_1080 (O_1080,N_23772,N_24630);
or UO_1081 (O_1081,N_22435,N_22263);
and UO_1082 (O_1082,N_22106,N_23649);
nor UO_1083 (O_1083,N_22304,N_22552);
nand UO_1084 (O_1084,N_24540,N_24583);
nor UO_1085 (O_1085,N_21967,N_23719);
and UO_1086 (O_1086,N_22377,N_22235);
nand UO_1087 (O_1087,N_22178,N_22886);
nor UO_1088 (O_1088,N_22356,N_23117);
or UO_1089 (O_1089,N_24097,N_22399);
nand UO_1090 (O_1090,N_24144,N_24719);
and UO_1091 (O_1091,N_24668,N_23048);
and UO_1092 (O_1092,N_23061,N_22839);
or UO_1093 (O_1093,N_24064,N_24559);
or UO_1094 (O_1094,N_22648,N_24043);
nand UO_1095 (O_1095,N_22890,N_23101);
and UO_1096 (O_1096,N_24196,N_24256);
nor UO_1097 (O_1097,N_24181,N_21925);
or UO_1098 (O_1098,N_23224,N_23154);
nor UO_1099 (O_1099,N_22128,N_23800);
xnor UO_1100 (O_1100,N_24872,N_21896);
and UO_1101 (O_1101,N_23486,N_22535);
or UO_1102 (O_1102,N_22543,N_23054);
nor UO_1103 (O_1103,N_24581,N_24912);
nor UO_1104 (O_1104,N_22997,N_24212);
or UO_1105 (O_1105,N_23739,N_23945);
xor UO_1106 (O_1106,N_24565,N_22338);
or UO_1107 (O_1107,N_21887,N_21985);
nand UO_1108 (O_1108,N_22262,N_22286);
xor UO_1109 (O_1109,N_22800,N_22421);
nand UO_1110 (O_1110,N_24135,N_24270);
or UO_1111 (O_1111,N_24626,N_23878);
xnor UO_1112 (O_1112,N_24392,N_23155);
nor UO_1113 (O_1113,N_23807,N_22343);
or UO_1114 (O_1114,N_23399,N_24061);
or UO_1115 (O_1115,N_24134,N_22925);
or UO_1116 (O_1116,N_23183,N_22834);
nand UO_1117 (O_1117,N_22599,N_23819);
xor UO_1118 (O_1118,N_21891,N_24637);
or UO_1119 (O_1119,N_22932,N_23636);
or UO_1120 (O_1120,N_22663,N_21943);
nand UO_1121 (O_1121,N_24069,N_22374);
and UO_1122 (O_1122,N_24847,N_22720);
nor UO_1123 (O_1123,N_22245,N_22707);
nor UO_1124 (O_1124,N_22829,N_22560);
xor UO_1125 (O_1125,N_23191,N_23107);
and UO_1126 (O_1126,N_24964,N_24794);
or UO_1127 (O_1127,N_24209,N_23213);
or UO_1128 (O_1128,N_24239,N_24968);
nor UO_1129 (O_1129,N_23426,N_23840);
nand UO_1130 (O_1130,N_22634,N_22139);
or UO_1131 (O_1131,N_23114,N_22853);
nor UO_1132 (O_1132,N_23685,N_24693);
nor UO_1133 (O_1133,N_22401,N_24450);
nand UO_1134 (O_1134,N_22652,N_23633);
or UO_1135 (O_1135,N_24697,N_22006);
or UO_1136 (O_1136,N_23934,N_22688);
or UO_1137 (O_1137,N_22946,N_23145);
and UO_1138 (O_1138,N_21917,N_24625);
nand UO_1139 (O_1139,N_22671,N_23290);
and UO_1140 (O_1140,N_24482,N_21910);
or UO_1141 (O_1141,N_23548,N_23892);
nor UO_1142 (O_1142,N_23572,N_24589);
or UO_1143 (O_1143,N_24145,N_24326);
nor UO_1144 (O_1144,N_24699,N_23782);
or UO_1145 (O_1145,N_24644,N_24880);
nand UO_1146 (O_1146,N_24506,N_23116);
nand UO_1147 (O_1147,N_23024,N_22559);
xnor UO_1148 (O_1148,N_23577,N_23641);
nor UO_1149 (O_1149,N_22479,N_21922);
nand UO_1150 (O_1150,N_22769,N_23632);
nand UO_1151 (O_1151,N_22788,N_24054);
and UO_1152 (O_1152,N_23802,N_22410);
nor UO_1153 (O_1153,N_24394,N_24173);
nand UO_1154 (O_1154,N_24749,N_21954);
and UO_1155 (O_1155,N_22322,N_23701);
nand UO_1156 (O_1156,N_23320,N_24875);
and UO_1157 (O_1157,N_22137,N_22937);
xor UO_1158 (O_1158,N_24492,N_24360);
nand UO_1159 (O_1159,N_22302,N_22945);
or UO_1160 (O_1160,N_23961,N_23184);
and UO_1161 (O_1161,N_22311,N_22923);
or UO_1162 (O_1162,N_22360,N_23019);
nor UO_1163 (O_1163,N_23085,N_23317);
nand UO_1164 (O_1164,N_23974,N_23332);
or UO_1165 (O_1165,N_23898,N_23194);
nand UO_1166 (O_1166,N_24900,N_23583);
and UO_1167 (O_1167,N_22586,N_24601);
nor UO_1168 (O_1168,N_23429,N_23498);
and UO_1169 (O_1169,N_23727,N_24836);
nor UO_1170 (O_1170,N_24763,N_24783);
and UO_1171 (O_1171,N_23964,N_24608);
and UO_1172 (O_1172,N_24996,N_23938);
or UO_1173 (O_1173,N_23045,N_23460);
and UO_1174 (O_1174,N_23278,N_24999);
xor UO_1175 (O_1175,N_23708,N_23454);
nor UO_1176 (O_1176,N_24292,N_24977);
nand UO_1177 (O_1177,N_23427,N_22523);
nand UO_1178 (O_1178,N_22200,N_23418);
nand UO_1179 (O_1179,N_24658,N_23305);
nand UO_1180 (O_1180,N_23862,N_23311);
nand UO_1181 (O_1181,N_22728,N_22310);
or UO_1182 (O_1182,N_23715,N_23846);
nor UO_1183 (O_1183,N_24349,N_24689);
and UO_1184 (O_1184,N_24858,N_22759);
nand UO_1185 (O_1185,N_23796,N_24745);
nor UO_1186 (O_1186,N_22165,N_23694);
and UO_1187 (O_1187,N_22331,N_24297);
nand UO_1188 (O_1188,N_24079,N_24410);
nand UO_1189 (O_1189,N_24191,N_23897);
nand UO_1190 (O_1190,N_22135,N_23933);
nor UO_1191 (O_1191,N_24548,N_24320);
or UO_1192 (O_1192,N_23931,N_22012);
nor UO_1193 (O_1193,N_22077,N_22828);
nand UO_1194 (O_1194,N_23808,N_24870);
nand UO_1195 (O_1195,N_23226,N_24021);
or UO_1196 (O_1196,N_22427,N_22915);
nor UO_1197 (O_1197,N_22387,N_23929);
nor UO_1198 (O_1198,N_22836,N_24308);
nor UO_1199 (O_1199,N_24933,N_22059);
nand UO_1200 (O_1200,N_22370,N_24227);
and UO_1201 (O_1201,N_24117,N_24686);
or UO_1202 (O_1202,N_24444,N_24104);
and UO_1203 (O_1203,N_23124,N_22959);
nor UO_1204 (O_1204,N_24110,N_24351);
and UO_1205 (O_1205,N_24688,N_22742);
or UO_1206 (O_1206,N_24119,N_23062);
nand UO_1207 (O_1207,N_23348,N_23926);
xor UO_1208 (O_1208,N_22714,N_21980);
and UO_1209 (O_1209,N_24271,N_24909);
and UO_1210 (O_1210,N_22379,N_23390);
nand UO_1211 (O_1211,N_22281,N_22295);
or UO_1212 (O_1212,N_24640,N_22031);
xor UO_1213 (O_1213,N_21886,N_22639);
and UO_1214 (O_1214,N_22520,N_22023);
nor UO_1215 (O_1215,N_24828,N_22472);
nor UO_1216 (O_1216,N_24575,N_22476);
nand UO_1217 (O_1217,N_23094,N_23986);
nand UO_1218 (O_1218,N_23082,N_23316);
or UO_1219 (O_1219,N_23575,N_23848);
or UO_1220 (O_1220,N_24662,N_23371);
or UO_1221 (O_1221,N_24025,N_23872);
nand UO_1222 (O_1222,N_22811,N_23504);
nor UO_1223 (O_1223,N_23832,N_22841);
or UO_1224 (O_1224,N_22679,N_22587);
and UO_1225 (O_1225,N_23248,N_24305);
nor UO_1226 (O_1226,N_24939,N_24019);
and UO_1227 (O_1227,N_22051,N_24001);
and UO_1228 (O_1228,N_22971,N_23510);
nor UO_1229 (O_1229,N_23515,N_22616);
nand UO_1230 (O_1230,N_24677,N_24831);
and UO_1231 (O_1231,N_23983,N_23525);
nand UO_1232 (O_1232,N_22279,N_23884);
and UO_1233 (O_1233,N_22463,N_23910);
nor UO_1234 (O_1234,N_22888,N_23047);
and UO_1235 (O_1235,N_22275,N_24205);
and UO_1236 (O_1236,N_22349,N_22038);
xor UO_1237 (O_1237,N_22968,N_23595);
nand UO_1238 (O_1238,N_23497,N_22396);
and UO_1239 (O_1239,N_24812,N_22974);
nand UO_1240 (O_1240,N_24837,N_23250);
xor UO_1241 (O_1241,N_22704,N_23488);
and UO_1242 (O_1242,N_24357,N_24087);
nor UO_1243 (O_1243,N_23385,N_24682);
nand UO_1244 (O_1244,N_23387,N_24701);
nand UO_1245 (O_1245,N_22508,N_22291);
or UO_1246 (O_1246,N_24111,N_24545);
and UO_1247 (O_1247,N_24645,N_22837);
or UO_1248 (O_1248,N_23319,N_24868);
nor UO_1249 (O_1249,N_23607,N_24463);
nor UO_1250 (O_1250,N_23223,N_22011);
nor UO_1251 (O_1251,N_22264,N_24538);
nor UO_1252 (O_1252,N_22276,N_23006);
nand UO_1253 (O_1253,N_24230,N_23258);
nor UO_1254 (O_1254,N_24895,N_23482);
nand UO_1255 (O_1255,N_23338,N_23941);
xor UO_1256 (O_1256,N_22772,N_23570);
xor UO_1257 (O_1257,N_24105,N_22664);
nor UO_1258 (O_1258,N_22464,N_23474);
nor UO_1259 (O_1259,N_23729,N_24915);
or UO_1260 (O_1260,N_22538,N_22112);
nor UO_1261 (O_1261,N_22324,N_22175);
nand UO_1262 (O_1262,N_22375,N_23587);
and UO_1263 (O_1263,N_22034,N_23675);
nand UO_1264 (O_1264,N_24798,N_24574);
nor UO_1265 (O_1265,N_22317,N_24014);
nand UO_1266 (O_1266,N_24460,N_24445);
nor UO_1267 (O_1267,N_23582,N_22922);
or UO_1268 (O_1268,N_22208,N_22373);
and UO_1269 (O_1269,N_23673,N_22860);
nand UO_1270 (O_1270,N_24584,N_23919);
nand UO_1271 (O_1271,N_23070,N_24279);
or UO_1272 (O_1272,N_23393,N_23657);
nor UO_1273 (O_1273,N_24114,N_22594);
and UO_1274 (O_1274,N_23647,N_24720);
and UO_1275 (O_1275,N_23304,N_22986);
and UO_1276 (O_1276,N_24424,N_23763);
nand UO_1277 (O_1277,N_24468,N_21961);
nor UO_1278 (O_1278,N_24992,N_23365);
and UO_1279 (O_1279,N_23549,N_23350);
or UO_1280 (O_1280,N_21977,N_22064);
or UO_1281 (O_1281,N_23766,N_24488);
nand UO_1282 (O_1282,N_23301,N_22827);
nor UO_1283 (O_1283,N_24006,N_23535);
xnor UO_1284 (O_1284,N_22503,N_22691);
and UO_1285 (O_1285,N_23899,N_24881);
or UO_1286 (O_1286,N_22453,N_24218);
or UO_1287 (O_1287,N_22091,N_23130);
nand UO_1288 (O_1288,N_22502,N_22989);
nor UO_1289 (O_1289,N_24932,N_24984);
xnor UO_1290 (O_1290,N_22995,N_24288);
nand UO_1291 (O_1291,N_21950,N_24907);
nand UO_1292 (O_1292,N_22572,N_22490);
and UO_1293 (O_1293,N_22146,N_24974);
nor UO_1294 (O_1294,N_23565,N_23682);
or UO_1295 (O_1295,N_22003,N_23589);
nand UO_1296 (O_1296,N_23671,N_22071);
nand UO_1297 (O_1297,N_23780,N_22867);
nand UO_1298 (O_1298,N_22638,N_24768);
nor UO_1299 (O_1299,N_23536,N_22743);
and UO_1300 (O_1300,N_22712,N_23631);
or UO_1301 (O_1301,N_22884,N_23134);
or UO_1302 (O_1302,N_22877,N_24760);
or UO_1303 (O_1303,N_23293,N_22515);
and UO_1304 (O_1304,N_23767,N_24776);
nor UO_1305 (O_1305,N_22962,N_24217);
or UO_1306 (O_1306,N_23886,N_22214);
or UO_1307 (O_1307,N_24995,N_22212);
or UO_1308 (O_1308,N_24945,N_24376);
or UO_1309 (O_1309,N_22070,N_24481);
nor UO_1310 (O_1310,N_24576,N_24634);
nor UO_1311 (O_1311,N_22987,N_22348);
and UO_1312 (O_1312,N_22422,N_24982);
nand UO_1313 (O_1313,N_22555,N_24222);
and UO_1314 (O_1314,N_23750,N_24150);
or UO_1315 (O_1315,N_22950,N_23710);
and UO_1316 (O_1316,N_23256,N_22269);
or UO_1317 (O_1317,N_22473,N_22238);
nand UO_1318 (O_1318,N_24491,N_21982);
and UO_1319 (O_1319,N_21939,N_24817);
nand UO_1320 (O_1320,N_22306,N_24245);
or UO_1321 (O_1321,N_24302,N_23303);
or UO_1322 (O_1322,N_23198,N_24350);
xnor UO_1323 (O_1323,N_24062,N_23799);
nor UO_1324 (O_1324,N_23790,N_22942);
xnor UO_1325 (O_1325,N_24269,N_21972);
nor UO_1326 (O_1326,N_23368,N_24206);
nand UO_1327 (O_1327,N_24694,N_22801);
or UO_1328 (O_1328,N_24705,N_22904);
or UO_1329 (O_1329,N_24383,N_24551);
nor UO_1330 (O_1330,N_21960,N_23251);
and UO_1331 (O_1331,N_24586,N_24942);
or UO_1332 (O_1332,N_24781,N_24730);
or UO_1333 (O_1333,N_22241,N_23783);
or UO_1334 (O_1334,N_24258,N_23177);
and UO_1335 (O_1335,N_22448,N_22428);
or UO_1336 (O_1336,N_21941,N_22497);
nor UO_1337 (O_1337,N_22074,N_21906);
or UO_1338 (O_1338,N_23989,N_22431);
nand UO_1339 (O_1339,N_24455,N_22655);
nor UO_1340 (O_1340,N_23239,N_22068);
or UO_1341 (O_1341,N_24676,N_22926);
xnor UO_1342 (O_1342,N_24159,N_22417);
and UO_1343 (O_1343,N_23824,N_23723);
nor UO_1344 (O_1344,N_22964,N_23099);
or UO_1345 (O_1345,N_24380,N_24893);
nor UO_1346 (O_1346,N_22651,N_22067);
nor UO_1347 (O_1347,N_22293,N_21940);
xnor UO_1348 (O_1348,N_23027,N_24708);
or UO_1349 (O_1349,N_22685,N_23943);
and UO_1350 (O_1350,N_24886,N_24727);
and UO_1351 (O_1351,N_24164,N_23760);
and UO_1352 (O_1352,N_23501,N_21888);
xnor UO_1353 (O_1353,N_24406,N_24202);
and UO_1354 (O_1354,N_23801,N_23724);
nor UO_1355 (O_1355,N_23606,N_23443);
or UO_1356 (O_1356,N_23280,N_23529);
nor UO_1357 (O_1357,N_23026,N_22780);
or UO_1358 (O_1358,N_23356,N_22980);
and UO_1359 (O_1359,N_22630,N_24494);
and UO_1360 (O_1360,N_22779,N_23804);
nor UO_1361 (O_1361,N_23925,N_22065);
and UO_1362 (O_1362,N_22136,N_22036);
nor UO_1363 (O_1363,N_23052,N_22524);
nor UO_1364 (O_1364,N_23567,N_23252);
xor UO_1365 (O_1365,N_22247,N_24808);
and UO_1366 (O_1366,N_24295,N_22665);
and UO_1367 (O_1367,N_24030,N_24580);
nand UO_1368 (O_1368,N_23838,N_24606);
and UO_1369 (O_1369,N_24855,N_23181);
and UO_1370 (O_1370,N_23081,N_24421);
or UO_1371 (O_1371,N_24857,N_23855);
nor UO_1372 (O_1372,N_23995,N_23851);
or UO_1373 (O_1373,N_23521,N_23140);
and UO_1374 (O_1374,N_23817,N_22564);
or UO_1375 (O_1375,N_23634,N_22848);
xor UO_1376 (O_1376,N_22390,N_22069);
nand UO_1377 (O_1377,N_24619,N_23032);
and UO_1378 (O_1378,N_23882,N_24882);
or UO_1379 (O_1379,N_24726,N_22121);
nand UO_1380 (O_1380,N_24620,N_21900);
or UO_1381 (O_1381,N_24123,N_23680);
and UO_1382 (O_1382,N_24833,N_24358);
and UO_1383 (O_1383,N_24573,N_23716);
nand UO_1384 (O_1384,N_24632,N_23912);
xor UO_1385 (O_1385,N_22593,N_21942);
nand UO_1386 (O_1386,N_24966,N_24791);
nand UO_1387 (O_1387,N_23965,N_24085);
or UO_1388 (O_1388,N_23351,N_23997);
nor UO_1389 (O_1389,N_24199,N_24081);
nand UO_1390 (O_1390,N_23972,N_22733);
and UO_1391 (O_1391,N_24971,N_22546);
nor UO_1392 (O_1392,N_24555,N_23158);
or UO_1393 (O_1393,N_22181,N_24211);
or UO_1394 (O_1394,N_24773,N_24072);
nand UO_1395 (O_1395,N_24963,N_24229);
nand UO_1396 (O_1396,N_22907,N_24412);
and UO_1397 (O_1397,N_24055,N_23388);
nor UO_1398 (O_1398,N_24821,N_22363);
and UO_1399 (O_1399,N_24894,N_23539);
and UO_1400 (O_1400,N_22354,N_23666);
or UO_1401 (O_1401,N_23440,N_24936);
nor UO_1402 (O_1402,N_24127,N_24554);
and UO_1403 (O_1403,N_24082,N_23295);
nor UO_1404 (O_1404,N_23004,N_22845);
nor UO_1405 (O_1405,N_22673,N_22046);
nor UO_1406 (O_1406,N_23262,N_22290);
nand UO_1407 (O_1407,N_24092,N_24591);
nand UO_1408 (O_1408,N_22217,N_22224);
nor UO_1409 (O_1409,N_23000,N_22149);
nand UO_1410 (O_1410,N_22296,N_23870);
or UO_1411 (O_1411,N_23017,N_24161);
and UO_1412 (O_1412,N_23588,N_23161);
nand UO_1413 (O_1413,N_21893,N_22754);
nand UO_1414 (O_1414,N_23859,N_24314);
nor UO_1415 (O_1415,N_22534,N_22300);
nor UO_1416 (O_1416,N_22483,N_24729);
xor UO_1417 (O_1417,N_23896,N_22708);
xor UO_1418 (O_1418,N_22303,N_24426);
nor UO_1419 (O_1419,N_22496,N_22082);
or UO_1420 (O_1420,N_23106,N_23533);
and UO_1421 (O_1421,N_22976,N_23098);
xnor UO_1422 (O_1422,N_24108,N_22975);
nand UO_1423 (O_1423,N_22752,N_24260);
nor UO_1424 (O_1424,N_22777,N_24736);
nand UO_1425 (O_1425,N_24024,N_24796);
nor UO_1426 (O_1426,N_24800,N_22977);
nor UO_1427 (O_1427,N_23468,N_22649);
nor UO_1428 (O_1428,N_22994,N_22551);
or UO_1429 (O_1429,N_23690,N_24372);
xor UO_1430 (O_1430,N_22694,N_23493);
nor UO_1431 (O_1431,N_23111,N_24422);
and UO_1432 (O_1432,N_24259,N_24611);
nor UO_1433 (O_1433,N_24298,N_24433);
and UO_1434 (O_1434,N_24028,N_24503);
and UO_1435 (O_1435,N_22782,N_22597);
nand UO_1436 (O_1436,N_24663,N_22646);
nand UO_1437 (O_1437,N_23008,N_22854);
and UO_1438 (O_1438,N_24052,N_23269);
or UO_1439 (O_1439,N_22345,N_24391);
nor UO_1440 (O_1440,N_24254,N_24756);
nor UO_1441 (O_1441,N_23056,N_22042);
nand UO_1442 (O_1442,N_22172,N_24973);
nand UO_1443 (O_1443,N_24107,N_23410);
nor UO_1444 (O_1444,N_24787,N_22596);
xnor UO_1445 (O_1445,N_22207,N_23475);
and UO_1446 (O_1446,N_24070,N_21955);
nor UO_1447 (O_1447,N_22737,N_22033);
or UO_1448 (O_1448,N_24388,N_22723);
xnor UO_1449 (O_1449,N_24331,N_22415);
or UO_1450 (O_1450,N_23699,N_22763);
xnor UO_1451 (O_1451,N_23274,N_24378);
or UO_1452 (O_1452,N_24546,N_21880);
or UO_1453 (O_1453,N_23695,N_22900);
nand UO_1454 (O_1454,N_22781,N_22722);
or UO_1455 (O_1455,N_23275,N_24710);
or UO_1456 (O_1456,N_22255,N_22204);
nor UO_1457 (O_1457,N_22227,N_22094);
nor UO_1458 (O_1458,N_23035,N_22541);
and UO_1459 (O_1459,N_24778,N_24456);
and UO_1460 (O_1460,N_24508,N_24988);
and UO_1461 (O_1461,N_23187,N_24646);
nor UO_1462 (O_1462,N_22142,N_22642);
nand UO_1463 (O_1463,N_23253,N_22292);
or UO_1464 (O_1464,N_23425,N_22645);
and UO_1465 (O_1465,N_22391,N_22056);
or UO_1466 (O_1466,N_22901,N_24558);
nand UO_1467 (O_1467,N_23395,N_23779);
and UO_1468 (O_1468,N_22605,N_23216);
or UO_1469 (O_1469,N_24178,N_23166);
and UO_1470 (O_1470,N_22882,N_22881);
nor UO_1471 (O_1471,N_23190,N_23297);
nand UO_1472 (O_1472,N_22613,N_22368);
and UO_1473 (O_1473,N_22037,N_24169);
and UO_1474 (O_1474,N_22716,N_23652);
nand UO_1475 (O_1475,N_22335,N_24041);
nand UO_1476 (O_1476,N_23720,N_21895);
and UO_1477 (O_1477,N_23578,N_24255);
or UO_1478 (O_1478,N_24003,N_24944);
xor UO_1479 (O_1479,N_24300,N_22734);
nor UO_1480 (O_1480,N_24579,N_22228);
nor UO_1481 (O_1481,N_23881,N_23867);
nor UO_1482 (O_1482,N_24466,N_24312);
and UO_1483 (O_1483,N_24472,N_23063);
nor UO_1484 (O_1484,N_23639,N_23619);
xnor UO_1485 (O_1485,N_24453,N_22487);
nand UO_1486 (O_1486,N_23670,N_21903);
nor UO_1487 (O_1487,N_23353,N_22090);
nor UO_1488 (O_1488,N_23433,N_22696);
xnor UO_1489 (O_1489,N_23144,N_23656);
nand UO_1490 (O_1490,N_23970,N_22341);
xnor UO_1491 (O_1491,N_23922,N_24863);
nor UO_1492 (O_1492,N_22967,N_23465);
or UO_1493 (O_1493,N_22202,N_21882);
xnor UO_1494 (O_1494,N_24368,N_23364);
or UO_1495 (O_1495,N_22445,N_23472);
nor UO_1496 (O_1496,N_23458,N_22388);
and UO_1497 (O_1497,N_23741,N_23883);
and UO_1498 (O_1498,N_22499,N_22537);
and UO_1499 (O_1499,N_23617,N_22584);
nor UO_1500 (O_1500,N_24208,N_22232);
or UO_1501 (O_1501,N_24197,N_22229);
nand UO_1502 (O_1502,N_24152,N_22385);
nand UO_1503 (O_1503,N_24530,N_24451);
and UO_1504 (O_1504,N_21986,N_24723);
and UO_1505 (O_1505,N_23516,N_22342);
nand UO_1506 (O_1506,N_22797,N_22730);
and UO_1507 (O_1507,N_22063,N_23627);
nand UO_1508 (O_1508,N_21933,N_22252);
nor UO_1509 (O_1509,N_24755,N_23936);
nor UO_1510 (O_1510,N_22514,N_24659);
nor UO_1511 (O_1511,N_24628,N_24088);
nor UO_1512 (O_1512,N_24911,N_23477);
xnor UO_1513 (O_1513,N_22481,N_24480);
or UO_1514 (O_1514,N_22549,N_22832);
nor UO_1515 (O_1515,N_22459,N_24304);
nor UO_1516 (O_1516,N_23622,N_24673);
and UO_1517 (O_1517,N_24286,N_22423);
and UO_1518 (O_1518,N_24744,N_24809);
or UO_1519 (O_1519,N_24272,N_23971);
nand UO_1520 (O_1520,N_22821,N_22746);
xor UO_1521 (O_1521,N_22718,N_23837);
nor UO_1522 (O_1522,N_24511,N_23374);
nor UO_1523 (O_1523,N_22933,N_24607);
and UO_1524 (O_1524,N_21929,N_23149);
or UO_1525 (O_1525,N_23812,N_22055);
nor UO_1526 (O_1526,N_24143,N_23090);
or UO_1527 (O_1527,N_24732,N_21911);
nand UO_1528 (O_1528,N_22700,N_23148);
xor UO_1529 (O_1529,N_22266,N_24264);
nand UO_1530 (O_1530,N_24027,N_23740);
and UO_1531 (O_1531,N_22595,N_23384);
nor UO_1532 (O_1532,N_23981,N_22109);
and UO_1533 (O_1533,N_24990,N_23640);
and UO_1534 (O_1534,N_23413,N_24643);
and UO_1535 (O_1535,N_24100,N_23571);
nor UO_1536 (O_1536,N_23402,N_22313);
nand UO_1537 (O_1537,N_23452,N_22686);
nor UO_1538 (O_1538,N_22825,N_22156);
nor UO_1539 (O_1539,N_22748,N_23436);
and UO_1540 (O_1540,N_22426,N_21947);
and UO_1541 (O_1541,N_24521,N_22948);
nor UO_1542 (O_1542,N_22025,N_24562);
or UO_1543 (O_1543,N_24207,N_22066);
nor UO_1544 (O_1544,N_24802,N_23982);
nand UO_1545 (O_1545,N_22817,N_24496);
nor UO_1546 (O_1546,N_22219,N_23470);
xor UO_1547 (O_1547,N_24313,N_22504);
or UO_1548 (O_1548,N_23267,N_22862);
nor UO_1549 (O_1549,N_23209,N_24170);
and UO_1550 (O_1550,N_23887,N_24226);
or UO_1551 (O_1551,N_23244,N_22369);
nor UO_1552 (O_1552,N_24587,N_22577);
nor UO_1553 (O_1553,N_23420,N_22280);
nor UO_1554 (O_1554,N_22710,N_22661);
nor UO_1555 (O_1555,N_22477,N_24434);
and UO_1556 (O_1556,N_23646,N_24823);
and UO_1557 (O_1557,N_23168,N_22943);
or UO_1558 (O_1558,N_24441,N_24531);
or UO_1559 (O_1559,N_24588,N_24031);
and UO_1560 (O_1560,N_23266,N_23118);
and UO_1561 (O_1561,N_24283,N_24921);
and UO_1562 (O_1562,N_21988,N_22824);
nand UO_1563 (O_1563,N_23187,N_23177);
nand UO_1564 (O_1564,N_23005,N_24559);
or UO_1565 (O_1565,N_24049,N_23606);
or UO_1566 (O_1566,N_23633,N_24408);
xnor UO_1567 (O_1567,N_24612,N_22479);
nor UO_1568 (O_1568,N_23164,N_23461);
xnor UO_1569 (O_1569,N_23276,N_22931);
xnor UO_1570 (O_1570,N_22031,N_22460);
and UO_1571 (O_1571,N_22974,N_22705);
or UO_1572 (O_1572,N_24819,N_22752);
or UO_1573 (O_1573,N_24215,N_22878);
or UO_1574 (O_1574,N_23952,N_23515);
nand UO_1575 (O_1575,N_21938,N_22982);
or UO_1576 (O_1576,N_22090,N_23271);
and UO_1577 (O_1577,N_22239,N_24443);
nand UO_1578 (O_1578,N_22092,N_22620);
and UO_1579 (O_1579,N_21901,N_23065);
xnor UO_1580 (O_1580,N_24005,N_22233);
and UO_1581 (O_1581,N_23922,N_22429);
xnor UO_1582 (O_1582,N_23663,N_24771);
and UO_1583 (O_1583,N_23760,N_22776);
nand UO_1584 (O_1584,N_23268,N_22556);
nor UO_1585 (O_1585,N_23371,N_23770);
and UO_1586 (O_1586,N_22492,N_23755);
nor UO_1587 (O_1587,N_22433,N_21939);
nor UO_1588 (O_1588,N_22968,N_23301);
xor UO_1589 (O_1589,N_24052,N_24144);
nor UO_1590 (O_1590,N_23141,N_22011);
nor UO_1591 (O_1591,N_22840,N_22306);
nand UO_1592 (O_1592,N_23278,N_23976);
or UO_1593 (O_1593,N_23687,N_22150);
nand UO_1594 (O_1594,N_22077,N_22756);
or UO_1595 (O_1595,N_24093,N_21947);
xnor UO_1596 (O_1596,N_24145,N_21888);
or UO_1597 (O_1597,N_22429,N_23840);
or UO_1598 (O_1598,N_22715,N_24369);
nand UO_1599 (O_1599,N_22916,N_23547);
and UO_1600 (O_1600,N_23834,N_23485);
nor UO_1601 (O_1601,N_23673,N_24343);
or UO_1602 (O_1602,N_22335,N_24858);
nor UO_1603 (O_1603,N_24802,N_24625);
or UO_1604 (O_1604,N_23611,N_22931);
or UO_1605 (O_1605,N_22584,N_23937);
nand UO_1606 (O_1606,N_22037,N_22376);
xor UO_1607 (O_1607,N_23115,N_21987);
and UO_1608 (O_1608,N_23885,N_22986);
and UO_1609 (O_1609,N_23917,N_24112);
or UO_1610 (O_1610,N_24544,N_23201);
xor UO_1611 (O_1611,N_24806,N_24367);
and UO_1612 (O_1612,N_23061,N_23472);
nand UO_1613 (O_1613,N_23382,N_24564);
nor UO_1614 (O_1614,N_24348,N_24527);
nand UO_1615 (O_1615,N_23037,N_22016);
nor UO_1616 (O_1616,N_22175,N_22657);
or UO_1617 (O_1617,N_24858,N_23094);
nor UO_1618 (O_1618,N_24008,N_24238);
xnor UO_1619 (O_1619,N_23385,N_23984);
nand UO_1620 (O_1620,N_24581,N_23697);
nand UO_1621 (O_1621,N_22795,N_24643);
and UO_1622 (O_1622,N_24444,N_23456);
and UO_1623 (O_1623,N_24550,N_23362);
nand UO_1624 (O_1624,N_22084,N_23375);
xor UO_1625 (O_1625,N_24344,N_21976);
nor UO_1626 (O_1626,N_21937,N_22591);
or UO_1627 (O_1627,N_24254,N_23592);
and UO_1628 (O_1628,N_22350,N_22035);
or UO_1629 (O_1629,N_23215,N_23514);
nand UO_1630 (O_1630,N_22778,N_22268);
nor UO_1631 (O_1631,N_21915,N_22758);
nand UO_1632 (O_1632,N_23440,N_23781);
nand UO_1633 (O_1633,N_24395,N_23963);
and UO_1634 (O_1634,N_22935,N_24801);
nand UO_1635 (O_1635,N_24626,N_24738);
and UO_1636 (O_1636,N_22746,N_24568);
nand UO_1637 (O_1637,N_24907,N_22311);
and UO_1638 (O_1638,N_24906,N_23171);
nand UO_1639 (O_1639,N_23499,N_24536);
and UO_1640 (O_1640,N_22125,N_24801);
nand UO_1641 (O_1641,N_22137,N_24443);
xnor UO_1642 (O_1642,N_24806,N_24020);
xnor UO_1643 (O_1643,N_23717,N_23467);
nor UO_1644 (O_1644,N_23079,N_23524);
nand UO_1645 (O_1645,N_22813,N_22474);
nor UO_1646 (O_1646,N_24765,N_24278);
and UO_1647 (O_1647,N_21964,N_24307);
nor UO_1648 (O_1648,N_24024,N_23334);
xor UO_1649 (O_1649,N_24364,N_22102);
or UO_1650 (O_1650,N_24255,N_23415);
and UO_1651 (O_1651,N_22859,N_22673);
nand UO_1652 (O_1652,N_24882,N_23073);
nand UO_1653 (O_1653,N_24332,N_23738);
nand UO_1654 (O_1654,N_23062,N_24149);
xor UO_1655 (O_1655,N_22987,N_22456);
or UO_1656 (O_1656,N_24968,N_22578);
and UO_1657 (O_1657,N_22868,N_22442);
or UO_1658 (O_1658,N_22467,N_23110);
nand UO_1659 (O_1659,N_23736,N_23244);
or UO_1660 (O_1660,N_24162,N_23792);
or UO_1661 (O_1661,N_22311,N_22693);
and UO_1662 (O_1662,N_23089,N_24817);
nor UO_1663 (O_1663,N_24395,N_23755);
xnor UO_1664 (O_1664,N_23821,N_21956);
or UO_1665 (O_1665,N_23802,N_23139);
nor UO_1666 (O_1666,N_24053,N_22493);
or UO_1667 (O_1667,N_22816,N_22209);
and UO_1668 (O_1668,N_23926,N_21986);
or UO_1669 (O_1669,N_23947,N_24764);
nand UO_1670 (O_1670,N_22225,N_24328);
nand UO_1671 (O_1671,N_22363,N_22683);
xnor UO_1672 (O_1672,N_23729,N_23786);
or UO_1673 (O_1673,N_24916,N_22746);
and UO_1674 (O_1674,N_24408,N_23180);
or UO_1675 (O_1675,N_22967,N_22890);
nand UO_1676 (O_1676,N_24757,N_24202);
xnor UO_1677 (O_1677,N_24945,N_23191);
and UO_1678 (O_1678,N_23699,N_23406);
nand UO_1679 (O_1679,N_22687,N_23356);
and UO_1680 (O_1680,N_24367,N_22034);
and UO_1681 (O_1681,N_24252,N_21916);
nor UO_1682 (O_1682,N_24175,N_24558);
or UO_1683 (O_1683,N_22716,N_23961);
nand UO_1684 (O_1684,N_24486,N_24679);
nor UO_1685 (O_1685,N_24017,N_24362);
nand UO_1686 (O_1686,N_22984,N_22096);
or UO_1687 (O_1687,N_23330,N_22804);
and UO_1688 (O_1688,N_22941,N_23013);
and UO_1689 (O_1689,N_22440,N_22528);
or UO_1690 (O_1690,N_21918,N_22514);
nand UO_1691 (O_1691,N_21984,N_22845);
nor UO_1692 (O_1692,N_23927,N_23690);
nand UO_1693 (O_1693,N_22430,N_22775);
nor UO_1694 (O_1694,N_23146,N_24031);
nor UO_1695 (O_1695,N_22305,N_24735);
nand UO_1696 (O_1696,N_22215,N_23319);
nand UO_1697 (O_1697,N_23398,N_24664);
nand UO_1698 (O_1698,N_23046,N_23403);
nand UO_1699 (O_1699,N_23336,N_24599);
or UO_1700 (O_1700,N_23884,N_24664);
or UO_1701 (O_1701,N_23399,N_22385);
nand UO_1702 (O_1702,N_24417,N_22282);
nand UO_1703 (O_1703,N_22079,N_23377);
nand UO_1704 (O_1704,N_24148,N_22060);
or UO_1705 (O_1705,N_22143,N_22585);
nor UO_1706 (O_1706,N_22380,N_24219);
nor UO_1707 (O_1707,N_23803,N_22106);
xnor UO_1708 (O_1708,N_22242,N_24959);
nor UO_1709 (O_1709,N_22742,N_23500);
xnor UO_1710 (O_1710,N_22201,N_22093);
xnor UO_1711 (O_1711,N_24075,N_23162);
or UO_1712 (O_1712,N_22173,N_23784);
and UO_1713 (O_1713,N_23937,N_24682);
nor UO_1714 (O_1714,N_22211,N_22005);
and UO_1715 (O_1715,N_22879,N_23745);
or UO_1716 (O_1716,N_24598,N_23162);
nand UO_1717 (O_1717,N_23258,N_24410);
and UO_1718 (O_1718,N_24716,N_22758);
nand UO_1719 (O_1719,N_22148,N_22401);
or UO_1720 (O_1720,N_24030,N_22024);
nand UO_1721 (O_1721,N_23957,N_22890);
and UO_1722 (O_1722,N_23852,N_23355);
nor UO_1723 (O_1723,N_21903,N_24304);
and UO_1724 (O_1724,N_24849,N_22857);
or UO_1725 (O_1725,N_24854,N_23570);
or UO_1726 (O_1726,N_23662,N_22678);
nor UO_1727 (O_1727,N_23909,N_23475);
nor UO_1728 (O_1728,N_23575,N_22664);
xnor UO_1729 (O_1729,N_22328,N_22863);
and UO_1730 (O_1730,N_24741,N_23449);
nand UO_1731 (O_1731,N_21881,N_21909);
nor UO_1732 (O_1732,N_24512,N_22169);
nor UO_1733 (O_1733,N_22522,N_24988);
or UO_1734 (O_1734,N_24864,N_22820);
xor UO_1735 (O_1735,N_23116,N_23870);
nor UO_1736 (O_1736,N_23092,N_24195);
and UO_1737 (O_1737,N_24700,N_24145);
nor UO_1738 (O_1738,N_23416,N_24853);
and UO_1739 (O_1739,N_24283,N_22861);
or UO_1740 (O_1740,N_22912,N_24071);
and UO_1741 (O_1741,N_24485,N_23721);
nor UO_1742 (O_1742,N_22293,N_23310);
nand UO_1743 (O_1743,N_22039,N_22948);
nand UO_1744 (O_1744,N_24987,N_23756);
and UO_1745 (O_1745,N_23176,N_21880);
and UO_1746 (O_1746,N_23578,N_23661);
and UO_1747 (O_1747,N_22742,N_23149);
nand UO_1748 (O_1748,N_24110,N_23845);
nand UO_1749 (O_1749,N_24573,N_22595);
or UO_1750 (O_1750,N_22229,N_22818);
nor UO_1751 (O_1751,N_22609,N_24979);
and UO_1752 (O_1752,N_23492,N_23065);
or UO_1753 (O_1753,N_22741,N_22556);
nand UO_1754 (O_1754,N_23272,N_23133);
nand UO_1755 (O_1755,N_24338,N_22316);
and UO_1756 (O_1756,N_24451,N_23860);
nand UO_1757 (O_1757,N_24304,N_22868);
nor UO_1758 (O_1758,N_24325,N_24121);
nand UO_1759 (O_1759,N_23480,N_24279);
or UO_1760 (O_1760,N_22137,N_24940);
or UO_1761 (O_1761,N_24211,N_22763);
and UO_1762 (O_1762,N_23885,N_24980);
or UO_1763 (O_1763,N_23579,N_23347);
and UO_1764 (O_1764,N_24596,N_24277);
nor UO_1765 (O_1765,N_23624,N_24344);
xnor UO_1766 (O_1766,N_22951,N_23892);
nand UO_1767 (O_1767,N_24159,N_24346);
nand UO_1768 (O_1768,N_24546,N_23146);
nand UO_1769 (O_1769,N_24998,N_24337);
nand UO_1770 (O_1770,N_24095,N_24448);
nor UO_1771 (O_1771,N_22049,N_22555);
nand UO_1772 (O_1772,N_24582,N_24025);
or UO_1773 (O_1773,N_24829,N_22451);
or UO_1774 (O_1774,N_23032,N_23870);
nor UO_1775 (O_1775,N_23107,N_22783);
xor UO_1776 (O_1776,N_23538,N_22340);
xor UO_1777 (O_1777,N_22227,N_23213);
nor UO_1778 (O_1778,N_24061,N_22008);
nor UO_1779 (O_1779,N_23402,N_21877);
and UO_1780 (O_1780,N_22489,N_22237);
or UO_1781 (O_1781,N_22517,N_22479);
nand UO_1782 (O_1782,N_23582,N_23051);
nor UO_1783 (O_1783,N_22578,N_23588);
nand UO_1784 (O_1784,N_23425,N_24677);
nand UO_1785 (O_1785,N_24009,N_22507);
nand UO_1786 (O_1786,N_23242,N_24055);
or UO_1787 (O_1787,N_22202,N_22447);
xor UO_1788 (O_1788,N_21904,N_21919);
and UO_1789 (O_1789,N_24004,N_22281);
nor UO_1790 (O_1790,N_21921,N_23247);
nand UO_1791 (O_1791,N_22228,N_23550);
or UO_1792 (O_1792,N_23315,N_23835);
and UO_1793 (O_1793,N_23695,N_24008);
nor UO_1794 (O_1794,N_24134,N_23278);
nor UO_1795 (O_1795,N_24006,N_24051);
nor UO_1796 (O_1796,N_23524,N_22909);
or UO_1797 (O_1797,N_24314,N_24548);
nor UO_1798 (O_1798,N_22880,N_24184);
xor UO_1799 (O_1799,N_24176,N_22715);
nor UO_1800 (O_1800,N_23952,N_23312);
nand UO_1801 (O_1801,N_22100,N_24109);
or UO_1802 (O_1802,N_22745,N_24607);
nand UO_1803 (O_1803,N_23835,N_23926);
or UO_1804 (O_1804,N_22706,N_23304);
or UO_1805 (O_1805,N_22304,N_24397);
xnor UO_1806 (O_1806,N_23922,N_21875);
nor UO_1807 (O_1807,N_22390,N_21891);
nor UO_1808 (O_1808,N_24253,N_23921);
or UO_1809 (O_1809,N_23260,N_22815);
or UO_1810 (O_1810,N_23459,N_23882);
nand UO_1811 (O_1811,N_24642,N_24496);
or UO_1812 (O_1812,N_22331,N_24743);
or UO_1813 (O_1813,N_23581,N_23359);
nand UO_1814 (O_1814,N_22765,N_23439);
nand UO_1815 (O_1815,N_24122,N_22111);
nand UO_1816 (O_1816,N_22187,N_24897);
nand UO_1817 (O_1817,N_24116,N_23545);
or UO_1818 (O_1818,N_23494,N_22352);
nor UO_1819 (O_1819,N_24665,N_23536);
or UO_1820 (O_1820,N_24323,N_24957);
nand UO_1821 (O_1821,N_23387,N_24986);
nor UO_1822 (O_1822,N_23602,N_24012);
nand UO_1823 (O_1823,N_22908,N_24704);
or UO_1824 (O_1824,N_24137,N_23010);
or UO_1825 (O_1825,N_22297,N_23275);
nand UO_1826 (O_1826,N_24508,N_22271);
xor UO_1827 (O_1827,N_22711,N_23668);
nor UO_1828 (O_1828,N_23362,N_22797);
or UO_1829 (O_1829,N_22411,N_22552);
nor UO_1830 (O_1830,N_23880,N_22817);
nor UO_1831 (O_1831,N_23904,N_24821);
and UO_1832 (O_1832,N_24902,N_23686);
and UO_1833 (O_1833,N_22001,N_24372);
or UO_1834 (O_1834,N_24455,N_24956);
and UO_1835 (O_1835,N_24949,N_23707);
nand UO_1836 (O_1836,N_22105,N_23371);
or UO_1837 (O_1837,N_22158,N_23471);
nor UO_1838 (O_1838,N_22029,N_23823);
nor UO_1839 (O_1839,N_23696,N_22470);
and UO_1840 (O_1840,N_23047,N_22574);
nand UO_1841 (O_1841,N_22505,N_21908);
and UO_1842 (O_1842,N_22771,N_24916);
and UO_1843 (O_1843,N_23049,N_24094);
or UO_1844 (O_1844,N_22282,N_23587);
and UO_1845 (O_1845,N_22930,N_22986);
nor UO_1846 (O_1846,N_24823,N_23349);
nor UO_1847 (O_1847,N_22241,N_23730);
or UO_1848 (O_1848,N_22582,N_22978);
or UO_1849 (O_1849,N_24117,N_24544);
and UO_1850 (O_1850,N_23332,N_22459);
nand UO_1851 (O_1851,N_22253,N_22959);
xnor UO_1852 (O_1852,N_23324,N_24102);
and UO_1853 (O_1853,N_24788,N_23478);
nand UO_1854 (O_1854,N_23591,N_21963);
or UO_1855 (O_1855,N_24743,N_24439);
nand UO_1856 (O_1856,N_24857,N_23254);
and UO_1857 (O_1857,N_24574,N_22991);
and UO_1858 (O_1858,N_22940,N_24803);
nor UO_1859 (O_1859,N_22699,N_24627);
nor UO_1860 (O_1860,N_24489,N_23957);
nand UO_1861 (O_1861,N_22870,N_24115);
nand UO_1862 (O_1862,N_22531,N_23318);
and UO_1863 (O_1863,N_24003,N_24926);
nand UO_1864 (O_1864,N_22547,N_22316);
nor UO_1865 (O_1865,N_23046,N_22643);
nand UO_1866 (O_1866,N_23654,N_22758);
and UO_1867 (O_1867,N_23921,N_23142);
or UO_1868 (O_1868,N_24930,N_22092);
nand UO_1869 (O_1869,N_24403,N_23838);
nor UO_1870 (O_1870,N_23636,N_22039);
nand UO_1871 (O_1871,N_24007,N_22201);
nand UO_1872 (O_1872,N_23626,N_24469);
nand UO_1873 (O_1873,N_23744,N_23010);
nor UO_1874 (O_1874,N_23009,N_23903);
nand UO_1875 (O_1875,N_24494,N_24811);
and UO_1876 (O_1876,N_24308,N_23629);
xnor UO_1877 (O_1877,N_24769,N_24755);
nor UO_1878 (O_1878,N_23565,N_23337);
xor UO_1879 (O_1879,N_22549,N_22252);
nand UO_1880 (O_1880,N_24972,N_23423);
and UO_1881 (O_1881,N_22219,N_24516);
nor UO_1882 (O_1882,N_22036,N_23337);
nor UO_1883 (O_1883,N_22220,N_23396);
and UO_1884 (O_1884,N_22332,N_24675);
nand UO_1885 (O_1885,N_23297,N_23910);
and UO_1886 (O_1886,N_23915,N_23417);
nor UO_1887 (O_1887,N_22722,N_24535);
xnor UO_1888 (O_1888,N_22116,N_23261);
nand UO_1889 (O_1889,N_23898,N_24406);
xor UO_1890 (O_1890,N_24258,N_23551);
and UO_1891 (O_1891,N_21894,N_23762);
and UO_1892 (O_1892,N_24298,N_22206);
or UO_1893 (O_1893,N_24328,N_24663);
nor UO_1894 (O_1894,N_24897,N_22071);
and UO_1895 (O_1895,N_22393,N_23870);
nor UO_1896 (O_1896,N_22692,N_23680);
and UO_1897 (O_1897,N_24997,N_22701);
xor UO_1898 (O_1898,N_24073,N_23410);
and UO_1899 (O_1899,N_22766,N_23133);
nand UO_1900 (O_1900,N_22828,N_24016);
nand UO_1901 (O_1901,N_22275,N_23455);
and UO_1902 (O_1902,N_21944,N_24090);
and UO_1903 (O_1903,N_24845,N_22127);
or UO_1904 (O_1904,N_24216,N_24761);
nand UO_1905 (O_1905,N_24550,N_23625);
nand UO_1906 (O_1906,N_24036,N_21892);
nand UO_1907 (O_1907,N_22322,N_23538);
and UO_1908 (O_1908,N_22815,N_22974);
and UO_1909 (O_1909,N_24097,N_22663);
and UO_1910 (O_1910,N_23319,N_23967);
nand UO_1911 (O_1911,N_22813,N_24604);
xnor UO_1912 (O_1912,N_24658,N_23933);
or UO_1913 (O_1913,N_24971,N_22077);
and UO_1914 (O_1914,N_24103,N_22788);
nand UO_1915 (O_1915,N_24399,N_23326);
nand UO_1916 (O_1916,N_22196,N_24434);
nor UO_1917 (O_1917,N_23691,N_24661);
and UO_1918 (O_1918,N_22370,N_22239);
nor UO_1919 (O_1919,N_24352,N_24626);
nor UO_1920 (O_1920,N_23827,N_22644);
or UO_1921 (O_1921,N_23308,N_24754);
nor UO_1922 (O_1922,N_24627,N_22385);
nor UO_1923 (O_1923,N_22032,N_23077);
nand UO_1924 (O_1924,N_23146,N_23273);
or UO_1925 (O_1925,N_22961,N_22965);
nand UO_1926 (O_1926,N_23972,N_22659);
and UO_1927 (O_1927,N_22627,N_22269);
xnor UO_1928 (O_1928,N_23244,N_21906);
or UO_1929 (O_1929,N_23698,N_23794);
nand UO_1930 (O_1930,N_23235,N_24992);
nand UO_1931 (O_1931,N_22801,N_24302);
and UO_1932 (O_1932,N_24219,N_23180);
and UO_1933 (O_1933,N_24434,N_24777);
nand UO_1934 (O_1934,N_21952,N_22415);
or UO_1935 (O_1935,N_22107,N_24649);
and UO_1936 (O_1936,N_22039,N_23251);
nand UO_1937 (O_1937,N_23362,N_21978);
or UO_1938 (O_1938,N_24762,N_23704);
nor UO_1939 (O_1939,N_23899,N_24337);
nor UO_1940 (O_1940,N_22153,N_22421);
or UO_1941 (O_1941,N_23134,N_24579);
or UO_1942 (O_1942,N_23000,N_24834);
nor UO_1943 (O_1943,N_24104,N_22971);
nor UO_1944 (O_1944,N_22681,N_22399);
nand UO_1945 (O_1945,N_24975,N_22539);
nor UO_1946 (O_1946,N_24010,N_22897);
nand UO_1947 (O_1947,N_22197,N_22104);
or UO_1948 (O_1948,N_24550,N_24657);
or UO_1949 (O_1949,N_23973,N_23453);
nand UO_1950 (O_1950,N_23915,N_24557);
and UO_1951 (O_1951,N_23153,N_24175);
and UO_1952 (O_1952,N_23346,N_22833);
and UO_1953 (O_1953,N_22796,N_22970);
nor UO_1954 (O_1954,N_23738,N_22208);
nand UO_1955 (O_1955,N_23003,N_24212);
nor UO_1956 (O_1956,N_22084,N_22589);
nor UO_1957 (O_1957,N_22422,N_23536);
xnor UO_1958 (O_1958,N_24974,N_24573);
and UO_1959 (O_1959,N_23861,N_22855);
and UO_1960 (O_1960,N_21876,N_24947);
nand UO_1961 (O_1961,N_23119,N_24581);
nand UO_1962 (O_1962,N_24704,N_22695);
nand UO_1963 (O_1963,N_22504,N_22730);
nand UO_1964 (O_1964,N_22526,N_22740);
and UO_1965 (O_1965,N_23679,N_23585);
or UO_1966 (O_1966,N_22063,N_22224);
and UO_1967 (O_1967,N_22365,N_24789);
nor UO_1968 (O_1968,N_23053,N_23083);
and UO_1969 (O_1969,N_22090,N_24344);
or UO_1970 (O_1970,N_23515,N_23553);
and UO_1971 (O_1971,N_22989,N_23144);
or UO_1972 (O_1972,N_23223,N_23141);
nand UO_1973 (O_1973,N_24987,N_24105);
nand UO_1974 (O_1974,N_23481,N_22861);
nor UO_1975 (O_1975,N_23290,N_23526);
nor UO_1976 (O_1976,N_23951,N_23756);
nand UO_1977 (O_1977,N_24803,N_23921);
nor UO_1978 (O_1978,N_23599,N_24809);
and UO_1979 (O_1979,N_24559,N_24135);
nand UO_1980 (O_1980,N_24469,N_24168);
or UO_1981 (O_1981,N_21904,N_24211);
nor UO_1982 (O_1982,N_23096,N_24358);
and UO_1983 (O_1983,N_24234,N_24091);
or UO_1984 (O_1984,N_24631,N_23472);
and UO_1985 (O_1985,N_24751,N_24602);
xor UO_1986 (O_1986,N_24252,N_24816);
xnor UO_1987 (O_1987,N_24931,N_22056);
and UO_1988 (O_1988,N_22054,N_24574);
nor UO_1989 (O_1989,N_21999,N_24711);
nor UO_1990 (O_1990,N_22108,N_22841);
nor UO_1991 (O_1991,N_23363,N_22259);
and UO_1992 (O_1992,N_23861,N_24062);
and UO_1993 (O_1993,N_22030,N_23201);
or UO_1994 (O_1994,N_24451,N_24765);
nor UO_1995 (O_1995,N_23049,N_22514);
nor UO_1996 (O_1996,N_22729,N_24810);
or UO_1997 (O_1997,N_22188,N_24147);
or UO_1998 (O_1998,N_23442,N_23647);
nand UO_1999 (O_1999,N_24248,N_23240);
nor UO_2000 (O_2000,N_22608,N_22209);
or UO_2001 (O_2001,N_24851,N_23698);
nand UO_2002 (O_2002,N_22429,N_23537);
nor UO_2003 (O_2003,N_23508,N_24344);
or UO_2004 (O_2004,N_22598,N_22875);
and UO_2005 (O_2005,N_24897,N_23121);
nand UO_2006 (O_2006,N_24649,N_22363);
xor UO_2007 (O_2007,N_24029,N_21952);
or UO_2008 (O_2008,N_23306,N_24126);
nand UO_2009 (O_2009,N_24642,N_23245);
and UO_2010 (O_2010,N_24818,N_23094);
and UO_2011 (O_2011,N_22381,N_24243);
nand UO_2012 (O_2012,N_24073,N_24178);
nor UO_2013 (O_2013,N_22504,N_22079);
and UO_2014 (O_2014,N_22805,N_23263);
nand UO_2015 (O_2015,N_23302,N_21993);
nor UO_2016 (O_2016,N_22179,N_24145);
nor UO_2017 (O_2017,N_23686,N_24761);
or UO_2018 (O_2018,N_24617,N_24682);
or UO_2019 (O_2019,N_22892,N_24982);
nor UO_2020 (O_2020,N_22723,N_23740);
nor UO_2021 (O_2021,N_22373,N_23929);
or UO_2022 (O_2022,N_23963,N_24834);
or UO_2023 (O_2023,N_22902,N_22716);
and UO_2024 (O_2024,N_24862,N_22843);
and UO_2025 (O_2025,N_23782,N_23508);
nor UO_2026 (O_2026,N_23319,N_22686);
or UO_2027 (O_2027,N_22459,N_24084);
nand UO_2028 (O_2028,N_22300,N_23090);
nand UO_2029 (O_2029,N_23536,N_23676);
xor UO_2030 (O_2030,N_23833,N_22093);
or UO_2031 (O_2031,N_22055,N_24872);
nand UO_2032 (O_2032,N_24275,N_24604);
nand UO_2033 (O_2033,N_23991,N_24497);
xor UO_2034 (O_2034,N_23989,N_22626);
and UO_2035 (O_2035,N_24660,N_22420);
nor UO_2036 (O_2036,N_23945,N_23703);
nor UO_2037 (O_2037,N_23979,N_24337);
or UO_2038 (O_2038,N_24918,N_24977);
xor UO_2039 (O_2039,N_24888,N_24984);
nand UO_2040 (O_2040,N_22826,N_21973);
nor UO_2041 (O_2041,N_23973,N_22492);
nand UO_2042 (O_2042,N_24886,N_23361);
and UO_2043 (O_2043,N_22828,N_24699);
or UO_2044 (O_2044,N_23318,N_22211);
or UO_2045 (O_2045,N_24468,N_22151);
nand UO_2046 (O_2046,N_23598,N_23913);
nor UO_2047 (O_2047,N_22643,N_22674);
nor UO_2048 (O_2048,N_23433,N_23875);
and UO_2049 (O_2049,N_23193,N_22917);
xor UO_2050 (O_2050,N_22838,N_22126);
nor UO_2051 (O_2051,N_23837,N_22119);
nor UO_2052 (O_2052,N_23947,N_22809);
nor UO_2053 (O_2053,N_24842,N_22559);
and UO_2054 (O_2054,N_22963,N_23403);
nor UO_2055 (O_2055,N_24762,N_23168);
nand UO_2056 (O_2056,N_24765,N_24797);
nand UO_2057 (O_2057,N_23597,N_24340);
and UO_2058 (O_2058,N_24297,N_23579);
and UO_2059 (O_2059,N_24431,N_23445);
and UO_2060 (O_2060,N_23011,N_24568);
nor UO_2061 (O_2061,N_22379,N_24433);
nand UO_2062 (O_2062,N_23295,N_23061);
or UO_2063 (O_2063,N_23299,N_24540);
and UO_2064 (O_2064,N_22811,N_24566);
nand UO_2065 (O_2065,N_24480,N_23500);
nand UO_2066 (O_2066,N_24761,N_24770);
nand UO_2067 (O_2067,N_24606,N_24643);
or UO_2068 (O_2068,N_24303,N_22961);
nand UO_2069 (O_2069,N_22820,N_23773);
and UO_2070 (O_2070,N_23220,N_24477);
nand UO_2071 (O_2071,N_23256,N_21914);
nor UO_2072 (O_2072,N_22092,N_21999);
or UO_2073 (O_2073,N_24571,N_22687);
nand UO_2074 (O_2074,N_22942,N_23384);
nor UO_2075 (O_2075,N_24104,N_23534);
or UO_2076 (O_2076,N_23404,N_22567);
or UO_2077 (O_2077,N_22447,N_22472);
or UO_2078 (O_2078,N_24138,N_22272);
nor UO_2079 (O_2079,N_22315,N_22862);
nor UO_2080 (O_2080,N_22060,N_23193);
xnor UO_2081 (O_2081,N_24051,N_24453);
and UO_2082 (O_2082,N_23305,N_24634);
xnor UO_2083 (O_2083,N_22612,N_24284);
xnor UO_2084 (O_2084,N_23686,N_21947);
xnor UO_2085 (O_2085,N_24407,N_24770);
or UO_2086 (O_2086,N_23627,N_24027);
and UO_2087 (O_2087,N_23714,N_23431);
nor UO_2088 (O_2088,N_24449,N_24320);
nor UO_2089 (O_2089,N_22023,N_24334);
or UO_2090 (O_2090,N_23982,N_24175);
and UO_2091 (O_2091,N_23235,N_24472);
or UO_2092 (O_2092,N_23137,N_23256);
nor UO_2093 (O_2093,N_24077,N_22711);
and UO_2094 (O_2094,N_22156,N_22445);
nor UO_2095 (O_2095,N_24161,N_22446);
nor UO_2096 (O_2096,N_22033,N_24011);
or UO_2097 (O_2097,N_22505,N_23019);
or UO_2098 (O_2098,N_24274,N_23466);
xnor UO_2099 (O_2099,N_24624,N_24630);
nand UO_2100 (O_2100,N_22421,N_24561);
and UO_2101 (O_2101,N_22348,N_24028);
nor UO_2102 (O_2102,N_22228,N_22324);
or UO_2103 (O_2103,N_22630,N_23788);
and UO_2104 (O_2104,N_24410,N_24024);
and UO_2105 (O_2105,N_23704,N_22663);
and UO_2106 (O_2106,N_24576,N_24734);
or UO_2107 (O_2107,N_22939,N_24918);
nand UO_2108 (O_2108,N_24229,N_23529);
xor UO_2109 (O_2109,N_24635,N_21918);
and UO_2110 (O_2110,N_22056,N_23035);
and UO_2111 (O_2111,N_24165,N_22182);
nand UO_2112 (O_2112,N_21905,N_22187);
nand UO_2113 (O_2113,N_24050,N_24911);
nor UO_2114 (O_2114,N_22747,N_23196);
or UO_2115 (O_2115,N_23386,N_23660);
or UO_2116 (O_2116,N_22034,N_23972);
nor UO_2117 (O_2117,N_23240,N_22875);
and UO_2118 (O_2118,N_24731,N_22584);
and UO_2119 (O_2119,N_21997,N_24557);
nand UO_2120 (O_2120,N_22639,N_22087);
and UO_2121 (O_2121,N_22498,N_23026);
xor UO_2122 (O_2122,N_24507,N_24715);
nor UO_2123 (O_2123,N_22463,N_23183);
and UO_2124 (O_2124,N_23808,N_24828);
nor UO_2125 (O_2125,N_24836,N_22422);
or UO_2126 (O_2126,N_23540,N_22078);
or UO_2127 (O_2127,N_22756,N_24641);
or UO_2128 (O_2128,N_22795,N_23189);
or UO_2129 (O_2129,N_24466,N_22791);
nor UO_2130 (O_2130,N_21917,N_22010);
and UO_2131 (O_2131,N_24621,N_24554);
or UO_2132 (O_2132,N_24773,N_22523);
xor UO_2133 (O_2133,N_22326,N_24331);
and UO_2134 (O_2134,N_24301,N_23010);
or UO_2135 (O_2135,N_24466,N_22422);
and UO_2136 (O_2136,N_24509,N_24900);
and UO_2137 (O_2137,N_23037,N_24314);
nor UO_2138 (O_2138,N_24916,N_24664);
nor UO_2139 (O_2139,N_24602,N_23285);
and UO_2140 (O_2140,N_24365,N_24446);
or UO_2141 (O_2141,N_22765,N_23202);
or UO_2142 (O_2142,N_24446,N_23778);
or UO_2143 (O_2143,N_22660,N_22643);
and UO_2144 (O_2144,N_24441,N_24870);
and UO_2145 (O_2145,N_24966,N_23240);
nor UO_2146 (O_2146,N_23908,N_23708);
nand UO_2147 (O_2147,N_23898,N_23646);
nand UO_2148 (O_2148,N_24132,N_22381);
and UO_2149 (O_2149,N_22370,N_23842);
or UO_2150 (O_2150,N_24584,N_24571);
or UO_2151 (O_2151,N_24004,N_22452);
nand UO_2152 (O_2152,N_23202,N_23284);
nand UO_2153 (O_2153,N_23394,N_21878);
and UO_2154 (O_2154,N_23766,N_24194);
and UO_2155 (O_2155,N_24924,N_23682);
and UO_2156 (O_2156,N_24843,N_23152);
and UO_2157 (O_2157,N_22861,N_21989);
nand UO_2158 (O_2158,N_22766,N_22990);
nor UO_2159 (O_2159,N_22497,N_23380);
or UO_2160 (O_2160,N_24170,N_23893);
nand UO_2161 (O_2161,N_24575,N_23568);
and UO_2162 (O_2162,N_22744,N_24346);
and UO_2163 (O_2163,N_24660,N_24956);
xor UO_2164 (O_2164,N_23153,N_22286);
and UO_2165 (O_2165,N_24606,N_24425);
nor UO_2166 (O_2166,N_22301,N_22514);
and UO_2167 (O_2167,N_24972,N_21900);
nor UO_2168 (O_2168,N_24371,N_23850);
and UO_2169 (O_2169,N_23013,N_23440);
nand UO_2170 (O_2170,N_22008,N_22425);
nand UO_2171 (O_2171,N_24487,N_23156);
and UO_2172 (O_2172,N_24354,N_22386);
and UO_2173 (O_2173,N_23352,N_22509);
or UO_2174 (O_2174,N_22656,N_23359);
nor UO_2175 (O_2175,N_22196,N_24394);
and UO_2176 (O_2176,N_24518,N_24418);
and UO_2177 (O_2177,N_23677,N_24120);
and UO_2178 (O_2178,N_22708,N_24291);
and UO_2179 (O_2179,N_23138,N_22191);
nand UO_2180 (O_2180,N_22004,N_23881);
nand UO_2181 (O_2181,N_21955,N_23262);
nand UO_2182 (O_2182,N_24911,N_24667);
nand UO_2183 (O_2183,N_23714,N_24468);
nor UO_2184 (O_2184,N_24507,N_24738);
and UO_2185 (O_2185,N_23635,N_23996);
nor UO_2186 (O_2186,N_23455,N_23074);
or UO_2187 (O_2187,N_24093,N_23817);
or UO_2188 (O_2188,N_24367,N_22599);
or UO_2189 (O_2189,N_22051,N_22269);
xor UO_2190 (O_2190,N_23169,N_24894);
nor UO_2191 (O_2191,N_23978,N_23894);
xor UO_2192 (O_2192,N_24567,N_24455);
and UO_2193 (O_2193,N_23877,N_23056);
and UO_2194 (O_2194,N_22701,N_24921);
or UO_2195 (O_2195,N_23560,N_23166);
nand UO_2196 (O_2196,N_24176,N_24366);
nor UO_2197 (O_2197,N_24407,N_22638);
nor UO_2198 (O_2198,N_22495,N_24339);
nor UO_2199 (O_2199,N_22482,N_22132);
xnor UO_2200 (O_2200,N_23123,N_22692);
and UO_2201 (O_2201,N_23282,N_24241);
nor UO_2202 (O_2202,N_24037,N_23930);
and UO_2203 (O_2203,N_22116,N_23320);
and UO_2204 (O_2204,N_24559,N_22298);
xnor UO_2205 (O_2205,N_23083,N_22963);
and UO_2206 (O_2206,N_23634,N_22030);
nor UO_2207 (O_2207,N_24280,N_24705);
nand UO_2208 (O_2208,N_23663,N_24559);
and UO_2209 (O_2209,N_23554,N_23296);
nand UO_2210 (O_2210,N_24437,N_24187);
nand UO_2211 (O_2211,N_22725,N_24304);
nand UO_2212 (O_2212,N_24343,N_24101);
or UO_2213 (O_2213,N_24544,N_22121);
and UO_2214 (O_2214,N_22131,N_23360);
or UO_2215 (O_2215,N_23631,N_23783);
nand UO_2216 (O_2216,N_22765,N_23357);
and UO_2217 (O_2217,N_22708,N_22784);
nor UO_2218 (O_2218,N_23941,N_22085);
xnor UO_2219 (O_2219,N_22113,N_23602);
and UO_2220 (O_2220,N_23015,N_22468);
and UO_2221 (O_2221,N_23565,N_24559);
and UO_2222 (O_2222,N_22856,N_24277);
nand UO_2223 (O_2223,N_22223,N_24702);
or UO_2224 (O_2224,N_23239,N_24741);
and UO_2225 (O_2225,N_24129,N_22366);
xnor UO_2226 (O_2226,N_23331,N_24660);
and UO_2227 (O_2227,N_24415,N_22119);
nor UO_2228 (O_2228,N_21944,N_24796);
or UO_2229 (O_2229,N_21991,N_22970);
or UO_2230 (O_2230,N_24101,N_22975);
and UO_2231 (O_2231,N_22204,N_23542);
nor UO_2232 (O_2232,N_22435,N_23185);
xnor UO_2233 (O_2233,N_23069,N_24102);
nor UO_2234 (O_2234,N_22648,N_23916);
nand UO_2235 (O_2235,N_22249,N_24648);
nand UO_2236 (O_2236,N_22055,N_24208);
xnor UO_2237 (O_2237,N_23393,N_22102);
or UO_2238 (O_2238,N_23577,N_23307);
nor UO_2239 (O_2239,N_22270,N_23787);
nand UO_2240 (O_2240,N_24188,N_23002);
and UO_2241 (O_2241,N_22201,N_23561);
and UO_2242 (O_2242,N_24698,N_24738);
nor UO_2243 (O_2243,N_21978,N_23277);
xor UO_2244 (O_2244,N_22139,N_24033);
nand UO_2245 (O_2245,N_23877,N_21958);
nor UO_2246 (O_2246,N_21935,N_24740);
and UO_2247 (O_2247,N_22919,N_24164);
and UO_2248 (O_2248,N_21889,N_22840);
and UO_2249 (O_2249,N_22816,N_22663);
and UO_2250 (O_2250,N_21935,N_24268);
nor UO_2251 (O_2251,N_22210,N_22028);
and UO_2252 (O_2252,N_24578,N_24447);
nor UO_2253 (O_2253,N_22637,N_24859);
nor UO_2254 (O_2254,N_24680,N_23038);
or UO_2255 (O_2255,N_24168,N_22034);
and UO_2256 (O_2256,N_24381,N_24047);
and UO_2257 (O_2257,N_23585,N_24892);
and UO_2258 (O_2258,N_24409,N_23900);
nor UO_2259 (O_2259,N_22322,N_22877);
or UO_2260 (O_2260,N_23241,N_21961);
xnor UO_2261 (O_2261,N_24830,N_22278);
nand UO_2262 (O_2262,N_23109,N_23320);
nor UO_2263 (O_2263,N_24218,N_22343);
nand UO_2264 (O_2264,N_24747,N_23891);
and UO_2265 (O_2265,N_24088,N_24643);
nand UO_2266 (O_2266,N_22778,N_23394);
and UO_2267 (O_2267,N_22832,N_24617);
and UO_2268 (O_2268,N_23969,N_22532);
xor UO_2269 (O_2269,N_23038,N_23569);
xor UO_2270 (O_2270,N_23278,N_24298);
or UO_2271 (O_2271,N_24827,N_22130);
xnor UO_2272 (O_2272,N_22301,N_22098);
or UO_2273 (O_2273,N_22467,N_24160);
nand UO_2274 (O_2274,N_22002,N_23313);
nor UO_2275 (O_2275,N_22835,N_23214);
xor UO_2276 (O_2276,N_24467,N_24578);
or UO_2277 (O_2277,N_23560,N_24093);
nand UO_2278 (O_2278,N_23838,N_22285);
or UO_2279 (O_2279,N_24513,N_23665);
and UO_2280 (O_2280,N_24686,N_22804);
nand UO_2281 (O_2281,N_24165,N_22927);
nor UO_2282 (O_2282,N_22233,N_22214);
nand UO_2283 (O_2283,N_24648,N_24254);
and UO_2284 (O_2284,N_23807,N_24179);
and UO_2285 (O_2285,N_22784,N_22102);
or UO_2286 (O_2286,N_22765,N_24012);
and UO_2287 (O_2287,N_23610,N_22352);
xor UO_2288 (O_2288,N_24163,N_24964);
and UO_2289 (O_2289,N_21989,N_23230);
nand UO_2290 (O_2290,N_21935,N_23525);
or UO_2291 (O_2291,N_24164,N_22953);
nand UO_2292 (O_2292,N_24746,N_22638);
nand UO_2293 (O_2293,N_24542,N_23255);
nand UO_2294 (O_2294,N_23922,N_23025);
xnor UO_2295 (O_2295,N_23628,N_22798);
or UO_2296 (O_2296,N_22342,N_22305);
or UO_2297 (O_2297,N_24569,N_22898);
or UO_2298 (O_2298,N_22021,N_22058);
nor UO_2299 (O_2299,N_24918,N_22313);
xor UO_2300 (O_2300,N_23180,N_24414);
nand UO_2301 (O_2301,N_22026,N_24702);
nor UO_2302 (O_2302,N_22582,N_23037);
xor UO_2303 (O_2303,N_24476,N_24019);
nand UO_2304 (O_2304,N_22101,N_22285);
nand UO_2305 (O_2305,N_22278,N_22694);
nor UO_2306 (O_2306,N_22190,N_22143);
or UO_2307 (O_2307,N_23627,N_23494);
and UO_2308 (O_2308,N_24931,N_24407);
nand UO_2309 (O_2309,N_24888,N_23857);
nor UO_2310 (O_2310,N_24494,N_22227);
nor UO_2311 (O_2311,N_22416,N_23843);
nand UO_2312 (O_2312,N_24282,N_23758);
or UO_2313 (O_2313,N_23877,N_22441);
nand UO_2314 (O_2314,N_24927,N_24109);
or UO_2315 (O_2315,N_22026,N_22206);
or UO_2316 (O_2316,N_22385,N_23987);
xor UO_2317 (O_2317,N_23376,N_23428);
and UO_2318 (O_2318,N_21938,N_24348);
or UO_2319 (O_2319,N_22101,N_24784);
nand UO_2320 (O_2320,N_22644,N_24341);
and UO_2321 (O_2321,N_22027,N_23766);
nor UO_2322 (O_2322,N_24068,N_24011);
nor UO_2323 (O_2323,N_24665,N_23614);
or UO_2324 (O_2324,N_24267,N_22058);
nor UO_2325 (O_2325,N_22316,N_24287);
xor UO_2326 (O_2326,N_22038,N_24711);
nor UO_2327 (O_2327,N_22483,N_21926);
nor UO_2328 (O_2328,N_24870,N_24020);
nor UO_2329 (O_2329,N_22638,N_24408);
or UO_2330 (O_2330,N_24580,N_24133);
xnor UO_2331 (O_2331,N_22187,N_23549);
or UO_2332 (O_2332,N_23674,N_22786);
and UO_2333 (O_2333,N_23310,N_23524);
and UO_2334 (O_2334,N_23612,N_24232);
nor UO_2335 (O_2335,N_22535,N_24325);
nand UO_2336 (O_2336,N_23261,N_23975);
and UO_2337 (O_2337,N_22993,N_23028);
nor UO_2338 (O_2338,N_21985,N_24836);
nand UO_2339 (O_2339,N_22036,N_24745);
or UO_2340 (O_2340,N_24226,N_24480);
and UO_2341 (O_2341,N_24777,N_22432);
and UO_2342 (O_2342,N_24329,N_23587);
and UO_2343 (O_2343,N_24595,N_24598);
nor UO_2344 (O_2344,N_24365,N_23954);
or UO_2345 (O_2345,N_24139,N_24973);
nand UO_2346 (O_2346,N_24731,N_22019);
nor UO_2347 (O_2347,N_23420,N_23945);
nor UO_2348 (O_2348,N_24026,N_23208);
or UO_2349 (O_2349,N_24247,N_24026);
nor UO_2350 (O_2350,N_24689,N_23410);
nand UO_2351 (O_2351,N_24494,N_22849);
and UO_2352 (O_2352,N_23025,N_22128);
xor UO_2353 (O_2353,N_22794,N_22857);
or UO_2354 (O_2354,N_23227,N_22224);
and UO_2355 (O_2355,N_22907,N_22541);
xnor UO_2356 (O_2356,N_24958,N_22388);
or UO_2357 (O_2357,N_22416,N_22103);
nor UO_2358 (O_2358,N_24598,N_22460);
and UO_2359 (O_2359,N_23471,N_23618);
or UO_2360 (O_2360,N_23696,N_22997);
and UO_2361 (O_2361,N_23364,N_22026);
and UO_2362 (O_2362,N_22894,N_22775);
and UO_2363 (O_2363,N_22200,N_24103);
nand UO_2364 (O_2364,N_22649,N_22228);
and UO_2365 (O_2365,N_23672,N_24461);
nand UO_2366 (O_2366,N_23423,N_24323);
nor UO_2367 (O_2367,N_23566,N_23839);
nor UO_2368 (O_2368,N_23809,N_24891);
and UO_2369 (O_2369,N_23816,N_23773);
nor UO_2370 (O_2370,N_23786,N_22856);
or UO_2371 (O_2371,N_24371,N_23031);
nand UO_2372 (O_2372,N_22086,N_22919);
nand UO_2373 (O_2373,N_24169,N_23167);
xnor UO_2374 (O_2374,N_22933,N_24433);
nor UO_2375 (O_2375,N_22477,N_21905);
nor UO_2376 (O_2376,N_23169,N_22092);
and UO_2377 (O_2377,N_22523,N_24578);
nand UO_2378 (O_2378,N_23270,N_23967);
and UO_2379 (O_2379,N_23454,N_23386);
or UO_2380 (O_2380,N_21890,N_22685);
nor UO_2381 (O_2381,N_22673,N_22553);
nand UO_2382 (O_2382,N_23930,N_22023);
xor UO_2383 (O_2383,N_22818,N_23585);
and UO_2384 (O_2384,N_24401,N_22131);
nor UO_2385 (O_2385,N_24423,N_24723);
nor UO_2386 (O_2386,N_22857,N_22497);
nand UO_2387 (O_2387,N_23148,N_22770);
nor UO_2388 (O_2388,N_22294,N_23718);
nand UO_2389 (O_2389,N_22005,N_24996);
nor UO_2390 (O_2390,N_23543,N_24980);
or UO_2391 (O_2391,N_24620,N_22933);
nand UO_2392 (O_2392,N_24840,N_22861);
nand UO_2393 (O_2393,N_23824,N_23453);
nor UO_2394 (O_2394,N_24317,N_22891);
and UO_2395 (O_2395,N_22610,N_22603);
nor UO_2396 (O_2396,N_23162,N_24824);
nand UO_2397 (O_2397,N_23887,N_24124);
nand UO_2398 (O_2398,N_24469,N_24829);
or UO_2399 (O_2399,N_24744,N_22975);
nor UO_2400 (O_2400,N_22682,N_24595);
nor UO_2401 (O_2401,N_23920,N_23876);
or UO_2402 (O_2402,N_22679,N_22416);
nand UO_2403 (O_2403,N_23728,N_22396);
xnor UO_2404 (O_2404,N_24126,N_22679);
nor UO_2405 (O_2405,N_23606,N_24629);
or UO_2406 (O_2406,N_22181,N_22377);
nand UO_2407 (O_2407,N_22479,N_22212);
xnor UO_2408 (O_2408,N_22755,N_24739);
nand UO_2409 (O_2409,N_24669,N_24267);
xor UO_2410 (O_2410,N_24455,N_24784);
or UO_2411 (O_2411,N_24937,N_23870);
or UO_2412 (O_2412,N_22375,N_23075);
and UO_2413 (O_2413,N_24667,N_24793);
nor UO_2414 (O_2414,N_21923,N_22310);
and UO_2415 (O_2415,N_23322,N_24633);
nand UO_2416 (O_2416,N_24047,N_23287);
nand UO_2417 (O_2417,N_23924,N_22130);
nor UO_2418 (O_2418,N_24790,N_23284);
and UO_2419 (O_2419,N_24732,N_24985);
or UO_2420 (O_2420,N_21964,N_23003);
or UO_2421 (O_2421,N_23625,N_23413);
or UO_2422 (O_2422,N_22512,N_24820);
or UO_2423 (O_2423,N_22117,N_24919);
and UO_2424 (O_2424,N_24727,N_22860);
nand UO_2425 (O_2425,N_24276,N_22585);
nand UO_2426 (O_2426,N_23408,N_22326);
or UO_2427 (O_2427,N_21882,N_22626);
and UO_2428 (O_2428,N_24131,N_23834);
nand UO_2429 (O_2429,N_23110,N_23851);
nand UO_2430 (O_2430,N_24924,N_22704);
or UO_2431 (O_2431,N_24842,N_22481);
nand UO_2432 (O_2432,N_24333,N_23265);
and UO_2433 (O_2433,N_22472,N_23440);
nand UO_2434 (O_2434,N_22264,N_22189);
nor UO_2435 (O_2435,N_22222,N_22801);
or UO_2436 (O_2436,N_23734,N_22667);
nand UO_2437 (O_2437,N_22579,N_23328);
nand UO_2438 (O_2438,N_23003,N_24331);
xor UO_2439 (O_2439,N_22629,N_23289);
nand UO_2440 (O_2440,N_22114,N_23784);
nor UO_2441 (O_2441,N_22191,N_23405);
or UO_2442 (O_2442,N_24995,N_22442);
xor UO_2443 (O_2443,N_24001,N_21889);
or UO_2444 (O_2444,N_24785,N_22282);
nor UO_2445 (O_2445,N_24692,N_22694);
nor UO_2446 (O_2446,N_24244,N_24504);
nand UO_2447 (O_2447,N_23041,N_23286);
nor UO_2448 (O_2448,N_24065,N_22855);
and UO_2449 (O_2449,N_24522,N_24674);
nor UO_2450 (O_2450,N_24290,N_24303);
xnor UO_2451 (O_2451,N_24945,N_23217);
or UO_2452 (O_2452,N_22231,N_24167);
nand UO_2453 (O_2453,N_23619,N_22914);
nor UO_2454 (O_2454,N_24627,N_22801);
and UO_2455 (O_2455,N_23565,N_23881);
and UO_2456 (O_2456,N_22020,N_23686);
and UO_2457 (O_2457,N_24024,N_24189);
nand UO_2458 (O_2458,N_22367,N_21977);
nor UO_2459 (O_2459,N_22563,N_22687);
xor UO_2460 (O_2460,N_24518,N_22692);
nor UO_2461 (O_2461,N_23972,N_24780);
nor UO_2462 (O_2462,N_24163,N_22987);
nand UO_2463 (O_2463,N_22636,N_23257);
nor UO_2464 (O_2464,N_22603,N_23782);
and UO_2465 (O_2465,N_23274,N_23943);
nor UO_2466 (O_2466,N_24040,N_22353);
nor UO_2467 (O_2467,N_22149,N_23633);
and UO_2468 (O_2468,N_22219,N_24247);
nand UO_2469 (O_2469,N_23198,N_24667);
xnor UO_2470 (O_2470,N_22552,N_21953);
xnor UO_2471 (O_2471,N_22577,N_23399);
or UO_2472 (O_2472,N_24566,N_24254);
nor UO_2473 (O_2473,N_22331,N_22377);
nor UO_2474 (O_2474,N_24358,N_23877);
and UO_2475 (O_2475,N_24532,N_22667);
nand UO_2476 (O_2476,N_24810,N_24310);
or UO_2477 (O_2477,N_24600,N_22836);
nand UO_2478 (O_2478,N_24612,N_23561);
or UO_2479 (O_2479,N_22962,N_24021);
xor UO_2480 (O_2480,N_22461,N_22888);
nand UO_2481 (O_2481,N_22464,N_23997);
nor UO_2482 (O_2482,N_24767,N_24397);
and UO_2483 (O_2483,N_24205,N_22589);
or UO_2484 (O_2484,N_23868,N_23851);
nand UO_2485 (O_2485,N_24692,N_22519);
and UO_2486 (O_2486,N_24740,N_23569);
or UO_2487 (O_2487,N_24913,N_22804);
nor UO_2488 (O_2488,N_24222,N_24908);
or UO_2489 (O_2489,N_23065,N_22742);
nand UO_2490 (O_2490,N_24993,N_24856);
nand UO_2491 (O_2491,N_22784,N_22910);
or UO_2492 (O_2492,N_23047,N_23238);
or UO_2493 (O_2493,N_22516,N_21930);
and UO_2494 (O_2494,N_22696,N_24584);
nor UO_2495 (O_2495,N_24343,N_22326);
nand UO_2496 (O_2496,N_22975,N_24244);
and UO_2497 (O_2497,N_23604,N_22326);
and UO_2498 (O_2498,N_24765,N_23957);
nor UO_2499 (O_2499,N_24832,N_23065);
and UO_2500 (O_2500,N_24330,N_23515);
and UO_2501 (O_2501,N_24974,N_24097);
xor UO_2502 (O_2502,N_21972,N_21875);
or UO_2503 (O_2503,N_23767,N_21876);
and UO_2504 (O_2504,N_22261,N_23069);
and UO_2505 (O_2505,N_21895,N_24403);
nor UO_2506 (O_2506,N_22914,N_23773);
and UO_2507 (O_2507,N_24479,N_22574);
nor UO_2508 (O_2508,N_22858,N_22604);
and UO_2509 (O_2509,N_24264,N_24241);
or UO_2510 (O_2510,N_22371,N_22191);
nand UO_2511 (O_2511,N_23976,N_23343);
nand UO_2512 (O_2512,N_24240,N_23217);
nor UO_2513 (O_2513,N_24030,N_23680);
and UO_2514 (O_2514,N_24057,N_22529);
xor UO_2515 (O_2515,N_23520,N_22434);
xor UO_2516 (O_2516,N_22538,N_22493);
and UO_2517 (O_2517,N_24501,N_23025);
and UO_2518 (O_2518,N_23315,N_24524);
nor UO_2519 (O_2519,N_22403,N_21926);
and UO_2520 (O_2520,N_22398,N_24286);
nor UO_2521 (O_2521,N_24283,N_22116);
nor UO_2522 (O_2522,N_23823,N_22187);
nand UO_2523 (O_2523,N_22746,N_23160);
nand UO_2524 (O_2524,N_23374,N_23284);
xnor UO_2525 (O_2525,N_22217,N_23605);
and UO_2526 (O_2526,N_22987,N_22785);
and UO_2527 (O_2527,N_24106,N_24071);
xnor UO_2528 (O_2528,N_23421,N_23298);
and UO_2529 (O_2529,N_21957,N_22518);
and UO_2530 (O_2530,N_23268,N_24287);
or UO_2531 (O_2531,N_24246,N_22923);
and UO_2532 (O_2532,N_24375,N_22057);
nand UO_2533 (O_2533,N_24743,N_22250);
and UO_2534 (O_2534,N_22210,N_23985);
and UO_2535 (O_2535,N_24108,N_22684);
nand UO_2536 (O_2536,N_24473,N_22607);
nand UO_2537 (O_2537,N_23549,N_23275);
and UO_2538 (O_2538,N_24417,N_21890);
nor UO_2539 (O_2539,N_22484,N_23934);
nor UO_2540 (O_2540,N_24820,N_22215);
or UO_2541 (O_2541,N_24397,N_22268);
nand UO_2542 (O_2542,N_23100,N_23740);
and UO_2543 (O_2543,N_24190,N_23472);
and UO_2544 (O_2544,N_24643,N_21995);
and UO_2545 (O_2545,N_22744,N_22022);
and UO_2546 (O_2546,N_24271,N_24120);
and UO_2547 (O_2547,N_22776,N_24146);
nor UO_2548 (O_2548,N_23842,N_24050);
nand UO_2549 (O_2549,N_24814,N_23109);
xor UO_2550 (O_2550,N_21958,N_24787);
nor UO_2551 (O_2551,N_23055,N_22779);
and UO_2552 (O_2552,N_22070,N_22841);
nand UO_2553 (O_2553,N_22818,N_23589);
nor UO_2554 (O_2554,N_24929,N_23238);
or UO_2555 (O_2555,N_24798,N_21944);
xor UO_2556 (O_2556,N_23250,N_24883);
and UO_2557 (O_2557,N_23069,N_23302);
xnor UO_2558 (O_2558,N_22031,N_22430);
xor UO_2559 (O_2559,N_22636,N_22355);
xor UO_2560 (O_2560,N_24014,N_23798);
and UO_2561 (O_2561,N_22632,N_22149);
nor UO_2562 (O_2562,N_24636,N_24765);
xor UO_2563 (O_2563,N_24671,N_22775);
nand UO_2564 (O_2564,N_24618,N_22179);
and UO_2565 (O_2565,N_24606,N_23735);
nor UO_2566 (O_2566,N_23211,N_21929);
or UO_2567 (O_2567,N_24141,N_23724);
nand UO_2568 (O_2568,N_24957,N_24213);
nor UO_2569 (O_2569,N_23492,N_23121);
or UO_2570 (O_2570,N_23474,N_23753);
nand UO_2571 (O_2571,N_24717,N_22377);
and UO_2572 (O_2572,N_22691,N_22866);
xor UO_2573 (O_2573,N_24813,N_24057);
nor UO_2574 (O_2574,N_22902,N_24284);
nand UO_2575 (O_2575,N_22953,N_21895);
and UO_2576 (O_2576,N_24568,N_24672);
nor UO_2577 (O_2577,N_23641,N_22170);
and UO_2578 (O_2578,N_22733,N_24089);
xnor UO_2579 (O_2579,N_23428,N_22727);
and UO_2580 (O_2580,N_22434,N_22677);
nand UO_2581 (O_2581,N_24172,N_22691);
nand UO_2582 (O_2582,N_22524,N_22678);
or UO_2583 (O_2583,N_22950,N_23010);
nor UO_2584 (O_2584,N_24398,N_24300);
nand UO_2585 (O_2585,N_23166,N_23813);
and UO_2586 (O_2586,N_24400,N_24892);
or UO_2587 (O_2587,N_21970,N_24641);
nor UO_2588 (O_2588,N_23190,N_22801);
nor UO_2589 (O_2589,N_22047,N_22033);
or UO_2590 (O_2590,N_24190,N_22570);
and UO_2591 (O_2591,N_23774,N_24724);
nand UO_2592 (O_2592,N_24695,N_22413);
and UO_2593 (O_2593,N_23580,N_24387);
nor UO_2594 (O_2594,N_23913,N_22559);
nand UO_2595 (O_2595,N_23312,N_24575);
nor UO_2596 (O_2596,N_22338,N_24270);
xor UO_2597 (O_2597,N_22515,N_22112);
nor UO_2598 (O_2598,N_24883,N_23102);
and UO_2599 (O_2599,N_22487,N_24611);
or UO_2600 (O_2600,N_23933,N_23678);
or UO_2601 (O_2601,N_23818,N_22472);
xnor UO_2602 (O_2602,N_24421,N_22753);
nand UO_2603 (O_2603,N_23073,N_22155);
and UO_2604 (O_2604,N_23569,N_24043);
nor UO_2605 (O_2605,N_23860,N_22477);
nor UO_2606 (O_2606,N_23367,N_23440);
nor UO_2607 (O_2607,N_23544,N_22362);
nand UO_2608 (O_2608,N_21891,N_23999);
nor UO_2609 (O_2609,N_24070,N_23511);
and UO_2610 (O_2610,N_23860,N_22241);
xor UO_2611 (O_2611,N_24053,N_23984);
nor UO_2612 (O_2612,N_22461,N_24768);
or UO_2613 (O_2613,N_23550,N_23989);
nor UO_2614 (O_2614,N_22450,N_23777);
nand UO_2615 (O_2615,N_24441,N_22011);
and UO_2616 (O_2616,N_22238,N_22113);
nor UO_2617 (O_2617,N_24739,N_24574);
nor UO_2618 (O_2618,N_23948,N_22682);
or UO_2619 (O_2619,N_22501,N_22600);
nor UO_2620 (O_2620,N_22596,N_24261);
and UO_2621 (O_2621,N_24568,N_24015);
nor UO_2622 (O_2622,N_23950,N_22301);
nand UO_2623 (O_2623,N_22820,N_22623);
or UO_2624 (O_2624,N_24426,N_22657);
and UO_2625 (O_2625,N_22476,N_24910);
nor UO_2626 (O_2626,N_23210,N_24689);
nor UO_2627 (O_2627,N_23939,N_23745);
nand UO_2628 (O_2628,N_21919,N_24308);
nand UO_2629 (O_2629,N_22140,N_24028);
xnor UO_2630 (O_2630,N_24195,N_24570);
and UO_2631 (O_2631,N_22169,N_22764);
or UO_2632 (O_2632,N_22349,N_24213);
and UO_2633 (O_2633,N_23283,N_23670);
or UO_2634 (O_2634,N_23792,N_24451);
nor UO_2635 (O_2635,N_22523,N_22577);
and UO_2636 (O_2636,N_22602,N_22306);
or UO_2637 (O_2637,N_22267,N_23659);
nor UO_2638 (O_2638,N_22544,N_22360);
and UO_2639 (O_2639,N_23058,N_22679);
nand UO_2640 (O_2640,N_22526,N_22927);
nor UO_2641 (O_2641,N_23637,N_22101);
or UO_2642 (O_2642,N_24603,N_23737);
and UO_2643 (O_2643,N_22143,N_24586);
nor UO_2644 (O_2644,N_24693,N_22749);
nor UO_2645 (O_2645,N_24575,N_24048);
nand UO_2646 (O_2646,N_23012,N_22461);
and UO_2647 (O_2647,N_23900,N_23616);
nand UO_2648 (O_2648,N_24097,N_22021);
nor UO_2649 (O_2649,N_22497,N_23339);
or UO_2650 (O_2650,N_23458,N_23157);
or UO_2651 (O_2651,N_24070,N_22522);
xor UO_2652 (O_2652,N_22458,N_24072);
or UO_2653 (O_2653,N_22663,N_24475);
nand UO_2654 (O_2654,N_24882,N_23061);
and UO_2655 (O_2655,N_22233,N_22415);
or UO_2656 (O_2656,N_23911,N_23816);
or UO_2657 (O_2657,N_24669,N_24577);
nand UO_2658 (O_2658,N_23019,N_22430);
and UO_2659 (O_2659,N_23334,N_22399);
or UO_2660 (O_2660,N_22675,N_22710);
xnor UO_2661 (O_2661,N_23820,N_22487);
xor UO_2662 (O_2662,N_24947,N_22496);
xnor UO_2663 (O_2663,N_24828,N_24733);
or UO_2664 (O_2664,N_22253,N_24633);
nand UO_2665 (O_2665,N_22079,N_22104);
xnor UO_2666 (O_2666,N_22452,N_23525);
or UO_2667 (O_2667,N_22285,N_22830);
nor UO_2668 (O_2668,N_22366,N_22443);
nand UO_2669 (O_2669,N_23231,N_23244);
or UO_2670 (O_2670,N_22033,N_24909);
or UO_2671 (O_2671,N_21935,N_24004);
or UO_2672 (O_2672,N_22385,N_21985);
nor UO_2673 (O_2673,N_24956,N_22161);
and UO_2674 (O_2674,N_24364,N_23451);
nand UO_2675 (O_2675,N_22897,N_23121);
or UO_2676 (O_2676,N_23447,N_22402);
or UO_2677 (O_2677,N_21981,N_22403);
or UO_2678 (O_2678,N_24793,N_22485);
or UO_2679 (O_2679,N_23016,N_23853);
and UO_2680 (O_2680,N_22285,N_22437);
nand UO_2681 (O_2681,N_22816,N_24321);
and UO_2682 (O_2682,N_22732,N_24343);
or UO_2683 (O_2683,N_24440,N_22336);
or UO_2684 (O_2684,N_21982,N_22327);
and UO_2685 (O_2685,N_23033,N_23066);
or UO_2686 (O_2686,N_23353,N_23205);
or UO_2687 (O_2687,N_23730,N_24904);
or UO_2688 (O_2688,N_24193,N_21945);
nand UO_2689 (O_2689,N_24868,N_22531);
nor UO_2690 (O_2690,N_24785,N_23051);
nor UO_2691 (O_2691,N_24541,N_24576);
and UO_2692 (O_2692,N_22996,N_24150);
xnor UO_2693 (O_2693,N_22526,N_24563);
and UO_2694 (O_2694,N_24337,N_24673);
and UO_2695 (O_2695,N_23309,N_22790);
and UO_2696 (O_2696,N_23910,N_22738);
nor UO_2697 (O_2697,N_24253,N_24016);
or UO_2698 (O_2698,N_23110,N_22436);
or UO_2699 (O_2699,N_24513,N_24746);
nand UO_2700 (O_2700,N_22669,N_22621);
nand UO_2701 (O_2701,N_22065,N_23633);
and UO_2702 (O_2702,N_22179,N_21942);
or UO_2703 (O_2703,N_23760,N_24175);
and UO_2704 (O_2704,N_24483,N_23308);
xor UO_2705 (O_2705,N_23207,N_23495);
or UO_2706 (O_2706,N_24100,N_23732);
nor UO_2707 (O_2707,N_24514,N_23493);
nor UO_2708 (O_2708,N_23815,N_24411);
and UO_2709 (O_2709,N_23922,N_24906);
and UO_2710 (O_2710,N_22279,N_22463);
and UO_2711 (O_2711,N_23468,N_23464);
or UO_2712 (O_2712,N_23375,N_24683);
nor UO_2713 (O_2713,N_23238,N_24439);
nand UO_2714 (O_2714,N_24611,N_23219);
and UO_2715 (O_2715,N_24397,N_22217);
and UO_2716 (O_2716,N_22238,N_23921);
nor UO_2717 (O_2717,N_24979,N_24920);
or UO_2718 (O_2718,N_22323,N_24849);
nor UO_2719 (O_2719,N_23955,N_22586);
nor UO_2720 (O_2720,N_22088,N_22513);
or UO_2721 (O_2721,N_23254,N_22063);
nand UO_2722 (O_2722,N_22868,N_24539);
or UO_2723 (O_2723,N_24258,N_23244);
or UO_2724 (O_2724,N_24388,N_23408);
or UO_2725 (O_2725,N_23495,N_24744);
nand UO_2726 (O_2726,N_23603,N_23009);
xor UO_2727 (O_2727,N_22068,N_23928);
nor UO_2728 (O_2728,N_23341,N_24564);
or UO_2729 (O_2729,N_22200,N_23049);
nor UO_2730 (O_2730,N_22093,N_24771);
and UO_2731 (O_2731,N_22693,N_22266);
or UO_2732 (O_2732,N_22933,N_24937);
or UO_2733 (O_2733,N_22449,N_23933);
nand UO_2734 (O_2734,N_24121,N_22327);
nand UO_2735 (O_2735,N_22885,N_24497);
and UO_2736 (O_2736,N_23003,N_24057);
and UO_2737 (O_2737,N_22204,N_22112);
xnor UO_2738 (O_2738,N_22851,N_23036);
nor UO_2739 (O_2739,N_23630,N_21954);
nand UO_2740 (O_2740,N_24557,N_23814);
or UO_2741 (O_2741,N_23332,N_24631);
or UO_2742 (O_2742,N_24739,N_22561);
nor UO_2743 (O_2743,N_22513,N_23798);
nand UO_2744 (O_2744,N_22324,N_23497);
or UO_2745 (O_2745,N_24886,N_24347);
or UO_2746 (O_2746,N_22739,N_24013);
or UO_2747 (O_2747,N_24070,N_24683);
nand UO_2748 (O_2748,N_22533,N_23694);
and UO_2749 (O_2749,N_22887,N_22821);
nor UO_2750 (O_2750,N_22266,N_22460);
and UO_2751 (O_2751,N_24351,N_22484);
nand UO_2752 (O_2752,N_24542,N_23640);
nand UO_2753 (O_2753,N_21962,N_24172);
nor UO_2754 (O_2754,N_24172,N_21977);
xnor UO_2755 (O_2755,N_22213,N_24295);
nand UO_2756 (O_2756,N_24394,N_23160);
or UO_2757 (O_2757,N_23382,N_24867);
nand UO_2758 (O_2758,N_22649,N_24444);
nand UO_2759 (O_2759,N_23243,N_22653);
and UO_2760 (O_2760,N_24033,N_22278);
and UO_2761 (O_2761,N_24877,N_23114);
and UO_2762 (O_2762,N_22776,N_23075);
and UO_2763 (O_2763,N_23692,N_24410);
nor UO_2764 (O_2764,N_24506,N_22926);
and UO_2765 (O_2765,N_22709,N_22262);
nor UO_2766 (O_2766,N_24714,N_23507);
nor UO_2767 (O_2767,N_23818,N_22811);
nand UO_2768 (O_2768,N_22835,N_23619);
and UO_2769 (O_2769,N_21966,N_24813);
or UO_2770 (O_2770,N_24901,N_24508);
nand UO_2771 (O_2771,N_22678,N_24368);
nand UO_2772 (O_2772,N_24252,N_22407);
nor UO_2773 (O_2773,N_22168,N_22532);
nand UO_2774 (O_2774,N_24754,N_23776);
nor UO_2775 (O_2775,N_23371,N_23856);
nor UO_2776 (O_2776,N_24107,N_23645);
and UO_2777 (O_2777,N_24896,N_23538);
and UO_2778 (O_2778,N_22640,N_22012);
nand UO_2779 (O_2779,N_22864,N_24637);
nor UO_2780 (O_2780,N_23108,N_24577);
nand UO_2781 (O_2781,N_22030,N_23968);
nand UO_2782 (O_2782,N_24566,N_22416);
and UO_2783 (O_2783,N_22992,N_24662);
and UO_2784 (O_2784,N_24314,N_22612);
or UO_2785 (O_2785,N_23949,N_22089);
nand UO_2786 (O_2786,N_22942,N_23821);
nor UO_2787 (O_2787,N_22251,N_23887);
xnor UO_2788 (O_2788,N_22974,N_23168);
and UO_2789 (O_2789,N_24233,N_23167);
and UO_2790 (O_2790,N_24225,N_23333);
or UO_2791 (O_2791,N_23077,N_23152);
or UO_2792 (O_2792,N_22718,N_24478);
nand UO_2793 (O_2793,N_22817,N_23826);
or UO_2794 (O_2794,N_24170,N_22186);
nand UO_2795 (O_2795,N_21943,N_22262);
or UO_2796 (O_2796,N_24650,N_22255);
nor UO_2797 (O_2797,N_24998,N_22306);
nor UO_2798 (O_2798,N_23219,N_22648);
nor UO_2799 (O_2799,N_22438,N_24418);
xnor UO_2800 (O_2800,N_22573,N_23520);
and UO_2801 (O_2801,N_22060,N_24469);
nand UO_2802 (O_2802,N_24666,N_22358);
or UO_2803 (O_2803,N_24927,N_22203);
and UO_2804 (O_2804,N_22471,N_22513);
or UO_2805 (O_2805,N_24350,N_22175);
xor UO_2806 (O_2806,N_23429,N_22369);
xor UO_2807 (O_2807,N_24179,N_24140);
nor UO_2808 (O_2808,N_24350,N_23506);
and UO_2809 (O_2809,N_22560,N_21880);
or UO_2810 (O_2810,N_23384,N_22277);
nand UO_2811 (O_2811,N_23343,N_22823);
or UO_2812 (O_2812,N_22790,N_22749);
nand UO_2813 (O_2813,N_24455,N_22566);
nand UO_2814 (O_2814,N_24139,N_23103);
or UO_2815 (O_2815,N_23118,N_22688);
and UO_2816 (O_2816,N_23843,N_23650);
and UO_2817 (O_2817,N_22932,N_23149);
nor UO_2818 (O_2818,N_21936,N_24723);
nand UO_2819 (O_2819,N_23342,N_23113);
or UO_2820 (O_2820,N_22736,N_24290);
or UO_2821 (O_2821,N_24002,N_23279);
or UO_2822 (O_2822,N_21918,N_24079);
or UO_2823 (O_2823,N_24578,N_22935);
nand UO_2824 (O_2824,N_22441,N_23690);
and UO_2825 (O_2825,N_24762,N_23910);
nand UO_2826 (O_2826,N_24731,N_23563);
nand UO_2827 (O_2827,N_23344,N_23809);
or UO_2828 (O_2828,N_23918,N_22219);
xnor UO_2829 (O_2829,N_24950,N_23859);
nor UO_2830 (O_2830,N_22477,N_22408);
nand UO_2831 (O_2831,N_22894,N_24400);
or UO_2832 (O_2832,N_24119,N_24365);
nand UO_2833 (O_2833,N_23340,N_23261);
or UO_2834 (O_2834,N_22594,N_24668);
xnor UO_2835 (O_2835,N_23206,N_22707);
or UO_2836 (O_2836,N_22972,N_21942);
nor UO_2837 (O_2837,N_23848,N_24755);
xor UO_2838 (O_2838,N_24474,N_21975);
nand UO_2839 (O_2839,N_23704,N_22800);
nor UO_2840 (O_2840,N_24222,N_24402);
nor UO_2841 (O_2841,N_22095,N_22043);
nor UO_2842 (O_2842,N_24313,N_24227);
nor UO_2843 (O_2843,N_22567,N_24789);
nor UO_2844 (O_2844,N_23953,N_23105);
and UO_2845 (O_2845,N_24804,N_22696);
and UO_2846 (O_2846,N_22924,N_21945);
nor UO_2847 (O_2847,N_22350,N_23478);
nor UO_2848 (O_2848,N_23941,N_24504);
or UO_2849 (O_2849,N_23292,N_24144);
or UO_2850 (O_2850,N_23779,N_24395);
nor UO_2851 (O_2851,N_22988,N_24958);
nand UO_2852 (O_2852,N_22596,N_22773);
xor UO_2853 (O_2853,N_23832,N_22019);
or UO_2854 (O_2854,N_22686,N_22721);
nor UO_2855 (O_2855,N_22946,N_24780);
xor UO_2856 (O_2856,N_23678,N_24074);
nor UO_2857 (O_2857,N_23806,N_23961);
nor UO_2858 (O_2858,N_24327,N_23921);
nor UO_2859 (O_2859,N_22825,N_23899);
xnor UO_2860 (O_2860,N_24398,N_23145);
nor UO_2861 (O_2861,N_22259,N_22944);
nor UO_2862 (O_2862,N_24890,N_22696);
nand UO_2863 (O_2863,N_24958,N_22037);
and UO_2864 (O_2864,N_24956,N_23376);
xor UO_2865 (O_2865,N_23101,N_24669);
nor UO_2866 (O_2866,N_22502,N_22122);
nand UO_2867 (O_2867,N_23389,N_22530);
or UO_2868 (O_2868,N_24926,N_24331);
and UO_2869 (O_2869,N_22965,N_22906);
xnor UO_2870 (O_2870,N_21928,N_24638);
nor UO_2871 (O_2871,N_24775,N_22381);
and UO_2872 (O_2872,N_22512,N_23972);
nor UO_2873 (O_2873,N_22475,N_22778);
xnor UO_2874 (O_2874,N_22602,N_23362);
xnor UO_2875 (O_2875,N_23170,N_23883);
or UO_2876 (O_2876,N_24100,N_22556);
nand UO_2877 (O_2877,N_24829,N_24342);
and UO_2878 (O_2878,N_24393,N_23692);
xnor UO_2879 (O_2879,N_23265,N_22917);
xnor UO_2880 (O_2880,N_23863,N_23952);
xor UO_2881 (O_2881,N_22881,N_22636);
nand UO_2882 (O_2882,N_23423,N_23893);
or UO_2883 (O_2883,N_23752,N_21970);
and UO_2884 (O_2884,N_23576,N_23617);
nand UO_2885 (O_2885,N_23203,N_24754);
and UO_2886 (O_2886,N_22256,N_22968);
or UO_2887 (O_2887,N_22575,N_24584);
and UO_2888 (O_2888,N_23325,N_22600);
or UO_2889 (O_2889,N_22442,N_23401);
nand UO_2890 (O_2890,N_23242,N_23290);
nand UO_2891 (O_2891,N_24947,N_22535);
or UO_2892 (O_2892,N_23965,N_22820);
nand UO_2893 (O_2893,N_22410,N_23754);
or UO_2894 (O_2894,N_23122,N_23715);
and UO_2895 (O_2895,N_23417,N_23517);
and UO_2896 (O_2896,N_24799,N_23761);
nor UO_2897 (O_2897,N_23207,N_22434);
nor UO_2898 (O_2898,N_23628,N_23694);
or UO_2899 (O_2899,N_22838,N_23564);
and UO_2900 (O_2900,N_23706,N_23876);
or UO_2901 (O_2901,N_22284,N_23460);
nand UO_2902 (O_2902,N_23565,N_24218);
nor UO_2903 (O_2903,N_23442,N_22919);
nor UO_2904 (O_2904,N_23988,N_23777);
or UO_2905 (O_2905,N_21907,N_23439);
nand UO_2906 (O_2906,N_22213,N_21940);
and UO_2907 (O_2907,N_23868,N_22179);
nor UO_2908 (O_2908,N_23225,N_22322);
nand UO_2909 (O_2909,N_22498,N_24908);
nor UO_2910 (O_2910,N_22503,N_23764);
nor UO_2911 (O_2911,N_24405,N_22389);
nand UO_2912 (O_2912,N_24801,N_23401);
or UO_2913 (O_2913,N_23247,N_22919);
nor UO_2914 (O_2914,N_22019,N_22222);
and UO_2915 (O_2915,N_24880,N_23411);
nor UO_2916 (O_2916,N_23067,N_23787);
nor UO_2917 (O_2917,N_24064,N_24528);
nor UO_2918 (O_2918,N_24771,N_21994);
nor UO_2919 (O_2919,N_23055,N_24036);
nor UO_2920 (O_2920,N_24169,N_23723);
and UO_2921 (O_2921,N_22283,N_23088);
or UO_2922 (O_2922,N_23167,N_23721);
nand UO_2923 (O_2923,N_22493,N_22190);
xnor UO_2924 (O_2924,N_22977,N_24573);
or UO_2925 (O_2925,N_24376,N_23872);
and UO_2926 (O_2926,N_24203,N_23134);
nor UO_2927 (O_2927,N_23264,N_22985);
nand UO_2928 (O_2928,N_23631,N_22364);
nor UO_2929 (O_2929,N_22853,N_24601);
nand UO_2930 (O_2930,N_24615,N_24411);
nand UO_2931 (O_2931,N_24219,N_23186);
xnor UO_2932 (O_2932,N_22518,N_23994);
nor UO_2933 (O_2933,N_23900,N_24918);
or UO_2934 (O_2934,N_22213,N_23516);
nand UO_2935 (O_2935,N_23653,N_23461);
or UO_2936 (O_2936,N_23106,N_23685);
nor UO_2937 (O_2937,N_22074,N_24935);
and UO_2938 (O_2938,N_23712,N_22872);
or UO_2939 (O_2939,N_24593,N_22049);
nor UO_2940 (O_2940,N_24891,N_23464);
nand UO_2941 (O_2941,N_23904,N_22704);
and UO_2942 (O_2942,N_24178,N_23847);
and UO_2943 (O_2943,N_24259,N_23797);
and UO_2944 (O_2944,N_22653,N_23079);
and UO_2945 (O_2945,N_24123,N_23662);
nand UO_2946 (O_2946,N_22675,N_22535);
xnor UO_2947 (O_2947,N_22542,N_22836);
or UO_2948 (O_2948,N_22867,N_22025);
nor UO_2949 (O_2949,N_22391,N_24708);
nor UO_2950 (O_2950,N_22491,N_22712);
nor UO_2951 (O_2951,N_22343,N_24017);
or UO_2952 (O_2952,N_22043,N_22071);
and UO_2953 (O_2953,N_24464,N_23128);
or UO_2954 (O_2954,N_24994,N_23653);
and UO_2955 (O_2955,N_24394,N_24511);
and UO_2956 (O_2956,N_21914,N_24415);
or UO_2957 (O_2957,N_23863,N_22541);
nand UO_2958 (O_2958,N_24659,N_23604);
nor UO_2959 (O_2959,N_22916,N_23071);
nor UO_2960 (O_2960,N_24261,N_24443);
nor UO_2961 (O_2961,N_23247,N_23580);
nand UO_2962 (O_2962,N_24779,N_24188);
and UO_2963 (O_2963,N_23028,N_22394);
or UO_2964 (O_2964,N_22328,N_22911);
or UO_2965 (O_2965,N_23164,N_23555);
nand UO_2966 (O_2966,N_24200,N_23834);
xor UO_2967 (O_2967,N_24927,N_23262);
nor UO_2968 (O_2968,N_22064,N_24041);
or UO_2969 (O_2969,N_22953,N_22919);
and UO_2970 (O_2970,N_22198,N_23051);
and UO_2971 (O_2971,N_24576,N_24360);
nor UO_2972 (O_2972,N_24133,N_22006);
nor UO_2973 (O_2973,N_22025,N_24257);
nand UO_2974 (O_2974,N_22479,N_24563);
and UO_2975 (O_2975,N_22630,N_24881);
or UO_2976 (O_2976,N_22816,N_23953);
nand UO_2977 (O_2977,N_24273,N_21902);
nor UO_2978 (O_2978,N_22697,N_24192);
xnor UO_2979 (O_2979,N_24096,N_22695);
nand UO_2980 (O_2980,N_22921,N_24229);
nand UO_2981 (O_2981,N_23282,N_22663);
nor UO_2982 (O_2982,N_22432,N_23879);
xor UO_2983 (O_2983,N_24596,N_24891);
or UO_2984 (O_2984,N_23162,N_22326);
and UO_2985 (O_2985,N_22905,N_24213);
nand UO_2986 (O_2986,N_24486,N_22310);
and UO_2987 (O_2987,N_24541,N_23642);
nor UO_2988 (O_2988,N_22029,N_24148);
nor UO_2989 (O_2989,N_24071,N_23663);
nand UO_2990 (O_2990,N_24339,N_24507);
nand UO_2991 (O_2991,N_23960,N_23016);
nor UO_2992 (O_2992,N_22842,N_24203);
nor UO_2993 (O_2993,N_23895,N_24460);
nor UO_2994 (O_2994,N_22439,N_23407);
and UO_2995 (O_2995,N_24832,N_24144);
and UO_2996 (O_2996,N_24476,N_24825);
or UO_2997 (O_2997,N_23033,N_24906);
and UO_2998 (O_2998,N_23153,N_24649);
nand UO_2999 (O_2999,N_24459,N_23423);
endmodule