module basic_500_3000_500_4_levels_1xor_2(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999;
nand U0 (N_0,In_274,In_230);
nand U1 (N_1,In_14,In_325);
and U2 (N_2,In_370,In_116);
nand U3 (N_3,In_278,In_33);
or U4 (N_4,In_125,In_267);
and U5 (N_5,In_65,In_234);
nor U6 (N_6,In_218,In_24);
or U7 (N_7,In_489,In_382);
or U8 (N_8,In_432,In_239);
or U9 (N_9,In_290,In_266);
and U10 (N_10,In_331,In_77);
nand U11 (N_11,In_244,In_42);
or U12 (N_12,In_294,In_292);
or U13 (N_13,In_420,In_51);
nor U14 (N_14,In_126,In_206);
or U15 (N_15,In_149,In_313);
nor U16 (N_16,In_473,In_401);
and U17 (N_17,In_487,In_198);
or U18 (N_18,In_312,In_207);
nor U19 (N_19,In_475,In_383);
nand U20 (N_20,In_106,In_256);
nor U21 (N_21,In_483,In_78);
nand U22 (N_22,In_273,In_480);
nand U23 (N_23,In_237,In_260);
or U24 (N_24,In_486,In_10);
nand U25 (N_25,In_213,In_227);
nor U26 (N_26,In_64,In_195);
or U27 (N_27,In_264,In_171);
nand U28 (N_28,In_317,In_62);
or U29 (N_29,In_339,In_481);
or U30 (N_30,In_414,In_61);
and U31 (N_31,In_177,In_238);
nand U32 (N_32,In_38,In_143);
nand U33 (N_33,In_87,In_377);
nand U34 (N_34,In_375,In_69);
or U35 (N_35,In_479,In_499);
nand U36 (N_36,In_393,In_21);
nor U37 (N_37,In_380,In_115);
or U38 (N_38,In_347,In_85);
and U39 (N_39,In_202,In_424);
and U40 (N_40,In_271,In_166);
and U41 (N_41,In_5,In_185);
nor U42 (N_42,In_163,In_193);
nand U43 (N_43,In_41,In_83);
and U44 (N_44,In_300,In_397);
nand U45 (N_45,In_385,In_427);
and U46 (N_46,In_31,In_450);
or U47 (N_47,In_173,In_406);
nand U48 (N_48,In_66,In_212);
nand U49 (N_49,In_330,In_444);
and U50 (N_50,In_47,In_362);
and U51 (N_51,In_351,In_469);
xnor U52 (N_52,In_29,In_392);
or U53 (N_53,In_257,In_229);
nor U54 (N_54,In_410,In_67);
and U55 (N_55,In_90,In_215);
or U56 (N_56,In_386,In_56);
or U57 (N_57,In_426,In_326);
nor U58 (N_58,In_224,In_361);
and U59 (N_59,In_18,In_68);
xor U60 (N_60,In_291,In_399);
nor U61 (N_61,In_390,In_219);
xnor U62 (N_62,In_463,In_357);
or U63 (N_63,In_153,In_54);
nor U64 (N_64,In_395,In_295);
nand U65 (N_65,In_169,In_13);
nand U66 (N_66,In_335,In_328);
and U67 (N_67,In_280,In_409);
or U68 (N_68,In_498,In_378);
nor U69 (N_69,In_263,In_270);
or U70 (N_70,In_232,In_387);
nor U71 (N_71,In_248,In_461);
and U72 (N_72,In_225,In_289);
and U73 (N_73,In_400,In_268);
nand U74 (N_74,In_293,In_184);
and U75 (N_75,In_287,In_320);
and U76 (N_76,In_452,In_358);
nand U77 (N_77,In_44,In_345);
nor U78 (N_78,In_415,In_316);
and U79 (N_79,In_297,In_497);
nor U80 (N_80,In_306,In_130);
and U81 (N_81,In_19,In_451);
and U82 (N_82,In_236,In_298);
and U83 (N_83,In_301,In_318);
nand U84 (N_84,In_190,In_307);
or U85 (N_85,In_348,In_200);
nand U86 (N_86,In_0,In_203);
nand U87 (N_87,In_168,In_91);
and U88 (N_88,In_104,In_346);
nand U89 (N_89,In_124,In_354);
nand U90 (N_90,In_102,In_440);
or U91 (N_91,In_416,In_407);
nand U92 (N_92,In_194,In_141);
xnor U93 (N_93,In_155,In_419);
nand U94 (N_94,In_223,In_144);
nor U95 (N_95,In_228,In_465);
and U96 (N_96,In_1,In_477);
and U97 (N_97,In_118,In_30);
nand U98 (N_98,In_205,In_250);
nand U99 (N_99,In_276,In_23);
and U100 (N_100,In_46,In_459);
or U101 (N_101,In_492,In_495);
and U102 (N_102,In_448,In_27);
or U103 (N_103,In_7,In_379);
and U104 (N_104,In_182,In_350);
or U105 (N_105,In_269,In_11);
nand U106 (N_106,In_366,In_389);
or U107 (N_107,In_97,In_75);
or U108 (N_108,In_468,In_132);
or U109 (N_109,In_360,In_26);
nor U110 (N_110,In_394,In_333);
and U111 (N_111,In_285,In_398);
nand U112 (N_112,In_183,In_32);
nor U113 (N_113,In_445,In_95);
nand U114 (N_114,In_288,In_137);
and U115 (N_115,In_93,In_249);
nand U116 (N_116,In_433,In_176);
or U117 (N_117,In_405,In_437);
xnor U118 (N_118,In_175,In_57);
nand U119 (N_119,In_253,In_343);
nand U120 (N_120,In_304,In_157);
nand U121 (N_121,In_337,In_167);
or U122 (N_122,In_135,In_88);
nor U123 (N_123,In_147,In_455);
nor U124 (N_124,In_36,In_16);
and U125 (N_125,In_60,In_80);
nand U126 (N_126,In_191,In_73);
nand U127 (N_127,In_281,In_423);
nor U128 (N_128,In_340,In_122);
nand U129 (N_129,In_243,In_277);
or U130 (N_130,In_111,In_404);
and U131 (N_131,In_82,In_247);
or U132 (N_132,In_45,In_128);
and U133 (N_133,In_364,In_187);
or U134 (N_134,In_96,In_282);
nand U135 (N_135,In_179,In_216);
nor U136 (N_136,In_327,In_4);
and U137 (N_137,In_208,In_431);
nor U138 (N_138,In_321,In_160);
and U139 (N_139,In_439,In_9);
nand U140 (N_140,In_210,In_48);
nor U141 (N_141,In_279,In_454);
nand U142 (N_142,In_418,In_456);
nand U143 (N_143,In_186,In_71);
and U144 (N_144,In_140,In_453);
nor U145 (N_145,In_412,In_367);
nand U146 (N_146,In_79,In_365);
nor U147 (N_147,In_22,In_472);
or U148 (N_148,In_161,In_8);
nor U149 (N_149,In_245,In_92);
nand U150 (N_150,In_484,In_403);
or U151 (N_151,In_356,In_408);
and U152 (N_152,In_478,In_52);
and U153 (N_153,In_123,In_467);
and U154 (N_154,In_188,In_302);
nand U155 (N_155,In_158,In_12);
nor U156 (N_156,In_81,In_430);
nand U157 (N_157,In_258,In_251);
nand U158 (N_158,In_127,In_252);
and U159 (N_159,In_209,In_283);
nand U160 (N_160,In_15,In_272);
nand U161 (N_161,In_152,In_222);
nand U162 (N_162,In_226,In_233);
nor U163 (N_163,In_314,In_329);
nand U164 (N_164,In_491,In_165);
or U165 (N_165,In_142,In_164);
nand U166 (N_166,In_436,In_310);
nor U167 (N_167,In_121,In_180);
xor U168 (N_168,In_107,In_113);
and U169 (N_169,In_324,In_221);
nor U170 (N_170,In_2,In_131);
and U171 (N_171,In_355,In_34);
and U172 (N_172,In_336,In_63);
nor U173 (N_173,In_50,In_76);
nor U174 (N_174,In_352,In_6);
nor U175 (N_175,In_349,In_58);
nor U176 (N_176,In_110,In_134);
or U177 (N_177,In_199,In_402);
and U178 (N_178,In_374,In_438);
or U179 (N_179,In_211,In_55);
nor U180 (N_180,In_334,In_315);
nand U181 (N_181,In_396,In_25);
and U182 (N_182,In_372,In_363);
nand U183 (N_183,In_369,In_39);
nor U184 (N_184,In_43,In_98);
nor U185 (N_185,In_490,In_296);
xor U186 (N_186,In_470,In_485);
or U187 (N_187,In_368,In_474);
nand U188 (N_188,In_482,In_162);
xor U189 (N_189,In_94,In_240);
xnor U190 (N_190,In_447,In_53);
or U191 (N_191,In_99,In_20);
or U192 (N_192,In_133,In_119);
nand U193 (N_193,In_422,In_105);
or U194 (N_194,In_265,In_100);
nand U195 (N_195,In_460,In_108);
and U196 (N_196,In_413,In_181);
nand U197 (N_197,In_442,In_196);
nor U198 (N_198,In_72,In_464);
nand U199 (N_199,In_139,In_308);
nor U200 (N_200,In_84,In_197);
nand U201 (N_201,In_217,In_172);
and U202 (N_202,In_204,In_476);
and U203 (N_203,In_255,In_471);
or U204 (N_204,In_388,In_103);
nor U205 (N_205,In_458,In_154);
and U206 (N_206,In_286,In_443);
or U207 (N_207,In_284,In_373);
nand U208 (N_208,In_242,In_466);
or U209 (N_209,In_112,In_359);
nand U210 (N_210,In_3,In_303);
and U211 (N_211,In_381,In_417);
and U212 (N_212,In_156,In_159);
and U213 (N_213,In_214,In_254);
nand U214 (N_214,In_129,In_40);
or U215 (N_215,In_189,In_435);
nor U216 (N_216,In_441,In_170);
nor U217 (N_217,In_28,In_494);
and U218 (N_218,In_151,In_89);
and U219 (N_219,In_262,In_428);
nor U220 (N_220,In_311,In_421);
or U221 (N_221,In_86,In_371);
nor U222 (N_222,In_138,In_299);
nor U223 (N_223,In_114,In_220);
nand U224 (N_224,In_344,In_101);
and U225 (N_225,In_446,In_35);
or U226 (N_226,In_148,In_319);
and U227 (N_227,In_353,In_178);
and U228 (N_228,In_59,In_434);
or U229 (N_229,In_109,In_462);
nor U230 (N_230,In_338,In_174);
and U231 (N_231,In_411,In_17);
and U232 (N_232,In_235,In_246);
and U233 (N_233,In_49,In_74);
or U234 (N_234,In_231,In_488);
and U235 (N_235,In_201,In_376);
nor U236 (N_236,In_117,In_332);
nand U237 (N_237,In_136,In_457);
nand U238 (N_238,In_309,In_259);
or U239 (N_239,In_342,In_391);
nand U240 (N_240,In_150,In_145);
or U241 (N_241,In_275,In_192);
nand U242 (N_242,In_341,In_496);
or U243 (N_243,In_146,In_429);
or U244 (N_244,In_322,In_261);
nor U245 (N_245,In_37,In_241);
nand U246 (N_246,In_449,In_493);
nand U247 (N_247,In_305,In_425);
nor U248 (N_248,In_384,In_70);
nand U249 (N_249,In_323,In_120);
and U250 (N_250,In_333,In_119);
and U251 (N_251,In_79,In_398);
or U252 (N_252,In_305,In_310);
and U253 (N_253,In_414,In_355);
or U254 (N_254,In_230,In_99);
and U255 (N_255,In_454,In_327);
nor U256 (N_256,In_192,In_177);
and U257 (N_257,In_188,In_388);
nand U258 (N_258,In_299,In_179);
or U259 (N_259,In_92,In_256);
or U260 (N_260,In_78,In_169);
or U261 (N_261,In_374,In_268);
or U262 (N_262,In_322,In_101);
nand U263 (N_263,In_232,In_460);
or U264 (N_264,In_227,In_141);
or U265 (N_265,In_261,In_33);
nand U266 (N_266,In_293,In_449);
nor U267 (N_267,In_423,In_465);
or U268 (N_268,In_258,In_91);
or U269 (N_269,In_89,In_184);
nand U270 (N_270,In_340,In_372);
nor U271 (N_271,In_295,In_309);
nand U272 (N_272,In_167,In_17);
nand U273 (N_273,In_15,In_236);
nand U274 (N_274,In_499,In_4);
or U275 (N_275,In_192,In_357);
nand U276 (N_276,In_322,In_367);
or U277 (N_277,In_189,In_283);
nor U278 (N_278,In_334,In_372);
and U279 (N_279,In_154,In_276);
nor U280 (N_280,In_343,In_65);
or U281 (N_281,In_462,In_160);
nand U282 (N_282,In_46,In_208);
nor U283 (N_283,In_411,In_26);
nand U284 (N_284,In_147,In_406);
and U285 (N_285,In_446,In_319);
or U286 (N_286,In_375,In_72);
and U287 (N_287,In_291,In_402);
or U288 (N_288,In_358,In_289);
nand U289 (N_289,In_435,In_482);
and U290 (N_290,In_168,In_417);
nand U291 (N_291,In_426,In_198);
nand U292 (N_292,In_41,In_406);
nand U293 (N_293,In_472,In_346);
nand U294 (N_294,In_370,In_49);
and U295 (N_295,In_283,In_118);
nor U296 (N_296,In_67,In_334);
and U297 (N_297,In_422,In_364);
and U298 (N_298,In_48,In_340);
xnor U299 (N_299,In_265,In_113);
and U300 (N_300,In_384,In_343);
nand U301 (N_301,In_258,In_359);
or U302 (N_302,In_372,In_384);
and U303 (N_303,In_162,In_328);
nor U304 (N_304,In_418,In_278);
nand U305 (N_305,In_302,In_323);
nand U306 (N_306,In_226,In_445);
nand U307 (N_307,In_167,In_400);
nor U308 (N_308,In_93,In_173);
or U309 (N_309,In_119,In_288);
nand U310 (N_310,In_471,In_366);
nand U311 (N_311,In_92,In_205);
or U312 (N_312,In_264,In_350);
or U313 (N_313,In_351,In_451);
and U314 (N_314,In_152,In_325);
and U315 (N_315,In_452,In_262);
or U316 (N_316,In_33,In_290);
nor U317 (N_317,In_446,In_396);
or U318 (N_318,In_493,In_91);
or U319 (N_319,In_167,In_276);
nand U320 (N_320,In_206,In_163);
and U321 (N_321,In_98,In_185);
nand U322 (N_322,In_89,In_133);
and U323 (N_323,In_359,In_331);
or U324 (N_324,In_422,In_44);
or U325 (N_325,In_240,In_290);
or U326 (N_326,In_11,In_170);
nand U327 (N_327,In_314,In_105);
or U328 (N_328,In_57,In_413);
nand U329 (N_329,In_312,In_418);
and U330 (N_330,In_389,In_287);
nand U331 (N_331,In_23,In_145);
nand U332 (N_332,In_387,In_425);
or U333 (N_333,In_277,In_233);
nand U334 (N_334,In_152,In_193);
nor U335 (N_335,In_403,In_61);
and U336 (N_336,In_51,In_261);
nand U337 (N_337,In_237,In_122);
and U338 (N_338,In_379,In_68);
nor U339 (N_339,In_353,In_219);
nand U340 (N_340,In_312,In_274);
nor U341 (N_341,In_3,In_4);
or U342 (N_342,In_352,In_371);
nand U343 (N_343,In_346,In_355);
and U344 (N_344,In_188,In_288);
nand U345 (N_345,In_489,In_200);
or U346 (N_346,In_253,In_387);
and U347 (N_347,In_150,In_43);
and U348 (N_348,In_165,In_264);
nand U349 (N_349,In_129,In_264);
nand U350 (N_350,In_323,In_150);
nand U351 (N_351,In_349,In_31);
nand U352 (N_352,In_423,In_431);
or U353 (N_353,In_175,In_70);
and U354 (N_354,In_157,In_226);
or U355 (N_355,In_309,In_445);
nor U356 (N_356,In_140,In_291);
nor U357 (N_357,In_164,In_331);
nand U358 (N_358,In_48,In_138);
xor U359 (N_359,In_470,In_97);
nor U360 (N_360,In_425,In_148);
nand U361 (N_361,In_312,In_485);
nor U362 (N_362,In_406,In_140);
or U363 (N_363,In_86,In_53);
or U364 (N_364,In_466,In_334);
or U365 (N_365,In_447,In_129);
nor U366 (N_366,In_302,In_392);
and U367 (N_367,In_165,In_445);
or U368 (N_368,In_291,In_416);
or U369 (N_369,In_334,In_236);
or U370 (N_370,In_181,In_387);
nand U371 (N_371,In_5,In_220);
nand U372 (N_372,In_99,In_411);
or U373 (N_373,In_292,In_377);
nand U374 (N_374,In_133,In_165);
nand U375 (N_375,In_18,In_117);
and U376 (N_376,In_325,In_441);
nor U377 (N_377,In_488,In_306);
nor U378 (N_378,In_373,In_279);
or U379 (N_379,In_331,In_27);
nor U380 (N_380,In_451,In_53);
and U381 (N_381,In_248,In_51);
nor U382 (N_382,In_440,In_324);
nand U383 (N_383,In_489,In_146);
or U384 (N_384,In_490,In_25);
nor U385 (N_385,In_225,In_367);
or U386 (N_386,In_123,In_111);
nand U387 (N_387,In_149,In_245);
nor U388 (N_388,In_238,In_112);
nand U389 (N_389,In_418,In_371);
and U390 (N_390,In_39,In_338);
or U391 (N_391,In_346,In_179);
nand U392 (N_392,In_263,In_242);
nor U393 (N_393,In_355,In_84);
nand U394 (N_394,In_289,In_6);
or U395 (N_395,In_408,In_250);
xnor U396 (N_396,In_80,In_236);
nor U397 (N_397,In_162,In_216);
and U398 (N_398,In_299,In_259);
or U399 (N_399,In_90,In_345);
nand U400 (N_400,In_166,In_66);
or U401 (N_401,In_0,In_76);
nand U402 (N_402,In_196,In_42);
nand U403 (N_403,In_11,In_431);
and U404 (N_404,In_291,In_64);
and U405 (N_405,In_437,In_479);
or U406 (N_406,In_38,In_474);
or U407 (N_407,In_210,In_385);
or U408 (N_408,In_386,In_347);
nand U409 (N_409,In_204,In_188);
or U410 (N_410,In_89,In_353);
or U411 (N_411,In_384,In_95);
and U412 (N_412,In_335,In_480);
or U413 (N_413,In_326,In_477);
nand U414 (N_414,In_29,In_108);
or U415 (N_415,In_333,In_237);
nor U416 (N_416,In_498,In_319);
nand U417 (N_417,In_222,In_138);
or U418 (N_418,In_471,In_12);
and U419 (N_419,In_388,In_44);
nand U420 (N_420,In_10,In_216);
and U421 (N_421,In_333,In_147);
nor U422 (N_422,In_11,In_436);
nor U423 (N_423,In_229,In_58);
nand U424 (N_424,In_198,In_367);
xor U425 (N_425,In_113,In_53);
nand U426 (N_426,In_70,In_254);
or U427 (N_427,In_276,In_30);
nor U428 (N_428,In_63,In_66);
or U429 (N_429,In_196,In_10);
and U430 (N_430,In_458,In_212);
nand U431 (N_431,In_396,In_487);
nand U432 (N_432,In_161,In_495);
or U433 (N_433,In_68,In_55);
or U434 (N_434,In_316,In_388);
and U435 (N_435,In_157,In_144);
and U436 (N_436,In_243,In_477);
or U437 (N_437,In_387,In_179);
nor U438 (N_438,In_382,In_66);
nor U439 (N_439,In_23,In_464);
and U440 (N_440,In_375,In_251);
nor U441 (N_441,In_318,In_447);
nand U442 (N_442,In_210,In_259);
nor U443 (N_443,In_316,In_378);
and U444 (N_444,In_452,In_88);
and U445 (N_445,In_339,In_375);
or U446 (N_446,In_87,In_239);
and U447 (N_447,In_31,In_189);
and U448 (N_448,In_92,In_110);
nor U449 (N_449,In_432,In_253);
and U450 (N_450,In_433,In_211);
or U451 (N_451,In_70,In_338);
or U452 (N_452,In_365,In_215);
nand U453 (N_453,In_473,In_368);
or U454 (N_454,In_306,In_292);
and U455 (N_455,In_351,In_163);
and U456 (N_456,In_158,In_488);
nor U457 (N_457,In_366,In_131);
nand U458 (N_458,In_257,In_344);
nor U459 (N_459,In_367,In_374);
nor U460 (N_460,In_389,In_244);
nand U461 (N_461,In_170,In_301);
nand U462 (N_462,In_123,In_378);
nor U463 (N_463,In_199,In_76);
nand U464 (N_464,In_171,In_263);
nand U465 (N_465,In_498,In_120);
and U466 (N_466,In_203,In_401);
nand U467 (N_467,In_262,In_276);
nor U468 (N_468,In_265,In_14);
or U469 (N_469,In_149,In_466);
nor U470 (N_470,In_450,In_24);
nand U471 (N_471,In_355,In_68);
nand U472 (N_472,In_213,In_494);
or U473 (N_473,In_362,In_273);
and U474 (N_474,In_125,In_310);
or U475 (N_475,In_20,In_19);
nand U476 (N_476,In_438,In_440);
nand U477 (N_477,In_401,In_348);
or U478 (N_478,In_467,In_483);
and U479 (N_479,In_141,In_290);
and U480 (N_480,In_371,In_98);
or U481 (N_481,In_56,In_488);
or U482 (N_482,In_445,In_391);
nand U483 (N_483,In_208,In_118);
nor U484 (N_484,In_340,In_211);
nand U485 (N_485,In_457,In_12);
and U486 (N_486,In_326,In_384);
nand U487 (N_487,In_496,In_206);
and U488 (N_488,In_324,In_91);
xor U489 (N_489,In_385,In_383);
nand U490 (N_490,In_452,In_379);
or U491 (N_491,In_236,In_416);
nand U492 (N_492,In_45,In_366);
nand U493 (N_493,In_407,In_441);
or U494 (N_494,In_223,In_176);
nand U495 (N_495,In_12,In_436);
nand U496 (N_496,In_305,In_477);
and U497 (N_497,In_445,In_146);
nor U498 (N_498,In_175,In_337);
and U499 (N_499,In_371,In_329);
or U500 (N_500,In_109,In_54);
nor U501 (N_501,In_131,In_178);
nor U502 (N_502,In_185,In_131);
and U503 (N_503,In_291,In_80);
or U504 (N_504,In_76,In_119);
and U505 (N_505,In_419,In_400);
or U506 (N_506,In_472,In_45);
nor U507 (N_507,In_14,In_106);
nand U508 (N_508,In_314,In_51);
nor U509 (N_509,In_216,In_369);
nand U510 (N_510,In_138,In_325);
or U511 (N_511,In_398,In_225);
nand U512 (N_512,In_17,In_177);
and U513 (N_513,In_201,In_191);
or U514 (N_514,In_485,In_413);
or U515 (N_515,In_164,In_353);
or U516 (N_516,In_315,In_415);
nand U517 (N_517,In_63,In_445);
or U518 (N_518,In_477,In_158);
or U519 (N_519,In_173,In_255);
and U520 (N_520,In_136,In_271);
and U521 (N_521,In_45,In_12);
or U522 (N_522,In_234,In_150);
or U523 (N_523,In_140,In_431);
nand U524 (N_524,In_368,In_271);
nor U525 (N_525,In_51,In_212);
or U526 (N_526,In_425,In_191);
or U527 (N_527,In_285,In_94);
or U528 (N_528,In_171,In_63);
and U529 (N_529,In_225,In_192);
nor U530 (N_530,In_120,In_360);
nand U531 (N_531,In_111,In_104);
or U532 (N_532,In_416,In_57);
nand U533 (N_533,In_40,In_210);
and U534 (N_534,In_254,In_170);
or U535 (N_535,In_234,In_487);
nor U536 (N_536,In_75,In_203);
or U537 (N_537,In_438,In_28);
nand U538 (N_538,In_405,In_283);
xnor U539 (N_539,In_119,In_385);
and U540 (N_540,In_112,In_102);
nand U541 (N_541,In_420,In_379);
nand U542 (N_542,In_381,In_326);
or U543 (N_543,In_105,In_351);
nor U544 (N_544,In_329,In_30);
or U545 (N_545,In_136,In_261);
or U546 (N_546,In_145,In_387);
and U547 (N_547,In_478,In_20);
or U548 (N_548,In_236,In_468);
xor U549 (N_549,In_113,In_455);
or U550 (N_550,In_310,In_66);
nand U551 (N_551,In_199,In_498);
nor U552 (N_552,In_385,In_305);
nand U553 (N_553,In_19,In_136);
xor U554 (N_554,In_280,In_254);
or U555 (N_555,In_222,In_134);
nand U556 (N_556,In_136,In_92);
or U557 (N_557,In_82,In_332);
nand U558 (N_558,In_478,In_196);
or U559 (N_559,In_488,In_31);
and U560 (N_560,In_263,In_41);
or U561 (N_561,In_361,In_152);
and U562 (N_562,In_156,In_261);
nand U563 (N_563,In_143,In_352);
or U564 (N_564,In_401,In_256);
or U565 (N_565,In_40,In_430);
nor U566 (N_566,In_416,In_183);
nor U567 (N_567,In_20,In_346);
nand U568 (N_568,In_306,In_309);
or U569 (N_569,In_196,In_394);
or U570 (N_570,In_288,In_481);
nand U571 (N_571,In_369,In_245);
or U572 (N_572,In_262,In_336);
and U573 (N_573,In_5,In_281);
or U574 (N_574,In_384,In_422);
nand U575 (N_575,In_207,In_227);
and U576 (N_576,In_213,In_486);
nand U577 (N_577,In_300,In_100);
nand U578 (N_578,In_328,In_280);
nor U579 (N_579,In_268,In_357);
or U580 (N_580,In_32,In_112);
and U581 (N_581,In_77,In_427);
nor U582 (N_582,In_42,In_496);
nor U583 (N_583,In_289,In_88);
nor U584 (N_584,In_130,In_362);
or U585 (N_585,In_389,In_310);
nand U586 (N_586,In_234,In_140);
and U587 (N_587,In_98,In_126);
nor U588 (N_588,In_390,In_345);
nand U589 (N_589,In_372,In_465);
or U590 (N_590,In_383,In_185);
and U591 (N_591,In_9,In_163);
or U592 (N_592,In_195,In_250);
or U593 (N_593,In_131,In_475);
nand U594 (N_594,In_69,In_354);
and U595 (N_595,In_50,In_441);
or U596 (N_596,In_417,In_109);
nand U597 (N_597,In_378,In_223);
nand U598 (N_598,In_212,In_15);
nand U599 (N_599,In_206,In_489);
or U600 (N_600,In_429,In_366);
nor U601 (N_601,In_322,In_410);
and U602 (N_602,In_72,In_441);
nor U603 (N_603,In_239,In_461);
or U604 (N_604,In_44,In_275);
and U605 (N_605,In_264,In_489);
or U606 (N_606,In_456,In_311);
nand U607 (N_607,In_401,In_206);
and U608 (N_608,In_127,In_466);
nor U609 (N_609,In_91,In_459);
nand U610 (N_610,In_190,In_446);
nand U611 (N_611,In_308,In_59);
or U612 (N_612,In_27,In_467);
nand U613 (N_613,In_358,In_260);
nand U614 (N_614,In_176,In_49);
or U615 (N_615,In_330,In_53);
nor U616 (N_616,In_422,In_21);
xnor U617 (N_617,In_441,In_472);
nand U618 (N_618,In_153,In_240);
and U619 (N_619,In_393,In_435);
or U620 (N_620,In_185,In_438);
nor U621 (N_621,In_478,In_429);
and U622 (N_622,In_166,In_377);
or U623 (N_623,In_375,In_427);
nand U624 (N_624,In_400,In_450);
xor U625 (N_625,In_398,In_90);
nor U626 (N_626,In_383,In_464);
and U627 (N_627,In_157,In_215);
nand U628 (N_628,In_101,In_217);
and U629 (N_629,In_190,In_30);
and U630 (N_630,In_312,In_273);
nor U631 (N_631,In_206,In_498);
or U632 (N_632,In_431,In_3);
or U633 (N_633,In_288,In_363);
or U634 (N_634,In_36,In_226);
or U635 (N_635,In_43,In_418);
or U636 (N_636,In_372,In_245);
nand U637 (N_637,In_158,In_323);
nand U638 (N_638,In_149,In_88);
and U639 (N_639,In_440,In_264);
and U640 (N_640,In_145,In_280);
nor U641 (N_641,In_282,In_350);
nor U642 (N_642,In_127,In_8);
xnor U643 (N_643,In_233,In_69);
nand U644 (N_644,In_246,In_143);
or U645 (N_645,In_105,In_333);
xor U646 (N_646,In_101,In_90);
and U647 (N_647,In_347,In_72);
nor U648 (N_648,In_287,In_309);
or U649 (N_649,In_328,In_389);
xor U650 (N_650,In_336,In_38);
nor U651 (N_651,In_128,In_9);
nor U652 (N_652,In_126,In_186);
and U653 (N_653,In_274,In_352);
nor U654 (N_654,In_194,In_14);
or U655 (N_655,In_1,In_224);
and U656 (N_656,In_335,In_302);
nor U657 (N_657,In_204,In_113);
or U658 (N_658,In_300,In_439);
or U659 (N_659,In_36,In_47);
or U660 (N_660,In_361,In_128);
nor U661 (N_661,In_206,In_298);
nand U662 (N_662,In_217,In_204);
and U663 (N_663,In_451,In_437);
and U664 (N_664,In_384,In_169);
nand U665 (N_665,In_127,In_297);
nor U666 (N_666,In_81,In_255);
or U667 (N_667,In_7,In_34);
or U668 (N_668,In_59,In_498);
and U669 (N_669,In_349,In_481);
and U670 (N_670,In_21,In_454);
and U671 (N_671,In_8,In_51);
nand U672 (N_672,In_40,In_35);
or U673 (N_673,In_263,In_220);
nor U674 (N_674,In_2,In_442);
nand U675 (N_675,In_394,In_324);
and U676 (N_676,In_339,In_116);
nand U677 (N_677,In_202,In_412);
nand U678 (N_678,In_115,In_281);
nor U679 (N_679,In_477,In_119);
and U680 (N_680,In_92,In_453);
or U681 (N_681,In_1,In_470);
and U682 (N_682,In_94,In_486);
or U683 (N_683,In_322,In_27);
nor U684 (N_684,In_313,In_174);
nand U685 (N_685,In_167,In_223);
nand U686 (N_686,In_404,In_92);
nor U687 (N_687,In_363,In_216);
or U688 (N_688,In_269,In_419);
nor U689 (N_689,In_403,In_17);
or U690 (N_690,In_343,In_439);
or U691 (N_691,In_257,In_340);
nor U692 (N_692,In_115,In_311);
nand U693 (N_693,In_89,In_401);
or U694 (N_694,In_179,In_91);
nor U695 (N_695,In_153,In_466);
and U696 (N_696,In_253,In_456);
nor U697 (N_697,In_238,In_331);
or U698 (N_698,In_100,In_499);
and U699 (N_699,In_320,In_422);
and U700 (N_700,In_107,In_241);
and U701 (N_701,In_371,In_242);
nand U702 (N_702,In_488,In_18);
nor U703 (N_703,In_457,In_431);
or U704 (N_704,In_196,In_491);
nand U705 (N_705,In_149,In_216);
or U706 (N_706,In_420,In_125);
nand U707 (N_707,In_356,In_463);
or U708 (N_708,In_118,In_133);
or U709 (N_709,In_129,In_360);
nor U710 (N_710,In_1,In_261);
or U711 (N_711,In_310,In_401);
or U712 (N_712,In_57,In_314);
or U713 (N_713,In_256,In_0);
or U714 (N_714,In_237,In_270);
and U715 (N_715,In_79,In_158);
or U716 (N_716,In_322,In_460);
and U717 (N_717,In_413,In_334);
nand U718 (N_718,In_298,In_380);
nor U719 (N_719,In_276,In_141);
nand U720 (N_720,In_304,In_349);
xnor U721 (N_721,In_237,In_410);
nand U722 (N_722,In_384,In_99);
nand U723 (N_723,In_241,In_400);
and U724 (N_724,In_18,In_442);
or U725 (N_725,In_453,In_169);
and U726 (N_726,In_312,In_279);
nor U727 (N_727,In_493,In_485);
nand U728 (N_728,In_10,In_342);
or U729 (N_729,In_321,In_483);
nor U730 (N_730,In_18,In_309);
or U731 (N_731,In_155,In_270);
nor U732 (N_732,In_454,In_282);
nor U733 (N_733,In_5,In_236);
and U734 (N_734,In_417,In_324);
nor U735 (N_735,In_250,In_295);
or U736 (N_736,In_214,In_303);
nand U737 (N_737,In_225,In_170);
nor U738 (N_738,In_271,In_219);
nand U739 (N_739,In_101,In_108);
nor U740 (N_740,In_51,In_288);
and U741 (N_741,In_341,In_79);
nor U742 (N_742,In_36,In_192);
or U743 (N_743,In_351,In_78);
or U744 (N_744,In_395,In_328);
nor U745 (N_745,In_178,In_488);
nand U746 (N_746,In_210,In_475);
nand U747 (N_747,In_477,In_202);
xnor U748 (N_748,In_203,In_486);
or U749 (N_749,In_422,In_230);
nor U750 (N_750,N_13,N_313);
nor U751 (N_751,N_715,N_252);
nor U752 (N_752,N_301,N_343);
and U753 (N_753,N_534,N_472);
nand U754 (N_754,N_373,N_102);
and U755 (N_755,N_505,N_174);
nor U756 (N_756,N_443,N_464);
and U757 (N_757,N_440,N_219);
nor U758 (N_758,N_749,N_577);
or U759 (N_759,N_541,N_173);
nand U760 (N_760,N_168,N_478);
nand U761 (N_761,N_142,N_309);
nand U762 (N_762,N_385,N_531);
and U763 (N_763,N_466,N_50);
nand U764 (N_764,N_570,N_631);
and U765 (N_765,N_590,N_650);
or U766 (N_766,N_361,N_295);
nand U767 (N_767,N_399,N_459);
nor U768 (N_768,N_308,N_639);
or U769 (N_769,N_109,N_282);
and U770 (N_770,N_341,N_100);
or U771 (N_771,N_38,N_406);
and U772 (N_772,N_351,N_193);
nor U773 (N_773,N_20,N_1);
and U774 (N_774,N_186,N_331);
and U775 (N_775,N_365,N_288);
and U776 (N_776,N_729,N_407);
nand U777 (N_777,N_22,N_571);
or U778 (N_778,N_118,N_511);
and U779 (N_779,N_708,N_504);
nand U780 (N_780,N_84,N_356);
nand U781 (N_781,N_528,N_388);
nand U782 (N_782,N_600,N_368);
nor U783 (N_783,N_414,N_322);
nor U784 (N_784,N_603,N_371);
and U785 (N_785,N_349,N_702);
nand U786 (N_786,N_294,N_265);
or U787 (N_787,N_196,N_101);
or U788 (N_788,N_576,N_587);
nor U789 (N_789,N_649,N_474);
nor U790 (N_790,N_648,N_699);
and U791 (N_791,N_81,N_350);
or U792 (N_792,N_524,N_564);
nor U793 (N_793,N_311,N_192);
or U794 (N_794,N_659,N_215);
and U795 (N_795,N_501,N_745);
nand U796 (N_796,N_691,N_610);
nand U797 (N_797,N_253,N_289);
and U798 (N_798,N_409,N_739);
nor U799 (N_799,N_494,N_55);
and U800 (N_800,N_134,N_404);
nor U801 (N_801,N_139,N_278);
nand U802 (N_802,N_463,N_697);
nand U803 (N_803,N_632,N_557);
nor U804 (N_804,N_329,N_232);
nor U805 (N_805,N_608,N_519);
nor U806 (N_806,N_347,N_605);
nand U807 (N_807,N_65,N_653);
nor U808 (N_808,N_444,N_680);
and U809 (N_809,N_185,N_255);
or U810 (N_810,N_310,N_179);
nor U811 (N_811,N_116,N_562);
nor U812 (N_812,N_107,N_147);
nor U813 (N_813,N_269,N_470);
and U814 (N_814,N_279,N_86);
and U815 (N_815,N_489,N_162);
nor U816 (N_816,N_197,N_513);
nand U817 (N_817,N_446,N_18);
or U818 (N_818,N_130,N_630);
nor U819 (N_819,N_296,N_140);
nor U820 (N_820,N_517,N_31);
nand U821 (N_821,N_302,N_54);
nand U822 (N_822,N_285,N_19);
and U823 (N_823,N_423,N_437);
nor U824 (N_824,N_203,N_607);
and U825 (N_825,N_551,N_67);
nor U826 (N_826,N_496,N_63);
nor U827 (N_827,N_121,N_432);
nand U828 (N_828,N_195,N_272);
nand U829 (N_829,N_676,N_231);
nand U830 (N_830,N_293,N_125);
or U831 (N_831,N_149,N_9);
nor U832 (N_832,N_224,N_448);
and U833 (N_833,N_667,N_359);
or U834 (N_834,N_122,N_317);
and U835 (N_835,N_159,N_613);
and U836 (N_836,N_730,N_623);
and U837 (N_837,N_334,N_549);
and U838 (N_838,N_438,N_495);
nand U839 (N_839,N_312,N_469);
nand U840 (N_840,N_320,N_479);
and U841 (N_841,N_737,N_628);
nor U842 (N_842,N_290,N_403);
and U843 (N_843,N_286,N_204);
or U844 (N_844,N_565,N_327);
or U845 (N_845,N_182,N_257);
or U846 (N_846,N_580,N_383);
and U847 (N_847,N_304,N_636);
nor U848 (N_848,N_180,N_2);
and U849 (N_849,N_53,N_574);
nand U850 (N_850,N_270,N_337);
or U851 (N_851,N_572,N_324);
nor U852 (N_852,N_129,N_170);
nand U853 (N_853,N_358,N_71);
or U854 (N_854,N_94,N_635);
or U855 (N_855,N_546,N_143);
nand U856 (N_856,N_679,N_740);
and U857 (N_857,N_412,N_240);
and U858 (N_858,N_451,N_410);
and U859 (N_859,N_105,N_675);
nand U860 (N_860,N_484,N_201);
or U861 (N_861,N_238,N_573);
nor U862 (N_862,N_742,N_644);
nand U863 (N_863,N_428,N_281);
nor U864 (N_864,N_357,N_160);
nor U865 (N_865,N_5,N_633);
and U866 (N_866,N_473,N_372);
and U867 (N_867,N_326,N_264);
nor U868 (N_868,N_123,N_236);
and U869 (N_869,N_533,N_391);
nand U870 (N_870,N_626,N_567);
and U871 (N_871,N_651,N_468);
and U872 (N_872,N_457,N_223);
or U873 (N_873,N_42,N_529);
or U874 (N_874,N_181,N_548);
nand U875 (N_875,N_332,N_543);
or U876 (N_876,N_674,N_604);
or U877 (N_877,N_425,N_330);
nand U878 (N_878,N_28,N_376);
or U879 (N_879,N_141,N_589);
and U880 (N_880,N_268,N_554);
nand U881 (N_881,N_601,N_111);
nor U882 (N_882,N_10,N_427);
and U883 (N_883,N_569,N_660);
nor U884 (N_884,N_396,N_58);
or U885 (N_885,N_559,N_335);
nor U886 (N_886,N_138,N_178);
nor U887 (N_887,N_612,N_115);
or U888 (N_888,N_200,N_266);
nor U889 (N_889,N_669,N_536);
nand U890 (N_890,N_202,N_538);
xor U891 (N_891,N_362,N_619);
and U892 (N_892,N_621,N_614);
and U893 (N_893,N_490,N_720);
nand U894 (N_894,N_685,N_70);
and U895 (N_895,N_360,N_422);
nand U896 (N_896,N_599,N_507);
nand U897 (N_897,N_678,N_526);
nand U898 (N_898,N_62,N_33);
or U899 (N_899,N_237,N_460);
nand U900 (N_900,N_104,N_378);
nand U901 (N_901,N_690,N_61);
nor U902 (N_902,N_500,N_712);
or U903 (N_903,N_39,N_634);
nor U904 (N_904,N_401,N_161);
nand U905 (N_905,N_655,N_390);
nor U906 (N_906,N_207,N_420);
xor U907 (N_907,N_728,N_214);
nor U908 (N_908,N_277,N_59);
or U909 (N_909,N_283,N_540);
or U910 (N_910,N_512,N_6);
nor U911 (N_911,N_527,N_492);
nand U912 (N_912,N_263,N_208);
nor U913 (N_913,N_688,N_213);
nand U914 (N_914,N_108,N_389);
and U915 (N_915,N_498,N_306);
nor U916 (N_916,N_627,N_319);
and U917 (N_917,N_439,N_611);
or U918 (N_918,N_411,N_618);
and U919 (N_919,N_561,N_346);
or U920 (N_920,N_449,N_128);
and U921 (N_921,N_689,N_416);
or U922 (N_922,N_27,N_355);
nor U923 (N_923,N_719,N_471);
nand U924 (N_924,N_731,N_344);
nand U925 (N_925,N_661,N_191);
nor U926 (N_926,N_336,N_397);
or U927 (N_927,N_638,N_458);
nand U928 (N_928,N_687,N_476);
nor U929 (N_929,N_502,N_522);
or U930 (N_930,N_683,N_694);
or U931 (N_931,N_624,N_64);
nor U932 (N_932,N_593,N_707);
xnor U933 (N_933,N_657,N_692);
nor U934 (N_934,N_35,N_227);
and U935 (N_935,N_384,N_247);
and U936 (N_936,N_426,N_76);
and U937 (N_937,N_26,N_436);
nand U938 (N_938,N_199,N_66);
nor U939 (N_939,N_413,N_441);
nor U940 (N_940,N_508,N_226);
nand U941 (N_941,N_155,N_321);
nand U942 (N_942,N_56,N_733);
nor U943 (N_943,N_176,N_251);
and U944 (N_944,N_563,N_617);
nor U945 (N_945,N_582,N_465);
nor U946 (N_946,N_291,N_609);
nand U947 (N_947,N_225,N_475);
nor U948 (N_948,N_395,N_732);
and U949 (N_949,N_189,N_110);
nand U950 (N_950,N_12,N_339);
or U951 (N_951,N_695,N_175);
or U952 (N_952,N_656,N_21);
xnor U953 (N_953,N_73,N_14);
and U954 (N_954,N_398,N_566);
nand U955 (N_955,N_434,N_724);
nor U956 (N_956,N_284,N_684);
nand U957 (N_957,N_620,N_113);
and U958 (N_958,N_408,N_568);
nand U959 (N_959,N_698,N_598);
and U960 (N_960,N_664,N_442);
nor U961 (N_961,N_514,N_169);
nor U962 (N_962,N_43,N_177);
nand U963 (N_963,N_467,N_297);
nor U964 (N_964,N_154,N_153);
nand U965 (N_965,N_616,N_435);
or U966 (N_966,N_69,N_455);
and U967 (N_967,N_499,N_523);
or U968 (N_968,N_700,N_323);
or U969 (N_969,N_642,N_3);
or U970 (N_970,N_520,N_183);
nand U971 (N_971,N_220,N_235);
and U972 (N_972,N_743,N_550);
or U973 (N_973,N_652,N_119);
or U974 (N_974,N_194,N_338);
and U975 (N_975,N_97,N_274);
nand U976 (N_976,N_723,N_352);
and U977 (N_977,N_672,N_133);
nand U978 (N_978,N_405,N_144);
nor U979 (N_979,N_454,N_30);
nand U980 (N_980,N_646,N_509);
or U981 (N_981,N_386,N_245);
nand U982 (N_982,N_595,N_705);
or U983 (N_983,N_671,N_682);
or U984 (N_984,N_452,N_273);
or U985 (N_985,N_711,N_99);
nand U986 (N_986,N_516,N_229);
or U987 (N_987,N_131,N_187);
nand U988 (N_988,N_585,N_222);
or U989 (N_989,N_462,N_83);
or U990 (N_990,N_544,N_537);
nand U991 (N_991,N_184,N_556);
nor U992 (N_992,N_261,N_665);
nor U993 (N_993,N_98,N_241);
nor U994 (N_994,N_419,N_267);
and U995 (N_995,N_300,N_606);
or U996 (N_996,N_521,N_239);
nor U997 (N_997,N_276,N_328);
and U998 (N_998,N_552,N_741);
and U999 (N_999,N_578,N_166);
and U1000 (N_1000,N_450,N_34);
and U1001 (N_1001,N_393,N_379);
nand U1002 (N_1002,N_553,N_367);
nand U1003 (N_1003,N_287,N_318);
or U1004 (N_1004,N_164,N_198);
nand U1005 (N_1005,N_738,N_275);
or U1006 (N_1006,N_486,N_721);
nor U1007 (N_1007,N_7,N_17);
nand U1008 (N_1008,N_271,N_342);
or U1009 (N_1009,N_497,N_369);
and U1010 (N_1010,N_588,N_668);
or U1011 (N_1011,N_256,N_431);
nand U1012 (N_1012,N_171,N_654);
and U1013 (N_1013,N_32,N_461);
or U1014 (N_1014,N_480,N_666);
nor U1015 (N_1015,N_246,N_72);
nor U1016 (N_1016,N_584,N_79);
nand U1017 (N_1017,N_11,N_15);
nor U1018 (N_1018,N_262,N_244);
or U1019 (N_1019,N_124,N_228);
or U1020 (N_1020,N_44,N_647);
nor U1021 (N_1021,N_353,N_430);
nand U1022 (N_1022,N_127,N_4);
nand U1023 (N_1023,N_392,N_316);
and U1024 (N_1024,N_686,N_47);
or U1025 (N_1025,N_243,N_303);
nand U1026 (N_1026,N_93,N_90);
xor U1027 (N_1027,N_530,N_539);
nand U1028 (N_1028,N_146,N_75);
nor U1029 (N_1029,N_96,N_421);
nor U1030 (N_1030,N_453,N_744);
nand U1031 (N_1031,N_88,N_41);
nand U1032 (N_1032,N_48,N_701);
or U1033 (N_1033,N_447,N_52);
nand U1034 (N_1034,N_429,N_40);
nand U1035 (N_1035,N_233,N_307);
or U1036 (N_1036,N_673,N_218);
nor U1037 (N_1037,N_91,N_709);
and U1038 (N_1038,N_112,N_481);
nor U1039 (N_1039,N_260,N_503);
nand U1040 (N_1040,N_456,N_693);
nand U1041 (N_1041,N_80,N_375);
nand U1042 (N_1042,N_525,N_488);
or U1043 (N_1043,N_746,N_558);
or U1044 (N_1044,N_625,N_298);
or U1045 (N_1045,N_29,N_25);
or U1046 (N_1046,N_670,N_77);
nor U1047 (N_1047,N_209,N_103);
xnor U1048 (N_1048,N_487,N_493);
nor U1049 (N_1049,N_583,N_254);
or U1050 (N_1050,N_82,N_114);
nor U1051 (N_1051,N_706,N_586);
nor U1052 (N_1052,N_417,N_363);
nor U1053 (N_1053,N_637,N_736);
nor U1054 (N_1054,N_36,N_314);
or U1055 (N_1055,N_158,N_591);
nor U1056 (N_1056,N_211,N_234);
nor U1057 (N_1057,N_190,N_710);
nor U1058 (N_1058,N_394,N_483);
nand U1059 (N_1059,N_560,N_718);
or U1060 (N_1060,N_16,N_51);
and U1061 (N_1061,N_89,N_354);
nand U1062 (N_1062,N_402,N_663);
nand U1063 (N_1063,N_210,N_597);
or U1064 (N_1064,N_643,N_703);
or U1065 (N_1065,N_370,N_532);
and U1066 (N_1066,N_615,N_87);
nor U1067 (N_1067,N_315,N_137);
and U1068 (N_1068,N_340,N_545);
and U1069 (N_1069,N_23,N_136);
and U1070 (N_1070,N_325,N_132);
and U1071 (N_1071,N_482,N_152);
nor U1072 (N_1072,N_151,N_380);
or U1073 (N_1073,N_212,N_415);
xor U1074 (N_1074,N_148,N_640);
nor U1075 (N_1075,N_333,N_156);
nand U1076 (N_1076,N_299,N_713);
nor U1077 (N_1077,N_92,N_382);
and U1078 (N_1078,N_305,N_106);
or U1079 (N_1079,N_734,N_216);
or U1080 (N_1080,N_575,N_259);
nor U1081 (N_1081,N_0,N_717);
or U1082 (N_1082,N_217,N_418);
nand U1083 (N_1083,N_381,N_491);
and U1084 (N_1084,N_150,N_230);
nand U1085 (N_1085,N_258,N_46);
nand U1086 (N_1086,N_206,N_485);
nand U1087 (N_1087,N_188,N_681);
nor U1088 (N_1088,N_120,N_542);
nand U1089 (N_1089,N_85,N_57);
and U1090 (N_1090,N_49,N_581);
or U1091 (N_1091,N_726,N_400);
nor U1092 (N_1092,N_579,N_662);
nand U1093 (N_1093,N_445,N_165);
and U1094 (N_1094,N_250,N_677);
nand U1095 (N_1095,N_242,N_629);
nand U1096 (N_1096,N_45,N_602);
or U1097 (N_1097,N_704,N_377);
nor U1098 (N_1098,N_248,N_60);
or U1099 (N_1099,N_74,N_78);
or U1100 (N_1100,N_596,N_424);
and U1101 (N_1101,N_387,N_366);
and U1102 (N_1102,N_658,N_374);
xnor U1103 (N_1103,N_477,N_37);
and U1104 (N_1104,N_515,N_518);
nor U1105 (N_1105,N_535,N_345);
nor U1106 (N_1106,N_364,N_163);
nand U1107 (N_1107,N_735,N_292);
nand U1108 (N_1108,N_622,N_348);
or U1109 (N_1109,N_135,N_510);
nor U1110 (N_1110,N_8,N_280);
nand U1111 (N_1111,N_722,N_645);
or U1112 (N_1112,N_747,N_716);
and U1113 (N_1113,N_641,N_117);
or U1114 (N_1114,N_727,N_555);
and U1115 (N_1115,N_145,N_24);
and U1116 (N_1116,N_68,N_594);
or U1117 (N_1117,N_592,N_725);
nor U1118 (N_1118,N_221,N_172);
nand U1119 (N_1119,N_167,N_748);
and U1120 (N_1120,N_433,N_696);
or U1121 (N_1121,N_205,N_249);
nor U1122 (N_1122,N_547,N_157);
or U1123 (N_1123,N_95,N_126);
or U1124 (N_1124,N_506,N_714);
or U1125 (N_1125,N_520,N_628);
and U1126 (N_1126,N_413,N_648);
or U1127 (N_1127,N_294,N_398);
nand U1128 (N_1128,N_645,N_284);
and U1129 (N_1129,N_18,N_721);
nor U1130 (N_1130,N_693,N_329);
nor U1131 (N_1131,N_579,N_205);
nand U1132 (N_1132,N_163,N_535);
nand U1133 (N_1133,N_629,N_483);
or U1134 (N_1134,N_252,N_62);
and U1135 (N_1135,N_521,N_314);
nor U1136 (N_1136,N_124,N_165);
nand U1137 (N_1137,N_484,N_478);
nand U1138 (N_1138,N_749,N_331);
or U1139 (N_1139,N_141,N_244);
or U1140 (N_1140,N_388,N_373);
nand U1141 (N_1141,N_646,N_156);
and U1142 (N_1142,N_644,N_74);
xnor U1143 (N_1143,N_628,N_265);
nand U1144 (N_1144,N_245,N_252);
or U1145 (N_1145,N_382,N_579);
nor U1146 (N_1146,N_665,N_26);
and U1147 (N_1147,N_44,N_549);
and U1148 (N_1148,N_313,N_383);
and U1149 (N_1149,N_569,N_472);
or U1150 (N_1150,N_651,N_539);
nand U1151 (N_1151,N_242,N_15);
and U1152 (N_1152,N_337,N_588);
nand U1153 (N_1153,N_5,N_27);
and U1154 (N_1154,N_13,N_342);
or U1155 (N_1155,N_669,N_336);
nor U1156 (N_1156,N_198,N_317);
nand U1157 (N_1157,N_553,N_651);
and U1158 (N_1158,N_106,N_668);
or U1159 (N_1159,N_197,N_371);
and U1160 (N_1160,N_486,N_203);
nor U1161 (N_1161,N_387,N_170);
or U1162 (N_1162,N_737,N_548);
nand U1163 (N_1163,N_50,N_153);
or U1164 (N_1164,N_237,N_190);
nor U1165 (N_1165,N_638,N_513);
nand U1166 (N_1166,N_365,N_27);
or U1167 (N_1167,N_260,N_392);
nand U1168 (N_1168,N_60,N_400);
and U1169 (N_1169,N_248,N_380);
nand U1170 (N_1170,N_202,N_323);
nor U1171 (N_1171,N_726,N_184);
nand U1172 (N_1172,N_282,N_684);
and U1173 (N_1173,N_739,N_571);
nand U1174 (N_1174,N_480,N_165);
nand U1175 (N_1175,N_586,N_58);
and U1176 (N_1176,N_540,N_440);
or U1177 (N_1177,N_151,N_729);
nand U1178 (N_1178,N_611,N_402);
and U1179 (N_1179,N_365,N_119);
and U1180 (N_1180,N_185,N_474);
or U1181 (N_1181,N_507,N_292);
nor U1182 (N_1182,N_640,N_498);
nand U1183 (N_1183,N_708,N_525);
nor U1184 (N_1184,N_640,N_730);
nand U1185 (N_1185,N_243,N_314);
and U1186 (N_1186,N_327,N_685);
or U1187 (N_1187,N_302,N_68);
nor U1188 (N_1188,N_291,N_124);
nand U1189 (N_1189,N_654,N_160);
nor U1190 (N_1190,N_9,N_467);
nand U1191 (N_1191,N_124,N_495);
and U1192 (N_1192,N_12,N_271);
or U1193 (N_1193,N_643,N_624);
or U1194 (N_1194,N_267,N_302);
nand U1195 (N_1195,N_485,N_312);
nor U1196 (N_1196,N_738,N_377);
or U1197 (N_1197,N_326,N_52);
or U1198 (N_1198,N_217,N_489);
or U1199 (N_1199,N_612,N_92);
and U1200 (N_1200,N_590,N_596);
or U1201 (N_1201,N_258,N_268);
or U1202 (N_1202,N_309,N_491);
nor U1203 (N_1203,N_47,N_238);
or U1204 (N_1204,N_674,N_361);
or U1205 (N_1205,N_413,N_408);
nand U1206 (N_1206,N_275,N_63);
nor U1207 (N_1207,N_486,N_639);
nor U1208 (N_1208,N_419,N_132);
or U1209 (N_1209,N_556,N_0);
nand U1210 (N_1210,N_607,N_340);
and U1211 (N_1211,N_300,N_527);
or U1212 (N_1212,N_115,N_632);
nand U1213 (N_1213,N_307,N_193);
nor U1214 (N_1214,N_272,N_512);
or U1215 (N_1215,N_679,N_141);
nor U1216 (N_1216,N_738,N_499);
or U1217 (N_1217,N_63,N_216);
nand U1218 (N_1218,N_246,N_308);
nand U1219 (N_1219,N_588,N_206);
and U1220 (N_1220,N_476,N_380);
nor U1221 (N_1221,N_412,N_317);
nand U1222 (N_1222,N_381,N_341);
or U1223 (N_1223,N_689,N_724);
or U1224 (N_1224,N_80,N_519);
nor U1225 (N_1225,N_115,N_725);
nor U1226 (N_1226,N_518,N_449);
nor U1227 (N_1227,N_661,N_514);
nand U1228 (N_1228,N_472,N_350);
and U1229 (N_1229,N_738,N_6);
and U1230 (N_1230,N_253,N_425);
nand U1231 (N_1231,N_540,N_398);
and U1232 (N_1232,N_237,N_395);
nor U1233 (N_1233,N_469,N_346);
and U1234 (N_1234,N_256,N_416);
or U1235 (N_1235,N_668,N_172);
nor U1236 (N_1236,N_379,N_135);
nand U1237 (N_1237,N_61,N_642);
or U1238 (N_1238,N_472,N_425);
nor U1239 (N_1239,N_91,N_707);
or U1240 (N_1240,N_27,N_603);
nand U1241 (N_1241,N_124,N_596);
nor U1242 (N_1242,N_597,N_194);
nor U1243 (N_1243,N_701,N_282);
nand U1244 (N_1244,N_615,N_587);
or U1245 (N_1245,N_326,N_422);
and U1246 (N_1246,N_19,N_145);
or U1247 (N_1247,N_554,N_569);
nand U1248 (N_1248,N_149,N_519);
nor U1249 (N_1249,N_706,N_238);
nand U1250 (N_1250,N_162,N_568);
nand U1251 (N_1251,N_564,N_123);
nor U1252 (N_1252,N_617,N_511);
and U1253 (N_1253,N_331,N_7);
nor U1254 (N_1254,N_596,N_692);
or U1255 (N_1255,N_134,N_749);
and U1256 (N_1256,N_309,N_144);
nor U1257 (N_1257,N_669,N_667);
or U1258 (N_1258,N_240,N_2);
or U1259 (N_1259,N_351,N_81);
nand U1260 (N_1260,N_202,N_493);
and U1261 (N_1261,N_571,N_228);
nor U1262 (N_1262,N_108,N_614);
nand U1263 (N_1263,N_210,N_214);
or U1264 (N_1264,N_670,N_233);
nand U1265 (N_1265,N_517,N_748);
or U1266 (N_1266,N_562,N_318);
and U1267 (N_1267,N_379,N_251);
and U1268 (N_1268,N_125,N_702);
and U1269 (N_1269,N_748,N_213);
and U1270 (N_1270,N_637,N_8);
and U1271 (N_1271,N_430,N_647);
nand U1272 (N_1272,N_327,N_120);
nand U1273 (N_1273,N_429,N_190);
nor U1274 (N_1274,N_632,N_499);
nand U1275 (N_1275,N_743,N_185);
and U1276 (N_1276,N_374,N_212);
nand U1277 (N_1277,N_289,N_8);
and U1278 (N_1278,N_565,N_197);
nand U1279 (N_1279,N_702,N_315);
or U1280 (N_1280,N_321,N_34);
nand U1281 (N_1281,N_105,N_438);
nand U1282 (N_1282,N_712,N_449);
or U1283 (N_1283,N_205,N_6);
nand U1284 (N_1284,N_404,N_528);
and U1285 (N_1285,N_362,N_119);
and U1286 (N_1286,N_501,N_198);
or U1287 (N_1287,N_108,N_369);
and U1288 (N_1288,N_289,N_434);
and U1289 (N_1289,N_296,N_42);
or U1290 (N_1290,N_156,N_93);
or U1291 (N_1291,N_122,N_443);
nand U1292 (N_1292,N_628,N_568);
or U1293 (N_1293,N_459,N_363);
nand U1294 (N_1294,N_80,N_532);
and U1295 (N_1295,N_545,N_99);
or U1296 (N_1296,N_395,N_111);
and U1297 (N_1297,N_563,N_103);
and U1298 (N_1298,N_503,N_448);
and U1299 (N_1299,N_143,N_383);
or U1300 (N_1300,N_664,N_374);
nand U1301 (N_1301,N_162,N_702);
nor U1302 (N_1302,N_86,N_1);
and U1303 (N_1303,N_118,N_532);
and U1304 (N_1304,N_145,N_260);
or U1305 (N_1305,N_291,N_131);
and U1306 (N_1306,N_552,N_213);
or U1307 (N_1307,N_519,N_590);
and U1308 (N_1308,N_454,N_457);
nor U1309 (N_1309,N_590,N_507);
nor U1310 (N_1310,N_598,N_195);
nand U1311 (N_1311,N_423,N_344);
and U1312 (N_1312,N_80,N_182);
or U1313 (N_1313,N_8,N_174);
or U1314 (N_1314,N_730,N_287);
nand U1315 (N_1315,N_719,N_243);
and U1316 (N_1316,N_656,N_165);
nor U1317 (N_1317,N_733,N_415);
nand U1318 (N_1318,N_650,N_168);
nand U1319 (N_1319,N_423,N_533);
nand U1320 (N_1320,N_713,N_182);
or U1321 (N_1321,N_116,N_534);
nor U1322 (N_1322,N_23,N_168);
nand U1323 (N_1323,N_260,N_200);
nor U1324 (N_1324,N_396,N_659);
nand U1325 (N_1325,N_518,N_418);
nor U1326 (N_1326,N_332,N_426);
nand U1327 (N_1327,N_498,N_674);
nor U1328 (N_1328,N_272,N_194);
nand U1329 (N_1329,N_681,N_131);
nor U1330 (N_1330,N_183,N_686);
nor U1331 (N_1331,N_216,N_367);
nor U1332 (N_1332,N_496,N_449);
nand U1333 (N_1333,N_181,N_658);
or U1334 (N_1334,N_22,N_403);
nand U1335 (N_1335,N_292,N_394);
and U1336 (N_1336,N_116,N_13);
nand U1337 (N_1337,N_492,N_14);
or U1338 (N_1338,N_89,N_83);
or U1339 (N_1339,N_198,N_327);
or U1340 (N_1340,N_41,N_652);
and U1341 (N_1341,N_700,N_658);
xor U1342 (N_1342,N_645,N_459);
nand U1343 (N_1343,N_0,N_3);
nor U1344 (N_1344,N_44,N_642);
nor U1345 (N_1345,N_85,N_267);
and U1346 (N_1346,N_113,N_745);
or U1347 (N_1347,N_46,N_182);
nand U1348 (N_1348,N_50,N_689);
nand U1349 (N_1349,N_256,N_254);
nor U1350 (N_1350,N_146,N_85);
or U1351 (N_1351,N_702,N_280);
and U1352 (N_1352,N_498,N_585);
or U1353 (N_1353,N_550,N_320);
and U1354 (N_1354,N_151,N_711);
nor U1355 (N_1355,N_587,N_422);
and U1356 (N_1356,N_726,N_696);
nor U1357 (N_1357,N_428,N_283);
nand U1358 (N_1358,N_467,N_68);
nand U1359 (N_1359,N_403,N_261);
nand U1360 (N_1360,N_256,N_298);
and U1361 (N_1361,N_177,N_235);
or U1362 (N_1362,N_598,N_471);
and U1363 (N_1363,N_223,N_622);
nor U1364 (N_1364,N_199,N_244);
nor U1365 (N_1365,N_235,N_27);
nor U1366 (N_1366,N_288,N_445);
and U1367 (N_1367,N_296,N_72);
or U1368 (N_1368,N_681,N_376);
nor U1369 (N_1369,N_53,N_189);
and U1370 (N_1370,N_553,N_301);
or U1371 (N_1371,N_553,N_659);
or U1372 (N_1372,N_410,N_318);
and U1373 (N_1373,N_703,N_533);
or U1374 (N_1374,N_720,N_737);
and U1375 (N_1375,N_474,N_493);
nand U1376 (N_1376,N_715,N_439);
or U1377 (N_1377,N_717,N_169);
and U1378 (N_1378,N_201,N_439);
or U1379 (N_1379,N_79,N_350);
nand U1380 (N_1380,N_170,N_103);
and U1381 (N_1381,N_667,N_276);
nor U1382 (N_1382,N_529,N_624);
or U1383 (N_1383,N_569,N_173);
nor U1384 (N_1384,N_122,N_524);
or U1385 (N_1385,N_722,N_100);
and U1386 (N_1386,N_63,N_272);
and U1387 (N_1387,N_234,N_736);
and U1388 (N_1388,N_37,N_703);
nor U1389 (N_1389,N_383,N_542);
nor U1390 (N_1390,N_164,N_315);
nor U1391 (N_1391,N_489,N_78);
nor U1392 (N_1392,N_399,N_598);
or U1393 (N_1393,N_301,N_498);
and U1394 (N_1394,N_579,N_736);
nor U1395 (N_1395,N_536,N_463);
nand U1396 (N_1396,N_344,N_48);
nor U1397 (N_1397,N_523,N_393);
nor U1398 (N_1398,N_342,N_181);
nor U1399 (N_1399,N_529,N_306);
and U1400 (N_1400,N_550,N_527);
or U1401 (N_1401,N_545,N_748);
nand U1402 (N_1402,N_339,N_478);
nand U1403 (N_1403,N_655,N_368);
and U1404 (N_1404,N_386,N_4);
nand U1405 (N_1405,N_238,N_581);
or U1406 (N_1406,N_726,N_251);
nor U1407 (N_1407,N_346,N_655);
nand U1408 (N_1408,N_509,N_245);
nor U1409 (N_1409,N_78,N_351);
nand U1410 (N_1410,N_708,N_10);
nand U1411 (N_1411,N_580,N_105);
nor U1412 (N_1412,N_36,N_159);
nand U1413 (N_1413,N_668,N_178);
nand U1414 (N_1414,N_311,N_682);
or U1415 (N_1415,N_126,N_553);
nand U1416 (N_1416,N_337,N_334);
and U1417 (N_1417,N_594,N_744);
or U1418 (N_1418,N_218,N_72);
nand U1419 (N_1419,N_4,N_708);
nor U1420 (N_1420,N_407,N_447);
nor U1421 (N_1421,N_456,N_282);
nor U1422 (N_1422,N_252,N_650);
nor U1423 (N_1423,N_430,N_77);
nand U1424 (N_1424,N_670,N_433);
nor U1425 (N_1425,N_487,N_298);
nand U1426 (N_1426,N_107,N_286);
nand U1427 (N_1427,N_692,N_295);
nand U1428 (N_1428,N_356,N_572);
or U1429 (N_1429,N_201,N_657);
and U1430 (N_1430,N_439,N_551);
nor U1431 (N_1431,N_476,N_177);
nand U1432 (N_1432,N_671,N_626);
or U1433 (N_1433,N_452,N_311);
and U1434 (N_1434,N_512,N_52);
nor U1435 (N_1435,N_142,N_247);
nor U1436 (N_1436,N_566,N_492);
and U1437 (N_1437,N_512,N_35);
nand U1438 (N_1438,N_244,N_486);
nor U1439 (N_1439,N_57,N_369);
nand U1440 (N_1440,N_529,N_648);
or U1441 (N_1441,N_61,N_367);
nor U1442 (N_1442,N_256,N_42);
nand U1443 (N_1443,N_364,N_428);
or U1444 (N_1444,N_496,N_319);
nand U1445 (N_1445,N_741,N_244);
and U1446 (N_1446,N_524,N_673);
and U1447 (N_1447,N_297,N_84);
nor U1448 (N_1448,N_373,N_354);
nand U1449 (N_1449,N_424,N_406);
nor U1450 (N_1450,N_108,N_251);
and U1451 (N_1451,N_306,N_447);
or U1452 (N_1452,N_671,N_350);
or U1453 (N_1453,N_629,N_487);
nand U1454 (N_1454,N_657,N_224);
nand U1455 (N_1455,N_605,N_240);
nand U1456 (N_1456,N_79,N_642);
nor U1457 (N_1457,N_389,N_168);
or U1458 (N_1458,N_578,N_193);
nor U1459 (N_1459,N_688,N_424);
nand U1460 (N_1460,N_366,N_57);
and U1461 (N_1461,N_71,N_60);
nand U1462 (N_1462,N_592,N_362);
nor U1463 (N_1463,N_601,N_474);
nand U1464 (N_1464,N_456,N_434);
nor U1465 (N_1465,N_713,N_288);
nor U1466 (N_1466,N_663,N_731);
nand U1467 (N_1467,N_343,N_406);
nand U1468 (N_1468,N_532,N_38);
nand U1469 (N_1469,N_404,N_225);
or U1470 (N_1470,N_150,N_29);
nand U1471 (N_1471,N_578,N_695);
or U1472 (N_1472,N_204,N_285);
nand U1473 (N_1473,N_547,N_143);
and U1474 (N_1474,N_355,N_704);
nor U1475 (N_1475,N_482,N_638);
nor U1476 (N_1476,N_662,N_659);
nor U1477 (N_1477,N_62,N_428);
and U1478 (N_1478,N_607,N_701);
and U1479 (N_1479,N_234,N_443);
and U1480 (N_1480,N_702,N_529);
nor U1481 (N_1481,N_569,N_391);
nor U1482 (N_1482,N_232,N_510);
and U1483 (N_1483,N_725,N_15);
nor U1484 (N_1484,N_671,N_653);
and U1485 (N_1485,N_301,N_257);
or U1486 (N_1486,N_442,N_545);
nand U1487 (N_1487,N_278,N_309);
and U1488 (N_1488,N_643,N_336);
or U1489 (N_1489,N_138,N_22);
and U1490 (N_1490,N_89,N_252);
and U1491 (N_1491,N_702,N_522);
nor U1492 (N_1492,N_7,N_73);
or U1493 (N_1493,N_701,N_622);
and U1494 (N_1494,N_118,N_707);
and U1495 (N_1495,N_450,N_247);
nand U1496 (N_1496,N_25,N_448);
or U1497 (N_1497,N_545,N_389);
nor U1498 (N_1498,N_739,N_565);
nor U1499 (N_1499,N_404,N_214);
nand U1500 (N_1500,N_1173,N_1136);
nand U1501 (N_1501,N_1307,N_941);
nor U1502 (N_1502,N_982,N_1343);
nand U1503 (N_1503,N_1061,N_882);
or U1504 (N_1504,N_769,N_1110);
nor U1505 (N_1505,N_816,N_1432);
and U1506 (N_1506,N_1243,N_1284);
nand U1507 (N_1507,N_1032,N_1232);
nand U1508 (N_1508,N_1141,N_946);
or U1509 (N_1509,N_1049,N_857);
nand U1510 (N_1510,N_1121,N_950);
nor U1511 (N_1511,N_1286,N_873);
nand U1512 (N_1512,N_1437,N_1490);
and U1513 (N_1513,N_845,N_1287);
or U1514 (N_1514,N_1394,N_1108);
or U1515 (N_1515,N_1280,N_1208);
nand U1516 (N_1516,N_1444,N_761);
and U1517 (N_1517,N_1309,N_1400);
nor U1518 (N_1518,N_1326,N_977);
nand U1519 (N_1519,N_1460,N_848);
nand U1520 (N_1520,N_965,N_752);
nor U1521 (N_1521,N_1306,N_1419);
nand U1522 (N_1522,N_869,N_1072);
nor U1523 (N_1523,N_1001,N_1106);
and U1524 (N_1524,N_1476,N_993);
or U1525 (N_1525,N_1092,N_1347);
nor U1526 (N_1526,N_1127,N_1491);
or U1527 (N_1527,N_753,N_1204);
nand U1528 (N_1528,N_992,N_1494);
nand U1529 (N_1529,N_1041,N_874);
and U1530 (N_1530,N_1148,N_971);
nor U1531 (N_1531,N_1089,N_922);
nand U1532 (N_1532,N_1448,N_1354);
nand U1533 (N_1533,N_1051,N_1132);
and U1534 (N_1534,N_1469,N_1150);
nor U1535 (N_1535,N_1238,N_1087);
nand U1536 (N_1536,N_1395,N_1119);
nor U1537 (N_1537,N_859,N_1158);
nand U1538 (N_1538,N_1386,N_885);
nand U1539 (N_1539,N_1194,N_1384);
and U1540 (N_1540,N_1240,N_1359);
or U1541 (N_1541,N_1472,N_1095);
nand U1542 (N_1542,N_1477,N_961);
nand U1543 (N_1543,N_1278,N_1063);
and U1544 (N_1544,N_959,N_1192);
and U1545 (N_1545,N_1486,N_1048);
nand U1546 (N_1546,N_853,N_1461);
or U1547 (N_1547,N_1138,N_1376);
xor U1548 (N_1548,N_870,N_956);
and U1549 (N_1549,N_773,N_1038);
and U1550 (N_1550,N_823,N_1266);
and U1551 (N_1551,N_804,N_1126);
or U1552 (N_1552,N_1210,N_1454);
or U1553 (N_1553,N_779,N_902);
nor U1554 (N_1554,N_1449,N_1219);
nor U1555 (N_1555,N_967,N_948);
nor U1556 (N_1556,N_962,N_1164);
and U1557 (N_1557,N_1157,N_1231);
nand U1558 (N_1558,N_1319,N_973);
and U1559 (N_1559,N_1271,N_1047);
and U1560 (N_1560,N_1004,N_1393);
xor U1561 (N_1561,N_847,N_1062);
nor U1562 (N_1562,N_1371,N_796);
nand U1563 (N_1563,N_807,N_891);
and U1564 (N_1564,N_999,N_1383);
nand U1565 (N_1565,N_1305,N_972);
or U1566 (N_1566,N_760,N_924);
nor U1567 (N_1567,N_1470,N_1482);
nand U1568 (N_1568,N_1235,N_1170);
or U1569 (N_1569,N_1188,N_1429);
nand U1570 (N_1570,N_1058,N_1211);
or U1571 (N_1571,N_1073,N_822);
and U1572 (N_1572,N_1253,N_875);
nand U1573 (N_1573,N_1064,N_783);
nor U1574 (N_1574,N_1369,N_1060);
or U1575 (N_1575,N_1279,N_1205);
and U1576 (N_1576,N_1338,N_1233);
nor U1577 (N_1577,N_1222,N_1292);
nor U1578 (N_1578,N_1328,N_888);
and U1579 (N_1579,N_1070,N_1435);
nand U1580 (N_1580,N_1375,N_996);
nand U1581 (N_1581,N_839,N_1399);
or U1582 (N_1582,N_981,N_878);
nand U1583 (N_1583,N_1056,N_871);
and U1584 (N_1584,N_815,N_1427);
nor U1585 (N_1585,N_887,N_1464);
nor U1586 (N_1586,N_1252,N_1363);
and U1587 (N_1587,N_945,N_889);
nand U1588 (N_1588,N_810,N_1090);
nor U1589 (N_1589,N_1273,N_1000);
nor U1590 (N_1590,N_1116,N_884);
or U1591 (N_1591,N_1496,N_813);
nand U1592 (N_1592,N_1011,N_1484);
nor U1593 (N_1593,N_1183,N_883);
nand U1594 (N_1594,N_1290,N_1250);
or U1595 (N_1595,N_1167,N_1411);
and U1596 (N_1596,N_792,N_1327);
nand U1597 (N_1597,N_952,N_830);
nand U1598 (N_1598,N_1337,N_1050);
nand U1599 (N_1599,N_890,N_1123);
nor U1600 (N_1600,N_1076,N_1035);
and U1601 (N_1601,N_1341,N_1228);
nor U1602 (N_1602,N_1163,N_997);
nand U1603 (N_1603,N_897,N_1313);
nand U1604 (N_1604,N_1080,N_1220);
and U1605 (N_1605,N_1331,N_886);
and U1606 (N_1606,N_1362,N_1440);
nor U1607 (N_1607,N_949,N_877);
or U1608 (N_1608,N_867,N_1016);
and U1609 (N_1609,N_1459,N_1356);
or U1610 (N_1610,N_1350,N_1390);
or U1611 (N_1611,N_1332,N_1109);
or U1612 (N_1612,N_1002,N_1206);
and U1613 (N_1613,N_1247,N_798);
and U1614 (N_1614,N_833,N_855);
nand U1615 (N_1615,N_940,N_1033);
nand U1616 (N_1616,N_1014,N_800);
nand U1617 (N_1617,N_1291,N_1135);
or U1618 (N_1618,N_1401,N_844);
nor U1619 (N_1619,N_821,N_942);
or U1620 (N_1620,N_1245,N_1415);
nor U1621 (N_1621,N_789,N_842);
xnor U1622 (N_1622,N_1254,N_1387);
and U1623 (N_1623,N_1042,N_1052);
nor U1624 (N_1624,N_976,N_817);
and U1625 (N_1625,N_1093,N_1137);
nor U1626 (N_1626,N_1006,N_918);
xor U1627 (N_1627,N_1368,N_768);
and U1628 (N_1628,N_1181,N_812);
or U1629 (N_1629,N_1406,N_1277);
or U1630 (N_1630,N_1430,N_963);
nand U1631 (N_1631,N_1264,N_814);
nand U1632 (N_1632,N_1481,N_1352);
and U1633 (N_1633,N_1385,N_1068);
or U1634 (N_1634,N_980,N_1324);
or U1635 (N_1635,N_1217,N_1404);
nor U1636 (N_1636,N_767,N_849);
nor U1637 (N_1637,N_958,N_1340);
nor U1638 (N_1638,N_966,N_1353);
nand U1639 (N_1639,N_1334,N_1071);
nand U1640 (N_1640,N_1227,N_1021);
or U1641 (N_1641,N_1096,N_1160);
nand U1642 (N_1642,N_910,N_876);
nor U1643 (N_1643,N_1423,N_1298);
and U1644 (N_1644,N_1100,N_1312);
or U1645 (N_1645,N_1237,N_1045);
nor U1646 (N_1646,N_818,N_1480);
and U1647 (N_1647,N_1151,N_868);
nand U1648 (N_1648,N_1224,N_1314);
and U1649 (N_1649,N_1302,N_1012);
nor U1650 (N_1650,N_1413,N_943);
and U1651 (N_1651,N_1318,N_1294);
nor U1652 (N_1652,N_1445,N_906);
nand U1653 (N_1653,N_947,N_1226);
nand U1654 (N_1654,N_1107,N_1007);
and U1655 (N_1655,N_793,N_1300);
or U1656 (N_1656,N_933,N_1200);
nor U1657 (N_1657,N_1149,N_1124);
xnor U1658 (N_1658,N_1169,N_791);
nor U1659 (N_1659,N_1357,N_1410);
and U1660 (N_1660,N_1140,N_819);
nand U1661 (N_1661,N_1317,N_1172);
nand U1662 (N_1662,N_954,N_1147);
nor U1663 (N_1663,N_923,N_1408);
or U1664 (N_1664,N_851,N_1168);
nand U1665 (N_1665,N_1251,N_1407);
or U1666 (N_1666,N_829,N_1133);
or U1667 (N_1667,N_892,N_1130);
or U1668 (N_1668,N_1055,N_916);
and U1669 (N_1669,N_1479,N_998);
xnor U1670 (N_1670,N_802,N_1207);
and U1671 (N_1671,N_1161,N_1420);
and U1672 (N_1672,N_1417,N_1308);
nor U1673 (N_1673,N_1255,N_1203);
and U1674 (N_1674,N_1462,N_1199);
nor U1675 (N_1675,N_1295,N_1128);
or U1676 (N_1676,N_785,N_1179);
nand U1677 (N_1677,N_1180,N_856);
and U1678 (N_1678,N_1463,N_1370);
or U1679 (N_1679,N_935,N_1493);
nand U1680 (N_1680,N_1256,N_1483);
or U1681 (N_1681,N_836,N_979);
and U1682 (N_1682,N_1025,N_1081);
nand U1683 (N_1683,N_1209,N_1225);
and U1684 (N_1684,N_903,N_852);
or U1685 (N_1685,N_824,N_1113);
or U1686 (N_1686,N_1084,N_939);
or U1687 (N_1687,N_860,N_1325);
nor U1688 (N_1688,N_809,N_1036);
nor U1689 (N_1689,N_1003,N_1452);
or U1690 (N_1690,N_1330,N_1391);
nand U1691 (N_1691,N_1186,N_975);
or U1692 (N_1692,N_1193,N_983);
nor U1693 (N_1693,N_1174,N_1441);
nand U1694 (N_1694,N_1187,N_1043);
nand U1695 (N_1695,N_1182,N_1131);
nand U1696 (N_1696,N_1274,N_1178);
or U1697 (N_1697,N_919,N_896);
nor U1698 (N_1698,N_1453,N_1165);
nor U1699 (N_1699,N_1267,N_1372);
nor U1700 (N_1700,N_994,N_901);
nand U1701 (N_1701,N_1336,N_1289);
nand U1702 (N_1702,N_1465,N_854);
or U1703 (N_1703,N_1241,N_1458);
and U1704 (N_1704,N_895,N_827);
nor U1705 (N_1705,N_1351,N_1299);
nor U1706 (N_1706,N_1120,N_1424);
and U1707 (N_1707,N_808,N_1425);
or U1708 (N_1708,N_970,N_1190);
nor U1709 (N_1709,N_1310,N_1059);
nand U1710 (N_1710,N_1155,N_1077);
or U1711 (N_1711,N_1360,N_1366);
and U1712 (N_1712,N_1497,N_1322);
nor U1713 (N_1713,N_1022,N_850);
or U1714 (N_1714,N_762,N_1345);
or U1715 (N_1715,N_1349,N_930);
and U1716 (N_1716,N_1171,N_1177);
or U1717 (N_1717,N_1303,N_1297);
or U1718 (N_1718,N_1339,N_825);
nor U1719 (N_1719,N_1456,N_913);
nor U1720 (N_1720,N_1378,N_1379);
nand U1721 (N_1721,N_1214,N_898);
or U1722 (N_1722,N_1315,N_838);
nand U1723 (N_1723,N_938,N_1083);
nor U1724 (N_1724,N_1159,N_1134);
and U1725 (N_1725,N_1422,N_1196);
or U1726 (N_1726,N_1215,N_1078);
nand U1727 (N_1727,N_1099,N_828);
and U1728 (N_1728,N_1288,N_1398);
xor U1729 (N_1729,N_832,N_1474);
nor U1730 (N_1730,N_757,N_861);
nor U1731 (N_1731,N_840,N_879);
nand U1732 (N_1732,N_1487,N_778);
and U1733 (N_1733,N_1154,N_1005);
or U1734 (N_1734,N_784,N_986);
or U1735 (N_1735,N_1402,N_968);
and U1736 (N_1736,N_863,N_1097);
and U1737 (N_1737,N_912,N_835);
nor U1738 (N_1738,N_1129,N_1023);
and U1739 (N_1739,N_1018,N_1248);
and U1740 (N_1740,N_1365,N_1166);
or U1741 (N_1741,N_1316,N_1443);
or U1742 (N_1742,N_1189,N_881);
nand U1743 (N_1743,N_786,N_1020);
and U1744 (N_1744,N_990,N_771);
or U1745 (N_1745,N_1091,N_758);
nor U1746 (N_1746,N_1367,N_1355);
nand U1747 (N_1747,N_843,N_1028);
or U1748 (N_1748,N_1431,N_1320);
or U1749 (N_1749,N_900,N_1030);
nand U1750 (N_1750,N_1088,N_1094);
nand U1751 (N_1751,N_894,N_1201);
nor U1752 (N_1752,N_1118,N_1105);
or U1753 (N_1753,N_1466,N_1333);
or U1754 (N_1754,N_1008,N_1373);
and U1755 (N_1755,N_1115,N_1162);
nor U1756 (N_1756,N_989,N_1428);
or U1757 (N_1757,N_1074,N_1268);
nand U1758 (N_1758,N_905,N_1475);
and U1759 (N_1759,N_806,N_1037);
nor U1760 (N_1760,N_775,N_1382);
nor U1761 (N_1761,N_770,N_907);
and U1762 (N_1762,N_1156,N_788);
nand U1763 (N_1763,N_1184,N_1457);
nand U1764 (N_1764,N_1380,N_1066);
or U1765 (N_1765,N_1467,N_1344);
or U1766 (N_1766,N_1485,N_1389);
nand U1767 (N_1767,N_826,N_1010);
nor U1768 (N_1768,N_1489,N_936);
nor U1769 (N_1769,N_801,N_1293);
or U1770 (N_1770,N_1381,N_974);
and U1771 (N_1771,N_858,N_1450);
and U1772 (N_1772,N_820,N_1392);
or U1773 (N_1773,N_797,N_1143);
and U1774 (N_1774,N_1262,N_1122);
nor U1775 (N_1775,N_991,N_1447);
and U1776 (N_1776,N_1239,N_1438);
and U1777 (N_1777,N_1009,N_1054);
nor U1778 (N_1778,N_1285,N_1434);
or U1779 (N_1779,N_1259,N_764);
nand U1780 (N_1780,N_1451,N_1125);
or U1781 (N_1781,N_787,N_925);
or U1782 (N_1782,N_834,N_1348);
nor U1783 (N_1783,N_1471,N_1246);
and U1784 (N_1784,N_1195,N_799);
and U1785 (N_1785,N_1202,N_1358);
nand U1786 (N_1786,N_1436,N_1213);
nand U1787 (N_1787,N_777,N_1034);
nor U1788 (N_1788,N_1269,N_1258);
nand U1789 (N_1789,N_1283,N_1426);
or U1790 (N_1790,N_1153,N_987);
nand U1791 (N_1791,N_759,N_1185);
nor U1792 (N_1792,N_1176,N_926);
and U1793 (N_1793,N_1495,N_1396);
and U1794 (N_1794,N_751,N_1017);
or U1795 (N_1795,N_1191,N_951);
or U1796 (N_1796,N_1069,N_1364);
or U1797 (N_1797,N_1329,N_1029);
nand U1798 (N_1798,N_1242,N_1103);
or U1799 (N_1799,N_1142,N_795);
or U1800 (N_1800,N_774,N_1044);
nor U1801 (N_1801,N_1403,N_1152);
or U1802 (N_1802,N_846,N_1114);
nand U1803 (N_1803,N_780,N_776);
nor U1804 (N_1804,N_1374,N_1388);
and U1805 (N_1805,N_1412,N_1230);
nor U1806 (N_1806,N_1019,N_927);
nor U1807 (N_1807,N_955,N_1272);
or U1808 (N_1808,N_929,N_1229);
and U1809 (N_1809,N_1085,N_964);
or U1810 (N_1810,N_1102,N_969);
nand U1811 (N_1811,N_1296,N_862);
nand U1812 (N_1812,N_1473,N_1468);
and U1813 (N_1813,N_1053,N_1065);
and U1814 (N_1814,N_1104,N_1086);
nand U1815 (N_1815,N_932,N_756);
nor U1816 (N_1816,N_937,N_1197);
and U1817 (N_1817,N_957,N_914);
and U1818 (N_1818,N_934,N_931);
and U1819 (N_1819,N_1175,N_1079);
or U1820 (N_1820,N_1488,N_803);
and U1821 (N_1821,N_754,N_1498);
nor U1822 (N_1822,N_995,N_1244);
nand U1823 (N_1823,N_1478,N_1027);
nand U1824 (N_1824,N_1263,N_1015);
and U1825 (N_1825,N_921,N_1013);
and U1826 (N_1826,N_1433,N_1101);
nand U1827 (N_1827,N_872,N_1311);
nor U1828 (N_1828,N_1067,N_899);
nand U1829 (N_1829,N_1026,N_1144);
xor U1830 (N_1830,N_1046,N_837);
nor U1831 (N_1831,N_1346,N_1075);
and U1832 (N_1832,N_765,N_1323);
or U1833 (N_1833,N_790,N_865);
or U1834 (N_1834,N_1057,N_1377);
xor U1835 (N_1835,N_1282,N_1216);
nand U1836 (N_1836,N_1098,N_953);
or U1837 (N_1837,N_1117,N_1223);
or U1838 (N_1838,N_1261,N_831);
nor U1839 (N_1839,N_1257,N_984);
and U1840 (N_1840,N_1301,N_794);
and U1841 (N_1841,N_1418,N_1236);
xnor U1842 (N_1842,N_1146,N_1342);
and U1843 (N_1843,N_782,N_1335);
nor U1844 (N_1844,N_1024,N_755);
or U1845 (N_1845,N_1275,N_928);
and U1846 (N_1846,N_1492,N_909);
nand U1847 (N_1847,N_1499,N_1397);
or U1848 (N_1848,N_1260,N_1031);
nor U1849 (N_1849,N_960,N_763);
and U1850 (N_1850,N_985,N_920);
or U1851 (N_1851,N_1361,N_1455);
nand U1852 (N_1852,N_911,N_1270);
and U1853 (N_1853,N_880,N_1304);
nor U1854 (N_1854,N_1416,N_1139);
and U1855 (N_1855,N_750,N_1112);
nor U1856 (N_1856,N_841,N_944);
nand U1857 (N_1857,N_893,N_864);
nand U1858 (N_1858,N_772,N_1409);
and U1859 (N_1859,N_1145,N_1321);
and U1860 (N_1860,N_1446,N_1218);
or U1861 (N_1861,N_781,N_1198);
and U1862 (N_1862,N_1265,N_1442);
nand U1863 (N_1863,N_1111,N_766);
nor U1864 (N_1864,N_1234,N_1405);
or U1865 (N_1865,N_1249,N_805);
nor U1866 (N_1866,N_1212,N_988);
nor U1867 (N_1867,N_1421,N_1414);
nor U1868 (N_1868,N_1082,N_908);
nand U1869 (N_1869,N_978,N_1276);
or U1870 (N_1870,N_917,N_1039);
xor U1871 (N_1871,N_1040,N_866);
nor U1872 (N_1872,N_1221,N_1281);
and U1873 (N_1873,N_915,N_904);
and U1874 (N_1874,N_1439,N_811);
nand U1875 (N_1875,N_830,N_1277);
nor U1876 (N_1876,N_1189,N_1018);
nand U1877 (N_1877,N_1353,N_1470);
nor U1878 (N_1878,N_875,N_831);
xor U1879 (N_1879,N_963,N_932);
nand U1880 (N_1880,N_1484,N_1176);
or U1881 (N_1881,N_971,N_1016);
nor U1882 (N_1882,N_1096,N_1080);
and U1883 (N_1883,N_794,N_1119);
nand U1884 (N_1884,N_1249,N_1008);
nor U1885 (N_1885,N_846,N_1280);
or U1886 (N_1886,N_1230,N_1415);
nand U1887 (N_1887,N_1340,N_1319);
nor U1888 (N_1888,N_864,N_1286);
and U1889 (N_1889,N_864,N_968);
or U1890 (N_1890,N_891,N_1443);
nor U1891 (N_1891,N_994,N_1127);
or U1892 (N_1892,N_1165,N_1129);
or U1893 (N_1893,N_1132,N_1047);
or U1894 (N_1894,N_1157,N_1362);
nor U1895 (N_1895,N_830,N_960);
nand U1896 (N_1896,N_892,N_987);
nand U1897 (N_1897,N_1300,N_1385);
and U1898 (N_1898,N_798,N_1352);
nor U1899 (N_1899,N_1328,N_958);
or U1900 (N_1900,N_805,N_1042);
or U1901 (N_1901,N_1318,N_938);
and U1902 (N_1902,N_794,N_1490);
nor U1903 (N_1903,N_986,N_1023);
or U1904 (N_1904,N_1091,N_920);
and U1905 (N_1905,N_1298,N_915);
nand U1906 (N_1906,N_862,N_1442);
nor U1907 (N_1907,N_1336,N_1176);
nor U1908 (N_1908,N_830,N_945);
nor U1909 (N_1909,N_837,N_1400);
nor U1910 (N_1910,N_1292,N_975);
and U1911 (N_1911,N_1363,N_974);
and U1912 (N_1912,N_1374,N_906);
and U1913 (N_1913,N_1428,N_1150);
nor U1914 (N_1914,N_1460,N_777);
nor U1915 (N_1915,N_1464,N_864);
and U1916 (N_1916,N_1184,N_1245);
nor U1917 (N_1917,N_1190,N_1059);
or U1918 (N_1918,N_1212,N_1029);
nand U1919 (N_1919,N_1188,N_804);
nand U1920 (N_1920,N_1429,N_1063);
and U1921 (N_1921,N_988,N_1159);
nor U1922 (N_1922,N_762,N_1333);
or U1923 (N_1923,N_1177,N_900);
nor U1924 (N_1924,N_831,N_1183);
nor U1925 (N_1925,N_1449,N_939);
or U1926 (N_1926,N_1116,N_1018);
or U1927 (N_1927,N_944,N_1197);
and U1928 (N_1928,N_1447,N_851);
and U1929 (N_1929,N_1100,N_1471);
or U1930 (N_1930,N_1436,N_1158);
nand U1931 (N_1931,N_1162,N_974);
nand U1932 (N_1932,N_1408,N_1280);
nand U1933 (N_1933,N_1339,N_1426);
and U1934 (N_1934,N_1275,N_810);
and U1935 (N_1935,N_861,N_881);
or U1936 (N_1936,N_1414,N_798);
and U1937 (N_1937,N_1427,N_1012);
nand U1938 (N_1938,N_902,N_1169);
nand U1939 (N_1939,N_1485,N_880);
nand U1940 (N_1940,N_1224,N_1380);
nor U1941 (N_1941,N_1210,N_1411);
or U1942 (N_1942,N_1377,N_1093);
or U1943 (N_1943,N_884,N_1150);
or U1944 (N_1944,N_1326,N_1099);
and U1945 (N_1945,N_1339,N_947);
nand U1946 (N_1946,N_871,N_1244);
nor U1947 (N_1947,N_912,N_1058);
nor U1948 (N_1948,N_1352,N_799);
nor U1949 (N_1949,N_1257,N_1024);
nand U1950 (N_1950,N_1006,N_1058);
nand U1951 (N_1951,N_1470,N_1352);
and U1952 (N_1952,N_1419,N_833);
nor U1953 (N_1953,N_1295,N_1473);
nor U1954 (N_1954,N_1459,N_904);
nor U1955 (N_1955,N_1337,N_1262);
and U1956 (N_1956,N_1345,N_837);
or U1957 (N_1957,N_1071,N_1429);
nand U1958 (N_1958,N_1013,N_1296);
nor U1959 (N_1959,N_968,N_1193);
or U1960 (N_1960,N_1024,N_1258);
or U1961 (N_1961,N_1180,N_1444);
or U1962 (N_1962,N_1098,N_1040);
and U1963 (N_1963,N_1375,N_1157);
nor U1964 (N_1964,N_1101,N_1082);
and U1965 (N_1965,N_1300,N_1050);
or U1966 (N_1966,N_762,N_858);
nor U1967 (N_1967,N_1212,N_1274);
and U1968 (N_1968,N_973,N_910);
or U1969 (N_1969,N_1199,N_1402);
or U1970 (N_1970,N_812,N_856);
nor U1971 (N_1971,N_913,N_1497);
nand U1972 (N_1972,N_970,N_1368);
nor U1973 (N_1973,N_809,N_893);
or U1974 (N_1974,N_1199,N_846);
and U1975 (N_1975,N_1211,N_869);
nand U1976 (N_1976,N_861,N_1354);
or U1977 (N_1977,N_1468,N_866);
or U1978 (N_1978,N_1014,N_920);
or U1979 (N_1979,N_988,N_1219);
and U1980 (N_1980,N_1115,N_822);
nand U1981 (N_1981,N_838,N_1328);
xnor U1982 (N_1982,N_1443,N_1465);
nand U1983 (N_1983,N_1031,N_1001);
or U1984 (N_1984,N_1010,N_1175);
nand U1985 (N_1985,N_1409,N_758);
nand U1986 (N_1986,N_1255,N_840);
nor U1987 (N_1987,N_1453,N_941);
nor U1988 (N_1988,N_1370,N_971);
nor U1989 (N_1989,N_867,N_866);
or U1990 (N_1990,N_1300,N_1258);
nor U1991 (N_1991,N_755,N_815);
or U1992 (N_1992,N_1442,N_1223);
nand U1993 (N_1993,N_1257,N_1345);
nor U1994 (N_1994,N_1280,N_1309);
or U1995 (N_1995,N_824,N_1056);
nand U1996 (N_1996,N_854,N_755);
xor U1997 (N_1997,N_1378,N_1084);
nor U1998 (N_1998,N_785,N_766);
and U1999 (N_1999,N_753,N_1293);
nand U2000 (N_2000,N_1022,N_1027);
nor U2001 (N_2001,N_1107,N_1185);
nand U2002 (N_2002,N_1087,N_1444);
nor U2003 (N_2003,N_1168,N_774);
and U2004 (N_2004,N_1214,N_1216);
or U2005 (N_2005,N_1418,N_881);
nor U2006 (N_2006,N_1417,N_944);
or U2007 (N_2007,N_1229,N_877);
nor U2008 (N_2008,N_1178,N_1444);
nor U2009 (N_2009,N_1296,N_908);
or U2010 (N_2010,N_1009,N_877);
nand U2011 (N_2011,N_1285,N_985);
and U2012 (N_2012,N_1170,N_791);
nand U2013 (N_2013,N_1377,N_967);
nand U2014 (N_2014,N_1404,N_850);
or U2015 (N_2015,N_811,N_934);
or U2016 (N_2016,N_997,N_1089);
or U2017 (N_2017,N_1470,N_1064);
and U2018 (N_2018,N_904,N_1071);
nand U2019 (N_2019,N_1312,N_947);
nand U2020 (N_2020,N_1095,N_857);
nor U2021 (N_2021,N_1325,N_835);
nor U2022 (N_2022,N_851,N_1397);
and U2023 (N_2023,N_1490,N_1387);
or U2024 (N_2024,N_1225,N_992);
nand U2025 (N_2025,N_915,N_1218);
or U2026 (N_2026,N_1088,N_991);
or U2027 (N_2027,N_918,N_778);
nand U2028 (N_2028,N_1219,N_880);
or U2029 (N_2029,N_1106,N_812);
xor U2030 (N_2030,N_972,N_1473);
and U2031 (N_2031,N_755,N_866);
or U2032 (N_2032,N_1387,N_1364);
or U2033 (N_2033,N_1219,N_1304);
nor U2034 (N_2034,N_1456,N_1372);
nand U2035 (N_2035,N_1099,N_1291);
or U2036 (N_2036,N_1248,N_1392);
nor U2037 (N_2037,N_1408,N_1095);
or U2038 (N_2038,N_857,N_1211);
or U2039 (N_2039,N_1219,N_962);
or U2040 (N_2040,N_1242,N_819);
nor U2041 (N_2041,N_1436,N_1476);
or U2042 (N_2042,N_1251,N_888);
and U2043 (N_2043,N_1240,N_1499);
nand U2044 (N_2044,N_1326,N_925);
nor U2045 (N_2045,N_986,N_1393);
nand U2046 (N_2046,N_957,N_852);
and U2047 (N_2047,N_1160,N_1303);
nor U2048 (N_2048,N_1009,N_788);
nand U2049 (N_2049,N_1476,N_966);
or U2050 (N_2050,N_1188,N_915);
and U2051 (N_2051,N_1191,N_1209);
or U2052 (N_2052,N_835,N_1182);
or U2053 (N_2053,N_1048,N_1401);
or U2054 (N_2054,N_1062,N_756);
and U2055 (N_2055,N_1218,N_932);
nand U2056 (N_2056,N_1054,N_1362);
or U2057 (N_2057,N_1037,N_1469);
or U2058 (N_2058,N_861,N_1286);
and U2059 (N_2059,N_1177,N_1354);
nand U2060 (N_2060,N_1199,N_1389);
or U2061 (N_2061,N_1397,N_978);
and U2062 (N_2062,N_1197,N_841);
and U2063 (N_2063,N_1076,N_1409);
and U2064 (N_2064,N_1069,N_913);
nand U2065 (N_2065,N_1054,N_1099);
or U2066 (N_2066,N_853,N_787);
nand U2067 (N_2067,N_1418,N_1378);
nor U2068 (N_2068,N_934,N_1176);
or U2069 (N_2069,N_1407,N_1393);
nor U2070 (N_2070,N_1384,N_801);
nor U2071 (N_2071,N_1419,N_1116);
nor U2072 (N_2072,N_1267,N_1493);
and U2073 (N_2073,N_1298,N_855);
nand U2074 (N_2074,N_1119,N_1493);
or U2075 (N_2075,N_1231,N_1305);
and U2076 (N_2076,N_1491,N_872);
nor U2077 (N_2077,N_1221,N_1429);
nor U2078 (N_2078,N_814,N_1080);
nand U2079 (N_2079,N_1283,N_1112);
nor U2080 (N_2080,N_1092,N_851);
or U2081 (N_2081,N_813,N_1308);
or U2082 (N_2082,N_911,N_1224);
nor U2083 (N_2083,N_1410,N_1134);
nand U2084 (N_2084,N_1292,N_753);
nand U2085 (N_2085,N_1390,N_1245);
or U2086 (N_2086,N_1351,N_950);
or U2087 (N_2087,N_1322,N_945);
or U2088 (N_2088,N_1486,N_1024);
and U2089 (N_2089,N_1417,N_1492);
and U2090 (N_2090,N_1264,N_1215);
and U2091 (N_2091,N_1422,N_1344);
nor U2092 (N_2092,N_1117,N_1086);
nand U2093 (N_2093,N_993,N_939);
and U2094 (N_2094,N_962,N_1382);
nand U2095 (N_2095,N_958,N_955);
nand U2096 (N_2096,N_1323,N_1005);
or U2097 (N_2097,N_1350,N_786);
or U2098 (N_2098,N_1282,N_1086);
nand U2099 (N_2099,N_1426,N_764);
or U2100 (N_2100,N_1321,N_945);
nor U2101 (N_2101,N_1032,N_1088);
and U2102 (N_2102,N_836,N_864);
nor U2103 (N_2103,N_1318,N_1088);
nand U2104 (N_2104,N_840,N_1224);
nand U2105 (N_2105,N_803,N_1100);
or U2106 (N_2106,N_1271,N_916);
and U2107 (N_2107,N_988,N_1272);
nor U2108 (N_2108,N_1148,N_862);
and U2109 (N_2109,N_1367,N_956);
nor U2110 (N_2110,N_1301,N_1361);
and U2111 (N_2111,N_1283,N_1480);
and U2112 (N_2112,N_785,N_1243);
nor U2113 (N_2113,N_1178,N_1086);
or U2114 (N_2114,N_918,N_1257);
or U2115 (N_2115,N_1049,N_1132);
nor U2116 (N_2116,N_1265,N_1234);
nor U2117 (N_2117,N_1415,N_1148);
nor U2118 (N_2118,N_925,N_1101);
and U2119 (N_2119,N_1208,N_873);
nand U2120 (N_2120,N_796,N_1170);
or U2121 (N_2121,N_1204,N_1402);
or U2122 (N_2122,N_1099,N_1445);
nor U2123 (N_2123,N_1292,N_810);
and U2124 (N_2124,N_1095,N_1262);
nor U2125 (N_2125,N_1015,N_972);
and U2126 (N_2126,N_1312,N_807);
or U2127 (N_2127,N_1127,N_1135);
nor U2128 (N_2128,N_1446,N_781);
nor U2129 (N_2129,N_1098,N_1298);
or U2130 (N_2130,N_1105,N_1158);
and U2131 (N_2131,N_1438,N_1414);
or U2132 (N_2132,N_1262,N_1265);
nand U2133 (N_2133,N_1142,N_909);
and U2134 (N_2134,N_987,N_936);
nand U2135 (N_2135,N_897,N_1464);
or U2136 (N_2136,N_1149,N_1448);
and U2137 (N_2137,N_1475,N_1411);
nor U2138 (N_2138,N_1208,N_1342);
nand U2139 (N_2139,N_1368,N_817);
or U2140 (N_2140,N_1276,N_1490);
nor U2141 (N_2141,N_1148,N_1498);
and U2142 (N_2142,N_851,N_974);
nor U2143 (N_2143,N_1427,N_1205);
nand U2144 (N_2144,N_1214,N_1171);
nand U2145 (N_2145,N_1026,N_1330);
or U2146 (N_2146,N_769,N_839);
nor U2147 (N_2147,N_1309,N_1023);
nand U2148 (N_2148,N_910,N_965);
and U2149 (N_2149,N_976,N_948);
nand U2150 (N_2150,N_761,N_1014);
nor U2151 (N_2151,N_1211,N_1193);
nand U2152 (N_2152,N_1063,N_1306);
and U2153 (N_2153,N_768,N_866);
and U2154 (N_2154,N_1042,N_1278);
nor U2155 (N_2155,N_1008,N_1486);
nand U2156 (N_2156,N_1086,N_1276);
nand U2157 (N_2157,N_1214,N_1481);
nor U2158 (N_2158,N_1496,N_1394);
and U2159 (N_2159,N_775,N_1002);
and U2160 (N_2160,N_1264,N_872);
and U2161 (N_2161,N_1250,N_1368);
and U2162 (N_2162,N_874,N_1258);
nor U2163 (N_2163,N_862,N_1173);
and U2164 (N_2164,N_876,N_1044);
nand U2165 (N_2165,N_1040,N_1124);
and U2166 (N_2166,N_1255,N_1017);
nor U2167 (N_2167,N_1000,N_1021);
or U2168 (N_2168,N_997,N_1432);
and U2169 (N_2169,N_1291,N_909);
or U2170 (N_2170,N_1066,N_900);
or U2171 (N_2171,N_1058,N_1226);
nand U2172 (N_2172,N_1170,N_949);
and U2173 (N_2173,N_1031,N_1202);
and U2174 (N_2174,N_1180,N_788);
nand U2175 (N_2175,N_1421,N_1194);
nand U2176 (N_2176,N_982,N_981);
nand U2177 (N_2177,N_903,N_779);
nor U2178 (N_2178,N_1221,N_1422);
or U2179 (N_2179,N_1116,N_1156);
nor U2180 (N_2180,N_876,N_1388);
nand U2181 (N_2181,N_1199,N_1114);
and U2182 (N_2182,N_1485,N_1436);
nor U2183 (N_2183,N_1435,N_883);
and U2184 (N_2184,N_899,N_1320);
nor U2185 (N_2185,N_1254,N_1279);
nand U2186 (N_2186,N_784,N_911);
nand U2187 (N_2187,N_1458,N_895);
nand U2188 (N_2188,N_1351,N_1284);
nand U2189 (N_2189,N_1451,N_1397);
and U2190 (N_2190,N_1120,N_959);
nor U2191 (N_2191,N_1013,N_1154);
nand U2192 (N_2192,N_1368,N_898);
or U2193 (N_2193,N_1106,N_955);
nor U2194 (N_2194,N_1283,N_1280);
nor U2195 (N_2195,N_1350,N_839);
or U2196 (N_2196,N_1208,N_1428);
nor U2197 (N_2197,N_1339,N_763);
or U2198 (N_2198,N_1313,N_1180);
nand U2199 (N_2199,N_892,N_1343);
or U2200 (N_2200,N_797,N_1463);
or U2201 (N_2201,N_895,N_1033);
or U2202 (N_2202,N_945,N_761);
nor U2203 (N_2203,N_1429,N_1109);
or U2204 (N_2204,N_1375,N_979);
nand U2205 (N_2205,N_1108,N_1445);
nand U2206 (N_2206,N_1219,N_1253);
nor U2207 (N_2207,N_1179,N_1330);
nor U2208 (N_2208,N_858,N_1473);
or U2209 (N_2209,N_1242,N_1209);
and U2210 (N_2210,N_1199,N_860);
nor U2211 (N_2211,N_959,N_802);
and U2212 (N_2212,N_1375,N_1342);
and U2213 (N_2213,N_1133,N_867);
or U2214 (N_2214,N_1336,N_954);
and U2215 (N_2215,N_1090,N_1259);
nor U2216 (N_2216,N_1288,N_1480);
nand U2217 (N_2217,N_1283,N_797);
or U2218 (N_2218,N_1195,N_1068);
and U2219 (N_2219,N_812,N_951);
nand U2220 (N_2220,N_1059,N_912);
nor U2221 (N_2221,N_1040,N_1266);
nor U2222 (N_2222,N_892,N_765);
or U2223 (N_2223,N_1051,N_1208);
and U2224 (N_2224,N_779,N_1398);
nand U2225 (N_2225,N_777,N_1470);
and U2226 (N_2226,N_888,N_828);
nand U2227 (N_2227,N_891,N_1078);
xnor U2228 (N_2228,N_1109,N_1031);
or U2229 (N_2229,N_1356,N_1329);
or U2230 (N_2230,N_1254,N_1397);
and U2231 (N_2231,N_1388,N_1405);
nor U2232 (N_2232,N_1468,N_1297);
and U2233 (N_2233,N_853,N_1203);
and U2234 (N_2234,N_1179,N_1222);
and U2235 (N_2235,N_1335,N_963);
or U2236 (N_2236,N_1383,N_1172);
nor U2237 (N_2237,N_1335,N_1349);
nand U2238 (N_2238,N_1439,N_1193);
nand U2239 (N_2239,N_794,N_996);
and U2240 (N_2240,N_1114,N_1266);
nand U2241 (N_2241,N_957,N_1339);
and U2242 (N_2242,N_759,N_1435);
and U2243 (N_2243,N_1281,N_1107);
nor U2244 (N_2244,N_807,N_1424);
or U2245 (N_2245,N_1178,N_1342);
or U2246 (N_2246,N_1049,N_1322);
or U2247 (N_2247,N_759,N_938);
nand U2248 (N_2248,N_1261,N_1472);
nor U2249 (N_2249,N_1349,N_818);
or U2250 (N_2250,N_1997,N_1562);
and U2251 (N_2251,N_2133,N_1594);
xnor U2252 (N_2252,N_2087,N_2051);
or U2253 (N_2253,N_2234,N_1753);
or U2254 (N_2254,N_1855,N_1954);
or U2255 (N_2255,N_1588,N_2139);
nor U2256 (N_2256,N_1648,N_1731);
nand U2257 (N_2257,N_1536,N_2205);
or U2258 (N_2258,N_1981,N_2023);
and U2259 (N_2259,N_1698,N_1689);
nor U2260 (N_2260,N_1608,N_1852);
and U2261 (N_2261,N_2142,N_1882);
nor U2262 (N_2262,N_2215,N_1835);
nor U2263 (N_2263,N_1825,N_2081);
and U2264 (N_2264,N_2084,N_2210);
and U2265 (N_2265,N_2120,N_1858);
or U2266 (N_2266,N_2020,N_1820);
nor U2267 (N_2267,N_1958,N_1741);
and U2268 (N_2268,N_1650,N_1752);
or U2269 (N_2269,N_1826,N_1661);
nand U2270 (N_2270,N_1716,N_2116);
nand U2271 (N_2271,N_1868,N_1847);
nand U2272 (N_2272,N_2074,N_1514);
and U2273 (N_2273,N_1695,N_2201);
nand U2274 (N_2274,N_1842,N_2102);
nor U2275 (N_2275,N_1757,N_2016);
nand U2276 (N_2276,N_1808,N_2062);
nor U2277 (N_2277,N_2165,N_1590);
nand U2278 (N_2278,N_1509,N_2245);
or U2279 (N_2279,N_1887,N_1705);
nor U2280 (N_2280,N_1974,N_1722);
and U2281 (N_2281,N_1611,N_2071);
or U2282 (N_2282,N_1863,N_2127);
and U2283 (N_2283,N_1680,N_1549);
and U2284 (N_2284,N_2197,N_1920);
nand U2285 (N_2285,N_2046,N_1559);
nor U2286 (N_2286,N_2209,N_2041);
or U2287 (N_2287,N_1723,N_2214);
nand U2288 (N_2288,N_1940,N_1918);
nor U2289 (N_2289,N_1782,N_1658);
or U2290 (N_2290,N_2146,N_1836);
and U2291 (N_2291,N_2222,N_1881);
and U2292 (N_2292,N_1865,N_1980);
nor U2293 (N_2293,N_2105,N_1572);
and U2294 (N_2294,N_1553,N_1596);
nor U2295 (N_2295,N_1631,N_1665);
and U2296 (N_2296,N_2160,N_1970);
and U2297 (N_2297,N_1829,N_1949);
or U2298 (N_2298,N_2176,N_1864);
nor U2299 (N_2299,N_1990,N_1651);
nor U2300 (N_2300,N_2244,N_1925);
nor U2301 (N_2301,N_2104,N_1856);
and U2302 (N_2302,N_1643,N_1555);
and U2303 (N_2303,N_1520,N_2153);
nand U2304 (N_2304,N_2191,N_2013);
nand U2305 (N_2305,N_1804,N_1908);
nor U2306 (N_2306,N_1971,N_1500);
and U2307 (N_2307,N_2189,N_1806);
or U2308 (N_2308,N_2048,N_1937);
nor U2309 (N_2309,N_1807,N_1953);
and U2310 (N_2310,N_1917,N_1668);
or U2311 (N_2311,N_1535,N_1973);
nor U2312 (N_2312,N_1686,N_1542);
nand U2313 (N_2313,N_2075,N_1923);
nand U2314 (N_2314,N_2027,N_2098);
and U2315 (N_2315,N_1606,N_1713);
nor U2316 (N_2316,N_1816,N_2158);
nor U2317 (N_2317,N_2175,N_2125);
nand U2318 (N_2318,N_2179,N_1595);
or U2319 (N_2319,N_1541,N_1916);
nor U2320 (N_2320,N_2178,N_2243);
or U2321 (N_2321,N_1607,N_1899);
nor U2322 (N_2322,N_2093,N_1831);
nand U2323 (N_2323,N_1646,N_1724);
or U2324 (N_2324,N_1503,N_2052);
or U2325 (N_2325,N_1991,N_1884);
nor U2326 (N_2326,N_1837,N_2216);
nor U2327 (N_2327,N_2157,N_1736);
nor U2328 (N_2328,N_1708,N_2237);
and U2329 (N_2329,N_2114,N_1687);
or U2330 (N_2330,N_2221,N_1720);
nor U2331 (N_2331,N_2026,N_1960);
nand U2332 (N_2332,N_1756,N_2100);
nor U2333 (N_2333,N_2110,N_1690);
or U2334 (N_2334,N_1662,N_1507);
xor U2335 (N_2335,N_1580,N_2091);
nand U2336 (N_2336,N_2092,N_1879);
nand U2337 (N_2337,N_2140,N_2060);
or U2338 (N_2338,N_2031,N_1929);
and U2339 (N_2339,N_1567,N_1630);
and U2340 (N_2340,N_2180,N_1853);
and U2341 (N_2341,N_1578,N_2218);
nor U2342 (N_2342,N_1944,N_1934);
nand U2343 (N_2343,N_2049,N_2053);
nor U2344 (N_2344,N_1823,N_2144);
or U2345 (N_2345,N_1563,N_2067);
or U2346 (N_2346,N_1739,N_2128);
or U2347 (N_2347,N_1778,N_2111);
nand U2348 (N_2348,N_1926,N_2231);
nand U2349 (N_2349,N_1721,N_1706);
nor U2350 (N_2350,N_1692,N_1815);
nand U2351 (N_2351,N_1604,N_1565);
nor U2352 (N_2352,N_1955,N_2090);
nor U2353 (N_2353,N_1583,N_1560);
or U2354 (N_2354,N_2055,N_2159);
and U2355 (N_2355,N_1784,N_1964);
and U2356 (N_2356,N_2012,N_2112);
nor U2357 (N_2357,N_1667,N_1691);
nor U2358 (N_2358,N_2036,N_1638);
and U2359 (N_2359,N_1593,N_1652);
nor U2360 (N_2360,N_1781,N_1709);
nor U2361 (N_2361,N_1699,N_2192);
and U2362 (N_2362,N_1543,N_1527);
or U2363 (N_2363,N_1532,N_1821);
nor U2364 (N_2364,N_1874,N_1615);
nand U2365 (N_2365,N_1810,N_1552);
nor U2366 (N_2366,N_1905,N_1927);
nand U2367 (N_2367,N_1576,N_1670);
or U2368 (N_2368,N_2109,N_2138);
or U2369 (N_2369,N_1663,N_1601);
nor U2370 (N_2370,N_1620,N_1566);
xor U2371 (N_2371,N_1712,N_1632);
and U2372 (N_2372,N_1759,N_1888);
nor U2373 (N_2373,N_1965,N_1840);
nand U2374 (N_2374,N_1586,N_2001);
and U2375 (N_2375,N_1894,N_2045);
or U2376 (N_2376,N_1945,N_2149);
or U2377 (N_2377,N_1575,N_2249);
and U2378 (N_2378,N_1569,N_1525);
nand U2379 (N_2379,N_2220,N_1733);
nor U2380 (N_2380,N_2141,N_1700);
nand U2381 (N_2381,N_1946,N_2219);
and U2382 (N_2382,N_1857,N_2009);
nand U2383 (N_2383,N_2029,N_2204);
and U2384 (N_2384,N_1963,N_2212);
nor U2385 (N_2385,N_2008,N_2166);
and U2386 (N_2386,N_2014,N_1775);
nor U2387 (N_2387,N_1785,N_1762);
and U2388 (N_2388,N_2145,N_2011);
nand U2389 (N_2389,N_1561,N_1589);
nand U2390 (N_2390,N_2163,N_2118);
or U2391 (N_2391,N_2068,N_1996);
or U2392 (N_2392,N_2078,N_1719);
nor U2393 (N_2393,N_1798,N_2208);
nor U2394 (N_2394,N_2037,N_2129);
or U2395 (N_2395,N_1635,N_1780);
xor U2396 (N_2396,N_1906,N_2030);
nor U2397 (N_2397,N_1904,N_1893);
and U2398 (N_2398,N_1627,N_1701);
nand U2399 (N_2399,N_1773,N_2168);
and U2400 (N_2400,N_1763,N_1967);
or U2401 (N_2401,N_2228,N_1506);
and U2402 (N_2402,N_1793,N_1743);
nand U2403 (N_2403,N_2079,N_1637);
nor U2404 (N_2404,N_1938,N_1833);
or U2405 (N_2405,N_2123,N_2136);
and U2406 (N_2406,N_2150,N_1523);
nand U2407 (N_2407,N_1735,N_1614);
nand U2408 (N_2408,N_1745,N_1693);
and U2409 (N_2409,N_1896,N_2240);
and U2410 (N_2410,N_1948,N_1554);
or U2411 (N_2411,N_1598,N_1516);
or U2412 (N_2412,N_1790,N_1626);
or U2413 (N_2413,N_1921,N_1851);
nor U2414 (N_2414,N_2061,N_2181);
nand U2415 (N_2415,N_1966,N_1765);
nor U2416 (N_2416,N_1750,N_1504);
and U2417 (N_2417,N_2038,N_1729);
or U2418 (N_2418,N_1633,N_1911);
nor U2419 (N_2419,N_2238,N_1546);
or U2420 (N_2420,N_1848,N_1922);
nand U2421 (N_2421,N_1886,N_1818);
or U2422 (N_2422,N_1803,N_1792);
nand U2423 (N_2423,N_1738,N_1714);
and U2424 (N_2424,N_1629,N_1915);
or U2425 (N_2425,N_1975,N_1682);
or U2426 (N_2426,N_1641,N_1900);
nor U2427 (N_2427,N_1732,N_2230);
and U2428 (N_2428,N_1664,N_1794);
nand U2429 (N_2429,N_1557,N_2135);
nor U2430 (N_2430,N_1844,N_2021);
nand U2431 (N_2431,N_1850,N_2151);
and U2432 (N_2432,N_1571,N_1909);
and U2433 (N_2433,N_1933,N_2132);
nand U2434 (N_2434,N_1564,N_1924);
nand U2435 (N_2435,N_1612,N_1801);
and U2436 (N_2436,N_2226,N_1534);
nor U2437 (N_2437,N_1969,N_1984);
or U2438 (N_2438,N_2198,N_2007);
nor U2439 (N_2439,N_1769,N_1528);
and U2440 (N_2440,N_1617,N_1849);
or U2441 (N_2441,N_1702,N_2088);
or U2442 (N_2442,N_2034,N_2134);
nor U2443 (N_2443,N_2119,N_2115);
or U2444 (N_2444,N_1895,N_1995);
nand U2445 (N_2445,N_2184,N_1545);
or U2446 (N_2446,N_1602,N_1809);
nor U2447 (N_2447,N_1889,N_1843);
nand U2448 (N_2448,N_2217,N_2235);
nand U2449 (N_2449,N_2099,N_2019);
and U2450 (N_2450,N_2069,N_2035);
nor U2451 (N_2451,N_1581,N_2170);
and U2452 (N_2452,N_1530,N_2039);
xor U2453 (N_2453,N_1869,N_1547);
nor U2454 (N_2454,N_1987,N_1715);
nand U2455 (N_2455,N_1846,N_2182);
and U2456 (N_2456,N_1574,N_2033);
nand U2457 (N_2457,N_1622,N_1685);
or U2458 (N_2458,N_1795,N_1951);
nand U2459 (N_2459,N_1678,N_2130);
nor U2460 (N_2460,N_1616,N_1704);
nand U2461 (N_2461,N_1587,N_1548);
or U2462 (N_2462,N_1737,N_2089);
nor U2463 (N_2463,N_1619,N_1813);
or U2464 (N_2464,N_1977,N_1524);
xnor U2465 (N_2465,N_2147,N_2076);
and U2466 (N_2466,N_2117,N_2101);
and U2467 (N_2467,N_1600,N_2174);
and U2468 (N_2468,N_2095,N_2167);
or U2469 (N_2469,N_1505,N_2143);
and U2470 (N_2470,N_2017,N_1799);
xnor U2471 (N_2471,N_1861,N_1989);
nand U2472 (N_2472,N_1754,N_2002);
nor U2473 (N_2473,N_1533,N_1928);
or U2474 (N_2474,N_1515,N_2018);
nor U2475 (N_2475,N_1772,N_1728);
or U2476 (N_2476,N_2070,N_1718);
and U2477 (N_2477,N_2108,N_1625);
or U2478 (N_2478,N_1746,N_1779);
or U2479 (N_2479,N_1994,N_1513);
nand U2480 (N_2480,N_1654,N_1866);
nor U2481 (N_2481,N_1675,N_2248);
nand U2482 (N_2482,N_2207,N_1788);
nand U2483 (N_2483,N_1556,N_1812);
nand U2484 (N_2484,N_1783,N_1898);
nand U2485 (N_2485,N_1609,N_1679);
and U2486 (N_2486,N_1824,N_1684);
and U2487 (N_2487,N_1657,N_1982);
and U2488 (N_2488,N_1747,N_1791);
nand U2489 (N_2489,N_2073,N_1742);
nor U2490 (N_2490,N_1901,N_1942);
or U2491 (N_2491,N_1907,N_1755);
nand U2492 (N_2492,N_2225,N_1777);
and U2493 (N_2493,N_1544,N_2096);
or U2494 (N_2494,N_1734,N_1903);
or U2495 (N_2495,N_2000,N_1919);
or U2496 (N_2496,N_1789,N_1870);
and U2497 (N_2497,N_1621,N_2004);
nand U2498 (N_2498,N_2113,N_1988);
nor U2499 (N_2499,N_1860,N_2195);
nor U2500 (N_2500,N_2164,N_1592);
nand U2501 (N_2501,N_2187,N_2241);
nor U2502 (N_2502,N_1885,N_2094);
xor U2503 (N_2503,N_1673,N_1914);
or U2504 (N_2504,N_1683,N_2010);
or U2505 (N_2505,N_1797,N_1510);
and U2506 (N_2506,N_1710,N_1947);
nand U2507 (N_2507,N_2015,N_1717);
nor U2508 (N_2508,N_2177,N_2124);
and U2509 (N_2509,N_1822,N_1838);
and U2510 (N_2510,N_1599,N_1744);
and U2511 (N_2511,N_1986,N_1760);
and U2512 (N_2512,N_2203,N_1992);
and U2513 (N_2513,N_2155,N_1636);
nor U2514 (N_2514,N_1669,N_1819);
and U2515 (N_2515,N_1913,N_1579);
nor U2516 (N_2516,N_2211,N_2044);
nand U2517 (N_2517,N_2050,N_1644);
nor U2518 (N_2518,N_1501,N_2224);
nand U2519 (N_2519,N_1883,N_1688);
or U2520 (N_2520,N_1800,N_1660);
nor U2521 (N_2521,N_1591,N_2233);
or U2522 (N_2522,N_1539,N_2003);
xor U2523 (N_2523,N_1956,N_2196);
and U2524 (N_2524,N_2242,N_2040);
and U2525 (N_2525,N_2152,N_1962);
nand U2526 (N_2526,N_2156,N_1570);
nand U2527 (N_2527,N_1845,N_1985);
and U2528 (N_2528,N_2172,N_1897);
nand U2529 (N_2529,N_1758,N_1518);
nor U2530 (N_2530,N_1711,N_1568);
nor U2531 (N_2531,N_1841,N_2103);
nor U2532 (N_2532,N_1979,N_2199);
nor U2533 (N_2533,N_1610,N_1936);
nor U2534 (N_2534,N_1707,N_2131);
and U2535 (N_2535,N_1828,N_2006);
and U2536 (N_2536,N_1943,N_1511);
nand U2537 (N_2537,N_2185,N_1508);
or U2538 (N_2538,N_1584,N_1978);
and U2539 (N_2539,N_2107,N_2042);
nor U2540 (N_2540,N_1659,N_1976);
and U2541 (N_2541,N_1618,N_2057);
nand U2542 (N_2542,N_1912,N_2054);
nand U2543 (N_2543,N_2229,N_1878);
and U2544 (N_2544,N_1655,N_1537);
nor U2545 (N_2545,N_1827,N_1639);
nor U2546 (N_2546,N_2126,N_1697);
nor U2547 (N_2547,N_1726,N_1573);
or U2548 (N_2548,N_2077,N_1939);
nor U2549 (N_2549,N_1730,N_1681);
nand U2550 (N_2550,N_1993,N_1748);
nand U2551 (N_2551,N_1634,N_1802);
nand U2552 (N_2552,N_1672,N_1876);
or U2553 (N_2553,N_2169,N_1774);
nor U2554 (N_2554,N_1613,N_1931);
xnor U2555 (N_2555,N_1968,N_1649);
nand U2556 (N_2556,N_1832,N_2085);
nor U2557 (N_2557,N_1666,N_1623);
nor U2558 (N_2558,N_1749,N_2148);
and U2559 (N_2559,N_2188,N_2183);
nand U2560 (N_2560,N_2239,N_1959);
nor U2561 (N_2561,N_2080,N_1877);
and U2562 (N_2562,N_2223,N_1817);
or U2563 (N_2563,N_2247,N_1740);
or U2564 (N_2564,N_1767,N_2005);
and U2565 (N_2565,N_1932,N_2121);
or U2566 (N_2566,N_1577,N_1558);
nor U2567 (N_2567,N_2137,N_1902);
and U2568 (N_2568,N_1854,N_1952);
and U2569 (N_2569,N_1764,N_2200);
and U2570 (N_2570,N_1770,N_1941);
or U2571 (N_2571,N_1696,N_1538);
nand U2572 (N_2572,N_1642,N_1502);
nor U2573 (N_2573,N_2072,N_2206);
nor U2574 (N_2574,N_2236,N_1891);
nand U2575 (N_2575,N_1582,N_1890);
and U2576 (N_2576,N_2173,N_1796);
and U2577 (N_2577,N_1873,N_1998);
nor U2578 (N_2578,N_2232,N_1859);
and U2579 (N_2579,N_2025,N_1972);
or U2580 (N_2580,N_2097,N_1526);
and U2581 (N_2581,N_1540,N_1653);
nor U2582 (N_2582,N_2047,N_1771);
and U2583 (N_2583,N_1531,N_1871);
nor U2584 (N_2584,N_1550,N_2032);
or U2585 (N_2585,N_2194,N_1597);
nand U2586 (N_2586,N_1880,N_1603);
and U2587 (N_2587,N_1787,N_2213);
and U2588 (N_2588,N_2043,N_2190);
and U2589 (N_2589,N_2056,N_2024);
nor U2590 (N_2590,N_1892,N_1839);
and U2591 (N_2591,N_1999,N_2063);
and U2592 (N_2592,N_2066,N_1811);
xor U2593 (N_2593,N_2246,N_1814);
nor U2594 (N_2594,N_1766,N_1830);
nand U2595 (N_2595,N_1862,N_1910);
and U2596 (N_2596,N_2227,N_2082);
xor U2597 (N_2597,N_1935,N_2122);
nor U2598 (N_2598,N_1647,N_1930);
or U2599 (N_2599,N_1551,N_1694);
and U2600 (N_2600,N_1522,N_2064);
and U2601 (N_2601,N_2202,N_1776);
nand U2602 (N_2602,N_2154,N_1677);
nor U2603 (N_2603,N_2059,N_2086);
nand U2604 (N_2604,N_1983,N_1867);
and U2605 (N_2605,N_1768,N_1628);
or U2606 (N_2606,N_1751,N_1961);
or U2607 (N_2607,N_1725,N_2083);
nor U2608 (N_2608,N_1957,N_1585);
nand U2609 (N_2609,N_1761,N_1950);
nor U2610 (N_2610,N_2058,N_2028);
and U2611 (N_2611,N_1727,N_1834);
and U2612 (N_2612,N_1521,N_2193);
or U2613 (N_2613,N_1529,N_2022);
or U2614 (N_2614,N_1703,N_1656);
nand U2615 (N_2615,N_1605,N_2171);
or U2616 (N_2616,N_1872,N_2106);
nor U2617 (N_2617,N_1786,N_1676);
or U2618 (N_2618,N_1624,N_2161);
or U2619 (N_2619,N_1875,N_1674);
nor U2620 (N_2620,N_1512,N_1519);
nor U2621 (N_2621,N_1671,N_2186);
nand U2622 (N_2622,N_1645,N_1640);
or U2623 (N_2623,N_2065,N_2162);
or U2624 (N_2624,N_1805,N_1517);
or U2625 (N_2625,N_2072,N_2099);
and U2626 (N_2626,N_1599,N_1669);
or U2627 (N_2627,N_1628,N_1778);
or U2628 (N_2628,N_1939,N_1767);
nand U2629 (N_2629,N_2164,N_2038);
nor U2630 (N_2630,N_1748,N_1502);
nor U2631 (N_2631,N_2062,N_1938);
and U2632 (N_2632,N_1655,N_2183);
or U2633 (N_2633,N_1998,N_1749);
nor U2634 (N_2634,N_2118,N_1553);
or U2635 (N_2635,N_2107,N_1778);
nor U2636 (N_2636,N_2108,N_1681);
and U2637 (N_2637,N_1793,N_1772);
nand U2638 (N_2638,N_1761,N_1943);
or U2639 (N_2639,N_1561,N_2172);
nand U2640 (N_2640,N_2075,N_1732);
nor U2641 (N_2641,N_1536,N_1604);
and U2642 (N_2642,N_1643,N_2080);
nor U2643 (N_2643,N_1832,N_1974);
nor U2644 (N_2644,N_1679,N_1509);
nor U2645 (N_2645,N_2036,N_1814);
or U2646 (N_2646,N_1907,N_1703);
or U2647 (N_2647,N_2243,N_1776);
and U2648 (N_2648,N_1780,N_2130);
or U2649 (N_2649,N_1616,N_1706);
nand U2650 (N_2650,N_1559,N_1873);
nand U2651 (N_2651,N_1755,N_2051);
or U2652 (N_2652,N_2208,N_1579);
or U2653 (N_2653,N_1633,N_2163);
and U2654 (N_2654,N_1933,N_2146);
nand U2655 (N_2655,N_1996,N_1536);
and U2656 (N_2656,N_1868,N_1716);
or U2657 (N_2657,N_1922,N_2134);
or U2658 (N_2658,N_1572,N_1776);
nor U2659 (N_2659,N_2127,N_1994);
nor U2660 (N_2660,N_2060,N_1981);
nand U2661 (N_2661,N_2053,N_1563);
or U2662 (N_2662,N_1785,N_1714);
and U2663 (N_2663,N_2048,N_2185);
nor U2664 (N_2664,N_2036,N_2110);
or U2665 (N_2665,N_1667,N_2113);
nor U2666 (N_2666,N_1580,N_1778);
and U2667 (N_2667,N_1833,N_1804);
and U2668 (N_2668,N_1964,N_1645);
and U2669 (N_2669,N_1636,N_1705);
or U2670 (N_2670,N_2242,N_1871);
nor U2671 (N_2671,N_1872,N_1685);
nor U2672 (N_2672,N_1645,N_1949);
or U2673 (N_2673,N_1799,N_1507);
nor U2674 (N_2674,N_2157,N_1976);
nor U2675 (N_2675,N_1992,N_1825);
and U2676 (N_2676,N_1716,N_1534);
xnor U2677 (N_2677,N_1962,N_1622);
nor U2678 (N_2678,N_1925,N_1734);
nor U2679 (N_2679,N_2085,N_2199);
or U2680 (N_2680,N_1716,N_1517);
or U2681 (N_2681,N_2103,N_1607);
and U2682 (N_2682,N_1651,N_2217);
or U2683 (N_2683,N_1759,N_1990);
nor U2684 (N_2684,N_2050,N_2216);
nand U2685 (N_2685,N_1589,N_2221);
nor U2686 (N_2686,N_1504,N_2183);
or U2687 (N_2687,N_2087,N_2115);
or U2688 (N_2688,N_1898,N_1558);
nor U2689 (N_2689,N_2079,N_1820);
nand U2690 (N_2690,N_1750,N_1894);
and U2691 (N_2691,N_2127,N_2124);
nand U2692 (N_2692,N_1503,N_2081);
nor U2693 (N_2693,N_1652,N_1901);
nor U2694 (N_2694,N_1854,N_1772);
or U2695 (N_2695,N_2033,N_1729);
nor U2696 (N_2696,N_1966,N_1580);
or U2697 (N_2697,N_1830,N_2094);
nand U2698 (N_2698,N_1853,N_2205);
or U2699 (N_2699,N_2030,N_2244);
or U2700 (N_2700,N_1942,N_1842);
or U2701 (N_2701,N_1861,N_1628);
xnor U2702 (N_2702,N_2145,N_2031);
or U2703 (N_2703,N_2116,N_2217);
nor U2704 (N_2704,N_1554,N_1936);
or U2705 (N_2705,N_2156,N_1583);
or U2706 (N_2706,N_1921,N_1606);
xnor U2707 (N_2707,N_2095,N_1611);
and U2708 (N_2708,N_1565,N_2070);
nor U2709 (N_2709,N_1956,N_1802);
and U2710 (N_2710,N_1541,N_2192);
or U2711 (N_2711,N_2164,N_1933);
nand U2712 (N_2712,N_1899,N_1671);
and U2713 (N_2713,N_1574,N_1882);
nor U2714 (N_2714,N_1812,N_1863);
and U2715 (N_2715,N_1911,N_1512);
or U2716 (N_2716,N_1554,N_1548);
and U2717 (N_2717,N_2192,N_2159);
nor U2718 (N_2718,N_1889,N_1729);
nand U2719 (N_2719,N_2049,N_1893);
nand U2720 (N_2720,N_1504,N_1591);
and U2721 (N_2721,N_1522,N_1786);
nand U2722 (N_2722,N_2174,N_1777);
nor U2723 (N_2723,N_2109,N_1738);
or U2724 (N_2724,N_2187,N_2016);
nor U2725 (N_2725,N_1818,N_1863);
nand U2726 (N_2726,N_1614,N_1693);
or U2727 (N_2727,N_1783,N_1743);
and U2728 (N_2728,N_2132,N_1614);
nor U2729 (N_2729,N_2173,N_1802);
nand U2730 (N_2730,N_1896,N_2121);
nor U2731 (N_2731,N_1727,N_1736);
or U2732 (N_2732,N_2113,N_1607);
and U2733 (N_2733,N_1956,N_2008);
and U2734 (N_2734,N_1741,N_2219);
nor U2735 (N_2735,N_1668,N_2043);
nor U2736 (N_2736,N_1765,N_1885);
and U2737 (N_2737,N_2175,N_1502);
nand U2738 (N_2738,N_2025,N_1570);
or U2739 (N_2739,N_1577,N_1590);
or U2740 (N_2740,N_1966,N_1973);
nor U2741 (N_2741,N_2128,N_1785);
nand U2742 (N_2742,N_2139,N_2010);
nand U2743 (N_2743,N_1804,N_2233);
nand U2744 (N_2744,N_2226,N_1747);
and U2745 (N_2745,N_2163,N_1630);
xnor U2746 (N_2746,N_1629,N_1979);
nor U2747 (N_2747,N_1760,N_2231);
or U2748 (N_2748,N_1997,N_2239);
nand U2749 (N_2749,N_2070,N_1714);
nand U2750 (N_2750,N_1989,N_2222);
and U2751 (N_2751,N_2020,N_1537);
nor U2752 (N_2752,N_2085,N_1600);
and U2753 (N_2753,N_1822,N_2105);
or U2754 (N_2754,N_1939,N_1640);
and U2755 (N_2755,N_1897,N_1666);
or U2756 (N_2756,N_1913,N_2175);
or U2757 (N_2757,N_1659,N_1536);
or U2758 (N_2758,N_1999,N_1824);
and U2759 (N_2759,N_2041,N_2206);
nand U2760 (N_2760,N_1963,N_1505);
or U2761 (N_2761,N_1548,N_2088);
and U2762 (N_2762,N_1735,N_1715);
nand U2763 (N_2763,N_1989,N_1799);
nand U2764 (N_2764,N_2173,N_1933);
and U2765 (N_2765,N_1928,N_1558);
or U2766 (N_2766,N_1505,N_1732);
nor U2767 (N_2767,N_1714,N_1922);
or U2768 (N_2768,N_2186,N_2039);
or U2769 (N_2769,N_2077,N_2006);
or U2770 (N_2770,N_1577,N_2079);
and U2771 (N_2771,N_1800,N_1725);
and U2772 (N_2772,N_1793,N_1770);
nand U2773 (N_2773,N_1980,N_1905);
nor U2774 (N_2774,N_1822,N_1911);
and U2775 (N_2775,N_1691,N_1671);
nand U2776 (N_2776,N_1791,N_2110);
nor U2777 (N_2777,N_2158,N_1905);
and U2778 (N_2778,N_2024,N_1673);
or U2779 (N_2779,N_2158,N_1985);
or U2780 (N_2780,N_1605,N_2201);
nand U2781 (N_2781,N_1666,N_1503);
and U2782 (N_2782,N_1622,N_2194);
and U2783 (N_2783,N_1992,N_1549);
nor U2784 (N_2784,N_2216,N_1614);
and U2785 (N_2785,N_1872,N_2145);
nand U2786 (N_2786,N_1965,N_1500);
nor U2787 (N_2787,N_2162,N_2050);
nor U2788 (N_2788,N_1651,N_1979);
or U2789 (N_2789,N_1890,N_2134);
or U2790 (N_2790,N_1700,N_1630);
nor U2791 (N_2791,N_1778,N_1904);
or U2792 (N_2792,N_1600,N_1582);
nand U2793 (N_2793,N_1527,N_2043);
and U2794 (N_2794,N_1563,N_1659);
nand U2795 (N_2795,N_1945,N_1810);
and U2796 (N_2796,N_1563,N_2023);
and U2797 (N_2797,N_2160,N_1672);
nor U2798 (N_2798,N_2056,N_2249);
nand U2799 (N_2799,N_2097,N_2110);
and U2800 (N_2800,N_1525,N_1703);
or U2801 (N_2801,N_1823,N_1894);
and U2802 (N_2802,N_2033,N_1819);
nor U2803 (N_2803,N_1542,N_1587);
or U2804 (N_2804,N_1820,N_1704);
nand U2805 (N_2805,N_2090,N_1829);
and U2806 (N_2806,N_1951,N_1979);
nand U2807 (N_2807,N_1893,N_1580);
or U2808 (N_2808,N_2218,N_1706);
or U2809 (N_2809,N_1564,N_1810);
nor U2810 (N_2810,N_1729,N_1994);
or U2811 (N_2811,N_2057,N_1827);
nor U2812 (N_2812,N_1581,N_1684);
or U2813 (N_2813,N_1585,N_2128);
nor U2814 (N_2814,N_2148,N_2165);
nor U2815 (N_2815,N_1507,N_2121);
xnor U2816 (N_2816,N_2092,N_2017);
nor U2817 (N_2817,N_1687,N_1876);
and U2818 (N_2818,N_1867,N_2041);
or U2819 (N_2819,N_2207,N_1934);
xor U2820 (N_2820,N_2077,N_1927);
nand U2821 (N_2821,N_1894,N_1951);
or U2822 (N_2822,N_1572,N_1946);
and U2823 (N_2823,N_1950,N_1654);
and U2824 (N_2824,N_1575,N_2061);
nor U2825 (N_2825,N_1814,N_1805);
and U2826 (N_2826,N_1606,N_2136);
and U2827 (N_2827,N_1913,N_2148);
nand U2828 (N_2828,N_1509,N_1765);
and U2829 (N_2829,N_2087,N_1530);
or U2830 (N_2830,N_1735,N_1742);
nor U2831 (N_2831,N_2108,N_2187);
nor U2832 (N_2832,N_1591,N_1681);
nor U2833 (N_2833,N_2204,N_1537);
and U2834 (N_2834,N_1699,N_1626);
nor U2835 (N_2835,N_1990,N_1596);
or U2836 (N_2836,N_1639,N_2089);
xor U2837 (N_2837,N_2170,N_2211);
and U2838 (N_2838,N_1565,N_1672);
or U2839 (N_2839,N_1923,N_2170);
nor U2840 (N_2840,N_1859,N_1810);
or U2841 (N_2841,N_1981,N_1615);
or U2842 (N_2842,N_2119,N_1745);
nand U2843 (N_2843,N_1810,N_1762);
nand U2844 (N_2844,N_1622,N_1908);
xor U2845 (N_2845,N_1575,N_2073);
and U2846 (N_2846,N_1992,N_1836);
and U2847 (N_2847,N_1817,N_2189);
and U2848 (N_2848,N_1990,N_1692);
nor U2849 (N_2849,N_1717,N_2239);
or U2850 (N_2850,N_1881,N_2225);
or U2851 (N_2851,N_1521,N_1563);
or U2852 (N_2852,N_1583,N_1636);
and U2853 (N_2853,N_1685,N_1673);
or U2854 (N_2854,N_2241,N_1677);
nor U2855 (N_2855,N_1537,N_2181);
xnor U2856 (N_2856,N_1626,N_1919);
and U2857 (N_2857,N_1509,N_1875);
and U2858 (N_2858,N_1924,N_1556);
or U2859 (N_2859,N_1564,N_2215);
or U2860 (N_2860,N_1712,N_2183);
nand U2861 (N_2861,N_2146,N_2022);
nor U2862 (N_2862,N_1830,N_1502);
nor U2863 (N_2863,N_1540,N_1749);
and U2864 (N_2864,N_2068,N_1862);
nor U2865 (N_2865,N_1941,N_1994);
and U2866 (N_2866,N_1658,N_1566);
xor U2867 (N_2867,N_1680,N_1684);
nand U2868 (N_2868,N_2177,N_1644);
and U2869 (N_2869,N_1577,N_1579);
nor U2870 (N_2870,N_1708,N_1854);
or U2871 (N_2871,N_1981,N_2102);
or U2872 (N_2872,N_1582,N_1807);
nand U2873 (N_2873,N_1599,N_2025);
or U2874 (N_2874,N_1665,N_2023);
or U2875 (N_2875,N_1647,N_1576);
or U2876 (N_2876,N_1544,N_1857);
and U2877 (N_2877,N_1863,N_1959);
nand U2878 (N_2878,N_1946,N_2090);
nand U2879 (N_2879,N_1983,N_1974);
and U2880 (N_2880,N_1544,N_2245);
nor U2881 (N_2881,N_1941,N_1922);
and U2882 (N_2882,N_1702,N_1912);
nor U2883 (N_2883,N_1881,N_1627);
or U2884 (N_2884,N_2208,N_2065);
and U2885 (N_2885,N_1536,N_1668);
nand U2886 (N_2886,N_1644,N_2090);
nor U2887 (N_2887,N_1667,N_1663);
or U2888 (N_2888,N_2097,N_2245);
nand U2889 (N_2889,N_1922,N_1726);
or U2890 (N_2890,N_2063,N_1839);
and U2891 (N_2891,N_1566,N_1806);
nand U2892 (N_2892,N_1710,N_1743);
nand U2893 (N_2893,N_1694,N_2158);
or U2894 (N_2894,N_2163,N_2150);
or U2895 (N_2895,N_1631,N_1678);
or U2896 (N_2896,N_1643,N_1554);
nand U2897 (N_2897,N_2082,N_1544);
nor U2898 (N_2898,N_2002,N_2089);
nand U2899 (N_2899,N_2163,N_1732);
nand U2900 (N_2900,N_1898,N_2248);
or U2901 (N_2901,N_2004,N_1765);
and U2902 (N_2902,N_1856,N_1849);
nor U2903 (N_2903,N_1603,N_2048);
nand U2904 (N_2904,N_1952,N_2192);
or U2905 (N_2905,N_1617,N_1640);
or U2906 (N_2906,N_1833,N_1882);
nand U2907 (N_2907,N_1707,N_1693);
nand U2908 (N_2908,N_2194,N_2173);
and U2909 (N_2909,N_1781,N_2098);
nor U2910 (N_2910,N_1904,N_1586);
nand U2911 (N_2911,N_1976,N_1663);
nor U2912 (N_2912,N_1892,N_2129);
and U2913 (N_2913,N_1596,N_1986);
nor U2914 (N_2914,N_1841,N_1784);
nand U2915 (N_2915,N_1637,N_1925);
nor U2916 (N_2916,N_1594,N_2109);
or U2917 (N_2917,N_1627,N_1831);
or U2918 (N_2918,N_1723,N_1937);
nor U2919 (N_2919,N_1766,N_1730);
and U2920 (N_2920,N_2177,N_1551);
and U2921 (N_2921,N_1581,N_2184);
and U2922 (N_2922,N_2132,N_1998);
or U2923 (N_2923,N_2181,N_1940);
or U2924 (N_2924,N_1799,N_1653);
nor U2925 (N_2925,N_2172,N_2070);
and U2926 (N_2926,N_2042,N_1682);
nor U2927 (N_2927,N_1607,N_2085);
nor U2928 (N_2928,N_1563,N_1793);
nand U2929 (N_2929,N_2215,N_1659);
nand U2930 (N_2930,N_2230,N_1915);
nand U2931 (N_2931,N_2058,N_1639);
and U2932 (N_2932,N_1828,N_1870);
or U2933 (N_2933,N_1542,N_1920);
and U2934 (N_2934,N_2148,N_1639);
nor U2935 (N_2935,N_2106,N_1650);
or U2936 (N_2936,N_1981,N_2169);
nor U2937 (N_2937,N_1741,N_1795);
nand U2938 (N_2938,N_1884,N_1759);
nor U2939 (N_2939,N_1912,N_1731);
nand U2940 (N_2940,N_2099,N_1572);
nor U2941 (N_2941,N_1767,N_2079);
or U2942 (N_2942,N_1850,N_1716);
and U2943 (N_2943,N_2116,N_1600);
or U2944 (N_2944,N_2055,N_1958);
nand U2945 (N_2945,N_1576,N_1901);
nor U2946 (N_2946,N_1549,N_2188);
or U2947 (N_2947,N_1621,N_2126);
or U2948 (N_2948,N_1821,N_1573);
nand U2949 (N_2949,N_1696,N_1726);
or U2950 (N_2950,N_1548,N_1507);
nand U2951 (N_2951,N_1591,N_1952);
or U2952 (N_2952,N_1542,N_1855);
nor U2953 (N_2953,N_1510,N_1532);
or U2954 (N_2954,N_1528,N_1545);
xnor U2955 (N_2955,N_1637,N_1669);
nand U2956 (N_2956,N_1555,N_2220);
or U2957 (N_2957,N_2156,N_1926);
nand U2958 (N_2958,N_2036,N_2229);
or U2959 (N_2959,N_1908,N_2208);
or U2960 (N_2960,N_1853,N_1973);
or U2961 (N_2961,N_1822,N_1652);
and U2962 (N_2962,N_2146,N_1695);
or U2963 (N_2963,N_2091,N_1564);
nor U2964 (N_2964,N_1990,N_2141);
xor U2965 (N_2965,N_1842,N_1763);
nand U2966 (N_2966,N_1835,N_1847);
nor U2967 (N_2967,N_2139,N_1778);
nand U2968 (N_2968,N_1989,N_2078);
or U2969 (N_2969,N_2056,N_1524);
nor U2970 (N_2970,N_1807,N_2098);
nand U2971 (N_2971,N_2192,N_1889);
and U2972 (N_2972,N_1846,N_1748);
nor U2973 (N_2973,N_2230,N_1584);
nand U2974 (N_2974,N_1829,N_1521);
and U2975 (N_2975,N_1906,N_1745);
nor U2976 (N_2976,N_1623,N_2126);
nor U2977 (N_2977,N_1664,N_2236);
or U2978 (N_2978,N_1884,N_2238);
nand U2979 (N_2979,N_2100,N_1648);
nand U2980 (N_2980,N_1943,N_1726);
nor U2981 (N_2981,N_1806,N_1882);
or U2982 (N_2982,N_1577,N_2077);
nand U2983 (N_2983,N_2087,N_1633);
xor U2984 (N_2984,N_1570,N_1734);
and U2985 (N_2985,N_1920,N_1505);
or U2986 (N_2986,N_2166,N_1853);
and U2987 (N_2987,N_2097,N_1590);
nor U2988 (N_2988,N_2036,N_1637);
or U2989 (N_2989,N_2004,N_1743);
and U2990 (N_2990,N_1676,N_1976);
nand U2991 (N_2991,N_2023,N_2224);
nand U2992 (N_2992,N_2071,N_1562);
nand U2993 (N_2993,N_2122,N_2166);
nor U2994 (N_2994,N_1920,N_1698);
or U2995 (N_2995,N_2168,N_1906);
nor U2996 (N_2996,N_2177,N_1517);
and U2997 (N_2997,N_1831,N_1908);
or U2998 (N_2998,N_1991,N_1867);
nand U2999 (N_2999,N_1816,N_1909);
nand UO_0 (O_0,N_2319,N_2626);
nand UO_1 (O_1,N_2273,N_2337);
nor UO_2 (O_2,N_2706,N_2350);
xor UO_3 (O_3,N_2748,N_2871);
or UO_4 (O_4,N_2405,N_2901);
or UO_5 (O_5,N_2975,N_2549);
xor UO_6 (O_6,N_2996,N_2945);
nand UO_7 (O_7,N_2821,N_2278);
and UO_8 (O_8,N_2606,N_2963);
and UO_9 (O_9,N_2588,N_2538);
nand UO_10 (O_10,N_2299,N_2364);
or UO_11 (O_11,N_2305,N_2446);
and UO_12 (O_12,N_2516,N_2995);
or UO_13 (O_13,N_2585,N_2433);
or UO_14 (O_14,N_2367,N_2641);
or UO_15 (O_15,N_2680,N_2518);
and UO_16 (O_16,N_2991,N_2862);
nor UO_17 (O_17,N_2979,N_2852);
nor UO_18 (O_18,N_2455,N_2958);
nor UO_19 (O_19,N_2725,N_2489);
and UO_20 (O_20,N_2677,N_2726);
and UO_21 (O_21,N_2263,N_2481);
or UO_22 (O_22,N_2863,N_2339);
or UO_23 (O_23,N_2969,N_2389);
and UO_24 (O_24,N_2378,N_2357);
and UO_25 (O_25,N_2492,N_2262);
or UO_26 (O_26,N_2929,N_2987);
nand UO_27 (O_27,N_2272,N_2829);
nor UO_28 (O_28,N_2815,N_2940);
nor UO_29 (O_29,N_2794,N_2279);
nand UO_30 (O_30,N_2457,N_2832);
and UO_31 (O_31,N_2326,N_2632);
and UO_32 (O_32,N_2509,N_2539);
nand UO_33 (O_33,N_2698,N_2611);
or UO_34 (O_34,N_2296,N_2345);
and UO_35 (O_35,N_2406,N_2898);
or UO_36 (O_36,N_2351,N_2540);
and UO_37 (O_37,N_2820,N_2582);
nand UO_38 (O_38,N_2445,N_2301);
xor UO_39 (O_39,N_2847,N_2573);
nand UO_40 (O_40,N_2695,N_2724);
and UO_41 (O_41,N_2946,N_2289);
nand UO_42 (O_42,N_2255,N_2789);
or UO_43 (O_43,N_2572,N_2924);
and UO_44 (O_44,N_2383,N_2978);
or UO_45 (O_45,N_2436,N_2541);
nor UO_46 (O_46,N_2998,N_2435);
nor UO_47 (O_47,N_2989,N_2330);
nor UO_48 (O_48,N_2905,N_2561);
nor UO_49 (O_49,N_2268,N_2935);
nor UO_50 (O_50,N_2684,N_2407);
and UO_51 (O_51,N_2605,N_2896);
or UO_52 (O_52,N_2661,N_2762);
nand UO_53 (O_53,N_2625,N_2997);
and UO_54 (O_54,N_2798,N_2557);
or UO_55 (O_55,N_2964,N_2738);
or UO_56 (O_56,N_2442,N_2884);
xor UO_57 (O_57,N_2633,N_2918);
and UO_58 (O_58,N_2437,N_2379);
and UO_59 (O_59,N_2697,N_2463);
and UO_60 (O_60,N_2645,N_2913);
or UO_61 (O_61,N_2439,N_2259);
or UO_62 (O_62,N_2276,N_2535);
and UO_63 (O_63,N_2347,N_2285);
and UO_64 (O_64,N_2309,N_2552);
and UO_65 (O_65,N_2889,N_2258);
nor UO_66 (O_66,N_2709,N_2895);
xor UO_67 (O_67,N_2551,N_2643);
and UO_68 (O_68,N_2571,N_2728);
and UO_69 (O_69,N_2876,N_2949);
or UO_70 (O_70,N_2513,N_2515);
or UO_71 (O_71,N_2425,N_2747);
nand UO_72 (O_72,N_2479,N_2358);
and UO_73 (O_73,N_2560,N_2317);
nor UO_74 (O_74,N_2784,N_2772);
and UO_75 (O_75,N_2683,N_2360);
and UO_76 (O_76,N_2685,N_2976);
nand UO_77 (O_77,N_2736,N_2927);
and UO_78 (O_78,N_2498,N_2699);
or UO_79 (O_79,N_2939,N_2893);
nand UO_80 (O_80,N_2682,N_2866);
nand UO_81 (O_81,N_2835,N_2271);
or UO_82 (O_82,N_2579,N_2444);
nor UO_83 (O_83,N_2938,N_2542);
nor UO_84 (O_84,N_2912,N_2475);
nor UO_85 (O_85,N_2381,N_2600);
nor UO_86 (O_86,N_2374,N_2909);
nand UO_87 (O_87,N_2877,N_2595);
and UO_88 (O_88,N_2526,N_2828);
nor UO_89 (O_89,N_2752,N_2416);
nor UO_90 (O_90,N_2776,N_2274);
and UO_91 (O_91,N_2315,N_2947);
nand UO_92 (O_92,N_2759,N_2369);
and UO_93 (O_93,N_2570,N_2723);
nor UO_94 (O_94,N_2868,N_2521);
or UO_95 (O_95,N_2713,N_2950);
xnor UO_96 (O_96,N_2854,N_2373);
and UO_97 (O_97,N_2659,N_2966);
nand UO_98 (O_98,N_2607,N_2785);
or UO_99 (O_99,N_2779,N_2756);
and UO_100 (O_100,N_2720,N_2742);
nor UO_101 (O_101,N_2769,N_2393);
and UO_102 (O_102,N_2657,N_2660);
or UO_103 (O_103,N_2801,N_2974);
or UO_104 (O_104,N_2331,N_2994);
nand UO_105 (O_105,N_2848,N_2972);
or UO_106 (O_106,N_2608,N_2496);
and UO_107 (O_107,N_2456,N_2627);
nand UO_108 (O_108,N_2290,N_2493);
and UO_109 (O_109,N_2688,N_2412);
and UO_110 (O_110,N_2970,N_2257);
and UO_111 (O_111,N_2294,N_2454);
and UO_112 (O_112,N_2870,N_2715);
nor UO_113 (O_113,N_2780,N_2525);
and UO_114 (O_114,N_2327,N_2316);
and UO_115 (O_115,N_2527,N_2808);
nand UO_116 (O_116,N_2533,N_2420);
nand UO_117 (O_117,N_2477,N_2928);
and UO_118 (O_118,N_2624,N_2658);
and UO_119 (O_119,N_2623,N_2587);
and UO_120 (O_120,N_2662,N_2298);
or UO_121 (O_121,N_2593,N_2286);
nand UO_122 (O_122,N_2512,N_2691);
or UO_123 (O_123,N_2622,N_2719);
and UO_124 (O_124,N_2644,N_2517);
nor UO_125 (O_125,N_2550,N_2265);
and UO_126 (O_126,N_2615,N_2790);
or UO_127 (O_127,N_2745,N_2771);
nand UO_128 (O_128,N_2630,N_2892);
nor UO_129 (O_129,N_2348,N_2599);
and UO_130 (O_130,N_2921,N_2578);
or UO_131 (O_131,N_2450,N_2910);
or UO_132 (O_132,N_2459,N_2890);
and UO_133 (O_133,N_2440,N_2781);
nand UO_134 (O_134,N_2583,N_2911);
and UO_135 (O_135,N_2341,N_2831);
nand UO_136 (O_136,N_2320,N_2499);
nand UO_137 (O_137,N_2313,N_2386);
or UO_138 (O_138,N_2874,N_2734);
or UO_139 (O_139,N_2902,N_2618);
nand UO_140 (O_140,N_2842,N_2594);
nor UO_141 (O_141,N_2923,N_2311);
nand UO_142 (O_142,N_2400,N_2344);
nor UO_143 (O_143,N_2277,N_2312);
nand UO_144 (O_144,N_2300,N_2730);
or UO_145 (O_145,N_2639,N_2295);
nor UO_146 (O_146,N_2569,N_2554);
or UO_147 (O_147,N_2894,N_2335);
and UO_148 (O_148,N_2325,N_2384);
nand UO_149 (O_149,N_2729,N_2749);
nand UO_150 (O_150,N_2792,N_2447);
and UO_151 (O_151,N_2992,N_2774);
nor UO_152 (O_152,N_2291,N_2708);
nor UO_153 (O_153,N_2318,N_2967);
and UO_154 (O_154,N_2655,N_2601);
or UO_155 (O_155,N_2673,N_2401);
or UO_156 (O_156,N_2956,N_2507);
and UO_157 (O_157,N_2944,N_2636);
or UO_158 (O_158,N_2710,N_2960);
and UO_159 (O_159,N_2452,N_2332);
and UO_160 (O_160,N_2328,N_2553);
nor UO_161 (O_161,N_2778,N_2472);
or UO_162 (O_162,N_2506,N_2423);
nor UO_163 (O_163,N_2620,N_2505);
nand UO_164 (O_164,N_2687,N_2448);
and UO_165 (O_165,N_2765,N_2564);
or UO_166 (O_166,N_2767,N_2284);
nand UO_167 (O_167,N_2414,N_2413);
nor UO_168 (O_168,N_2656,N_2873);
and UO_169 (O_169,N_2418,N_2390);
nor UO_170 (O_170,N_2260,N_2635);
nand UO_171 (O_171,N_2322,N_2329);
nor UO_172 (O_172,N_2797,N_2908);
and UO_173 (O_173,N_2536,N_2629);
nand UO_174 (O_174,N_2486,N_2796);
nor UO_175 (O_175,N_2654,N_2899);
nand UO_176 (O_176,N_2356,N_2398);
nor UO_177 (O_177,N_2649,N_2529);
nand UO_178 (O_178,N_2597,N_2547);
or UO_179 (O_179,N_2504,N_2880);
nand UO_180 (O_180,N_2566,N_2668);
and UO_181 (O_181,N_2634,N_2758);
nand UO_182 (O_182,N_2856,N_2495);
or UO_183 (O_183,N_2882,N_2942);
and UO_184 (O_184,N_2665,N_2368);
nor UO_185 (O_185,N_2592,N_2333);
nand UO_186 (O_186,N_2689,N_2867);
nand UO_187 (O_187,N_2510,N_2556);
or UO_188 (O_188,N_2421,N_2482);
and UO_189 (O_189,N_2500,N_2469);
or UO_190 (O_190,N_2642,N_2371);
nand UO_191 (O_191,N_2883,N_2352);
and UO_192 (O_192,N_2380,N_2490);
nor UO_193 (O_193,N_2891,N_2844);
and UO_194 (O_194,N_2631,N_2543);
and UO_195 (O_195,N_2760,N_2650);
nor UO_196 (O_196,N_2932,N_2961);
nor UO_197 (O_197,N_2647,N_2993);
nor UO_198 (O_198,N_2256,N_2834);
nor UO_199 (O_199,N_2563,N_2596);
and UO_200 (O_200,N_2711,N_2814);
or UO_201 (O_201,N_2532,N_2805);
nand UO_202 (O_202,N_2838,N_2565);
and UO_203 (O_203,N_2669,N_2886);
nand UO_204 (O_204,N_2885,N_2735);
nor UO_205 (O_205,N_2485,N_2411);
and UO_206 (O_206,N_2743,N_2361);
or UO_207 (O_207,N_2422,N_2269);
or UO_208 (O_208,N_2514,N_2984);
or UO_209 (O_209,N_2755,N_2394);
nor UO_210 (O_210,N_2581,N_2840);
nor UO_211 (O_211,N_2354,N_2342);
nand UO_212 (O_212,N_2737,N_2845);
nor UO_213 (O_213,N_2793,N_2399);
nor UO_214 (O_214,N_2718,N_2590);
nand UO_215 (O_215,N_2451,N_2764);
and UO_216 (O_216,N_2846,N_2476);
and UO_217 (O_217,N_2519,N_2334);
nor UO_218 (O_218,N_2777,N_2283);
and UO_219 (O_219,N_2859,N_2251);
and UO_220 (O_220,N_2548,N_2621);
nor UO_221 (O_221,N_2810,N_2408);
or UO_222 (O_222,N_2403,N_2732);
and UO_223 (O_223,N_2575,N_2458);
nand UO_224 (O_224,N_2503,N_2474);
nand UO_225 (O_225,N_2799,N_2744);
nor UO_226 (O_226,N_2340,N_2520);
nor UO_227 (O_227,N_2302,N_2310);
xnor UO_228 (O_228,N_2982,N_2293);
or UO_229 (O_229,N_2919,N_2686);
or UO_230 (O_230,N_2707,N_2757);
or UO_231 (O_231,N_2468,N_2637);
nand UO_232 (O_232,N_2926,N_2449);
or UO_233 (O_233,N_2971,N_2395);
nor UO_234 (O_234,N_2851,N_2850);
nand UO_235 (O_235,N_2349,N_2679);
or UO_236 (O_236,N_2692,N_2544);
nor UO_237 (O_237,N_2574,N_2986);
nand UO_238 (O_238,N_2951,N_2343);
nand UO_239 (O_239,N_2616,N_2941);
nand UO_240 (O_240,N_2802,N_2487);
and UO_241 (O_241,N_2336,N_2836);
or UO_242 (O_242,N_2822,N_2775);
and UO_243 (O_243,N_2250,N_2528);
and UO_244 (O_244,N_2990,N_2973);
and UO_245 (O_245,N_2434,N_2537);
or UO_246 (O_246,N_2981,N_2702);
nor UO_247 (O_247,N_2304,N_2653);
nand UO_248 (O_248,N_2853,N_2717);
or UO_249 (O_249,N_2559,N_2704);
xor UO_250 (O_250,N_2488,N_2640);
nand UO_251 (O_251,N_2353,N_2672);
and UO_252 (O_252,N_2432,N_2508);
or UO_253 (O_253,N_2419,N_2524);
nand UO_254 (O_254,N_2453,N_2841);
nor UO_255 (O_255,N_2471,N_2746);
nand UO_256 (O_256,N_2827,N_2365);
nand UO_257 (O_257,N_2930,N_2462);
nor UO_258 (O_258,N_2470,N_2999);
or UO_259 (O_259,N_2270,N_2791);
or UO_260 (O_260,N_2813,N_2768);
nor UO_261 (O_261,N_2324,N_2965);
nor UO_262 (O_262,N_2690,N_2603);
nor UO_263 (O_263,N_2985,N_2703);
or UO_264 (O_264,N_2281,N_2617);
nor UO_265 (O_265,N_2375,N_2721);
nor UO_266 (O_266,N_2807,N_2376);
and UO_267 (O_267,N_2392,N_2288);
nand UO_268 (O_268,N_2555,N_2959);
or UO_269 (O_269,N_2604,N_2651);
nor UO_270 (O_270,N_2917,N_2819);
nand UO_271 (O_271,N_2837,N_2287);
or UO_272 (O_272,N_2962,N_2900);
or UO_273 (O_273,N_2700,N_2638);
and UO_274 (O_274,N_2714,N_2937);
nand UO_275 (O_275,N_2696,N_2598);
or UO_276 (O_276,N_2522,N_2646);
and UO_277 (O_277,N_2591,N_2580);
nor UO_278 (O_278,N_2740,N_2491);
nor UO_279 (O_279,N_2954,N_2830);
nand UO_280 (O_280,N_2786,N_2429);
and UO_281 (O_281,N_2292,N_2678);
or UO_282 (O_282,N_2465,N_2438);
or UO_283 (O_283,N_2417,N_2427);
and UO_284 (O_284,N_2818,N_2523);
and UO_285 (O_285,N_2410,N_2681);
or UO_286 (O_286,N_2826,N_2303);
or UO_287 (O_287,N_2428,N_2861);
nor UO_288 (O_288,N_2875,N_2614);
or UO_289 (O_289,N_2282,N_2473);
nor UO_290 (O_290,N_2731,N_2931);
nor UO_291 (O_291,N_2806,N_2602);
nor UO_292 (O_292,N_2359,N_2855);
nand UO_293 (O_293,N_2577,N_2860);
xor UO_294 (O_294,N_2628,N_2857);
and UO_295 (O_295,N_2788,N_2934);
or UO_296 (O_296,N_2671,N_2907);
and UO_297 (O_297,N_2568,N_2546);
nor UO_298 (O_298,N_2534,N_2693);
nor UO_299 (O_299,N_2409,N_2530);
and UO_300 (O_300,N_2576,N_2663);
xor UO_301 (O_301,N_2675,N_2988);
or UO_302 (O_302,N_2562,N_2253);
or UO_303 (O_303,N_2897,N_2906);
nor UO_304 (O_304,N_2297,N_2664);
or UO_305 (O_305,N_2402,N_2670);
nor UO_306 (O_306,N_2824,N_2502);
and UO_307 (O_307,N_2275,N_2957);
or UO_308 (O_308,N_2254,N_2461);
nand UO_309 (O_309,N_2694,N_2727);
and UO_310 (O_310,N_2404,N_2948);
nor UO_311 (O_311,N_2478,N_2466);
nand UO_312 (O_312,N_2610,N_2415);
nor UO_313 (O_313,N_2497,N_2494);
nand UO_314 (O_314,N_2612,N_2484);
and UO_315 (O_315,N_2916,N_2823);
and UO_316 (O_316,N_2952,N_2983);
nor UO_317 (O_317,N_2914,N_2722);
nand UO_318 (O_318,N_2280,N_2397);
and UO_319 (O_319,N_2346,N_2881);
or UO_320 (O_320,N_2589,N_2441);
nor UO_321 (O_321,N_2955,N_2266);
or UO_322 (O_322,N_2652,N_2787);
nand UO_323 (O_323,N_2980,N_2804);
nor UO_324 (O_324,N_2667,N_2306);
nor UO_325 (O_325,N_2531,N_2953);
and UO_326 (O_326,N_2977,N_2936);
or UO_327 (O_327,N_2872,N_2426);
and UO_328 (O_328,N_2716,N_2609);
nand UO_329 (O_329,N_2920,N_2878);
nor UO_330 (O_330,N_2809,N_2586);
nand UO_331 (O_331,N_2887,N_2362);
and UO_332 (O_332,N_2833,N_2812);
nor UO_333 (O_333,N_2323,N_2733);
or UO_334 (O_334,N_2584,N_2467);
and UO_335 (O_335,N_2355,N_2674);
or UO_336 (O_336,N_2267,N_2431);
or UO_337 (O_337,N_2825,N_2396);
nand UO_338 (O_338,N_2782,N_2869);
nor UO_339 (O_339,N_2858,N_2864);
or UO_340 (O_340,N_2558,N_2751);
or UO_341 (O_341,N_2816,N_2264);
or UO_342 (O_342,N_2314,N_2712);
nand UO_343 (O_343,N_2705,N_2372);
nand UO_344 (O_344,N_2922,N_2770);
and UO_345 (O_345,N_2308,N_2370);
nand UO_346 (O_346,N_2676,N_2817);
nor UO_347 (O_347,N_2803,N_2338);
nand UO_348 (O_348,N_2460,N_2753);
or UO_349 (O_349,N_2613,N_2511);
and UO_350 (O_350,N_2943,N_2501);
nor UO_351 (O_351,N_2619,N_2424);
xnor UO_352 (O_352,N_2391,N_2701);
nand UO_353 (O_353,N_2773,N_2443);
nand UO_354 (O_354,N_2795,N_2387);
nor UO_355 (O_355,N_2915,N_2483);
nand UO_356 (O_356,N_2933,N_2750);
or UO_357 (O_357,N_2366,N_2968);
or UO_358 (O_358,N_2567,N_2843);
or UO_359 (O_359,N_2363,N_2307);
and UO_360 (O_360,N_2925,N_2903);
nor UO_361 (O_361,N_2879,N_2763);
or UO_362 (O_362,N_2741,N_2261);
nand UO_363 (O_363,N_2464,N_2321);
and UO_364 (O_364,N_2252,N_2904);
nor UO_365 (O_365,N_2545,N_2480);
nand UO_366 (O_366,N_2839,N_2382);
or UO_367 (O_367,N_2388,N_2648);
nand UO_368 (O_368,N_2865,N_2783);
nor UO_369 (O_369,N_2888,N_2811);
nor UO_370 (O_370,N_2739,N_2849);
and UO_371 (O_371,N_2800,N_2430);
nor UO_372 (O_372,N_2766,N_2377);
or UO_373 (O_373,N_2761,N_2385);
or UO_374 (O_374,N_2754,N_2666);
nor UO_375 (O_375,N_2772,N_2595);
nand UO_376 (O_376,N_2606,N_2471);
and UO_377 (O_377,N_2857,N_2960);
nand UO_378 (O_378,N_2908,N_2752);
nor UO_379 (O_379,N_2644,N_2472);
or UO_380 (O_380,N_2874,N_2896);
xnor UO_381 (O_381,N_2279,N_2429);
and UO_382 (O_382,N_2342,N_2353);
nand UO_383 (O_383,N_2250,N_2681);
nand UO_384 (O_384,N_2802,N_2388);
or UO_385 (O_385,N_2808,N_2416);
nand UO_386 (O_386,N_2543,N_2376);
and UO_387 (O_387,N_2652,N_2259);
or UO_388 (O_388,N_2366,N_2986);
and UO_389 (O_389,N_2942,N_2296);
and UO_390 (O_390,N_2548,N_2671);
or UO_391 (O_391,N_2464,N_2651);
and UO_392 (O_392,N_2588,N_2667);
nand UO_393 (O_393,N_2406,N_2824);
nor UO_394 (O_394,N_2726,N_2810);
or UO_395 (O_395,N_2589,N_2629);
nor UO_396 (O_396,N_2753,N_2786);
nor UO_397 (O_397,N_2273,N_2546);
nand UO_398 (O_398,N_2416,N_2982);
nor UO_399 (O_399,N_2514,N_2481);
and UO_400 (O_400,N_2600,N_2989);
xor UO_401 (O_401,N_2324,N_2539);
nor UO_402 (O_402,N_2957,N_2701);
nand UO_403 (O_403,N_2377,N_2641);
nor UO_404 (O_404,N_2661,N_2494);
nand UO_405 (O_405,N_2699,N_2883);
and UO_406 (O_406,N_2797,N_2371);
nor UO_407 (O_407,N_2450,N_2830);
or UO_408 (O_408,N_2475,N_2385);
and UO_409 (O_409,N_2524,N_2710);
and UO_410 (O_410,N_2552,N_2693);
or UO_411 (O_411,N_2795,N_2440);
xnor UO_412 (O_412,N_2496,N_2556);
nand UO_413 (O_413,N_2487,N_2733);
nor UO_414 (O_414,N_2475,N_2921);
and UO_415 (O_415,N_2411,N_2496);
nor UO_416 (O_416,N_2373,N_2590);
nand UO_417 (O_417,N_2847,N_2699);
nor UO_418 (O_418,N_2655,N_2886);
nor UO_419 (O_419,N_2703,N_2643);
or UO_420 (O_420,N_2382,N_2568);
nor UO_421 (O_421,N_2499,N_2987);
nand UO_422 (O_422,N_2420,N_2696);
nand UO_423 (O_423,N_2266,N_2743);
and UO_424 (O_424,N_2690,N_2960);
or UO_425 (O_425,N_2869,N_2636);
and UO_426 (O_426,N_2596,N_2722);
nor UO_427 (O_427,N_2340,N_2578);
nor UO_428 (O_428,N_2392,N_2492);
nor UO_429 (O_429,N_2585,N_2639);
or UO_430 (O_430,N_2732,N_2825);
and UO_431 (O_431,N_2998,N_2394);
xor UO_432 (O_432,N_2571,N_2538);
or UO_433 (O_433,N_2619,N_2660);
and UO_434 (O_434,N_2695,N_2288);
nor UO_435 (O_435,N_2545,N_2713);
nor UO_436 (O_436,N_2450,N_2837);
or UO_437 (O_437,N_2765,N_2674);
or UO_438 (O_438,N_2399,N_2708);
nand UO_439 (O_439,N_2965,N_2276);
or UO_440 (O_440,N_2643,N_2980);
nand UO_441 (O_441,N_2890,N_2559);
and UO_442 (O_442,N_2662,N_2924);
or UO_443 (O_443,N_2517,N_2375);
nand UO_444 (O_444,N_2744,N_2675);
or UO_445 (O_445,N_2488,N_2870);
nor UO_446 (O_446,N_2279,N_2446);
and UO_447 (O_447,N_2986,N_2724);
nor UO_448 (O_448,N_2777,N_2871);
nand UO_449 (O_449,N_2796,N_2421);
and UO_450 (O_450,N_2426,N_2817);
nor UO_451 (O_451,N_2336,N_2539);
and UO_452 (O_452,N_2881,N_2397);
nand UO_453 (O_453,N_2913,N_2842);
nor UO_454 (O_454,N_2589,N_2701);
nand UO_455 (O_455,N_2848,N_2433);
and UO_456 (O_456,N_2361,N_2619);
nor UO_457 (O_457,N_2684,N_2783);
and UO_458 (O_458,N_2495,N_2646);
nand UO_459 (O_459,N_2664,N_2372);
nand UO_460 (O_460,N_2709,N_2711);
nor UO_461 (O_461,N_2492,N_2837);
nor UO_462 (O_462,N_2360,N_2886);
nor UO_463 (O_463,N_2932,N_2443);
and UO_464 (O_464,N_2632,N_2972);
nor UO_465 (O_465,N_2486,N_2844);
nor UO_466 (O_466,N_2546,N_2401);
nand UO_467 (O_467,N_2286,N_2500);
or UO_468 (O_468,N_2263,N_2368);
nand UO_469 (O_469,N_2255,N_2960);
nor UO_470 (O_470,N_2759,N_2747);
nor UO_471 (O_471,N_2800,N_2649);
nor UO_472 (O_472,N_2468,N_2635);
and UO_473 (O_473,N_2739,N_2484);
or UO_474 (O_474,N_2305,N_2336);
nand UO_475 (O_475,N_2278,N_2405);
nand UO_476 (O_476,N_2425,N_2522);
nand UO_477 (O_477,N_2365,N_2535);
or UO_478 (O_478,N_2822,N_2574);
nor UO_479 (O_479,N_2609,N_2332);
nand UO_480 (O_480,N_2272,N_2765);
nand UO_481 (O_481,N_2919,N_2578);
nand UO_482 (O_482,N_2999,N_2808);
nor UO_483 (O_483,N_2426,N_2463);
nor UO_484 (O_484,N_2658,N_2466);
nor UO_485 (O_485,N_2993,N_2865);
and UO_486 (O_486,N_2268,N_2661);
and UO_487 (O_487,N_2883,N_2570);
or UO_488 (O_488,N_2660,N_2937);
or UO_489 (O_489,N_2965,N_2635);
nor UO_490 (O_490,N_2990,N_2282);
or UO_491 (O_491,N_2363,N_2875);
nor UO_492 (O_492,N_2468,N_2872);
or UO_493 (O_493,N_2513,N_2722);
or UO_494 (O_494,N_2904,N_2264);
and UO_495 (O_495,N_2462,N_2796);
nand UO_496 (O_496,N_2997,N_2980);
and UO_497 (O_497,N_2896,N_2900);
nand UO_498 (O_498,N_2586,N_2672);
xnor UO_499 (O_499,N_2829,N_2521);
endmodule