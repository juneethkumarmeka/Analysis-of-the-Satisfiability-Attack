module basic_750_5000_1000_25_levels_5xor_8(In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749,O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999);
input In_0,In_1,In_2,In_3,In_4,In_5,In_6,In_7,In_8,In_9,In_10,In_11,In_12,In_13,In_14,In_15,In_16,In_17,In_18,In_19,In_20,In_21,In_22,In_23,In_24,In_25,In_26,In_27,In_28,In_29,In_30,In_31,In_32,In_33,In_34,In_35,In_36,In_37,In_38,In_39,In_40,In_41,In_42,In_43,In_44,In_45,In_46,In_47,In_48,In_49,In_50,In_51,In_52,In_53,In_54,In_55,In_56,In_57,In_58,In_59,In_60,In_61,In_62,In_63,In_64,In_65,In_66,In_67,In_68,In_69,In_70,In_71,In_72,In_73,In_74,In_75,In_76,In_77,In_78,In_79,In_80,In_81,In_82,In_83,In_84,In_85,In_86,In_87,In_88,In_89,In_90,In_91,In_92,In_93,In_94,In_95,In_96,In_97,In_98,In_99,In_100,In_101,In_102,In_103,In_104,In_105,In_106,In_107,In_108,In_109,In_110,In_111,In_112,In_113,In_114,In_115,In_116,In_117,In_118,In_119,In_120,In_121,In_122,In_123,In_124,In_125,In_126,In_127,In_128,In_129,In_130,In_131,In_132,In_133,In_134,In_135,In_136,In_137,In_138,In_139,In_140,In_141,In_142,In_143,In_144,In_145,In_146,In_147,In_148,In_149,In_150,In_151,In_152,In_153,In_154,In_155,In_156,In_157,In_158,In_159,In_160,In_161,In_162,In_163,In_164,In_165,In_166,In_167,In_168,In_169,In_170,In_171,In_172,In_173,In_174,In_175,In_176,In_177,In_178,In_179,In_180,In_181,In_182,In_183,In_184,In_185,In_186,In_187,In_188,In_189,In_190,In_191,In_192,In_193,In_194,In_195,In_196,In_197,In_198,In_199,In_200,In_201,In_202,In_203,In_204,In_205,In_206,In_207,In_208,In_209,In_210,In_211,In_212,In_213,In_214,In_215,In_216,In_217,In_218,In_219,In_220,In_221,In_222,In_223,In_224,In_225,In_226,In_227,In_228,In_229,In_230,In_231,In_232,In_233,In_234,In_235,In_236,In_237,In_238,In_239,In_240,In_241,In_242,In_243,In_244,In_245,In_246,In_247,In_248,In_249,In_250,In_251,In_252,In_253,In_254,In_255,In_256,In_257,In_258,In_259,In_260,In_261,In_262,In_263,In_264,In_265,In_266,In_267,In_268,In_269,In_270,In_271,In_272,In_273,In_274,In_275,In_276,In_277,In_278,In_279,In_280,In_281,In_282,In_283,In_284,In_285,In_286,In_287,In_288,In_289,In_290,In_291,In_292,In_293,In_294,In_295,In_296,In_297,In_298,In_299,In_300,In_301,In_302,In_303,In_304,In_305,In_306,In_307,In_308,In_309,In_310,In_311,In_312,In_313,In_314,In_315,In_316,In_317,In_318,In_319,In_320,In_321,In_322,In_323,In_324,In_325,In_326,In_327,In_328,In_329,In_330,In_331,In_332,In_333,In_334,In_335,In_336,In_337,In_338,In_339,In_340,In_341,In_342,In_343,In_344,In_345,In_346,In_347,In_348,In_349,In_350,In_351,In_352,In_353,In_354,In_355,In_356,In_357,In_358,In_359,In_360,In_361,In_362,In_363,In_364,In_365,In_366,In_367,In_368,In_369,In_370,In_371,In_372,In_373,In_374,In_375,In_376,In_377,In_378,In_379,In_380,In_381,In_382,In_383,In_384,In_385,In_386,In_387,In_388,In_389,In_390,In_391,In_392,In_393,In_394,In_395,In_396,In_397,In_398,In_399,In_400,In_401,In_402,In_403,In_404,In_405,In_406,In_407,In_408,In_409,In_410,In_411,In_412,In_413,In_414,In_415,In_416,In_417,In_418,In_419,In_420,In_421,In_422,In_423,In_424,In_425,In_426,In_427,In_428,In_429,In_430,In_431,In_432,In_433,In_434,In_435,In_436,In_437,In_438,In_439,In_440,In_441,In_442,In_443,In_444,In_445,In_446,In_447,In_448,In_449,In_450,In_451,In_452,In_453,In_454,In_455,In_456,In_457,In_458,In_459,In_460,In_461,In_462,In_463,In_464,In_465,In_466,In_467,In_468,In_469,In_470,In_471,In_472,In_473,In_474,In_475,In_476,In_477,In_478,In_479,In_480,In_481,In_482,In_483,In_484,In_485,In_486,In_487,In_488,In_489,In_490,In_491,In_492,In_493,In_494,In_495,In_496,In_497,In_498,In_499,In_500,In_501,In_502,In_503,In_504,In_505,In_506,In_507,In_508,In_509,In_510,In_511,In_512,In_513,In_514,In_515,In_516,In_517,In_518,In_519,In_520,In_521,In_522,In_523,In_524,In_525,In_526,In_527,In_528,In_529,In_530,In_531,In_532,In_533,In_534,In_535,In_536,In_537,In_538,In_539,In_540,In_541,In_542,In_543,In_544,In_545,In_546,In_547,In_548,In_549,In_550,In_551,In_552,In_553,In_554,In_555,In_556,In_557,In_558,In_559,In_560,In_561,In_562,In_563,In_564,In_565,In_566,In_567,In_568,In_569,In_570,In_571,In_572,In_573,In_574,In_575,In_576,In_577,In_578,In_579,In_580,In_581,In_582,In_583,In_584,In_585,In_586,In_587,In_588,In_589,In_590,In_591,In_592,In_593,In_594,In_595,In_596,In_597,In_598,In_599,In_600,In_601,In_602,In_603,In_604,In_605,In_606,In_607,In_608,In_609,In_610,In_611,In_612,In_613,In_614,In_615,In_616,In_617,In_618,In_619,In_620,In_621,In_622,In_623,In_624,In_625,In_626,In_627,In_628,In_629,In_630,In_631,In_632,In_633,In_634,In_635,In_636,In_637,In_638,In_639,In_640,In_641,In_642,In_643,In_644,In_645,In_646,In_647,In_648,In_649,In_650,In_651,In_652,In_653,In_654,In_655,In_656,In_657,In_658,In_659,In_660,In_661,In_662,In_663,In_664,In_665,In_666,In_667,In_668,In_669,In_670,In_671,In_672,In_673,In_674,In_675,In_676,In_677,In_678,In_679,In_680,In_681,In_682,In_683,In_684,In_685,In_686,In_687,In_688,In_689,In_690,In_691,In_692,In_693,In_694,In_695,In_696,In_697,In_698,In_699,In_700,In_701,In_702,In_703,In_704,In_705,In_706,In_707,In_708,In_709,In_710,In_711,In_712,In_713,In_714,In_715,In_716,In_717,In_718,In_719,In_720,In_721,In_722,In_723,In_724,In_725,In_726,In_727,In_728,In_729,In_730,In_731,In_732,In_733,In_734,In_735,In_736,In_737,In_738,In_739,In_740,In_741,In_742,In_743,In_744,In_745,In_746,In_747,In_748,In_749;
output O_0,O_1,O_2,O_3,O_4,O_5,O_6,O_7,O_8,O_9,O_10,O_11,O_12,O_13,O_14,O_15,O_16,O_17,O_18,O_19,O_20,O_21,O_22,O_23,O_24,O_25,O_26,O_27,O_28,O_29,O_30,O_31,O_32,O_33,O_34,O_35,O_36,O_37,O_38,O_39,O_40,O_41,O_42,O_43,O_44,O_45,O_46,O_47,O_48,O_49,O_50,O_51,O_52,O_53,O_54,O_55,O_56,O_57,O_58,O_59,O_60,O_61,O_62,O_63,O_64,O_65,O_66,O_67,O_68,O_69,O_70,O_71,O_72,O_73,O_74,O_75,O_76,O_77,O_78,O_79,O_80,O_81,O_82,O_83,O_84,O_85,O_86,O_87,O_88,O_89,O_90,O_91,O_92,O_93,O_94,O_95,O_96,O_97,O_98,O_99,O_100,O_101,O_102,O_103,O_104,O_105,O_106,O_107,O_108,O_109,O_110,O_111,O_112,O_113,O_114,O_115,O_116,O_117,O_118,O_119,O_120,O_121,O_122,O_123,O_124,O_125,O_126,O_127,O_128,O_129,O_130,O_131,O_132,O_133,O_134,O_135,O_136,O_137,O_138,O_139,O_140,O_141,O_142,O_143,O_144,O_145,O_146,O_147,O_148,O_149,O_150,O_151,O_152,O_153,O_154,O_155,O_156,O_157,O_158,O_159,O_160,O_161,O_162,O_163,O_164,O_165,O_166,O_167,O_168,O_169,O_170,O_171,O_172,O_173,O_174,O_175,O_176,O_177,O_178,O_179,O_180,O_181,O_182,O_183,O_184,O_185,O_186,O_187,O_188,O_189,O_190,O_191,O_192,O_193,O_194,O_195,O_196,O_197,O_198,O_199,O_200,O_201,O_202,O_203,O_204,O_205,O_206,O_207,O_208,O_209,O_210,O_211,O_212,O_213,O_214,O_215,O_216,O_217,O_218,O_219,O_220,O_221,O_222,O_223,O_224,O_225,O_226,O_227,O_228,O_229,O_230,O_231,O_232,O_233,O_234,O_235,O_236,O_237,O_238,O_239,O_240,O_241,O_242,O_243,O_244,O_245,O_246,O_247,O_248,O_249,O_250,O_251,O_252,O_253,O_254,O_255,O_256,O_257,O_258,O_259,O_260,O_261,O_262,O_263,O_264,O_265,O_266,O_267,O_268,O_269,O_270,O_271,O_272,O_273,O_274,O_275,O_276,O_277,O_278,O_279,O_280,O_281,O_282,O_283,O_284,O_285,O_286,O_287,O_288,O_289,O_290,O_291,O_292,O_293,O_294,O_295,O_296,O_297,O_298,O_299,O_300,O_301,O_302,O_303,O_304,O_305,O_306,O_307,O_308,O_309,O_310,O_311,O_312,O_313,O_314,O_315,O_316,O_317,O_318,O_319,O_320,O_321,O_322,O_323,O_324,O_325,O_326,O_327,O_328,O_329,O_330,O_331,O_332,O_333,O_334,O_335,O_336,O_337,O_338,O_339,O_340,O_341,O_342,O_343,O_344,O_345,O_346,O_347,O_348,O_349,O_350,O_351,O_352,O_353,O_354,O_355,O_356,O_357,O_358,O_359,O_360,O_361,O_362,O_363,O_364,O_365,O_366,O_367,O_368,O_369,O_370,O_371,O_372,O_373,O_374,O_375,O_376,O_377,O_378,O_379,O_380,O_381,O_382,O_383,O_384,O_385,O_386,O_387,O_388,O_389,O_390,O_391,O_392,O_393,O_394,O_395,O_396,O_397,O_398,O_399,O_400,O_401,O_402,O_403,O_404,O_405,O_406,O_407,O_408,O_409,O_410,O_411,O_412,O_413,O_414,O_415,O_416,O_417,O_418,O_419,O_420,O_421,O_422,O_423,O_424,O_425,O_426,O_427,O_428,O_429,O_430,O_431,O_432,O_433,O_434,O_435,O_436,O_437,O_438,O_439,O_440,O_441,O_442,O_443,O_444,O_445,O_446,O_447,O_448,O_449,O_450,O_451,O_452,O_453,O_454,O_455,O_456,O_457,O_458,O_459,O_460,O_461,O_462,O_463,O_464,O_465,O_466,O_467,O_468,O_469,O_470,O_471,O_472,O_473,O_474,O_475,O_476,O_477,O_478,O_479,O_480,O_481,O_482,O_483,O_484,O_485,O_486,O_487,O_488,O_489,O_490,O_491,O_492,O_493,O_494,O_495,O_496,O_497,O_498,O_499,O_500,O_501,O_502,O_503,O_504,O_505,O_506,O_507,O_508,O_509,O_510,O_511,O_512,O_513,O_514,O_515,O_516,O_517,O_518,O_519,O_520,O_521,O_522,O_523,O_524,O_525,O_526,O_527,O_528,O_529,O_530,O_531,O_532,O_533,O_534,O_535,O_536,O_537,O_538,O_539,O_540,O_541,O_542,O_543,O_544,O_545,O_546,O_547,O_548,O_549,O_550,O_551,O_552,O_553,O_554,O_555,O_556,O_557,O_558,O_559,O_560,O_561,O_562,O_563,O_564,O_565,O_566,O_567,O_568,O_569,O_570,O_571,O_572,O_573,O_574,O_575,O_576,O_577,O_578,O_579,O_580,O_581,O_582,O_583,O_584,O_585,O_586,O_587,O_588,O_589,O_590,O_591,O_592,O_593,O_594,O_595,O_596,O_597,O_598,O_599,O_600,O_601,O_602,O_603,O_604,O_605,O_606,O_607,O_608,O_609,O_610,O_611,O_612,O_613,O_614,O_615,O_616,O_617,O_618,O_619,O_620,O_621,O_622,O_623,O_624,O_625,O_626,O_627,O_628,O_629,O_630,O_631,O_632,O_633,O_634,O_635,O_636,O_637,O_638,O_639,O_640,O_641,O_642,O_643,O_644,O_645,O_646,O_647,O_648,O_649,O_650,O_651,O_652,O_653,O_654,O_655,O_656,O_657,O_658,O_659,O_660,O_661,O_662,O_663,O_664,O_665,O_666,O_667,O_668,O_669,O_670,O_671,O_672,O_673,O_674,O_675,O_676,O_677,O_678,O_679,O_680,O_681,O_682,O_683,O_684,O_685,O_686,O_687,O_688,O_689,O_690,O_691,O_692,O_693,O_694,O_695,O_696,O_697,O_698,O_699,O_700,O_701,O_702,O_703,O_704,O_705,O_706,O_707,O_708,O_709,O_710,O_711,O_712,O_713,O_714,O_715,O_716,O_717,O_718,O_719,O_720,O_721,O_722,O_723,O_724,O_725,O_726,O_727,O_728,O_729,O_730,O_731,O_732,O_733,O_734,O_735,O_736,O_737,O_738,O_739,O_740,O_741,O_742,O_743,O_744,O_745,O_746,O_747,O_748,O_749,O_750,O_751,O_752,O_753,O_754,O_755,O_756,O_757,O_758,O_759,O_760,O_761,O_762,O_763,O_764,O_765,O_766,O_767,O_768,O_769,O_770,O_771,O_772,O_773,O_774,O_775,O_776,O_777,O_778,O_779,O_780,O_781,O_782,O_783,O_784,O_785,O_786,O_787,O_788,O_789,O_790,O_791,O_792,O_793,O_794,O_795,O_796,O_797,O_798,O_799,O_800,O_801,O_802,O_803,O_804,O_805,O_806,O_807,O_808,O_809,O_810,O_811,O_812,O_813,O_814,O_815,O_816,O_817,O_818,O_819,O_820,O_821,O_822,O_823,O_824,O_825,O_826,O_827,O_828,O_829,O_830,O_831,O_832,O_833,O_834,O_835,O_836,O_837,O_838,O_839,O_840,O_841,O_842,O_843,O_844,O_845,O_846,O_847,O_848,O_849,O_850,O_851,O_852,O_853,O_854,O_855,O_856,O_857,O_858,O_859,O_860,O_861,O_862,O_863,O_864,O_865,O_866,O_867,O_868,O_869,O_870,O_871,O_872,O_873,O_874,O_875,O_876,O_877,O_878,O_879,O_880,O_881,O_882,O_883,O_884,O_885,O_886,O_887,O_888,O_889,O_890,O_891,O_892,O_893,O_894,O_895,O_896,O_897,O_898,O_899,O_900,O_901,O_902,O_903,O_904,O_905,O_906,O_907,O_908,O_909,O_910,O_911,O_912,O_913,O_914,O_915,O_916,O_917,O_918,O_919,O_920,O_921,O_922,O_923,O_924,O_925,O_926,O_927,O_928,O_929,O_930,O_931,O_932,O_933,O_934,O_935,O_936,O_937,O_938,O_939,O_940,O_941,O_942,O_943,O_944,O_945,O_946,O_947,O_948,O_949,O_950,O_951,O_952,O_953,O_954,O_955,O_956,O_957,O_958,O_959,O_960,O_961,O_962,O_963,O_964,O_965,O_966,O_967,O_968,O_969,O_970,O_971,O_972,O_973,O_974,O_975,O_976,O_977,O_978,O_979,O_980,O_981,O_982,O_983,O_984,O_985,O_986,O_987,O_988,O_989,O_990,O_991,O_992,O_993,O_994,O_995,O_996,O_997,O_998,O_999;
wire N_0,N_1,N_2,N_3,N_4,N_5,N_6,N_7,N_8,N_9,N_10,N_11,N_12,N_13,N_14,N_15,N_16,N_17,N_18,N_19,N_20,N_21,N_22,N_23,N_24,N_25,N_26,N_27,N_28,N_29,N_30,N_31,N_32,N_33,N_34,N_35,N_36,N_37,N_38,N_39,N_40,N_41,N_42,N_43,N_44,N_45,N_46,N_47,N_48,N_49,N_50,N_51,N_52,N_53,N_54,N_55,N_56,N_57,N_58,N_59,N_60,N_61,N_62,N_63,N_64,N_65,N_66,N_67,N_68,N_69,N_70,N_71,N_72,N_73,N_74,N_75,N_76,N_77,N_78,N_79,N_80,N_81,N_82,N_83,N_84,N_85,N_86,N_87,N_88,N_89,N_90,N_91,N_92,N_93,N_94,N_95,N_96,N_97,N_98,N_99,N_100,N_101,N_102,N_103,N_104,N_105,N_106,N_107,N_108,N_109,N_110,N_111,N_112,N_113,N_114,N_115,N_116,N_117,N_118,N_119,N_120,N_121,N_122,N_123,N_124,N_125,N_126,N_127,N_128,N_129,N_130,N_131,N_132,N_133,N_134,N_135,N_136,N_137,N_138,N_139,N_140,N_141,N_142,N_143,N_144,N_145,N_146,N_147,N_148,N_149,N_150,N_151,N_152,N_153,N_154,N_155,N_156,N_157,N_158,N_159,N_160,N_161,N_162,N_163,N_164,N_165,N_166,N_167,N_168,N_169,N_170,N_171,N_172,N_173,N_174,N_175,N_176,N_177,N_178,N_179,N_180,N_181,N_182,N_183,N_184,N_185,N_186,N_187,N_188,N_189,N_190,N_191,N_192,N_193,N_194,N_195,N_196,N_197,N_198,N_199,N_200,N_201,N_202,N_203,N_204,N_205,N_206,N_207,N_208,N_209,N_210,N_211,N_212,N_213,N_214,N_215,N_216,N_217,N_218,N_219,N_220,N_221,N_222,N_223,N_224,N_225,N_226,N_227,N_228,N_229,N_230,N_231,N_232,N_233,N_234,N_235,N_236,N_237,N_238,N_239,N_240,N_241,N_242,N_243,N_244,N_245,N_246,N_247,N_248,N_249,N_250,N_251,N_252,N_253,N_254,N_255,N_256,N_257,N_258,N_259,N_260,N_261,N_262,N_263,N_264,N_265,N_266,N_267,N_268,N_269,N_270,N_271,N_272,N_273,N_274,N_275,N_276,N_277,N_278,N_279,N_280,N_281,N_282,N_283,N_284,N_285,N_286,N_287,N_288,N_289,N_290,N_291,N_292,N_293,N_294,N_295,N_296,N_297,N_298,N_299,N_300,N_301,N_302,N_303,N_304,N_305,N_306,N_307,N_308,N_309,N_310,N_311,N_312,N_313,N_314,N_315,N_316,N_317,N_318,N_319,N_320,N_321,N_322,N_323,N_324,N_325,N_326,N_327,N_328,N_329,N_330,N_331,N_332,N_333,N_334,N_335,N_336,N_337,N_338,N_339,N_340,N_341,N_342,N_343,N_344,N_345,N_346,N_347,N_348,N_349,N_350,N_351,N_352,N_353,N_354,N_355,N_356,N_357,N_358,N_359,N_360,N_361,N_362,N_363,N_364,N_365,N_366,N_367,N_368,N_369,N_370,N_371,N_372,N_373,N_374,N_375,N_376,N_377,N_378,N_379,N_380,N_381,N_382,N_383,N_384,N_385,N_386,N_387,N_388,N_389,N_390,N_391,N_392,N_393,N_394,N_395,N_396,N_397,N_398,N_399,N_400,N_401,N_402,N_403,N_404,N_405,N_406,N_407,N_408,N_409,N_410,N_411,N_412,N_413,N_414,N_415,N_416,N_417,N_418,N_419,N_420,N_421,N_422,N_423,N_424,N_425,N_426,N_427,N_428,N_429,N_430,N_431,N_432,N_433,N_434,N_435,N_436,N_437,N_438,N_439,N_440,N_441,N_442,N_443,N_444,N_445,N_446,N_447,N_448,N_449,N_450,N_451,N_452,N_453,N_454,N_455,N_456,N_457,N_458,N_459,N_460,N_461,N_462,N_463,N_464,N_465,N_466,N_467,N_468,N_469,N_470,N_471,N_472,N_473,N_474,N_475,N_476,N_477,N_478,N_479,N_480,N_481,N_482,N_483,N_484,N_485,N_486,N_487,N_488,N_489,N_490,N_491,N_492,N_493,N_494,N_495,N_496,N_497,N_498,N_499,N_500,N_501,N_502,N_503,N_504,N_505,N_506,N_507,N_508,N_509,N_510,N_511,N_512,N_513,N_514,N_515,N_516,N_517,N_518,N_519,N_520,N_521,N_522,N_523,N_524,N_525,N_526,N_527,N_528,N_529,N_530,N_531,N_532,N_533,N_534,N_535,N_536,N_537,N_538,N_539,N_540,N_541,N_542,N_543,N_544,N_545,N_546,N_547,N_548,N_549,N_550,N_551,N_552,N_553,N_554,N_555,N_556,N_557,N_558,N_559,N_560,N_561,N_562,N_563,N_564,N_565,N_566,N_567,N_568,N_569,N_570,N_571,N_572,N_573,N_574,N_575,N_576,N_577,N_578,N_579,N_580,N_581,N_582,N_583,N_584,N_585,N_586,N_587,N_588,N_589,N_590,N_591,N_592,N_593,N_594,N_595,N_596,N_597,N_598,N_599,N_600,N_601,N_602,N_603,N_604,N_605,N_606,N_607,N_608,N_609,N_610,N_611,N_612,N_613,N_614,N_615,N_616,N_617,N_618,N_619,N_620,N_621,N_622,N_623,N_624,N_625,N_626,N_627,N_628,N_629,N_630,N_631,N_632,N_633,N_634,N_635,N_636,N_637,N_638,N_639,N_640,N_641,N_642,N_643,N_644,N_645,N_646,N_647,N_648,N_649,N_650,N_651,N_652,N_653,N_654,N_655,N_656,N_657,N_658,N_659,N_660,N_661,N_662,N_663,N_664,N_665,N_666,N_667,N_668,N_669,N_670,N_671,N_672,N_673,N_674,N_675,N_676,N_677,N_678,N_679,N_680,N_681,N_682,N_683,N_684,N_685,N_686,N_687,N_688,N_689,N_690,N_691,N_692,N_693,N_694,N_695,N_696,N_697,N_698,N_699,N_700,N_701,N_702,N_703,N_704,N_705,N_706,N_707,N_708,N_709,N_710,N_711,N_712,N_713,N_714,N_715,N_716,N_717,N_718,N_719,N_720,N_721,N_722,N_723,N_724,N_725,N_726,N_727,N_728,N_729,N_730,N_731,N_732,N_733,N_734,N_735,N_736,N_737,N_738,N_739,N_740,N_741,N_742,N_743,N_744,N_745,N_746,N_747,N_748,N_749,N_750,N_751,N_752,N_753,N_754,N_755,N_756,N_757,N_758,N_759,N_760,N_761,N_762,N_763,N_764,N_765,N_766,N_767,N_768,N_769,N_770,N_771,N_772,N_773,N_774,N_775,N_776,N_777,N_778,N_779,N_780,N_781,N_782,N_783,N_784,N_785,N_786,N_787,N_788,N_789,N_790,N_791,N_792,N_793,N_794,N_795,N_796,N_797,N_798,N_799,N_800,N_801,N_802,N_803,N_804,N_805,N_806,N_807,N_808,N_809,N_810,N_811,N_812,N_813,N_814,N_815,N_816,N_817,N_818,N_819,N_820,N_821,N_822,N_823,N_824,N_825,N_826,N_827,N_828,N_829,N_830,N_831,N_832,N_833,N_834,N_835,N_836,N_837,N_838,N_839,N_840,N_841,N_842,N_843,N_844,N_845,N_846,N_847,N_848,N_849,N_850,N_851,N_852,N_853,N_854,N_855,N_856,N_857,N_858,N_859,N_860,N_861,N_862,N_863,N_864,N_865,N_866,N_867,N_868,N_869,N_870,N_871,N_872,N_873,N_874,N_875,N_876,N_877,N_878,N_879,N_880,N_881,N_882,N_883,N_884,N_885,N_886,N_887,N_888,N_889,N_890,N_891,N_892,N_893,N_894,N_895,N_896,N_897,N_898,N_899,N_900,N_901,N_902,N_903,N_904,N_905,N_906,N_907,N_908,N_909,N_910,N_911,N_912,N_913,N_914,N_915,N_916,N_917,N_918,N_919,N_920,N_921,N_922,N_923,N_924,N_925,N_926,N_927,N_928,N_929,N_930,N_931,N_932,N_933,N_934,N_935,N_936,N_937,N_938,N_939,N_940,N_941,N_942,N_943,N_944,N_945,N_946,N_947,N_948,N_949,N_950,N_951,N_952,N_953,N_954,N_955,N_956,N_957,N_958,N_959,N_960,N_961,N_962,N_963,N_964,N_965,N_966,N_967,N_968,N_969,N_970,N_971,N_972,N_973,N_974,N_975,N_976,N_977,N_978,N_979,N_980,N_981,N_982,N_983,N_984,N_985,N_986,N_987,N_988,N_989,N_990,N_991,N_992,N_993,N_994,N_995,N_996,N_997,N_998,N_999,N_1000,N_1001,N_1002,N_1003,N_1004,N_1005,N_1006,N_1007,N_1008,N_1009,N_1010,N_1011,N_1012,N_1013,N_1014,N_1015,N_1016,N_1017,N_1018,N_1019,N_1020,N_1021,N_1022,N_1023,N_1024,N_1025,N_1026,N_1027,N_1028,N_1029,N_1030,N_1031,N_1032,N_1033,N_1034,N_1035,N_1036,N_1037,N_1038,N_1039,N_1040,N_1041,N_1042,N_1043,N_1044,N_1045,N_1046,N_1047,N_1048,N_1049,N_1050,N_1051,N_1052,N_1053,N_1054,N_1055,N_1056,N_1057,N_1058,N_1059,N_1060,N_1061,N_1062,N_1063,N_1064,N_1065,N_1066,N_1067,N_1068,N_1069,N_1070,N_1071,N_1072,N_1073,N_1074,N_1075,N_1076,N_1077,N_1078,N_1079,N_1080,N_1081,N_1082,N_1083,N_1084,N_1085,N_1086,N_1087,N_1088,N_1089,N_1090,N_1091,N_1092,N_1093,N_1094,N_1095,N_1096,N_1097,N_1098,N_1099,N_1100,N_1101,N_1102,N_1103,N_1104,N_1105,N_1106,N_1107,N_1108,N_1109,N_1110,N_1111,N_1112,N_1113,N_1114,N_1115,N_1116,N_1117,N_1118,N_1119,N_1120,N_1121,N_1122,N_1123,N_1124,N_1125,N_1126,N_1127,N_1128,N_1129,N_1130,N_1131,N_1132,N_1133,N_1134,N_1135,N_1136,N_1137,N_1138,N_1139,N_1140,N_1141,N_1142,N_1143,N_1144,N_1145,N_1146,N_1147,N_1148,N_1149,N_1150,N_1151,N_1152,N_1153,N_1154,N_1155,N_1156,N_1157,N_1158,N_1159,N_1160,N_1161,N_1162,N_1163,N_1164,N_1165,N_1166,N_1167,N_1168,N_1169,N_1170,N_1171,N_1172,N_1173,N_1174,N_1175,N_1176,N_1177,N_1178,N_1179,N_1180,N_1181,N_1182,N_1183,N_1184,N_1185,N_1186,N_1187,N_1188,N_1189,N_1190,N_1191,N_1192,N_1193,N_1194,N_1195,N_1196,N_1197,N_1198,N_1199,N_1200,N_1201,N_1202,N_1203,N_1204,N_1205,N_1206,N_1207,N_1208,N_1209,N_1210,N_1211,N_1212,N_1213,N_1214,N_1215,N_1216,N_1217,N_1218,N_1219,N_1220,N_1221,N_1222,N_1223,N_1224,N_1225,N_1226,N_1227,N_1228,N_1229,N_1230,N_1231,N_1232,N_1233,N_1234,N_1235,N_1236,N_1237,N_1238,N_1239,N_1240,N_1241,N_1242,N_1243,N_1244,N_1245,N_1246,N_1247,N_1248,N_1249,N_1250,N_1251,N_1252,N_1253,N_1254,N_1255,N_1256,N_1257,N_1258,N_1259,N_1260,N_1261,N_1262,N_1263,N_1264,N_1265,N_1266,N_1267,N_1268,N_1269,N_1270,N_1271,N_1272,N_1273,N_1274,N_1275,N_1276,N_1277,N_1278,N_1279,N_1280,N_1281,N_1282,N_1283,N_1284,N_1285,N_1286,N_1287,N_1288,N_1289,N_1290,N_1291,N_1292,N_1293,N_1294,N_1295,N_1296,N_1297,N_1298,N_1299,N_1300,N_1301,N_1302,N_1303,N_1304,N_1305,N_1306,N_1307,N_1308,N_1309,N_1310,N_1311,N_1312,N_1313,N_1314,N_1315,N_1316,N_1317,N_1318,N_1319,N_1320,N_1321,N_1322,N_1323,N_1324,N_1325,N_1326,N_1327,N_1328,N_1329,N_1330,N_1331,N_1332,N_1333,N_1334,N_1335,N_1336,N_1337,N_1338,N_1339,N_1340,N_1341,N_1342,N_1343,N_1344,N_1345,N_1346,N_1347,N_1348,N_1349,N_1350,N_1351,N_1352,N_1353,N_1354,N_1355,N_1356,N_1357,N_1358,N_1359,N_1360,N_1361,N_1362,N_1363,N_1364,N_1365,N_1366,N_1367,N_1368,N_1369,N_1370,N_1371,N_1372,N_1373,N_1374,N_1375,N_1376,N_1377,N_1378,N_1379,N_1380,N_1381,N_1382,N_1383,N_1384,N_1385,N_1386,N_1387,N_1388,N_1389,N_1390,N_1391,N_1392,N_1393,N_1394,N_1395,N_1396,N_1397,N_1398,N_1399,N_1400,N_1401,N_1402,N_1403,N_1404,N_1405,N_1406,N_1407,N_1408,N_1409,N_1410,N_1411,N_1412,N_1413,N_1414,N_1415,N_1416,N_1417,N_1418,N_1419,N_1420,N_1421,N_1422,N_1423,N_1424,N_1425,N_1426,N_1427,N_1428,N_1429,N_1430,N_1431,N_1432,N_1433,N_1434,N_1435,N_1436,N_1437,N_1438,N_1439,N_1440,N_1441,N_1442,N_1443,N_1444,N_1445,N_1446,N_1447,N_1448,N_1449,N_1450,N_1451,N_1452,N_1453,N_1454,N_1455,N_1456,N_1457,N_1458,N_1459,N_1460,N_1461,N_1462,N_1463,N_1464,N_1465,N_1466,N_1467,N_1468,N_1469,N_1470,N_1471,N_1472,N_1473,N_1474,N_1475,N_1476,N_1477,N_1478,N_1479,N_1480,N_1481,N_1482,N_1483,N_1484,N_1485,N_1486,N_1487,N_1488,N_1489,N_1490,N_1491,N_1492,N_1493,N_1494,N_1495,N_1496,N_1497,N_1498,N_1499,N_1500,N_1501,N_1502,N_1503,N_1504,N_1505,N_1506,N_1507,N_1508,N_1509,N_1510,N_1511,N_1512,N_1513,N_1514,N_1515,N_1516,N_1517,N_1518,N_1519,N_1520,N_1521,N_1522,N_1523,N_1524,N_1525,N_1526,N_1527,N_1528,N_1529,N_1530,N_1531,N_1532,N_1533,N_1534,N_1535,N_1536,N_1537,N_1538,N_1539,N_1540,N_1541,N_1542,N_1543,N_1544,N_1545,N_1546,N_1547,N_1548,N_1549,N_1550,N_1551,N_1552,N_1553,N_1554,N_1555,N_1556,N_1557,N_1558,N_1559,N_1560,N_1561,N_1562,N_1563,N_1564,N_1565,N_1566,N_1567,N_1568,N_1569,N_1570,N_1571,N_1572,N_1573,N_1574,N_1575,N_1576,N_1577,N_1578,N_1579,N_1580,N_1581,N_1582,N_1583,N_1584,N_1585,N_1586,N_1587,N_1588,N_1589,N_1590,N_1591,N_1592,N_1593,N_1594,N_1595,N_1596,N_1597,N_1598,N_1599,N_1600,N_1601,N_1602,N_1603,N_1604,N_1605,N_1606,N_1607,N_1608,N_1609,N_1610,N_1611,N_1612,N_1613,N_1614,N_1615,N_1616,N_1617,N_1618,N_1619,N_1620,N_1621,N_1622,N_1623,N_1624,N_1625,N_1626,N_1627,N_1628,N_1629,N_1630,N_1631,N_1632,N_1633,N_1634,N_1635,N_1636,N_1637,N_1638,N_1639,N_1640,N_1641,N_1642,N_1643,N_1644,N_1645,N_1646,N_1647,N_1648,N_1649,N_1650,N_1651,N_1652,N_1653,N_1654,N_1655,N_1656,N_1657,N_1658,N_1659,N_1660,N_1661,N_1662,N_1663,N_1664,N_1665,N_1666,N_1667,N_1668,N_1669,N_1670,N_1671,N_1672,N_1673,N_1674,N_1675,N_1676,N_1677,N_1678,N_1679,N_1680,N_1681,N_1682,N_1683,N_1684,N_1685,N_1686,N_1687,N_1688,N_1689,N_1690,N_1691,N_1692,N_1693,N_1694,N_1695,N_1696,N_1697,N_1698,N_1699,N_1700,N_1701,N_1702,N_1703,N_1704,N_1705,N_1706,N_1707,N_1708,N_1709,N_1710,N_1711,N_1712,N_1713,N_1714,N_1715,N_1716,N_1717,N_1718,N_1719,N_1720,N_1721,N_1722,N_1723,N_1724,N_1725,N_1726,N_1727,N_1728,N_1729,N_1730,N_1731,N_1732,N_1733,N_1734,N_1735,N_1736,N_1737,N_1738,N_1739,N_1740,N_1741,N_1742,N_1743,N_1744,N_1745,N_1746,N_1747,N_1748,N_1749,N_1750,N_1751,N_1752,N_1753,N_1754,N_1755,N_1756,N_1757,N_1758,N_1759,N_1760,N_1761,N_1762,N_1763,N_1764,N_1765,N_1766,N_1767,N_1768,N_1769,N_1770,N_1771,N_1772,N_1773,N_1774,N_1775,N_1776,N_1777,N_1778,N_1779,N_1780,N_1781,N_1782,N_1783,N_1784,N_1785,N_1786,N_1787,N_1788,N_1789,N_1790,N_1791,N_1792,N_1793,N_1794,N_1795,N_1796,N_1797,N_1798,N_1799,N_1800,N_1801,N_1802,N_1803,N_1804,N_1805,N_1806,N_1807,N_1808,N_1809,N_1810,N_1811,N_1812,N_1813,N_1814,N_1815,N_1816,N_1817,N_1818,N_1819,N_1820,N_1821,N_1822,N_1823,N_1824,N_1825,N_1826,N_1827,N_1828,N_1829,N_1830,N_1831,N_1832,N_1833,N_1834,N_1835,N_1836,N_1837,N_1838,N_1839,N_1840,N_1841,N_1842,N_1843,N_1844,N_1845,N_1846,N_1847,N_1848,N_1849,N_1850,N_1851,N_1852,N_1853,N_1854,N_1855,N_1856,N_1857,N_1858,N_1859,N_1860,N_1861,N_1862,N_1863,N_1864,N_1865,N_1866,N_1867,N_1868,N_1869,N_1870,N_1871,N_1872,N_1873,N_1874,N_1875,N_1876,N_1877,N_1878,N_1879,N_1880,N_1881,N_1882,N_1883,N_1884,N_1885,N_1886,N_1887,N_1888,N_1889,N_1890,N_1891,N_1892,N_1893,N_1894,N_1895,N_1896,N_1897,N_1898,N_1899,N_1900,N_1901,N_1902,N_1903,N_1904,N_1905,N_1906,N_1907,N_1908,N_1909,N_1910,N_1911,N_1912,N_1913,N_1914,N_1915,N_1916,N_1917,N_1918,N_1919,N_1920,N_1921,N_1922,N_1923,N_1924,N_1925,N_1926,N_1927,N_1928,N_1929,N_1930,N_1931,N_1932,N_1933,N_1934,N_1935,N_1936,N_1937,N_1938,N_1939,N_1940,N_1941,N_1942,N_1943,N_1944,N_1945,N_1946,N_1947,N_1948,N_1949,N_1950,N_1951,N_1952,N_1953,N_1954,N_1955,N_1956,N_1957,N_1958,N_1959,N_1960,N_1961,N_1962,N_1963,N_1964,N_1965,N_1966,N_1967,N_1968,N_1969,N_1970,N_1971,N_1972,N_1973,N_1974,N_1975,N_1976,N_1977,N_1978,N_1979,N_1980,N_1981,N_1982,N_1983,N_1984,N_1985,N_1986,N_1987,N_1988,N_1989,N_1990,N_1991,N_1992,N_1993,N_1994,N_1995,N_1996,N_1997,N_1998,N_1999,N_2000,N_2001,N_2002,N_2003,N_2004,N_2005,N_2006,N_2007,N_2008,N_2009,N_2010,N_2011,N_2012,N_2013,N_2014,N_2015,N_2016,N_2017,N_2018,N_2019,N_2020,N_2021,N_2022,N_2023,N_2024,N_2025,N_2026,N_2027,N_2028,N_2029,N_2030,N_2031,N_2032,N_2033,N_2034,N_2035,N_2036,N_2037,N_2038,N_2039,N_2040,N_2041,N_2042,N_2043,N_2044,N_2045,N_2046,N_2047,N_2048,N_2049,N_2050,N_2051,N_2052,N_2053,N_2054,N_2055,N_2056,N_2057,N_2058,N_2059,N_2060,N_2061,N_2062,N_2063,N_2064,N_2065,N_2066,N_2067,N_2068,N_2069,N_2070,N_2071,N_2072,N_2073,N_2074,N_2075,N_2076,N_2077,N_2078,N_2079,N_2080,N_2081,N_2082,N_2083,N_2084,N_2085,N_2086,N_2087,N_2088,N_2089,N_2090,N_2091,N_2092,N_2093,N_2094,N_2095,N_2096,N_2097,N_2098,N_2099,N_2100,N_2101,N_2102,N_2103,N_2104,N_2105,N_2106,N_2107,N_2108,N_2109,N_2110,N_2111,N_2112,N_2113,N_2114,N_2115,N_2116,N_2117,N_2118,N_2119,N_2120,N_2121,N_2122,N_2123,N_2124,N_2125,N_2126,N_2127,N_2128,N_2129,N_2130,N_2131,N_2132,N_2133,N_2134,N_2135,N_2136,N_2137,N_2138,N_2139,N_2140,N_2141,N_2142,N_2143,N_2144,N_2145,N_2146,N_2147,N_2148,N_2149,N_2150,N_2151,N_2152,N_2153,N_2154,N_2155,N_2156,N_2157,N_2158,N_2159,N_2160,N_2161,N_2162,N_2163,N_2164,N_2165,N_2166,N_2167,N_2168,N_2169,N_2170,N_2171,N_2172,N_2173,N_2174,N_2175,N_2176,N_2177,N_2178,N_2179,N_2180,N_2181,N_2182,N_2183,N_2184,N_2185,N_2186,N_2187,N_2188,N_2189,N_2190,N_2191,N_2192,N_2193,N_2194,N_2195,N_2196,N_2197,N_2198,N_2199,N_2200,N_2201,N_2202,N_2203,N_2204,N_2205,N_2206,N_2207,N_2208,N_2209,N_2210,N_2211,N_2212,N_2213,N_2214,N_2215,N_2216,N_2217,N_2218,N_2219,N_2220,N_2221,N_2222,N_2223,N_2224,N_2225,N_2226,N_2227,N_2228,N_2229,N_2230,N_2231,N_2232,N_2233,N_2234,N_2235,N_2236,N_2237,N_2238,N_2239,N_2240,N_2241,N_2242,N_2243,N_2244,N_2245,N_2246,N_2247,N_2248,N_2249,N_2250,N_2251,N_2252,N_2253,N_2254,N_2255,N_2256,N_2257,N_2258,N_2259,N_2260,N_2261,N_2262,N_2263,N_2264,N_2265,N_2266,N_2267,N_2268,N_2269,N_2270,N_2271,N_2272,N_2273,N_2274,N_2275,N_2276,N_2277,N_2278,N_2279,N_2280,N_2281,N_2282,N_2283,N_2284,N_2285,N_2286,N_2287,N_2288,N_2289,N_2290,N_2291,N_2292,N_2293,N_2294,N_2295,N_2296,N_2297,N_2298,N_2299,N_2300,N_2301,N_2302,N_2303,N_2304,N_2305,N_2306,N_2307,N_2308,N_2309,N_2310,N_2311,N_2312,N_2313,N_2314,N_2315,N_2316,N_2317,N_2318,N_2319,N_2320,N_2321,N_2322,N_2323,N_2324,N_2325,N_2326,N_2327,N_2328,N_2329,N_2330,N_2331,N_2332,N_2333,N_2334,N_2335,N_2336,N_2337,N_2338,N_2339,N_2340,N_2341,N_2342,N_2343,N_2344,N_2345,N_2346,N_2347,N_2348,N_2349,N_2350,N_2351,N_2352,N_2353,N_2354,N_2355,N_2356,N_2357,N_2358,N_2359,N_2360,N_2361,N_2362,N_2363,N_2364,N_2365,N_2366,N_2367,N_2368,N_2369,N_2370,N_2371,N_2372,N_2373,N_2374,N_2375,N_2376,N_2377,N_2378,N_2379,N_2380,N_2381,N_2382,N_2383,N_2384,N_2385,N_2386,N_2387,N_2388,N_2389,N_2390,N_2391,N_2392,N_2393,N_2394,N_2395,N_2396,N_2397,N_2398,N_2399,N_2400,N_2401,N_2402,N_2403,N_2404,N_2405,N_2406,N_2407,N_2408,N_2409,N_2410,N_2411,N_2412,N_2413,N_2414,N_2415,N_2416,N_2417,N_2418,N_2419,N_2420,N_2421,N_2422,N_2423,N_2424,N_2425,N_2426,N_2427,N_2428,N_2429,N_2430,N_2431,N_2432,N_2433,N_2434,N_2435,N_2436,N_2437,N_2438,N_2439,N_2440,N_2441,N_2442,N_2443,N_2444,N_2445,N_2446,N_2447,N_2448,N_2449,N_2450,N_2451,N_2452,N_2453,N_2454,N_2455,N_2456,N_2457,N_2458,N_2459,N_2460,N_2461,N_2462,N_2463,N_2464,N_2465,N_2466,N_2467,N_2468,N_2469,N_2470,N_2471,N_2472,N_2473,N_2474,N_2475,N_2476,N_2477,N_2478,N_2479,N_2480,N_2481,N_2482,N_2483,N_2484,N_2485,N_2486,N_2487,N_2488,N_2489,N_2490,N_2491,N_2492,N_2493,N_2494,N_2495,N_2496,N_2497,N_2498,N_2499,N_2500,N_2501,N_2502,N_2503,N_2504,N_2505,N_2506,N_2507,N_2508,N_2509,N_2510,N_2511,N_2512,N_2513,N_2514,N_2515,N_2516,N_2517,N_2518,N_2519,N_2520,N_2521,N_2522,N_2523,N_2524,N_2525,N_2526,N_2527,N_2528,N_2529,N_2530,N_2531,N_2532,N_2533,N_2534,N_2535,N_2536,N_2537,N_2538,N_2539,N_2540,N_2541,N_2542,N_2543,N_2544,N_2545,N_2546,N_2547,N_2548,N_2549,N_2550,N_2551,N_2552,N_2553,N_2554,N_2555,N_2556,N_2557,N_2558,N_2559,N_2560,N_2561,N_2562,N_2563,N_2564,N_2565,N_2566,N_2567,N_2568,N_2569,N_2570,N_2571,N_2572,N_2573,N_2574,N_2575,N_2576,N_2577,N_2578,N_2579,N_2580,N_2581,N_2582,N_2583,N_2584,N_2585,N_2586,N_2587,N_2588,N_2589,N_2590,N_2591,N_2592,N_2593,N_2594,N_2595,N_2596,N_2597,N_2598,N_2599,N_2600,N_2601,N_2602,N_2603,N_2604,N_2605,N_2606,N_2607,N_2608,N_2609,N_2610,N_2611,N_2612,N_2613,N_2614,N_2615,N_2616,N_2617,N_2618,N_2619,N_2620,N_2621,N_2622,N_2623,N_2624,N_2625,N_2626,N_2627,N_2628,N_2629,N_2630,N_2631,N_2632,N_2633,N_2634,N_2635,N_2636,N_2637,N_2638,N_2639,N_2640,N_2641,N_2642,N_2643,N_2644,N_2645,N_2646,N_2647,N_2648,N_2649,N_2650,N_2651,N_2652,N_2653,N_2654,N_2655,N_2656,N_2657,N_2658,N_2659,N_2660,N_2661,N_2662,N_2663,N_2664,N_2665,N_2666,N_2667,N_2668,N_2669,N_2670,N_2671,N_2672,N_2673,N_2674,N_2675,N_2676,N_2677,N_2678,N_2679,N_2680,N_2681,N_2682,N_2683,N_2684,N_2685,N_2686,N_2687,N_2688,N_2689,N_2690,N_2691,N_2692,N_2693,N_2694,N_2695,N_2696,N_2697,N_2698,N_2699,N_2700,N_2701,N_2702,N_2703,N_2704,N_2705,N_2706,N_2707,N_2708,N_2709,N_2710,N_2711,N_2712,N_2713,N_2714,N_2715,N_2716,N_2717,N_2718,N_2719,N_2720,N_2721,N_2722,N_2723,N_2724,N_2725,N_2726,N_2727,N_2728,N_2729,N_2730,N_2731,N_2732,N_2733,N_2734,N_2735,N_2736,N_2737,N_2738,N_2739,N_2740,N_2741,N_2742,N_2743,N_2744,N_2745,N_2746,N_2747,N_2748,N_2749,N_2750,N_2751,N_2752,N_2753,N_2754,N_2755,N_2756,N_2757,N_2758,N_2759,N_2760,N_2761,N_2762,N_2763,N_2764,N_2765,N_2766,N_2767,N_2768,N_2769,N_2770,N_2771,N_2772,N_2773,N_2774,N_2775,N_2776,N_2777,N_2778,N_2779,N_2780,N_2781,N_2782,N_2783,N_2784,N_2785,N_2786,N_2787,N_2788,N_2789,N_2790,N_2791,N_2792,N_2793,N_2794,N_2795,N_2796,N_2797,N_2798,N_2799,N_2800,N_2801,N_2802,N_2803,N_2804,N_2805,N_2806,N_2807,N_2808,N_2809,N_2810,N_2811,N_2812,N_2813,N_2814,N_2815,N_2816,N_2817,N_2818,N_2819,N_2820,N_2821,N_2822,N_2823,N_2824,N_2825,N_2826,N_2827,N_2828,N_2829,N_2830,N_2831,N_2832,N_2833,N_2834,N_2835,N_2836,N_2837,N_2838,N_2839,N_2840,N_2841,N_2842,N_2843,N_2844,N_2845,N_2846,N_2847,N_2848,N_2849,N_2850,N_2851,N_2852,N_2853,N_2854,N_2855,N_2856,N_2857,N_2858,N_2859,N_2860,N_2861,N_2862,N_2863,N_2864,N_2865,N_2866,N_2867,N_2868,N_2869,N_2870,N_2871,N_2872,N_2873,N_2874,N_2875,N_2876,N_2877,N_2878,N_2879,N_2880,N_2881,N_2882,N_2883,N_2884,N_2885,N_2886,N_2887,N_2888,N_2889,N_2890,N_2891,N_2892,N_2893,N_2894,N_2895,N_2896,N_2897,N_2898,N_2899,N_2900,N_2901,N_2902,N_2903,N_2904,N_2905,N_2906,N_2907,N_2908,N_2909,N_2910,N_2911,N_2912,N_2913,N_2914,N_2915,N_2916,N_2917,N_2918,N_2919,N_2920,N_2921,N_2922,N_2923,N_2924,N_2925,N_2926,N_2927,N_2928,N_2929,N_2930,N_2931,N_2932,N_2933,N_2934,N_2935,N_2936,N_2937,N_2938,N_2939,N_2940,N_2941,N_2942,N_2943,N_2944,N_2945,N_2946,N_2947,N_2948,N_2949,N_2950,N_2951,N_2952,N_2953,N_2954,N_2955,N_2956,N_2957,N_2958,N_2959,N_2960,N_2961,N_2962,N_2963,N_2964,N_2965,N_2966,N_2967,N_2968,N_2969,N_2970,N_2971,N_2972,N_2973,N_2974,N_2975,N_2976,N_2977,N_2978,N_2979,N_2980,N_2981,N_2982,N_2983,N_2984,N_2985,N_2986,N_2987,N_2988,N_2989,N_2990,N_2991,N_2992,N_2993,N_2994,N_2995,N_2996,N_2997,N_2998,N_2999,N_3000,N_3001,N_3002,N_3003,N_3004,N_3005,N_3006,N_3007,N_3008,N_3009,N_3010,N_3011,N_3012,N_3013,N_3014,N_3015,N_3016,N_3017,N_3018,N_3019,N_3020,N_3021,N_3022,N_3023,N_3024,N_3025,N_3026,N_3027,N_3028,N_3029,N_3030,N_3031,N_3032,N_3033,N_3034,N_3035,N_3036,N_3037,N_3038,N_3039,N_3040,N_3041,N_3042,N_3043,N_3044,N_3045,N_3046,N_3047,N_3048,N_3049,N_3050,N_3051,N_3052,N_3053,N_3054,N_3055,N_3056,N_3057,N_3058,N_3059,N_3060,N_3061,N_3062,N_3063,N_3064,N_3065,N_3066,N_3067,N_3068,N_3069,N_3070,N_3071,N_3072,N_3073,N_3074,N_3075,N_3076,N_3077,N_3078,N_3079,N_3080,N_3081,N_3082,N_3083,N_3084,N_3085,N_3086,N_3087,N_3088,N_3089,N_3090,N_3091,N_3092,N_3093,N_3094,N_3095,N_3096,N_3097,N_3098,N_3099,N_3100,N_3101,N_3102,N_3103,N_3104,N_3105,N_3106,N_3107,N_3108,N_3109,N_3110,N_3111,N_3112,N_3113,N_3114,N_3115,N_3116,N_3117,N_3118,N_3119,N_3120,N_3121,N_3122,N_3123,N_3124,N_3125,N_3126,N_3127,N_3128,N_3129,N_3130,N_3131,N_3132,N_3133,N_3134,N_3135,N_3136,N_3137,N_3138,N_3139,N_3140,N_3141,N_3142,N_3143,N_3144,N_3145,N_3146,N_3147,N_3148,N_3149,N_3150,N_3151,N_3152,N_3153,N_3154,N_3155,N_3156,N_3157,N_3158,N_3159,N_3160,N_3161,N_3162,N_3163,N_3164,N_3165,N_3166,N_3167,N_3168,N_3169,N_3170,N_3171,N_3172,N_3173,N_3174,N_3175,N_3176,N_3177,N_3178,N_3179,N_3180,N_3181,N_3182,N_3183,N_3184,N_3185,N_3186,N_3187,N_3188,N_3189,N_3190,N_3191,N_3192,N_3193,N_3194,N_3195,N_3196,N_3197,N_3198,N_3199,N_3200,N_3201,N_3202,N_3203,N_3204,N_3205,N_3206,N_3207,N_3208,N_3209,N_3210,N_3211,N_3212,N_3213,N_3214,N_3215,N_3216,N_3217,N_3218,N_3219,N_3220,N_3221,N_3222,N_3223,N_3224,N_3225,N_3226,N_3227,N_3228,N_3229,N_3230,N_3231,N_3232,N_3233,N_3234,N_3235,N_3236,N_3237,N_3238,N_3239,N_3240,N_3241,N_3242,N_3243,N_3244,N_3245,N_3246,N_3247,N_3248,N_3249,N_3250,N_3251,N_3252,N_3253,N_3254,N_3255,N_3256,N_3257,N_3258,N_3259,N_3260,N_3261,N_3262,N_3263,N_3264,N_3265,N_3266,N_3267,N_3268,N_3269,N_3270,N_3271,N_3272,N_3273,N_3274,N_3275,N_3276,N_3277,N_3278,N_3279,N_3280,N_3281,N_3282,N_3283,N_3284,N_3285,N_3286,N_3287,N_3288,N_3289,N_3290,N_3291,N_3292,N_3293,N_3294,N_3295,N_3296,N_3297,N_3298,N_3299,N_3300,N_3301,N_3302,N_3303,N_3304,N_3305,N_3306,N_3307,N_3308,N_3309,N_3310,N_3311,N_3312,N_3313,N_3314,N_3315,N_3316,N_3317,N_3318,N_3319,N_3320,N_3321,N_3322,N_3323,N_3324,N_3325,N_3326,N_3327,N_3328,N_3329,N_3330,N_3331,N_3332,N_3333,N_3334,N_3335,N_3336,N_3337,N_3338,N_3339,N_3340,N_3341,N_3342,N_3343,N_3344,N_3345,N_3346,N_3347,N_3348,N_3349,N_3350,N_3351,N_3352,N_3353,N_3354,N_3355,N_3356,N_3357,N_3358,N_3359,N_3360,N_3361,N_3362,N_3363,N_3364,N_3365,N_3366,N_3367,N_3368,N_3369,N_3370,N_3371,N_3372,N_3373,N_3374,N_3375,N_3376,N_3377,N_3378,N_3379,N_3380,N_3381,N_3382,N_3383,N_3384,N_3385,N_3386,N_3387,N_3388,N_3389,N_3390,N_3391,N_3392,N_3393,N_3394,N_3395,N_3396,N_3397,N_3398,N_3399,N_3400,N_3401,N_3402,N_3403,N_3404,N_3405,N_3406,N_3407,N_3408,N_3409,N_3410,N_3411,N_3412,N_3413,N_3414,N_3415,N_3416,N_3417,N_3418,N_3419,N_3420,N_3421,N_3422,N_3423,N_3424,N_3425,N_3426,N_3427,N_3428,N_3429,N_3430,N_3431,N_3432,N_3433,N_3434,N_3435,N_3436,N_3437,N_3438,N_3439,N_3440,N_3441,N_3442,N_3443,N_3444,N_3445,N_3446,N_3447,N_3448,N_3449,N_3450,N_3451,N_3452,N_3453,N_3454,N_3455,N_3456,N_3457,N_3458,N_3459,N_3460,N_3461,N_3462,N_3463,N_3464,N_3465,N_3466,N_3467,N_3468,N_3469,N_3470,N_3471,N_3472,N_3473,N_3474,N_3475,N_3476,N_3477,N_3478,N_3479,N_3480,N_3481,N_3482,N_3483,N_3484,N_3485,N_3486,N_3487,N_3488,N_3489,N_3490,N_3491,N_3492,N_3493,N_3494,N_3495,N_3496,N_3497,N_3498,N_3499,N_3500,N_3501,N_3502,N_3503,N_3504,N_3505,N_3506,N_3507,N_3508,N_3509,N_3510,N_3511,N_3512,N_3513,N_3514,N_3515,N_3516,N_3517,N_3518,N_3519,N_3520,N_3521,N_3522,N_3523,N_3524,N_3525,N_3526,N_3527,N_3528,N_3529,N_3530,N_3531,N_3532,N_3533,N_3534,N_3535,N_3536,N_3537,N_3538,N_3539,N_3540,N_3541,N_3542,N_3543,N_3544,N_3545,N_3546,N_3547,N_3548,N_3549,N_3550,N_3551,N_3552,N_3553,N_3554,N_3555,N_3556,N_3557,N_3558,N_3559,N_3560,N_3561,N_3562,N_3563,N_3564,N_3565,N_3566,N_3567,N_3568,N_3569,N_3570,N_3571,N_3572,N_3573,N_3574,N_3575,N_3576,N_3577,N_3578,N_3579,N_3580,N_3581,N_3582,N_3583,N_3584,N_3585,N_3586,N_3587,N_3588,N_3589,N_3590,N_3591,N_3592,N_3593,N_3594,N_3595,N_3596,N_3597,N_3598,N_3599,N_3600,N_3601,N_3602,N_3603,N_3604,N_3605,N_3606,N_3607,N_3608,N_3609,N_3610,N_3611,N_3612,N_3613,N_3614,N_3615,N_3616,N_3617,N_3618,N_3619,N_3620,N_3621,N_3622,N_3623,N_3624,N_3625,N_3626,N_3627,N_3628,N_3629,N_3630,N_3631,N_3632,N_3633,N_3634,N_3635,N_3636,N_3637,N_3638,N_3639,N_3640,N_3641,N_3642,N_3643,N_3644,N_3645,N_3646,N_3647,N_3648,N_3649,N_3650,N_3651,N_3652,N_3653,N_3654,N_3655,N_3656,N_3657,N_3658,N_3659,N_3660,N_3661,N_3662,N_3663,N_3664,N_3665,N_3666,N_3667,N_3668,N_3669,N_3670,N_3671,N_3672,N_3673,N_3674,N_3675,N_3676,N_3677,N_3678,N_3679,N_3680,N_3681,N_3682,N_3683,N_3684,N_3685,N_3686,N_3687,N_3688,N_3689,N_3690,N_3691,N_3692,N_3693,N_3694,N_3695,N_3696,N_3697,N_3698,N_3699,N_3700,N_3701,N_3702,N_3703,N_3704,N_3705,N_3706,N_3707,N_3708,N_3709,N_3710,N_3711,N_3712,N_3713,N_3714,N_3715,N_3716,N_3717,N_3718,N_3719,N_3720,N_3721,N_3722,N_3723,N_3724,N_3725,N_3726,N_3727,N_3728,N_3729,N_3730,N_3731,N_3732,N_3733,N_3734,N_3735,N_3736,N_3737,N_3738,N_3739,N_3740,N_3741,N_3742,N_3743,N_3744,N_3745,N_3746,N_3747,N_3748,N_3749,N_3750,N_3751,N_3752,N_3753,N_3754,N_3755,N_3756,N_3757,N_3758,N_3759,N_3760,N_3761,N_3762,N_3763,N_3764,N_3765,N_3766,N_3767,N_3768,N_3769,N_3770,N_3771,N_3772,N_3773,N_3774,N_3775,N_3776,N_3777,N_3778,N_3779,N_3780,N_3781,N_3782,N_3783,N_3784,N_3785,N_3786,N_3787,N_3788,N_3789,N_3790,N_3791,N_3792,N_3793,N_3794,N_3795,N_3796,N_3797,N_3798,N_3799,N_3800,N_3801,N_3802,N_3803,N_3804,N_3805,N_3806,N_3807,N_3808,N_3809,N_3810,N_3811,N_3812,N_3813,N_3814,N_3815,N_3816,N_3817,N_3818,N_3819,N_3820,N_3821,N_3822,N_3823,N_3824,N_3825,N_3826,N_3827,N_3828,N_3829,N_3830,N_3831,N_3832,N_3833,N_3834,N_3835,N_3836,N_3837,N_3838,N_3839,N_3840,N_3841,N_3842,N_3843,N_3844,N_3845,N_3846,N_3847,N_3848,N_3849,N_3850,N_3851,N_3852,N_3853,N_3854,N_3855,N_3856,N_3857,N_3858,N_3859,N_3860,N_3861,N_3862,N_3863,N_3864,N_3865,N_3866,N_3867,N_3868,N_3869,N_3870,N_3871,N_3872,N_3873,N_3874,N_3875,N_3876,N_3877,N_3878,N_3879,N_3880,N_3881,N_3882,N_3883,N_3884,N_3885,N_3886,N_3887,N_3888,N_3889,N_3890,N_3891,N_3892,N_3893,N_3894,N_3895,N_3896,N_3897,N_3898,N_3899,N_3900,N_3901,N_3902,N_3903,N_3904,N_3905,N_3906,N_3907,N_3908,N_3909,N_3910,N_3911,N_3912,N_3913,N_3914,N_3915,N_3916,N_3917,N_3918,N_3919,N_3920,N_3921,N_3922,N_3923,N_3924,N_3925,N_3926,N_3927,N_3928,N_3929,N_3930,N_3931,N_3932,N_3933,N_3934,N_3935,N_3936,N_3937,N_3938,N_3939,N_3940,N_3941,N_3942,N_3943,N_3944,N_3945,N_3946,N_3947,N_3948,N_3949,N_3950,N_3951,N_3952,N_3953,N_3954,N_3955,N_3956,N_3957,N_3958,N_3959,N_3960,N_3961,N_3962,N_3963,N_3964,N_3965,N_3966,N_3967,N_3968,N_3969,N_3970,N_3971,N_3972,N_3973,N_3974,N_3975,N_3976,N_3977,N_3978,N_3979,N_3980,N_3981,N_3982,N_3983,N_3984,N_3985,N_3986,N_3987,N_3988,N_3989,N_3990,N_3991,N_3992,N_3993,N_3994,N_3995,N_3996,N_3997,N_3998,N_3999,N_4000,N_4001,N_4002,N_4003,N_4004,N_4005,N_4006,N_4007,N_4008,N_4009,N_4010,N_4011,N_4012,N_4013,N_4014,N_4015,N_4016,N_4017,N_4018,N_4019,N_4020,N_4021,N_4022,N_4023,N_4024,N_4025,N_4026,N_4027,N_4028,N_4029,N_4030,N_4031,N_4032,N_4033,N_4034,N_4035,N_4036,N_4037,N_4038,N_4039,N_4040,N_4041,N_4042,N_4043,N_4044,N_4045,N_4046,N_4047,N_4048,N_4049,N_4050,N_4051,N_4052,N_4053,N_4054,N_4055,N_4056,N_4057,N_4058,N_4059,N_4060,N_4061,N_4062,N_4063,N_4064,N_4065,N_4066,N_4067,N_4068,N_4069,N_4070,N_4071,N_4072,N_4073,N_4074,N_4075,N_4076,N_4077,N_4078,N_4079,N_4080,N_4081,N_4082,N_4083,N_4084,N_4085,N_4086,N_4087,N_4088,N_4089,N_4090,N_4091,N_4092,N_4093,N_4094,N_4095,N_4096,N_4097,N_4098,N_4099,N_4100,N_4101,N_4102,N_4103,N_4104,N_4105,N_4106,N_4107,N_4108,N_4109,N_4110,N_4111,N_4112,N_4113,N_4114,N_4115,N_4116,N_4117,N_4118,N_4119,N_4120,N_4121,N_4122,N_4123,N_4124,N_4125,N_4126,N_4127,N_4128,N_4129,N_4130,N_4131,N_4132,N_4133,N_4134,N_4135,N_4136,N_4137,N_4138,N_4139,N_4140,N_4141,N_4142,N_4143,N_4144,N_4145,N_4146,N_4147,N_4148,N_4149,N_4150,N_4151,N_4152,N_4153,N_4154,N_4155,N_4156,N_4157,N_4158,N_4159,N_4160,N_4161,N_4162,N_4163,N_4164,N_4165,N_4166,N_4167,N_4168,N_4169,N_4170,N_4171,N_4172,N_4173,N_4174,N_4175,N_4176,N_4177,N_4178,N_4179,N_4180,N_4181,N_4182,N_4183,N_4184,N_4185,N_4186,N_4187,N_4188,N_4189,N_4190,N_4191,N_4192,N_4193,N_4194,N_4195,N_4196,N_4197,N_4198,N_4199,N_4200,N_4201,N_4202,N_4203,N_4204,N_4205,N_4206,N_4207,N_4208,N_4209,N_4210,N_4211,N_4212,N_4213,N_4214,N_4215,N_4216,N_4217,N_4218,N_4219,N_4220,N_4221,N_4222,N_4223,N_4224,N_4225,N_4226,N_4227,N_4228,N_4229,N_4230,N_4231,N_4232,N_4233,N_4234,N_4235,N_4236,N_4237,N_4238,N_4239,N_4240,N_4241,N_4242,N_4243,N_4244,N_4245,N_4246,N_4247,N_4248,N_4249,N_4250,N_4251,N_4252,N_4253,N_4254,N_4255,N_4256,N_4257,N_4258,N_4259,N_4260,N_4261,N_4262,N_4263,N_4264,N_4265,N_4266,N_4267,N_4268,N_4269,N_4270,N_4271,N_4272,N_4273,N_4274,N_4275,N_4276,N_4277,N_4278,N_4279,N_4280,N_4281,N_4282,N_4283,N_4284,N_4285,N_4286,N_4287,N_4288,N_4289,N_4290,N_4291,N_4292,N_4293,N_4294,N_4295,N_4296,N_4297,N_4298,N_4299,N_4300,N_4301,N_4302,N_4303,N_4304,N_4305,N_4306,N_4307,N_4308,N_4309,N_4310,N_4311,N_4312,N_4313,N_4314,N_4315,N_4316,N_4317,N_4318,N_4319,N_4320,N_4321,N_4322,N_4323,N_4324,N_4325,N_4326,N_4327,N_4328,N_4329,N_4330,N_4331,N_4332,N_4333,N_4334,N_4335,N_4336,N_4337,N_4338,N_4339,N_4340,N_4341,N_4342,N_4343,N_4344,N_4345,N_4346,N_4347,N_4348,N_4349,N_4350,N_4351,N_4352,N_4353,N_4354,N_4355,N_4356,N_4357,N_4358,N_4359,N_4360,N_4361,N_4362,N_4363,N_4364,N_4365,N_4366,N_4367,N_4368,N_4369,N_4370,N_4371,N_4372,N_4373,N_4374,N_4375,N_4376,N_4377,N_4378,N_4379,N_4380,N_4381,N_4382,N_4383,N_4384,N_4385,N_4386,N_4387,N_4388,N_4389,N_4390,N_4391,N_4392,N_4393,N_4394,N_4395,N_4396,N_4397,N_4398,N_4399,N_4400,N_4401,N_4402,N_4403,N_4404,N_4405,N_4406,N_4407,N_4408,N_4409,N_4410,N_4411,N_4412,N_4413,N_4414,N_4415,N_4416,N_4417,N_4418,N_4419,N_4420,N_4421,N_4422,N_4423,N_4424,N_4425,N_4426,N_4427,N_4428,N_4429,N_4430,N_4431,N_4432,N_4433,N_4434,N_4435,N_4436,N_4437,N_4438,N_4439,N_4440,N_4441,N_4442,N_4443,N_4444,N_4445,N_4446,N_4447,N_4448,N_4449,N_4450,N_4451,N_4452,N_4453,N_4454,N_4455,N_4456,N_4457,N_4458,N_4459,N_4460,N_4461,N_4462,N_4463,N_4464,N_4465,N_4466,N_4467,N_4468,N_4469,N_4470,N_4471,N_4472,N_4473,N_4474,N_4475,N_4476,N_4477,N_4478,N_4479,N_4480,N_4481,N_4482,N_4483,N_4484,N_4485,N_4486,N_4487,N_4488,N_4489,N_4490,N_4491,N_4492,N_4493,N_4494,N_4495,N_4496,N_4497,N_4498,N_4499,N_4500,N_4501,N_4502,N_4503,N_4504,N_4505,N_4506,N_4507,N_4508,N_4509,N_4510,N_4511,N_4512,N_4513,N_4514,N_4515,N_4516,N_4517,N_4518,N_4519,N_4520,N_4521,N_4522,N_4523,N_4524,N_4525,N_4526,N_4527,N_4528,N_4529,N_4530,N_4531,N_4532,N_4533,N_4534,N_4535,N_4536,N_4537,N_4538,N_4539,N_4540,N_4541,N_4542,N_4543,N_4544,N_4545,N_4546,N_4547,N_4548,N_4549,N_4550,N_4551,N_4552,N_4553,N_4554,N_4555,N_4556,N_4557,N_4558,N_4559,N_4560,N_4561,N_4562,N_4563,N_4564,N_4565,N_4566,N_4567,N_4568,N_4569,N_4570,N_4571,N_4572,N_4573,N_4574,N_4575,N_4576,N_4577,N_4578,N_4579,N_4580,N_4581,N_4582,N_4583,N_4584,N_4585,N_4586,N_4587,N_4588,N_4589,N_4590,N_4591,N_4592,N_4593,N_4594,N_4595,N_4596,N_4597,N_4598,N_4599,N_4600,N_4601,N_4602,N_4603,N_4604,N_4605,N_4606,N_4607,N_4608,N_4609,N_4610,N_4611,N_4612,N_4613,N_4614,N_4615,N_4616,N_4617,N_4618,N_4619,N_4620,N_4621,N_4622,N_4623,N_4624,N_4625,N_4626,N_4627,N_4628,N_4629,N_4630,N_4631,N_4632,N_4633,N_4634,N_4635,N_4636,N_4637,N_4638,N_4639,N_4640,N_4641,N_4642,N_4643,N_4644,N_4645,N_4646,N_4647,N_4648,N_4649,N_4650,N_4651,N_4652,N_4653,N_4654,N_4655,N_4656,N_4657,N_4658,N_4659,N_4660,N_4661,N_4662,N_4663,N_4664,N_4665,N_4666,N_4667,N_4668,N_4669,N_4670,N_4671,N_4672,N_4673,N_4674,N_4675,N_4676,N_4677,N_4678,N_4679,N_4680,N_4681,N_4682,N_4683,N_4684,N_4685,N_4686,N_4687,N_4688,N_4689,N_4690,N_4691,N_4692,N_4693,N_4694,N_4695,N_4696,N_4697,N_4698,N_4699,N_4700,N_4701,N_4702,N_4703,N_4704,N_4705,N_4706,N_4707,N_4708,N_4709,N_4710,N_4711,N_4712,N_4713,N_4714,N_4715,N_4716,N_4717,N_4718,N_4719,N_4720,N_4721,N_4722,N_4723,N_4724,N_4725,N_4726,N_4727,N_4728,N_4729,N_4730,N_4731,N_4732,N_4733,N_4734,N_4735,N_4736,N_4737,N_4738,N_4739,N_4740,N_4741,N_4742,N_4743,N_4744,N_4745,N_4746,N_4747,N_4748,N_4749,N_4750,N_4751,N_4752,N_4753,N_4754,N_4755,N_4756,N_4757,N_4758,N_4759,N_4760,N_4761,N_4762,N_4763,N_4764,N_4765,N_4766,N_4767,N_4768,N_4769,N_4770,N_4771,N_4772,N_4773,N_4774,N_4775,N_4776,N_4777,N_4778,N_4779,N_4780,N_4781,N_4782,N_4783,N_4784,N_4785,N_4786,N_4787,N_4788,N_4789,N_4790,N_4791,N_4792,N_4793,N_4794,N_4795,N_4796,N_4797,N_4798,N_4799,N_4800,N_4801,N_4802,N_4803,N_4804,N_4805,N_4806,N_4807,N_4808,N_4809,N_4810,N_4811,N_4812,N_4813,N_4814,N_4815,N_4816,N_4817,N_4818,N_4819,N_4820,N_4821,N_4822,N_4823,N_4824,N_4825,N_4826,N_4827,N_4828,N_4829,N_4830,N_4831,N_4832,N_4833,N_4834,N_4835,N_4836,N_4837,N_4838,N_4839,N_4840,N_4841,N_4842,N_4843,N_4844,N_4845,N_4846,N_4847,N_4848,N_4849,N_4850,N_4851,N_4852,N_4853,N_4854,N_4855,N_4856,N_4857,N_4858,N_4859,N_4860,N_4861,N_4862,N_4863,N_4864,N_4865,N_4866,N_4867,N_4868,N_4869,N_4870,N_4871,N_4872,N_4873,N_4874,N_4875,N_4876,N_4877,N_4878,N_4879,N_4880,N_4881,N_4882,N_4883,N_4884,N_4885,N_4886,N_4887,N_4888,N_4889,N_4890,N_4891,N_4892,N_4893,N_4894,N_4895,N_4896,N_4897,N_4898,N_4899,N_4900,N_4901,N_4902,N_4903,N_4904,N_4905,N_4906,N_4907,N_4908,N_4909,N_4910,N_4911,N_4912,N_4913,N_4914,N_4915,N_4916,N_4917,N_4918,N_4919,N_4920,N_4921,N_4922,N_4923,N_4924,N_4925,N_4926,N_4927,N_4928,N_4929,N_4930,N_4931,N_4932,N_4933,N_4934,N_4935,N_4936,N_4937,N_4938,N_4939,N_4940,N_4941,N_4942,N_4943,N_4944,N_4945,N_4946,N_4947,N_4948,N_4949,N_4950,N_4951,N_4952,N_4953,N_4954,N_4955,N_4956,N_4957,N_4958,N_4959,N_4960,N_4961,N_4962,N_4963,N_4964,N_4965,N_4966,N_4967,N_4968,N_4969,N_4970,N_4971,N_4972,N_4973,N_4974,N_4975,N_4976,N_4977,N_4978,N_4979,N_4980,N_4981,N_4982,N_4983,N_4984,N_4985,N_4986,N_4987,N_4988,N_4989,N_4990,N_4991,N_4992,N_4993,N_4994,N_4995,N_4996,N_4997,N_4998,N_4999;
nand U0 (N_0,In_404,In_119);
nand U1 (N_1,In_695,In_371);
and U2 (N_2,In_48,In_659);
nand U3 (N_3,In_718,In_338);
nand U4 (N_4,In_256,In_378);
and U5 (N_5,In_152,In_442);
nand U6 (N_6,In_42,In_239);
nor U7 (N_7,In_41,In_12);
nor U8 (N_8,In_612,In_386);
nand U9 (N_9,In_545,In_615);
and U10 (N_10,In_490,In_45);
and U11 (N_11,In_308,In_491);
nor U12 (N_12,In_356,In_577);
or U13 (N_13,In_295,In_637);
or U14 (N_14,In_484,In_209);
and U15 (N_15,In_475,In_705);
and U16 (N_16,In_403,In_473);
or U17 (N_17,In_266,In_498);
nor U18 (N_18,In_642,In_696);
and U19 (N_19,In_14,In_325);
nand U20 (N_20,In_599,In_517);
nand U21 (N_21,In_293,In_16);
nand U22 (N_22,In_644,In_390);
or U23 (N_23,In_125,In_106);
xnor U24 (N_24,In_175,In_296);
nand U25 (N_25,In_510,In_117);
and U26 (N_26,In_465,In_204);
and U27 (N_27,In_508,In_749);
xnor U28 (N_28,In_206,In_722);
and U29 (N_29,In_529,In_99);
and U30 (N_30,In_76,In_411);
nand U31 (N_31,In_425,In_421);
nand U32 (N_32,In_747,In_423);
or U33 (N_33,In_246,In_51);
and U34 (N_34,In_302,In_536);
or U35 (N_35,In_522,In_310);
nor U36 (N_36,In_441,In_156);
nand U37 (N_37,In_252,In_200);
nor U38 (N_38,In_518,In_623);
or U39 (N_39,In_133,In_8);
nor U40 (N_40,In_311,In_512);
or U41 (N_41,In_461,In_19);
nand U42 (N_42,In_242,In_668);
and U43 (N_43,In_625,In_214);
or U44 (N_44,In_714,In_579);
nor U45 (N_45,In_107,In_726);
nor U46 (N_46,In_346,In_559);
or U47 (N_47,In_576,In_80);
and U48 (N_48,In_306,In_552);
nor U49 (N_49,In_56,In_660);
nor U50 (N_50,In_343,In_147);
nand U51 (N_51,In_5,In_217);
or U52 (N_52,In_740,In_263);
nand U53 (N_53,In_710,In_700);
or U54 (N_54,In_173,In_572);
nor U55 (N_55,In_192,In_128);
nand U56 (N_56,In_741,In_22);
xor U57 (N_57,In_514,In_245);
or U58 (N_58,In_591,In_13);
nand U59 (N_59,In_21,In_701);
nor U60 (N_60,In_163,In_391);
or U61 (N_61,In_291,In_419);
nand U62 (N_62,In_331,In_614);
nor U63 (N_63,In_400,In_113);
and U64 (N_64,In_342,In_20);
or U65 (N_65,In_432,In_344);
nand U66 (N_66,In_410,In_730);
nand U67 (N_67,In_723,In_176);
xnor U68 (N_68,In_732,In_187);
nor U69 (N_69,In_566,In_622);
or U70 (N_70,In_375,In_538);
or U71 (N_71,In_497,In_160);
nand U72 (N_72,In_715,In_406);
or U73 (N_73,In_127,In_57);
and U74 (N_74,In_408,In_624);
xor U75 (N_75,In_583,In_549);
xor U76 (N_76,In_570,In_348);
nor U77 (N_77,In_321,In_554);
or U78 (N_78,In_645,In_329);
nor U79 (N_79,In_9,In_435);
nand U80 (N_80,In_458,In_731);
nor U81 (N_81,In_420,In_301);
and U82 (N_82,In_560,In_505);
nor U83 (N_83,In_126,In_516);
and U84 (N_84,In_692,In_401);
and U85 (N_85,In_352,In_673);
nor U86 (N_86,In_734,In_537);
or U87 (N_87,In_221,In_687);
nor U88 (N_88,In_628,In_480);
nor U89 (N_89,In_184,In_122);
nor U90 (N_90,In_597,In_459);
nand U91 (N_91,In_494,In_65);
xor U92 (N_92,In_743,In_72);
nand U93 (N_93,In_626,In_121);
and U94 (N_94,In_150,In_259);
or U95 (N_95,In_728,In_273);
nor U96 (N_96,In_651,In_678);
nor U97 (N_97,In_100,In_546);
or U98 (N_98,In_499,In_573);
and U99 (N_99,In_229,In_190);
nand U100 (N_100,In_304,In_215);
xnor U101 (N_101,In_608,In_0);
and U102 (N_102,In_662,In_611);
or U103 (N_103,In_361,In_153);
nor U104 (N_104,In_527,In_297);
and U105 (N_105,In_254,In_157);
nand U106 (N_106,In_95,In_643);
xor U107 (N_107,In_519,In_558);
nor U108 (N_108,In_481,In_196);
and U109 (N_109,In_275,In_370);
nand U110 (N_110,In_82,In_682);
nor U111 (N_111,In_253,In_46);
and U112 (N_112,In_380,In_36);
nor U113 (N_113,In_564,In_300);
or U114 (N_114,In_198,In_716);
and U115 (N_115,In_276,In_199);
nor U116 (N_116,In_328,In_681);
and U117 (N_117,In_711,In_418);
nand U118 (N_118,In_249,In_413);
nand U119 (N_119,In_650,In_75);
xor U120 (N_120,In_197,In_142);
xor U121 (N_121,In_446,In_648);
nand U122 (N_122,In_78,In_399);
xnor U123 (N_123,In_208,In_213);
nor U124 (N_124,In_470,In_108);
nand U125 (N_125,In_81,In_621);
and U126 (N_126,In_704,In_424);
nor U127 (N_127,In_541,In_71);
nor U128 (N_128,In_589,In_504);
nand U129 (N_129,In_52,In_129);
and U130 (N_130,In_220,In_55);
and U131 (N_131,In_212,In_294);
xor U132 (N_132,In_193,In_454);
and U133 (N_133,In_702,In_202);
nand U134 (N_134,In_151,In_658);
nand U135 (N_135,In_556,In_70);
and U136 (N_136,In_647,In_224);
and U137 (N_137,In_154,In_322);
nand U138 (N_138,In_664,In_670);
or U139 (N_139,In_136,In_268);
nand U140 (N_140,In_267,In_675);
nor U141 (N_141,In_733,In_496);
or U142 (N_142,In_571,In_60);
nand U143 (N_143,In_610,In_737);
or U144 (N_144,In_284,In_607);
or U145 (N_145,In_677,In_241);
xor U146 (N_146,In_557,In_90);
or U147 (N_147,In_178,In_289);
nor U148 (N_148,In_563,In_398);
and U149 (N_149,In_205,In_86);
nor U150 (N_150,In_639,In_143);
nand U151 (N_151,In_238,In_598);
nand U152 (N_152,In_587,In_627);
or U153 (N_153,In_500,In_416);
nor U154 (N_154,In_62,In_316);
nor U155 (N_155,In_636,In_319);
nor U156 (N_156,In_307,In_233);
or U157 (N_157,In_596,In_164);
nor U158 (N_158,In_685,In_111);
nand U159 (N_159,In_616,In_464);
and U160 (N_160,In_593,In_148);
nor U161 (N_161,In_66,In_713);
nor U162 (N_162,In_326,In_368);
and U163 (N_163,In_472,In_92);
nor U164 (N_164,In_739,In_439);
or U165 (N_165,In_544,In_271);
or U166 (N_166,In_35,In_54);
nand U167 (N_167,In_260,In_699);
nand U168 (N_168,In_582,In_34);
nand U169 (N_169,In_149,In_452);
nor U170 (N_170,In_580,In_28);
nor U171 (N_171,In_394,In_262);
nand U172 (N_172,In_466,In_449);
xor U173 (N_173,In_186,In_179);
xor U174 (N_174,In_110,In_671);
and U175 (N_175,In_323,In_447);
nor U176 (N_176,In_376,In_548);
nor U177 (N_177,In_96,In_94);
or U178 (N_178,In_305,In_689);
nor U179 (N_179,In_58,In_59);
nor U180 (N_180,In_502,In_524);
nand U181 (N_181,In_247,In_520);
nor U182 (N_182,In_283,In_482);
nand U183 (N_183,In_725,In_155);
or U184 (N_184,In_287,In_535);
nor U185 (N_185,In_140,In_542);
and U186 (N_186,In_364,In_47);
or U187 (N_187,In_511,In_18);
or U188 (N_188,In_298,In_703);
or U189 (N_189,In_594,In_303);
and U190 (N_190,In_476,In_456);
nand U191 (N_191,In_333,In_581);
xor U192 (N_192,In_357,In_444);
or U193 (N_193,In_632,In_738);
nor U194 (N_194,In_667,In_431);
nand U195 (N_195,In_477,In_64);
and U196 (N_196,In_350,In_382);
nor U197 (N_197,In_201,In_251);
or U198 (N_198,In_244,In_162);
nand U199 (N_199,In_281,In_341);
and U200 (N_200,In_161,In_29);
and U201 (N_201,N_117,In_219);
and U202 (N_202,N_33,N_136);
and U203 (N_203,In_114,In_426);
nand U204 (N_204,In_440,N_130);
and U205 (N_205,N_61,In_25);
nor U206 (N_206,N_143,N_75);
nand U207 (N_207,N_42,In_513);
nand U208 (N_208,N_29,In_226);
nor U209 (N_209,N_178,In_609);
nand U210 (N_210,N_139,N_46);
nor U211 (N_211,N_19,N_10);
nor U212 (N_212,In_132,N_3);
or U213 (N_213,In_592,In_724);
nor U214 (N_214,N_170,In_665);
nand U215 (N_215,In_455,In_676);
xnor U216 (N_216,N_127,N_25);
and U217 (N_217,In_102,N_104);
nor U218 (N_218,In_169,N_173);
nand U219 (N_219,N_191,In_601);
or U220 (N_220,In_130,N_39);
nor U221 (N_221,In_116,In_124);
and U222 (N_222,In_474,In_77);
nor U223 (N_223,In_457,N_106);
nor U224 (N_224,N_159,In_282);
or U225 (N_225,In_415,N_135);
nand U226 (N_226,N_148,In_274);
and U227 (N_227,In_232,In_417);
and U228 (N_228,In_746,In_506);
nand U229 (N_229,In_377,N_193);
or U230 (N_230,In_223,N_121);
or U231 (N_231,N_20,In_84);
nand U232 (N_232,In_347,N_35);
or U233 (N_233,In_721,N_160);
and U234 (N_234,N_52,N_197);
nand U235 (N_235,In_652,In_278);
and U236 (N_236,N_198,In_412);
nand U237 (N_237,N_95,In_586);
xnor U238 (N_238,In_655,In_359);
nand U239 (N_239,In_141,In_392);
and U240 (N_240,In_686,In_37);
nor U241 (N_241,In_83,In_684);
and U242 (N_242,In_26,N_80);
and U243 (N_243,In_744,In_222);
nand U244 (N_244,N_141,In_286);
or U245 (N_245,N_70,In_174);
xnor U246 (N_246,In_332,In_430);
nor U247 (N_247,N_112,In_98);
nand U248 (N_248,N_140,In_330);
nand U249 (N_249,In_706,In_460);
nor U250 (N_250,In_363,In_30);
nand U251 (N_251,In_27,In_654);
nand U252 (N_252,In_495,In_194);
xnor U253 (N_253,N_100,N_67);
nand U254 (N_254,In_534,In_50);
nand U255 (N_255,In_729,In_409);
or U256 (N_256,N_120,N_122);
or U257 (N_257,In_89,N_172);
and U258 (N_258,N_71,In_33);
nand U259 (N_259,N_50,N_167);
and U260 (N_260,In_688,In_397);
or U261 (N_261,N_142,In_354);
and U262 (N_262,In_467,N_62);
nand U263 (N_263,In_462,In_468);
nor U264 (N_264,N_161,In_367);
or U265 (N_265,In_620,In_379);
nand U266 (N_266,N_175,N_74);
and U267 (N_267,In_146,In_340);
nor U268 (N_268,N_64,In_280);
nor U269 (N_269,In_335,In_451);
or U270 (N_270,In_641,In_39);
nor U271 (N_271,In_189,In_666);
or U272 (N_272,In_10,In_619);
nand U273 (N_273,In_530,In_235);
and U274 (N_274,In_182,N_81);
xor U275 (N_275,In_653,In_145);
nor U276 (N_276,N_181,In_49);
nand U277 (N_277,In_317,N_152);
and U278 (N_278,In_483,N_154);
nor U279 (N_279,N_156,In_68);
nand U280 (N_280,In_74,In_736);
xnor U281 (N_281,In_427,In_1);
and U282 (N_282,In_180,In_595);
nor U283 (N_283,In_661,In_159);
nand U284 (N_284,N_47,In_588);
and U285 (N_285,In_93,In_237);
xnor U286 (N_286,In_345,In_369);
nand U287 (N_287,N_72,N_88);
nor U288 (N_288,In_567,N_94);
nand U289 (N_289,In_463,In_191);
or U290 (N_290,N_65,N_79);
nor U291 (N_291,N_18,N_15);
xor U292 (N_292,In_657,N_133);
and U293 (N_293,In_562,In_312);
nor U294 (N_294,In_188,In_231);
xnor U295 (N_295,In_603,In_374);
nand U296 (N_296,N_128,In_584);
and U297 (N_297,In_358,N_83);
nand U298 (N_298,N_1,N_180);
or U299 (N_299,In_634,In_469);
nor U300 (N_300,N_158,In_38);
or U301 (N_301,In_503,In_745);
and U302 (N_302,N_92,N_189);
nand U303 (N_303,In_314,In_373);
xnor U304 (N_304,In_486,N_49);
or U305 (N_305,N_90,In_15);
xor U306 (N_306,In_574,In_539);
nand U307 (N_307,In_485,In_488);
and U308 (N_308,In_438,N_6);
and U309 (N_309,N_125,N_108);
nor U310 (N_310,N_27,N_165);
or U311 (N_311,In_327,In_309);
nor U312 (N_312,In_227,N_145);
nor U313 (N_313,In_509,In_261);
nor U314 (N_314,In_674,N_169);
xor U315 (N_315,In_167,In_450);
nand U316 (N_316,N_138,N_194);
nor U317 (N_317,In_493,In_393);
nor U318 (N_318,In_550,N_37);
or U319 (N_319,In_324,In_523);
and U320 (N_320,In_631,N_183);
nor U321 (N_321,In_396,N_51);
and U322 (N_322,In_288,In_349);
nor U323 (N_323,N_56,N_171);
xor U324 (N_324,In_735,In_228);
nand U325 (N_325,In_384,In_139);
or U326 (N_326,In_613,In_69);
or U327 (N_327,In_585,In_203);
nor U328 (N_328,In_561,In_181);
and U329 (N_329,N_182,In_183);
or U330 (N_330,N_119,In_590);
nand U331 (N_331,In_719,In_366);
nor U332 (N_332,N_114,In_445);
and U333 (N_333,In_690,N_4);
nand U334 (N_334,N_91,N_76);
and U335 (N_335,In_315,N_9);
nor U336 (N_336,In_551,In_656);
and U337 (N_337,N_54,In_540);
nand U338 (N_338,In_604,In_120);
and U339 (N_339,In_569,N_28);
and U340 (N_340,N_69,N_101);
nand U341 (N_341,N_21,In_712);
nor U342 (N_342,N_123,In_547);
or U343 (N_343,In_137,N_45);
or U344 (N_344,N_103,N_164);
xnor U345 (N_345,In_158,In_478);
or U346 (N_346,In_680,In_104);
nand U347 (N_347,In_693,N_17);
nand U348 (N_348,In_24,In_337);
and U349 (N_349,N_150,N_5);
nand U350 (N_350,In_362,In_290);
or U351 (N_351,N_34,N_111);
xor U352 (N_352,N_134,N_110);
or U353 (N_353,In_600,In_171);
and U354 (N_354,In_679,In_334);
or U355 (N_355,In_115,In_748);
xnor U356 (N_356,N_187,In_568);
or U357 (N_357,N_146,In_230);
or U358 (N_358,In_543,N_84);
nor U359 (N_359,In_53,In_525);
and U360 (N_360,In_265,N_2);
and U361 (N_361,N_11,In_85);
or U362 (N_362,In_389,N_137);
and U363 (N_363,N_31,N_0);
and U364 (N_364,In_299,N_144);
and U365 (N_365,N_55,In_553);
and U366 (N_366,N_77,In_105);
and U367 (N_367,In_618,In_727);
xor U368 (N_368,In_318,In_663);
or U369 (N_369,In_313,N_68);
nand U370 (N_370,N_53,N_30);
nor U371 (N_371,In_433,In_669);
or U372 (N_372,N_132,In_207);
nand U373 (N_373,In_177,In_694);
and U374 (N_374,In_292,In_138);
nand U375 (N_375,N_43,In_531);
nand U376 (N_376,N_157,In_32);
or U377 (N_377,In_507,N_151);
nand U378 (N_378,In_2,In_672);
nand U379 (N_379,In_23,N_177);
and U380 (N_380,N_40,In_277);
nand U381 (N_381,In_118,In_355);
and U382 (N_382,In_258,In_489);
and U383 (N_383,In_240,In_381);
nand U384 (N_384,In_285,In_492);
or U385 (N_385,In_629,N_162);
and U386 (N_386,N_115,N_107);
nor U387 (N_387,N_85,In_388);
nand U388 (N_388,In_646,N_8);
or U389 (N_389,N_66,In_63);
nor U390 (N_390,In_195,In_43);
and U391 (N_391,N_168,In_234);
nor U392 (N_392,N_176,In_257);
or U393 (N_393,In_135,N_60);
and U394 (N_394,In_360,In_269);
and U395 (N_395,N_24,In_387);
and U396 (N_396,In_4,In_40);
and U397 (N_397,N_26,In_339);
nand U398 (N_398,In_31,In_172);
nand U399 (N_399,In_720,In_270);
nor U400 (N_400,In_336,In_521);
or U401 (N_401,N_342,N_240);
nand U402 (N_402,In_395,N_208);
nand U403 (N_403,N_383,N_298);
and U404 (N_404,N_364,N_212);
xor U405 (N_405,N_291,In_635);
or U406 (N_406,In_533,N_371);
nor U407 (N_407,N_294,N_301);
nor U408 (N_408,In_264,N_41);
xor U409 (N_409,In_3,In_638);
and U410 (N_410,In_279,In_555);
nand U411 (N_411,N_231,N_210);
and U412 (N_412,In_73,In_640);
nand U413 (N_413,N_186,N_378);
nand U414 (N_414,In_255,N_201);
nor U415 (N_415,N_327,N_217);
nor U416 (N_416,In_44,N_385);
or U417 (N_417,N_174,In_372);
nand U418 (N_418,N_259,N_129);
and U419 (N_419,N_220,N_360);
and U420 (N_420,In_365,In_7);
nor U421 (N_421,In_248,N_63);
or U422 (N_422,N_243,In_414);
or U423 (N_423,N_23,N_376);
nand U424 (N_424,N_296,N_306);
xor U425 (N_425,N_275,In_170);
nor U426 (N_426,In_131,In_6);
nor U427 (N_427,In_742,In_717);
xnor U428 (N_428,N_264,In_144);
nor U429 (N_429,N_184,In_606);
and U430 (N_430,N_323,N_219);
or U431 (N_431,N_254,N_375);
nor U432 (N_432,N_271,N_356);
nand U433 (N_433,N_384,N_325);
nor U434 (N_434,N_310,In_165);
nor U435 (N_435,N_199,In_87);
or U436 (N_436,In_605,N_227);
or U437 (N_437,N_206,N_293);
nor U438 (N_438,In_443,N_82);
xnor U439 (N_439,N_337,N_14);
and U440 (N_440,N_299,N_339);
xor U441 (N_441,N_302,N_250);
nor U442 (N_442,N_363,N_328);
or U443 (N_443,N_304,In_385);
nand U444 (N_444,N_347,In_407);
or U445 (N_445,In_383,In_422);
nor U446 (N_446,N_391,N_244);
nand U447 (N_447,N_247,N_93);
and U448 (N_448,N_362,N_257);
or U449 (N_449,N_292,In_218);
nor U450 (N_450,N_399,In_501);
nand U451 (N_451,N_367,N_48);
nand U452 (N_452,N_326,N_396);
nor U453 (N_453,N_333,N_276);
nand U454 (N_454,N_290,N_269);
or U455 (N_455,N_267,In_210);
xnor U456 (N_456,N_248,N_279);
and U457 (N_457,In_707,N_359);
nand U458 (N_458,N_256,In_97);
nor U459 (N_459,N_222,In_101);
or U460 (N_460,N_149,N_349);
and U461 (N_461,N_12,N_204);
or U462 (N_462,N_377,N_32);
xor U463 (N_463,N_345,In_602);
and U464 (N_464,N_379,N_246);
nor U465 (N_465,N_365,N_211);
and U466 (N_466,N_270,N_98);
or U467 (N_467,N_251,N_372);
nand U468 (N_468,N_331,In_109);
xor U469 (N_469,In_453,In_91);
and U470 (N_470,In_448,N_397);
xnor U471 (N_471,N_366,N_36);
or U472 (N_472,N_223,N_253);
and U473 (N_473,N_245,N_338);
and U474 (N_474,N_321,In_112);
nand U475 (N_475,N_288,N_131);
nor U476 (N_476,N_382,N_57);
nor U477 (N_477,In_532,N_370);
nor U478 (N_478,N_280,N_96);
or U479 (N_479,In_578,N_285);
or U480 (N_480,N_188,In_272);
nor U481 (N_481,N_307,N_312);
and U482 (N_482,N_265,In_428);
xor U483 (N_483,N_316,N_289);
or U484 (N_484,N_281,N_319);
nor U485 (N_485,N_209,In_633);
or U486 (N_486,N_228,N_16);
and U487 (N_487,N_303,N_87);
and U488 (N_488,N_58,In_526);
or U489 (N_489,N_357,N_118);
or U490 (N_490,In_709,In_17);
or U491 (N_491,N_155,N_387);
and U492 (N_492,N_215,In_402);
nor U493 (N_493,N_354,In_236);
and U494 (N_494,N_341,N_196);
and U495 (N_495,In_67,N_226);
nand U496 (N_496,N_22,N_7);
nor U497 (N_497,In_351,In_630);
nand U498 (N_498,In_185,N_386);
or U499 (N_499,N_113,N_236);
nand U500 (N_500,In_429,N_335);
nor U501 (N_501,N_230,N_221);
and U502 (N_502,In_528,N_268);
nor U503 (N_503,N_203,N_320);
or U504 (N_504,N_284,N_179);
nand U505 (N_505,N_258,N_214);
and U506 (N_506,N_238,N_13);
nand U507 (N_507,N_239,N_252);
or U508 (N_508,N_346,N_274);
nor U509 (N_509,N_340,N_334);
or U510 (N_510,N_353,N_205);
and U511 (N_511,N_234,N_314);
and U512 (N_512,N_324,N_330);
nand U513 (N_513,In_708,N_361);
nor U514 (N_514,N_305,In_434);
nand U515 (N_515,N_393,N_286);
or U516 (N_516,In_649,In_698);
nand U517 (N_517,N_398,N_235);
nor U518 (N_518,In_565,N_329);
and U519 (N_519,N_218,N_190);
nor U520 (N_520,N_105,In_575);
and U521 (N_521,N_355,N_380);
nor U522 (N_522,In_697,N_272);
nand U523 (N_523,In_134,N_86);
nor U524 (N_524,N_124,N_392);
nor U525 (N_525,N_263,N_224);
nand U526 (N_526,In_61,In_79);
or U527 (N_527,N_300,N_237);
or U528 (N_528,N_295,N_395);
or U529 (N_529,N_229,N_59);
and U530 (N_530,In_243,N_287);
and U531 (N_531,In_123,In_436);
or U532 (N_532,In_216,In_225);
and U533 (N_533,N_374,N_225);
and U534 (N_534,In_617,N_261);
nor U535 (N_535,N_381,N_233);
nor U536 (N_536,N_318,N_358);
and U537 (N_537,N_352,N_368);
nor U538 (N_538,N_311,N_200);
nor U539 (N_539,N_216,N_350);
or U540 (N_540,N_373,N_44);
nand U541 (N_541,N_277,In_487);
nor U542 (N_542,N_73,In_320);
or U543 (N_543,N_109,N_241);
and U544 (N_544,N_192,N_185);
nand U545 (N_545,In_515,N_343);
nand U546 (N_546,N_313,N_38);
nand U547 (N_547,N_389,N_332);
nand U548 (N_548,In_250,N_394);
nor U549 (N_549,N_163,N_89);
nand U550 (N_550,N_232,In_437);
and U551 (N_551,In_683,In_11);
and U552 (N_552,N_390,N_166);
nand U553 (N_553,In_103,N_213);
nor U554 (N_554,In_479,N_242);
nor U555 (N_555,N_278,N_351);
nand U556 (N_556,In_166,N_116);
xnor U557 (N_557,N_207,N_348);
or U558 (N_558,N_336,In_405);
or U559 (N_559,N_322,N_309);
nand U560 (N_560,N_102,N_317);
nand U561 (N_561,N_260,N_266);
and U562 (N_562,N_78,In_691);
xor U563 (N_563,N_282,In_471);
nor U564 (N_564,N_97,In_168);
nor U565 (N_565,In_88,N_388);
and U566 (N_566,In_211,N_297);
or U567 (N_567,N_344,N_255);
or U568 (N_568,N_315,N_153);
nand U569 (N_569,N_369,N_249);
and U570 (N_570,N_262,N_202);
nand U571 (N_571,N_283,N_126);
nand U572 (N_572,N_99,N_308);
nor U573 (N_573,N_195,N_147);
or U574 (N_574,In_353,N_273);
nor U575 (N_575,N_399,N_184);
nor U576 (N_576,N_131,In_707);
nor U577 (N_577,N_377,In_630);
and U578 (N_578,N_320,N_383);
nand U579 (N_579,N_12,N_244);
or U580 (N_580,N_319,N_109);
or U581 (N_581,In_395,N_223);
and U582 (N_582,N_380,In_210);
nand U583 (N_583,In_528,N_355);
nor U584 (N_584,N_250,N_337);
xor U585 (N_585,N_363,N_59);
or U586 (N_586,N_233,N_82);
or U587 (N_587,In_17,N_329);
nand U588 (N_588,In_185,N_319);
or U589 (N_589,In_649,N_318);
nand U590 (N_590,N_311,N_44);
and U591 (N_591,N_381,In_264);
nand U592 (N_592,N_186,N_153);
or U593 (N_593,In_405,N_99);
xor U594 (N_594,N_340,N_381);
or U595 (N_595,N_113,N_89);
nand U596 (N_596,In_336,In_385);
xnor U597 (N_597,N_264,In_709);
and U598 (N_598,N_235,In_443);
xor U599 (N_599,N_270,N_299);
nor U600 (N_600,N_474,N_568);
or U601 (N_601,N_437,N_489);
nand U602 (N_602,N_405,N_435);
nor U603 (N_603,N_540,N_422);
xnor U604 (N_604,N_480,N_456);
nor U605 (N_605,N_570,N_493);
and U606 (N_606,N_484,N_502);
and U607 (N_607,N_460,N_504);
nor U608 (N_608,N_400,N_584);
nor U609 (N_609,N_466,N_598);
and U610 (N_610,N_458,N_461);
xnor U611 (N_611,N_587,N_416);
or U612 (N_612,N_462,N_589);
or U613 (N_613,N_535,N_527);
nand U614 (N_614,N_557,N_438);
and U615 (N_615,N_574,N_546);
nand U616 (N_616,N_430,N_596);
nand U617 (N_617,N_436,N_449);
and U618 (N_618,N_478,N_455);
or U619 (N_619,N_401,N_464);
or U620 (N_620,N_520,N_408);
and U621 (N_621,N_521,N_550);
xor U622 (N_622,N_450,N_413);
or U623 (N_623,N_441,N_439);
xor U624 (N_624,N_554,N_403);
nand U625 (N_625,N_523,N_530);
nor U626 (N_626,N_560,N_440);
and U627 (N_627,N_476,N_531);
or U628 (N_628,N_431,N_423);
or U629 (N_629,N_417,N_591);
nor U630 (N_630,N_513,N_432);
or U631 (N_631,N_418,N_515);
nor U632 (N_632,N_517,N_500);
xor U633 (N_633,N_522,N_412);
or U634 (N_634,N_507,N_564);
or U635 (N_635,N_511,N_424);
xor U636 (N_636,N_414,N_445);
nor U637 (N_637,N_410,N_468);
and U638 (N_638,N_573,N_490);
nor U639 (N_639,N_539,N_516);
or U640 (N_640,N_506,N_497);
xnor U641 (N_641,N_576,N_544);
and U642 (N_642,N_491,N_448);
or U643 (N_643,N_471,N_433);
nand U644 (N_644,N_538,N_402);
or U645 (N_645,N_404,N_585);
and U646 (N_646,N_518,N_525);
and U647 (N_647,N_465,N_529);
or U648 (N_648,N_426,N_453);
or U649 (N_649,N_483,N_467);
and U650 (N_650,N_588,N_503);
and U651 (N_651,N_498,N_572);
nand U652 (N_652,N_566,N_512);
or U653 (N_653,N_590,N_556);
nor U654 (N_654,N_519,N_594);
nand U655 (N_655,N_469,N_543);
or U656 (N_656,N_475,N_429);
and U657 (N_657,N_494,N_434);
xor U658 (N_658,N_420,N_597);
nand U659 (N_659,N_411,N_581);
nand U660 (N_660,N_537,N_495);
nand U661 (N_661,N_562,N_472);
nand U662 (N_662,N_508,N_463);
or U663 (N_663,N_419,N_509);
nor U664 (N_664,N_485,N_533);
or U665 (N_665,N_447,N_510);
and U666 (N_666,N_446,N_470);
or U667 (N_667,N_580,N_586);
or U668 (N_668,N_486,N_571);
or U669 (N_669,N_595,N_593);
nor U670 (N_670,N_553,N_555);
nand U671 (N_671,N_496,N_451);
or U672 (N_672,N_549,N_532);
nor U673 (N_673,N_427,N_407);
nor U674 (N_674,N_536,N_599);
and U675 (N_675,N_514,N_421);
and U676 (N_676,N_583,N_579);
nor U677 (N_677,N_524,N_487);
nor U678 (N_678,N_561,N_488);
nor U679 (N_679,N_552,N_457);
nand U680 (N_680,N_409,N_459);
or U681 (N_681,N_545,N_541);
nor U682 (N_682,N_428,N_425);
nand U683 (N_683,N_559,N_526);
and U684 (N_684,N_443,N_548);
xnor U685 (N_685,N_501,N_577);
nand U686 (N_686,N_477,N_567);
or U687 (N_687,N_563,N_452);
and U688 (N_688,N_444,N_505);
and U689 (N_689,N_473,N_499);
nor U690 (N_690,N_415,N_406);
nand U691 (N_691,N_558,N_592);
and U692 (N_692,N_578,N_479);
or U693 (N_693,N_582,N_547);
or U694 (N_694,N_442,N_528);
nor U695 (N_695,N_534,N_492);
or U696 (N_696,N_482,N_542);
nor U697 (N_697,N_575,N_569);
nor U698 (N_698,N_481,N_551);
and U699 (N_699,N_565,N_454);
nor U700 (N_700,N_514,N_442);
and U701 (N_701,N_592,N_514);
nor U702 (N_702,N_448,N_461);
and U703 (N_703,N_499,N_433);
nand U704 (N_704,N_507,N_517);
and U705 (N_705,N_480,N_580);
nand U706 (N_706,N_459,N_497);
or U707 (N_707,N_548,N_421);
xnor U708 (N_708,N_597,N_587);
nand U709 (N_709,N_598,N_552);
nor U710 (N_710,N_532,N_469);
and U711 (N_711,N_558,N_501);
or U712 (N_712,N_589,N_405);
nor U713 (N_713,N_545,N_457);
nand U714 (N_714,N_472,N_492);
or U715 (N_715,N_524,N_569);
and U716 (N_716,N_411,N_549);
or U717 (N_717,N_598,N_537);
nand U718 (N_718,N_475,N_588);
nor U719 (N_719,N_467,N_577);
xor U720 (N_720,N_424,N_419);
nand U721 (N_721,N_546,N_499);
nor U722 (N_722,N_420,N_594);
nand U723 (N_723,N_457,N_548);
xor U724 (N_724,N_599,N_587);
nor U725 (N_725,N_512,N_430);
nor U726 (N_726,N_575,N_586);
nand U727 (N_727,N_482,N_461);
nand U728 (N_728,N_597,N_562);
xnor U729 (N_729,N_426,N_476);
or U730 (N_730,N_473,N_428);
and U731 (N_731,N_480,N_499);
nand U732 (N_732,N_513,N_476);
nand U733 (N_733,N_474,N_453);
nand U734 (N_734,N_468,N_558);
nor U735 (N_735,N_483,N_577);
nor U736 (N_736,N_497,N_493);
nand U737 (N_737,N_571,N_566);
or U738 (N_738,N_436,N_469);
and U739 (N_739,N_483,N_443);
nand U740 (N_740,N_547,N_541);
xnor U741 (N_741,N_419,N_463);
nand U742 (N_742,N_577,N_416);
nor U743 (N_743,N_484,N_480);
and U744 (N_744,N_576,N_599);
or U745 (N_745,N_582,N_548);
and U746 (N_746,N_478,N_491);
and U747 (N_747,N_503,N_487);
or U748 (N_748,N_445,N_566);
nor U749 (N_749,N_592,N_459);
and U750 (N_750,N_469,N_552);
and U751 (N_751,N_592,N_443);
nand U752 (N_752,N_488,N_431);
or U753 (N_753,N_503,N_510);
xor U754 (N_754,N_587,N_424);
nand U755 (N_755,N_538,N_489);
or U756 (N_756,N_560,N_546);
nor U757 (N_757,N_457,N_427);
nor U758 (N_758,N_537,N_430);
or U759 (N_759,N_412,N_568);
and U760 (N_760,N_583,N_496);
nor U761 (N_761,N_437,N_411);
nand U762 (N_762,N_571,N_534);
nand U763 (N_763,N_513,N_410);
or U764 (N_764,N_581,N_478);
xor U765 (N_765,N_481,N_572);
and U766 (N_766,N_592,N_480);
or U767 (N_767,N_528,N_491);
and U768 (N_768,N_401,N_517);
nand U769 (N_769,N_445,N_576);
nand U770 (N_770,N_588,N_577);
nand U771 (N_771,N_551,N_512);
or U772 (N_772,N_523,N_505);
nor U773 (N_773,N_481,N_537);
nor U774 (N_774,N_500,N_564);
nor U775 (N_775,N_473,N_412);
nand U776 (N_776,N_503,N_522);
nor U777 (N_777,N_445,N_536);
nand U778 (N_778,N_422,N_487);
nand U779 (N_779,N_495,N_486);
or U780 (N_780,N_573,N_494);
nand U781 (N_781,N_558,N_464);
nor U782 (N_782,N_459,N_580);
or U783 (N_783,N_457,N_405);
or U784 (N_784,N_491,N_416);
and U785 (N_785,N_427,N_499);
nor U786 (N_786,N_488,N_407);
and U787 (N_787,N_405,N_429);
nor U788 (N_788,N_500,N_575);
nor U789 (N_789,N_565,N_471);
nor U790 (N_790,N_567,N_429);
nor U791 (N_791,N_447,N_456);
nor U792 (N_792,N_554,N_409);
nand U793 (N_793,N_489,N_584);
or U794 (N_794,N_582,N_468);
nor U795 (N_795,N_536,N_541);
nor U796 (N_796,N_475,N_519);
nand U797 (N_797,N_441,N_531);
nor U798 (N_798,N_437,N_520);
and U799 (N_799,N_422,N_464);
nand U800 (N_800,N_772,N_797);
or U801 (N_801,N_662,N_608);
xor U802 (N_802,N_759,N_735);
nor U803 (N_803,N_773,N_784);
nor U804 (N_804,N_730,N_721);
or U805 (N_805,N_648,N_639);
nor U806 (N_806,N_746,N_619);
or U807 (N_807,N_668,N_650);
or U808 (N_808,N_767,N_656);
and U809 (N_809,N_638,N_641);
nor U810 (N_810,N_686,N_763);
and U811 (N_811,N_622,N_676);
and U812 (N_812,N_614,N_713);
nor U813 (N_813,N_742,N_647);
xnor U814 (N_814,N_745,N_754);
nand U815 (N_815,N_760,N_620);
or U816 (N_816,N_634,N_645);
and U817 (N_817,N_642,N_774);
or U818 (N_818,N_690,N_611);
and U819 (N_819,N_621,N_702);
nand U820 (N_820,N_604,N_744);
and U821 (N_821,N_785,N_798);
nor U822 (N_822,N_661,N_795);
or U823 (N_823,N_728,N_709);
or U824 (N_824,N_779,N_740);
nand U825 (N_825,N_717,N_739);
or U826 (N_826,N_758,N_617);
nand U827 (N_827,N_747,N_749);
nand U828 (N_828,N_794,N_799);
nor U829 (N_829,N_724,N_697);
or U830 (N_830,N_601,N_748);
or U831 (N_831,N_653,N_729);
and U832 (N_832,N_658,N_751);
and U833 (N_833,N_616,N_663);
nand U834 (N_834,N_607,N_694);
nand U835 (N_835,N_723,N_714);
or U836 (N_836,N_768,N_726);
nor U837 (N_837,N_640,N_788);
nor U838 (N_838,N_674,N_673);
nand U839 (N_839,N_600,N_737);
nand U840 (N_840,N_769,N_793);
xor U841 (N_841,N_612,N_770);
and U842 (N_842,N_693,N_623);
nand U843 (N_843,N_630,N_776);
or U844 (N_844,N_766,N_734);
nor U845 (N_845,N_757,N_701);
nand U846 (N_846,N_711,N_736);
nor U847 (N_847,N_722,N_603);
nor U848 (N_848,N_627,N_672);
nor U849 (N_849,N_626,N_660);
or U850 (N_850,N_646,N_664);
and U851 (N_851,N_696,N_685);
and U852 (N_852,N_665,N_613);
or U853 (N_853,N_609,N_698);
or U854 (N_854,N_637,N_657);
nand U855 (N_855,N_689,N_781);
or U856 (N_856,N_715,N_688);
and U857 (N_857,N_692,N_705);
or U858 (N_858,N_700,N_629);
or U859 (N_859,N_606,N_738);
nor U860 (N_860,N_753,N_750);
xor U861 (N_861,N_624,N_786);
nand U862 (N_862,N_643,N_687);
nor U863 (N_863,N_778,N_743);
nand U864 (N_864,N_655,N_752);
or U865 (N_865,N_659,N_682);
and U866 (N_866,N_681,N_755);
xor U867 (N_867,N_602,N_695);
xnor U868 (N_868,N_679,N_710);
or U869 (N_869,N_651,N_771);
nor U870 (N_870,N_732,N_678);
nand U871 (N_871,N_741,N_733);
nor U872 (N_872,N_712,N_762);
and U873 (N_873,N_725,N_765);
xor U874 (N_874,N_605,N_691);
xnor U875 (N_875,N_628,N_731);
nor U876 (N_876,N_718,N_764);
or U877 (N_877,N_756,N_666);
or U878 (N_878,N_610,N_792);
nor U879 (N_879,N_652,N_633);
or U880 (N_880,N_654,N_706);
and U881 (N_881,N_684,N_707);
nand U882 (N_882,N_703,N_675);
and U883 (N_883,N_631,N_677);
xor U884 (N_884,N_720,N_669);
nor U885 (N_885,N_775,N_683);
or U886 (N_886,N_680,N_615);
or U887 (N_887,N_649,N_716);
and U888 (N_888,N_704,N_708);
or U889 (N_889,N_644,N_632);
nor U890 (N_890,N_783,N_777);
and U891 (N_891,N_761,N_670);
and U892 (N_892,N_790,N_780);
and U893 (N_893,N_618,N_782);
or U894 (N_894,N_671,N_719);
xnor U895 (N_895,N_787,N_636);
nand U896 (N_896,N_791,N_635);
or U897 (N_897,N_796,N_699);
or U898 (N_898,N_625,N_727);
and U899 (N_899,N_667,N_789);
and U900 (N_900,N_747,N_726);
and U901 (N_901,N_638,N_745);
nand U902 (N_902,N_613,N_796);
and U903 (N_903,N_658,N_770);
or U904 (N_904,N_690,N_667);
and U905 (N_905,N_763,N_717);
and U906 (N_906,N_764,N_646);
or U907 (N_907,N_663,N_676);
nor U908 (N_908,N_771,N_627);
or U909 (N_909,N_715,N_738);
xnor U910 (N_910,N_683,N_744);
xnor U911 (N_911,N_768,N_747);
nor U912 (N_912,N_703,N_660);
nand U913 (N_913,N_743,N_627);
and U914 (N_914,N_649,N_704);
or U915 (N_915,N_682,N_666);
nand U916 (N_916,N_780,N_653);
or U917 (N_917,N_634,N_733);
and U918 (N_918,N_622,N_617);
nor U919 (N_919,N_749,N_761);
and U920 (N_920,N_658,N_745);
nand U921 (N_921,N_686,N_751);
or U922 (N_922,N_793,N_609);
nand U923 (N_923,N_658,N_754);
and U924 (N_924,N_753,N_693);
or U925 (N_925,N_697,N_624);
and U926 (N_926,N_686,N_624);
nor U927 (N_927,N_619,N_648);
nand U928 (N_928,N_672,N_669);
nand U929 (N_929,N_640,N_668);
nand U930 (N_930,N_607,N_666);
and U931 (N_931,N_691,N_793);
or U932 (N_932,N_723,N_778);
and U933 (N_933,N_646,N_613);
and U934 (N_934,N_646,N_635);
or U935 (N_935,N_659,N_720);
nor U936 (N_936,N_658,N_758);
nand U937 (N_937,N_723,N_719);
or U938 (N_938,N_611,N_686);
and U939 (N_939,N_633,N_750);
nand U940 (N_940,N_644,N_608);
nor U941 (N_941,N_716,N_691);
nand U942 (N_942,N_768,N_706);
or U943 (N_943,N_764,N_768);
nand U944 (N_944,N_610,N_636);
nand U945 (N_945,N_741,N_644);
or U946 (N_946,N_761,N_643);
xnor U947 (N_947,N_637,N_755);
xor U948 (N_948,N_723,N_779);
and U949 (N_949,N_660,N_620);
nand U950 (N_950,N_798,N_653);
nor U951 (N_951,N_675,N_715);
or U952 (N_952,N_735,N_660);
nand U953 (N_953,N_758,N_776);
and U954 (N_954,N_790,N_644);
nand U955 (N_955,N_623,N_768);
nand U956 (N_956,N_698,N_729);
and U957 (N_957,N_649,N_761);
or U958 (N_958,N_720,N_663);
or U959 (N_959,N_620,N_699);
and U960 (N_960,N_646,N_741);
nor U961 (N_961,N_689,N_627);
nand U962 (N_962,N_735,N_609);
and U963 (N_963,N_677,N_663);
xor U964 (N_964,N_603,N_656);
or U965 (N_965,N_650,N_798);
or U966 (N_966,N_735,N_629);
or U967 (N_967,N_778,N_793);
nand U968 (N_968,N_796,N_610);
nand U969 (N_969,N_695,N_642);
or U970 (N_970,N_794,N_685);
nor U971 (N_971,N_661,N_776);
or U972 (N_972,N_613,N_617);
nor U973 (N_973,N_726,N_728);
nor U974 (N_974,N_735,N_614);
and U975 (N_975,N_776,N_772);
nor U976 (N_976,N_624,N_764);
and U977 (N_977,N_696,N_652);
and U978 (N_978,N_629,N_604);
nand U979 (N_979,N_791,N_683);
or U980 (N_980,N_686,N_655);
and U981 (N_981,N_726,N_609);
nand U982 (N_982,N_660,N_792);
nor U983 (N_983,N_616,N_728);
or U984 (N_984,N_796,N_740);
nor U985 (N_985,N_721,N_650);
nand U986 (N_986,N_680,N_636);
nor U987 (N_987,N_743,N_725);
and U988 (N_988,N_682,N_761);
and U989 (N_989,N_619,N_614);
or U990 (N_990,N_785,N_604);
nand U991 (N_991,N_668,N_677);
or U992 (N_992,N_764,N_793);
xnor U993 (N_993,N_628,N_676);
and U994 (N_994,N_675,N_601);
and U995 (N_995,N_722,N_775);
and U996 (N_996,N_649,N_799);
nor U997 (N_997,N_661,N_635);
or U998 (N_998,N_681,N_602);
nor U999 (N_999,N_753,N_770);
and U1000 (N_1000,N_913,N_910);
or U1001 (N_1001,N_859,N_896);
nor U1002 (N_1002,N_946,N_937);
nand U1003 (N_1003,N_933,N_990);
and U1004 (N_1004,N_911,N_941);
nand U1005 (N_1005,N_805,N_814);
nand U1006 (N_1006,N_828,N_848);
or U1007 (N_1007,N_889,N_852);
or U1008 (N_1008,N_867,N_986);
and U1009 (N_1009,N_938,N_829);
nand U1010 (N_1010,N_949,N_847);
nand U1011 (N_1011,N_860,N_849);
nor U1012 (N_1012,N_975,N_870);
or U1013 (N_1013,N_837,N_952);
nand U1014 (N_1014,N_871,N_991);
nor U1015 (N_1015,N_944,N_950);
and U1016 (N_1016,N_831,N_830);
or U1017 (N_1017,N_943,N_834);
and U1018 (N_1018,N_918,N_845);
xnor U1019 (N_1019,N_916,N_930);
or U1020 (N_1020,N_994,N_800);
nand U1021 (N_1021,N_935,N_957);
nor U1022 (N_1022,N_897,N_892);
nand U1023 (N_1023,N_971,N_978);
xnor U1024 (N_1024,N_904,N_864);
nand U1025 (N_1025,N_981,N_887);
nor U1026 (N_1026,N_818,N_858);
and U1027 (N_1027,N_806,N_825);
nand U1028 (N_1028,N_980,N_919);
nand U1029 (N_1029,N_842,N_813);
nor U1030 (N_1030,N_844,N_960);
nand U1031 (N_1031,N_861,N_921);
xor U1032 (N_1032,N_823,N_917);
nor U1033 (N_1033,N_951,N_906);
nand U1034 (N_1034,N_940,N_998);
nand U1035 (N_1035,N_958,N_999);
and U1036 (N_1036,N_816,N_934);
nor U1037 (N_1037,N_977,N_912);
nand U1038 (N_1038,N_835,N_926);
and U1039 (N_1039,N_964,N_922);
nand U1040 (N_1040,N_987,N_878);
xor U1041 (N_1041,N_840,N_970);
nor U1042 (N_1042,N_909,N_915);
and U1043 (N_1043,N_826,N_968);
or U1044 (N_1044,N_932,N_850);
nand U1045 (N_1045,N_979,N_804);
or U1046 (N_1046,N_945,N_963);
or U1047 (N_1047,N_819,N_961);
xor U1048 (N_1048,N_812,N_865);
nor U1049 (N_1049,N_841,N_827);
and U1050 (N_1050,N_851,N_993);
nand U1051 (N_1051,N_923,N_927);
and U1052 (N_1052,N_900,N_839);
and U1053 (N_1053,N_976,N_882);
nand U1054 (N_1054,N_939,N_832);
nor U1055 (N_1055,N_905,N_902);
nand U1056 (N_1056,N_868,N_821);
nor U1057 (N_1057,N_803,N_914);
nand U1058 (N_1058,N_824,N_886);
and U1059 (N_1059,N_925,N_972);
nor U1060 (N_1060,N_966,N_967);
nor U1061 (N_1061,N_989,N_836);
or U1062 (N_1062,N_924,N_953);
or U1063 (N_1063,N_810,N_862);
and U1064 (N_1064,N_920,N_936);
and U1065 (N_1065,N_853,N_815);
or U1066 (N_1066,N_954,N_874);
or U1067 (N_1067,N_885,N_872);
or U1068 (N_1068,N_947,N_802);
nor U1069 (N_1069,N_891,N_908);
nand U1070 (N_1070,N_883,N_948);
xor U1071 (N_1071,N_929,N_807);
and U1072 (N_1072,N_863,N_903);
nor U1073 (N_1073,N_974,N_898);
xnor U1074 (N_1074,N_959,N_955);
and U1075 (N_1075,N_869,N_881);
and U1076 (N_1076,N_846,N_931);
nand U1077 (N_1077,N_983,N_928);
or U1078 (N_1078,N_992,N_973);
nand U1079 (N_1079,N_855,N_985);
xor U1080 (N_1080,N_895,N_893);
and U1081 (N_1081,N_884,N_997);
and U1082 (N_1082,N_956,N_820);
and U1083 (N_1083,N_995,N_817);
nand U1084 (N_1084,N_996,N_866);
and U1085 (N_1085,N_942,N_879);
nand U1086 (N_1086,N_982,N_843);
and U1087 (N_1087,N_838,N_873);
and U1088 (N_1088,N_856,N_969);
xnor U1089 (N_1089,N_877,N_962);
or U1090 (N_1090,N_875,N_880);
xnor U1091 (N_1091,N_809,N_888);
or U1092 (N_1092,N_894,N_822);
nor U1093 (N_1093,N_801,N_833);
and U1094 (N_1094,N_890,N_808);
xor U1095 (N_1095,N_984,N_811);
nor U1096 (N_1096,N_901,N_854);
nand U1097 (N_1097,N_965,N_876);
nor U1098 (N_1098,N_988,N_857);
and U1099 (N_1099,N_899,N_907);
nor U1100 (N_1100,N_933,N_852);
or U1101 (N_1101,N_838,N_914);
and U1102 (N_1102,N_800,N_870);
and U1103 (N_1103,N_904,N_940);
or U1104 (N_1104,N_898,N_841);
and U1105 (N_1105,N_839,N_988);
xnor U1106 (N_1106,N_842,N_976);
nand U1107 (N_1107,N_906,N_924);
nand U1108 (N_1108,N_939,N_961);
or U1109 (N_1109,N_835,N_843);
or U1110 (N_1110,N_930,N_998);
nand U1111 (N_1111,N_833,N_863);
nand U1112 (N_1112,N_801,N_965);
nand U1113 (N_1113,N_986,N_977);
and U1114 (N_1114,N_980,N_982);
or U1115 (N_1115,N_982,N_914);
or U1116 (N_1116,N_928,N_885);
nand U1117 (N_1117,N_977,N_846);
xor U1118 (N_1118,N_919,N_823);
nor U1119 (N_1119,N_962,N_899);
nand U1120 (N_1120,N_883,N_886);
nand U1121 (N_1121,N_969,N_898);
nand U1122 (N_1122,N_990,N_960);
xor U1123 (N_1123,N_947,N_905);
and U1124 (N_1124,N_909,N_858);
and U1125 (N_1125,N_956,N_910);
and U1126 (N_1126,N_994,N_818);
nor U1127 (N_1127,N_871,N_811);
nand U1128 (N_1128,N_922,N_852);
nand U1129 (N_1129,N_852,N_833);
and U1130 (N_1130,N_843,N_918);
and U1131 (N_1131,N_993,N_835);
nand U1132 (N_1132,N_831,N_902);
nand U1133 (N_1133,N_899,N_987);
xor U1134 (N_1134,N_875,N_827);
and U1135 (N_1135,N_814,N_891);
nand U1136 (N_1136,N_837,N_985);
nand U1137 (N_1137,N_847,N_818);
xnor U1138 (N_1138,N_917,N_861);
nor U1139 (N_1139,N_864,N_860);
and U1140 (N_1140,N_873,N_839);
and U1141 (N_1141,N_916,N_850);
nor U1142 (N_1142,N_842,N_991);
nand U1143 (N_1143,N_875,N_911);
or U1144 (N_1144,N_940,N_906);
nor U1145 (N_1145,N_815,N_842);
and U1146 (N_1146,N_884,N_919);
and U1147 (N_1147,N_919,N_997);
nand U1148 (N_1148,N_910,N_851);
nor U1149 (N_1149,N_843,N_917);
nor U1150 (N_1150,N_945,N_915);
and U1151 (N_1151,N_866,N_807);
and U1152 (N_1152,N_849,N_803);
and U1153 (N_1153,N_929,N_808);
or U1154 (N_1154,N_924,N_879);
or U1155 (N_1155,N_956,N_812);
nand U1156 (N_1156,N_852,N_853);
and U1157 (N_1157,N_944,N_946);
and U1158 (N_1158,N_866,N_893);
nor U1159 (N_1159,N_955,N_875);
nor U1160 (N_1160,N_966,N_812);
nand U1161 (N_1161,N_844,N_828);
and U1162 (N_1162,N_939,N_914);
and U1163 (N_1163,N_957,N_901);
nor U1164 (N_1164,N_864,N_830);
or U1165 (N_1165,N_854,N_943);
and U1166 (N_1166,N_829,N_875);
and U1167 (N_1167,N_998,N_814);
nor U1168 (N_1168,N_930,N_904);
nor U1169 (N_1169,N_806,N_842);
and U1170 (N_1170,N_929,N_864);
and U1171 (N_1171,N_813,N_990);
xor U1172 (N_1172,N_813,N_858);
nor U1173 (N_1173,N_815,N_952);
xor U1174 (N_1174,N_914,N_883);
and U1175 (N_1175,N_998,N_970);
and U1176 (N_1176,N_881,N_864);
nand U1177 (N_1177,N_994,N_914);
nand U1178 (N_1178,N_956,N_960);
or U1179 (N_1179,N_885,N_932);
nand U1180 (N_1180,N_800,N_984);
xor U1181 (N_1181,N_931,N_845);
and U1182 (N_1182,N_805,N_800);
or U1183 (N_1183,N_865,N_831);
or U1184 (N_1184,N_930,N_986);
xor U1185 (N_1185,N_887,N_995);
nand U1186 (N_1186,N_989,N_814);
nor U1187 (N_1187,N_933,N_816);
xor U1188 (N_1188,N_881,N_846);
or U1189 (N_1189,N_800,N_900);
nor U1190 (N_1190,N_988,N_883);
nand U1191 (N_1191,N_873,N_934);
nand U1192 (N_1192,N_808,N_818);
nand U1193 (N_1193,N_990,N_988);
nand U1194 (N_1194,N_956,N_901);
xnor U1195 (N_1195,N_857,N_892);
xor U1196 (N_1196,N_970,N_978);
nor U1197 (N_1197,N_837,N_897);
nor U1198 (N_1198,N_820,N_907);
or U1199 (N_1199,N_915,N_858);
nor U1200 (N_1200,N_1061,N_1069);
nand U1201 (N_1201,N_1079,N_1020);
nand U1202 (N_1202,N_1107,N_1196);
and U1203 (N_1203,N_1100,N_1117);
xor U1204 (N_1204,N_1003,N_1029);
nand U1205 (N_1205,N_1006,N_1129);
and U1206 (N_1206,N_1092,N_1170);
nand U1207 (N_1207,N_1164,N_1177);
nand U1208 (N_1208,N_1059,N_1036);
xnor U1209 (N_1209,N_1044,N_1019);
nand U1210 (N_1210,N_1083,N_1128);
nand U1211 (N_1211,N_1081,N_1017);
nor U1212 (N_1212,N_1141,N_1115);
or U1213 (N_1213,N_1048,N_1031);
xnor U1214 (N_1214,N_1013,N_1178);
and U1215 (N_1215,N_1185,N_1000);
or U1216 (N_1216,N_1102,N_1009);
and U1217 (N_1217,N_1137,N_1037);
nor U1218 (N_1218,N_1111,N_1192);
and U1219 (N_1219,N_1086,N_1063);
and U1220 (N_1220,N_1058,N_1012);
and U1221 (N_1221,N_1130,N_1035);
and U1222 (N_1222,N_1011,N_1120);
xnor U1223 (N_1223,N_1176,N_1056);
or U1224 (N_1224,N_1018,N_1110);
nor U1225 (N_1225,N_1104,N_1190);
or U1226 (N_1226,N_1132,N_1184);
or U1227 (N_1227,N_1140,N_1123);
nand U1228 (N_1228,N_1133,N_1160);
and U1229 (N_1229,N_1103,N_1191);
and U1230 (N_1230,N_1121,N_1015);
nand U1231 (N_1231,N_1147,N_1051);
or U1232 (N_1232,N_1070,N_1023);
and U1233 (N_1233,N_1161,N_1085);
or U1234 (N_1234,N_1050,N_1150);
xor U1235 (N_1235,N_1088,N_1138);
or U1236 (N_1236,N_1074,N_1008);
or U1237 (N_1237,N_1146,N_1106);
nand U1238 (N_1238,N_1093,N_1022);
nand U1239 (N_1239,N_1149,N_1001);
and U1240 (N_1240,N_1135,N_1126);
nor U1241 (N_1241,N_1116,N_1041);
nand U1242 (N_1242,N_1096,N_1194);
or U1243 (N_1243,N_1142,N_1034);
nand U1244 (N_1244,N_1193,N_1172);
or U1245 (N_1245,N_1005,N_1040);
nor U1246 (N_1246,N_1122,N_1167);
nor U1247 (N_1247,N_1014,N_1109);
and U1248 (N_1248,N_1181,N_1077);
and U1249 (N_1249,N_1045,N_1024);
nor U1250 (N_1250,N_1156,N_1047);
nor U1251 (N_1251,N_1112,N_1025);
nor U1252 (N_1252,N_1113,N_1028);
or U1253 (N_1253,N_1002,N_1175);
and U1254 (N_1254,N_1007,N_1187);
and U1255 (N_1255,N_1134,N_1078);
or U1256 (N_1256,N_1065,N_1108);
or U1257 (N_1257,N_1091,N_1136);
and U1258 (N_1258,N_1188,N_1189);
and U1259 (N_1259,N_1046,N_1032);
or U1260 (N_1260,N_1021,N_1072);
and U1261 (N_1261,N_1197,N_1062);
xor U1262 (N_1262,N_1154,N_1076);
nor U1263 (N_1263,N_1052,N_1016);
xnor U1264 (N_1264,N_1105,N_1101);
or U1265 (N_1265,N_1162,N_1080);
or U1266 (N_1266,N_1097,N_1038);
xnor U1267 (N_1267,N_1186,N_1068);
xor U1268 (N_1268,N_1124,N_1098);
nor U1269 (N_1269,N_1151,N_1087);
or U1270 (N_1270,N_1064,N_1033);
nand U1271 (N_1271,N_1173,N_1071);
xnor U1272 (N_1272,N_1127,N_1148);
and U1273 (N_1273,N_1159,N_1174);
or U1274 (N_1274,N_1166,N_1179);
or U1275 (N_1275,N_1180,N_1143);
nand U1276 (N_1276,N_1073,N_1010);
nor U1277 (N_1277,N_1095,N_1075);
or U1278 (N_1278,N_1183,N_1195);
and U1279 (N_1279,N_1153,N_1145);
and U1280 (N_1280,N_1089,N_1067);
nand U1281 (N_1281,N_1094,N_1042);
nor U1282 (N_1282,N_1066,N_1055);
or U1283 (N_1283,N_1118,N_1039);
or U1284 (N_1284,N_1054,N_1169);
nor U1285 (N_1285,N_1060,N_1119);
nand U1286 (N_1286,N_1057,N_1026);
nor U1287 (N_1287,N_1158,N_1082);
or U1288 (N_1288,N_1090,N_1131);
and U1289 (N_1289,N_1198,N_1152);
nor U1290 (N_1290,N_1171,N_1182);
or U1291 (N_1291,N_1165,N_1157);
nor U1292 (N_1292,N_1168,N_1099);
xor U1293 (N_1293,N_1004,N_1199);
nor U1294 (N_1294,N_1049,N_1139);
and U1295 (N_1295,N_1144,N_1114);
nand U1296 (N_1296,N_1125,N_1027);
xor U1297 (N_1297,N_1053,N_1084);
and U1298 (N_1298,N_1155,N_1030);
or U1299 (N_1299,N_1163,N_1043);
and U1300 (N_1300,N_1135,N_1111);
nand U1301 (N_1301,N_1055,N_1069);
nor U1302 (N_1302,N_1068,N_1001);
and U1303 (N_1303,N_1178,N_1051);
nor U1304 (N_1304,N_1033,N_1093);
nor U1305 (N_1305,N_1111,N_1152);
and U1306 (N_1306,N_1169,N_1045);
nand U1307 (N_1307,N_1003,N_1113);
nor U1308 (N_1308,N_1126,N_1078);
and U1309 (N_1309,N_1064,N_1101);
and U1310 (N_1310,N_1125,N_1162);
nor U1311 (N_1311,N_1174,N_1152);
or U1312 (N_1312,N_1011,N_1175);
and U1313 (N_1313,N_1114,N_1138);
nor U1314 (N_1314,N_1033,N_1078);
and U1315 (N_1315,N_1085,N_1093);
xnor U1316 (N_1316,N_1047,N_1109);
or U1317 (N_1317,N_1184,N_1080);
and U1318 (N_1318,N_1141,N_1195);
and U1319 (N_1319,N_1159,N_1050);
or U1320 (N_1320,N_1117,N_1148);
or U1321 (N_1321,N_1030,N_1019);
nand U1322 (N_1322,N_1055,N_1139);
nor U1323 (N_1323,N_1137,N_1185);
and U1324 (N_1324,N_1059,N_1111);
xnor U1325 (N_1325,N_1152,N_1040);
nand U1326 (N_1326,N_1098,N_1134);
nand U1327 (N_1327,N_1118,N_1121);
or U1328 (N_1328,N_1192,N_1140);
and U1329 (N_1329,N_1020,N_1055);
or U1330 (N_1330,N_1148,N_1064);
and U1331 (N_1331,N_1059,N_1001);
nand U1332 (N_1332,N_1174,N_1132);
xnor U1333 (N_1333,N_1029,N_1080);
nor U1334 (N_1334,N_1111,N_1182);
nand U1335 (N_1335,N_1078,N_1059);
or U1336 (N_1336,N_1044,N_1061);
and U1337 (N_1337,N_1174,N_1196);
or U1338 (N_1338,N_1164,N_1139);
xor U1339 (N_1339,N_1041,N_1047);
nand U1340 (N_1340,N_1175,N_1181);
or U1341 (N_1341,N_1050,N_1005);
nor U1342 (N_1342,N_1100,N_1042);
and U1343 (N_1343,N_1118,N_1140);
or U1344 (N_1344,N_1101,N_1085);
nand U1345 (N_1345,N_1167,N_1062);
xor U1346 (N_1346,N_1112,N_1004);
or U1347 (N_1347,N_1049,N_1041);
xor U1348 (N_1348,N_1161,N_1060);
nor U1349 (N_1349,N_1083,N_1008);
xor U1350 (N_1350,N_1148,N_1025);
and U1351 (N_1351,N_1016,N_1011);
nor U1352 (N_1352,N_1017,N_1061);
or U1353 (N_1353,N_1144,N_1160);
and U1354 (N_1354,N_1092,N_1010);
or U1355 (N_1355,N_1160,N_1183);
and U1356 (N_1356,N_1137,N_1118);
or U1357 (N_1357,N_1116,N_1139);
nand U1358 (N_1358,N_1176,N_1002);
or U1359 (N_1359,N_1115,N_1138);
and U1360 (N_1360,N_1094,N_1046);
nor U1361 (N_1361,N_1134,N_1064);
nor U1362 (N_1362,N_1024,N_1042);
or U1363 (N_1363,N_1060,N_1109);
or U1364 (N_1364,N_1194,N_1028);
or U1365 (N_1365,N_1100,N_1036);
and U1366 (N_1366,N_1010,N_1170);
or U1367 (N_1367,N_1088,N_1169);
or U1368 (N_1368,N_1098,N_1069);
and U1369 (N_1369,N_1039,N_1017);
and U1370 (N_1370,N_1142,N_1047);
nor U1371 (N_1371,N_1027,N_1078);
nand U1372 (N_1372,N_1043,N_1052);
nand U1373 (N_1373,N_1017,N_1100);
xnor U1374 (N_1374,N_1090,N_1030);
and U1375 (N_1375,N_1177,N_1126);
and U1376 (N_1376,N_1028,N_1062);
and U1377 (N_1377,N_1137,N_1140);
xor U1378 (N_1378,N_1013,N_1019);
nor U1379 (N_1379,N_1161,N_1076);
or U1380 (N_1380,N_1089,N_1193);
xnor U1381 (N_1381,N_1120,N_1008);
and U1382 (N_1382,N_1067,N_1149);
nor U1383 (N_1383,N_1098,N_1036);
nand U1384 (N_1384,N_1018,N_1104);
nand U1385 (N_1385,N_1153,N_1096);
or U1386 (N_1386,N_1162,N_1184);
and U1387 (N_1387,N_1067,N_1084);
nand U1388 (N_1388,N_1195,N_1000);
xor U1389 (N_1389,N_1009,N_1026);
and U1390 (N_1390,N_1189,N_1089);
or U1391 (N_1391,N_1053,N_1161);
nand U1392 (N_1392,N_1161,N_1096);
xor U1393 (N_1393,N_1186,N_1025);
nand U1394 (N_1394,N_1025,N_1133);
or U1395 (N_1395,N_1059,N_1049);
or U1396 (N_1396,N_1182,N_1186);
nand U1397 (N_1397,N_1009,N_1096);
or U1398 (N_1398,N_1162,N_1014);
nand U1399 (N_1399,N_1024,N_1068);
xnor U1400 (N_1400,N_1356,N_1201);
nand U1401 (N_1401,N_1210,N_1380);
nand U1402 (N_1402,N_1397,N_1343);
nand U1403 (N_1403,N_1353,N_1249);
xor U1404 (N_1404,N_1332,N_1294);
nor U1405 (N_1405,N_1345,N_1290);
and U1406 (N_1406,N_1256,N_1318);
nor U1407 (N_1407,N_1339,N_1265);
or U1408 (N_1408,N_1347,N_1317);
xor U1409 (N_1409,N_1323,N_1218);
nand U1410 (N_1410,N_1331,N_1320);
nor U1411 (N_1411,N_1241,N_1221);
and U1412 (N_1412,N_1258,N_1319);
xor U1413 (N_1413,N_1292,N_1269);
nor U1414 (N_1414,N_1285,N_1222);
xor U1415 (N_1415,N_1350,N_1276);
and U1416 (N_1416,N_1229,N_1238);
and U1417 (N_1417,N_1307,N_1378);
nor U1418 (N_1418,N_1208,N_1223);
nor U1419 (N_1419,N_1302,N_1342);
or U1420 (N_1420,N_1361,N_1274);
nand U1421 (N_1421,N_1291,N_1263);
or U1422 (N_1422,N_1390,N_1384);
nand U1423 (N_1423,N_1227,N_1370);
and U1424 (N_1424,N_1388,N_1346);
or U1425 (N_1425,N_1209,N_1309);
and U1426 (N_1426,N_1219,N_1373);
nand U1427 (N_1427,N_1205,N_1359);
nor U1428 (N_1428,N_1298,N_1305);
or U1429 (N_1429,N_1243,N_1213);
and U1430 (N_1430,N_1293,N_1216);
nor U1431 (N_1431,N_1391,N_1341);
or U1432 (N_1432,N_1369,N_1286);
nor U1433 (N_1433,N_1396,N_1366);
nand U1434 (N_1434,N_1214,N_1364);
nor U1435 (N_1435,N_1280,N_1371);
or U1436 (N_1436,N_1299,N_1228);
nor U1437 (N_1437,N_1313,N_1338);
and U1438 (N_1438,N_1230,N_1275);
nand U1439 (N_1439,N_1304,N_1204);
nor U1440 (N_1440,N_1233,N_1224);
or U1441 (N_1441,N_1351,N_1267);
and U1442 (N_1442,N_1215,N_1310);
or U1443 (N_1443,N_1308,N_1301);
or U1444 (N_1444,N_1374,N_1277);
and U1445 (N_1445,N_1283,N_1245);
nor U1446 (N_1446,N_1336,N_1329);
nand U1447 (N_1447,N_1352,N_1273);
xor U1448 (N_1448,N_1225,N_1337);
and U1449 (N_1449,N_1255,N_1316);
or U1450 (N_1450,N_1251,N_1253);
or U1451 (N_1451,N_1385,N_1322);
and U1452 (N_1452,N_1232,N_1300);
nand U1453 (N_1453,N_1207,N_1247);
and U1454 (N_1454,N_1239,N_1279);
and U1455 (N_1455,N_1237,N_1379);
nand U1456 (N_1456,N_1288,N_1367);
or U1457 (N_1457,N_1262,N_1314);
xor U1458 (N_1458,N_1375,N_1268);
or U1459 (N_1459,N_1244,N_1200);
or U1460 (N_1460,N_1250,N_1387);
or U1461 (N_1461,N_1248,N_1303);
or U1462 (N_1462,N_1334,N_1335);
and U1463 (N_1463,N_1358,N_1321);
or U1464 (N_1464,N_1254,N_1312);
xnor U1465 (N_1465,N_1354,N_1257);
or U1466 (N_1466,N_1376,N_1372);
and U1467 (N_1467,N_1333,N_1355);
and U1468 (N_1468,N_1324,N_1392);
nor U1469 (N_1469,N_1377,N_1287);
nor U1470 (N_1470,N_1211,N_1281);
and U1471 (N_1471,N_1368,N_1252);
nand U1472 (N_1472,N_1278,N_1203);
or U1473 (N_1473,N_1226,N_1271);
or U1474 (N_1474,N_1217,N_1357);
nor U1475 (N_1475,N_1260,N_1289);
xnor U1476 (N_1476,N_1365,N_1297);
or U1477 (N_1477,N_1348,N_1315);
and U1478 (N_1478,N_1264,N_1246);
and U1479 (N_1479,N_1382,N_1270);
nand U1480 (N_1480,N_1235,N_1311);
and U1481 (N_1481,N_1326,N_1360);
nand U1482 (N_1482,N_1328,N_1242);
nand U1483 (N_1483,N_1330,N_1327);
or U1484 (N_1484,N_1325,N_1240);
nand U1485 (N_1485,N_1394,N_1381);
or U1486 (N_1486,N_1295,N_1220);
nand U1487 (N_1487,N_1236,N_1344);
or U1488 (N_1488,N_1383,N_1389);
nand U1489 (N_1489,N_1363,N_1362);
nor U1490 (N_1490,N_1296,N_1386);
and U1491 (N_1491,N_1234,N_1340);
nand U1492 (N_1492,N_1202,N_1261);
or U1493 (N_1493,N_1259,N_1282);
nand U1494 (N_1494,N_1306,N_1231);
xor U1495 (N_1495,N_1393,N_1399);
and U1496 (N_1496,N_1284,N_1266);
nand U1497 (N_1497,N_1212,N_1395);
and U1498 (N_1498,N_1206,N_1398);
nor U1499 (N_1499,N_1272,N_1349);
and U1500 (N_1500,N_1338,N_1279);
nor U1501 (N_1501,N_1305,N_1390);
nor U1502 (N_1502,N_1210,N_1391);
and U1503 (N_1503,N_1210,N_1259);
and U1504 (N_1504,N_1296,N_1329);
and U1505 (N_1505,N_1358,N_1365);
nor U1506 (N_1506,N_1221,N_1314);
or U1507 (N_1507,N_1291,N_1389);
or U1508 (N_1508,N_1282,N_1271);
and U1509 (N_1509,N_1270,N_1287);
or U1510 (N_1510,N_1351,N_1248);
nor U1511 (N_1511,N_1399,N_1329);
nand U1512 (N_1512,N_1340,N_1296);
xor U1513 (N_1513,N_1342,N_1244);
nor U1514 (N_1514,N_1385,N_1367);
and U1515 (N_1515,N_1256,N_1310);
nor U1516 (N_1516,N_1339,N_1270);
nor U1517 (N_1517,N_1275,N_1352);
nor U1518 (N_1518,N_1374,N_1279);
nand U1519 (N_1519,N_1253,N_1367);
nor U1520 (N_1520,N_1325,N_1376);
or U1521 (N_1521,N_1391,N_1202);
or U1522 (N_1522,N_1336,N_1237);
nand U1523 (N_1523,N_1367,N_1279);
nand U1524 (N_1524,N_1245,N_1239);
nand U1525 (N_1525,N_1375,N_1264);
or U1526 (N_1526,N_1393,N_1367);
nor U1527 (N_1527,N_1376,N_1331);
or U1528 (N_1528,N_1362,N_1375);
nand U1529 (N_1529,N_1278,N_1271);
or U1530 (N_1530,N_1277,N_1249);
or U1531 (N_1531,N_1316,N_1357);
or U1532 (N_1532,N_1381,N_1292);
and U1533 (N_1533,N_1233,N_1211);
or U1534 (N_1534,N_1205,N_1243);
nor U1535 (N_1535,N_1358,N_1227);
nand U1536 (N_1536,N_1383,N_1242);
or U1537 (N_1537,N_1349,N_1220);
or U1538 (N_1538,N_1208,N_1235);
nor U1539 (N_1539,N_1227,N_1368);
or U1540 (N_1540,N_1338,N_1335);
nand U1541 (N_1541,N_1274,N_1227);
and U1542 (N_1542,N_1380,N_1299);
or U1543 (N_1543,N_1393,N_1375);
or U1544 (N_1544,N_1388,N_1291);
and U1545 (N_1545,N_1348,N_1332);
nand U1546 (N_1546,N_1372,N_1369);
and U1547 (N_1547,N_1356,N_1255);
nand U1548 (N_1548,N_1328,N_1307);
and U1549 (N_1549,N_1377,N_1372);
and U1550 (N_1550,N_1246,N_1206);
or U1551 (N_1551,N_1338,N_1229);
or U1552 (N_1552,N_1394,N_1334);
or U1553 (N_1553,N_1294,N_1377);
nand U1554 (N_1554,N_1298,N_1323);
and U1555 (N_1555,N_1356,N_1212);
and U1556 (N_1556,N_1309,N_1397);
and U1557 (N_1557,N_1295,N_1254);
or U1558 (N_1558,N_1387,N_1383);
nor U1559 (N_1559,N_1334,N_1390);
nor U1560 (N_1560,N_1222,N_1227);
or U1561 (N_1561,N_1300,N_1206);
or U1562 (N_1562,N_1381,N_1319);
nor U1563 (N_1563,N_1349,N_1362);
and U1564 (N_1564,N_1372,N_1215);
and U1565 (N_1565,N_1353,N_1323);
or U1566 (N_1566,N_1288,N_1220);
and U1567 (N_1567,N_1312,N_1393);
or U1568 (N_1568,N_1250,N_1200);
and U1569 (N_1569,N_1267,N_1239);
nand U1570 (N_1570,N_1363,N_1350);
and U1571 (N_1571,N_1319,N_1207);
nand U1572 (N_1572,N_1290,N_1237);
nand U1573 (N_1573,N_1251,N_1313);
and U1574 (N_1574,N_1363,N_1320);
nand U1575 (N_1575,N_1255,N_1249);
or U1576 (N_1576,N_1239,N_1248);
or U1577 (N_1577,N_1262,N_1269);
or U1578 (N_1578,N_1326,N_1244);
and U1579 (N_1579,N_1313,N_1345);
or U1580 (N_1580,N_1310,N_1377);
or U1581 (N_1581,N_1203,N_1210);
and U1582 (N_1582,N_1254,N_1308);
or U1583 (N_1583,N_1382,N_1346);
and U1584 (N_1584,N_1319,N_1242);
or U1585 (N_1585,N_1299,N_1272);
or U1586 (N_1586,N_1214,N_1277);
and U1587 (N_1587,N_1204,N_1303);
nor U1588 (N_1588,N_1203,N_1394);
or U1589 (N_1589,N_1332,N_1399);
xnor U1590 (N_1590,N_1299,N_1251);
or U1591 (N_1591,N_1219,N_1277);
or U1592 (N_1592,N_1212,N_1336);
or U1593 (N_1593,N_1306,N_1307);
nand U1594 (N_1594,N_1265,N_1232);
or U1595 (N_1595,N_1308,N_1379);
nor U1596 (N_1596,N_1316,N_1281);
nand U1597 (N_1597,N_1222,N_1232);
nand U1598 (N_1598,N_1304,N_1235);
nor U1599 (N_1599,N_1243,N_1207);
or U1600 (N_1600,N_1400,N_1560);
and U1601 (N_1601,N_1475,N_1563);
nand U1602 (N_1602,N_1558,N_1582);
nor U1603 (N_1603,N_1439,N_1430);
nand U1604 (N_1604,N_1568,N_1588);
xor U1605 (N_1605,N_1519,N_1492);
nor U1606 (N_1606,N_1442,N_1455);
xor U1607 (N_1607,N_1459,N_1498);
nand U1608 (N_1608,N_1411,N_1522);
xor U1609 (N_1609,N_1458,N_1594);
or U1610 (N_1610,N_1420,N_1580);
and U1611 (N_1611,N_1443,N_1518);
nor U1612 (N_1612,N_1462,N_1567);
and U1613 (N_1613,N_1461,N_1510);
nand U1614 (N_1614,N_1431,N_1419);
nand U1615 (N_1615,N_1493,N_1495);
nor U1616 (N_1616,N_1465,N_1441);
or U1617 (N_1617,N_1479,N_1422);
nand U1618 (N_1618,N_1526,N_1482);
and U1619 (N_1619,N_1547,N_1586);
nand U1620 (N_1620,N_1546,N_1432);
xnor U1621 (N_1621,N_1515,N_1486);
nand U1622 (N_1622,N_1483,N_1406);
nor U1623 (N_1623,N_1589,N_1418);
xor U1624 (N_1624,N_1545,N_1485);
nand U1625 (N_1625,N_1478,N_1573);
nor U1626 (N_1626,N_1408,N_1529);
nand U1627 (N_1627,N_1579,N_1550);
nand U1628 (N_1628,N_1513,N_1543);
nand U1629 (N_1629,N_1593,N_1481);
nor U1630 (N_1630,N_1544,N_1596);
nand U1631 (N_1631,N_1409,N_1554);
nand U1632 (N_1632,N_1464,N_1444);
xnor U1633 (N_1633,N_1553,N_1427);
nor U1634 (N_1634,N_1506,N_1583);
nor U1635 (N_1635,N_1562,N_1440);
or U1636 (N_1636,N_1565,N_1435);
and U1637 (N_1637,N_1433,N_1404);
and U1638 (N_1638,N_1574,N_1595);
nor U1639 (N_1639,N_1477,N_1488);
nor U1640 (N_1640,N_1533,N_1448);
nand U1641 (N_1641,N_1437,N_1598);
and U1642 (N_1642,N_1502,N_1561);
nand U1643 (N_1643,N_1436,N_1512);
xnor U1644 (N_1644,N_1552,N_1487);
or U1645 (N_1645,N_1538,N_1523);
nand U1646 (N_1646,N_1555,N_1549);
nand U1647 (N_1647,N_1508,N_1514);
or U1648 (N_1648,N_1470,N_1524);
nor U1649 (N_1649,N_1410,N_1457);
nor U1650 (N_1650,N_1467,N_1413);
or U1651 (N_1651,N_1445,N_1532);
nand U1652 (N_1652,N_1490,N_1402);
and U1653 (N_1653,N_1489,N_1438);
xor U1654 (N_1654,N_1536,N_1497);
nand U1655 (N_1655,N_1539,N_1548);
nor U1656 (N_1656,N_1591,N_1599);
or U1657 (N_1657,N_1521,N_1585);
and U1658 (N_1658,N_1511,N_1575);
and U1659 (N_1659,N_1429,N_1405);
xor U1660 (N_1660,N_1449,N_1452);
nor U1661 (N_1661,N_1557,N_1572);
and U1662 (N_1662,N_1531,N_1463);
nand U1663 (N_1663,N_1499,N_1484);
nand U1664 (N_1664,N_1480,N_1507);
nor U1665 (N_1665,N_1423,N_1525);
and U1666 (N_1666,N_1581,N_1504);
nand U1667 (N_1667,N_1447,N_1451);
or U1668 (N_1668,N_1450,N_1414);
nand U1669 (N_1669,N_1453,N_1428);
and U1670 (N_1670,N_1576,N_1584);
nand U1671 (N_1671,N_1520,N_1412);
and U1672 (N_1672,N_1476,N_1540);
or U1673 (N_1673,N_1434,N_1571);
nand U1674 (N_1674,N_1403,N_1541);
or U1675 (N_1675,N_1542,N_1534);
and U1676 (N_1676,N_1517,N_1577);
and U1677 (N_1677,N_1407,N_1415);
nand U1678 (N_1678,N_1425,N_1417);
nand U1679 (N_1679,N_1466,N_1421);
nor U1680 (N_1680,N_1491,N_1509);
nand U1681 (N_1681,N_1474,N_1468);
nand U1682 (N_1682,N_1416,N_1469);
nor U1683 (N_1683,N_1592,N_1535);
nand U1684 (N_1684,N_1446,N_1460);
and U1685 (N_1685,N_1503,N_1473);
nand U1686 (N_1686,N_1527,N_1426);
or U1687 (N_1687,N_1551,N_1530);
and U1688 (N_1688,N_1454,N_1501);
or U1689 (N_1689,N_1556,N_1472);
nand U1690 (N_1690,N_1566,N_1456);
xor U1691 (N_1691,N_1401,N_1564);
and U1692 (N_1692,N_1578,N_1597);
nor U1693 (N_1693,N_1505,N_1587);
nand U1694 (N_1694,N_1570,N_1424);
and U1695 (N_1695,N_1471,N_1569);
and U1696 (N_1696,N_1496,N_1590);
nand U1697 (N_1697,N_1559,N_1494);
nand U1698 (N_1698,N_1516,N_1500);
or U1699 (N_1699,N_1528,N_1537);
nor U1700 (N_1700,N_1483,N_1518);
nand U1701 (N_1701,N_1597,N_1415);
or U1702 (N_1702,N_1558,N_1538);
xor U1703 (N_1703,N_1486,N_1535);
xor U1704 (N_1704,N_1475,N_1436);
and U1705 (N_1705,N_1507,N_1422);
and U1706 (N_1706,N_1599,N_1499);
xnor U1707 (N_1707,N_1468,N_1423);
nand U1708 (N_1708,N_1463,N_1451);
nand U1709 (N_1709,N_1424,N_1575);
and U1710 (N_1710,N_1551,N_1406);
and U1711 (N_1711,N_1567,N_1423);
nand U1712 (N_1712,N_1547,N_1543);
nor U1713 (N_1713,N_1454,N_1585);
nor U1714 (N_1714,N_1422,N_1518);
or U1715 (N_1715,N_1448,N_1512);
and U1716 (N_1716,N_1401,N_1434);
or U1717 (N_1717,N_1541,N_1563);
xnor U1718 (N_1718,N_1412,N_1434);
nand U1719 (N_1719,N_1549,N_1515);
nand U1720 (N_1720,N_1422,N_1481);
and U1721 (N_1721,N_1446,N_1567);
or U1722 (N_1722,N_1520,N_1415);
nor U1723 (N_1723,N_1504,N_1595);
nand U1724 (N_1724,N_1420,N_1460);
nand U1725 (N_1725,N_1465,N_1516);
or U1726 (N_1726,N_1517,N_1462);
or U1727 (N_1727,N_1566,N_1542);
nor U1728 (N_1728,N_1412,N_1410);
and U1729 (N_1729,N_1564,N_1508);
nand U1730 (N_1730,N_1445,N_1461);
nor U1731 (N_1731,N_1511,N_1419);
or U1732 (N_1732,N_1587,N_1522);
and U1733 (N_1733,N_1512,N_1502);
nor U1734 (N_1734,N_1467,N_1409);
nor U1735 (N_1735,N_1583,N_1442);
xnor U1736 (N_1736,N_1549,N_1593);
xnor U1737 (N_1737,N_1540,N_1474);
xnor U1738 (N_1738,N_1494,N_1411);
and U1739 (N_1739,N_1420,N_1555);
nand U1740 (N_1740,N_1573,N_1453);
and U1741 (N_1741,N_1497,N_1460);
or U1742 (N_1742,N_1437,N_1401);
nand U1743 (N_1743,N_1548,N_1421);
and U1744 (N_1744,N_1415,N_1504);
or U1745 (N_1745,N_1502,N_1407);
and U1746 (N_1746,N_1590,N_1488);
and U1747 (N_1747,N_1528,N_1439);
nand U1748 (N_1748,N_1507,N_1417);
and U1749 (N_1749,N_1494,N_1546);
nor U1750 (N_1750,N_1558,N_1571);
nor U1751 (N_1751,N_1468,N_1465);
nor U1752 (N_1752,N_1538,N_1524);
and U1753 (N_1753,N_1425,N_1430);
nand U1754 (N_1754,N_1458,N_1507);
nand U1755 (N_1755,N_1498,N_1437);
nand U1756 (N_1756,N_1569,N_1580);
nand U1757 (N_1757,N_1559,N_1434);
xor U1758 (N_1758,N_1550,N_1408);
nand U1759 (N_1759,N_1482,N_1582);
nand U1760 (N_1760,N_1579,N_1557);
and U1761 (N_1761,N_1511,N_1423);
and U1762 (N_1762,N_1473,N_1596);
nand U1763 (N_1763,N_1480,N_1590);
nand U1764 (N_1764,N_1422,N_1510);
or U1765 (N_1765,N_1515,N_1400);
nand U1766 (N_1766,N_1431,N_1535);
nand U1767 (N_1767,N_1598,N_1537);
and U1768 (N_1768,N_1591,N_1458);
nand U1769 (N_1769,N_1590,N_1531);
nor U1770 (N_1770,N_1533,N_1414);
nand U1771 (N_1771,N_1562,N_1473);
xor U1772 (N_1772,N_1451,N_1472);
nor U1773 (N_1773,N_1526,N_1488);
or U1774 (N_1774,N_1443,N_1566);
or U1775 (N_1775,N_1583,N_1585);
or U1776 (N_1776,N_1407,N_1587);
nor U1777 (N_1777,N_1468,N_1512);
or U1778 (N_1778,N_1551,N_1509);
and U1779 (N_1779,N_1595,N_1424);
nor U1780 (N_1780,N_1500,N_1454);
nor U1781 (N_1781,N_1420,N_1554);
nand U1782 (N_1782,N_1427,N_1512);
nand U1783 (N_1783,N_1415,N_1565);
nand U1784 (N_1784,N_1512,N_1487);
xor U1785 (N_1785,N_1506,N_1537);
nor U1786 (N_1786,N_1492,N_1432);
nand U1787 (N_1787,N_1528,N_1409);
nor U1788 (N_1788,N_1598,N_1488);
nor U1789 (N_1789,N_1416,N_1419);
and U1790 (N_1790,N_1412,N_1498);
or U1791 (N_1791,N_1466,N_1449);
nand U1792 (N_1792,N_1518,N_1427);
nand U1793 (N_1793,N_1559,N_1413);
nor U1794 (N_1794,N_1420,N_1597);
and U1795 (N_1795,N_1580,N_1582);
nor U1796 (N_1796,N_1527,N_1594);
or U1797 (N_1797,N_1506,N_1469);
nand U1798 (N_1798,N_1420,N_1474);
or U1799 (N_1799,N_1487,N_1546);
xnor U1800 (N_1800,N_1694,N_1773);
or U1801 (N_1801,N_1741,N_1665);
xnor U1802 (N_1802,N_1639,N_1631);
nor U1803 (N_1803,N_1727,N_1737);
or U1804 (N_1804,N_1764,N_1740);
nand U1805 (N_1805,N_1643,N_1797);
nand U1806 (N_1806,N_1771,N_1689);
or U1807 (N_1807,N_1774,N_1610);
xor U1808 (N_1808,N_1707,N_1698);
nand U1809 (N_1809,N_1730,N_1726);
or U1810 (N_1810,N_1677,N_1735);
or U1811 (N_1811,N_1786,N_1780);
and U1812 (N_1812,N_1678,N_1632);
or U1813 (N_1813,N_1603,N_1746);
and U1814 (N_1814,N_1782,N_1785);
nor U1815 (N_1815,N_1719,N_1650);
xnor U1816 (N_1816,N_1614,N_1648);
or U1817 (N_1817,N_1647,N_1630);
nand U1818 (N_1818,N_1700,N_1655);
nor U1819 (N_1819,N_1680,N_1695);
xnor U1820 (N_1820,N_1792,N_1673);
nand U1821 (N_1821,N_1754,N_1667);
and U1822 (N_1822,N_1616,N_1653);
nand U1823 (N_1823,N_1795,N_1783);
and U1824 (N_1824,N_1659,N_1765);
and U1825 (N_1825,N_1621,N_1779);
xor U1826 (N_1826,N_1704,N_1758);
nor U1827 (N_1827,N_1745,N_1715);
nand U1828 (N_1828,N_1657,N_1656);
nand U1829 (N_1829,N_1766,N_1784);
and U1830 (N_1830,N_1768,N_1674);
and U1831 (N_1831,N_1775,N_1710);
nand U1832 (N_1832,N_1636,N_1761);
or U1833 (N_1833,N_1663,N_1602);
or U1834 (N_1834,N_1609,N_1660);
nor U1835 (N_1835,N_1666,N_1608);
or U1836 (N_1836,N_1791,N_1717);
and U1837 (N_1837,N_1635,N_1624);
and U1838 (N_1838,N_1645,N_1777);
nand U1839 (N_1839,N_1778,N_1601);
or U1840 (N_1840,N_1709,N_1699);
and U1841 (N_1841,N_1607,N_1628);
and U1842 (N_1842,N_1734,N_1749);
nor U1843 (N_1843,N_1685,N_1649);
nor U1844 (N_1844,N_1759,N_1733);
nand U1845 (N_1845,N_1613,N_1747);
or U1846 (N_1846,N_1728,N_1760);
xnor U1847 (N_1847,N_1713,N_1738);
nor U1848 (N_1848,N_1723,N_1744);
and U1849 (N_1849,N_1763,N_1637);
nor U1850 (N_1850,N_1725,N_1661);
and U1851 (N_1851,N_1789,N_1686);
xor U1852 (N_1852,N_1756,N_1757);
nand U1853 (N_1853,N_1794,N_1634);
and U1854 (N_1854,N_1625,N_1642);
or U1855 (N_1855,N_1753,N_1638);
nor U1856 (N_1856,N_1619,N_1743);
or U1857 (N_1857,N_1620,N_1742);
or U1858 (N_1858,N_1711,N_1702);
nand U1859 (N_1859,N_1683,N_1669);
or U1860 (N_1860,N_1676,N_1688);
nor U1861 (N_1861,N_1622,N_1796);
and U1862 (N_1862,N_1776,N_1705);
nor U1863 (N_1863,N_1605,N_1633);
nor U1864 (N_1864,N_1681,N_1793);
nand U1865 (N_1865,N_1668,N_1626);
nor U1866 (N_1866,N_1751,N_1755);
nand U1867 (N_1867,N_1684,N_1644);
xor U1868 (N_1868,N_1798,N_1722);
nor U1869 (N_1869,N_1675,N_1732);
or U1870 (N_1870,N_1623,N_1721);
nor U1871 (N_1871,N_1770,N_1662);
nand U1872 (N_1872,N_1627,N_1720);
xnor U1873 (N_1873,N_1731,N_1652);
nor U1874 (N_1874,N_1712,N_1682);
and U1875 (N_1875,N_1790,N_1629);
nand U1876 (N_1876,N_1724,N_1618);
and U1877 (N_1877,N_1748,N_1658);
and U1878 (N_1878,N_1718,N_1640);
nand U1879 (N_1879,N_1604,N_1703);
or U1880 (N_1880,N_1701,N_1615);
nand U1881 (N_1881,N_1691,N_1611);
nor U1882 (N_1882,N_1696,N_1664);
and U1883 (N_1883,N_1672,N_1772);
xor U1884 (N_1884,N_1690,N_1679);
xnor U1885 (N_1885,N_1693,N_1750);
nor U1886 (N_1886,N_1708,N_1670);
and U1887 (N_1887,N_1752,N_1600);
nor U1888 (N_1888,N_1729,N_1788);
and U1889 (N_1889,N_1671,N_1739);
or U1890 (N_1890,N_1716,N_1687);
or U1891 (N_1891,N_1762,N_1697);
nor U1892 (N_1892,N_1651,N_1799);
nand U1893 (N_1893,N_1612,N_1606);
nor U1894 (N_1894,N_1617,N_1767);
nor U1895 (N_1895,N_1736,N_1787);
nand U1896 (N_1896,N_1641,N_1769);
nand U1897 (N_1897,N_1706,N_1654);
or U1898 (N_1898,N_1714,N_1646);
or U1899 (N_1899,N_1781,N_1692);
nor U1900 (N_1900,N_1777,N_1740);
nor U1901 (N_1901,N_1663,N_1694);
or U1902 (N_1902,N_1673,N_1701);
or U1903 (N_1903,N_1765,N_1605);
nor U1904 (N_1904,N_1719,N_1682);
nor U1905 (N_1905,N_1705,N_1643);
nand U1906 (N_1906,N_1627,N_1797);
or U1907 (N_1907,N_1648,N_1771);
nor U1908 (N_1908,N_1682,N_1618);
nand U1909 (N_1909,N_1632,N_1702);
or U1910 (N_1910,N_1759,N_1611);
nand U1911 (N_1911,N_1612,N_1628);
and U1912 (N_1912,N_1662,N_1648);
nor U1913 (N_1913,N_1732,N_1799);
and U1914 (N_1914,N_1711,N_1647);
nand U1915 (N_1915,N_1659,N_1607);
nand U1916 (N_1916,N_1655,N_1650);
and U1917 (N_1917,N_1788,N_1629);
xor U1918 (N_1918,N_1605,N_1771);
nand U1919 (N_1919,N_1761,N_1744);
and U1920 (N_1920,N_1670,N_1661);
and U1921 (N_1921,N_1787,N_1671);
or U1922 (N_1922,N_1652,N_1628);
and U1923 (N_1923,N_1606,N_1677);
nand U1924 (N_1924,N_1624,N_1726);
or U1925 (N_1925,N_1784,N_1760);
and U1926 (N_1926,N_1677,N_1682);
or U1927 (N_1927,N_1746,N_1715);
or U1928 (N_1928,N_1761,N_1690);
nor U1929 (N_1929,N_1600,N_1660);
and U1930 (N_1930,N_1618,N_1671);
or U1931 (N_1931,N_1669,N_1771);
or U1932 (N_1932,N_1630,N_1765);
nor U1933 (N_1933,N_1684,N_1615);
nand U1934 (N_1934,N_1671,N_1716);
nor U1935 (N_1935,N_1787,N_1691);
or U1936 (N_1936,N_1784,N_1775);
and U1937 (N_1937,N_1666,N_1782);
and U1938 (N_1938,N_1609,N_1785);
nor U1939 (N_1939,N_1648,N_1690);
and U1940 (N_1940,N_1764,N_1665);
nor U1941 (N_1941,N_1619,N_1684);
nor U1942 (N_1942,N_1652,N_1603);
nor U1943 (N_1943,N_1784,N_1671);
and U1944 (N_1944,N_1718,N_1783);
nor U1945 (N_1945,N_1769,N_1735);
nor U1946 (N_1946,N_1626,N_1623);
and U1947 (N_1947,N_1735,N_1698);
or U1948 (N_1948,N_1702,N_1767);
nand U1949 (N_1949,N_1672,N_1683);
xnor U1950 (N_1950,N_1768,N_1642);
or U1951 (N_1951,N_1678,N_1637);
nor U1952 (N_1952,N_1600,N_1797);
xnor U1953 (N_1953,N_1659,N_1753);
or U1954 (N_1954,N_1751,N_1756);
and U1955 (N_1955,N_1606,N_1714);
and U1956 (N_1956,N_1633,N_1673);
or U1957 (N_1957,N_1780,N_1682);
or U1958 (N_1958,N_1673,N_1737);
xor U1959 (N_1959,N_1739,N_1686);
nand U1960 (N_1960,N_1650,N_1717);
or U1961 (N_1961,N_1768,N_1790);
xnor U1962 (N_1962,N_1604,N_1729);
or U1963 (N_1963,N_1658,N_1651);
and U1964 (N_1964,N_1640,N_1767);
nand U1965 (N_1965,N_1788,N_1751);
nor U1966 (N_1966,N_1797,N_1698);
and U1967 (N_1967,N_1679,N_1749);
nor U1968 (N_1968,N_1727,N_1640);
or U1969 (N_1969,N_1692,N_1615);
or U1970 (N_1970,N_1641,N_1672);
nand U1971 (N_1971,N_1768,N_1661);
nor U1972 (N_1972,N_1768,N_1718);
nor U1973 (N_1973,N_1763,N_1727);
or U1974 (N_1974,N_1654,N_1637);
or U1975 (N_1975,N_1604,N_1708);
nor U1976 (N_1976,N_1721,N_1644);
xnor U1977 (N_1977,N_1779,N_1687);
and U1978 (N_1978,N_1668,N_1741);
nor U1979 (N_1979,N_1608,N_1662);
xor U1980 (N_1980,N_1652,N_1619);
or U1981 (N_1981,N_1711,N_1782);
and U1982 (N_1982,N_1653,N_1607);
nand U1983 (N_1983,N_1739,N_1748);
nand U1984 (N_1984,N_1781,N_1690);
nand U1985 (N_1985,N_1734,N_1765);
nand U1986 (N_1986,N_1780,N_1793);
nand U1987 (N_1987,N_1650,N_1792);
nor U1988 (N_1988,N_1654,N_1790);
or U1989 (N_1989,N_1681,N_1607);
nand U1990 (N_1990,N_1660,N_1735);
or U1991 (N_1991,N_1666,N_1679);
xnor U1992 (N_1992,N_1621,N_1799);
or U1993 (N_1993,N_1603,N_1642);
nor U1994 (N_1994,N_1686,N_1661);
nand U1995 (N_1995,N_1600,N_1610);
and U1996 (N_1996,N_1625,N_1727);
xor U1997 (N_1997,N_1672,N_1736);
xnor U1998 (N_1998,N_1778,N_1678);
xnor U1999 (N_1999,N_1776,N_1640);
or U2000 (N_2000,N_1984,N_1900);
nor U2001 (N_2001,N_1965,N_1807);
and U2002 (N_2002,N_1870,N_1891);
and U2003 (N_2003,N_1836,N_1842);
and U2004 (N_2004,N_1887,N_1893);
and U2005 (N_2005,N_1915,N_1960);
and U2006 (N_2006,N_1908,N_1844);
and U2007 (N_2007,N_1888,N_1952);
or U2008 (N_2008,N_1948,N_1904);
and U2009 (N_2009,N_1875,N_1851);
nand U2010 (N_2010,N_1994,N_1881);
nor U2011 (N_2011,N_1884,N_1862);
or U2012 (N_2012,N_1961,N_1889);
nor U2013 (N_2013,N_1897,N_1976);
nand U2014 (N_2014,N_1934,N_1967);
nor U2015 (N_2015,N_1947,N_1895);
and U2016 (N_2016,N_1920,N_1944);
nand U2017 (N_2017,N_1854,N_1800);
or U2018 (N_2018,N_1864,N_1973);
nor U2019 (N_2019,N_1993,N_1931);
or U2020 (N_2020,N_1855,N_1823);
and U2021 (N_2021,N_1914,N_1865);
xor U2022 (N_2022,N_1917,N_1905);
nor U2023 (N_2023,N_1938,N_1820);
or U2024 (N_2024,N_1860,N_1958);
or U2025 (N_2025,N_1843,N_1953);
nand U2026 (N_2026,N_1968,N_1912);
nor U2027 (N_2027,N_1939,N_1959);
nand U2028 (N_2028,N_1833,N_1829);
or U2029 (N_2029,N_1809,N_1954);
nand U2030 (N_2030,N_1998,N_1879);
xor U2031 (N_2031,N_1841,N_1966);
nor U2032 (N_2032,N_1817,N_1831);
or U2033 (N_2033,N_1988,N_1838);
nand U2034 (N_2034,N_1813,N_1804);
xnor U2035 (N_2035,N_1996,N_1981);
nor U2036 (N_2036,N_1972,N_1977);
and U2037 (N_2037,N_1827,N_1882);
nor U2038 (N_2038,N_1835,N_1986);
xor U2039 (N_2039,N_1922,N_1970);
nand U2040 (N_2040,N_1877,N_1815);
nor U2041 (N_2041,N_1847,N_1909);
or U2042 (N_2042,N_1899,N_1856);
or U2043 (N_2043,N_1982,N_1987);
nand U2044 (N_2044,N_1980,N_1828);
and U2045 (N_2045,N_1866,N_1883);
and U2046 (N_2046,N_1937,N_1814);
or U2047 (N_2047,N_1999,N_1857);
nor U2048 (N_2048,N_1949,N_1818);
or U2049 (N_2049,N_1845,N_1929);
nand U2050 (N_2050,N_1907,N_1846);
or U2051 (N_2051,N_1990,N_1859);
nand U2052 (N_2052,N_1849,N_1853);
and U2053 (N_2053,N_1941,N_1918);
nor U2054 (N_2054,N_1906,N_1816);
nand U2055 (N_2055,N_1890,N_1940);
nand U2056 (N_2056,N_1808,N_1927);
nand U2057 (N_2057,N_1801,N_1943);
or U2058 (N_2058,N_1956,N_1894);
nand U2059 (N_2059,N_1848,N_1926);
and U2060 (N_2060,N_1837,N_1867);
nor U2061 (N_2061,N_1928,N_1892);
xor U2062 (N_2062,N_1810,N_1840);
and U2063 (N_2063,N_1910,N_1876);
nor U2064 (N_2064,N_1869,N_1950);
and U2065 (N_2065,N_1936,N_1834);
or U2066 (N_2066,N_1992,N_1916);
or U2067 (N_2067,N_1805,N_1880);
or U2068 (N_2068,N_1957,N_1852);
or U2069 (N_2069,N_1951,N_1896);
nand U2070 (N_2070,N_1932,N_1969);
nor U2071 (N_2071,N_1822,N_1985);
xnor U2072 (N_2072,N_1919,N_1868);
nor U2073 (N_2073,N_1911,N_1902);
or U2074 (N_2074,N_1826,N_1885);
nor U2075 (N_2075,N_1913,N_1979);
or U2076 (N_2076,N_1811,N_1878);
nand U2077 (N_2077,N_1975,N_1989);
nor U2078 (N_2078,N_1819,N_1830);
nand U2079 (N_2079,N_1858,N_1983);
nand U2080 (N_2080,N_1901,N_1946);
xnor U2081 (N_2081,N_1863,N_1995);
or U2082 (N_2082,N_1886,N_1832);
and U2083 (N_2083,N_1962,N_1812);
or U2084 (N_2084,N_1839,N_1921);
and U2085 (N_2085,N_1903,N_1978);
or U2086 (N_2086,N_1930,N_1871);
and U2087 (N_2087,N_1925,N_1850);
nor U2088 (N_2088,N_1997,N_1898);
xnor U2089 (N_2089,N_1942,N_1924);
and U2090 (N_2090,N_1971,N_1874);
nand U2091 (N_2091,N_1861,N_1935);
nand U2092 (N_2092,N_1945,N_1802);
and U2093 (N_2093,N_1872,N_1825);
nand U2094 (N_2094,N_1955,N_1963);
nand U2095 (N_2095,N_1991,N_1964);
and U2096 (N_2096,N_1824,N_1803);
or U2097 (N_2097,N_1873,N_1974);
or U2098 (N_2098,N_1933,N_1821);
nor U2099 (N_2099,N_1923,N_1806);
nand U2100 (N_2100,N_1940,N_1888);
nor U2101 (N_2101,N_1880,N_1874);
nor U2102 (N_2102,N_1880,N_1818);
xor U2103 (N_2103,N_1861,N_1820);
nand U2104 (N_2104,N_1880,N_1956);
xnor U2105 (N_2105,N_1833,N_1906);
nand U2106 (N_2106,N_1979,N_1952);
nor U2107 (N_2107,N_1815,N_1802);
xor U2108 (N_2108,N_1927,N_1999);
nand U2109 (N_2109,N_1891,N_1842);
xor U2110 (N_2110,N_1873,N_1981);
or U2111 (N_2111,N_1844,N_1824);
xor U2112 (N_2112,N_1956,N_1884);
nor U2113 (N_2113,N_1847,N_1927);
or U2114 (N_2114,N_1926,N_1905);
xnor U2115 (N_2115,N_1980,N_1978);
nand U2116 (N_2116,N_1979,N_1941);
and U2117 (N_2117,N_1804,N_1844);
and U2118 (N_2118,N_1923,N_1952);
nand U2119 (N_2119,N_1845,N_1820);
or U2120 (N_2120,N_1953,N_1874);
or U2121 (N_2121,N_1920,N_1924);
or U2122 (N_2122,N_1833,N_1949);
nor U2123 (N_2123,N_1988,N_1995);
and U2124 (N_2124,N_1975,N_1894);
xnor U2125 (N_2125,N_1981,N_1856);
nand U2126 (N_2126,N_1809,N_1946);
nor U2127 (N_2127,N_1844,N_1860);
nor U2128 (N_2128,N_1826,N_1817);
xor U2129 (N_2129,N_1980,N_1993);
xnor U2130 (N_2130,N_1925,N_1939);
and U2131 (N_2131,N_1831,N_1869);
or U2132 (N_2132,N_1926,N_1966);
or U2133 (N_2133,N_1936,N_1905);
nor U2134 (N_2134,N_1803,N_1876);
nor U2135 (N_2135,N_1995,N_1969);
and U2136 (N_2136,N_1943,N_1966);
nand U2137 (N_2137,N_1802,N_1925);
nor U2138 (N_2138,N_1996,N_1985);
xnor U2139 (N_2139,N_1809,N_1886);
nor U2140 (N_2140,N_1963,N_1980);
nor U2141 (N_2141,N_1902,N_1872);
nand U2142 (N_2142,N_1882,N_1811);
xor U2143 (N_2143,N_1824,N_1931);
nor U2144 (N_2144,N_1891,N_1850);
nand U2145 (N_2145,N_1884,N_1806);
or U2146 (N_2146,N_1891,N_1992);
nor U2147 (N_2147,N_1817,N_1888);
xnor U2148 (N_2148,N_1845,N_1937);
or U2149 (N_2149,N_1854,N_1931);
nor U2150 (N_2150,N_1948,N_1884);
nand U2151 (N_2151,N_1870,N_1883);
nand U2152 (N_2152,N_1848,N_1948);
nand U2153 (N_2153,N_1826,N_1877);
and U2154 (N_2154,N_1891,N_1867);
and U2155 (N_2155,N_1973,N_1902);
nor U2156 (N_2156,N_1843,N_1946);
or U2157 (N_2157,N_1815,N_1959);
and U2158 (N_2158,N_1824,N_1889);
nand U2159 (N_2159,N_1854,N_1831);
and U2160 (N_2160,N_1896,N_1965);
nand U2161 (N_2161,N_1905,N_1991);
nor U2162 (N_2162,N_1910,N_1833);
or U2163 (N_2163,N_1954,N_1854);
and U2164 (N_2164,N_1844,N_1981);
xor U2165 (N_2165,N_1926,N_1932);
nand U2166 (N_2166,N_1809,N_1901);
nor U2167 (N_2167,N_1819,N_1838);
nor U2168 (N_2168,N_1807,N_1806);
nand U2169 (N_2169,N_1860,N_1803);
or U2170 (N_2170,N_1806,N_1905);
nor U2171 (N_2171,N_1875,N_1991);
and U2172 (N_2172,N_1886,N_1833);
nand U2173 (N_2173,N_1925,N_1881);
nand U2174 (N_2174,N_1996,N_1956);
and U2175 (N_2175,N_1800,N_1822);
and U2176 (N_2176,N_1962,N_1883);
nand U2177 (N_2177,N_1815,N_1850);
and U2178 (N_2178,N_1960,N_1983);
and U2179 (N_2179,N_1962,N_1845);
or U2180 (N_2180,N_1939,N_1809);
nor U2181 (N_2181,N_1970,N_1895);
nor U2182 (N_2182,N_1840,N_1975);
nor U2183 (N_2183,N_1909,N_1960);
and U2184 (N_2184,N_1856,N_1933);
or U2185 (N_2185,N_1935,N_1893);
nor U2186 (N_2186,N_1942,N_1872);
and U2187 (N_2187,N_1899,N_1949);
or U2188 (N_2188,N_1817,N_1891);
nor U2189 (N_2189,N_1912,N_1988);
xnor U2190 (N_2190,N_1842,N_1826);
xor U2191 (N_2191,N_1967,N_1819);
and U2192 (N_2192,N_1825,N_1803);
or U2193 (N_2193,N_1974,N_1847);
xor U2194 (N_2194,N_1867,N_1958);
nand U2195 (N_2195,N_1836,N_1877);
or U2196 (N_2196,N_1935,N_1851);
and U2197 (N_2197,N_1969,N_1879);
and U2198 (N_2198,N_1952,N_1871);
or U2199 (N_2199,N_1838,N_1812);
nand U2200 (N_2200,N_2156,N_2188);
nand U2201 (N_2201,N_2114,N_2033);
nand U2202 (N_2202,N_2009,N_2141);
nand U2203 (N_2203,N_2029,N_2035);
and U2204 (N_2204,N_2086,N_2112);
nand U2205 (N_2205,N_2129,N_2131);
and U2206 (N_2206,N_2026,N_2031);
and U2207 (N_2207,N_2117,N_2122);
nor U2208 (N_2208,N_2099,N_2014);
and U2209 (N_2209,N_2187,N_2028);
nor U2210 (N_2210,N_2170,N_2169);
nand U2211 (N_2211,N_2092,N_2036);
or U2212 (N_2212,N_2003,N_2042);
nand U2213 (N_2213,N_2077,N_2085);
and U2214 (N_2214,N_2037,N_2139);
or U2215 (N_2215,N_2019,N_2032);
nor U2216 (N_2216,N_2113,N_2124);
and U2217 (N_2217,N_2105,N_2055);
or U2218 (N_2218,N_2051,N_2175);
nand U2219 (N_2219,N_2178,N_2103);
or U2220 (N_2220,N_2094,N_2142);
nand U2221 (N_2221,N_2147,N_2118);
nand U2222 (N_2222,N_2180,N_2193);
and U2223 (N_2223,N_2177,N_2002);
nor U2224 (N_2224,N_2093,N_2107);
nor U2225 (N_2225,N_2174,N_2096);
and U2226 (N_2226,N_2063,N_2073);
nor U2227 (N_2227,N_2043,N_2120);
and U2228 (N_2228,N_2132,N_2184);
nand U2229 (N_2229,N_2087,N_2007);
nand U2230 (N_2230,N_2186,N_2140);
nand U2231 (N_2231,N_2168,N_2091);
nand U2232 (N_2232,N_2075,N_2136);
xor U2233 (N_2233,N_2015,N_2152);
and U2234 (N_2234,N_2115,N_2098);
and U2235 (N_2235,N_2133,N_2121);
nand U2236 (N_2236,N_2171,N_2176);
nand U2237 (N_2237,N_2155,N_2017);
xnor U2238 (N_2238,N_2018,N_2199);
xor U2239 (N_2239,N_2183,N_2054);
or U2240 (N_2240,N_2069,N_2083);
nor U2241 (N_2241,N_2061,N_2046);
xor U2242 (N_2242,N_2125,N_2135);
nor U2243 (N_2243,N_2010,N_2182);
or U2244 (N_2244,N_2194,N_2078);
and U2245 (N_2245,N_2104,N_2161);
or U2246 (N_2246,N_2151,N_2082);
nand U2247 (N_2247,N_2192,N_2145);
nand U2248 (N_2248,N_2181,N_2079);
nor U2249 (N_2249,N_2158,N_2040);
or U2250 (N_2250,N_2076,N_2106);
or U2251 (N_2251,N_2039,N_2144);
nor U2252 (N_2252,N_2025,N_2008);
and U2253 (N_2253,N_2097,N_2137);
nor U2254 (N_2254,N_2149,N_2047);
and U2255 (N_2255,N_2068,N_2001);
nor U2256 (N_2256,N_2164,N_2020);
xor U2257 (N_2257,N_2011,N_2004);
nor U2258 (N_2258,N_2130,N_2023);
and U2259 (N_2259,N_2196,N_2100);
or U2260 (N_2260,N_2024,N_2070);
and U2261 (N_2261,N_2123,N_2146);
nor U2262 (N_2262,N_2116,N_2134);
nor U2263 (N_2263,N_2165,N_2030);
nor U2264 (N_2264,N_2005,N_2034);
nor U2265 (N_2265,N_2160,N_2050);
xor U2266 (N_2266,N_2071,N_2143);
nand U2267 (N_2267,N_2006,N_2044);
xor U2268 (N_2268,N_2159,N_2128);
nor U2269 (N_2269,N_2119,N_2058);
nor U2270 (N_2270,N_2110,N_2163);
or U2271 (N_2271,N_2189,N_2045);
or U2272 (N_2272,N_2049,N_2066);
or U2273 (N_2273,N_2172,N_2162);
and U2274 (N_2274,N_2179,N_2062);
or U2275 (N_2275,N_2041,N_2190);
and U2276 (N_2276,N_2157,N_2148);
and U2277 (N_2277,N_2138,N_2198);
nor U2278 (N_2278,N_2173,N_2053);
nor U2279 (N_2279,N_2154,N_2126);
xor U2280 (N_2280,N_2111,N_2027);
nand U2281 (N_2281,N_2064,N_2048);
nand U2282 (N_2282,N_2016,N_2052);
nand U2283 (N_2283,N_2000,N_2109);
xor U2284 (N_2284,N_2074,N_2012);
nand U2285 (N_2285,N_2191,N_2195);
xnor U2286 (N_2286,N_2095,N_2166);
and U2287 (N_2287,N_2185,N_2057);
nand U2288 (N_2288,N_2088,N_2089);
and U2289 (N_2289,N_2065,N_2108);
xor U2290 (N_2290,N_2090,N_2150);
nand U2291 (N_2291,N_2101,N_2081);
xor U2292 (N_2292,N_2084,N_2072);
nor U2293 (N_2293,N_2059,N_2153);
nor U2294 (N_2294,N_2022,N_2197);
xnor U2295 (N_2295,N_2038,N_2056);
nand U2296 (N_2296,N_2167,N_2127);
nand U2297 (N_2297,N_2102,N_2060);
xnor U2298 (N_2298,N_2013,N_2021);
nor U2299 (N_2299,N_2067,N_2080);
nand U2300 (N_2300,N_2084,N_2013);
xor U2301 (N_2301,N_2104,N_2114);
nor U2302 (N_2302,N_2132,N_2072);
and U2303 (N_2303,N_2119,N_2051);
nor U2304 (N_2304,N_2152,N_2180);
nand U2305 (N_2305,N_2196,N_2045);
nand U2306 (N_2306,N_2027,N_2113);
nor U2307 (N_2307,N_2025,N_2009);
xor U2308 (N_2308,N_2087,N_2040);
nand U2309 (N_2309,N_2105,N_2145);
or U2310 (N_2310,N_2132,N_2015);
or U2311 (N_2311,N_2041,N_2152);
and U2312 (N_2312,N_2044,N_2069);
nand U2313 (N_2313,N_2093,N_2024);
or U2314 (N_2314,N_2068,N_2004);
or U2315 (N_2315,N_2179,N_2149);
or U2316 (N_2316,N_2096,N_2030);
and U2317 (N_2317,N_2098,N_2192);
xor U2318 (N_2318,N_2158,N_2105);
nor U2319 (N_2319,N_2104,N_2142);
and U2320 (N_2320,N_2013,N_2018);
or U2321 (N_2321,N_2013,N_2054);
and U2322 (N_2322,N_2006,N_2159);
nor U2323 (N_2323,N_2081,N_2022);
or U2324 (N_2324,N_2190,N_2081);
nand U2325 (N_2325,N_2094,N_2124);
nor U2326 (N_2326,N_2160,N_2158);
and U2327 (N_2327,N_2077,N_2133);
xor U2328 (N_2328,N_2053,N_2119);
nor U2329 (N_2329,N_2082,N_2095);
nor U2330 (N_2330,N_2181,N_2059);
xor U2331 (N_2331,N_2077,N_2103);
and U2332 (N_2332,N_2068,N_2071);
and U2333 (N_2333,N_2196,N_2079);
nor U2334 (N_2334,N_2145,N_2186);
nor U2335 (N_2335,N_2088,N_2114);
and U2336 (N_2336,N_2011,N_2044);
and U2337 (N_2337,N_2159,N_2190);
nand U2338 (N_2338,N_2092,N_2014);
nand U2339 (N_2339,N_2020,N_2004);
nor U2340 (N_2340,N_2127,N_2081);
nor U2341 (N_2341,N_2013,N_2190);
nor U2342 (N_2342,N_2107,N_2079);
nand U2343 (N_2343,N_2095,N_2002);
nand U2344 (N_2344,N_2032,N_2093);
or U2345 (N_2345,N_2191,N_2000);
or U2346 (N_2346,N_2079,N_2180);
and U2347 (N_2347,N_2030,N_2127);
nand U2348 (N_2348,N_2097,N_2181);
xor U2349 (N_2349,N_2024,N_2003);
nor U2350 (N_2350,N_2161,N_2143);
or U2351 (N_2351,N_2017,N_2198);
or U2352 (N_2352,N_2018,N_2110);
and U2353 (N_2353,N_2039,N_2017);
nand U2354 (N_2354,N_2188,N_2134);
or U2355 (N_2355,N_2138,N_2104);
xor U2356 (N_2356,N_2114,N_2039);
or U2357 (N_2357,N_2122,N_2181);
nor U2358 (N_2358,N_2072,N_2148);
or U2359 (N_2359,N_2066,N_2150);
or U2360 (N_2360,N_2167,N_2132);
nor U2361 (N_2361,N_2133,N_2159);
nand U2362 (N_2362,N_2131,N_2080);
nor U2363 (N_2363,N_2052,N_2021);
xor U2364 (N_2364,N_2047,N_2038);
nand U2365 (N_2365,N_2072,N_2189);
nand U2366 (N_2366,N_2104,N_2068);
or U2367 (N_2367,N_2078,N_2062);
or U2368 (N_2368,N_2096,N_2145);
and U2369 (N_2369,N_2054,N_2153);
and U2370 (N_2370,N_2119,N_2121);
or U2371 (N_2371,N_2112,N_2065);
or U2372 (N_2372,N_2179,N_2114);
xor U2373 (N_2373,N_2083,N_2099);
and U2374 (N_2374,N_2178,N_2120);
and U2375 (N_2375,N_2099,N_2123);
and U2376 (N_2376,N_2126,N_2189);
xnor U2377 (N_2377,N_2103,N_2063);
nand U2378 (N_2378,N_2070,N_2116);
or U2379 (N_2379,N_2119,N_2024);
nor U2380 (N_2380,N_2145,N_2133);
nand U2381 (N_2381,N_2062,N_2073);
and U2382 (N_2382,N_2138,N_2015);
and U2383 (N_2383,N_2127,N_2040);
xor U2384 (N_2384,N_2189,N_2007);
or U2385 (N_2385,N_2033,N_2019);
nand U2386 (N_2386,N_2009,N_2177);
xnor U2387 (N_2387,N_2082,N_2124);
and U2388 (N_2388,N_2189,N_2119);
or U2389 (N_2389,N_2189,N_2176);
or U2390 (N_2390,N_2143,N_2130);
and U2391 (N_2391,N_2088,N_2063);
nand U2392 (N_2392,N_2151,N_2127);
or U2393 (N_2393,N_2143,N_2113);
nor U2394 (N_2394,N_2145,N_2051);
nand U2395 (N_2395,N_2004,N_2106);
or U2396 (N_2396,N_2072,N_2190);
and U2397 (N_2397,N_2189,N_2100);
nor U2398 (N_2398,N_2177,N_2145);
and U2399 (N_2399,N_2140,N_2018);
nand U2400 (N_2400,N_2272,N_2375);
nand U2401 (N_2401,N_2304,N_2269);
xnor U2402 (N_2402,N_2217,N_2307);
and U2403 (N_2403,N_2349,N_2209);
nand U2404 (N_2404,N_2330,N_2323);
and U2405 (N_2405,N_2387,N_2221);
or U2406 (N_2406,N_2282,N_2252);
nand U2407 (N_2407,N_2374,N_2345);
and U2408 (N_2408,N_2225,N_2296);
and U2409 (N_2409,N_2250,N_2280);
nand U2410 (N_2410,N_2343,N_2348);
or U2411 (N_2411,N_2396,N_2376);
nand U2412 (N_2412,N_2310,N_2373);
nor U2413 (N_2413,N_2268,N_2288);
or U2414 (N_2414,N_2210,N_2226);
and U2415 (N_2415,N_2244,N_2356);
or U2416 (N_2416,N_2352,N_2227);
and U2417 (N_2417,N_2367,N_2295);
nor U2418 (N_2418,N_2372,N_2264);
or U2419 (N_2419,N_2338,N_2294);
nor U2420 (N_2420,N_2283,N_2361);
and U2421 (N_2421,N_2340,N_2362);
nand U2422 (N_2422,N_2317,N_2350);
nor U2423 (N_2423,N_2257,N_2360);
nand U2424 (N_2424,N_2214,N_2392);
nor U2425 (N_2425,N_2298,N_2398);
nor U2426 (N_2426,N_2275,N_2251);
or U2427 (N_2427,N_2293,N_2364);
or U2428 (N_2428,N_2395,N_2236);
nand U2429 (N_2429,N_2386,N_2397);
and U2430 (N_2430,N_2385,N_2270);
nand U2431 (N_2431,N_2228,N_2303);
or U2432 (N_2432,N_2201,N_2239);
and U2433 (N_2433,N_2215,N_2207);
or U2434 (N_2434,N_2271,N_2290);
or U2435 (N_2435,N_2229,N_2313);
and U2436 (N_2436,N_2377,N_2224);
xnor U2437 (N_2437,N_2318,N_2233);
nor U2438 (N_2438,N_2285,N_2322);
and U2439 (N_2439,N_2266,N_2234);
nand U2440 (N_2440,N_2337,N_2289);
nor U2441 (N_2441,N_2208,N_2306);
and U2442 (N_2442,N_2390,N_2394);
nand U2443 (N_2443,N_2389,N_2248);
nor U2444 (N_2444,N_2202,N_2391);
nand U2445 (N_2445,N_2316,N_2219);
and U2446 (N_2446,N_2238,N_2355);
nor U2447 (N_2447,N_2276,N_2324);
nand U2448 (N_2448,N_2261,N_2299);
nand U2449 (N_2449,N_2274,N_2231);
or U2450 (N_2450,N_2254,N_2216);
nor U2451 (N_2451,N_2321,N_2309);
and U2452 (N_2452,N_2240,N_2383);
or U2453 (N_2453,N_2302,N_2382);
and U2454 (N_2454,N_2308,N_2326);
and U2455 (N_2455,N_2365,N_2287);
and U2456 (N_2456,N_2319,N_2301);
nor U2457 (N_2457,N_2399,N_2247);
and U2458 (N_2458,N_2205,N_2300);
and U2459 (N_2459,N_2388,N_2212);
or U2460 (N_2460,N_2245,N_2243);
nor U2461 (N_2461,N_2237,N_2206);
nor U2462 (N_2462,N_2347,N_2292);
nand U2463 (N_2463,N_2260,N_2325);
nand U2464 (N_2464,N_2278,N_2200);
or U2465 (N_2465,N_2384,N_2258);
or U2466 (N_2466,N_2393,N_2341);
and U2467 (N_2467,N_2259,N_2267);
and U2468 (N_2468,N_2346,N_2263);
nor U2469 (N_2469,N_2332,N_2333);
nor U2470 (N_2470,N_2336,N_2327);
nor U2471 (N_2471,N_2314,N_2256);
nand U2472 (N_2472,N_2218,N_2284);
nand U2473 (N_2473,N_2235,N_2213);
nor U2474 (N_2474,N_2342,N_2328);
or U2475 (N_2475,N_2334,N_2242);
or U2476 (N_2476,N_2329,N_2368);
or U2477 (N_2477,N_2305,N_2371);
nor U2478 (N_2478,N_2354,N_2344);
or U2479 (N_2479,N_2220,N_2265);
or U2480 (N_2480,N_2320,N_2378);
nor U2481 (N_2481,N_2255,N_2363);
or U2482 (N_2482,N_2253,N_2351);
nand U2483 (N_2483,N_2366,N_2249);
and U2484 (N_2484,N_2358,N_2370);
nor U2485 (N_2485,N_2369,N_2381);
nor U2486 (N_2486,N_2286,N_2279);
nand U2487 (N_2487,N_2246,N_2273);
and U2488 (N_2488,N_2312,N_2331);
nor U2489 (N_2489,N_2277,N_2204);
nand U2490 (N_2490,N_2297,N_2335);
xnor U2491 (N_2491,N_2315,N_2379);
xor U2492 (N_2492,N_2203,N_2339);
and U2493 (N_2493,N_2223,N_2262);
nand U2494 (N_2494,N_2222,N_2281);
nand U2495 (N_2495,N_2232,N_2357);
or U2496 (N_2496,N_2291,N_2380);
or U2497 (N_2497,N_2311,N_2353);
nor U2498 (N_2498,N_2211,N_2359);
nor U2499 (N_2499,N_2230,N_2241);
nand U2500 (N_2500,N_2309,N_2312);
or U2501 (N_2501,N_2260,N_2275);
and U2502 (N_2502,N_2392,N_2386);
nor U2503 (N_2503,N_2287,N_2244);
and U2504 (N_2504,N_2202,N_2316);
nor U2505 (N_2505,N_2345,N_2282);
nor U2506 (N_2506,N_2302,N_2284);
xor U2507 (N_2507,N_2286,N_2274);
and U2508 (N_2508,N_2272,N_2345);
or U2509 (N_2509,N_2200,N_2382);
xnor U2510 (N_2510,N_2313,N_2309);
nand U2511 (N_2511,N_2292,N_2279);
nor U2512 (N_2512,N_2236,N_2323);
or U2513 (N_2513,N_2237,N_2266);
or U2514 (N_2514,N_2324,N_2272);
or U2515 (N_2515,N_2341,N_2349);
nor U2516 (N_2516,N_2234,N_2205);
or U2517 (N_2517,N_2283,N_2223);
nor U2518 (N_2518,N_2205,N_2313);
and U2519 (N_2519,N_2250,N_2316);
or U2520 (N_2520,N_2203,N_2349);
and U2521 (N_2521,N_2296,N_2294);
nand U2522 (N_2522,N_2361,N_2267);
or U2523 (N_2523,N_2241,N_2210);
and U2524 (N_2524,N_2203,N_2251);
or U2525 (N_2525,N_2273,N_2233);
and U2526 (N_2526,N_2333,N_2303);
and U2527 (N_2527,N_2374,N_2379);
nor U2528 (N_2528,N_2210,N_2378);
nor U2529 (N_2529,N_2286,N_2371);
and U2530 (N_2530,N_2210,N_2235);
and U2531 (N_2531,N_2322,N_2301);
nor U2532 (N_2532,N_2255,N_2390);
nor U2533 (N_2533,N_2205,N_2276);
nand U2534 (N_2534,N_2217,N_2389);
or U2535 (N_2535,N_2273,N_2235);
or U2536 (N_2536,N_2329,N_2375);
or U2537 (N_2537,N_2300,N_2303);
nand U2538 (N_2538,N_2375,N_2320);
and U2539 (N_2539,N_2345,N_2333);
xnor U2540 (N_2540,N_2311,N_2374);
nand U2541 (N_2541,N_2359,N_2206);
nor U2542 (N_2542,N_2209,N_2371);
xor U2543 (N_2543,N_2243,N_2397);
or U2544 (N_2544,N_2374,N_2319);
xnor U2545 (N_2545,N_2268,N_2348);
nand U2546 (N_2546,N_2252,N_2369);
nand U2547 (N_2547,N_2305,N_2326);
and U2548 (N_2548,N_2217,N_2375);
or U2549 (N_2549,N_2347,N_2349);
nor U2550 (N_2550,N_2326,N_2365);
and U2551 (N_2551,N_2386,N_2278);
nand U2552 (N_2552,N_2345,N_2386);
and U2553 (N_2553,N_2335,N_2392);
nand U2554 (N_2554,N_2315,N_2350);
or U2555 (N_2555,N_2203,N_2313);
xnor U2556 (N_2556,N_2290,N_2343);
nor U2557 (N_2557,N_2204,N_2213);
or U2558 (N_2558,N_2343,N_2254);
or U2559 (N_2559,N_2398,N_2364);
nand U2560 (N_2560,N_2224,N_2203);
and U2561 (N_2561,N_2398,N_2324);
nand U2562 (N_2562,N_2278,N_2317);
nor U2563 (N_2563,N_2376,N_2317);
or U2564 (N_2564,N_2318,N_2290);
or U2565 (N_2565,N_2350,N_2297);
and U2566 (N_2566,N_2279,N_2305);
xor U2567 (N_2567,N_2361,N_2382);
and U2568 (N_2568,N_2296,N_2310);
nor U2569 (N_2569,N_2273,N_2346);
or U2570 (N_2570,N_2367,N_2286);
or U2571 (N_2571,N_2324,N_2310);
nand U2572 (N_2572,N_2230,N_2348);
nor U2573 (N_2573,N_2308,N_2321);
and U2574 (N_2574,N_2279,N_2296);
nor U2575 (N_2575,N_2200,N_2281);
nand U2576 (N_2576,N_2256,N_2319);
nor U2577 (N_2577,N_2201,N_2276);
nand U2578 (N_2578,N_2202,N_2329);
and U2579 (N_2579,N_2392,N_2366);
or U2580 (N_2580,N_2275,N_2279);
nand U2581 (N_2581,N_2263,N_2392);
and U2582 (N_2582,N_2319,N_2365);
and U2583 (N_2583,N_2305,N_2285);
nand U2584 (N_2584,N_2263,N_2204);
or U2585 (N_2585,N_2387,N_2386);
nor U2586 (N_2586,N_2355,N_2382);
nand U2587 (N_2587,N_2228,N_2344);
nand U2588 (N_2588,N_2309,N_2259);
or U2589 (N_2589,N_2369,N_2244);
nand U2590 (N_2590,N_2380,N_2266);
nor U2591 (N_2591,N_2223,N_2357);
nor U2592 (N_2592,N_2238,N_2353);
nor U2593 (N_2593,N_2395,N_2391);
and U2594 (N_2594,N_2251,N_2245);
nor U2595 (N_2595,N_2303,N_2360);
and U2596 (N_2596,N_2293,N_2353);
or U2597 (N_2597,N_2399,N_2329);
nor U2598 (N_2598,N_2290,N_2307);
nor U2599 (N_2599,N_2218,N_2262);
xor U2600 (N_2600,N_2478,N_2501);
or U2601 (N_2601,N_2515,N_2569);
and U2602 (N_2602,N_2437,N_2516);
and U2603 (N_2603,N_2456,N_2529);
and U2604 (N_2604,N_2590,N_2416);
nor U2605 (N_2605,N_2409,N_2421);
and U2606 (N_2606,N_2581,N_2495);
nand U2607 (N_2607,N_2431,N_2553);
nand U2608 (N_2608,N_2591,N_2432);
nand U2609 (N_2609,N_2461,N_2425);
and U2610 (N_2610,N_2457,N_2400);
and U2611 (N_2611,N_2537,N_2531);
and U2612 (N_2612,N_2471,N_2522);
xor U2613 (N_2613,N_2455,N_2496);
xnor U2614 (N_2614,N_2463,N_2442);
or U2615 (N_2615,N_2443,N_2564);
or U2616 (N_2616,N_2563,N_2404);
and U2617 (N_2617,N_2540,N_2511);
nand U2618 (N_2618,N_2582,N_2459);
xor U2619 (N_2619,N_2476,N_2423);
nand U2620 (N_2620,N_2528,N_2593);
nand U2621 (N_2621,N_2481,N_2574);
and U2622 (N_2622,N_2543,N_2486);
and U2623 (N_2623,N_2587,N_2592);
or U2624 (N_2624,N_2510,N_2527);
and U2625 (N_2625,N_2545,N_2458);
nand U2626 (N_2626,N_2534,N_2597);
nor U2627 (N_2627,N_2491,N_2507);
or U2628 (N_2628,N_2467,N_2468);
nand U2629 (N_2629,N_2562,N_2503);
nand U2630 (N_2630,N_2547,N_2584);
nand U2631 (N_2631,N_2517,N_2480);
nor U2632 (N_2632,N_2559,N_2482);
nand U2633 (N_2633,N_2525,N_2402);
nand U2634 (N_2634,N_2598,N_2557);
and U2635 (N_2635,N_2505,N_2586);
nand U2636 (N_2636,N_2492,N_2578);
or U2637 (N_2637,N_2552,N_2485);
nor U2638 (N_2638,N_2538,N_2469);
and U2639 (N_2639,N_2433,N_2556);
and U2640 (N_2640,N_2464,N_2453);
or U2641 (N_2641,N_2412,N_2407);
nor U2642 (N_2642,N_2558,N_2576);
and U2643 (N_2643,N_2494,N_2484);
nand U2644 (N_2644,N_2500,N_2445);
nor U2645 (N_2645,N_2438,N_2580);
or U2646 (N_2646,N_2405,N_2436);
or U2647 (N_2647,N_2465,N_2497);
or U2648 (N_2648,N_2483,N_2520);
and U2649 (N_2649,N_2583,N_2502);
and U2650 (N_2650,N_2439,N_2533);
nand U2651 (N_2651,N_2513,N_2474);
and U2652 (N_2652,N_2594,N_2477);
nor U2653 (N_2653,N_2401,N_2506);
and U2654 (N_2654,N_2460,N_2473);
and U2655 (N_2655,N_2499,N_2523);
nor U2656 (N_2656,N_2521,N_2488);
nand U2657 (N_2657,N_2512,N_2566);
nand U2658 (N_2658,N_2429,N_2541);
and U2659 (N_2659,N_2560,N_2414);
and U2660 (N_2660,N_2408,N_2588);
and U2661 (N_2661,N_2504,N_2568);
nor U2662 (N_2662,N_2532,N_2470);
or U2663 (N_2663,N_2424,N_2447);
nor U2664 (N_2664,N_2452,N_2410);
nor U2665 (N_2665,N_2428,N_2487);
or U2666 (N_2666,N_2514,N_2403);
or U2667 (N_2667,N_2542,N_2449);
xor U2668 (N_2668,N_2422,N_2536);
nand U2669 (N_2669,N_2446,N_2595);
or U2670 (N_2670,N_2585,N_2475);
nand U2671 (N_2671,N_2508,N_2571);
nor U2672 (N_2672,N_2539,N_2417);
xor U2673 (N_2673,N_2518,N_2567);
or U2674 (N_2674,N_2589,N_2462);
or U2675 (N_2675,N_2509,N_2565);
or U2676 (N_2676,N_2554,N_2415);
or U2677 (N_2677,N_2546,N_2530);
nand U2678 (N_2678,N_2406,N_2572);
or U2679 (N_2679,N_2535,N_2444);
or U2680 (N_2680,N_2544,N_2579);
or U2681 (N_2681,N_2526,N_2427);
or U2682 (N_2682,N_2426,N_2493);
or U2683 (N_2683,N_2479,N_2561);
and U2684 (N_2684,N_2498,N_2524);
and U2685 (N_2685,N_2489,N_2435);
nor U2686 (N_2686,N_2577,N_2434);
nor U2687 (N_2687,N_2430,N_2596);
xnor U2688 (N_2688,N_2575,N_2419);
or U2689 (N_2689,N_2450,N_2599);
nor U2690 (N_2690,N_2413,N_2549);
nand U2691 (N_2691,N_2454,N_2570);
nor U2692 (N_2692,N_2519,N_2441);
and U2693 (N_2693,N_2411,N_2440);
nor U2694 (N_2694,N_2448,N_2555);
nor U2695 (N_2695,N_2472,N_2548);
nand U2696 (N_2696,N_2550,N_2573);
and U2697 (N_2697,N_2490,N_2551);
xor U2698 (N_2698,N_2466,N_2418);
nor U2699 (N_2699,N_2420,N_2451);
xnor U2700 (N_2700,N_2408,N_2528);
or U2701 (N_2701,N_2512,N_2552);
nor U2702 (N_2702,N_2436,N_2516);
and U2703 (N_2703,N_2473,N_2528);
xnor U2704 (N_2704,N_2405,N_2498);
nand U2705 (N_2705,N_2537,N_2403);
nor U2706 (N_2706,N_2547,N_2481);
and U2707 (N_2707,N_2490,N_2425);
or U2708 (N_2708,N_2421,N_2423);
nand U2709 (N_2709,N_2439,N_2501);
nand U2710 (N_2710,N_2543,N_2530);
nor U2711 (N_2711,N_2454,N_2589);
xor U2712 (N_2712,N_2554,N_2561);
and U2713 (N_2713,N_2575,N_2468);
or U2714 (N_2714,N_2542,N_2434);
nor U2715 (N_2715,N_2434,N_2562);
or U2716 (N_2716,N_2560,N_2536);
nor U2717 (N_2717,N_2587,N_2466);
nand U2718 (N_2718,N_2598,N_2540);
nand U2719 (N_2719,N_2552,N_2470);
nor U2720 (N_2720,N_2491,N_2476);
xnor U2721 (N_2721,N_2563,N_2559);
nand U2722 (N_2722,N_2507,N_2521);
or U2723 (N_2723,N_2458,N_2572);
or U2724 (N_2724,N_2519,N_2506);
and U2725 (N_2725,N_2509,N_2512);
nor U2726 (N_2726,N_2437,N_2573);
or U2727 (N_2727,N_2424,N_2509);
nand U2728 (N_2728,N_2580,N_2522);
or U2729 (N_2729,N_2411,N_2576);
nand U2730 (N_2730,N_2568,N_2423);
and U2731 (N_2731,N_2449,N_2476);
nor U2732 (N_2732,N_2555,N_2515);
or U2733 (N_2733,N_2542,N_2424);
or U2734 (N_2734,N_2502,N_2566);
or U2735 (N_2735,N_2549,N_2541);
nand U2736 (N_2736,N_2527,N_2440);
nor U2737 (N_2737,N_2564,N_2582);
nor U2738 (N_2738,N_2494,N_2535);
or U2739 (N_2739,N_2492,N_2579);
nor U2740 (N_2740,N_2415,N_2462);
nand U2741 (N_2741,N_2530,N_2590);
nor U2742 (N_2742,N_2589,N_2468);
nor U2743 (N_2743,N_2534,N_2503);
nor U2744 (N_2744,N_2562,N_2582);
nor U2745 (N_2745,N_2481,N_2420);
nand U2746 (N_2746,N_2579,N_2549);
and U2747 (N_2747,N_2428,N_2488);
and U2748 (N_2748,N_2447,N_2484);
nand U2749 (N_2749,N_2470,N_2568);
nor U2750 (N_2750,N_2593,N_2410);
or U2751 (N_2751,N_2595,N_2499);
xor U2752 (N_2752,N_2427,N_2420);
nand U2753 (N_2753,N_2401,N_2551);
and U2754 (N_2754,N_2503,N_2547);
and U2755 (N_2755,N_2539,N_2415);
nand U2756 (N_2756,N_2419,N_2415);
xor U2757 (N_2757,N_2593,N_2547);
and U2758 (N_2758,N_2409,N_2553);
and U2759 (N_2759,N_2401,N_2517);
nand U2760 (N_2760,N_2418,N_2493);
nand U2761 (N_2761,N_2560,N_2490);
and U2762 (N_2762,N_2567,N_2413);
nor U2763 (N_2763,N_2410,N_2575);
and U2764 (N_2764,N_2597,N_2459);
nor U2765 (N_2765,N_2445,N_2449);
nor U2766 (N_2766,N_2530,N_2582);
nand U2767 (N_2767,N_2441,N_2544);
and U2768 (N_2768,N_2591,N_2565);
xor U2769 (N_2769,N_2514,N_2497);
and U2770 (N_2770,N_2404,N_2540);
xor U2771 (N_2771,N_2552,N_2585);
or U2772 (N_2772,N_2594,N_2432);
or U2773 (N_2773,N_2456,N_2455);
nand U2774 (N_2774,N_2572,N_2484);
xor U2775 (N_2775,N_2567,N_2464);
or U2776 (N_2776,N_2566,N_2421);
and U2777 (N_2777,N_2563,N_2570);
and U2778 (N_2778,N_2497,N_2402);
or U2779 (N_2779,N_2457,N_2407);
nor U2780 (N_2780,N_2430,N_2575);
nor U2781 (N_2781,N_2431,N_2519);
nand U2782 (N_2782,N_2517,N_2488);
nand U2783 (N_2783,N_2457,N_2417);
xnor U2784 (N_2784,N_2535,N_2429);
nand U2785 (N_2785,N_2440,N_2510);
nand U2786 (N_2786,N_2450,N_2539);
or U2787 (N_2787,N_2530,N_2410);
and U2788 (N_2788,N_2412,N_2478);
and U2789 (N_2789,N_2599,N_2443);
and U2790 (N_2790,N_2572,N_2416);
and U2791 (N_2791,N_2500,N_2471);
nand U2792 (N_2792,N_2425,N_2510);
or U2793 (N_2793,N_2485,N_2450);
nor U2794 (N_2794,N_2538,N_2584);
and U2795 (N_2795,N_2563,N_2582);
or U2796 (N_2796,N_2562,N_2501);
or U2797 (N_2797,N_2459,N_2542);
nor U2798 (N_2798,N_2435,N_2522);
xor U2799 (N_2799,N_2545,N_2463);
xor U2800 (N_2800,N_2674,N_2744);
nand U2801 (N_2801,N_2619,N_2791);
nor U2802 (N_2802,N_2681,N_2730);
or U2803 (N_2803,N_2793,N_2666);
nor U2804 (N_2804,N_2659,N_2690);
nor U2805 (N_2805,N_2651,N_2604);
nor U2806 (N_2806,N_2646,N_2625);
xor U2807 (N_2807,N_2695,N_2778);
and U2808 (N_2808,N_2628,N_2785);
or U2809 (N_2809,N_2656,N_2622);
nand U2810 (N_2810,N_2623,N_2618);
nor U2811 (N_2811,N_2776,N_2712);
nand U2812 (N_2812,N_2749,N_2678);
nand U2813 (N_2813,N_2613,N_2707);
nand U2814 (N_2814,N_2731,N_2654);
nand U2815 (N_2815,N_2753,N_2643);
nor U2816 (N_2816,N_2772,N_2696);
and U2817 (N_2817,N_2600,N_2663);
and U2818 (N_2818,N_2692,N_2649);
nor U2819 (N_2819,N_2669,N_2718);
nor U2820 (N_2820,N_2679,N_2773);
nand U2821 (N_2821,N_2665,N_2766);
or U2822 (N_2822,N_2675,N_2637);
or U2823 (N_2823,N_2779,N_2781);
xnor U2824 (N_2824,N_2787,N_2699);
and U2825 (N_2825,N_2719,N_2631);
or U2826 (N_2826,N_2794,N_2762);
xnor U2827 (N_2827,N_2709,N_2689);
or U2828 (N_2828,N_2769,N_2615);
nor U2829 (N_2829,N_2752,N_2700);
nand U2830 (N_2830,N_2655,N_2759);
or U2831 (N_2831,N_2751,N_2677);
nand U2832 (N_2832,N_2612,N_2782);
or U2833 (N_2833,N_2605,N_2632);
and U2834 (N_2834,N_2614,N_2742);
or U2835 (N_2835,N_2662,N_2610);
or U2836 (N_2836,N_2790,N_2763);
nand U2837 (N_2837,N_2722,N_2720);
nand U2838 (N_2838,N_2682,N_2713);
or U2839 (N_2839,N_2676,N_2797);
and U2840 (N_2840,N_2765,N_2638);
or U2841 (N_2841,N_2795,N_2657);
or U2842 (N_2842,N_2647,N_2741);
or U2843 (N_2843,N_2634,N_2739);
or U2844 (N_2844,N_2672,N_2694);
nand U2845 (N_2845,N_2667,N_2653);
and U2846 (N_2846,N_2664,N_2608);
nor U2847 (N_2847,N_2764,N_2650);
nor U2848 (N_2848,N_2697,N_2774);
nand U2849 (N_2849,N_2792,N_2606);
xor U2850 (N_2850,N_2705,N_2607);
or U2851 (N_2851,N_2645,N_2685);
xnor U2852 (N_2852,N_2734,N_2726);
or U2853 (N_2853,N_2748,N_2771);
or U2854 (N_2854,N_2629,N_2740);
nor U2855 (N_2855,N_2721,N_2636);
or U2856 (N_2856,N_2783,N_2683);
or U2857 (N_2857,N_2671,N_2788);
nand U2858 (N_2858,N_2691,N_2728);
nor U2859 (N_2859,N_2796,N_2693);
nand U2860 (N_2860,N_2641,N_2703);
nor U2861 (N_2861,N_2789,N_2747);
nand U2862 (N_2862,N_2661,N_2601);
or U2863 (N_2863,N_2715,N_2743);
xor U2864 (N_2864,N_2711,N_2640);
and U2865 (N_2865,N_2799,N_2750);
nor U2866 (N_2866,N_2755,N_2770);
nand U2867 (N_2867,N_2745,N_2708);
or U2868 (N_2868,N_2777,N_2626);
or U2869 (N_2869,N_2768,N_2727);
nor U2870 (N_2870,N_2686,N_2648);
or U2871 (N_2871,N_2736,N_2684);
and U2872 (N_2872,N_2660,N_2784);
nor U2873 (N_2873,N_2746,N_2698);
xor U2874 (N_2874,N_2627,N_2609);
nor U2875 (N_2875,N_2644,N_2621);
and U2876 (N_2876,N_2658,N_2639);
and U2877 (N_2877,N_2775,N_2617);
nand U2878 (N_2878,N_2603,N_2716);
nor U2879 (N_2879,N_2602,N_2706);
or U2880 (N_2880,N_2729,N_2780);
and U2881 (N_2881,N_2760,N_2717);
xor U2882 (N_2882,N_2670,N_2668);
nor U2883 (N_2883,N_2723,N_2732);
and U2884 (N_2884,N_2767,N_2635);
nand U2885 (N_2885,N_2701,N_2761);
nand U2886 (N_2886,N_2798,N_2633);
or U2887 (N_2887,N_2786,N_2687);
nor U2888 (N_2888,N_2756,N_2738);
and U2889 (N_2889,N_2733,N_2757);
or U2890 (N_2890,N_2652,N_2737);
nor U2891 (N_2891,N_2688,N_2710);
and U2892 (N_2892,N_2754,N_2680);
nand U2893 (N_2893,N_2611,N_2624);
nand U2894 (N_2894,N_2714,N_2724);
nor U2895 (N_2895,N_2735,N_2758);
and U2896 (N_2896,N_2725,N_2702);
or U2897 (N_2897,N_2642,N_2704);
and U2898 (N_2898,N_2673,N_2630);
nor U2899 (N_2899,N_2616,N_2620);
nand U2900 (N_2900,N_2798,N_2717);
or U2901 (N_2901,N_2716,N_2647);
nand U2902 (N_2902,N_2717,N_2692);
or U2903 (N_2903,N_2761,N_2764);
and U2904 (N_2904,N_2705,N_2750);
xnor U2905 (N_2905,N_2799,N_2669);
nand U2906 (N_2906,N_2754,N_2738);
nand U2907 (N_2907,N_2693,N_2620);
nor U2908 (N_2908,N_2656,N_2671);
nand U2909 (N_2909,N_2644,N_2706);
nor U2910 (N_2910,N_2797,N_2760);
or U2911 (N_2911,N_2778,N_2687);
and U2912 (N_2912,N_2615,N_2774);
or U2913 (N_2913,N_2710,N_2612);
nand U2914 (N_2914,N_2725,N_2653);
and U2915 (N_2915,N_2660,N_2752);
or U2916 (N_2916,N_2643,N_2663);
nand U2917 (N_2917,N_2623,N_2727);
and U2918 (N_2918,N_2648,N_2627);
nor U2919 (N_2919,N_2694,N_2735);
nor U2920 (N_2920,N_2602,N_2668);
or U2921 (N_2921,N_2771,N_2638);
or U2922 (N_2922,N_2717,N_2728);
nor U2923 (N_2923,N_2729,N_2643);
xor U2924 (N_2924,N_2684,N_2635);
nand U2925 (N_2925,N_2771,N_2709);
or U2926 (N_2926,N_2619,N_2797);
or U2927 (N_2927,N_2651,N_2674);
nor U2928 (N_2928,N_2782,N_2750);
or U2929 (N_2929,N_2639,N_2757);
or U2930 (N_2930,N_2625,N_2794);
xor U2931 (N_2931,N_2695,N_2708);
and U2932 (N_2932,N_2698,N_2620);
nand U2933 (N_2933,N_2656,N_2629);
nor U2934 (N_2934,N_2734,N_2787);
or U2935 (N_2935,N_2618,N_2773);
xor U2936 (N_2936,N_2765,N_2779);
nand U2937 (N_2937,N_2759,N_2764);
xor U2938 (N_2938,N_2690,N_2744);
and U2939 (N_2939,N_2739,N_2777);
xor U2940 (N_2940,N_2721,N_2781);
nand U2941 (N_2941,N_2683,N_2735);
and U2942 (N_2942,N_2703,N_2772);
or U2943 (N_2943,N_2715,N_2681);
or U2944 (N_2944,N_2762,N_2651);
nand U2945 (N_2945,N_2779,N_2797);
nand U2946 (N_2946,N_2750,N_2714);
and U2947 (N_2947,N_2783,N_2641);
nand U2948 (N_2948,N_2704,N_2604);
nand U2949 (N_2949,N_2734,N_2753);
or U2950 (N_2950,N_2620,N_2653);
xnor U2951 (N_2951,N_2646,N_2635);
and U2952 (N_2952,N_2760,N_2682);
nor U2953 (N_2953,N_2635,N_2619);
or U2954 (N_2954,N_2774,N_2721);
nor U2955 (N_2955,N_2764,N_2659);
and U2956 (N_2956,N_2665,N_2755);
nor U2957 (N_2957,N_2607,N_2637);
nand U2958 (N_2958,N_2766,N_2672);
nor U2959 (N_2959,N_2742,N_2704);
nand U2960 (N_2960,N_2642,N_2758);
nor U2961 (N_2961,N_2762,N_2753);
nand U2962 (N_2962,N_2774,N_2786);
xnor U2963 (N_2963,N_2616,N_2781);
or U2964 (N_2964,N_2600,N_2712);
or U2965 (N_2965,N_2723,N_2770);
nor U2966 (N_2966,N_2631,N_2659);
nor U2967 (N_2967,N_2797,N_2678);
nor U2968 (N_2968,N_2762,N_2777);
nand U2969 (N_2969,N_2691,N_2719);
nor U2970 (N_2970,N_2686,N_2665);
and U2971 (N_2971,N_2640,N_2666);
and U2972 (N_2972,N_2636,N_2790);
nand U2973 (N_2973,N_2722,N_2701);
and U2974 (N_2974,N_2696,N_2678);
nor U2975 (N_2975,N_2621,N_2714);
nor U2976 (N_2976,N_2764,N_2766);
nand U2977 (N_2977,N_2631,N_2692);
nor U2978 (N_2978,N_2622,N_2772);
nor U2979 (N_2979,N_2606,N_2782);
nand U2980 (N_2980,N_2700,N_2630);
or U2981 (N_2981,N_2620,N_2703);
nor U2982 (N_2982,N_2695,N_2646);
xor U2983 (N_2983,N_2718,N_2628);
nor U2984 (N_2984,N_2643,N_2719);
and U2985 (N_2985,N_2770,N_2649);
and U2986 (N_2986,N_2628,N_2715);
nor U2987 (N_2987,N_2687,N_2689);
nor U2988 (N_2988,N_2745,N_2757);
xor U2989 (N_2989,N_2632,N_2665);
nand U2990 (N_2990,N_2695,N_2686);
or U2991 (N_2991,N_2621,N_2793);
nor U2992 (N_2992,N_2672,N_2795);
or U2993 (N_2993,N_2696,N_2610);
or U2994 (N_2994,N_2611,N_2648);
nand U2995 (N_2995,N_2635,N_2755);
and U2996 (N_2996,N_2788,N_2755);
or U2997 (N_2997,N_2768,N_2623);
nor U2998 (N_2998,N_2663,N_2607);
nor U2999 (N_2999,N_2695,N_2714);
or U3000 (N_3000,N_2952,N_2963);
nor U3001 (N_3001,N_2956,N_2808);
or U3002 (N_3002,N_2865,N_2837);
nor U3003 (N_3003,N_2847,N_2942);
xnor U3004 (N_3004,N_2899,N_2998);
nor U3005 (N_3005,N_2980,N_2997);
nand U3006 (N_3006,N_2844,N_2932);
or U3007 (N_3007,N_2981,N_2845);
nand U3008 (N_3008,N_2810,N_2850);
nand U3009 (N_3009,N_2831,N_2870);
nor U3010 (N_3010,N_2886,N_2950);
nand U3011 (N_3011,N_2922,N_2918);
and U3012 (N_3012,N_2924,N_2945);
or U3013 (N_3013,N_2839,N_2993);
nor U3014 (N_3014,N_2902,N_2852);
or U3015 (N_3015,N_2943,N_2809);
and U3016 (N_3016,N_2824,N_2987);
or U3017 (N_3017,N_2897,N_2879);
and U3018 (N_3018,N_2894,N_2919);
nand U3019 (N_3019,N_2921,N_2923);
nor U3020 (N_3020,N_2971,N_2884);
or U3021 (N_3021,N_2906,N_2848);
nand U3022 (N_3022,N_2977,N_2881);
xnor U3023 (N_3023,N_2937,N_2860);
nor U3024 (N_3024,N_2869,N_2927);
and U3025 (N_3025,N_2901,N_2815);
nand U3026 (N_3026,N_2889,N_2895);
nand U3027 (N_3027,N_2826,N_2841);
xnor U3028 (N_3028,N_2846,N_2917);
nand U3029 (N_3029,N_2802,N_2866);
nand U3030 (N_3030,N_2962,N_2887);
xor U3031 (N_3031,N_2991,N_2903);
or U3032 (N_3032,N_2931,N_2948);
nor U3033 (N_3033,N_2816,N_2909);
xnor U3034 (N_3034,N_2856,N_2957);
or U3035 (N_3035,N_2867,N_2925);
and U3036 (N_3036,N_2955,N_2842);
or U3037 (N_3037,N_2872,N_2905);
or U3038 (N_3038,N_2965,N_2936);
or U3039 (N_3039,N_2960,N_2910);
and U3040 (N_3040,N_2811,N_2983);
nand U3041 (N_3041,N_2933,N_2883);
nand U3042 (N_3042,N_2900,N_2882);
or U3043 (N_3043,N_2996,N_2949);
nor U3044 (N_3044,N_2953,N_2941);
xnor U3045 (N_3045,N_2877,N_2893);
and U3046 (N_3046,N_2836,N_2973);
nand U3047 (N_3047,N_2873,N_2911);
or U3048 (N_3048,N_2885,N_2888);
xor U3049 (N_3049,N_2859,N_2986);
or U3050 (N_3050,N_2978,N_2892);
nand U3051 (N_3051,N_2875,N_2858);
nand U3052 (N_3052,N_2995,N_2823);
nand U3053 (N_3053,N_2862,N_2999);
and U3054 (N_3054,N_2814,N_2817);
and U3055 (N_3055,N_2891,N_2840);
nor U3056 (N_3056,N_2935,N_2982);
or U3057 (N_3057,N_2807,N_2947);
or U3058 (N_3058,N_2994,N_2944);
xor U3059 (N_3059,N_2806,N_2954);
nand U3060 (N_3060,N_2857,N_2966);
xor U3061 (N_3061,N_2904,N_2861);
nor U3062 (N_3062,N_2992,N_2880);
or U3063 (N_3063,N_2908,N_2961);
nor U3064 (N_3064,N_2804,N_2812);
nor U3065 (N_3065,N_2946,N_2929);
and U3066 (N_3066,N_2827,N_2822);
or U3067 (N_3067,N_2985,N_2928);
nor U3068 (N_3068,N_2876,N_2813);
and U3069 (N_3069,N_2972,N_2926);
or U3070 (N_3070,N_2820,N_2939);
nand U3071 (N_3071,N_2851,N_2805);
and U3072 (N_3072,N_2970,N_2830);
and U3073 (N_3073,N_2801,N_2984);
and U3074 (N_3074,N_2990,N_2803);
nand U3075 (N_3075,N_2854,N_2818);
or U3076 (N_3076,N_2938,N_2969);
and U3077 (N_3077,N_2959,N_2975);
nand U3078 (N_3078,N_2915,N_2934);
nand U3079 (N_3079,N_2849,N_2920);
nor U3080 (N_3080,N_2913,N_2988);
xor U3081 (N_3081,N_2974,N_2819);
and U3082 (N_3082,N_2951,N_2958);
nor U3083 (N_3083,N_2890,N_2976);
nand U3084 (N_3084,N_2940,N_2829);
or U3085 (N_3085,N_2800,N_2989);
xor U3086 (N_3086,N_2828,N_2930);
nand U3087 (N_3087,N_2898,N_2832);
xor U3088 (N_3088,N_2964,N_2863);
and U3089 (N_3089,N_2896,N_2838);
nor U3090 (N_3090,N_2907,N_2825);
and U3091 (N_3091,N_2843,N_2835);
nand U3092 (N_3092,N_2979,N_2871);
nor U3093 (N_3093,N_2968,N_2864);
nor U3094 (N_3094,N_2914,N_2916);
or U3095 (N_3095,N_2821,N_2868);
nand U3096 (N_3096,N_2878,N_2874);
nand U3097 (N_3097,N_2853,N_2834);
or U3098 (N_3098,N_2855,N_2833);
or U3099 (N_3099,N_2967,N_2912);
nor U3100 (N_3100,N_2913,N_2859);
nand U3101 (N_3101,N_2916,N_2891);
nor U3102 (N_3102,N_2892,N_2833);
or U3103 (N_3103,N_2960,N_2851);
xnor U3104 (N_3104,N_2848,N_2901);
nor U3105 (N_3105,N_2875,N_2898);
and U3106 (N_3106,N_2910,N_2900);
nor U3107 (N_3107,N_2904,N_2869);
xnor U3108 (N_3108,N_2820,N_2941);
and U3109 (N_3109,N_2873,N_2899);
and U3110 (N_3110,N_2998,N_2842);
nor U3111 (N_3111,N_2851,N_2999);
nand U3112 (N_3112,N_2879,N_2844);
or U3113 (N_3113,N_2939,N_2840);
nand U3114 (N_3114,N_2889,N_2862);
and U3115 (N_3115,N_2812,N_2891);
or U3116 (N_3116,N_2862,N_2978);
nand U3117 (N_3117,N_2806,N_2832);
nor U3118 (N_3118,N_2839,N_2983);
nor U3119 (N_3119,N_2880,N_2862);
and U3120 (N_3120,N_2879,N_2920);
or U3121 (N_3121,N_2957,N_2824);
xor U3122 (N_3122,N_2839,N_2940);
xnor U3123 (N_3123,N_2912,N_2814);
or U3124 (N_3124,N_2850,N_2904);
and U3125 (N_3125,N_2965,N_2845);
nand U3126 (N_3126,N_2899,N_2836);
nand U3127 (N_3127,N_2952,N_2864);
nor U3128 (N_3128,N_2894,N_2845);
nand U3129 (N_3129,N_2947,N_2953);
nor U3130 (N_3130,N_2917,N_2984);
or U3131 (N_3131,N_2997,N_2877);
or U3132 (N_3132,N_2802,N_2804);
xor U3133 (N_3133,N_2816,N_2841);
and U3134 (N_3134,N_2924,N_2903);
nor U3135 (N_3135,N_2927,N_2848);
xnor U3136 (N_3136,N_2856,N_2814);
nor U3137 (N_3137,N_2860,N_2882);
and U3138 (N_3138,N_2823,N_2907);
nand U3139 (N_3139,N_2860,N_2831);
nor U3140 (N_3140,N_2816,N_2804);
nor U3141 (N_3141,N_2979,N_2875);
nor U3142 (N_3142,N_2874,N_2942);
or U3143 (N_3143,N_2973,N_2805);
and U3144 (N_3144,N_2913,N_2818);
xor U3145 (N_3145,N_2887,N_2874);
or U3146 (N_3146,N_2889,N_2884);
or U3147 (N_3147,N_2862,N_2897);
nand U3148 (N_3148,N_2885,N_2960);
nand U3149 (N_3149,N_2839,N_2815);
nand U3150 (N_3150,N_2876,N_2935);
nand U3151 (N_3151,N_2877,N_2814);
nand U3152 (N_3152,N_2991,N_2902);
nor U3153 (N_3153,N_2895,N_2810);
and U3154 (N_3154,N_2997,N_2943);
or U3155 (N_3155,N_2995,N_2863);
or U3156 (N_3156,N_2977,N_2937);
nor U3157 (N_3157,N_2909,N_2894);
and U3158 (N_3158,N_2942,N_2992);
xor U3159 (N_3159,N_2808,N_2866);
nor U3160 (N_3160,N_2915,N_2976);
nand U3161 (N_3161,N_2864,N_2946);
nor U3162 (N_3162,N_2824,N_2898);
and U3163 (N_3163,N_2934,N_2824);
and U3164 (N_3164,N_2893,N_2928);
xor U3165 (N_3165,N_2852,N_2910);
or U3166 (N_3166,N_2834,N_2888);
and U3167 (N_3167,N_2937,N_2945);
nand U3168 (N_3168,N_2835,N_2811);
and U3169 (N_3169,N_2801,N_2805);
nand U3170 (N_3170,N_2836,N_2904);
nand U3171 (N_3171,N_2853,N_2981);
nand U3172 (N_3172,N_2849,N_2851);
xor U3173 (N_3173,N_2984,N_2863);
nand U3174 (N_3174,N_2975,N_2829);
nor U3175 (N_3175,N_2897,N_2982);
nor U3176 (N_3176,N_2817,N_2892);
or U3177 (N_3177,N_2844,N_2856);
or U3178 (N_3178,N_2952,N_2878);
or U3179 (N_3179,N_2892,N_2886);
nor U3180 (N_3180,N_2915,N_2962);
and U3181 (N_3181,N_2826,N_2866);
or U3182 (N_3182,N_2905,N_2949);
nand U3183 (N_3183,N_2802,N_2812);
nor U3184 (N_3184,N_2805,N_2850);
nor U3185 (N_3185,N_2911,N_2804);
or U3186 (N_3186,N_2930,N_2884);
or U3187 (N_3187,N_2855,N_2992);
nand U3188 (N_3188,N_2939,N_2989);
and U3189 (N_3189,N_2986,N_2913);
xnor U3190 (N_3190,N_2851,N_2886);
xnor U3191 (N_3191,N_2977,N_2942);
nor U3192 (N_3192,N_2857,N_2889);
and U3193 (N_3193,N_2842,N_2870);
nand U3194 (N_3194,N_2950,N_2951);
xnor U3195 (N_3195,N_2841,N_2839);
nand U3196 (N_3196,N_2955,N_2857);
and U3197 (N_3197,N_2927,N_2895);
nor U3198 (N_3198,N_2806,N_2882);
xor U3199 (N_3199,N_2927,N_2901);
nand U3200 (N_3200,N_3194,N_3112);
nand U3201 (N_3201,N_3094,N_3044);
and U3202 (N_3202,N_3026,N_3166);
or U3203 (N_3203,N_3143,N_3134);
and U3204 (N_3204,N_3197,N_3199);
or U3205 (N_3205,N_3139,N_3122);
xnor U3206 (N_3206,N_3085,N_3058);
or U3207 (N_3207,N_3130,N_3108);
and U3208 (N_3208,N_3072,N_3086);
xnor U3209 (N_3209,N_3078,N_3135);
and U3210 (N_3210,N_3103,N_3019);
nand U3211 (N_3211,N_3041,N_3158);
nor U3212 (N_3212,N_3080,N_3119);
nand U3213 (N_3213,N_3152,N_3113);
nor U3214 (N_3214,N_3154,N_3123);
nand U3215 (N_3215,N_3181,N_3017);
nand U3216 (N_3216,N_3193,N_3136);
nand U3217 (N_3217,N_3046,N_3030);
xnor U3218 (N_3218,N_3020,N_3021);
xor U3219 (N_3219,N_3115,N_3024);
xor U3220 (N_3220,N_3079,N_3138);
or U3221 (N_3221,N_3065,N_3124);
and U3222 (N_3222,N_3137,N_3096);
xnor U3223 (N_3223,N_3029,N_3189);
or U3224 (N_3224,N_3184,N_3173);
nor U3225 (N_3225,N_3150,N_3081);
xnor U3226 (N_3226,N_3049,N_3155);
xor U3227 (N_3227,N_3187,N_3125);
nand U3228 (N_3228,N_3025,N_3090);
nor U3229 (N_3229,N_3045,N_3012);
nand U3230 (N_3230,N_3153,N_3027);
nand U3231 (N_3231,N_3056,N_3190);
nand U3232 (N_3232,N_3177,N_3164);
xor U3233 (N_3233,N_3013,N_3182);
nor U3234 (N_3234,N_3069,N_3148);
or U3235 (N_3235,N_3036,N_3057);
nor U3236 (N_3236,N_3088,N_3171);
nand U3237 (N_3237,N_3098,N_3104);
and U3238 (N_3238,N_3028,N_3099);
nor U3239 (N_3239,N_3120,N_3168);
nor U3240 (N_3240,N_3174,N_3077);
nand U3241 (N_3241,N_3083,N_3109);
nor U3242 (N_3242,N_3140,N_3059);
nand U3243 (N_3243,N_3198,N_3014);
or U3244 (N_3244,N_3070,N_3003);
nand U3245 (N_3245,N_3052,N_3195);
and U3246 (N_3246,N_3073,N_3087);
or U3247 (N_3247,N_3053,N_3179);
nand U3248 (N_3248,N_3048,N_3178);
nand U3249 (N_3249,N_3196,N_3102);
and U3250 (N_3250,N_3091,N_3031);
and U3251 (N_3251,N_3006,N_3009);
nand U3252 (N_3252,N_3071,N_3180);
nand U3253 (N_3253,N_3142,N_3082);
and U3254 (N_3254,N_3131,N_3110);
nand U3255 (N_3255,N_3067,N_3133);
nand U3256 (N_3256,N_3001,N_3097);
xnor U3257 (N_3257,N_3105,N_3183);
nor U3258 (N_3258,N_3114,N_3092);
nand U3259 (N_3259,N_3062,N_3100);
nand U3260 (N_3260,N_3037,N_3061);
or U3261 (N_3261,N_3132,N_3186);
nand U3262 (N_3262,N_3089,N_3165);
and U3263 (N_3263,N_3170,N_3188);
or U3264 (N_3264,N_3022,N_3167);
xor U3265 (N_3265,N_3162,N_3121);
or U3266 (N_3266,N_3007,N_3172);
and U3267 (N_3267,N_3068,N_3141);
and U3268 (N_3268,N_3005,N_3107);
or U3269 (N_3269,N_3160,N_3191);
or U3270 (N_3270,N_3128,N_3018);
nand U3271 (N_3271,N_3035,N_3163);
nand U3272 (N_3272,N_3000,N_3118);
or U3273 (N_3273,N_3146,N_3175);
nor U3274 (N_3274,N_3051,N_3159);
nand U3275 (N_3275,N_3008,N_3064);
and U3276 (N_3276,N_3033,N_3032);
nor U3277 (N_3277,N_3169,N_3116);
or U3278 (N_3278,N_3050,N_3117);
and U3279 (N_3279,N_3076,N_3156);
or U3280 (N_3280,N_3063,N_3111);
or U3281 (N_3281,N_3144,N_3043);
nand U3282 (N_3282,N_3034,N_3185);
or U3283 (N_3283,N_3047,N_3145);
nor U3284 (N_3284,N_3101,N_3147);
nor U3285 (N_3285,N_3161,N_3151);
nor U3286 (N_3286,N_3016,N_3010);
and U3287 (N_3287,N_3149,N_3054);
nor U3288 (N_3288,N_3126,N_3055);
nand U3289 (N_3289,N_3129,N_3038);
xnor U3290 (N_3290,N_3095,N_3002);
and U3291 (N_3291,N_3040,N_3176);
and U3292 (N_3292,N_3039,N_3074);
and U3293 (N_3293,N_3075,N_3042);
nand U3294 (N_3294,N_3004,N_3157);
nand U3295 (N_3295,N_3127,N_3015);
or U3296 (N_3296,N_3192,N_3066);
and U3297 (N_3297,N_3106,N_3060);
xnor U3298 (N_3298,N_3011,N_3084);
nand U3299 (N_3299,N_3023,N_3093);
xnor U3300 (N_3300,N_3196,N_3101);
xor U3301 (N_3301,N_3065,N_3125);
or U3302 (N_3302,N_3108,N_3084);
xor U3303 (N_3303,N_3033,N_3000);
and U3304 (N_3304,N_3122,N_3044);
nand U3305 (N_3305,N_3136,N_3074);
and U3306 (N_3306,N_3128,N_3082);
nand U3307 (N_3307,N_3177,N_3168);
nor U3308 (N_3308,N_3006,N_3041);
or U3309 (N_3309,N_3110,N_3087);
or U3310 (N_3310,N_3046,N_3189);
and U3311 (N_3311,N_3012,N_3119);
nor U3312 (N_3312,N_3173,N_3182);
xnor U3313 (N_3313,N_3186,N_3127);
and U3314 (N_3314,N_3032,N_3087);
xor U3315 (N_3315,N_3052,N_3083);
or U3316 (N_3316,N_3064,N_3025);
nand U3317 (N_3317,N_3080,N_3021);
nand U3318 (N_3318,N_3064,N_3041);
nor U3319 (N_3319,N_3144,N_3195);
nor U3320 (N_3320,N_3012,N_3150);
or U3321 (N_3321,N_3127,N_3181);
nand U3322 (N_3322,N_3161,N_3092);
and U3323 (N_3323,N_3074,N_3132);
nor U3324 (N_3324,N_3064,N_3114);
xnor U3325 (N_3325,N_3166,N_3105);
and U3326 (N_3326,N_3176,N_3086);
nor U3327 (N_3327,N_3134,N_3115);
or U3328 (N_3328,N_3026,N_3049);
or U3329 (N_3329,N_3014,N_3082);
or U3330 (N_3330,N_3126,N_3194);
nor U3331 (N_3331,N_3006,N_3190);
or U3332 (N_3332,N_3096,N_3011);
nand U3333 (N_3333,N_3135,N_3136);
nand U3334 (N_3334,N_3033,N_3138);
or U3335 (N_3335,N_3141,N_3185);
or U3336 (N_3336,N_3189,N_3113);
xnor U3337 (N_3337,N_3152,N_3038);
or U3338 (N_3338,N_3127,N_3128);
nand U3339 (N_3339,N_3025,N_3063);
nor U3340 (N_3340,N_3056,N_3171);
nor U3341 (N_3341,N_3162,N_3166);
nand U3342 (N_3342,N_3091,N_3197);
nand U3343 (N_3343,N_3002,N_3091);
and U3344 (N_3344,N_3003,N_3054);
and U3345 (N_3345,N_3038,N_3080);
nor U3346 (N_3346,N_3100,N_3073);
nand U3347 (N_3347,N_3115,N_3192);
nor U3348 (N_3348,N_3115,N_3147);
and U3349 (N_3349,N_3042,N_3056);
nand U3350 (N_3350,N_3062,N_3180);
nand U3351 (N_3351,N_3179,N_3011);
and U3352 (N_3352,N_3185,N_3100);
nand U3353 (N_3353,N_3049,N_3013);
or U3354 (N_3354,N_3132,N_3053);
or U3355 (N_3355,N_3042,N_3124);
and U3356 (N_3356,N_3034,N_3143);
and U3357 (N_3357,N_3149,N_3007);
nand U3358 (N_3358,N_3118,N_3134);
and U3359 (N_3359,N_3076,N_3019);
and U3360 (N_3360,N_3093,N_3187);
and U3361 (N_3361,N_3184,N_3020);
nand U3362 (N_3362,N_3073,N_3146);
or U3363 (N_3363,N_3149,N_3064);
nand U3364 (N_3364,N_3071,N_3189);
xnor U3365 (N_3365,N_3042,N_3156);
and U3366 (N_3366,N_3012,N_3189);
or U3367 (N_3367,N_3170,N_3078);
xor U3368 (N_3368,N_3029,N_3049);
xnor U3369 (N_3369,N_3054,N_3050);
or U3370 (N_3370,N_3186,N_3060);
nor U3371 (N_3371,N_3154,N_3116);
nand U3372 (N_3372,N_3029,N_3042);
nor U3373 (N_3373,N_3022,N_3132);
and U3374 (N_3374,N_3190,N_3164);
nor U3375 (N_3375,N_3141,N_3026);
nand U3376 (N_3376,N_3056,N_3086);
nor U3377 (N_3377,N_3109,N_3195);
nor U3378 (N_3378,N_3154,N_3000);
nand U3379 (N_3379,N_3146,N_3115);
nor U3380 (N_3380,N_3164,N_3005);
and U3381 (N_3381,N_3144,N_3080);
and U3382 (N_3382,N_3187,N_3131);
or U3383 (N_3383,N_3093,N_3140);
nand U3384 (N_3384,N_3146,N_3195);
or U3385 (N_3385,N_3102,N_3041);
nor U3386 (N_3386,N_3022,N_3112);
or U3387 (N_3387,N_3059,N_3045);
nor U3388 (N_3388,N_3152,N_3102);
or U3389 (N_3389,N_3139,N_3163);
nor U3390 (N_3390,N_3048,N_3198);
nand U3391 (N_3391,N_3046,N_3099);
nor U3392 (N_3392,N_3047,N_3040);
nand U3393 (N_3393,N_3159,N_3021);
and U3394 (N_3394,N_3068,N_3095);
nor U3395 (N_3395,N_3055,N_3121);
xor U3396 (N_3396,N_3033,N_3065);
and U3397 (N_3397,N_3025,N_3004);
nand U3398 (N_3398,N_3037,N_3180);
and U3399 (N_3399,N_3144,N_3177);
nand U3400 (N_3400,N_3306,N_3227);
nand U3401 (N_3401,N_3290,N_3216);
nor U3402 (N_3402,N_3369,N_3389);
nand U3403 (N_3403,N_3336,N_3264);
nand U3404 (N_3404,N_3343,N_3209);
nor U3405 (N_3405,N_3329,N_3318);
nor U3406 (N_3406,N_3279,N_3355);
or U3407 (N_3407,N_3303,N_3297);
and U3408 (N_3408,N_3273,N_3339);
or U3409 (N_3409,N_3294,N_3392);
nor U3410 (N_3410,N_3348,N_3221);
nor U3411 (N_3411,N_3345,N_3344);
and U3412 (N_3412,N_3299,N_3352);
nor U3413 (N_3413,N_3338,N_3398);
nor U3414 (N_3414,N_3202,N_3287);
and U3415 (N_3415,N_3375,N_3214);
nor U3416 (N_3416,N_3206,N_3301);
or U3417 (N_3417,N_3249,N_3233);
nor U3418 (N_3418,N_3260,N_3263);
or U3419 (N_3419,N_3333,N_3374);
and U3420 (N_3420,N_3365,N_3331);
nand U3421 (N_3421,N_3208,N_3228);
nor U3422 (N_3422,N_3242,N_3342);
or U3423 (N_3423,N_3388,N_3218);
or U3424 (N_3424,N_3371,N_3212);
nand U3425 (N_3425,N_3222,N_3230);
nor U3426 (N_3426,N_3235,N_3312);
nand U3427 (N_3427,N_3321,N_3267);
or U3428 (N_3428,N_3243,N_3391);
nand U3429 (N_3429,N_3353,N_3223);
xnor U3430 (N_3430,N_3354,N_3236);
or U3431 (N_3431,N_3275,N_3272);
and U3432 (N_3432,N_3368,N_3281);
and U3433 (N_3433,N_3350,N_3237);
and U3434 (N_3434,N_3399,N_3386);
and U3435 (N_3435,N_3238,N_3325);
and U3436 (N_3436,N_3359,N_3319);
or U3437 (N_3437,N_3362,N_3284);
nand U3438 (N_3438,N_3364,N_3349);
nor U3439 (N_3439,N_3367,N_3360);
and U3440 (N_3440,N_3200,N_3324);
and U3441 (N_3441,N_3278,N_3385);
nor U3442 (N_3442,N_3314,N_3210);
nor U3443 (N_3443,N_3397,N_3395);
nand U3444 (N_3444,N_3327,N_3320);
or U3445 (N_3445,N_3255,N_3310);
nor U3446 (N_3446,N_3302,N_3335);
nand U3447 (N_3447,N_3373,N_3358);
and U3448 (N_3448,N_3363,N_3239);
or U3449 (N_3449,N_3265,N_3381);
nand U3450 (N_3450,N_3262,N_3213);
or U3451 (N_3451,N_3293,N_3271);
and U3452 (N_3452,N_3309,N_3288);
and U3453 (N_3453,N_3308,N_3207);
nand U3454 (N_3454,N_3316,N_3323);
and U3455 (N_3455,N_3337,N_3377);
and U3456 (N_3456,N_3383,N_3311);
nand U3457 (N_3457,N_3245,N_3322);
or U3458 (N_3458,N_3250,N_3231);
or U3459 (N_3459,N_3379,N_3387);
nor U3460 (N_3460,N_3292,N_3240);
nor U3461 (N_3461,N_3330,N_3246);
nand U3462 (N_3462,N_3347,N_3219);
nor U3463 (N_3463,N_3285,N_3346);
nand U3464 (N_3464,N_3384,N_3203);
nand U3465 (N_3465,N_3226,N_3296);
and U3466 (N_3466,N_3276,N_3282);
nand U3467 (N_3467,N_3201,N_3370);
and U3468 (N_3468,N_3215,N_3225);
nand U3469 (N_3469,N_3289,N_3378);
and U3470 (N_3470,N_3291,N_3286);
and U3471 (N_3471,N_3252,N_3205);
nor U3472 (N_3472,N_3253,N_3328);
xor U3473 (N_3473,N_3351,N_3270);
or U3474 (N_3474,N_3393,N_3247);
or U3475 (N_3475,N_3341,N_3251);
or U3476 (N_3476,N_3266,N_3241);
or U3477 (N_3477,N_3300,N_3256);
nor U3478 (N_3478,N_3356,N_3298);
nor U3479 (N_3479,N_3269,N_3244);
nand U3480 (N_3480,N_3396,N_3234);
and U3481 (N_3481,N_3382,N_3332);
nor U3482 (N_3482,N_3357,N_3394);
nor U3483 (N_3483,N_3274,N_3261);
nor U3484 (N_3484,N_3305,N_3390);
nor U3485 (N_3485,N_3258,N_3340);
nand U3486 (N_3486,N_3268,N_3277);
or U3487 (N_3487,N_3257,N_3224);
and U3488 (N_3488,N_3204,N_3307);
nand U3489 (N_3489,N_3315,N_3304);
or U3490 (N_3490,N_3254,N_3376);
xor U3491 (N_3491,N_3280,N_3361);
or U3492 (N_3492,N_3317,N_3326);
xnor U3493 (N_3493,N_3229,N_3248);
nand U3494 (N_3494,N_3295,N_3334);
xor U3495 (N_3495,N_3232,N_3366);
nand U3496 (N_3496,N_3372,N_3211);
nand U3497 (N_3497,N_3217,N_3380);
and U3498 (N_3498,N_3220,N_3313);
xor U3499 (N_3499,N_3259,N_3283);
or U3500 (N_3500,N_3201,N_3390);
xnor U3501 (N_3501,N_3327,N_3360);
nand U3502 (N_3502,N_3382,N_3267);
nand U3503 (N_3503,N_3247,N_3201);
and U3504 (N_3504,N_3313,N_3377);
nand U3505 (N_3505,N_3294,N_3353);
nor U3506 (N_3506,N_3297,N_3273);
nand U3507 (N_3507,N_3283,N_3331);
xor U3508 (N_3508,N_3374,N_3253);
and U3509 (N_3509,N_3339,N_3201);
or U3510 (N_3510,N_3257,N_3223);
nand U3511 (N_3511,N_3293,N_3338);
and U3512 (N_3512,N_3339,N_3343);
nand U3513 (N_3513,N_3298,N_3258);
or U3514 (N_3514,N_3287,N_3318);
nand U3515 (N_3515,N_3393,N_3322);
nand U3516 (N_3516,N_3321,N_3203);
and U3517 (N_3517,N_3392,N_3221);
or U3518 (N_3518,N_3276,N_3359);
nor U3519 (N_3519,N_3379,N_3209);
and U3520 (N_3520,N_3226,N_3337);
xor U3521 (N_3521,N_3281,N_3235);
or U3522 (N_3522,N_3395,N_3215);
nand U3523 (N_3523,N_3343,N_3346);
nand U3524 (N_3524,N_3293,N_3289);
nor U3525 (N_3525,N_3393,N_3366);
nor U3526 (N_3526,N_3287,N_3292);
and U3527 (N_3527,N_3376,N_3287);
nor U3528 (N_3528,N_3202,N_3277);
and U3529 (N_3529,N_3374,N_3239);
nor U3530 (N_3530,N_3376,N_3205);
or U3531 (N_3531,N_3260,N_3269);
nor U3532 (N_3532,N_3261,N_3212);
and U3533 (N_3533,N_3258,N_3391);
or U3534 (N_3534,N_3215,N_3350);
nor U3535 (N_3535,N_3286,N_3231);
xor U3536 (N_3536,N_3205,N_3307);
xor U3537 (N_3537,N_3258,N_3315);
nor U3538 (N_3538,N_3311,N_3298);
nor U3539 (N_3539,N_3283,N_3267);
nor U3540 (N_3540,N_3269,N_3281);
xor U3541 (N_3541,N_3368,N_3312);
and U3542 (N_3542,N_3295,N_3280);
and U3543 (N_3543,N_3329,N_3357);
or U3544 (N_3544,N_3339,N_3223);
or U3545 (N_3545,N_3231,N_3279);
nand U3546 (N_3546,N_3209,N_3345);
xnor U3547 (N_3547,N_3205,N_3361);
nor U3548 (N_3548,N_3354,N_3367);
xnor U3549 (N_3549,N_3290,N_3248);
and U3550 (N_3550,N_3363,N_3248);
nor U3551 (N_3551,N_3216,N_3375);
or U3552 (N_3552,N_3241,N_3323);
nor U3553 (N_3553,N_3327,N_3392);
or U3554 (N_3554,N_3307,N_3381);
nand U3555 (N_3555,N_3266,N_3344);
nor U3556 (N_3556,N_3276,N_3366);
nand U3557 (N_3557,N_3245,N_3324);
nor U3558 (N_3558,N_3318,N_3301);
nor U3559 (N_3559,N_3340,N_3240);
and U3560 (N_3560,N_3329,N_3326);
nor U3561 (N_3561,N_3348,N_3327);
or U3562 (N_3562,N_3374,N_3323);
or U3563 (N_3563,N_3342,N_3275);
nor U3564 (N_3564,N_3233,N_3306);
nand U3565 (N_3565,N_3335,N_3380);
nor U3566 (N_3566,N_3288,N_3217);
or U3567 (N_3567,N_3325,N_3331);
and U3568 (N_3568,N_3330,N_3253);
nor U3569 (N_3569,N_3211,N_3271);
or U3570 (N_3570,N_3294,N_3334);
nor U3571 (N_3571,N_3270,N_3322);
nor U3572 (N_3572,N_3299,N_3264);
and U3573 (N_3573,N_3296,N_3267);
or U3574 (N_3574,N_3363,N_3207);
or U3575 (N_3575,N_3287,N_3290);
nand U3576 (N_3576,N_3309,N_3241);
nor U3577 (N_3577,N_3288,N_3280);
or U3578 (N_3578,N_3207,N_3373);
or U3579 (N_3579,N_3306,N_3364);
or U3580 (N_3580,N_3245,N_3330);
nor U3581 (N_3581,N_3220,N_3361);
and U3582 (N_3582,N_3358,N_3203);
nor U3583 (N_3583,N_3324,N_3352);
xnor U3584 (N_3584,N_3259,N_3394);
xor U3585 (N_3585,N_3391,N_3216);
or U3586 (N_3586,N_3336,N_3235);
or U3587 (N_3587,N_3251,N_3358);
nand U3588 (N_3588,N_3226,N_3230);
nand U3589 (N_3589,N_3219,N_3369);
or U3590 (N_3590,N_3288,N_3353);
nand U3591 (N_3591,N_3306,N_3230);
nor U3592 (N_3592,N_3213,N_3236);
or U3593 (N_3593,N_3274,N_3361);
or U3594 (N_3594,N_3375,N_3221);
and U3595 (N_3595,N_3258,N_3347);
nand U3596 (N_3596,N_3374,N_3317);
or U3597 (N_3597,N_3204,N_3332);
nand U3598 (N_3598,N_3293,N_3209);
or U3599 (N_3599,N_3299,N_3271);
nand U3600 (N_3600,N_3436,N_3542);
or U3601 (N_3601,N_3512,N_3441);
or U3602 (N_3602,N_3539,N_3432);
and U3603 (N_3603,N_3556,N_3427);
xnor U3604 (N_3604,N_3507,N_3494);
nand U3605 (N_3605,N_3425,N_3469);
xnor U3606 (N_3606,N_3531,N_3574);
and U3607 (N_3607,N_3440,N_3503);
nor U3608 (N_3608,N_3578,N_3567);
or U3609 (N_3609,N_3497,N_3499);
and U3610 (N_3610,N_3589,N_3517);
nor U3611 (N_3611,N_3423,N_3478);
nor U3612 (N_3612,N_3446,N_3546);
nor U3613 (N_3613,N_3450,N_3487);
nand U3614 (N_3614,N_3411,N_3434);
and U3615 (N_3615,N_3513,N_3516);
nor U3616 (N_3616,N_3420,N_3493);
nor U3617 (N_3617,N_3460,N_3581);
or U3618 (N_3618,N_3518,N_3476);
or U3619 (N_3619,N_3575,N_3596);
xor U3620 (N_3620,N_3402,N_3551);
xnor U3621 (N_3621,N_3412,N_3569);
and U3622 (N_3622,N_3571,N_3439);
or U3623 (N_3623,N_3520,N_3501);
or U3624 (N_3624,N_3403,N_3552);
nor U3625 (N_3625,N_3470,N_3593);
nand U3626 (N_3626,N_3522,N_3413);
or U3627 (N_3627,N_3532,N_3481);
and U3628 (N_3628,N_3486,N_3442);
and U3629 (N_3629,N_3489,N_3484);
nand U3630 (N_3630,N_3594,N_3409);
and U3631 (N_3631,N_3563,N_3529);
nand U3632 (N_3632,N_3406,N_3428);
xnor U3633 (N_3633,N_3500,N_3421);
nor U3634 (N_3634,N_3566,N_3465);
nand U3635 (N_3635,N_3579,N_3416);
and U3636 (N_3636,N_3467,N_3472);
nand U3637 (N_3637,N_3521,N_3457);
and U3638 (N_3638,N_3570,N_3559);
and U3639 (N_3639,N_3536,N_3519);
nor U3640 (N_3640,N_3400,N_3414);
and U3641 (N_3641,N_3550,N_3491);
nor U3642 (N_3642,N_3495,N_3514);
nand U3643 (N_3643,N_3511,N_3561);
xor U3644 (N_3644,N_3463,N_3528);
nand U3645 (N_3645,N_3419,N_3431);
nand U3646 (N_3646,N_3525,N_3451);
nor U3647 (N_3647,N_3498,N_3461);
nor U3648 (N_3648,N_3454,N_3543);
nand U3649 (N_3649,N_3558,N_3568);
nor U3650 (N_3650,N_3417,N_3599);
nor U3651 (N_3651,N_3438,N_3549);
xnor U3652 (N_3652,N_3401,N_3523);
and U3653 (N_3653,N_3560,N_3557);
nor U3654 (N_3654,N_3537,N_3535);
nor U3655 (N_3655,N_3429,N_3591);
nand U3656 (N_3656,N_3508,N_3488);
nor U3657 (N_3657,N_3505,N_3464);
nor U3658 (N_3658,N_3527,N_3443);
nor U3659 (N_3659,N_3598,N_3584);
or U3660 (N_3660,N_3415,N_3405);
and U3661 (N_3661,N_3471,N_3453);
and U3662 (N_3662,N_3482,N_3477);
nand U3663 (N_3663,N_3466,N_3404);
nor U3664 (N_3664,N_3479,N_3506);
nand U3665 (N_3665,N_3510,N_3424);
nand U3666 (N_3666,N_3583,N_3435);
and U3667 (N_3667,N_3492,N_3562);
and U3668 (N_3668,N_3555,N_3509);
nand U3669 (N_3669,N_3496,N_3540);
and U3670 (N_3670,N_3545,N_3455);
nor U3671 (N_3671,N_3445,N_3585);
or U3672 (N_3672,N_3408,N_3504);
nand U3673 (N_3673,N_3418,N_3582);
nand U3674 (N_3674,N_3422,N_3553);
or U3675 (N_3675,N_3592,N_3586);
xnor U3676 (N_3676,N_3447,N_3480);
nor U3677 (N_3677,N_3433,N_3547);
or U3678 (N_3678,N_3452,N_3533);
and U3679 (N_3679,N_3524,N_3573);
nand U3680 (N_3680,N_3468,N_3597);
and U3681 (N_3681,N_3459,N_3534);
and U3682 (N_3682,N_3407,N_3448);
nor U3683 (N_3683,N_3538,N_3595);
or U3684 (N_3684,N_3473,N_3572);
nor U3685 (N_3685,N_3430,N_3515);
nand U3686 (N_3686,N_3530,N_3410);
and U3687 (N_3687,N_3426,N_3564);
nor U3688 (N_3688,N_3548,N_3588);
or U3689 (N_3689,N_3490,N_3485);
and U3690 (N_3690,N_3475,N_3456);
xor U3691 (N_3691,N_3437,N_3541);
and U3692 (N_3692,N_3544,N_3580);
xnor U3693 (N_3693,N_3554,N_3526);
nor U3694 (N_3694,N_3577,N_3565);
nor U3695 (N_3695,N_3502,N_3444);
nand U3696 (N_3696,N_3462,N_3590);
and U3697 (N_3697,N_3474,N_3449);
or U3698 (N_3698,N_3458,N_3587);
xnor U3699 (N_3699,N_3483,N_3576);
xnor U3700 (N_3700,N_3502,N_3529);
nand U3701 (N_3701,N_3569,N_3578);
and U3702 (N_3702,N_3456,N_3506);
or U3703 (N_3703,N_3475,N_3443);
or U3704 (N_3704,N_3545,N_3446);
xor U3705 (N_3705,N_3487,N_3468);
xnor U3706 (N_3706,N_3578,N_3414);
nand U3707 (N_3707,N_3506,N_3568);
nand U3708 (N_3708,N_3464,N_3521);
or U3709 (N_3709,N_3478,N_3532);
and U3710 (N_3710,N_3493,N_3566);
or U3711 (N_3711,N_3577,N_3416);
or U3712 (N_3712,N_3469,N_3574);
or U3713 (N_3713,N_3541,N_3430);
nor U3714 (N_3714,N_3411,N_3460);
or U3715 (N_3715,N_3411,N_3566);
and U3716 (N_3716,N_3568,N_3452);
nor U3717 (N_3717,N_3574,N_3550);
nor U3718 (N_3718,N_3525,N_3463);
nand U3719 (N_3719,N_3446,N_3591);
nand U3720 (N_3720,N_3403,N_3451);
xor U3721 (N_3721,N_3535,N_3444);
xor U3722 (N_3722,N_3480,N_3523);
nor U3723 (N_3723,N_3448,N_3528);
nor U3724 (N_3724,N_3561,N_3473);
or U3725 (N_3725,N_3511,N_3576);
or U3726 (N_3726,N_3417,N_3595);
xor U3727 (N_3727,N_3476,N_3496);
or U3728 (N_3728,N_3452,N_3583);
nand U3729 (N_3729,N_3476,N_3503);
nand U3730 (N_3730,N_3405,N_3555);
and U3731 (N_3731,N_3474,N_3594);
nand U3732 (N_3732,N_3414,N_3598);
nand U3733 (N_3733,N_3470,N_3474);
and U3734 (N_3734,N_3417,N_3455);
nand U3735 (N_3735,N_3409,N_3565);
and U3736 (N_3736,N_3496,N_3576);
and U3737 (N_3737,N_3446,N_3406);
nand U3738 (N_3738,N_3581,N_3406);
nor U3739 (N_3739,N_3555,N_3469);
and U3740 (N_3740,N_3516,N_3453);
or U3741 (N_3741,N_3459,N_3549);
and U3742 (N_3742,N_3480,N_3491);
nor U3743 (N_3743,N_3452,N_3477);
or U3744 (N_3744,N_3504,N_3578);
nand U3745 (N_3745,N_3488,N_3413);
nand U3746 (N_3746,N_3400,N_3553);
and U3747 (N_3747,N_3580,N_3437);
nand U3748 (N_3748,N_3582,N_3532);
nor U3749 (N_3749,N_3453,N_3408);
and U3750 (N_3750,N_3593,N_3419);
nor U3751 (N_3751,N_3523,N_3482);
or U3752 (N_3752,N_3442,N_3531);
and U3753 (N_3753,N_3557,N_3554);
and U3754 (N_3754,N_3544,N_3462);
nand U3755 (N_3755,N_3486,N_3566);
nand U3756 (N_3756,N_3551,N_3569);
nand U3757 (N_3757,N_3446,N_3566);
nand U3758 (N_3758,N_3504,N_3593);
nand U3759 (N_3759,N_3509,N_3520);
or U3760 (N_3760,N_3551,N_3428);
nand U3761 (N_3761,N_3453,N_3466);
xor U3762 (N_3762,N_3441,N_3403);
or U3763 (N_3763,N_3494,N_3560);
nor U3764 (N_3764,N_3445,N_3415);
nor U3765 (N_3765,N_3512,N_3481);
nor U3766 (N_3766,N_3592,N_3421);
nor U3767 (N_3767,N_3549,N_3547);
nor U3768 (N_3768,N_3579,N_3589);
nand U3769 (N_3769,N_3448,N_3465);
nor U3770 (N_3770,N_3546,N_3581);
nor U3771 (N_3771,N_3462,N_3481);
nor U3772 (N_3772,N_3442,N_3427);
or U3773 (N_3773,N_3549,N_3491);
and U3774 (N_3774,N_3567,N_3511);
and U3775 (N_3775,N_3590,N_3571);
nand U3776 (N_3776,N_3587,N_3429);
nor U3777 (N_3777,N_3576,N_3527);
nor U3778 (N_3778,N_3513,N_3471);
and U3779 (N_3779,N_3584,N_3475);
nand U3780 (N_3780,N_3514,N_3576);
or U3781 (N_3781,N_3470,N_3426);
and U3782 (N_3782,N_3560,N_3545);
and U3783 (N_3783,N_3427,N_3455);
nand U3784 (N_3784,N_3467,N_3417);
and U3785 (N_3785,N_3503,N_3416);
or U3786 (N_3786,N_3479,N_3469);
xnor U3787 (N_3787,N_3559,N_3499);
nand U3788 (N_3788,N_3488,N_3422);
xor U3789 (N_3789,N_3545,N_3511);
or U3790 (N_3790,N_3441,N_3549);
and U3791 (N_3791,N_3471,N_3511);
nand U3792 (N_3792,N_3561,N_3407);
and U3793 (N_3793,N_3581,N_3466);
nor U3794 (N_3794,N_3566,N_3423);
and U3795 (N_3795,N_3560,N_3475);
xor U3796 (N_3796,N_3587,N_3566);
nor U3797 (N_3797,N_3463,N_3535);
nand U3798 (N_3798,N_3533,N_3416);
and U3799 (N_3799,N_3538,N_3592);
or U3800 (N_3800,N_3773,N_3720);
or U3801 (N_3801,N_3629,N_3618);
or U3802 (N_3802,N_3734,N_3605);
and U3803 (N_3803,N_3779,N_3755);
nor U3804 (N_3804,N_3692,N_3751);
nand U3805 (N_3805,N_3765,N_3694);
and U3806 (N_3806,N_3680,N_3706);
nor U3807 (N_3807,N_3645,N_3601);
or U3808 (N_3808,N_3620,N_3619);
nor U3809 (N_3809,N_3721,N_3713);
or U3810 (N_3810,N_3639,N_3738);
nand U3811 (N_3811,N_3743,N_3678);
xnor U3812 (N_3812,N_3625,N_3776);
nor U3813 (N_3813,N_3780,N_3668);
and U3814 (N_3814,N_3607,N_3650);
nand U3815 (N_3815,N_3675,N_3715);
or U3816 (N_3816,N_3689,N_3770);
nand U3817 (N_3817,N_3700,N_3719);
nor U3818 (N_3818,N_3767,N_3774);
and U3819 (N_3819,N_3617,N_3728);
nor U3820 (N_3820,N_3695,N_3760);
nand U3821 (N_3821,N_3624,N_3753);
nor U3822 (N_3822,N_3792,N_3679);
nand U3823 (N_3823,N_3662,N_3641);
or U3824 (N_3824,N_3615,N_3756);
and U3825 (N_3825,N_3784,N_3637);
xor U3826 (N_3826,N_3798,N_3785);
or U3827 (N_3827,N_3712,N_3766);
nor U3828 (N_3828,N_3684,N_3772);
and U3829 (N_3829,N_3777,N_3663);
nand U3830 (N_3830,N_3793,N_3718);
nor U3831 (N_3831,N_3716,N_3795);
nand U3832 (N_3832,N_3748,N_3652);
nand U3833 (N_3833,N_3616,N_3758);
xnor U3834 (N_3834,N_3705,N_3764);
nor U3835 (N_3835,N_3640,N_3646);
or U3836 (N_3836,N_3672,N_3649);
or U3837 (N_3837,N_3763,N_3782);
and U3838 (N_3838,N_3709,N_3606);
nor U3839 (N_3839,N_3653,N_3697);
nor U3840 (N_3840,N_3744,N_3673);
and U3841 (N_3841,N_3769,N_3703);
or U3842 (N_3842,N_3740,N_3790);
xnor U3843 (N_3843,N_3724,N_3600);
or U3844 (N_3844,N_3690,N_3737);
nor U3845 (N_3845,N_3656,N_3741);
nor U3846 (N_3846,N_3754,N_3685);
or U3847 (N_3847,N_3632,N_3613);
or U3848 (N_3848,N_3608,N_3638);
and U3849 (N_3849,N_3723,N_3621);
nand U3850 (N_3850,N_3627,N_3686);
xor U3851 (N_3851,N_3768,N_3670);
or U3852 (N_3852,N_3603,N_3749);
and U3853 (N_3853,N_3671,N_3722);
or U3854 (N_3854,N_3711,N_3794);
nand U3855 (N_3855,N_3628,N_3714);
nand U3856 (N_3856,N_3698,N_3666);
or U3857 (N_3857,N_3702,N_3732);
or U3858 (N_3858,N_3726,N_3664);
and U3859 (N_3859,N_3696,N_3750);
nand U3860 (N_3860,N_3677,N_3704);
nor U3861 (N_3861,N_3659,N_3701);
or U3862 (N_3862,N_3717,N_3682);
nor U3863 (N_3863,N_3791,N_3727);
nand U3864 (N_3864,N_3759,N_3742);
nand U3865 (N_3865,N_3746,N_3636);
nand U3866 (N_3866,N_3681,N_3655);
nor U3867 (N_3867,N_3783,N_3731);
or U3868 (N_3868,N_3658,N_3611);
and U3869 (N_3869,N_3683,N_3623);
nand U3870 (N_3870,N_3604,N_3693);
or U3871 (N_3871,N_3687,N_3739);
and U3872 (N_3872,N_3661,N_3725);
or U3873 (N_3873,N_3778,N_3797);
nand U3874 (N_3874,N_3635,N_3612);
or U3875 (N_3875,N_3633,N_3752);
xnor U3876 (N_3876,N_3762,N_3651);
or U3877 (N_3877,N_3642,N_3781);
and U3878 (N_3878,N_3609,N_3699);
and U3879 (N_3879,N_3626,N_3799);
nand U3880 (N_3880,N_3775,N_3657);
or U3881 (N_3881,N_3710,N_3735);
and U3882 (N_3882,N_3665,N_3648);
nor U3883 (N_3883,N_3631,N_3708);
nand U3884 (N_3884,N_3736,N_3634);
nand U3885 (N_3885,N_3669,N_3788);
nor U3886 (N_3886,N_3787,N_3733);
nand U3887 (N_3887,N_3667,N_3761);
nor U3888 (N_3888,N_3691,N_3771);
xor U3889 (N_3889,N_3602,N_3757);
or U3890 (N_3890,N_3614,N_3610);
or U3891 (N_3891,N_3676,N_3630);
nor U3892 (N_3892,N_3688,N_3660);
nor U3893 (N_3893,N_3789,N_3747);
nand U3894 (N_3894,N_3643,N_3674);
nand U3895 (N_3895,N_3647,N_3707);
or U3896 (N_3896,N_3786,N_3745);
nor U3897 (N_3897,N_3644,N_3796);
xor U3898 (N_3898,N_3730,N_3622);
and U3899 (N_3899,N_3654,N_3729);
or U3900 (N_3900,N_3786,N_3727);
and U3901 (N_3901,N_3743,N_3648);
nor U3902 (N_3902,N_3661,N_3677);
nand U3903 (N_3903,N_3636,N_3797);
nand U3904 (N_3904,N_3683,N_3740);
nor U3905 (N_3905,N_3607,N_3710);
and U3906 (N_3906,N_3724,N_3699);
and U3907 (N_3907,N_3701,N_3657);
or U3908 (N_3908,N_3649,N_3647);
nand U3909 (N_3909,N_3777,N_3711);
xnor U3910 (N_3910,N_3675,N_3693);
nor U3911 (N_3911,N_3664,N_3735);
nand U3912 (N_3912,N_3737,N_3745);
nand U3913 (N_3913,N_3756,N_3668);
and U3914 (N_3914,N_3795,N_3714);
nor U3915 (N_3915,N_3777,N_3644);
or U3916 (N_3916,N_3682,N_3683);
nor U3917 (N_3917,N_3760,N_3675);
nor U3918 (N_3918,N_3772,N_3765);
or U3919 (N_3919,N_3688,N_3744);
or U3920 (N_3920,N_3795,N_3718);
nand U3921 (N_3921,N_3680,N_3640);
or U3922 (N_3922,N_3701,N_3784);
and U3923 (N_3923,N_3619,N_3634);
nand U3924 (N_3924,N_3700,N_3704);
nor U3925 (N_3925,N_3756,N_3626);
and U3926 (N_3926,N_3700,N_3753);
and U3927 (N_3927,N_3696,N_3710);
or U3928 (N_3928,N_3788,N_3739);
or U3929 (N_3929,N_3623,N_3757);
or U3930 (N_3930,N_3627,N_3793);
nor U3931 (N_3931,N_3635,N_3692);
nor U3932 (N_3932,N_3643,N_3640);
nand U3933 (N_3933,N_3764,N_3621);
xor U3934 (N_3934,N_3744,N_3629);
nor U3935 (N_3935,N_3757,N_3790);
nand U3936 (N_3936,N_3629,N_3630);
nand U3937 (N_3937,N_3613,N_3642);
or U3938 (N_3938,N_3661,N_3678);
nor U3939 (N_3939,N_3742,N_3647);
or U3940 (N_3940,N_3648,N_3760);
and U3941 (N_3941,N_3793,N_3738);
xnor U3942 (N_3942,N_3761,N_3798);
nand U3943 (N_3943,N_3792,N_3734);
and U3944 (N_3944,N_3691,N_3714);
and U3945 (N_3945,N_3665,N_3664);
nand U3946 (N_3946,N_3688,N_3661);
and U3947 (N_3947,N_3678,N_3702);
or U3948 (N_3948,N_3715,N_3603);
nand U3949 (N_3949,N_3683,N_3727);
nand U3950 (N_3950,N_3695,N_3787);
and U3951 (N_3951,N_3771,N_3693);
nor U3952 (N_3952,N_3793,N_3602);
and U3953 (N_3953,N_3660,N_3755);
or U3954 (N_3954,N_3733,N_3619);
nor U3955 (N_3955,N_3765,N_3666);
nand U3956 (N_3956,N_3610,N_3796);
nand U3957 (N_3957,N_3751,N_3700);
nor U3958 (N_3958,N_3780,N_3689);
or U3959 (N_3959,N_3775,N_3642);
nand U3960 (N_3960,N_3713,N_3724);
and U3961 (N_3961,N_3685,N_3759);
and U3962 (N_3962,N_3622,N_3657);
nand U3963 (N_3963,N_3741,N_3710);
xor U3964 (N_3964,N_3620,N_3688);
xnor U3965 (N_3965,N_3768,N_3616);
nand U3966 (N_3966,N_3611,N_3704);
nand U3967 (N_3967,N_3727,N_3701);
or U3968 (N_3968,N_3689,N_3624);
nor U3969 (N_3969,N_3634,N_3669);
nand U3970 (N_3970,N_3757,N_3646);
nand U3971 (N_3971,N_3652,N_3713);
and U3972 (N_3972,N_3665,N_3631);
xor U3973 (N_3973,N_3733,N_3625);
and U3974 (N_3974,N_3787,N_3669);
nor U3975 (N_3975,N_3774,N_3768);
nand U3976 (N_3976,N_3676,N_3719);
nand U3977 (N_3977,N_3616,N_3780);
nor U3978 (N_3978,N_3672,N_3618);
or U3979 (N_3979,N_3701,N_3700);
nor U3980 (N_3980,N_3656,N_3758);
and U3981 (N_3981,N_3782,N_3747);
and U3982 (N_3982,N_3647,N_3656);
nand U3983 (N_3983,N_3751,N_3670);
and U3984 (N_3984,N_3735,N_3665);
or U3985 (N_3985,N_3792,N_3643);
nor U3986 (N_3986,N_3696,N_3793);
nor U3987 (N_3987,N_3680,N_3638);
and U3988 (N_3988,N_3781,N_3783);
xor U3989 (N_3989,N_3703,N_3654);
xnor U3990 (N_3990,N_3698,N_3646);
nor U3991 (N_3991,N_3694,N_3712);
and U3992 (N_3992,N_3703,N_3723);
or U3993 (N_3993,N_3783,N_3669);
nand U3994 (N_3994,N_3720,N_3780);
or U3995 (N_3995,N_3660,N_3796);
and U3996 (N_3996,N_3639,N_3712);
or U3997 (N_3997,N_3694,N_3633);
or U3998 (N_3998,N_3710,N_3684);
nand U3999 (N_3999,N_3692,N_3655);
and U4000 (N_4000,N_3829,N_3922);
nor U4001 (N_4001,N_3896,N_3988);
nor U4002 (N_4002,N_3886,N_3912);
and U4003 (N_4003,N_3814,N_3889);
and U4004 (N_4004,N_3946,N_3810);
or U4005 (N_4005,N_3824,N_3813);
nand U4006 (N_4006,N_3854,N_3942);
or U4007 (N_4007,N_3973,N_3866);
and U4008 (N_4008,N_3858,N_3982);
or U4009 (N_4009,N_3938,N_3803);
and U4010 (N_4010,N_3885,N_3914);
or U4011 (N_4011,N_3978,N_3871);
or U4012 (N_4012,N_3873,N_3997);
nor U4013 (N_4013,N_3985,N_3940);
nand U4014 (N_4014,N_3860,N_3848);
or U4015 (N_4015,N_3881,N_3929);
or U4016 (N_4016,N_3899,N_3840);
nand U4017 (N_4017,N_3882,N_3880);
nor U4018 (N_4018,N_3838,N_3841);
nor U4019 (N_4019,N_3987,N_3927);
nand U4020 (N_4020,N_3844,N_3893);
or U4021 (N_4021,N_3977,N_3902);
nand U4022 (N_4022,N_3924,N_3937);
nand U4023 (N_4023,N_3801,N_3864);
nor U4024 (N_4024,N_3976,N_3818);
and U4025 (N_4025,N_3898,N_3846);
nand U4026 (N_4026,N_3925,N_3996);
nor U4027 (N_4027,N_3954,N_3990);
xnor U4028 (N_4028,N_3883,N_3943);
nand U4029 (N_4029,N_3835,N_3804);
xor U4030 (N_4030,N_3931,N_3830);
or U4031 (N_4031,N_3932,N_3939);
and U4032 (N_4032,N_3822,N_3984);
and U4033 (N_4033,N_3934,N_3811);
and U4034 (N_4034,N_3979,N_3888);
nor U4035 (N_4035,N_3819,N_3917);
nand U4036 (N_4036,N_3855,N_3923);
and U4037 (N_4037,N_3817,N_3843);
xor U4038 (N_4038,N_3870,N_3849);
nor U4039 (N_4039,N_3809,N_3834);
or U4040 (N_4040,N_3933,N_3981);
or U4041 (N_4041,N_3930,N_3832);
xnor U4042 (N_4042,N_3968,N_3936);
nand U4043 (N_4043,N_3994,N_3874);
nor U4044 (N_4044,N_3993,N_3891);
or U4045 (N_4045,N_3957,N_3837);
nand U4046 (N_4046,N_3862,N_3913);
xor U4047 (N_4047,N_3950,N_3876);
nand U4048 (N_4048,N_3851,N_3820);
nand U4049 (N_4049,N_3875,N_3825);
nor U4050 (N_4050,N_3836,N_3918);
and U4051 (N_4051,N_3958,N_3833);
nor U4052 (N_4052,N_3863,N_3872);
nand U4053 (N_4053,N_3907,N_3831);
and U4054 (N_4054,N_3948,N_3847);
nor U4055 (N_4055,N_3901,N_3903);
nor U4056 (N_4056,N_3869,N_3992);
nor U4057 (N_4057,N_3920,N_3800);
nand U4058 (N_4058,N_3900,N_3963);
and U4059 (N_4059,N_3850,N_3859);
or U4060 (N_4060,N_3964,N_3989);
xnor U4061 (N_4061,N_3951,N_3909);
nor U4062 (N_4062,N_3812,N_3944);
nor U4063 (N_4063,N_3919,N_3805);
or U4064 (N_4064,N_3975,N_3960);
and U4065 (N_4065,N_3906,N_3905);
nor U4066 (N_4066,N_3941,N_3953);
and U4067 (N_4067,N_3897,N_3956);
or U4068 (N_4068,N_3853,N_3865);
nor U4069 (N_4069,N_3845,N_3867);
or U4070 (N_4070,N_3887,N_3890);
or U4071 (N_4071,N_3856,N_3955);
nand U4072 (N_4072,N_3999,N_3969);
or U4073 (N_4073,N_3808,N_3971);
or U4074 (N_4074,N_3959,N_3879);
and U4075 (N_4075,N_3970,N_3892);
or U4076 (N_4076,N_3821,N_3823);
nor U4077 (N_4077,N_3911,N_3878);
or U4078 (N_4078,N_3842,N_3945);
or U4079 (N_4079,N_3949,N_3884);
nor U4080 (N_4080,N_3857,N_3962);
or U4081 (N_4081,N_3966,N_3998);
xnor U4082 (N_4082,N_3952,N_3828);
nand U4083 (N_4083,N_3965,N_3839);
nor U4084 (N_4084,N_3868,N_3995);
xor U4085 (N_4085,N_3972,N_3961);
nand U4086 (N_4086,N_3974,N_3947);
nand U4087 (N_4087,N_3806,N_3826);
or U4088 (N_4088,N_3802,N_3908);
and U4089 (N_4089,N_3928,N_3915);
nand U4090 (N_4090,N_3921,N_3827);
xor U4091 (N_4091,N_3935,N_3983);
and U4092 (N_4092,N_3894,N_3877);
and U4093 (N_4093,N_3910,N_3861);
and U4094 (N_4094,N_3916,N_3926);
and U4095 (N_4095,N_3852,N_3980);
and U4096 (N_4096,N_3967,N_3807);
or U4097 (N_4097,N_3904,N_3815);
and U4098 (N_4098,N_3895,N_3816);
nand U4099 (N_4099,N_3991,N_3986);
nand U4100 (N_4100,N_3886,N_3874);
nand U4101 (N_4101,N_3959,N_3813);
and U4102 (N_4102,N_3804,N_3890);
xor U4103 (N_4103,N_3962,N_3868);
or U4104 (N_4104,N_3802,N_3933);
or U4105 (N_4105,N_3964,N_3899);
and U4106 (N_4106,N_3956,N_3979);
and U4107 (N_4107,N_3881,N_3833);
or U4108 (N_4108,N_3825,N_3912);
nand U4109 (N_4109,N_3998,N_3805);
nand U4110 (N_4110,N_3817,N_3879);
or U4111 (N_4111,N_3905,N_3817);
nor U4112 (N_4112,N_3901,N_3942);
or U4113 (N_4113,N_3959,N_3859);
nor U4114 (N_4114,N_3943,N_3910);
or U4115 (N_4115,N_3874,N_3833);
or U4116 (N_4116,N_3852,N_3974);
nand U4117 (N_4117,N_3859,N_3995);
xor U4118 (N_4118,N_3890,N_3968);
or U4119 (N_4119,N_3803,N_3910);
nor U4120 (N_4120,N_3909,N_3919);
nand U4121 (N_4121,N_3975,N_3846);
nor U4122 (N_4122,N_3839,N_3963);
nand U4123 (N_4123,N_3908,N_3996);
nand U4124 (N_4124,N_3928,N_3980);
or U4125 (N_4125,N_3896,N_3926);
nor U4126 (N_4126,N_3906,N_3821);
or U4127 (N_4127,N_3914,N_3834);
and U4128 (N_4128,N_3861,N_3983);
and U4129 (N_4129,N_3942,N_3984);
or U4130 (N_4130,N_3844,N_3965);
nor U4131 (N_4131,N_3851,N_3927);
nor U4132 (N_4132,N_3864,N_3894);
nor U4133 (N_4133,N_3972,N_3958);
nor U4134 (N_4134,N_3993,N_3990);
nor U4135 (N_4135,N_3923,N_3915);
nor U4136 (N_4136,N_3934,N_3904);
or U4137 (N_4137,N_3912,N_3830);
and U4138 (N_4138,N_3883,N_3858);
nand U4139 (N_4139,N_3963,N_3933);
and U4140 (N_4140,N_3831,N_3939);
or U4141 (N_4141,N_3900,N_3879);
or U4142 (N_4142,N_3816,N_3887);
and U4143 (N_4143,N_3862,N_3802);
and U4144 (N_4144,N_3928,N_3927);
and U4145 (N_4145,N_3807,N_3836);
nor U4146 (N_4146,N_3998,N_3975);
xnor U4147 (N_4147,N_3827,N_3911);
nand U4148 (N_4148,N_3972,N_3966);
nor U4149 (N_4149,N_3929,N_3957);
or U4150 (N_4150,N_3853,N_3923);
nand U4151 (N_4151,N_3990,N_3983);
and U4152 (N_4152,N_3913,N_3880);
and U4153 (N_4153,N_3904,N_3807);
or U4154 (N_4154,N_3937,N_3886);
xnor U4155 (N_4155,N_3852,N_3992);
nor U4156 (N_4156,N_3980,N_3803);
and U4157 (N_4157,N_3950,N_3995);
xor U4158 (N_4158,N_3897,N_3851);
nor U4159 (N_4159,N_3887,N_3877);
nand U4160 (N_4160,N_3881,N_3854);
nor U4161 (N_4161,N_3876,N_3842);
xnor U4162 (N_4162,N_3944,N_3892);
and U4163 (N_4163,N_3946,N_3805);
nor U4164 (N_4164,N_3821,N_3900);
nand U4165 (N_4165,N_3998,N_3953);
or U4166 (N_4166,N_3971,N_3874);
nor U4167 (N_4167,N_3898,N_3951);
nand U4168 (N_4168,N_3956,N_3975);
nor U4169 (N_4169,N_3897,N_3884);
or U4170 (N_4170,N_3849,N_3846);
and U4171 (N_4171,N_3927,N_3986);
xnor U4172 (N_4172,N_3860,N_3875);
nor U4173 (N_4173,N_3826,N_3855);
or U4174 (N_4174,N_3884,N_3849);
and U4175 (N_4175,N_3963,N_3803);
nand U4176 (N_4176,N_3850,N_3986);
or U4177 (N_4177,N_3902,N_3975);
xor U4178 (N_4178,N_3894,N_3814);
nor U4179 (N_4179,N_3852,N_3932);
or U4180 (N_4180,N_3982,N_3843);
and U4181 (N_4181,N_3852,N_3910);
or U4182 (N_4182,N_3822,N_3923);
nand U4183 (N_4183,N_3872,N_3864);
nand U4184 (N_4184,N_3833,N_3937);
xor U4185 (N_4185,N_3993,N_3938);
xor U4186 (N_4186,N_3967,N_3852);
nor U4187 (N_4187,N_3966,N_3802);
or U4188 (N_4188,N_3895,N_3901);
nand U4189 (N_4189,N_3893,N_3837);
nor U4190 (N_4190,N_3898,N_3858);
or U4191 (N_4191,N_3877,N_3888);
or U4192 (N_4192,N_3983,N_3856);
and U4193 (N_4193,N_3981,N_3972);
or U4194 (N_4194,N_3970,N_3876);
or U4195 (N_4195,N_3887,N_3888);
nor U4196 (N_4196,N_3975,N_3806);
nand U4197 (N_4197,N_3956,N_3939);
nor U4198 (N_4198,N_3848,N_3969);
nor U4199 (N_4199,N_3862,N_3860);
nor U4200 (N_4200,N_4158,N_4095);
and U4201 (N_4201,N_4040,N_4101);
and U4202 (N_4202,N_4154,N_4003);
and U4203 (N_4203,N_4026,N_4093);
or U4204 (N_4204,N_4016,N_4060);
and U4205 (N_4205,N_4067,N_4122);
nor U4206 (N_4206,N_4028,N_4110);
nor U4207 (N_4207,N_4098,N_4164);
or U4208 (N_4208,N_4139,N_4001);
or U4209 (N_4209,N_4037,N_4163);
nand U4210 (N_4210,N_4054,N_4077);
nor U4211 (N_4211,N_4073,N_4050);
and U4212 (N_4212,N_4128,N_4052);
nand U4213 (N_4213,N_4057,N_4085);
or U4214 (N_4214,N_4083,N_4113);
nor U4215 (N_4215,N_4103,N_4051);
and U4216 (N_4216,N_4055,N_4120);
and U4217 (N_4217,N_4102,N_4109);
nor U4218 (N_4218,N_4081,N_4089);
nand U4219 (N_4219,N_4173,N_4127);
and U4220 (N_4220,N_4135,N_4141);
or U4221 (N_4221,N_4070,N_4167);
nand U4222 (N_4222,N_4086,N_4177);
and U4223 (N_4223,N_4180,N_4088);
nand U4224 (N_4224,N_4191,N_4025);
or U4225 (N_4225,N_4182,N_4186);
xnor U4226 (N_4226,N_4075,N_4157);
and U4227 (N_4227,N_4005,N_4034);
and U4228 (N_4228,N_4046,N_4129);
and U4229 (N_4229,N_4118,N_4045);
or U4230 (N_4230,N_4064,N_4043);
nand U4231 (N_4231,N_4160,N_4063);
xnor U4232 (N_4232,N_4197,N_4123);
or U4233 (N_4233,N_4195,N_4189);
nand U4234 (N_4234,N_4159,N_4148);
or U4235 (N_4235,N_4048,N_4008);
or U4236 (N_4236,N_4019,N_4074);
or U4237 (N_4237,N_4111,N_4017);
nor U4238 (N_4238,N_4092,N_4184);
and U4239 (N_4239,N_4169,N_4134);
nor U4240 (N_4240,N_4112,N_4150);
nand U4241 (N_4241,N_4143,N_4193);
nor U4242 (N_4242,N_4072,N_4030);
and U4243 (N_4243,N_4031,N_4176);
nand U4244 (N_4244,N_4115,N_4002);
and U4245 (N_4245,N_4145,N_4199);
nand U4246 (N_4246,N_4061,N_4059);
nand U4247 (N_4247,N_4185,N_4042);
or U4248 (N_4248,N_4170,N_4062);
nor U4249 (N_4249,N_4178,N_4079);
nor U4250 (N_4250,N_4172,N_4099);
nand U4251 (N_4251,N_4084,N_4187);
xnor U4252 (N_4252,N_4039,N_4151);
and U4253 (N_4253,N_4020,N_4027);
and U4254 (N_4254,N_4012,N_4024);
or U4255 (N_4255,N_4107,N_4010);
or U4256 (N_4256,N_4156,N_4144);
and U4257 (N_4257,N_4198,N_4011);
nand U4258 (N_4258,N_4142,N_4036);
nor U4259 (N_4259,N_4175,N_4021);
nor U4260 (N_4260,N_4125,N_4116);
and U4261 (N_4261,N_4058,N_4104);
or U4262 (N_4262,N_4004,N_4165);
nor U4263 (N_4263,N_4196,N_4090);
or U4264 (N_4264,N_4171,N_4168);
nand U4265 (N_4265,N_4138,N_4018);
nor U4266 (N_4266,N_4044,N_4194);
and U4267 (N_4267,N_4126,N_4078);
or U4268 (N_4268,N_4114,N_4162);
nand U4269 (N_4269,N_4119,N_4091);
and U4270 (N_4270,N_4032,N_4188);
and U4271 (N_4271,N_4068,N_4131);
nand U4272 (N_4272,N_4013,N_4097);
xor U4273 (N_4273,N_4009,N_4130);
nand U4274 (N_4274,N_4181,N_4035);
and U4275 (N_4275,N_4049,N_4015);
and U4276 (N_4276,N_4146,N_4183);
or U4277 (N_4277,N_4071,N_4137);
and U4278 (N_4278,N_4047,N_4080);
nor U4279 (N_4279,N_4149,N_4152);
nor U4280 (N_4280,N_4069,N_4174);
or U4281 (N_4281,N_4161,N_4147);
nor U4282 (N_4282,N_4056,N_4117);
or U4283 (N_4283,N_4041,N_4094);
nor U4284 (N_4284,N_4082,N_4105);
nor U4285 (N_4285,N_4000,N_4140);
and U4286 (N_4286,N_4053,N_4007);
or U4287 (N_4287,N_4029,N_4132);
nand U4288 (N_4288,N_4038,N_4033);
nand U4289 (N_4289,N_4190,N_4153);
nand U4290 (N_4290,N_4192,N_4166);
nand U4291 (N_4291,N_4133,N_4106);
nor U4292 (N_4292,N_4155,N_4066);
and U4293 (N_4293,N_4087,N_4108);
nor U4294 (N_4294,N_4100,N_4096);
nand U4295 (N_4295,N_4022,N_4124);
nand U4296 (N_4296,N_4136,N_4014);
nor U4297 (N_4297,N_4076,N_4023);
xor U4298 (N_4298,N_4006,N_4179);
and U4299 (N_4299,N_4121,N_4065);
xnor U4300 (N_4300,N_4183,N_4088);
nor U4301 (N_4301,N_4054,N_4139);
and U4302 (N_4302,N_4075,N_4145);
nand U4303 (N_4303,N_4106,N_4149);
and U4304 (N_4304,N_4193,N_4074);
and U4305 (N_4305,N_4183,N_4163);
nand U4306 (N_4306,N_4072,N_4124);
or U4307 (N_4307,N_4190,N_4041);
xor U4308 (N_4308,N_4080,N_4106);
nor U4309 (N_4309,N_4094,N_4071);
xor U4310 (N_4310,N_4010,N_4118);
and U4311 (N_4311,N_4136,N_4097);
and U4312 (N_4312,N_4015,N_4131);
nor U4313 (N_4313,N_4159,N_4092);
or U4314 (N_4314,N_4129,N_4197);
nand U4315 (N_4315,N_4126,N_4002);
and U4316 (N_4316,N_4115,N_4150);
nor U4317 (N_4317,N_4085,N_4181);
nor U4318 (N_4318,N_4100,N_4104);
and U4319 (N_4319,N_4176,N_4077);
nand U4320 (N_4320,N_4107,N_4030);
xnor U4321 (N_4321,N_4133,N_4104);
nand U4322 (N_4322,N_4109,N_4068);
nor U4323 (N_4323,N_4081,N_4147);
nand U4324 (N_4324,N_4186,N_4168);
nor U4325 (N_4325,N_4056,N_4122);
and U4326 (N_4326,N_4177,N_4002);
nand U4327 (N_4327,N_4011,N_4159);
or U4328 (N_4328,N_4183,N_4102);
and U4329 (N_4329,N_4003,N_4125);
or U4330 (N_4330,N_4151,N_4011);
and U4331 (N_4331,N_4177,N_4036);
and U4332 (N_4332,N_4110,N_4189);
and U4333 (N_4333,N_4184,N_4018);
nand U4334 (N_4334,N_4043,N_4186);
nor U4335 (N_4335,N_4182,N_4031);
or U4336 (N_4336,N_4127,N_4008);
nor U4337 (N_4337,N_4090,N_4095);
nand U4338 (N_4338,N_4161,N_4046);
nor U4339 (N_4339,N_4153,N_4034);
nor U4340 (N_4340,N_4197,N_4174);
or U4341 (N_4341,N_4092,N_4123);
xor U4342 (N_4342,N_4017,N_4142);
nor U4343 (N_4343,N_4034,N_4111);
xnor U4344 (N_4344,N_4088,N_4092);
nor U4345 (N_4345,N_4135,N_4192);
nand U4346 (N_4346,N_4192,N_4137);
and U4347 (N_4347,N_4116,N_4190);
nor U4348 (N_4348,N_4015,N_4176);
and U4349 (N_4349,N_4023,N_4059);
nor U4350 (N_4350,N_4050,N_4190);
and U4351 (N_4351,N_4055,N_4085);
nor U4352 (N_4352,N_4124,N_4102);
and U4353 (N_4353,N_4103,N_4042);
nand U4354 (N_4354,N_4103,N_4070);
nand U4355 (N_4355,N_4014,N_4074);
or U4356 (N_4356,N_4014,N_4025);
and U4357 (N_4357,N_4013,N_4088);
or U4358 (N_4358,N_4130,N_4155);
xor U4359 (N_4359,N_4121,N_4154);
nand U4360 (N_4360,N_4050,N_4051);
xor U4361 (N_4361,N_4002,N_4023);
nor U4362 (N_4362,N_4128,N_4177);
and U4363 (N_4363,N_4188,N_4170);
nand U4364 (N_4364,N_4056,N_4161);
and U4365 (N_4365,N_4120,N_4151);
nand U4366 (N_4366,N_4158,N_4140);
or U4367 (N_4367,N_4131,N_4107);
nor U4368 (N_4368,N_4126,N_4094);
and U4369 (N_4369,N_4168,N_4187);
and U4370 (N_4370,N_4079,N_4167);
and U4371 (N_4371,N_4113,N_4069);
and U4372 (N_4372,N_4121,N_4007);
and U4373 (N_4373,N_4067,N_4005);
nand U4374 (N_4374,N_4060,N_4138);
nand U4375 (N_4375,N_4196,N_4160);
and U4376 (N_4376,N_4041,N_4015);
and U4377 (N_4377,N_4174,N_4156);
and U4378 (N_4378,N_4118,N_4182);
nand U4379 (N_4379,N_4026,N_4191);
nand U4380 (N_4380,N_4027,N_4157);
or U4381 (N_4381,N_4090,N_4120);
nor U4382 (N_4382,N_4164,N_4060);
xnor U4383 (N_4383,N_4149,N_4176);
or U4384 (N_4384,N_4057,N_4168);
nand U4385 (N_4385,N_4080,N_4134);
nand U4386 (N_4386,N_4108,N_4046);
xnor U4387 (N_4387,N_4064,N_4004);
or U4388 (N_4388,N_4048,N_4076);
nor U4389 (N_4389,N_4112,N_4033);
and U4390 (N_4390,N_4101,N_4038);
nor U4391 (N_4391,N_4156,N_4027);
and U4392 (N_4392,N_4107,N_4051);
or U4393 (N_4393,N_4194,N_4038);
and U4394 (N_4394,N_4176,N_4119);
and U4395 (N_4395,N_4145,N_4138);
and U4396 (N_4396,N_4058,N_4099);
xnor U4397 (N_4397,N_4187,N_4005);
and U4398 (N_4398,N_4172,N_4160);
or U4399 (N_4399,N_4149,N_4196);
nand U4400 (N_4400,N_4217,N_4321);
nor U4401 (N_4401,N_4328,N_4246);
xnor U4402 (N_4402,N_4352,N_4273);
or U4403 (N_4403,N_4208,N_4390);
and U4404 (N_4404,N_4232,N_4214);
or U4405 (N_4405,N_4283,N_4366);
nor U4406 (N_4406,N_4327,N_4386);
or U4407 (N_4407,N_4357,N_4395);
or U4408 (N_4408,N_4236,N_4201);
and U4409 (N_4409,N_4221,N_4385);
and U4410 (N_4410,N_4392,N_4346);
nand U4411 (N_4411,N_4314,N_4340);
or U4412 (N_4412,N_4375,N_4234);
or U4413 (N_4413,N_4229,N_4317);
nor U4414 (N_4414,N_4339,N_4311);
nand U4415 (N_4415,N_4396,N_4342);
nor U4416 (N_4416,N_4387,N_4359);
nand U4417 (N_4417,N_4367,N_4245);
nor U4418 (N_4418,N_4279,N_4253);
nor U4419 (N_4419,N_4393,N_4225);
and U4420 (N_4420,N_4384,N_4290);
and U4421 (N_4421,N_4312,N_4356);
xnor U4422 (N_4422,N_4293,N_4333);
nor U4423 (N_4423,N_4382,N_4228);
nor U4424 (N_4424,N_4376,N_4336);
or U4425 (N_4425,N_4291,N_4389);
or U4426 (N_4426,N_4200,N_4275);
nor U4427 (N_4427,N_4238,N_4285);
nor U4428 (N_4428,N_4269,N_4324);
xnor U4429 (N_4429,N_4300,N_4237);
and U4430 (N_4430,N_4358,N_4364);
or U4431 (N_4431,N_4368,N_4256);
or U4432 (N_4432,N_4315,N_4383);
or U4433 (N_4433,N_4202,N_4276);
or U4434 (N_4434,N_4260,N_4298);
and U4435 (N_4435,N_4353,N_4394);
nor U4436 (N_4436,N_4391,N_4306);
nand U4437 (N_4437,N_4272,N_4329);
nor U4438 (N_4438,N_4313,N_4205);
nand U4439 (N_4439,N_4226,N_4363);
nand U4440 (N_4440,N_4277,N_4207);
nand U4441 (N_4441,N_4224,N_4255);
xnor U4442 (N_4442,N_4223,N_4295);
or U4443 (N_4443,N_4380,N_4398);
or U4444 (N_4444,N_4247,N_4233);
nor U4445 (N_4445,N_4284,N_4203);
or U4446 (N_4446,N_4369,N_4362);
or U4447 (N_4447,N_4319,N_4209);
nor U4448 (N_4448,N_4219,N_4282);
or U4449 (N_4449,N_4211,N_4280);
nor U4450 (N_4450,N_4250,N_4302);
and U4451 (N_4451,N_4216,N_4240);
and U4452 (N_4452,N_4331,N_4265);
and U4453 (N_4453,N_4373,N_4325);
or U4454 (N_4454,N_4281,N_4239);
xor U4455 (N_4455,N_4278,N_4289);
nor U4456 (N_4456,N_4299,N_4347);
xor U4457 (N_4457,N_4274,N_4341);
nand U4458 (N_4458,N_4294,N_4220);
nor U4459 (N_4459,N_4215,N_4303);
or U4460 (N_4460,N_4349,N_4268);
nand U4461 (N_4461,N_4377,N_4355);
or U4462 (N_4462,N_4337,N_4263);
nor U4463 (N_4463,N_4379,N_4242);
or U4464 (N_4464,N_4243,N_4251);
nand U4465 (N_4465,N_4388,N_4248);
nand U4466 (N_4466,N_4305,N_4332);
and U4467 (N_4467,N_4212,N_4345);
nand U4468 (N_4468,N_4399,N_4267);
nand U4469 (N_4469,N_4227,N_4288);
or U4470 (N_4470,N_4286,N_4261);
nand U4471 (N_4471,N_4222,N_4213);
nand U4472 (N_4472,N_4316,N_4231);
xor U4473 (N_4473,N_4309,N_4370);
nand U4474 (N_4474,N_4264,N_4343);
nor U4475 (N_4475,N_4230,N_4361);
and U4476 (N_4476,N_4301,N_4257);
or U4477 (N_4477,N_4335,N_4320);
or U4478 (N_4478,N_4287,N_4365);
xnor U4479 (N_4479,N_4262,N_4378);
nor U4480 (N_4480,N_4259,N_4350);
or U4481 (N_4481,N_4360,N_4249);
or U4482 (N_4482,N_4344,N_4297);
nand U4483 (N_4483,N_4308,N_4304);
and U4484 (N_4484,N_4252,N_4323);
nand U4485 (N_4485,N_4235,N_4296);
nor U4486 (N_4486,N_4266,N_4310);
nor U4487 (N_4487,N_4292,N_4351);
and U4488 (N_4488,N_4330,N_4322);
nand U4489 (N_4489,N_4338,N_4354);
or U4490 (N_4490,N_4218,N_4307);
nand U4491 (N_4491,N_4334,N_4371);
nor U4492 (N_4492,N_4206,N_4318);
and U4493 (N_4493,N_4204,N_4254);
xor U4494 (N_4494,N_4244,N_4258);
nand U4495 (N_4495,N_4326,N_4270);
nand U4496 (N_4496,N_4271,N_4397);
and U4497 (N_4497,N_4372,N_4348);
and U4498 (N_4498,N_4241,N_4374);
nand U4499 (N_4499,N_4210,N_4381);
or U4500 (N_4500,N_4255,N_4284);
nor U4501 (N_4501,N_4243,N_4377);
and U4502 (N_4502,N_4259,N_4335);
and U4503 (N_4503,N_4383,N_4379);
or U4504 (N_4504,N_4240,N_4202);
or U4505 (N_4505,N_4253,N_4321);
nor U4506 (N_4506,N_4333,N_4289);
or U4507 (N_4507,N_4299,N_4263);
nor U4508 (N_4508,N_4327,N_4321);
nor U4509 (N_4509,N_4386,N_4273);
nand U4510 (N_4510,N_4343,N_4390);
nor U4511 (N_4511,N_4358,N_4245);
xnor U4512 (N_4512,N_4344,N_4223);
and U4513 (N_4513,N_4285,N_4354);
or U4514 (N_4514,N_4399,N_4323);
and U4515 (N_4515,N_4257,N_4386);
and U4516 (N_4516,N_4236,N_4282);
xnor U4517 (N_4517,N_4249,N_4221);
or U4518 (N_4518,N_4202,N_4304);
nor U4519 (N_4519,N_4208,N_4223);
or U4520 (N_4520,N_4321,N_4385);
and U4521 (N_4521,N_4230,N_4311);
nor U4522 (N_4522,N_4364,N_4229);
nor U4523 (N_4523,N_4296,N_4298);
nor U4524 (N_4524,N_4384,N_4253);
nand U4525 (N_4525,N_4293,N_4265);
and U4526 (N_4526,N_4379,N_4388);
xnor U4527 (N_4527,N_4336,N_4369);
and U4528 (N_4528,N_4386,N_4377);
nor U4529 (N_4529,N_4213,N_4342);
nand U4530 (N_4530,N_4205,N_4367);
or U4531 (N_4531,N_4268,N_4280);
xnor U4532 (N_4532,N_4262,N_4232);
and U4533 (N_4533,N_4309,N_4246);
or U4534 (N_4534,N_4335,N_4358);
nor U4535 (N_4535,N_4345,N_4253);
nor U4536 (N_4536,N_4358,N_4305);
or U4537 (N_4537,N_4321,N_4243);
or U4538 (N_4538,N_4368,N_4212);
and U4539 (N_4539,N_4341,N_4251);
nand U4540 (N_4540,N_4276,N_4298);
and U4541 (N_4541,N_4270,N_4283);
or U4542 (N_4542,N_4349,N_4395);
and U4543 (N_4543,N_4362,N_4233);
nor U4544 (N_4544,N_4259,N_4301);
nand U4545 (N_4545,N_4265,N_4313);
or U4546 (N_4546,N_4307,N_4294);
nor U4547 (N_4547,N_4324,N_4325);
nand U4548 (N_4548,N_4304,N_4367);
or U4549 (N_4549,N_4226,N_4355);
and U4550 (N_4550,N_4351,N_4242);
xnor U4551 (N_4551,N_4317,N_4224);
and U4552 (N_4552,N_4317,N_4222);
xor U4553 (N_4553,N_4294,N_4246);
nand U4554 (N_4554,N_4300,N_4219);
and U4555 (N_4555,N_4288,N_4259);
nand U4556 (N_4556,N_4216,N_4303);
nor U4557 (N_4557,N_4220,N_4325);
and U4558 (N_4558,N_4208,N_4328);
and U4559 (N_4559,N_4367,N_4273);
nand U4560 (N_4560,N_4321,N_4211);
or U4561 (N_4561,N_4268,N_4228);
or U4562 (N_4562,N_4204,N_4234);
nor U4563 (N_4563,N_4375,N_4325);
nor U4564 (N_4564,N_4283,N_4297);
nor U4565 (N_4565,N_4362,N_4382);
and U4566 (N_4566,N_4263,N_4305);
or U4567 (N_4567,N_4339,N_4325);
and U4568 (N_4568,N_4368,N_4233);
nand U4569 (N_4569,N_4252,N_4221);
nor U4570 (N_4570,N_4367,N_4215);
or U4571 (N_4571,N_4393,N_4213);
nand U4572 (N_4572,N_4312,N_4317);
nand U4573 (N_4573,N_4322,N_4368);
or U4574 (N_4574,N_4213,N_4244);
and U4575 (N_4575,N_4346,N_4269);
nor U4576 (N_4576,N_4352,N_4292);
or U4577 (N_4577,N_4226,N_4351);
or U4578 (N_4578,N_4302,N_4364);
and U4579 (N_4579,N_4336,N_4215);
nor U4580 (N_4580,N_4260,N_4245);
xor U4581 (N_4581,N_4254,N_4346);
or U4582 (N_4582,N_4292,N_4263);
nor U4583 (N_4583,N_4354,N_4255);
or U4584 (N_4584,N_4382,N_4283);
or U4585 (N_4585,N_4226,N_4243);
nor U4586 (N_4586,N_4288,N_4258);
and U4587 (N_4587,N_4312,N_4310);
and U4588 (N_4588,N_4302,N_4284);
nor U4589 (N_4589,N_4325,N_4214);
or U4590 (N_4590,N_4345,N_4392);
or U4591 (N_4591,N_4367,N_4353);
nand U4592 (N_4592,N_4392,N_4336);
or U4593 (N_4593,N_4253,N_4348);
or U4594 (N_4594,N_4210,N_4370);
nand U4595 (N_4595,N_4293,N_4382);
or U4596 (N_4596,N_4209,N_4360);
or U4597 (N_4597,N_4301,N_4329);
nor U4598 (N_4598,N_4293,N_4350);
and U4599 (N_4599,N_4276,N_4255);
or U4600 (N_4600,N_4476,N_4534);
and U4601 (N_4601,N_4495,N_4592);
or U4602 (N_4602,N_4448,N_4522);
and U4603 (N_4603,N_4503,N_4593);
nand U4604 (N_4604,N_4435,N_4504);
nand U4605 (N_4605,N_4416,N_4402);
nand U4606 (N_4606,N_4472,N_4405);
and U4607 (N_4607,N_4479,N_4540);
or U4608 (N_4608,N_4509,N_4515);
nand U4609 (N_4609,N_4525,N_4417);
nand U4610 (N_4610,N_4488,N_4581);
and U4611 (N_4611,N_4501,N_4570);
xor U4612 (N_4612,N_4591,N_4452);
nand U4613 (N_4613,N_4572,N_4541);
nand U4614 (N_4614,N_4464,N_4524);
or U4615 (N_4615,N_4561,N_4573);
xor U4616 (N_4616,N_4533,N_4582);
or U4617 (N_4617,N_4461,N_4518);
and U4618 (N_4618,N_4446,N_4571);
xnor U4619 (N_4619,N_4489,N_4498);
nor U4620 (N_4620,N_4458,N_4440);
and U4621 (N_4621,N_4437,N_4460);
or U4622 (N_4622,N_4548,N_4547);
nor U4623 (N_4623,N_4493,N_4517);
nor U4624 (N_4624,N_4442,N_4411);
nand U4625 (N_4625,N_4466,N_4430);
nand U4626 (N_4626,N_4550,N_4595);
nor U4627 (N_4627,N_4559,N_4447);
and U4628 (N_4628,N_4563,N_4567);
nor U4629 (N_4629,N_4566,N_4409);
nand U4630 (N_4630,N_4484,N_4439);
nor U4631 (N_4631,N_4555,N_4404);
and U4632 (N_4632,N_4438,N_4485);
nand U4633 (N_4633,N_4478,N_4568);
and U4634 (N_4634,N_4575,N_4549);
or U4635 (N_4635,N_4450,N_4530);
or U4636 (N_4636,N_4401,N_4556);
nand U4637 (N_4637,N_4445,N_4414);
or U4638 (N_4638,N_4510,N_4507);
nand U4639 (N_4639,N_4418,N_4436);
or U4640 (N_4640,N_4463,N_4511);
and U4641 (N_4641,N_4456,N_4426);
and U4642 (N_4642,N_4521,N_4597);
nand U4643 (N_4643,N_4576,N_4429);
nor U4644 (N_4644,N_4529,N_4494);
xnor U4645 (N_4645,N_4403,N_4532);
or U4646 (N_4646,N_4574,N_4586);
nand U4647 (N_4647,N_4496,N_4543);
nand U4648 (N_4648,N_4523,N_4537);
and U4649 (N_4649,N_4470,N_4433);
or U4650 (N_4650,N_4474,N_4565);
nor U4651 (N_4651,N_4526,N_4406);
nor U4652 (N_4652,N_4560,N_4410);
nor U4653 (N_4653,N_4519,N_4455);
or U4654 (N_4654,N_4554,N_4457);
nor U4655 (N_4655,N_4468,N_4590);
or U4656 (N_4656,N_4531,N_4490);
or U4657 (N_4657,N_4588,N_4505);
nand U4658 (N_4658,N_4465,N_4546);
xnor U4659 (N_4659,N_4441,N_4587);
xnor U4660 (N_4660,N_4562,N_4598);
nor U4661 (N_4661,N_4473,N_4539);
nand U4662 (N_4662,N_4513,N_4512);
nor U4663 (N_4663,N_4449,N_4583);
and U4664 (N_4664,N_4594,N_4545);
and U4665 (N_4665,N_4538,N_4407);
and U4666 (N_4666,N_4506,N_4453);
or U4667 (N_4667,N_4502,N_4497);
xor U4668 (N_4668,N_4462,N_4542);
and U4669 (N_4669,N_4413,N_4412);
nand U4670 (N_4670,N_4599,N_4500);
or U4671 (N_4671,N_4508,N_4432);
nor U4672 (N_4672,N_4400,N_4528);
nor U4673 (N_4673,N_4408,N_4499);
or U4674 (N_4674,N_4577,N_4431);
or U4675 (N_4675,N_4454,N_4558);
nor U4676 (N_4676,N_4424,N_4444);
xnor U4677 (N_4677,N_4483,N_4423);
or U4678 (N_4678,N_4487,N_4584);
nor U4679 (N_4679,N_4578,N_4551);
and U4680 (N_4680,N_4527,N_4564);
nor U4681 (N_4681,N_4419,N_4579);
xnor U4682 (N_4682,N_4481,N_4569);
and U4683 (N_4683,N_4415,N_4585);
nor U4684 (N_4684,N_4459,N_4420);
nor U4685 (N_4685,N_4514,N_4552);
or U4686 (N_4686,N_4427,N_4434);
and U4687 (N_4687,N_4589,N_4544);
nor U4688 (N_4688,N_4491,N_4421);
nor U4689 (N_4689,N_4475,N_4553);
nor U4690 (N_4690,N_4477,N_4443);
or U4691 (N_4691,N_4428,N_4557);
or U4692 (N_4692,N_4516,N_4535);
or U4693 (N_4693,N_4520,N_4480);
nor U4694 (N_4694,N_4492,N_4536);
or U4695 (N_4695,N_4596,N_4422);
or U4696 (N_4696,N_4425,N_4486);
or U4697 (N_4697,N_4469,N_4467);
nand U4698 (N_4698,N_4580,N_4471);
or U4699 (N_4699,N_4451,N_4482);
xnor U4700 (N_4700,N_4589,N_4475);
or U4701 (N_4701,N_4505,N_4511);
and U4702 (N_4702,N_4431,N_4565);
nor U4703 (N_4703,N_4551,N_4425);
nor U4704 (N_4704,N_4507,N_4429);
or U4705 (N_4705,N_4581,N_4477);
or U4706 (N_4706,N_4598,N_4448);
xnor U4707 (N_4707,N_4561,N_4436);
and U4708 (N_4708,N_4540,N_4470);
xor U4709 (N_4709,N_4494,N_4414);
or U4710 (N_4710,N_4485,N_4528);
or U4711 (N_4711,N_4441,N_4422);
and U4712 (N_4712,N_4575,N_4531);
nor U4713 (N_4713,N_4501,N_4404);
nor U4714 (N_4714,N_4565,N_4477);
or U4715 (N_4715,N_4550,N_4405);
or U4716 (N_4716,N_4538,N_4427);
nor U4717 (N_4717,N_4581,N_4473);
xnor U4718 (N_4718,N_4406,N_4534);
or U4719 (N_4719,N_4421,N_4410);
or U4720 (N_4720,N_4567,N_4491);
and U4721 (N_4721,N_4435,N_4450);
nand U4722 (N_4722,N_4407,N_4400);
nor U4723 (N_4723,N_4536,N_4579);
and U4724 (N_4724,N_4405,N_4481);
or U4725 (N_4725,N_4429,N_4444);
or U4726 (N_4726,N_4583,N_4416);
nor U4727 (N_4727,N_4401,N_4479);
or U4728 (N_4728,N_4498,N_4567);
and U4729 (N_4729,N_4437,N_4467);
nor U4730 (N_4730,N_4599,N_4531);
xor U4731 (N_4731,N_4571,N_4419);
or U4732 (N_4732,N_4557,N_4556);
and U4733 (N_4733,N_4486,N_4417);
nor U4734 (N_4734,N_4572,N_4562);
xor U4735 (N_4735,N_4553,N_4523);
and U4736 (N_4736,N_4456,N_4435);
or U4737 (N_4737,N_4474,N_4567);
or U4738 (N_4738,N_4564,N_4510);
nand U4739 (N_4739,N_4545,N_4430);
nand U4740 (N_4740,N_4506,N_4406);
nand U4741 (N_4741,N_4535,N_4566);
and U4742 (N_4742,N_4568,N_4557);
or U4743 (N_4743,N_4423,N_4479);
nand U4744 (N_4744,N_4500,N_4520);
nor U4745 (N_4745,N_4592,N_4498);
or U4746 (N_4746,N_4537,N_4478);
or U4747 (N_4747,N_4562,N_4557);
or U4748 (N_4748,N_4404,N_4400);
nor U4749 (N_4749,N_4407,N_4586);
and U4750 (N_4750,N_4406,N_4470);
nand U4751 (N_4751,N_4575,N_4463);
and U4752 (N_4752,N_4494,N_4550);
and U4753 (N_4753,N_4564,N_4470);
nand U4754 (N_4754,N_4412,N_4594);
or U4755 (N_4755,N_4522,N_4550);
and U4756 (N_4756,N_4568,N_4442);
nand U4757 (N_4757,N_4452,N_4496);
or U4758 (N_4758,N_4531,N_4425);
or U4759 (N_4759,N_4481,N_4559);
xor U4760 (N_4760,N_4571,N_4598);
nor U4761 (N_4761,N_4543,N_4581);
nand U4762 (N_4762,N_4589,N_4505);
nor U4763 (N_4763,N_4587,N_4483);
or U4764 (N_4764,N_4515,N_4406);
nor U4765 (N_4765,N_4471,N_4431);
or U4766 (N_4766,N_4593,N_4553);
or U4767 (N_4767,N_4477,N_4525);
nand U4768 (N_4768,N_4534,N_4571);
xnor U4769 (N_4769,N_4471,N_4536);
nor U4770 (N_4770,N_4536,N_4476);
or U4771 (N_4771,N_4573,N_4599);
and U4772 (N_4772,N_4487,N_4571);
nand U4773 (N_4773,N_4415,N_4543);
or U4774 (N_4774,N_4531,N_4496);
or U4775 (N_4775,N_4516,N_4522);
or U4776 (N_4776,N_4557,N_4456);
nand U4777 (N_4777,N_4481,N_4499);
nor U4778 (N_4778,N_4494,N_4469);
or U4779 (N_4779,N_4464,N_4534);
and U4780 (N_4780,N_4539,N_4429);
nor U4781 (N_4781,N_4552,N_4574);
or U4782 (N_4782,N_4599,N_4461);
or U4783 (N_4783,N_4589,N_4540);
nor U4784 (N_4784,N_4563,N_4404);
or U4785 (N_4785,N_4482,N_4587);
or U4786 (N_4786,N_4567,N_4544);
and U4787 (N_4787,N_4585,N_4522);
nor U4788 (N_4788,N_4417,N_4564);
nor U4789 (N_4789,N_4508,N_4530);
xor U4790 (N_4790,N_4487,N_4588);
or U4791 (N_4791,N_4517,N_4577);
nand U4792 (N_4792,N_4599,N_4518);
nand U4793 (N_4793,N_4469,N_4432);
or U4794 (N_4794,N_4461,N_4551);
or U4795 (N_4795,N_4445,N_4413);
and U4796 (N_4796,N_4522,N_4554);
and U4797 (N_4797,N_4483,N_4504);
and U4798 (N_4798,N_4536,N_4578);
nor U4799 (N_4799,N_4549,N_4470);
xor U4800 (N_4800,N_4799,N_4779);
nand U4801 (N_4801,N_4694,N_4687);
nor U4802 (N_4802,N_4617,N_4757);
and U4803 (N_4803,N_4656,N_4625);
and U4804 (N_4804,N_4674,N_4790);
or U4805 (N_4805,N_4763,N_4608);
xnor U4806 (N_4806,N_4760,N_4715);
or U4807 (N_4807,N_4751,N_4690);
and U4808 (N_4808,N_4652,N_4786);
nand U4809 (N_4809,N_4713,N_4663);
nand U4810 (N_4810,N_4741,N_4791);
nand U4811 (N_4811,N_4645,N_4739);
nor U4812 (N_4812,N_4758,N_4701);
nand U4813 (N_4813,N_4734,N_4667);
nand U4814 (N_4814,N_4776,N_4771);
nor U4815 (N_4815,N_4628,N_4784);
or U4816 (N_4816,N_4736,N_4759);
or U4817 (N_4817,N_4721,N_4788);
nand U4818 (N_4818,N_4697,N_4660);
xnor U4819 (N_4819,N_4650,N_4699);
or U4820 (N_4820,N_4795,N_4621);
or U4821 (N_4821,N_4769,N_4724);
and U4822 (N_4822,N_4601,N_4752);
nor U4823 (N_4823,N_4657,N_4689);
and U4824 (N_4824,N_4731,N_4728);
or U4825 (N_4825,N_4710,N_4643);
and U4826 (N_4826,N_4793,N_4647);
xor U4827 (N_4827,N_4743,N_4716);
or U4828 (N_4828,N_4609,N_4677);
and U4829 (N_4829,N_4756,N_4633);
nand U4830 (N_4830,N_4631,N_4666);
or U4831 (N_4831,N_4700,N_4746);
nand U4832 (N_4832,N_4636,N_4673);
nand U4833 (N_4833,N_4698,N_4789);
nor U4834 (N_4834,N_4692,N_4745);
and U4835 (N_4835,N_4653,N_4671);
nor U4836 (N_4836,N_4618,N_4750);
and U4837 (N_4837,N_4717,N_4733);
nor U4838 (N_4838,N_4764,N_4642);
and U4839 (N_4839,N_4602,N_4670);
or U4840 (N_4840,N_4735,N_4794);
nand U4841 (N_4841,N_4708,N_4648);
and U4842 (N_4842,N_4744,N_4696);
nand U4843 (N_4843,N_4632,N_4600);
or U4844 (N_4844,N_4729,N_4668);
and U4845 (N_4845,N_4768,N_4691);
nor U4846 (N_4846,N_4611,N_4765);
and U4847 (N_4847,N_4635,N_4603);
or U4848 (N_4848,N_4669,N_4703);
and U4849 (N_4849,N_4641,N_4624);
or U4850 (N_4850,N_4615,N_4772);
or U4851 (N_4851,N_4678,N_4704);
nand U4852 (N_4852,N_4705,N_4792);
nand U4853 (N_4853,N_4798,N_4740);
xor U4854 (N_4854,N_4640,N_4655);
or U4855 (N_4855,N_4676,N_4762);
and U4856 (N_4856,N_4754,N_4679);
nor U4857 (N_4857,N_4723,N_4738);
xor U4858 (N_4858,N_4742,N_4714);
nor U4859 (N_4859,N_4658,N_4637);
nor U4860 (N_4860,N_4707,N_4665);
nand U4861 (N_4861,N_4630,N_4626);
nand U4862 (N_4862,N_4619,N_4718);
nand U4863 (N_4863,N_4712,N_4755);
or U4864 (N_4864,N_4646,N_4639);
and U4865 (N_4865,N_4681,N_4605);
nand U4866 (N_4866,N_4651,N_4782);
or U4867 (N_4867,N_4766,N_4607);
and U4868 (N_4868,N_4649,N_4616);
and U4869 (N_4869,N_4664,N_4706);
nand U4870 (N_4870,N_4622,N_4623);
and U4871 (N_4871,N_4761,N_4688);
nand U4872 (N_4872,N_4702,N_4680);
or U4873 (N_4873,N_4749,N_4737);
nor U4874 (N_4874,N_4777,N_4634);
or U4875 (N_4875,N_4725,N_4610);
xnor U4876 (N_4876,N_4797,N_4682);
nor U4877 (N_4877,N_4604,N_4662);
or U4878 (N_4878,N_4727,N_4770);
nand U4879 (N_4879,N_4659,N_4780);
nor U4880 (N_4880,N_4719,N_4614);
xnor U4881 (N_4881,N_4747,N_4695);
nand U4882 (N_4882,N_4774,N_4722);
or U4883 (N_4883,N_4709,N_4775);
or U4884 (N_4884,N_4675,N_4796);
or U4885 (N_4885,N_4606,N_4620);
and U4886 (N_4886,N_4785,N_4684);
nor U4887 (N_4887,N_4685,N_4753);
nor U4888 (N_4888,N_4720,N_4612);
nand U4889 (N_4889,N_4748,N_4773);
nand U4890 (N_4890,N_4732,N_4693);
or U4891 (N_4891,N_4661,N_4683);
nand U4892 (N_4892,N_4654,N_4787);
xnor U4893 (N_4893,N_4627,N_4686);
nand U4894 (N_4894,N_4638,N_4767);
nor U4895 (N_4895,N_4730,N_4783);
xnor U4896 (N_4896,N_4629,N_4726);
or U4897 (N_4897,N_4711,N_4781);
nor U4898 (N_4898,N_4672,N_4613);
or U4899 (N_4899,N_4644,N_4778);
nor U4900 (N_4900,N_4784,N_4780);
and U4901 (N_4901,N_4756,N_4751);
nor U4902 (N_4902,N_4658,N_4648);
or U4903 (N_4903,N_4762,N_4653);
nand U4904 (N_4904,N_4724,N_4673);
nand U4905 (N_4905,N_4710,N_4669);
nand U4906 (N_4906,N_4608,N_4722);
nor U4907 (N_4907,N_4738,N_4781);
or U4908 (N_4908,N_4627,N_4630);
and U4909 (N_4909,N_4736,N_4698);
nand U4910 (N_4910,N_4639,N_4694);
and U4911 (N_4911,N_4765,N_4787);
or U4912 (N_4912,N_4667,N_4639);
nor U4913 (N_4913,N_4603,N_4608);
nand U4914 (N_4914,N_4778,N_4711);
nand U4915 (N_4915,N_4703,N_4673);
or U4916 (N_4916,N_4748,N_4747);
nor U4917 (N_4917,N_4622,N_4692);
nor U4918 (N_4918,N_4676,N_4711);
nor U4919 (N_4919,N_4793,N_4682);
or U4920 (N_4920,N_4668,N_4796);
or U4921 (N_4921,N_4687,N_4799);
nor U4922 (N_4922,N_4790,N_4725);
nor U4923 (N_4923,N_4737,N_4668);
nor U4924 (N_4924,N_4787,N_4741);
and U4925 (N_4925,N_4661,N_4686);
nand U4926 (N_4926,N_4639,N_4720);
nor U4927 (N_4927,N_4641,N_4614);
or U4928 (N_4928,N_4635,N_4689);
xor U4929 (N_4929,N_4716,N_4640);
nor U4930 (N_4930,N_4627,N_4654);
and U4931 (N_4931,N_4684,N_4607);
nand U4932 (N_4932,N_4749,N_4761);
or U4933 (N_4933,N_4681,N_4785);
nand U4934 (N_4934,N_4652,N_4739);
xnor U4935 (N_4935,N_4643,N_4655);
nor U4936 (N_4936,N_4629,N_4770);
nor U4937 (N_4937,N_4721,N_4698);
and U4938 (N_4938,N_4664,N_4700);
nor U4939 (N_4939,N_4648,N_4713);
nand U4940 (N_4940,N_4644,N_4714);
nor U4941 (N_4941,N_4641,N_4667);
or U4942 (N_4942,N_4733,N_4687);
and U4943 (N_4943,N_4709,N_4761);
nand U4944 (N_4944,N_4611,N_4738);
nand U4945 (N_4945,N_4785,N_4702);
and U4946 (N_4946,N_4790,N_4630);
or U4947 (N_4947,N_4711,N_4643);
or U4948 (N_4948,N_4621,N_4712);
nor U4949 (N_4949,N_4672,N_4773);
or U4950 (N_4950,N_4686,N_4746);
and U4951 (N_4951,N_4610,N_4739);
or U4952 (N_4952,N_4605,N_4738);
nor U4953 (N_4953,N_4788,N_4772);
nand U4954 (N_4954,N_4653,N_4676);
or U4955 (N_4955,N_4657,N_4760);
or U4956 (N_4956,N_4647,N_4663);
nor U4957 (N_4957,N_4738,N_4774);
and U4958 (N_4958,N_4614,N_4715);
and U4959 (N_4959,N_4722,N_4651);
xor U4960 (N_4960,N_4717,N_4639);
nor U4961 (N_4961,N_4692,N_4738);
and U4962 (N_4962,N_4629,N_4710);
nor U4963 (N_4963,N_4639,N_4715);
nor U4964 (N_4964,N_4680,N_4748);
or U4965 (N_4965,N_4697,N_4774);
or U4966 (N_4966,N_4724,N_4672);
or U4967 (N_4967,N_4621,N_4766);
nand U4968 (N_4968,N_4775,N_4661);
and U4969 (N_4969,N_4730,N_4753);
nor U4970 (N_4970,N_4640,N_4686);
or U4971 (N_4971,N_4797,N_4795);
nor U4972 (N_4972,N_4774,N_4714);
nor U4973 (N_4973,N_4785,N_4652);
xor U4974 (N_4974,N_4719,N_4705);
nor U4975 (N_4975,N_4608,N_4757);
and U4976 (N_4976,N_4680,N_4699);
nand U4977 (N_4977,N_4614,N_4610);
nand U4978 (N_4978,N_4743,N_4679);
and U4979 (N_4979,N_4714,N_4778);
and U4980 (N_4980,N_4705,N_4768);
or U4981 (N_4981,N_4613,N_4706);
or U4982 (N_4982,N_4628,N_4794);
xnor U4983 (N_4983,N_4757,N_4611);
and U4984 (N_4984,N_4653,N_4770);
and U4985 (N_4985,N_4737,N_4660);
or U4986 (N_4986,N_4657,N_4621);
or U4987 (N_4987,N_4675,N_4606);
nand U4988 (N_4988,N_4637,N_4702);
nand U4989 (N_4989,N_4671,N_4636);
or U4990 (N_4990,N_4781,N_4735);
nor U4991 (N_4991,N_4759,N_4607);
nor U4992 (N_4992,N_4721,N_4691);
nand U4993 (N_4993,N_4759,N_4620);
and U4994 (N_4994,N_4796,N_4617);
and U4995 (N_4995,N_4626,N_4751);
and U4996 (N_4996,N_4735,N_4658);
xor U4997 (N_4997,N_4743,N_4726);
nand U4998 (N_4998,N_4731,N_4674);
and U4999 (N_4999,N_4728,N_4709);
or UO_0 (O_0,N_4913,N_4935);
nor UO_1 (O_1,N_4886,N_4863);
nor UO_2 (O_2,N_4979,N_4872);
or UO_3 (O_3,N_4989,N_4849);
or UO_4 (O_4,N_4919,N_4911);
xnor UO_5 (O_5,N_4998,N_4864);
xnor UO_6 (O_6,N_4865,N_4952);
nand UO_7 (O_7,N_4828,N_4895);
nor UO_8 (O_8,N_4986,N_4845);
or UO_9 (O_9,N_4967,N_4927);
or UO_10 (O_10,N_4889,N_4946);
and UO_11 (O_11,N_4902,N_4819);
nand UO_12 (O_12,N_4993,N_4947);
nor UO_13 (O_13,N_4892,N_4983);
nor UO_14 (O_14,N_4879,N_4851);
nor UO_15 (O_15,N_4970,N_4873);
nand UO_16 (O_16,N_4957,N_4977);
nand UO_17 (O_17,N_4976,N_4885);
nor UO_18 (O_18,N_4800,N_4971);
nand UO_19 (O_19,N_4887,N_4921);
and UO_20 (O_20,N_4988,N_4939);
or UO_21 (O_21,N_4918,N_4923);
nor UO_22 (O_22,N_4958,N_4909);
nor UO_23 (O_23,N_4848,N_4944);
and UO_24 (O_24,N_4920,N_4853);
xnor UO_25 (O_25,N_4890,N_4930);
or UO_26 (O_26,N_4928,N_4868);
and UO_27 (O_27,N_4994,N_4860);
nand UO_28 (O_28,N_4821,N_4884);
xor UO_29 (O_29,N_4999,N_4817);
nor UO_30 (O_30,N_4899,N_4869);
nor UO_31 (O_31,N_4840,N_4894);
xnor UO_32 (O_32,N_4896,N_4907);
nor UO_33 (O_33,N_4812,N_4905);
or UO_34 (O_34,N_4802,N_4975);
or UO_35 (O_35,N_4901,N_4950);
and UO_36 (O_36,N_4898,N_4910);
nand UO_37 (O_37,N_4831,N_4995);
nand UO_38 (O_38,N_4893,N_4839);
or UO_39 (O_39,N_4940,N_4938);
nor UO_40 (O_40,N_4991,N_4854);
and UO_41 (O_41,N_4941,N_4897);
nand UO_42 (O_42,N_4888,N_4980);
nor UO_43 (O_43,N_4933,N_4917);
and UO_44 (O_44,N_4875,N_4856);
or UO_45 (O_45,N_4847,N_4818);
xnor UO_46 (O_46,N_4814,N_4972);
and UO_47 (O_47,N_4992,N_4838);
nand UO_48 (O_48,N_4906,N_4969);
nor UO_49 (O_49,N_4841,N_4877);
or UO_50 (O_50,N_4951,N_4966);
nor UO_51 (O_51,N_4805,N_4945);
nand UO_52 (O_52,N_4830,N_4883);
and UO_53 (O_53,N_4843,N_4916);
and UO_54 (O_54,N_4891,N_4823);
or UO_55 (O_55,N_4937,N_4931);
or UO_56 (O_56,N_4810,N_4974);
nand UO_57 (O_57,N_4866,N_4852);
and UO_58 (O_58,N_4942,N_4981);
or UO_59 (O_59,N_4878,N_4908);
nor UO_60 (O_60,N_4973,N_4968);
and UO_61 (O_61,N_4929,N_4964);
or UO_62 (O_62,N_4903,N_4963);
nor UO_63 (O_63,N_4826,N_4804);
or UO_64 (O_64,N_4806,N_4962);
and UO_65 (O_65,N_4859,N_4850);
xor UO_66 (O_66,N_4961,N_4932);
or UO_67 (O_67,N_4936,N_4808);
or UO_68 (O_68,N_4811,N_4862);
nand UO_69 (O_69,N_4881,N_4978);
or UO_70 (O_70,N_4867,N_4824);
nor UO_71 (O_71,N_4985,N_4987);
and UO_72 (O_72,N_4801,N_4855);
and UO_73 (O_73,N_4904,N_4813);
or UO_74 (O_74,N_4825,N_4833);
or UO_75 (O_75,N_4857,N_4871);
or UO_76 (O_76,N_4829,N_4959);
nor UO_77 (O_77,N_4956,N_4925);
or UO_78 (O_78,N_4915,N_4832);
or UO_79 (O_79,N_4948,N_4820);
nor UO_80 (O_80,N_4990,N_4816);
or UO_81 (O_81,N_4827,N_4984);
nor UO_82 (O_82,N_4809,N_4996);
nor UO_83 (O_83,N_4842,N_4982);
or UO_84 (O_84,N_4844,N_4953);
and UO_85 (O_85,N_4954,N_4924);
nor UO_86 (O_86,N_4943,N_4880);
nor UO_87 (O_87,N_4858,N_4882);
or UO_88 (O_88,N_4965,N_4815);
nor UO_89 (O_89,N_4900,N_4870);
or UO_90 (O_90,N_4807,N_4874);
and UO_91 (O_91,N_4846,N_4837);
nand UO_92 (O_92,N_4997,N_4949);
nand UO_93 (O_93,N_4960,N_4912);
nand UO_94 (O_94,N_4876,N_4922);
or UO_95 (O_95,N_4803,N_4934);
nand UO_96 (O_96,N_4914,N_4861);
nor UO_97 (O_97,N_4926,N_4834);
nor UO_98 (O_98,N_4822,N_4955);
or UO_99 (O_99,N_4836,N_4835);
nor UO_100 (O_100,N_4840,N_4909);
or UO_101 (O_101,N_4914,N_4813);
nor UO_102 (O_102,N_4850,N_4952);
nand UO_103 (O_103,N_4887,N_4995);
nand UO_104 (O_104,N_4901,N_4888);
xor UO_105 (O_105,N_4904,N_4929);
and UO_106 (O_106,N_4866,N_4905);
or UO_107 (O_107,N_4934,N_4917);
xor UO_108 (O_108,N_4971,N_4936);
nor UO_109 (O_109,N_4817,N_4975);
and UO_110 (O_110,N_4936,N_4807);
nor UO_111 (O_111,N_4921,N_4947);
nand UO_112 (O_112,N_4814,N_4930);
or UO_113 (O_113,N_4818,N_4966);
nor UO_114 (O_114,N_4846,N_4973);
nand UO_115 (O_115,N_4930,N_4893);
nand UO_116 (O_116,N_4832,N_4897);
xnor UO_117 (O_117,N_4902,N_4938);
nand UO_118 (O_118,N_4907,N_4841);
nand UO_119 (O_119,N_4950,N_4825);
and UO_120 (O_120,N_4905,N_4918);
nor UO_121 (O_121,N_4828,N_4847);
nor UO_122 (O_122,N_4818,N_4898);
and UO_123 (O_123,N_4830,N_4999);
and UO_124 (O_124,N_4937,N_4858);
and UO_125 (O_125,N_4945,N_4909);
nand UO_126 (O_126,N_4942,N_4952);
nand UO_127 (O_127,N_4944,N_4971);
nor UO_128 (O_128,N_4807,N_4978);
nor UO_129 (O_129,N_4992,N_4859);
or UO_130 (O_130,N_4892,N_4870);
nor UO_131 (O_131,N_4950,N_4837);
nor UO_132 (O_132,N_4998,N_4820);
nand UO_133 (O_133,N_4916,N_4829);
nand UO_134 (O_134,N_4999,N_4875);
nand UO_135 (O_135,N_4902,N_4854);
nand UO_136 (O_136,N_4923,N_4938);
and UO_137 (O_137,N_4863,N_4998);
and UO_138 (O_138,N_4814,N_4984);
nand UO_139 (O_139,N_4964,N_4866);
or UO_140 (O_140,N_4903,N_4875);
nand UO_141 (O_141,N_4944,N_4812);
and UO_142 (O_142,N_4873,N_4801);
or UO_143 (O_143,N_4927,N_4833);
or UO_144 (O_144,N_4892,N_4994);
or UO_145 (O_145,N_4988,N_4904);
nand UO_146 (O_146,N_4973,N_4850);
xnor UO_147 (O_147,N_4904,N_4865);
or UO_148 (O_148,N_4844,N_4870);
and UO_149 (O_149,N_4891,N_4848);
nor UO_150 (O_150,N_4819,N_4805);
and UO_151 (O_151,N_4912,N_4819);
nor UO_152 (O_152,N_4841,N_4933);
nand UO_153 (O_153,N_4976,N_4994);
xor UO_154 (O_154,N_4870,N_4964);
nor UO_155 (O_155,N_4994,N_4959);
or UO_156 (O_156,N_4878,N_4826);
nand UO_157 (O_157,N_4834,N_4826);
and UO_158 (O_158,N_4964,N_4991);
or UO_159 (O_159,N_4802,N_4938);
nand UO_160 (O_160,N_4906,N_4884);
and UO_161 (O_161,N_4803,N_4953);
xnor UO_162 (O_162,N_4923,N_4819);
and UO_163 (O_163,N_4802,N_4922);
or UO_164 (O_164,N_4871,N_4888);
or UO_165 (O_165,N_4991,N_4969);
or UO_166 (O_166,N_4976,N_4986);
nand UO_167 (O_167,N_4843,N_4992);
or UO_168 (O_168,N_4815,N_4901);
or UO_169 (O_169,N_4984,N_4854);
nor UO_170 (O_170,N_4966,N_4968);
nor UO_171 (O_171,N_4906,N_4929);
or UO_172 (O_172,N_4986,N_4847);
nor UO_173 (O_173,N_4915,N_4943);
and UO_174 (O_174,N_4903,N_4939);
or UO_175 (O_175,N_4994,N_4856);
nand UO_176 (O_176,N_4927,N_4875);
or UO_177 (O_177,N_4918,N_4874);
xor UO_178 (O_178,N_4959,N_4808);
nand UO_179 (O_179,N_4969,N_4900);
or UO_180 (O_180,N_4820,N_4911);
nor UO_181 (O_181,N_4854,N_4976);
and UO_182 (O_182,N_4899,N_4855);
or UO_183 (O_183,N_4991,N_4859);
nand UO_184 (O_184,N_4969,N_4863);
xor UO_185 (O_185,N_4875,N_4842);
nand UO_186 (O_186,N_4800,N_4880);
nor UO_187 (O_187,N_4909,N_4952);
or UO_188 (O_188,N_4886,N_4936);
xnor UO_189 (O_189,N_4829,N_4821);
and UO_190 (O_190,N_4809,N_4933);
and UO_191 (O_191,N_4897,N_4983);
xnor UO_192 (O_192,N_4880,N_4841);
xnor UO_193 (O_193,N_4953,N_4829);
nand UO_194 (O_194,N_4873,N_4855);
and UO_195 (O_195,N_4919,N_4877);
xor UO_196 (O_196,N_4901,N_4915);
nand UO_197 (O_197,N_4801,N_4924);
xor UO_198 (O_198,N_4987,N_4807);
or UO_199 (O_199,N_4832,N_4845);
or UO_200 (O_200,N_4959,N_4997);
nand UO_201 (O_201,N_4868,N_4966);
nand UO_202 (O_202,N_4986,N_4945);
nand UO_203 (O_203,N_4902,N_4952);
xor UO_204 (O_204,N_4984,N_4818);
nor UO_205 (O_205,N_4821,N_4824);
or UO_206 (O_206,N_4967,N_4805);
nand UO_207 (O_207,N_4967,N_4866);
nor UO_208 (O_208,N_4862,N_4933);
nand UO_209 (O_209,N_4953,N_4938);
xnor UO_210 (O_210,N_4948,N_4807);
and UO_211 (O_211,N_4864,N_4895);
or UO_212 (O_212,N_4865,N_4893);
xnor UO_213 (O_213,N_4921,N_4932);
nand UO_214 (O_214,N_4877,N_4867);
or UO_215 (O_215,N_4834,N_4913);
nor UO_216 (O_216,N_4908,N_4996);
nor UO_217 (O_217,N_4817,N_4857);
xnor UO_218 (O_218,N_4959,N_4951);
nor UO_219 (O_219,N_4888,N_4917);
nand UO_220 (O_220,N_4925,N_4842);
nor UO_221 (O_221,N_4871,N_4879);
and UO_222 (O_222,N_4948,N_4995);
and UO_223 (O_223,N_4860,N_4911);
and UO_224 (O_224,N_4825,N_4927);
nand UO_225 (O_225,N_4970,N_4929);
nand UO_226 (O_226,N_4956,N_4997);
nor UO_227 (O_227,N_4904,N_4915);
nand UO_228 (O_228,N_4863,N_4872);
and UO_229 (O_229,N_4934,N_4921);
nand UO_230 (O_230,N_4855,N_4916);
xnor UO_231 (O_231,N_4868,N_4927);
or UO_232 (O_232,N_4969,N_4847);
and UO_233 (O_233,N_4959,N_4998);
nor UO_234 (O_234,N_4836,N_4846);
xor UO_235 (O_235,N_4923,N_4989);
and UO_236 (O_236,N_4932,N_4900);
and UO_237 (O_237,N_4870,N_4875);
nand UO_238 (O_238,N_4882,N_4914);
nand UO_239 (O_239,N_4996,N_4820);
nor UO_240 (O_240,N_4988,N_4854);
or UO_241 (O_241,N_4865,N_4858);
nand UO_242 (O_242,N_4808,N_4857);
nor UO_243 (O_243,N_4914,N_4863);
nand UO_244 (O_244,N_4807,N_4811);
and UO_245 (O_245,N_4800,N_4873);
nand UO_246 (O_246,N_4837,N_4854);
and UO_247 (O_247,N_4904,N_4960);
xnor UO_248 (O_248,N_4998,N_4939);
xor UO_249 (O_249,N_4866,N_4865);
nor UO_250 (O_250,N_4984,N_4934);
or UO_251 (O_251,N_4843,N_4949);
and UO_252 (O_252,N_4980,N_4806);
and UO_253 (O_253,N_4877,N_4846);
nor UO_254 (O_254,N_4852,N_4991);
and UO_255 (O_255,N_4977,N_4883);
or UO_256 (O_256,N_4818,N_4889);
nand UO_257 (O_257,N_4981,N_4960);
nor UO_258 (O_258,N_4803,N_4867);
nor UO_259 (O_259,N_4876,N_4893);
and UO_260 (O_260,N_4910,N_4934);
or UO_261 (O_261,N_4876,N_4918);
nor UO_262 (O_262,N_4918,N_4896);
nand UO_263 (O_263,N_4859,N_4875);
nand UO_264 (O_264,N_4818,N_4978);
nor UO_265 (O_265,N_4876,N_4925);
xor UO_266 (O_266,N_4811,N_4983);
or UO_267 (O_267,N_4950,N_4934);
nor UO_268 (O_268,N_4887,N_4959);
nand UO_269 (O_269,N_4950,N_4804);
and UO_270 (O_270,N_4993,N_4982);
or UO_271 (O_271,N_4921,N_4870);
or UO_272 (O_272,N_4802,N_4879);
nor UO_273 (O_273,N_4918,N_4867);
nand UO_274 (O_274,N_4863,N_4878);
nor UO_275 (O_275,N_4908,N_4881);
nor UO_276 (O_276,N_4870,N_4904);
or UO_277 (O_277,N_4928,N_4991);
or UO_278 (O_278,N_4890,N_4936);
or UO_279 (O_279,N_4915,N_4969);
nor UO_280 (O_280,N_4887,N_4996);
nand UO_281 (O_281,N_4855,N_4970);
nand UO_282 (O_282,N_4844,N_4950);
or UO_283 (O_283,N_4946,N_4896);
or UO_284 (O_284,N_4805,N_4904);
nand UO_285 (O_285,N_4874,N_4887);
nor UO_286 (O_286,N_4933,N_4919);
or UO_287 (O_287,N_4880,N_4986);
xor UO_288 (O_288,N_4819,N_4807);
nand UO_289 (O_289,N_4987,N_4989);
or UO_290 (O_290,N_4885,N_4895);
nand UO_291 (O_291,N_4894,N_4943);
nor UO_292 (O_292,N_4988,N_4862);
xnor UO_293 (O_293,N_4952,N_4853);
and UO_294 (O_294,N_4923,N_4887);
or UO_295 (O_295,N_4955,N_4865);
or UO_296 (O_296,N_4838,N_4976);
or UO_297 (O_297,N_4991,N_4930);
or UO_298 (O_298,N_4897,N_4830);
xnor UO_299 (O_299,N_4838,N_4860);
or UO_300 (O_300,N_4800,N_4818);
and UO_301 (O_301,N_4963,N_4921);
nand UO_302 (O_302,N_4893,N_4920);
nor UO_303 (O_303,N_4957,N_4921);
or UO_304 (O_304,N_4938,N_4996);
xor UO_305 (O_305,N_4997,N_4849);
and UO_306 (O_306,N_4955,N_4812);
nor UO_307 (O_307,N_4985,N_4837);
nor UO_308 (O_308,N_4943,N_4874);
and UO_309 (O_309,N_4892,N_4885);
nand UO_310 (O_310,N_4874,N_4825);
and UO_311 (O_311,N_4962,N_4988);
nor UO_312 (O_312,N_4844,N_4943);
nand UO_313 (O_313,N_4919,N_4848);
nor UO_314 (O_314,N_4991,N_4836);
and UO_315 (O_315,N_4950,N_4945);
nand UO_316 (O_316,N_4827,N_4956);
and UO_317 (O_317,N_4961,N_4977);
nor UO_318 (O_318,N_4975,N_4946);
nor UO_319 (O_319,N_4990,N_4876);
or UO_320 (O_320,N_4880,N_4983);
and UO_321 (O_321,N_4990,N_4852);
nand UO_322 (O_322,N_4977,N_4981);
nor UO_323 (O_323,N_4913,N_4838);
nand UO_324 (O_324,N_4878,N_4996);
nor UO_325 (O_325,N_4896,N_4804);
nand UO_326 (O_326,N_4952,N_4921);
xor UO_327 (O_327,N_4945,N_4976);
nor UO_328 (O_328,N_4806,N_4941);
nor UO_329 (O_329,N_4913,N_4914);
xor UO_330 (O_330,N_4908,N_4925);
and UO_331 (O_331,N_4875,N_4801);
nor UO_332 (O_332,N_4973,N_4897);
nand UO_333 (O_333,N_4880,N_4894);
nor UO_334 (O_334,N_4838,N_4890);
nor UO_335 (O_335,N_4987,N_4961);
or UO_336 (O_336,N_4886,N_4822);
nand UO_337 (O_337,N_4825,N_4997);
and UO_338 (O_338,N_4948,N_4899);
or UO_339 (O_339,N_4908,N_4970);
nor UO_340 (O_340,N_4829,N_4994);
and UO_341 (O_341,N_4825,N_4905);
nand UO_342 (O_342,N_4860,N_4877);
xnor UO_343 (O_343,N_4947,N_4909);
nor UO_344 (O_344,N_4896,N_4943);
or UO_345 (O_345,N_4862,N_4923);
nand UO_346 (O_346,N_4962,N_4842);
xor UO_347 (O_347,N_4922,N_4862);
nand UO_348 (O_348,N_4959,N_4832);
and UO_349 (O_349,N_4895,N_4916);
nor UO_350 (O_350,N_4819,N_4845);
and UO_351 (O_351,N_4877,N_4945);
nor UO_352 (O_352,N_4882,N_4869);
xnor UO_353 (O_353,N_4931,N_4895);
or UO_354 (O_354,N_4921,N_4966);
nor UO_355 (O_355,N_4899,N_4900);
or UO_356 (O_356,N_4869,N_4852);
or UO_357 (O_357,N_4884,N_4994);
nand UO_358 (O_358,N_4916,N_4899);
nor UO_359 (O_359,N_4920,N_4808);
nand UO_360 (O_360,N_4925,N_4867);
xor UO_361 (O_361,N_4845,N_4992);
nand UO_362 (O_362,N_4881,N_4819);
or UO_363 (O_363,N_4969,N_4862);
or UO_364 (O_364,N_4962,N_4953);
nand UO_365 (O_365,N_4843,N_4999);
or UO_366 (O_366,N_4818,N_4813);
nand UO_367 (O_367,N_4967,N_4852);
nor UO_368 (O_368,N_4935,N_4926);
nand UO_369 (O_369,N_4891,N_4909);
or UO_370 (O_370,N_4858,N_4956);
nand UO_371 (O_371,N_4810,N_4817);
and UO_372 (O_372,N_4820,N_4870);
and UO_373 (O_373,N_4909,N_4978);
or UO_374 (O_374,N_4986,N_4835);
nor UO_375 (O_375,N_4868,N_4904);
nor UO_376 (O_376,N_4851,N_4994);
xnor UO_377 (O_377,N_4932,N_4939);
and UO_378 (O_378,N_4984,N_4849);
nor UO_379 (O_379,N_4831,N_4956);
xor UO_380 (O_380,N_4830,N_4839);
or UO_381 (O_381,N_4848,N_4948);
nand UO_382 (O_382,N_4939,N_4827);
and UO_383 (O_383,N_4900,N_4882);
nor UO_384 (O_384,N_4957,N_4805);
nand UO_385 (O_385,N_4811,N_4975);
and UO_386 (O_386,N_4951,N_4842);
xor UO_387 (O_387,N_4859,N_4808);
xor UO_388 (O_388,N_4911,N_4967);
xor UO_389 (O_389,N_4982,N_4990);
nand UO_390 (O_390,N_4998,N_4942);
nor UO_391 (O_391,N_4808,N_4901);
nor UO_392 (O_392,N_4944,N_4988);
nand UO_393 (O_393,N_4933,N_4907);
xnor UO_394 (O_394,N_4946,N_4877);
and UO_395 (O_395,N_4842,N_4950);
nand UO_396 (O_396,N_4969,N_4825);
nand UO_397 (O_397,N_4841,N_4864);
and UO_398 (O_398,N_4922,N_4980);
nor UO_399 (O_399,N_4943,N_4831);
nor UO_400 (O_400,N_4859,N_4829);
nor UO_401 (O_401,N_4911,N_4822);
and UO_402 (O_402,N_4933,N_4921);
or UO_403 (O_403,N_4807,N_4989);
nand UO_404 (O_404,N_4890,N_4811);
and UO_405 (O_405,N_4802,N_4830);
or UO_406 (O_406,N_4840,N_4974);
and UO_407 (O_407,N_4909,N_4832);
xor UO_408 (O_408,N_4815,N_4961);
or UO_409 (O_409,N_4934,N_4953);
or UO_410 (O_410,N_4806,N_4971);
or UO_411 (O_411,N_4824,N_4862);
nor UO_412 (O_412,N_4822,N_4827);
or UO_413 (O_413,N_4838,N_4967);
or UO_414 (O_414,N_4976,N_4920);
nor UO_415 (O_415,N_4833,N_4985);
and UO_416 (O_416,N_4890,N_4974);
nand UO_417 (O_417,N_4901,N_4863);
and UO_418 (O_418,N_4875,N_4914);
xor UO_419 (O_419,N_4889,N_4801);
nand UO_420 (O_420,N_4889,N_4913);
nand UO_421 (O_421,N_4955,N_4845);
and UO_422 (O_422,N_4988,N_4826);
or UO_423 (O_423,N_4816,N_4897);
nor UO_424 (O_424,N_4905,N_4888);
or UO_425 (O_425,N_4866,N_4862);
or UO_426 (O_426,N_4911,N_4965);
or UO_427 (O_427,N_4876,N_4910);
nand UO_428 (O_428,N_4869,N_4945);
nand UO_429 (O_429,N_4804,N_4966);
or UO_430 (O_430,N_4978,N_4809);
nand UO_431 (O_431,N_4916,N_4950);
nand UO_432 (O_432,N_4939,N_4867);
or UO_433 (O_433,N_4850,N_4947);
and UO_434 (O_434,N_4893,N_4945);
xor UO_435 (O_435,N_4877,N_4986);
and UO_436 (O_436,N_4960,N_4918);
nand UO_437 (O_437,N_4883,N_4840);
and UO_438 (O_438,N_4840,N_4849);
or UO_439 (O_439,N_4810,N_4826);
or UO_440 (O_440,N_4985,N_4848);
and UO_441 (O_441,N_4970,N_4818);
or UO_442 (O_442,N_4868,N_4806);
or UO_443 (O_443,N_4917,N_4837);
nand UO_444 (O_444,N_4960,N_4965);
nor UO_445 (O_445,N_4976,N_4895);
or UO_446 (O_446,N_4819,N_4944);
nor UO_447 (O_447,N_4847,N_4841);
or UO_448 (O_448,N_4896,N_4924);
and UO_449 (O_449,N_4996,N_4930);
nor UO_450 (O_450,N_4962,N_4883);
and UO_451 (O_451,N_4887,N_4820);
nand UO_452 (O_452,N_4833,N_4883);
or UO_453 (O_453,N_4932,N_4839);
nor UO_454 (O_454,N_4859,N_4812);
and UO_455 (O_455,N_4942,N_4974);
or UO_456 (O_456,N_4827,N_4962);
and UO_457 (O_457,N_4996,N_4935);
nand UO_458 (O_458,N_4827,N_4944);
and UO_459 (O_459,N_4982,N_4974);
or UO_460 (O_460,N_4999,N_4951);
or UO_461 (O_461,N_4840,N_4913);
and UO_462 (O_462,N_4814,N_4928);
and UO_463 (O_463,N_4910,N_4951);
xor UO_464 (O_464,N_4968,N_4924);
nor UO_465 (O_465,N_4974,N_4937);
and UO_466 (O_466,N_4863,N_4850);
and UO_467 (O_467,N_4857,N_4936);
xnor UO_468 (O_468,N_4995,N_4801);
xor UO_469 (O_469,N_4945,N_4919);
nor UO_470 (O_470,N_4896,N_4976);
nor UO_471 (O_471,N_4860,N_4805);
nor UO_472 (O_472,N_4932,N_4898);
or UO_473 (O_473,N_4966,N_4825);
nor UO_474 (O_474,N_4963,N_4836);
nand UO_475 (O_475,N_4834,N_4901);
and UO_476 (O_476,N_4809,N_4983);
and UO_477 (O_477,N_4852,N_4847);
or UO_478 (O_478,N_4995,N_4998);
and UO_479 (O_479,N_4975,N_4884);
nand UO_480 (O_480,N_4995,N_4802);
nor UO_481 (O_481,N_4864,N_4968);
nor UO_482 (O_482,N_4824,N_4846);
or UO_483 (O_483,N_4856,N_4815);
nand UO_484 (O_484,N_4873,N_4937);
nand UO_485 (O_485,N_4977,N_4878);
and UO_486 (O_486,N_4889,N_4960);
or UO_487 (O_487,N_4972,N_4872);
and UO_488 (O_488,N_4988,N_4894);
and UO_489 (O_489,N_4912,N_4891);
nand UO_490 (O_490,N_4864,N_4819);
or UO_491 (O_491,N_4957,N_4997);
or UO_492 (O_492,N_4879,N_4950);
xnor UO_493 (O_493,N_4817,N_4979);
or UO_494 (O_494,N_4804,N_4846);
or UO_495 (O_495,N_4816,N_4992);
or UO_496 (O_496,N_4966,N_4900);
or UO_497 (O_497,N_4876,N_4878);
nor UO_498 (O_498,N_4854,N_4921);
and UO_499 (O_499,N_4984,N_4806);
and UO_500 (O_500,N_4956,N_4849);
nor UO_501 (O_501,N_4876,N_4861);
nand UO_502 (O_502,N_4980,N_4820);
nand UO_503 (O_503,N_4853,N_4939);
nor UO_504 (O_504,N_4867,N_4856);
nor UO_505 (O_505,N_4857,N_4983);
and UO_506 (O_506,N_4997,N_4976);
nand UO_507 (O_507,N_4974,N_4849);
or UO_508 (O_508,N_4886,N_4912);
or UO_509 (O_509,N_4819,N_4884);
or UO_510 (O_510,N_4980,N_4891);
nor UO_511 (O_511,N_4997,N_4830);
xor UO_512 (O_512,N_4949,N_4858);
and UO_513 (O_513,N_4923,N_4878);
and UO_514 (O_514,N_4881,N_4901);
nor UO_515 (O_515,N_4929,N_4946);
or UO_516 (O_516,N_4946,N_4865);
nand UO_517 (O_517,N_4896,N_4914);
or UO_518 (O_518,N_4993,N_4906);
nand UO_519 (O_519,N_4804,N_4924);
and UO_520 (O_520,N_4987,N_4944);
nor UO_521 (O_521,N_4929,N_4926);
or UO_522 (O_522,N_4861,N_4891);
nand UO_523 (O_523,N_4823,N_4825);
or UO_524 (O_524,N_4889,N_4834);
nor UO_525 (O_525,N_4928,N_4820);
nor UO_526 (O_526,N_4929,N_4876);
nor UO_527 (O_527,N_4808,N_4950);
xor UO_528 (O_528,N_4943,N_4981);
nand UO_529 (O_529,N_4830,N_4902);
nor UO_530 (O_530,N_4958,N_4941);
nor UO_531 (O_531,N_4902,N_4849);
and UO_532 (O_532,N_4854,N_4880);
nand UO_533 (O_533,N_4932,N_4906);
nand UO_534 (O_534,N_4931,N_4904);
and UO_535 (O_535,N_4801,N_4806);
xor UO_536 (O_536,N_4943,N_4925);
nand UO_537 (O_537,N_4939,N_4981);
and UO_538 (O_538,N_4952,N_4855);
nand UO_539 (O_539,N_4867,N_4876);
nand UO_540 (O_540,N_4861,N_4880);
nor UO_541 (O_541,N_4937,N_4956);
or UO_542 (O_542,N_4816,N_4996);
and UO_543 (O_543,N_4837,N_4965);
or UO_544 (O_544,N_4813,N_4837);
or UO_545 (O_545,N_4939,N_4942);
nand UO_546 (O_546,N_4901,N_4970);
and UO_547 (O_547,N_4855,N_4939);
nand UO_548 (O_548,N_4880,N_4989);
and UO_549 (O_549,N_4876,N_4969);
and UO_550 (O_550,N_4973,N_4892);
xor UO_551 (O_551,N_4992,N_4866);
or UO_552 (O_552,N_4898,N_4940);
nand UO_553 (O_553,N_4806,N_4925);
or UO_554 (O_554,N_4901,N_4962);
nor UO_555 (O_555,N_4957,N_4996);
and UO_556 (O_556,N_4904,N_4949);
xor UO_557 (O_557,N_4918,N_4822);
nor UO_558 (O_558,N_4830,N_4913);
nand UO_559 (O_559,N_4925,N_4823);
nand UO_560 (O_560,N_4923,N_4851);
and UO_561 (O_561,N_4913,N_4833);
nand UO_562 (O_562,N_4980,N_4927);
and UO_563 (O_563,N_4847,N_4945);
nor UO_564 (O_564,N_4847,N_4978);
or UO_565 (O_565,N_4861,N_4900);
xnor UO_566 (O_566,N_4930,N_4823);
or UO_567 (O_567,N_4847,N_4853);
and UO_568 (O_568,N_4944,N_4840);
or UO_569 (O_569,N_4966,N_4918);
or UO_570 (O_570,N_4981,N_4944);
and UO_571 (O_571,N_4895,N_4962);
and UO_572 (O_572,N_4957,N_4927);
and UO_573 (O_573,N_4924,N_4913);
and UO_574 (O_574,N_4971,N_4813);
nand UO_575 (O_575,N_4900,N_4947);
or UO_576 (O_576,N_4902,N_4931);
nand UO_577 (O_577,N_4929,N_4849);
nor UO_578 (O_578,N_4930,N_4877);
nand UO_579 (O_579,N_4817,N_4959);
or UO_580 (O_580,N_4987,N_4825);
and UO_581 (O_581,N_4980,N_4839);
and UO_582 (O_582,N_4939,N_4991);
nand UO_583 (O_583,N_4956,N_4812);
nor UO_584 (O_584,N_4982,N_4826);
nand UO_585 (O_585,N_4952,N_4809);
nand UO_586 (O_586,N_4864,N_4997);
and UO_587 (O_587,N_4925,N_4942);
or UO_588 (O_588,N_4963,N_4855);
nor UO_589 (O_589,N_4958,N_4899);
nor UO_590 (O_590,N_4902,N_4979);
and UO_591 (O_591,N_4947,N_4943);
nand UO_592 (O_592,N_4979,N_4873);
nand UO_593 (O_593,N_4820,N_4978);
nand UO_594 (O_594,N_4996,N_4800);
nand UO_595 (O_595,N_4900,N_4972);
nand UO_596 (O_596,N_4904,N_4983);
nor UO_597 (O_597,N_4889,N_4959);
and UO_598 (O_598,N_4850,N_4855);
or UO_599 (O_599,N_4899,N_4824);
nor UO_600 (O_600,N_4865,N_4832);
nand UO_601 (O_601,N_4843,N_4911);
or UO_602 (O_602,N_4919,N_4972);
nor UO_603 (O_603,N_4895,N_4883);
nor UO_604 (O_604,N_4981,N_4874);
xor UO_605 (O_605,N_4819,N_4871);
or UO_606 (O_606,N_4864,N_4930);
nor UO_607 (O_607,N_4804,N_4916);
or UO_608 (O_608,N_4823,N_4944);
xor UO_609 (O_609,N_4810,N_4878);
and UO_610 (O_610,N_4850,N_4807);
nor UO_611 (O_611,N_4993,N_4917);
xor UO_612 (O_612,N_4903,N_4805);
and UO_613 (O_613,N_4929,N_4805);
and UO_614 (O_614,N_4921,N_4979);
nor UO_615 (O_615,N_4912,N_4941);
and UO_616 (O_616,N_4913,N_4881);
and UO_617 (O_617,N_4826,N_4906);
or UO_618 (O_618,N_4982,N_4916);
or UO_619 (O_619,N_4849,N_4867);
nand UO_620 (O_620,N_4831,N_4826);
nand UO_621 (O_621,N_4932,N_4826);
or UO_622 (O_622,N_4858,N_4977);
or UO_623 (O_623,N_4930,N_4910);
or UO_624 (O_624,N_4878,N_4976);
or UO_625 (O_625,N_4968,N_4905);
xor UO_626 (O_626,N_4862,N_4821);
nor UO_627 (O_627,N_4808,N_4983);
and UO_628 (O_628,N_4830,N_4841);
and UO_629 (O_629,N_4811,N_4897);
nor UO_630 (O_630,N_4905,N_4841);
and UO_631 (O_631,N_4935,N_4964);
xnor UO_632 (O_632,N_4946,N_4801);
nor UO_633 (O_633,N_4993,N_4837);
nand UO_634 (O_634,N_4864,N_4926);
and UO_635 (O_635,N_4823,N_4844);
nand UO_636 (O_636,N_4801,N_4857);
and UO_637 (O_637,N_4856,N_4946);
or UO_638 (O_638,N_4905,N_4876);
or UO_639 (O_639,N_4861,N_4976);
nor UO_640 (O_640,N_4921,N_4896);
or UO_641 (O_641,N_4983,N_4837);
nand UO_642 (O_642,N_4945,N_4801);
nor UO_643 (O_643,N_4955,N_4814);
nor UO_644 (O_644,N_4825,N_4862);
and UO_645 (O_645,N_4995,N_4968);
or UO_646 (O_646,N_4855,N_4909);
nor UO_647 (O_647,N_4985,N_4964);
and UO_648 (O_648,N_4808,N_4977);
nand UO_649 (O_649,N_4800,N_4855);
xor UO_650 (O_650,N_4850,N_4894);
and UO_651 (O_651,N_4953,N_4875);
nor UO_652 (O_652,N_4876,N_4823);
or UO_653 (O_653,N_4807,N_4996);
xor UO_654 (O_654,N_4842,N_4990);
and UO_655 (O_655,N_4847,N_4906);
xnor UO_656 (O_656,N_4887,N_4833);
or UO_657 (O_657,N_4917,N_4816);
nor UO_658 (O_658,N_4912,N_4803);
nand UO_659 (O_659,N_4866,N_4972);
and UO_660 (O_660,N_4963,N_4962);
xor UO_661 (O_661,N_4813,N_4952);
or UO_662 (O_662,N_4961,N_4899);
nand UO_663 (O_663,N_4818,N_4944);
nand UO_664 (O_664,N_4827,N_4808);
nand UO_665 (O_665,N_4975,N_4954);
nor UO_666 (O_666,N_4963,N_4878);
nor UO_667 (O_667,N_4985,N_4868);
nor UO_668 (O_668,N_4982,N_4957);
nand UO_669 (O_669,N_4995,N_4986);
or UO_670 (O_670,N_4893,N_4940);
nand UO_671 (O_671,N_4838,N_4966);
or UO_672 (O_672,N_4984,N_4993);
and UO_673 (O_673,N_4970,N_4809);
or UO_674 (O_674,N_4972,N_4886);
or UO_675 (O_675,N_4966,N_4983);
and UO_676 (O_676,N_4987,N_4916);
and UO_677 (O_677,N_4813,N_4874);
nand UO_678 (O_678,N_4999,N_4811);
nand UO_679 (O_679,N_4909,N_4918);
xor UO_680 (O_680,N_4856,N_4919);
nor UO_681 (O_681,N_4904,N_4814);
and UO_682 (O_682,N_4896,N_4972);
nand UO_683 (O_683,N_4880,N_4851);
nor UO_684 (O_684,N_4982,N_4867);
xnor UO_685 (O_685,N_4988,N_4901);
or UO_686 (O_686,N_4968,N_4981);
and UO_687 (O_687,N_4922,N_4818);
xor UO_688 (O_688,N_4820,N_4862);
and UO_689 (O_689,N_4932,N_4948);
and UO_690 (O_690,N_4871,N_4940);
nor UO_691 (O_691,N_4808,N_4926);
nor UO_692 (O_692,N_4968,N_4811);
or UO_693 (O_693,N_4801,N_4808);
nand UO_694 (O_694,N_4943,N_4828);
nand UO_695 (O_695,N_4850,N_4857);
and UO_696 (O_696,N_4990,N_4870);
nor UO_697 (O_697,N_4882,N_4917);
and UO_698 (O_698,N_4931,N_4882);
and UO_699 (O_699,N_4989,N_4907);
or UO_700 (O_700,N_4804,N_4879);
and UO_701 (O_701,N_4990,N_4848);
nand UO_702 (O_702,N_4846,N_4947);
nor UO_703 (O_703,N_4812,N_4838);
nor UO_704 (O_704,N_4887,N_4871);
nand UO_705 (O_705,N_4806,N_4940);
nand UO_706 (O_706,N_4908,N_4895);
or UO_707 (O_707,N_4805,N_4869);
nor UO_708 (O_708,N_4832,N_4883);
nand UO_709 (O_709,N_4826,N_4912);
and UO_710 (O_710,N_4886,N_4828);
and UO_711 (O_711,N_4814,N_4923);
or UO_712 (O_712,N_4864,N_4889);
or UO_713 (O_713,N_4807,N_4802);
or UO_714 (O_714,N_4981,N_4867);
nand UO_715 (O_715,N_4913,N_4969);
or UO_716 (O_716,N_4860,N_4907);
nand UO_717 (O_717,N_4826,N_4968);
or UO_718 (O_718,N_4908,N_4945);
or UO_719 (O_719,N_4983,N_4975);
or UO_720 (O_720,N_4983,N_4858);
or UO_721 (O_721,N_4857,N_4946);
xnor UO_722 (O_722,N_4823,N_4802);
nor UO_723 (O_723,N_4961,N_4816);
nand UO_724 (O_724,N_4852,N_4819);
and UO_725 (O_725,N_4914,N_4983);
and UO_726 (O_726,N_4857,N_4831);
nand UO_727 (O_727,N_4855,N_4820);
and UO_728 (O_728,N_4855,N_4808);
nand UO_729 (O_729,N_4947,N_4868);
or UO_730 (O_730,N_4939,N_4929);
and UO_731 (O_731,N_4964,N_4976);
nor UO_732 (O_732,N_4938,N_4892);
nand UO_733 (O_733,N_4871,N_4860);
nor UO_734 (O_734,N_4801,N_4956);
nand UO_735 (O_735,N_4817,N_4926);
nand UO_736 (O_736,N_4993,N_4954);
nor UO_737 (O_737,N_4851,N_4811);
nor UO_738 (O_738,N_4903,N_4869);
xor UO_739 (O_739,N_4991,N_4872);
and UO_740 (O_740,N_4944,N_4825);
nor UO_741 (O_741,N_4993,N_4912);
nor UO_742 (O_742,N_4805,N_4858);
or UO_743 (O_743,N_4849,N_4829);
nand UO_744 (O_744,N_4809,N_4935);
or UO_745 (O_745,N_4973,N_4894);
and UO_746 (O_746,N_4844,N_4947);
and UO_747 (O_747,N_4878,N_4900);
xnor UO_748 (O_748,N_4961,N_4957);
nor UO_749 (O_749,N_4945,N_4806);
nand UO_750 (O_750,N_4941,N_4951);
or UO_751 (O_751,N_4943,N_4882);
nor UO_752 (O_752,N_4822,N_4939);
or UO_753 (O_753,N_4911,N_4904);
and UO_754 (O_754,N_4842,N_4868);
nor UO_755 (O_755,N_4948,N_4869);
or UO_756 (O_756,N_4895,N_4901);
or UO_757 (O_757,N_4947,N_4836);
xnor UO_758 (O_758,N_4897,N_4805);
xor UO_759 (O_759,N_4913,N_4810);
nand UO_760 (O_760,N_4947,N_4961);
or UO_761 (O_761,N_4808,N_4844);
and UO_762 (O_762,N_4872,N_4960);
or UO_763 (O_763,N_4962,N_4841);
and UO_764 (O_764,N_4959,N_4870);
or UO_765 (O_765,N_4866,N_4978);
or UO_766 (O_766,N_4847,N_4823);
nand UO_767 (O_767,N_4804,N_4817);
nand UO_768 (O_768,N_4826,N_4858);
nand UO_769 (O_769,N_4924,N_4840);
nor UO_770 (O_770,N_4857,N_4933);
xor UO_771 (O_771,N_4823,N_4869);
and UO_772 (O_772,N_4987,N_4872);
nor UO_773 (O_773,N_4840,N_4918);
and UO_774 (O_774,N_4937,N_4989);
nand UO_775 (O_775,N_4903,N_4931);
or UO_776 (O_776,N_4971,N_4910);
nor UO_777 (O_777,N_4992,N_4964);
nand UO_778 (O_778,N_4949,N_4863);
and UO_779 (O_779,N_4937,N_4908);
xnor UO_780 (O_780,N_4917,N_4921);
nand UO_781 (O_781,N_4880,N_4958);
nand UO_782 (O_782,N_4917,N_4949);
and UO_783 (O_783,N_4817,N_4809);
nand UO_784 (O_784,N_4915,N_4958);
nor UO_785 (O_785,N_4999,N_4860);
or UO_786 (O_786,N_4816,N_4984);
or UO_787 (O_787,N_4854,N_4932);
nand UO_788 (O_788,N_4956,N_4933);
and UO_789 (O_789,N_4967,N_4876);
or UO_790 (O_790,N_4866,N_4867);
nand UO_791 (O_791,N_4800,N_4925);
nor UO_792 (O_792,N_4975,N_4899);
and UO_793 (O_793,N_4997,N_4828);
xor UO_794 (O_794,N_4945,N_4866);
and UO_795 (O_795,N_4984,N_4850);
and UO_796 (O_796,N_4988,N_4975);
xnor UO_797 (O_797,N_4817,N_4963);
and UO_798 (O_798,N_4922,N_4954);
or UO_799 (O_799,N_4984,N_4899);
xnor UO_800 (O_800,N_4813,N_4897);
nor UO_801 (O_801,N_4905,N_4906);
and UO_802 (O_802,N_4827,N_4857);
and UO_803 (O_803,N_4810,N_4840);
nand UO_804 (O_804,N_4887,N_4958);
nand UO_805 (O_805,N_4922,N_4911);
xor UO_806 (O_806,N_4964,N_4952);
or UO_807 (O_807,N_4910,N_4800);
and UO_808 (O_808,N_4955,N_4995);
xnor UO_809 (O_809,N_4927,N_4911);
or UO_810 (O_810,N_4889,N_4956);
or UO_811 (O_811,N_4831,N_4897);
nor UO_812 (O_812,N_4952,N_4897);
nand UO_813 (O_813,N_4942,N_4905);
nor UO_814 (O_814,N_4965,N_4893);
nor UO_815 (O_815,N_4975,N_4920);
nor UO_816 (O_816,N_4957,N_4847);
or UO_817 (O_817,N_4819,N_4921);
nor UO_818 (O_818,N_4973,N_4937);
and UO_819 (O_819,N_4951,N_4840);
nor UO_820 (O_820,N_4850,N_4958);
nor UO_821 (O_821,N_4824,N_4857);
xnor UO_822 (O_822,N_4970,N_4835);
nor UO_823 (O_823,N_4886,N_4965);
or UO_824 (O_824,N_4804,N_4823);
and UO_825 (O_825,N_4905,N_4997);
nor UO_826 (O_826,N_4903,N_4971);
nand UO_827 (O_827,N_4850,N_4881);
nand UO_828 (O_828,N_4869,N_4802);
or UO_829 (O_829,N_4805,N_4912);
nor UO_830 (O_830,N_4819,N_4898);
or UO_831 (O_831,N_4986,N_4904);
nand UO_832 (O_832,N_4843,N_4908);
nor UO_833 (O_833,N_4802,N_4874);
or UO_834 (O_834,N_4960,N_4979);
nand UO_835 (O_835,N_4809,N_4917);
nor UO_836 (O_836,N_4959,N_4975);
and UO_837 (O_837,N_4841,N_4983);
or UO_838 (O_838,N_4867,N_4889);
nor UO_839 (O_839,N_4982,N_4933);
xor UO_840 (O_840,N_4928,N_4957);
and UO_841 (O_841,N_4871,N_4834);
or UO_842 (O_842,N_4857,N_4852);
nand UO_843 (O_843,N_4945,N_4914);
nor UO_844 (O_844,N_4856,N_4835);
or UO_845 (O_845,N_4860,N_4810);
nor UO_846 (O_846,N_4813,N_4912);
nand UO_847 (O_847,N_4838,N_4950);
xnor UO_848 (O_848,N_4830,N_4994);
nand UO_849 (O_849,N_4906,N_4914);
nor UO_850 (O_850,N_4899,N_4823);
nor UO_851 (O_851,N_4956,N_4901);
or UO_852 (O_852,N_4870,N_4884);
and UO_853 (O_853,N_4929,N_4993);
and UO_854 (O_854,N_4949,N_4894);
and UO_855 (O_855,N_4802,N_4954);
or UO_856 (O_856,N_4949,N_4833);
nor UO_857 (O_857,N_4816,N_4838);
nor UO_858 (O_858,N_4842,N_4970);
nor UO_859 (O_859,N_4816,N_4948);
nand UO_860 (O_860,N_4902,N_4939);
or UO_861 (O_861,N_4820,N_4923);
or UO_862 (O_862,N_4846,N_4911);
nor UO_863 (O_863,N_4803,N_4957);
and UO_864 (O_864,N_4800,N_4998);
nor UO_865 (O_865,N_4943,N_4809);
or UO_866 (O_866,N_4831,N_4990);
nand UO_867 (O_867,N_4910,N_4932);
nor UO_868 (O_868,N_4996,N_4981);
nand UO_869 (O_869,N_4982,N_4938);
nand UO_870 (O_870,N_4983,N_4855);
xnor UO_871 (O_871,N_4999,N_4849);
nor UO_872 (O_872,N_4922,N_4988);
nand UO_873 (O_873,N_4871,N_4999);
nor UO_874 (O_874,N_4963,N_4800);
nand UO_875 (O_875,N_4833,N_4907);
or UO_876 (O_876,N_4945,N_4904);
or UO_877 (O_877,N_4995,N_4850);
nor UO_878 (O_878,N_4965,N_4918);
nand UO_879 (O_879,N_4946,N_4902);
or UO_880 (O_880,N_4808,N_4867);
and UO_881 (O_881,N_4842,N_4939);
nand UO_882 (O_882,N_4838,N_4971);
nor UO_883 (O_883,N_4964,N_4900);
nor UO_884 (O_884,N_4842,N_4800);
nor UO_885 (O_885,N_4863,N_4923);
or UO_886 (O_886,N_4878,N_4842);
nor UO_887 (O_887,N_4868,N_4967);
nor UO_888 (O_888,N_4950,N_4860);
nand UO_889 (O_889,N_4854,N_4980);
or UO_890 (O_890,N_4862,N_4899);
or UO_891 (O_891,N_4923,N_4995);
or UO_892 (O_892,N_4809,N_4959);
nand UO_893 (O_893,N_4985,N_4828);
and UO_894 (O_894,N_4890,N_4849);
and UO_895 (O_895,N_4809,N_4930);
nor UO_896 (O_896,N_4969,N_4907);
nand UO_897 (O_897,N_4883,N_4885);
nor UO_898 (O_898,N_4840,N_4954);
or UO_899 (O_899,N_4934,N_4851);
nand UO_900 (O_900,N_4844,N_4879);
or UO_901 (O_901,N_4821,N_4929);
and UO_902 (O_902,N_4887,N_4849);
nand UO_903 (O_903,N_4980,N_4947);
nor UO_904 (O_904,N_4980,N_4814);
or UO_905 (O_905,N_4832,N_4916);
nor UO_906 (O_906,N_4808,N_4985);
and UO_907 (O_907,N_4921,N_4890);
nand UO_908 (O_908,N_4999,N_4876);
and UO_909 (O_909,N_4964,N_4873);
or UO_910 (O_910,N_4847,N_4904);
nor UO_911 (O_911,N_4983,N_4873);
and UO_912 (O_912,N_4826,N_4974);
and UO_913 (O_913,N_4868,N_4924);
and UO_914 (O_914,N_4937,N_4959);
nor UO_915 (O_915,N_4905,N_4904);
or UO_916 (O_916,N_4920,N_4880);
and UO_917 (O_917,N_4896,N_4965);
or UO_918 (O_918,N_4972,N_4882);
nor UO_919 (O_919,N_4913,N_4908);
nor UO_920 (O_920,N_4993,N_4962);
nand UO_921 (O_921,N_4947,N_4890);
and UO_922 (O_922,N_4963,N_4854);
nand UO_923 (O_923,N_4938,N_4891);
nand UO_924 (O_924,N_4950,N_4997);
or UO_925 (O_925,N_4882,N_4951);
and UO_926 (O_926,N_4945,N_4819);
or UO_927 (O_927,N_4921,N_4878);
or UO_928 (O_928,N_4894,N_4999);
and UO_929 (O_929,N_4899,N_4804);
nand UO_930 (O_930,N_4847,N_4881);
or UO_931 (O_931,N_4801,N_4803);
xnor UO_932 (O_932,N_4904,N_4818);
or UO_933 (O_933,N_4971,N_4886);
nor UO_934 (O_934,N_4911,N_4960);
or UO_935 (O_935,N_4801,N_4877);
and UO_936 (O_936,N_4837,N_4880);
nor UO_937 (O_937,N_4854,N_4944);
nand UO_938 (O_938,N_4871,N_4863);
or UO_939 (O_939,N_4877,N_4904);
and UO_940 (O_940,N_4891,N_4966);
xnor UO_941 (O_941,N_4895,N_4970);
and UO_942 (O_942,N_4881,N_4980);
nor UO_943 (O_943,N_4885,N_4929);
xnor UO_944 (O_944,N_4825,N_4902);
or UO_945 (O_945,N_4986,N_4825);
nand UO_946 (O_946,N_4962,N_4925);
nand UO_947 (O_947,N_4903,N_4801);
nor UO_948 (O_948,N_4836,N_4985);
nand UO_949 (O_949,N_4933,N_4872);
and UO_950 (O_950,N_4982,N_4903);
and UO_951 (O_951,N_4986,N_4907);
nand UO_952 (O_952,N_4898,N_4889);
nand UO_953 (O_953,N_4801,N_4869);
xor UO_954 (O_954,N_4907,N_4827);
nand UO_955 (O_955,N_4990,N_4955);
nor UO_956 (O_956,N_4803,N_4845);
nor UO_957 (O_957,N_4866,N_4843);
and UO_958 (O_958,N_4848,N_4898);
nor UO_959 (O_959,N_4848,N_4831);
nand UO_960 (O_960,N_4933,N_4904);
nand UO_961 (O_961,N_4895,N_4889);
and UO_962 (O_962,N_4986,N_4862);
or UO_963 (O_963,N_4891,N_4963);
or UO_964 (O_964,N_4980,N_4817);
xor UO_965 (O_965,N_4912,N_4842);
xor UO_966 (O_966,N_4845,N_4933);
nand UO_967 (O_967,N_4903,N_4812);
and UO_968 (O_968,N_4929,N_4994);
xor UO_969 (O_969,N_4805,N_4935);
or UO_970 (O_970,N_4918,N_4856);
or UO_971 (O_971,N_4897,N_4933);
and UO_972 (O_972,N_4800,N_4867);
and UO_973 (O_973,N_4860,N_4822);
nor UO_974 (O_974,N_4898,N_4944);
xnor UO_975 (O_975,N_4992,N_4949);
or UO_976 (O_976,N_4887,N_4865);
or UO_977 (O_977,N_4922,N_4999);
xnor UO_978 (O_978,N_4832,N_4964);
or UO_979 (O_979,N_4928,N_4813);
and UO_980 (O_980,N_4897,N_4979);
xnor UO_981 (O_981,N_4892,N_4937);
or UO_982 (O_982,N_4873,N_4899);
or UO_983 (O_983,N_4849,N_4963);
nand UO_984 (O_984,N_4994,N_4868);
or UO_985 (O_985,N_4836,N_4875);
nor UO_986 (O_986,N_4812,N_4827);
nor UO_987 (O_987,N_4924,N_4940);
nor UO_988 (O_988,N_4857,N_4848);
nor UO_989 (O_989,N_4856,N_4896);
and UO_990 (O_990,N_4835,N_4984);
nand UO_991 (O_991,N_4836,N_4853);
nor UO_992 (O_992,N_4937,N_4916);
nand UO_993 (O_993,N_4938,N_4853);
and UO_994 (O_994,N_4943,N_4907);
and UO_995 (O_995,N_4837,N_4910);
or UO_996 (O_996,N_4832,N_4892);
and UO_997 (O_997,N_4908,N_4821);
nand UO_998 (O_998,N_4823,N_4909);
and UO_999 (O_999,N_4955,N_4967);
endmodule